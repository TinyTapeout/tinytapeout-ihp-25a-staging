module tt_um_znah_vga_ca (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire clknet_leaf_0_clk;
 wire \cell_x[0] ;
 wire \cell_x[1] ;
 wire \cell_x[2] ;
 wire \cell_x[3] ;
 wire \cell_x[4] ;
 wire \cell_x[5] ;
 wire \cell_x[6] ;
 wire \cell_x[7] ;
 wire \cellsbuf_[0].A ;
 wire \cellsbuf_[100].A ;
 wire \cellsbuf_[101].A ;
 wire \cellsbuf_[102].A ;
 wire \cellsbuf_[103].A ;
 wire \cellsbuf_[104].A ;
 wire \cellsbuf_[105].A ;
 wire \cellsbuf_[106].A ;
 wire \cellsbuf_[107].A ;
 wire \cellsbuf_[108].A ;
 wire \cellsbuf_[109].A ;
 wire \cellsbuf_[10].A ;
 wire \cellsbuf_[110].A ;
 wire \cellsbuf_[111].A ;
 wire \cellsbuf_[112].A ;
 wire \cellsbuf_[113].A ;
 wire \cellsbuf_[114].A ;
 wire \cellsbuf_[115].A ;
 wire \cellsbuf_[116].A ;
 wire \cellsbuf_[117].A ;
 wire \cellsbuf_[118].A ;
 wire \cellsbuf_[119].A ;
 wire \cellsbuf_[11].A ;
 wire \cellsbuf_[120].A ;
 wire \cellsbuf_[121].A ;
 wire \cellsbuf_[122].A ;
 wire \cellsbuf_[123].A ;
 wire \cellsbuf_[124].A ;
 wire \cellsbuf_[125].A ;
 wire \cellsbuf_[126].A ;
 wire \cellsbuf_[127].A ;
 wire \cellsbuf_[128].A ;
 wire \cellsbuf_[129].A ;
 wire \cellsbuf_[12].A ;
 wire \cellsbuf_[130].A ;
 wire \cellsbuf_[131].A ;
 wire \cellsbuf_[132].A ;
 wire \cellsbuf_[133].A ;
 wire \cellsbuf_[134].A ;
 wire \cellsbuf_[135].A ;
 wire \cellsbuf_[136].A ;
 wire \cellsbuf_[137].A ;
 wire \cellsbuf_[138].A ;
 wire \cellsbuf_[139].A ;
 wire \cellsbuf_[13].A ;
 wire \cellsbuf_[140].A ;
 wire \cellsbuf_[141].A ;
 wire \cellsbuf_[142].A ;
 wire \cellsbuf_[143].A ;
 wire \cellsbuf_[144].A ;
 wire \cellsbuf_[145].A ;
 wire \cellsbuf_[146].A ;
 wire \cellsbuf_[147].A ;
 wire \cellsbuf_[148].A ;
 wire \cellsbuf_[149].A ;
 wire \cellsbuf_[14].A ;
 wire \cellsbuf_[150].A ;
 wire \cellsbuf_[151].A ;
 wire \cellsbuf_[152].A ;
 wire \cellsbuf_[153].A ;
 wire \cellsbuf_[154].A ;
 wire \cellsbuf_[155].A ;
 wire \cellsbuf_[156].A ;
 wire \cellsbuf_[157].A ;
 wire \cellsbuf_[158].A ;
 wire \cellsbuf_[159].A ;
 wire \cellsbuf_[15].A ;
 wire \cellsbuf_[16].A ;
 wire \cellsbuf_[17].A ;
 wire \cellsbuf_[18].A ;
 wire \cellsbuf_[19].A ;
 wire \cellsbuf_[1].A ;
 wire \cellsbuf_[20].A ;
 wire \cellsbuf_[21].A ;
 wire \cellsbuf_[22].A ;
 wire \cellsbuf_[23].A ;
 wire \cellsbuf_[24].A ;
 wire \cellsbuf_[25].A ;
 wire \cellsbuf_[26].A ;
 wire \cellsbuf_[27].A ;
 wire \cellsbuf_[28].A ;
 wire \cellsbuf_[29].A ;
 wire \cellsbuf_[2].A ;
 wire \cellsbuf_[30].A ;
 wire \cellsbuf_[31].A ;
 wire \cellsbuf_[32].A ;
 wire \cellsbuf_[33].A ;
 wire \cellsbuf_[34].A ;
 wire \cellsbuf_[35].A ;
 wire \cellsbuf_[36].A ;
 wire \cellsbuf_[37].A ;
 wire \cellsbuf_[38].A ;
 wire \cellsbuf_[39].A ;
 wire \cellsbuf_[3].A ;
 wire \cellsbuf_[40].A ;
 wire \cellsbuf_[41].A ;
 wire \cellsbuf_[42].A ;
 wire \cellsbuf_[43].A ;
 wire \cellsbuf_[44].A ;
 wire \cellsbuf_[45].A ;
 wire \cellsbuf_[46].A ;
 wire \cellsbuf_[47].A ;
 wire \cellsbuf_[48].A ;
 wire \cellsbuf_[49].A ;
 wire \cellsbuf_[4].A ;
 wire \cellsbuf_[50].A ;
 wire \cellsbuf_[51].A ;
 wire \cellsbuf_[52].A ;
 wire \cellsbuf_[53].A ;
 wire \cellsbuf_[54].A ;
 wire \cellsbuf_[55].A ;
 wire \cellsbuf_[56].A ;
 wire \cellsbuf_[57].A ;
 wire \cellsbuf_[58].A ;
 wire \cellsbuf_[59].A ;
 wire \cellsbuf_[5].A ;
 wire \cellsbuf_[60].A ;
 wire \cellsbuf_[61].A ;
 wire \cellsbuf_[62].A ;
 wire \cellsbuf_[63].A ;
 wire \cellsbuf_[64].A ;
 wire \cellsbuf_[65].A ;
 wire \cellsbuf_[66].A ;
 wire \cellsbuf_[67].A ;
 wire \cellsbuf_[68].A ;
 wire \cellsbuf_[69].A ;
 wire \cellsbuf_[6].A ;
 wire \cellsbuf_[70].A ;
 wire \cellsbuf_[71].A ;
 wire \cellsbuf_[72].A ;
 wire \cellsbuf_[73].A ;
 wire \cellsbuf_[74].A ;
 wire \cellsbuf_[75].A ;
 wire \cellsbuf_[76].A ;
 wire \cellsbuf_[77].A ;
 wire \cellsbuf_[78].A ;
 wire \cellsbuf_[79].A ;
 wire \cellsbuf_[7].A ;
 wire \cellsbuf_[80].A ;
 wire \cellsbuf_[81].A ;
 wire \cellsbuf_[82].A ;
 wire \cellsbuf_[83].A ;
 wire \cellsbuf_[84].A ;
 wire \cellsbuf_[85].A ;
 wire \cellsbuf_[86].A ;
 wire \cellsbuf_[87].A ;
 wire \cellsbuf_[88].A ;
 wire \cellsbuf_[89].A ;
 wire \cellsbuf_[8].A ;
 wire \cellsbuf_[90].A ;
 wire \cellsbuf_[91].A ;
 wire \cellsbuf_[92].A ;
 wire \cellsbuf_[93].A ;
 wire \cellsbuf_[94].A ;
 wire \cellsbuf_[95].A ;
 wire \cellsbuf_[96].A ;
 wire \cellsbuf_[97].A ;
 wire \cellsbuf_[98].A ;
 wire \cellsbuf_[99].A ;
 wire \cellsbuf_[9].A ;
 wire \fract_x[0] ;
 wire \fract_x[1] ;
 wire \fract_y[0] ;
 wire \fract_y[1] ;
 wire hsync;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \i[0] ;
 wire \i[1] ;
 wire \i[2] ;
 wire left;
 wire \next_cellsbuf_[0].A ;
 wire \next_cellsbuf_[100].A ;
 wire \next_cellsbuf_[101].A ;
 wire \next_cellsbuf_[102].A ;
 wire \next_cellsbuf_[103].A ;
 wire \next_cellsbuf_[104].A ;
 wire \next_cellsbuf_[105].A ;
 wire \next_cellsbuf_[106].A ;
 wire \next_cellsbuf_[107].A ;
 wire \next_cellsbuf_[108].A ;
 wire \next_cellsbuf_[109].A ;
 wire \next_cellsbuf_[10].A ;
 wire \next_cellsbuf_[110].A ;
 wire \next_cellsbuf_[111].A ;
 wire \next_cellsbuf_[112].A ;
 wire \next_cellsbuf_[113].A ;
 wire \next_cellsbuf_[114].A ;
 wire \next_cellsbuf_[115].A ;
 wire \next_cellsbuf_[116].A ;
 wire \next_cellsbuf_[117].A ;
 wire \next_cellsbuf_[118].A ;
 wire \next_cellsbuf_[119].A ;
 wire \next_cellsbuf_[11].A ;
 wire \next_cellsbuf_[120].A ;
 wire \next_cellsbuf_[121].A ;
 wire \next_cellsbuf_[122].A ;
 wire \next_cellsbuf_[123].A ;
 wire \next_cellsbuf_[124].A ;
 wire \next_cellsbuf_[125].A ;
 wire \next_cellsbuf_[126].A ;
 wire \next_cellsbuf_[127].A ;
 wire \next_cellsbuf_[128].A ;
 wire \next_cellsbuf_[129].A ;
 wire \next_cellsbuf_[12].A ;
 wire \next_cellsbuf_[130].A ;
 wire \next_cellsbuf_[131].A ;
 wire \next_cellsbuf_[132].A ;
 wire \next_cellsbuf_[133].A ;
 wire \next_cellsbuf_[134].A ;
 wire \next_cellsbuf_[135].A ;
 wire \next_cellsbuf_[136].A ;
 wire \next_cellsbuf_[137].A ;
 wire \next_cellsbuf_[138].A ;
 wire \next_cellsbuf_[139].A ;
 wire \next_cellsbuf_[13].A ;
 wire \next_cellsbuf_[140].A ;
 wire \next_cellsbuf_[141].A ;
 wire \next_cellsbuf_[142].A ;
 wire \next_cellsbuf_[143].A ;
 wire \next_cellsbuf_[144].A ;
 wire \next_cellsbuf_[145].A ;
 wire \next_cellsbuf_[146].A ;
 wire \next_cellsbuf_[147].A ;
 wire \next_cellsbuf_[148].A ;
 wire \next_cellsbuf_[149].A ;
 wire \next_cellsbuf_[14].A ;
 wire \next_cellsbuf_[150].A ;
 wire \next_cellsbuf_[151].A ;
 wire \next_cellsbuf_[152].A ;
 wire \next_cellsbuf_[153].A ;
 wire \next_cellsbuf_[154].A ;
 wire \next_cellsbuf_[155].A ;
 wire \next_cellsbuf_[156].A ;
 wire \next_cellsbuf_[157].A ;
 wire \next_cellsbuf_[158].A ;
 wire \next_cellsbuf_[159].A ;
 wire \next_cellsbuf_[15].A ;
 wire \next_cellsbuf_[16].A ;
 wire \next_cellsbuf_[17].A ;
 wire \next_cellsbuf_[18].A ;
 wire \next_cellsbuf_[19].A ;
 wire \next_cellsbuf_[1].A ;
 wire \next_cellsbuf_[20].A ;
 wire \next_cellsbuf_[21].A ;
 wire \next_cellsbuf_[22].A ;
 wire \next_cellsbuf_[23].A ;
 wire \next_cellsbuf_[24].A ;
 wire \next_cellsbuf_[25].A ;
 wire \next_cellsbuf_[26].A ;
 wire \next_cellsbuf_[27].A ;
 wire \next_cellsbuf_[28].A ;
 wire \next_cellsbuf_[29].A ;
 wire \next_cellsbuf_[2].A ;
 wire \next_cellsbuf_[30].A ;
 wire \next_cellsbuf_[31].A ;
 wire \next_cellsbuf_[32].A ;
 wire \next_cellsbuf_[33].A ;
 wire \next_cellsbuf_[34].A ;
 wire \next_cellsbuf_[35].A ;
 wire \next_cellsbuf_[36].A ;
 wire \next_cellsbuf_[37].A ;
 wire \next_cellsbuf_[38].A ;
 wire \next_cellsbuf_[39].A ;
 wire \next_cellsbuf_[3].A ;
 wire \next_cellsbuf_[40].A ;
 wire \next_cellsbuf_[41].A ;
 wire \next_cellsbuf_[42].A ;
 wire \next_cellsbuf_[43].A ;
 wire \next_cellsbuf_[44].A ;
 wire \next_cellsbuf_[45].A ;
 wire \next_cellsbuf_[46].A ;
 wire \next_cellsbuf_[47].A ;
 wire \next_cellsbuf_[48].A ;
 wire \next_cellsbuf_[49].A ;
 wire \next_cellsbuf_[4].A ;
 wire \next_cellsbuf_[50].A ;
 wire \next_cellsbuf_[51].A ;
 wire \next_cellsbuf_[52].A ;
 wire \next_cellsbuf_[53].A ;
 wire \next_cellsbuf_[54].A ;
 wire \next_cellsbuf_[55].A ;
 wire \next_cellsbuf_[56].A ;
 wire \next_cellsbuf_[57].A ;
 wire \next_cellsbuf_[58].A ;
 wire \next_cellsbuf_[59].A ;
 wire \next_cellsbuf_[5].A ;
 wire \next_cellsbuf_[60].A ;
 wire \next_cellsbuf_[61].A ;
 wire \next_cellsbuf_[62].A ;
 wire \next_cellsbuf_[63].A ;
 wire \next_cellsbuf_[64].A ;
 wire \next_cellsbuf_[65].A ;
 wire \next_cellsbuf_[66].A ;
 wire \next_cellsbuf_[67].A ;
 wire \next_cellsbuf_[68].A ;
 wire \next_cellsbuf_[69].A ;
 wire \next_cellsbuf_[6].A ;
 wire \next_cellsbuf_[70].A ;
 wire \next_cellsbuf_[71].A ;
 wire \next_cellsbuf_[72].A ;
 wire \next_cellsbuf_[73].A ;
 wire \next_cellsbuf_[74].A ;
 wire \next_cellsbuf_[75].A ;
 wire \next_cellsbuf_[76].A ;
 wire \next_cellsbuf_[77].A ;
 wire \next_cellsbuf_[78].A ;
 wire \next_cellsbuf_[79].A ;
 wire \next_cellsbuf_[7].A ;
 wire \next_cellsbuf_[80].A ;
 wire \next_cellsbuf_[81].A ;
 wire \next_cellsbuf_[82].A ;
 wire \next_cellsbuf_[83].A ;
 wire \next_cellsbuf_[84].A ;
 wire \next_cellsbuf_[85].A ;
 wire \next_cellsbuf_[86].A ;
 wire \next_cellsbuf_[87].A ;
 wire \next_cellsbuf_[88].A ;
 wire \next_cellsbuf_[89].A ;
 wire \next_cellsbuf_[8].A ;
 wire \next_cellsbuf_[90].A ;
 wire \next_cellsbuf_[91].A ;
 wire \next_cellsbuf_[92].A ;
 wire \next_cellsbuf_[93].A ;
 wire \next_cellsbuf_[94].A ;
 wire \next_cellsbuf_[95].A ;
 wire \next_cellsbuf_[96].A ;
 wire \next_cellsbuf_[97].A ;
 wire \next_cellsbuf_[98].A ;
 wire \next_cellsbuf_[99].A ;
 wire \next_cellsbuf_[9].A ;
 wire \row_count[0] ;
 wire \row_count[1] ;
 wire \row_count[2] ;
 wire \row_count[3] ;
 wire \row_count[4] ;
 wire \row_count[5] ;
 wire \row_count[6] ;
 wire \row_count[7] ;
 wire \rule[0] ;
 wire \rule[1] ;
 wire \rule[2] ;
 wire \rule[3] ;
 wire \rule[4] ;
 wire \rule[5] ;
 wire \rule[6] ;
 wire \rule[7] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net1;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;

 sg13g2_inv_1 _1248_ (.Y(_0434_),
    .A(net917));
 sg13g2_inv_1 _1249_ (.Y(_0435_),
    .A(\i[0] ));
 sg13g2_inv_1 _1250_ (.Y(_0436_),
    .A(net963));
 sg13g2_inv_1 _1251_ (.Y(_0437_),
    .A(net441));
 sg13g2_inv_1 _1252_ (.Y(_0438_),
    .A(\fract_y[0] ));
 sg13g2_inv_1 _1253_ (.Y(_0439_),
    .A(_0010_));
 sg13g2_inv_1 _1254_ (.Y(_0440_),
    .A(_0012_));
 sg13g2_inv_1 _1255_ (.Y(_0441_),
    .A(net252));
 sg13g2_inv_1 _1256_ (.Y(_0442_),
    .A(net440));
 sg13g2_nand4_1 _1257_ (.B(\hvsync_gen.vpos[7] ),
    .C(\hvsync_gen.vpos[6] ),
    .A(\hvsync_gen.vpos[8] ),
    .Y(_0443_),
    .D(\hvsync_gen.vpos[5] ));
 sg13g2_nor4_2 _1258_ (.A(\hvsync_gen.vpos[9] ),
    .B(\hvsync_gen.vpos[4] ),
    .C(\hvsync_gen.vpos[2] ),
    .Y(_0444_),
    .D(_0443_));
 sg13g2_and3_1 _1259_ (.X(_0008_),
    .A(\hvsync_gen.vpos[3] ),
    .B(net845),
    .C(_0444_));
 sg13g2_nor3_1 _1260_ (.A(net962),
    .B(net938),
    .C(net955),
    .Y(_0445_));
 sg13g2_and3_1 _1261_ (.X(_0446_),
    .A(net962),
    .B(net938),
    .C(net955));
 sg13g2_nand3b_1 _1262_ (.B(net957),
    .C(net959),
    .Y(_0447_),
    .A_N(net913));
 sg13g2_nor3_1 _1263_ (.A(_0445_),
    .B(_0446_),
    .C(_0447_),
    .Y(_0007_));
 sg13g2_nor2b_2 _1264_ (.A(\hvsync_gen.vpos[9] ),
    .B_N(_0443_),
    .Y(_0448_));
 sg13g2_o21ai_1 _1265_ (.B1(\cell_x[7] ),
    .Y(_0449_),
    .A1(\cell_x[5] ),
    .A2(\cell_x[6] ));
 sg13g2_and3_2 _1266_ (.X(_0450_),
    .A(\cellsbuf_[0].A ),
    .B(_0448_),
    .C(_0449_));
 sg13g2_and2_1 _1267_ (.A(\rule[1] ),
    .B(_0450_),
    .X(uo_out[6]));
 sg13g2_and2_1 _1268_ (.A(\rule[2] ),
    .B(_0450_),
    .X(uo_out[2]));
 sg13g2_and2_1 _1269_ (.A(\rule[3] ),
    .B(_0450_),
    .X(uo_out[5]));
 sg13g2_and2_1 _1270_ (.A(\rule[4] ),
    .B(_0450_),
    .X(uo_out[1]));
 sg13g2_and2_1 _1271_ (.A(\rule[5] ),
    .B(_0450_),
    .X(uo_out[4]));
 sg13g2_and2_1 _1272_ (.A(\rule[6] ),
    .B(_0450_),
    .X(uo_out[0]));
 sg13g2_or4_1 _1273_ (.A(\cell_x[2] ),
    .B(\cell_x[3] ),
    .C(\cell_x[1] ),
    .D(\cell_x[0] ),
    .X(_0451_));
 sg13g2_nor2_1 _1274_ (.A(\fract_x[0] ),
    .B(net969),
    .Y(_0452_));
 sg13g2_or2_1 _1275_ (.X(_0453_),
    .B(\fract_x[1] ),
    .A(\fract_x[0] ));
 sg13g2_nor4_2 _1276_ (.A(\cell_x[4] ),
    .B(_0447_),
    .C(_0451_),
    .Y(_0454_),
    .D(_0453_));
 sg13g2_and2_2 _1277_ (.A(\fract_y[1] ),
    .B(\fract_y[0] ),
    .X(_0455_));
 sg13g2_and3_1 _1278_ (.X(_0456_),
    .A(_0448_),
    .B(_0454_),
    .C(_0455_));
 sg13g2_nand3_1 _1279_ (.B(_0454_),
    .C(_0455_),
    .A(_0448_),
    .Y(_0457_));
 sg13g2_nor2_2 _1280_ (.A(\fract_y[1] ),
    .B(\fract_y[0] ),
    .Y(_0458_));
 sg13g2_nor3_1 _1281_ (.A(\hvsync_gen.vpos[3] ),
    .B(\fract_y[1] ),
    .C(\fract_y[0] ),
    .Y(_0459_));
 sg13g2_nand2b_1 _1282_ (.Y(_0460_),
    .B(_0458_),
    .A_N(\hvsync_gen.vpos[3] ));
 sg13g2_nand3_1 _1283_ (.B(_0454_),
    .C(_0459_),
    .A(_0444_),
    .Y(_0461_));
 sg13g2_nand2_2 _1284_ (.Y(_0462_),
    .A(_0457_),
    .B(_0461_));
 sg13g2_nand3_1 _1285_ (.B(_0454_),
    .C(_0455_),
    .A(_0448_),
    .Y(_0463_));
 sg13g2_nand3_1 _1286_ (.B(_0454_),
    .C(_0459_),
    .A(_0444_),
    .Y(_0464_));
 sg13g2_nand2_2 _1287_ (.Y(_0465_),
    .A(_0463_),
    .B(_0464_));
 sg13g2_and3_1 _1288_ (.X(_0466_),
    .A(net931),
    .B(net935),
    .C(\row_count[0] ));
 sg13g2_nand3_1 _1289_ (.B(\row_count[1] ),
    .C(\row_count[0] ),
    .A(\row_count[2] ),
    .Y(_0467_));
 sg13g2_o21ai_1 _1290_ (.B1(_0011_),
    .Y(_0468_),
    .A1(\row_count[3] ),
    .A2(_0467_));
 sg13g2_and3_1 _1291_ (.X(_0469_),
    .A(\row_count[6] ),
    .B(\row_count[5] ),
    .C(\row_count[4] ));
 sg13g2_nand3_1 _1292_ (.B(net929),
    .C(\row_count[4] ),
    .A(net924),
    .Y(_0470_));
 sg13g2_nor2_1 _1293_ (.A(\row_count[7] ),
    .B(_0470_),
    .Y(_0471_));
 sg13g2_a21oi_2 _1294_ (.B1(_0439_),
    .Y(_0472_),
    .A2(_0471_),
    .A1(_0468_));
 sg13g2_a21oi_2 _1295_ (.B1(_0456_),
    .Y(_0473_),
    .A2(_0472_),
    .A1(_0435_));
 sg13g2_nand2_1 _1296_ (.Y(_0474_),
    .A(\row_count[3] ),
    .B(_0466_));
 sg13g2_and4_2 _1297_ (.A(\row_count[7] ),
    .B(\row_count[3] ),
    .C(_0466_),
    .D(_0469_),
    .X(_0475_));
 sg13g2_a21oi_1 _1298_ (.A1(_0440_),
    .A2(_0475_),
    .Y(_0476_),
    .B1(_0457_));
 sg13g2_or3_1 _1299_ (.A(_0009_),
    .B(_0473_),
    .C(_0476_),
    .X(_0477_));
 sg13g2_o21ai_1 _1300_ (.B1(_0009_),
    .Y(_0478_),
    .A1(_0473_),
    .A2(_0476_));
 sg13g2_nand3_1 _1301_ (.B(_0477_),
    .C(_0478_),
    .A(_0465_),
    .Y(_0479_));
 sg13g2_o21ai_1 _1302_ (.B1(_0479_),
    .Y(_0480_),
    .A1(_0009_),
    .A2(_0462_));
 sg13g2_nor2_1 _1303_ (.A(_0013_),
    .B(_0462_),
    .Y(_0481_));
 sg13g2_nand3_1 _1304_ (.B(\i[0] ),
    .C(_0475_),
    .A(\i[1] ),
    .Y(_0482_));
 sg13g2_mux2_1 _1305_ (.A0(_0482_),
    .A1(\i[1] ),
    .S(_0463_),
    .X(_0483_));
 sg13g2_o21ai_1 _1306_ (.B1(_0013_),
    .Y(_0484_),
    .A1(_0473_),
    .A2(_0483_));
 sg13g2_or3_1 _1307_ (.A(_0013_),
    .B(_0473_),
    .C(_0483_),
    .X(_0485_));
 sg13g2_nand3_1 _1308_ (.B(_0484_),
    .C(_0485_),
    .A(_0465_),
    .Y(_0486_));
 sg13g2_nor2b_2 _1309_ (.A(_0481_),
    .B_N(_0486_),
    .Y(_0487_));
 sg13g2_nand2b_2 _1310_ (.Y(_0488_),
    .B(_0486_),
    .A_N(_0481_));
 sg13g2_nand2_1 _1311_ (.Y(_0489_),
    .A(net253),
    .B(_0488_));
 sg13g2_nor2_1 _1312_ (.A(_0012_),
    .B(_0462_),
    .Y(_0490_));
 sg13g2_nor2_1 _1313_ (.A(_0463_),
    .B(_0475_),
    .Y(_0491_));
 sg13g2_mux2_1 _1314_ (.A0(_0472_),
    .A1(_0475_),
    .S(_0456_),
    .X(_0492_));
 sg13g2_nand2b_1 _1315_ (.Y(_0493_),
    .B(_0012_),
    .A_N(_0492_));
 sg13g2_nand2_1 _1316_ (.Y(_0494_),
    .A(_0440_),
    .B(_0492_));
 sg13g2_nand3_1 _1317_ (.B(_0493_),
    .C(_0494_),
    .A(_0465_),
    .Y(_0495_));
 sg13g2_nor2b_2 _1318_ (.A(_0490_),
    .B_N(_0495_),
    .Y(_0496_));
 sg13g2_nand2b_1 _1319_ (.Y(_0497_),
    .B(_0495_),
    .A_N(_0490_));
 sg13g2_nor3_1 _1320_ (.A(net251),
    .B(_0487_),
    .C(_0496_),
    .Y(_0498_));
 sg13g2_nand3_1 _1321_ (.B(_0488_),
    .C(_0497_),
    .A(net253),
    .Y(_0499_));
 sg13g2_a21oi_2 _1322_ (.B1(net251),
    .Y(_0500_),
    .A2(_0496_),
    .A1(_0487_));
 sg13g2_o21ai_1 _1323_ (.B1(net252),
    .Y(_0501_),
    .A1(_0488_),
    .A2(_0497_));
 sg13g2_and3_1 _1324_ (.X(_0000_),
    .A(_0480_),
    .B(_0499_),
    .C(_0500_));
 sg13g2_nand3_1 _1325_ (.B(_0499_),
    .C(_0500_),
    .A(_0480_),
    .Y(_0001_));
 sg13g2_nand3_1 _1326_ (.B(_0480_),
    .C(_0497_),
    .A(net252),
    .Y(_0502_));
 sg13g2_mux2_1 _1327_ (.A0(_0488_),
    .A1(_0489_),
    .S(_0502_),
    .X(_0002_));
 sg13g2_nand4_1 _1328_ (.B(_0480_),
    .C(_0487_),
    .A(net252),
    .Y(_0503_),
    .D(_0496_));
 sg13g2_and2_1 _1329_ (.A(_0499_),
    .B(_0503_),
    .X(_0003_));
 sg13g2_nand2b_1 _1330_ (.Y(_0504_),
    .B(_0488_),
    .A_N(_0480_));
 sg13g2_nand2_1 _1331_ (.Y(_0004_),
    .A(_0500_),
    .B(_0504_));
 sg13g2_nand2_1 _1332_ (.Y(_0505_),
    .A(_0480_),
    .B(_0487_));
 sg13g2_and3_1 _1333_ (.X(_0005_),
    .A(_0500_),
    .B(_0504_),
    .C(_0505_));
 sg13g2_o21ai_1 _1334_ (.B1(_0502_),
    .Y(_0006_),
    .A1(_0498_),
    .A2(_0501_));
 sg13g2_nor2_1 _1335_ (.A(_0480_),
    .B(_0499_),
    .Y(_0018_));
 sg13g2_and4_2 _1336_ (.A(net252),
    .B(_0448_),
    .C(_0449_),
    .D(_0452_),
    .X(_0506_));
 sg13g2_nand4_1 _1337_ (.B(_0448_),
    .C(_0449_),
    .A(net252),
    .Y(_0507_),
    .D(_0452_));
 sg13g2_mux2_1 _1338_ (.A0(net943),
    .A1(left),
    .S(net250),
    .X(_0019_));
 sg13g2_nor2b_1 _1339_ (.A(\cellsbuf_[158].A ),
    .B_N(\rule[4] ),
    .Y(_0508_));
 sg13g2_a21oi_1 _1340_ (.A1(\cellsbuf_[158].A ),
    .A2(\rule[5] ),
    .Y(_0509_),
    .B1(_0508_));
 sg13g2_mux2_1 _1341_ (.A0(\rule[0] ),
    .A1(\rule[1] ),
    .S(\cellsbuf_[158].A ),
    .X(_0510_));
 sg13g2_o21ai_1 _1342_ (.B1(_0458_),
    .Y(_0511_),
    .A1(left),
    .A2(_0510_));
 sg13g2_a21oi_1 _1343_ (.A1(left),
    .A2(_0509_),
    .Y(_0512_),
    .B1(_0511_));
 sg13g2_nor2_1 _1344_ (.A(\hvsync_gen.vpos[8] ),
    .B(\hvsync_gen.vpos[7] ),
    .Y(_0513_));
 sg13g2_nor3_1 _1345_ (.A(\hvsync_gen.vpos[6] ),
    .B(\hvsync_gen.vpos[5] ),
    .C(\hvsync_gen.vpos[4] ),
    .Y(_0514_));
 sg13g2_nand2_1 _1346_ (.Y(_0515_),
    .A(_0513_),
    .B(_0514_));
 sg13g2_nor4_2 _1347_ (.A(\hvsync_gen.vpos[9] ),
    .B(\hvsync_gen.vpos[2] ),
    .C(_0460_),
    .Y(_0516_),
    .D(_0515_));
 sg13g2_mux4_1 _1348_ (.S0(\cellsbuf_[158].A ),
    .A0(\rule[2] ),
    .A1(\rule[3] ),
    .A2(\rule[6] ),
    .A3(\rule[7] ),
    .S1(left),
    .X(_0517_));
 sg13g2_nand3b_1 _1349_ (.B(_0458_),
    .C(\cellsbuf_[159].A ),
    .Y(_0518_),
    .A_N(_0517_));
 sg13g2_o21ai_1 _1350_ (.B1(_0518_),
    .Y(_0519_),
    .A1(\cellsbuf_[159].A ),
    .A2(_0512_));
 sg13g2_nor3_1 _1351_ (.A(\row_count[2] ),
    .B(\row_count[1] ),
    .C(\row_count[0] ),
    .Y(_0520_));
 sg13g2_nor4_1 _1352_ (.A(\row_count[6] ),
    .B(\row_count[5] ),
    .C(\row_count[4] ),
    .D(\row_count[3] ),
    .Y(_0521_));
 sg13g2_nor4_1 _1353_ (.A(\i[2] ),
    .B(\i[1] ),
    .C(\i[0] ),
    .D(\row_count[7] ),
    .Y(_0522_));
 sg13g2_nand3_1 _1354_ (.B(_0521_),
    .C(_0522_),
    .A(_0520_),
    .Y(_0523_));
 sg13g2_nor2b_1 _1355_ (.A(\cell_x[5] ),
    .B_N(\cell_x[6] ),
    .Y(_0524_));
 sg13g2_nand2_1 _1356_ (.Y(_0525_),
    .A(\cell_x[4] ),
    .B(_0524_));
 sg13g2_nor3_1 _1357_ (.A(\cell_x[7] ),
    .B(_0451_),
    .C(_0525_),
    .Y(_0526_));
 sg13g2_mux2_1 _1358_ (.A0(_0526_),
    .A1(\next_cellsbuf_[159].A ),
    .S(_0523_),
    .X(_0527_));
 sg13g2_nand2_1 _1359_ (.Y(_0528_),
    .A(_0516_),
    .B(_0527_));
 sg13g2_o21ai_1 _1360_ (.B1(_0528_),
    .Y(_0529_),
    .A1(_0516_),
    .A2(_0519_));
 sg13g2_nand2_1 _1361_ (.Y(_0530_),
    .A(_0506_),
    .B(_0529_));
 sg13g2_nand2_1 _1362_ (.Y(_0531_),
    .A(net254),
    .B(net876));
 sg13g2_o21ai_1 _1363_ (.B1(_0530_),
    .Y(_0020_),
    .A1(_0506_),
    .A2(_0531_));
 sg13g2_nor4_1 _1364_ (.A(\hvsync_gen.vpos[9] ),
    .B(_0460_),
    .C(net245),
    .D(_0515_),
    .Y(_0532_));
 sg13g2_mux2_1 _1365_ (.A0(net601),
    .A1(net798),
    .S(net218),
    .X(_0021_));
 sg13g2_mux2_1 _1366_ (.A0(\next_cellsbuf_[2].A ),
    .A1(net601),
    .S(net218),
    .X(_0022_));
 sg13g2_mux2_1 _1367_ (.A0(net618),
    .A1(\next_cellsbuf_[2].A ),
    .S(net218),
    .X(_0023_));
 sg13g2_mux2_1 _1368_ (.A0(net636),
    .A1(net618),
    .S(net218),
    .X(_0024_));
 sg13g2_mux2_1 _1369_ (.A0(net634),
    .A1(\next_cellsbuf_[4].A ),
    .S(net218),
    .X(_0025_));
 sg13g2_mux2_1 _1370_ (.A0(net525),
    .A1(net634),
    .S(net218),
    .X(_0026_));
 sg13g2_mux2_1 _1371_ (.A0(\next_cellsbuf_[7].A ),
    .A1(net525),
    .S(net216),
    .X(_0027_));
 sg13g2_mux2_1 _1372_ (.A0(net788),
    .A1(\next_cellsbuf_[7].A ),
    .S(net216),
    .X(_0028_));
 sg13g2_mux2_1 _1373_ (.A0(net891),
    .A1(net788),
    .S(net216),
    .X(_0029_));
 sg13g2_mux2_1 _1374_ (.A0(net774),
    .A1(\next_cellsbuf_[9].A ),
    .S(net216),
    .X(_0030_));
 sg13g2_mux2_1 _1375_ (.A0(net603),
    .A1(\next_cellsbuf_[10].A ),
    .S(net217),
    .X(_0031_));
 sg13g2_mux2_1 _1376_ (.A0(net805),
    .A1(net603),
    .S(net214),
    .X(_0032_));
 sg13g2_mux2_1 _1377_ (.A0(net810),
    .A1(net805),
    .S(net214),
    .X(_0033_));
 sg13g2_mux2_1 _1378_ (.A0(net887),
    .A1(net810),
    .S(net214),
    .X(_0034_));
 sg13g2_mux2_1 _1379_ (.A0(net885),
    .A1(\next_cellsbuf_[14].A ),
    .S(net219),
    .X(_0035_));
 sg13g2_mux2_1 _1380_ (.A0(net854),
    .A1(\next_cellsbuf_[15].A ),
    .S(net213),
    .X(_0036_));
 sg13g2_mux2_1 _1381_ (.A0(net915),
    .A1(net854),
    .S(net213),
    .X(_0037_));
 sg13g2_mux2_1 _1382_ (.A0(net720),
    .A1(\next_cellsbuf_[17].A ),
    .S(net212),
    .X(_0038_));
 sg13g2_mux2_1 _1383_ (.A0(net614),
    .A1(\next_cellsbuf_[18].A ),
    .S(net211),
    .X(_0039_));
 sg13g2_mux2_1 _1384_ (.A0(net508),
    .A1(\next_cellsbuf_[19].A ),
    .S(net211),
    .X(_0040_));
 sg13g2_mux2_1 _1385_ (.A0(net840),
    .A1(net508),
    .S(net211),
    .X(_0041_));
 sg13g2_mux2_1 _1386_ (.A0(net704),
    .A1(\next_cellsbuf_[21].A ),
    .S(net211),
    .X(_0042_));
 sg13g2_mux2_1 _1387_ (.A0(net764),
    .A1(net704),
    .S(net211),
    .X(_0043_));
 sg13g2_mux2_1 _1388_ (.A0(net487),
    .A1(\next_cellsbuf_[23].A ),
    .S(net211),
    .X(_0044_));
 sg13g2_mux2_1 _1389_ (.A0(net637),
    .A1(net487),
    .S(net212),
    .X(_0045_));
 sg13g2_mux2_1 _1390_ (.A0(net856),
    .A1(net637),
    .S(net211),
    .X(_0046_));
 sg13g2_mux2_1 _1391_ (.A0(net591),
    .A1(\next_cellsbuf_[26].A ),
    .S(net211),
    .X(_0047_));
 sg13g2_mux2_1 _1392_ (.A0(net666),
    .A1(net591),
    .S(net205),
    .X(_0048_));
 sg13g2_mux2_1 _1393_ (.A0(net595),
    .A1(\next_cellsbuf_[28].A ),
    .S(net204),
    .X(_0049_));
 sg13g2_mux2_1 _1394_ (.A0(net761),
    .A1(net595),
    .S(net205),
    .X(_0050_));
 sg13g2_mux2_1 _1395_ (.A0(net587),
    .A1(\next_cellsbuf_[30].A ),
    .S(net205),
    .X(_0051_));
 sg13g2_mux2_1 _1396_ (.A0(net841),
    .A1(net587),
    .S(net205),
    .X(_0052_));
 sg13g2_mux2_1 _1397_ (.A0(net880),
    .A1(net841),
    .S(net206),
    .X(_0053_));
 sg13g2_mux2_1 _1398_ (.A0(net567),
    .A1(\next_cellsbuf_[33].A ),
    .S(net206),
    .X(_0054_));
 sg13g2_mux2_1 _1399_ (.A0(net848),
    .A1(net567),
    .S(net206),
    .X(_0055_));
 sg13g2_mux2_1 _1400_ (.A0(net813),
    .A1(\next_cellsbuf_[35].A ),
    .S(net206),
    .X(_0056_));
 sg13g2_mux2_1 _1401_ (.A0(net808),
    .A1(\next_cellsbuf_[36].A ),
    .S(net206),
    .X(_0057_));
 sg13g2_mux2_1 _1402_ (.A0(net565),
    .A1(\next_cellsbuf_[37].A ),
    .S(net200),
    .X(_0058_));
 sg13g2_mux2_1 _1403_ (.A0(net739),
    .A1(net565),
    .S(net200),
    .X(_0059_));
 sg13g2_mux2_1 _1404_ (.A0(net499),
    .A1(\next_cellsbuf_[39].A ),
    .S(net199),
    .X(_0060_));
 sg13g2_mux2_1 _1405_ (.A0(net659),
    .A1(net499),
    .S(net199),
    .X(_0061_));
 sg13g2_mux2_1 _1406_ (.A0(net576),
    .A1(net659),
    .S(net199),
    .X(_0062_));
 sg13g2_mux2_1 _1407_ (.A0(net538),
    .A1(net576),
    .S(net199),
    .X(_0063_));
 sg13g2_mux2_1 _1408_ (.A0(\next_cellsbuf_[44].A ),
    .A1(net538),
    .S(net199),
    .X(_0064_));
 sg13g2_mux2_1 _1409_ (.A0(net857),
    .A1(\next_cellsbuf_[44].A ),
    .S(net197),
    .X(_0065_));
 sg13g2_mux2_1 _1410_ (.A0(net817),
    .A1(\next_cellsbuf_[45].A ),
    .S(net196),
    .X(_0066_));
 sg13g2_mux2_1 _1411_ (.A0(net709),
    .A1(\next_cellsbuf_[46].A ),
    .S(net197),
    .X(_0067_));
 sg13g2_mux2_1 _1412_ (.A0(net804),
    .A1(net709),
    .S(net201),
    .X(_0068_));
 sg13g2_mux2_1 _1413_ (.A0(net640),
    .A1(\next_cellsbuf_[48].A ),
    .S(net201),
    .X(_0069_));
 sg13g2_mux2_1 _1414_ (.A0(net665),
    .A1(net640),
    .S(net203),
    .X(_0070_));
 sg13g2_mux2_1 _1415_ (.A0(net822),
    .A1(net665),
    .S(net203),
    .X(_0071_));
 sg13g2_mux2_1 _1416_ (.A0(net649),
    .A1(\next_cellsbuf_[51].A ),
    .S(net203),
    .X(_0072_));
 sg13g2_mux2_1 _1417_ (.A0(net844),
    .A1(net649),
    .S(net202),
    .X(_0073_));
 sg13g2_mux2_1 _1418_ (.A0(net728),
    .A1(\next_cellsbuf_[53].A ),
    .S(net202),
    .X(_0074_));
 sg13g2_mux2_1 _1419_ (.A0(net765),
    .A1(net728),
    .S(net208),
    .X(_0075_));
 sg13g2_mux2_1 _1420_ (.A0(net655),
    .A1(\next_cellsbuf_[55].A ),
    .S(net208),
    .X(_0076_));
 sg13g2_mux2_1 _1421_ (.A0(net706),
    .A1(net655),
    .S(net209),
    .X(_0077_));
 sg13g2_mux2_1 _1422_ (.A0(net795),
    .A1(net706),
    .S(net210),
    .X(_0078_));
 sg13g2_mux2_1 _1423_ (.A0(net802),
    .A1(net795),
    .S(net210),
    .X(_0079_));
 sg13g2_mux2_1 _1424_ (.A0(net744),
    .A1(\next_cellsbuf_[59].A ),
    .S(net210),
    .X(_0080_));
 sg13g2_mux2_1 _1425_ (.A0(net702),
    .A1(\next_cellsbuf_[60].A ),
    .S(net217),
    .X(_0081_));
 sg13g2_mux2_1 _1426_ (.A0(net762),
    .A1(net702),
    .S(net217),
    .X(_0082_));
 sg13g2_mux2_1 _1427_ (.A0(net657),
    .A1(\next_cellsbuf_[62].A ),
    .S(net217),
    .X(_0083_));
 sg13g2_mux2_1 _1428_ (.A0(net527),
    .A1(net657),
    .S(net214),
    .X(_0084_));
 sg13g2_mux2_1 _1429_ (.A0(net459),
    .A1(net527),
    .S(net215),
    .X(_0085_));
 sg13g2_mux2_1 _1430_ (.A0(\next_cellsbuf_[66].A ),
    .A1(net459),
    .S(net215),
    .X(_0086_));
 sg13g2_mux2_1 _1431_ (.A0(net528),
    .A1(\next_cellsbuf_[66].A ),
    .S(net216),
    .X(_0087_));
 sg13g2_mux2_1 _1432_ (.A0(net849),
    .A1(net528),
    .S(net216),
    .X(_0088_));
 sg13g2_mux2_1 _1433_ (.A0(net833),
    .A1(\next_cellsbuf_[68].A ),
    .S(net215),
    .X(_0089_));
 sg13g2_mux2_1 _1434_ (.A0(net717),
    .A1(\next_cellsbuf_[69].A ),
    .S(net216),
    .X(_0090_));
 sg13g2_mux2_1 _1435_ (.A0(net889),
    .A1(net717),
    .S(net215),
    .X(_0091_));
 sg13g2_mux2_1 _1436_ (.A0(net890),
    .A1(net889),
    .S(net215),
    .X(_0092_));
 sg13g2_mux2_1 _1437_ (.A0(net756),
    .A1(\next_cellsbuf_[72].A ),
    .S(net215),
    .X(_0093_));
 sg13g2_mux2_1 _1438_ (.A0(net549),
    .A1(\next_cellsbuf_[73].A ),
    .S(net215),
    .X(_0094_));
 sg13g2_mux2_1 _1439_ (.A0(net667),
    .A1(net549),
    .S(net215),
    .X(_0095_));
 sg13g2_mux2_1 _1440_ (.A0(net581),
    .A1(\next_cellsbuf_[75].A ),
    .S(net214),
    .X(_0096_));
 sg13g2_mux2_1 _1441_ (.A0(net531),
    .A1(\next_cellsbuf_[76].A ),
    .S(net214),
    .X(_0097_));
 sg13g2_mux2_1 _1442_ (.A0(net700),
    .A1(net531),
    .S(net214),
    .X(_0098_));
 sg13g2_mux2_1 _1443_ (.A0(net675),
    .A1(\next_cellsbuf_[78].A ),
    .S(net214),
    .X(_0099_));
 sg13g2_mux2_1 _1444_ (.A0(net787),
    .A1(net675),
    .S(net210),
    .X(_0100_));
 sg13g2_mux2_1 _1445_ (.A0(net683),
    .A1(\next_cellsbuf_[80].A ),
    .S(net210),
    .X(_0101_));
 sg13g2_mux2_1 _1446_ (.A0(net807),
    .A1(net683),
    .S(net210),
    .X(_0102_));
 sg13g2_mux2_1 _1447_ (.A0(net647),
    .A1(\next_cellsbuf_[82].A ),
    .S(net213),
    .X(_0103_));
 sg13g2_mux2_1 _1448_ (.A0(net719),
    .A1(net647),
    .S(net208),
    .X(_0104_));
 sg13g2_mux2_1 _1449_ (.A0(net695),
    .A1(\next_cellsbuf_[84].A ),
    .S(net208),
    .X(_0105_));
 sg13g2_mux2_1 _1450_ (.A0(net671),
    .A1(\next_cellsbuf_[85].A ),
    .S(net208),
    .X(_0106_));
 sg13g2_mux2_1 _1451_ (.A0(net682),
    .A1(net671),
    .S(net208),
    .X(_0107_));
 sg13g2_mux2_1 _1452_ (.A0(net773),
    .A1(net682),
    .S(net208),
    .X(_0108_));
 sg13g2_mux2_1 _1453_ (.A0(net827),
    .A1(net773),
    .S(net202),
    .X(_0109_));
 sg13g2_mux2_1 _1454_ (.A0(net842),
    .A1(net827),
    .S(net202),
    .X(_0110_));
 sg13g2_mux2_1 _1455_ (.A0(net758),
    .A1(\next_cellsbuf_[90].A ),
    .S(net202),
    .X(_0111_));
 sg13g2_mux2_1 _1456_ (.A0(net792),
    .A1(net758),
    .S(net202),
    .X(_0112_));
 sg13g2_mux2_1 _1457_ (.A0(net815),
    .A1(net792),
    .S(net201),
    .X(_0113_));
 sg13g2_mux2_1 _1458_ (.A0(net642),
    .A1(\next_cellsbuf_[93].A ),
    .S(net201),
    .X(_0114_));
 sg13g2_mux2_1 _1459_ (.A0(net646),
    .A1(net642),
    .S(net201),
    .X(_0115_));
 sg13g2_mux2_1 _1460_ (.A0(net905),
    .A1(net646),
    .S(net201),
    .X(_0116_));
 sg13g2_mux2_1 _1461_ (.A0(net824),
    .A1(\next_cellsbuf_[96].A ),
    .S(net201),
    .X(_0117_));
 sg13g2_mux2_1 _1462_ (.A0(net869),
    .A1(net824),
    .S(net201),
    .X(_0118_));
 sg13g2_mux2_1 _1463_ (.A0(net725),
    .A1(\next_cellsbuf_[98].A ),
    .S(net196),
    .X(_0119_));
 sg13g2_mux2_1 _1464_ (.A0(net559),
    .A1(\next_cellsbuf_[99].A ),
    .S(net196),
    .X(_0120_));
 sg13g2_mux2_1 _1465_ (.A0(net898),
    .A1(net559),
    .S(net196),
    .X(_0121_));
 sg13g2_mux2_1 _1466_ (.A0(net573),
    .A1(\next_cellsbuf_[101].A ),
    .S(net196),
    .X(_0122_));
 sg13g2_mux2_1 _1467_ (.A0(net510),
    .A1(\next_cellsbuf_[102].A ),
    .S(net196),
    .X(_0123_));
 sg13g2_mux2_1 _1468_ (.A0(net537),
    .A1(net510),
    .S(net196),
    .X(_0124_));
 sg13g2_mux2_1 _1469_ (.A0(net850),
    .A1(net537),
    .S(net197),
    .X(_0125_));
 sg13g2_mux2_1 _1470_ (.A0(net777),
    .A1(\next_cellsbuf_[105].A ),
    .S(net196),
    .X(_0126_));
 sg13g2_mux2_1 _1471_ (.A0(net668),
    .A1(\next_cellsbuf_[106].A ),
    .S(net194),
    .X(_0127_));
 sg13g2_mux2_1 _1472_ (.A0(net515),
    .A1(\next_cellsbuf_[107].A ),
    .S(net194),
    .X(_0128_));
 sg13g2_mux2_1 _1473_ (.A0(net505),
    .A1(net515),
    .S(net194),
    .X(_0129_));
 sg13g2_mux2_1 _1474_ (.A0(net453),
    .A1(net505),
    .S(net194),
    .X(_0130_));
 sg13g2_mux2_1 _1475_ (.A0(\next_cellsbuf_[111].A ),
    .A1(net453),
    .S(net194),
    .X(_0131_));
 sg13g2_mux2_1 _1476_ (.A0(net691),
    .A1(\next_cellsbuf_[111].A ),
    .S(net194),
    .X(_0132_));
 sg13g2_mux2_1 _1477_ (.A0(net485),
    .A1(\next_cellsbuf_[112].A ),
    .S(net194),
    .X(_0133_));
 sg13g2_mux2_1 _1478_ (.A0(net514),
    .A1(net485),
    .S(net195),
    .X(_0134_));
 sg13g2_mux2_1 _1479_ (.A0(net506),
    .A1(\next_cellsbuf_[114].A ),
    .S(net195),
    .X(_0135_));
 sg13g2_mux2_1 _1480_ (.A0(net575),
    .A1(net506),
    .S(net195),
    .X(_0136_));
 sg13g2_mux2_1 _1481_ (.A0(net831),
    .A1(net575),
    .S(net195),
    .X(_0137_));
 sg13g2_mux2_1 _1482_ (.A0(net894),
    .A1(net831),
    .S(net195),
    .X(_0138_));
 sg13g2_mux2_1 _1483_ (.A0(net607),
    .A1(\next_cellsbuf_[118].A ),
    .S(net194),
    .X(_0139_));
 sg13g2_mux2_1 _1484_ (.A0(net801),
    .A1(net607),
    .S(net195),
    .X(_0140_));
 sg13g2_mux2_1 _1485_ (.A0(net839),
    .A1(net801),
    .S(net198),
    .X(_0141_));
 sg13g2_mux2_1 _1486_ (.A0(net632),
    .A1(\next_cellsbuf_[121].A ),
    .S(net198),
    .X(_0142_));
 sg13g2_mux2_1 _1487_ (.A0(net763),
    .A1(net632),
    .S(net198),
    .X(_0143_));
 sg13g2_mux2_1 _1488_ (.A0(net517),
    .A1(\next_cellsbuf_[123].A ),
    .S(net198),
    .X(_0144_));
 sg13g2_mux2_1 _1489_ (.A0(net681),
    .A1(net517),
    .S(net198),
    .X(_0145_));
 sg13g2_mux2_1 _1490_ (.A0(net463),
    .A1(net681),
    .S(net198),
    .X(_0146_));
 sg13g2_mux2_1 _1491_ (.A0(\next_cellsbuf_[127].A ),
    .A1(net463),
    .S(net200),
    .X(_0147_));
 sg13g2_mux2_1 _1492_ (.A0(net622),
    .A1(\next_cellsbuf_[127].A ),
    .S(net200),
    .X(_0148_));
 sg13g2_mux2_1 _1493_ (.A0(net791),
    .A1(net622),
    .S(net200),
    .X(_0149_));
 sg13g2_mux2_1 _1494_ (.A0(net697),
    .A1(\next_cellsbuf_[129].A ),
    .S(net198),
    .X(_0150_));
 sg13g2_mux2_1 _1495_ (.A0(net651),
    .A1(\next_cellsbuf_[130].A ),
    .S(net198),
    .X(_0151_));
 sg13g2_mux2_1 _1496_ (.A0(net624),
    .A1(\next_cellsbuf_[131].A ),
    .S(net199),
    .X(_0152_));
 sg13g2_mux2_1 _1497_ (.A0(net620),
    .A1(\next_cellsbuf_[132].A ),
    .S(net199),
    .X(_0153_));
 sg13g2_mux2_1 _1498_ (.A0(net598),
    .A1(\next_cellsbuf_[133].A ),
    .S(net199),
    .X(_0154_));
 sg13g2_mux2_1 _1499_ (.A0(net716),
    .A1(net598),
    .S(net206),
    .X(_0155_));
 sg13g2_mux2_1 _1500_ (.A0(net738),
    .A1(net716),
    .S(net206),
    .X(_0156_));
 sg13g2_mux2_1 _1501_ (.A0(net503),
    .A1(\next_cellsbuf_[136].A ),
    .S(net206),
    .X(_0157_));
 sg13g2_mux2_1 _1502_ (.A0(net501),
    .A1(\next_cellsbuf_[137].A ),
    .S(net205),
    .X(_0158_));
 sg13g2_mux2_1 _1503_ (.A0(net687),
    .A1(net501),
    .S(net204),
    .X(_0159_));
 sg13g2_mux2_1 _1504_ (.A0(net569),
    .A1(net687),
    .S(net204),
    .X(_0160_));
 sg13g2_mux2_1 _1505_ (.A0(\next_cellsbuf_[141].A ),
    .A1(net569),
    .S(net204),
    .X(_0161_));
 sg13g2_mux2_1 _1506_ (.A0(net811),
    .A1(\next_cellsbuf_[141].A ),
    .S(net204),
    .X(_0162_));
 sg13g2_mux2_1 _1507_ (.A0(net662),
    .A1(\next_cellsbuf_[142].A ),
    .S(net204),
    .X(_0163_));
 sg13g2_mux2_1 _1508_ (.A0(net670),
    .A1(net662),
    .S(net204),
    .X(_0164_));
 sg13g2_mux2_1 _1509_ (.A0(net806),
    .A1(net670),
    .S(net204),
    .X(_0165_));
 sg13g2_mux2_1 _1510_ (.A0(net884),
    .A1(net806),
    .S(net202),
    .X(_0166_));
 sg13g2_mux2_1 _1511_ (.A0(net779),
    .A1(\next_cellsbuf_[146].A ),
    .S(net203),
    .X(_0167_));
 sg13g2_mux2_1 _1512_ (.A0(net584),
    .A1(\next_cellsbuf_[147].A ),
    .S(net202),
    .X(_0168_));
 sg13g2_mux2_1 _1513_ (.A0(net753),
    .A1(net584),
    .S(net203),
    .X(_0169_));
 sg13g2_mux2_1 _1514_ (.A0(net751),
    .A1(\next_cellsbuf_[149].A ),
    .S(net209),
    .X(_0170_));
 sg13g2_mux2_1 _1515_ (.A0(net766),
    .A1(net751),
    .S(net209),
    .X(_0171_));
 sg13g2_mux2_1 _1516_ (.A0(net754),
    .A1(\next_cellsbuf_[151].A ),
    .S(net209),
    .X(_0172_));
 sg13g2_mux2_1 _1517_ (.A0(net713),
    .A1(\next_cellsbuf_[152].A ),
    .S(net209),
    .X(_0173_));
 sg13g2_mux2_1 _1518_ (.A0(net685),
    .A1(\next_cellsbuf_[153].A ),
    .S(net208),
    .X(_0174_));
 sg13g2_mux2_1 _1519_ (.A0(net616),
    .A1(\next_cellsbuf_[154].A ),
    .S(net212),
    .X(_0175_));
 sg13g2_mux2_1 _1520_ (.A0(net589),
    .A1(\next_cellsbuf_[155].A ),
    .S(net212),
    .X(_0176_));
 sg13g2_mux2_1 _1521_ (.A0(net512),
    .A1(\next_cellsbuf_[156].A ),
    .S(net212),
    .X(_0177_));
 sg13g2_mux2_1 _1522_ (.A0(net734),
    .A1(net512),
    .S(net212),
    .X(_0178_));
 sg13g2_mux2_1 _1523_ (.A0(\next_cellsbuf_[159].A ),
    .A1(net734),
    .S(net212),
    .X(_0179_));
 sg13g2_and2_1 _1524_ (.A(\fract_x[0] ),
    .B(net969),
    .X(_0371_));
 sg13g2_and4_2 _1525_ (.A(\fract_x[0] ),
    .B(net972),
    .C(net445),
    .D(\cell_x[0] ),
    .X(_0372_));
 sg13g2_nand2_1 _1526_ (.Y(_0373_),
    .A(net967),
    .B(_0372_));
 sg13g2_nor2_1 _1527_ (.A(\cell_x[3] ),
    .B(\cell_x[4] ),
    .Y(_0374_));
 sg13g2_nand3_1 _1528_ (.B(_0524_),
    .C(_0374_),
    .A(\cell_x[7] ),
    .Y(_0375_));
 sg13g2_o21ai_1 _1529_ (.B1(net252),
    .Y(_0376_),
    .A1(_0373_),
    .A2(_0375_));
 sg13g2_nor2_1 _1530_ (.A(_0442_),
    .B(net222),
    .Y(_0180_));
 sg13g2_nor3_1 _1531_ (.A(net970),
    .B(_0371_),
    .C(net221),
    .Y(_0181_));
 sg13g2_xnor2_1 _1532_ (.Y(_0377_),
    .A(net951),
    .B(_0371_));
 sg13g2_nor2_1 _1533_ (.A(net222),
    .B(net952),
    .Y(_0182_));
 sg13g2_a21oi_1 _1534_ (.A1(\cell_x[0] ),
    .A2(_0371_),
    .Y(_0378_),
    .B1(net445));
 sg13g2_nor3_1 _1535_ (.A(net251),
    .B(_0372_),
    .C(net446),
    .Y(_0183_));
 sg13g2_o21ai_1 _1536_ (.B1(net252),
    .Y(_0379_),
    .A1(net962),
    .A2(_0372_));
 sg13g2_nor2b_1 _1537_ (.A(_0379_),
    .B_N(_0373_),
    .Y(_0184_));
 sg13g2_and3_1 _1538_ (.X(_0380_),
    .A(\cell_x[2] ),
    .B(net938),
    .C(_0372_));
 sg13g2_a21oi_1 _1539_ (.A1(\cell_x[2] ),
    .A2(_0372_),
    .Y(_0381_),
    .B1(net938));
 sg13g2_nor3_1 _1540_ (.A(net222),
    .B(_0380_),
    .C(net939),
    .Y(_0185_));
 sg13g2_and2_1 _1541_ (.A(_0446_),
    .B(_0372_),
    .X(_0382_));
 sg13g2_nor2_1 _1542_ (.A(net955),
    .B(_0380_),
    .Y(_0383_));
 sg13g2_nor3_1 _1543_ (.A(net222),
    .B(_0382_),
    .C(net956),
    .Y(_0186_));
 sg13g2_xnor2_1 _1544_ (.Y(_0384_),
    .A(net959),
    .B(_0382_));
 sg13g2_nor2_1 _1545_ (.A(net222),
    .B(_0384_),
    .Y(_0187_));
 sg13g2_a21oi_1 _1546_ (.A1(\cell_x[5] ),
    .A2(_0382_),
    .Y(_0385_),
    .B1(net913));
 sg13g2_nand3_1 _1547_ (.B(net913),
    .C(_0382_),
    .A(net973),
    .Y(_0386_));
 sg13g2_nand2b_1 _1548_ (.Y(_0387_),
    .B(_0386_),
    .A_N(net222));
 sg13g2_nor2_1 _1549_ (.A(net914),
    .B(_0387_),
    .Y(_0188_));
 sg13g2_xor2_1 _1550_ (.B(_0386_),
    .A(net957),
    .X(_0388_));
 sg13g2_nor2_1 _1551_ (.A(net221),
    .B(net958),
    .Y(_0189_));
 sg13g2_mux2_1 _1552_ (.A0(net876),
    .A1(net465),
    .S(net239),
    .X(_0190_));
 sg13g2_mux2_1 _1553_ (.A0(net465),
    .A1(\cellsbuf_[2].A ),
    .S(net245),
    .X(_0191_));
 sg13g2_mux2_1 _1554_ (.A0(net912),
    .A1(net830),
    .S(net239),
    .X(_0192_));
 sg13g2_mux2_1 _1555_ (.A0(net830),
    .A1(net722),
    .S(net239),
    .X(_0193_));
 sg13g2_mux2_1 _1556_ (.A0(net722),
    .A1(net644),
    .S(net239),
    .X(_0194_));
 sg13g2_mux2_1 _1557_ (.A0(net644),
    .A1(\cellsbuf_[6].A ),
    .S(net239),
    .X(_0195_));
 sg13g2_mux2_1 _1558_ (.A0(net689),
    .A1(\cellsbuf_[7].A ),
    .S(net239),
    .X(_0196_));
 sg13g2_mux2_1 _1559_ (.A0(net879),
    .A1(net579),
    .S(net239),
    .X(_0197_));
 sg13g2_mux2_1 _1560_ (.A0(net579),
    .A1(\cellsbuf_[9].A ),
    .S(net239),
    .X(_0198_));
 sg13g2_mux2_1 _1561_ (.A0(net873),
    .A1(net586),
    .S(net240),
    .X(_0199_));
 sg13g2_mux2_1 _1562_ (.A0(net586),
    .A1(net489),
    .S(net240),
    .X(_0200_));
 sg13g2_mux2_1 _1563_ (.A0(net489),
    .A1(\cellsbuf_[12].A ),
    .S(net240),
    .X(_0201_));
 sg13g2_mux2_1 _1564_ (.A0(net853),
    .A1(net639),
    .S(net240),
    .X(_0202_));
 sg13g2_mux2_1 _1565_ (.A0(net639),
    .A1(net449),
    .S(net242),
    .X(_0203_));
 sg13g2_mux2_1 _1566_ (.A0(net449),
    .A1(\cellsbuf_[15].A ),
    .S(net242),
    .X(_0204_));
 sg13g2_mux2_1 _1567_ (.A0(net851),
    .A1(\cellsbuf_[16].A ),
    .S(net242),
    .X(_0205_));
 sg13g2_mux2_1 _1568_ (.A0(net882),
    .A1(net473),
    .S(net242),
    .X(_0206_));
 sg13g2_mux2_1 _1569_ (.A0(net473),
    .A1(\cellsbuf_[18].A ),
    .S(net246),
    .X(_0207_));
 sg13g2_mux2_1 _1570_ (.A0(net547),
    .A1(\cellsbuf_[19].A ),
    .S(net246),
    .X(_0208_));
 sg13g2_mux2_1 _1571_ (.A0(net900),
    .A1(\cellsbuf_[20].A ),
    .S(net246),
    .X(_0209_));
 sg13g2_mux2_1 _1572_ (.A0(net908),
    .A1(net749),
    .S(net249),
    .X(_0210_));
 sg13g2_mux2_1 _1573_ (.A0(net749),
    .A1(\cellsbuf_[22].A ),
    .S(net249),
    .X(_0211_));
 sg13g2_mux2_1 _1574_ (.A0(net907),
    .A1(net870),
    .S(net243),
    .X(_0212_));
 sg13g2_mux2_1 _1575_ (.A0(net870),
    .A1(\cellsbuf_[24].A ),
    .S(net243),
    .X(_0213_));
 sg13g2_mux2_1 _1576_ (.A0(net878),
    .A1(net630),
    .S(net242),
    .X(_0214_));
 sg13g2_mux2_1 _1577_ (.A0(net630),
    .A1(\cellsbuf_[26].A ),
    .S(net242),
    .X(_0215_));
 sg13g2_mux2_1 _1578_ (.A0(net797),
    .A1(net552),
    .S(net240),
    .X(_0216_));
 sg13g2_mux2_1 _1579_ (.A0(net552),
    .A1(\cellsbuf_[28].A ),
    .S(net240),
    .X(_0217_));
 sg13g2_mux2_1 _1580_ (.A0(net863),
    .A1(net715),
    .S(net240),
    .X(_0218_));
 sg13g2_mux2_1 _1581_ (.A0(net715),
    .A1(net711),
    .S(net240),
    .X(_0219_));
 sg13g2_mux2_1 _1582_ (.A0(net711),
    .A1(\cellsbuf_[31].A ),
    .S(net236),
    .X(_0220_));
 sg13g2_mux2_1 _1583_ (.A0(net828),
    .A1(net523),
    .S(net236),
    .X(_0221_));
 sg13g2_mux2_1 _1584_ (.A0(net523),
    .A1(\cellsbuf_[33].A ),
    .S(net236),
    .X(_0222_));
 sg13g2_mux2_1 _1585_ (.A0(net561),
    .A1(\cellsbuf_[34].A ),
    .S(net236),
    .X(_0223_));
 sg13g2_mux2_1 _1586_ (.A0(net731),
    .A1(\cellsbuf_[35].A ),
    .S(net236),
    .X(_0224_));
 sg13g2_mux2_1 _1587_ (.A0(net747),
    .A1(net493),
    .S(net235),
    .X(_0225_));
 sg13g2_mux2_1 _1588_ (.A0(net493),
    .A1(\cellsbuf_[37].A ),
    .S(net235),
    .X(_0226_));
 sg13g2_mux2_1 _1589_ (.A0(net664),
    .A1(net455),
    .S(net235),
    .X(_0227_));
 sg13g2_mux2_1 _1590_ (.A0(net455),
    .A1(\cellsbuf_[39].A ),
    .S(net235),
    .X(_0228_));
 sg13g2_mux2_1 _1591_ (.A0(net881),
    .A1(net860),
    .S(net237),
    .X(_0229_));
 sg13g2_mux2_1 _1592_ (.A0(net860),
    .A1(\cellsbuf_[41].A ),
    .S(net229),
    .X(_0230_));
 sg13g2_mux2_1 _1593_ (.A0(net866),
    .A1(net583),
    .S(net229),
    .X(_0231_));
 sg13g2_mux2_1 _1594_ (.A0(net583),
    .A1(net467),
    .S(net229),
    .X(_0232_));
 sg13g2_mux2_1 _1595_ (.A0(net467),
    .A1(\cellsbuf_[44].A ),
    .S(net229),
    .X(_0233_));
 sg13g2_mux2_1 _1596_ (.A0(net730),
    .A1(net564),
    .S(net227),
    .X(_0234_));
 sg13g2_mux2_1 _1597_ (.A0(net564),
    .A1(net555),
    .S(net227),
    .X(_0235_));
 sg13g2_mux2_1 _1598_ (.A0(net555),
    .A1(\cellsbuf_[47].A ),
    .S(net227),
    .X(_0236_));
 sg13g2_mux2_1 _1599_ (.A0(net688),
    .A1(net554),
    .S(net227),
    .X(_0237_));
 sg13g2_mux2_1 _1600_ (.A0(net554),
    .A1(net497),
    .S(net227),
    .X(_0238_));
 sg13g2_mux2_1 _1601_ (.A0(net497),
    .A1(\cellsbuf_[50].A ),
    .S(net227),
    .X(_0239_));
 sg13g2_mux2_1 _1602_ (.A0(net782),
    .A1(\cellsbuf_[51].A ),
    .S(net227),
    .X(_0240_));
 sg13g2_mux2_1 _1603_ (.A0(net875),
    .A1(net609),
    .S(net224),
    .X(_0241_));
 sg13g2_mux2_1 _1604_ (.A0(net609),
    .A1(\cellsbuf_[53].A ),
    .S(net224),
    .X(_0242_));
 sg13g2_mux2_1 _1605_ (.A0(net790),
    .A1(net769),
    .S(net224),
    .X(_0243_));
 sg13g2_mux2_1 _1606_ (.A0(net769),
    .A1(net542),
    .S(net224),
    .X(_0244_));
 sg13g2_mux2_1 _1607_ (.A0(net542),
    .A1(net461),
    .S(net224),
    .X(_0245_));
 sg13g2_mux2_1 _1608_ (.A0(net461),
    .A1(\cellsbuf_[57].A ),
    .S(net224),
    .X(_0246_));
 sg13g2_mux2_1 _1609_ (.A0(net893),
    .A1(net481),
    .S(net224),
    .X(_0247_));
 sg13g2_mux2_1 _1610_ (.A0(net481),
    .A1(\cellsbuf_[59].A ),
    .S(net223),
    .X(_0248_));
 sg13g2_mux2_1 _1611_ (.A0(net748),
    .A1(net626),
    .S(net223),
    .X(_0249_));
 sg13g2_mux2_1 _1612_ (.A0(net626),
    .A1(\cellsbuf_[61].A ),
    .S(net223),
    .X(_0250_));
 sg13g2_mux2_1 _1613_ (.A0(net660),
    .A1(\cellsbuf_[62].A ),
    .S(net223),
    .X(_0251_));
 sg13g2_mux2_1 _1614_ (.A0(net867),
    .A1(\cellsbuf_[63].A ),
    .S(net223),
    .X(_0252_));
 sg13g2_mux2_1 _1615_ (.A0(\cellsbuf_[63].A ),
    .A1(net736),
    .S(net223),
    .X(_0253_));
 sg13g2_mux2_1 _1616_ (.A0(net736),
    .A1(net829),
    .S(net223),
    .X(_0254_));
 sg13g2_mux2_1 _1617_ (.A0(net829),
    .A1(net823),
    .S(net223),
    .X(_0255_));
 sg13g2_mux2_1 _1618_ (.A0(net823),
    .A1(net457),
    .S(net225),
    .X(_0256_));
 sg13g2_mux2_1 _1619_ (.A0(net457),
    .A1(\cellsbuf_[68].A ),
    .S(net225),
    .X(_0257_));
 sg13g2_mux2_1 _1620_ (.A0(\cellsbuf_[68].A ),
    .A1(net785),
    .S(net225),
    .X(_0258_));
 sg13g2_mux2_1 _1621_ (.A0(net785),
    .A1(net557),
    .S(net225),
    .X(_0259_));
 sg13g2_mux2_1 _1622_ (.A0(net557),
    .A1(\cellsbuf_[71].A ),
    .S(net226),
    .X(_0260_));
 sg13g2_mux2_1 _1623_ (.A0(net593),
    .A1(\cellsbuf_[72].A ),
    .S(net226),
    .X(_0261_));
 sg13g2_mux2_1 _1624_ (.A0(net768),
    .A1(net540),
    .S(net225),
    .X(_0262_));
 sg13g2_mux2_1 _1625_ (.A0(net540),
    .A1(\cellsbuf_[74].A ),
    .S(net225),
    .X(_0263_));
 sg13g2_mux2_1 _1626_ (.A0(net611),
    .A1(\cellsbuf_[75].A ),
    .S(net225),
    .X(_0264_));
 sg13g2_mux2_1 _1627_ (.A0(net820),
    .A1(\cellsbuf_[76].A ),
    .S(net225),
    .X(_0265_));
 sg13g2_mux2_1 _1628_ (.A0(net837),
    .A1(\cellsbuf_[77].A ),
    .S(net231),
    .X(_0266_));
 sg13g2_mux2_1 _1629_ (.A0(net883),
    .A1(net874),
    .S(net234),
    .X(_0267_));
 sg13g2_mux2_1 _1630_ (.A0(net874),
    .A1(net862),
    .S(net231),
    .X(_0268_));
 sg13g2_mux2_1 _1631_ (.A0(net862),
    .A1(net447),
    .S(net231),
    .X(_0269_));
 sg13g2_mux2_1 _1632_ (.A0(net447),
    .A1(\cellsbuf_[81].A ),
    .S(net231),
    .X(_0270_));
 sg13g2_mux2_1 _1633_ (.A0(net832),
    .A1(net451),
    .S(net231),
    .X(_0271_));
 sg13g2_mux2_1 _1634_ (.A0(net451),
    .A1(\cellsbuf_[83].A ),
    .S(net231),
    .X(_0272_));
 sg13g2_mux2_1 _1635_ (.A0(net784),
    .A1(net563),
    .S(net231),
    .X(_0273_));
 sg13g2_mux2_1 _1636_ (.A0(net563),
    .A1(net530),
    .S(net231),
    .X(_0274_));
 sg13g2_mux2_1 _1637_ (.A0(net530),
    .A1(net519),
    .S(net232),
    .X(_0275_));
 sg13g2_mux2_1 _1638_ (.A0(net519),
    .A1(\cellsbuf_[87].A ),
    .S(net232),
    .X(_0276_));
 sg13g2_mux2_1 _1639_ (.A0(net693),
    .A1(\cellsbuf_[88].A ),
    .S(net232),
    .X(_0277_));
 sg13g2_mux2_1 _1640_ (.A0(net727),
    .A1(net479),
    .S(net232),
    .X(_0278_));
 sg13g2_mux2_1 _1641_ (.A0(net479),
    .A1(\cellsbuf_[90].A ),
    .S(net232),
    .X(_0279_));
 sg13g2_mux2_1 _1642_ (.A0(net902),
    .A1(net680),
    .S(net232),
    .X(_0280_));
 sg13g2_mux2_1 _1643_ (.A0(net680),
    .A1(net577),
    .S(net232),
    .X(_0281_));
 sg13g2_mux2_1 _1644_ (.A0(net577),
    .A1(\cellsbuf_[93].A ),
    .S(net232),
    .X(_0282_));
 sg13g2_mux2_1 _1645_ (.A0(net699),
    .A1(net533),
    .S(net233),
    .X(_0283_));
 sg13g2_mux2_1 _1646_ (.A0(net533),
    .A1(\cellsbuf_[95].A ),
    .S(net233),
    .X(_0284_));
 sg13g2_mux2_1 _1647_ (.A0(net826),
    .A1(net771),
    .S(net233),
    .X(_0285_));
 sg13g2_mux2_1 _1648_ (.A0(net771),
    .A1(\cellsbuf_[97].A ),
    .S(net233),
    .X(_0286_));
 sg13g2_mux2_1 _1649_ (.A0(net776),
    .A1(net495),
    .S(net233),
    .X(_0287_));
 sg13g2_mux2_1 _1650_ (.A0(net495),
    .A1(\cellsbuf_[99].A ),
    .S(net233),
    .X(_0288_));
 sg13g2_mux2_1 _1651_ (.A0(net673),
    .A1(\cellsbuf_[100].A ),
    .S(net236),
    .X(_0289_));
 sg13g2_mux2_1 _1652_ (.A0(net770),
    .A1(net491),
    .S(net235),
    .X(_0290_));
 sg13g2_mux2_1 _1653_ (.A0(net491),
    .A1(\cellsbuf_[102].A ),
    .S(net235),
    .X(_0291_));
 sg13g2_mux2_1 _1654_ (.A0(net746),
    .A1(net475),
    .S(net235),
    .X(_0292_));
 sg13g2_mux2_1 _1655_ (.A0(net475),
    .A1(\cellsbuf_[104].A ),
    .S(net229),
    .X(_0293_));
 sg13g2_mux2_1 _1656_ (.A0(net872),
    .A1(net816),
    .S(net229),
    .X(_0294_));
 sg13g2_mux2_1 _1657_ (.A0(net816),
    .A1(net760),
    .S(net229),
    .X(_0295_));
 sg13g2_mux2_1 _1658_ (.A0(net760),
    .A1(net551),
    .S(net227),
    .X(_0296_));
 sg13g2_mux2_1 _1659_ (.A0(net551),
    .A1(net477),
    .S(net228),
    .X(_0297_));
 sg13g2_mux2_1 _1660_ (.A0(net477),
    .A1(\cellsbuf_[109].A ),
    .S(net228),
    .X(_0298_));
 sg13g2_mux2_1 _1661_ (.A0(net793),
    .A1(\cellsbuf_[110].A ),
    .S(net228),
    .X(_0299_));
 sg13g2_mux2_1 _1662_ (.A0(net835),
    .A1(net613),
    .S(net228),
    .X(_0300_));
 sg13g2_mux2_1 _1663_ (.A0(net613),
    .A1(net597),
    .S(net228),
    .X(_0301_));
 sg13g2_mux2_1 _1664_ (.A0(net597),
    .A1(net471),
    .S(net228),
    .X(_0302_));
 sg13g2_mux2_1 _1665_ (.A0(net471),
    .A1(\cellsbuf_[114].A ),
    .S(net228),
    .X(_0303_));
 sg13g2_mux2_1 _1666_ (.A0(net707),
    .A1(\cellsbuf_[115].A ),
    .S(net228),
    .X(_0304_));
 sg13g2_mux2_1 _1667_ (.A0(net847),
    .A1(net796),
    .S(net229),
    .X(_0305_));
 sg13g2_mux2_1 _1668_ (.A0(net796),
    .A1(net743),
    .S(net230),
    .X(_0306_));
 sg13g2_mux2_1 _1669_ (.A0(net743),
    .A1(net535),
    .S(net230),
    .X(_0307_));
 sg13g2_mux2_1 _1670_ (.A0(net535),
    .A1(\cellsbuf_[119].A ),
    .S(net230),
    .X(_0308_));
 sg13g2_mux2_1 _1671_ (.A0(net859),
    .A1(net677),
    .S(net237),
    .X(_0309_));
 sg13g2_mux2_1 _1672_ (.A0(net677),
    .A1(net545),
    .S(net235),
    .X(_0310_));
 sg13g2_mux2_1 _1673_ (.A0(net545),
    .A1(\cellsbuf_[122].A ),
    .S(net237),
    .X(_0311_));
 sg13g2_mux2_1 _1674_ (.A0(net605),
    .A1(\cellsbuf_[123].A ),
    .S(net237),
    .X(_0312_));
 sg13g2_mux2_1 _1675_ (.A0(net899),
    .A1(net819),
    .S(net237),
    .X(_0313_));
 sg13g2_mux2_1 _1676_ (.A0(net819),
    .A1(net628),
    .S(net237),
    .X(_0314_));
 sg13g2_mux2_1 _1677_ (.A0(net628),
    .A1(\cellsbuf_[126].A ),
    .S(net236),
    .X(_0315_));
 sg13g2_mux2_1 _1678_ (.A0(net723),
    .A1(\cellsbuf_[127].A ),
    .S(net236),
    .X(_0316_));
 sg13g2_mux2_1 _1679_ (.A0(net892),
    .A1(net638),
    .S(net241),
    .X(_0317_));
 sg13g2_mux2_1 _1680_ (.A0(net638),
    .A1(net600),
    .S(net241),
    .X(_0318_));
 sg13g2_mux2_1 _1681_ (.A0(net600),
    .A1(net521),
    .S(net241),
    .X(_0319_));
 sg13g2_mux2_1 _1682_ (.A0(net521),
    .A1(\cellsbuf_[131].A ),
    .S(net241),
    .X(_0320_));
 sg13g2_mux2_1 _1683_ (.A0(net733),
    .A1(net443),
    .S(net243),
    .X(_0321_));
 sg13g2_mux2_1 _1684_ (.A0(net443),
    .A1(\cellsbuf_[133].A ),
    .S(net243),
    .X(_0322_));
 sg13g2_mux2_1 _1685_ (.A0(net877),
    .A1(net740),
    .S(net242),
    .X(_0323_));
 sg13g2_mux2_1 _1686_ (.A0(net740),
    .A1(net483),
    .S(net242),
    .X(_0324_));
 sg13g2_mux2_1 _1687_ (.A0(net483),
    .A1(\cellsbuf_[136].A ),
    .S(net246),
    .X(_0325_));
 sg13g2_mux2_1 _1688_ (.A0(net843),
    .A1(net781),
    .S(net246),
    .X(_0326_));
 sg13g2_mux2_1 _1689_ (.A0(net781),
    .A1(net767),
    .S(net246),
    .X(_0327_));
 sg13g2_mux2_1 _1690_ (.A0(net767),
    .A1(net678),
    .S(net246),
    .X(_0328_));
 sg13g2_mux2_1 _1691_ (.A0(net678),
    .A1(\cellsbuf_[140].A ),
    .S(net246),
    .X(_0329_));
 sg13g2_mux2_1 _1692_ (.A0(net888),
    .A1(net571),
    .S(net247),
    .X(_0330_));
 sg13g2_mux2_1 _1693_ (.A0(net571),
    .A1(\cellsbuf_[142].A ),
    .S(net247),
    .X(_0331_));
 sg13g2_mux2_1 _1694_ (.A0(net909),
    .A1(net741),
    .S(net247),
    .X(_0332_));
 sg13g2_mux2_1 _1695_ (.A0(net741),
    .A1(\cellsbuf_[144].A ),
    .S(net247),
    .X(_0333_));
 sg13g2_mux2_1 _1696_ (.A0(net896),
    .A1(net543),
    .S(net247),
    .X(_0334_));
 sg13g2_mux2_1 _1697_ (.A0(net543),
    .A1(\cellsbuf_[146].A ),
    .S(net249),
    .X(_0335_));
 sg13g2_mux2_1 _1698_ (.A0(net906),
    .A1(net897),
    .S(net247),
    .X(_0336_));
 sg13g2_mux2_1 _1699_ (.A0(net897),
    .A1(net799),
    .S(net247),
    .X(_0337_));
 sg13g2_mux2_1 _1700_ (.A0(net799),
    .A1(\cellsbuf_[149].A ),
    .S(net247),
    .X(_0338_));
 sg13g2_mux2_1 _1701_ (.A0(net895),
    .A1(net701),
    .S(net248),
    .X(_0339_));
 sg13g2_mux2_1 _1702_ (.A0(net701),
    .A1(net469),
    .S(net248),
    .X(_0340_));
 sg13g2_mux2_1 _1703_ (.A0(net469),
    .A1(\cellsbuf_[152].A ),
    .S(net248),
    .X(_0341_));
 sg13g2_mux2_1 _1704_ (.A0(net836),
    .A1(net803),
    .S(net248),
    .X(_0342_));
 sg13g2_mux2_1 _1705_ (.A0(net803),
    .A1(net653),
    .S(net248),
    .X(_0343_));
 sg13g2_mux2_1 _1706_ (.A0(net653),
    .A1(\cellsbuf_[155].A ),
    .S(net248),
    .X(_0344_));
 sg13g2_mux2_1 _1707_ (.A0(net864),
    .A1(\cellsbuf_[156].A ),
    .S(net248),
    .X(_0345_));
 sg13g2_mux2_1 _1708_ (.A0(net903),
    .A1(\cellsbuf_[157].A ),
    .S(net250),
    .X(_0346_));
 sg13g2_mux2_1 _1709_ (.A0(\cellsbuf_[158].A ),
    .A1(net933),
    .S(_0506_),
    .X(_0347_));
 sg13g2_mux2_1 _1710_ (.A0(net950),
    .A1(net943),
    .S(net250),
    .X(_0348_));
 sg13g2_nand2_1 _1711_ (.Y(_0389_),
    .A(net916),
    .B(net218));
 sg13g2_mux2_1 _1712_ (.A0(_0529_),
    .A1(net798),
    .S(_0389_),
    .X(_0349_));
 sg13g2_o21ai_1 _1713_ (.B1(net253),
    .Y(_0390_),
    .A1(\row_count[0] ),
    .A2(net220));
 sg13g2_a21oi_1 _1714_ (.A1(_0437_),
    .A2(net220),
    .Y(_0350_),
    .B1(_0390_));
 sg13g2_a21oi_1 _1715_ (.A1(\row_count[0] ),
    .A2(_0462_),
    .Y(_0391_),
    .B1(net935));
 sg13g2_and3_1 _1716_ (.X(_0392_),
    .A(net935),
    .B(\row_count[0] ),
    .C(_0462_));
 sg13g2_nor3_1 _1717_ (.A(_0441_),
    .B(net936),
    .C(_0392_),
    .Y(_0351_));
 sg13g2_o21ai_1 _1718_ (.B1(net253),
    .Y(_0393_),
    .A1(net931),
    .A2(_0392_));
 sg13g2_a21oi_1 _1719_ (.A1(net931),
    .A2(_0392_),
    .Y(_0352_),
    .B1(_0393_));
 sg13g2_mux2_1 _1720_ (.A0(\row_count[3] ),
    .A1(_0011_),
    .S(_0457_),
    .X(_0394_));
 sg13g2_o21ai_1 _1721_ (.B1(net254),
    .Y(_0395_),
    .A1(net965),
    .A2(net220));
 sg13g2_xnor2_1 _1722_ (.Y(_0396_),
    .A(_0466_),
    .B(_0394_));
 sg13g2_a21oi_1 _1723_ (.A1(net220),
    .A2(_0396_),
    .Y(_0353_),
    .B1(_0395_));
 sg13g2_nand2_1 _1724_ (.Y(_0397_),
    .A(_0457_),
    .B(_0468_));
 sg13g2_o21ai_1 _1725_ (.B1(_0397_),
    .Y(_0398_),
    .A1(_0457_),
    .A2(_0474_));
 sg13g2_xor2_1 _1726_ (.B(_0398_),
    .A(net910),
    .X(_0399_));
 sg13g2_o21ai_1 _1727_ (.B1(net254),
    .Y(_0400_),
    .A1(\row_count[4] ),
    .A2(net220));
 sg13g2_a21oi_1 _1728_ (.A1(net220),
    .A2(_0399_),
    .Y(_0354_),
    .B1(_0400_));
 sg13g2_and2_1 _1729_ (.A(\row_count[4] ),
    .B(_0462_),
    .X(_0401_));
 sg13g2_a21oi_1 _1730_ (.A1(_0398_),
    .A2(_0401_),
    .Y(_0402_),
    .B1(net929));
 sg13g2_and4_1 _1731_ (.A(net929),
    .B(\row_count[4] ),
    .C(_0462_),
    .D(_0398_),
    .X(_0403_));
 sg13g2_nor3_1 _1732_ (.A(net251),
    .B(net930),
    .C(_0403_),
    .Y(_0355_));
 sg13g2_o21ai_1 _1733_ (.B1(net254),
    .Y(_0404_),
    .A1(net924),
    .A2(_0403_));
 sg13g2_a21oi_1 _1734_ (.A1(net924),
    .A2(_0403_),
    .Y(_0356_),
    .B1(_0404_));
 sg13g2_o21ai_1 _1735_ (.B1(net254),
    .Y(_0405_),
    .A1(net963),
    .A2(net220));
 sg13g2_nand3_1 _1736_ (.B(_0468_),
    .C(_0469_),
    .A(_0010_),
    .Y(_0406_));
 sg13g2_a21oi_1 _1737_ (.A1(_0468_),
    .A2(_0469_),
    .Y(_0407_),
    .B1(_0010_));
 sg13g2_nor2_1 _1738_ (.A(_0456_),
    .B(_0407_),
    .Y(_0408_));
 sg13g2_o21ai_1 _1739_ (.B1(_0436_),
    .Y(_0409_),
    .A1(_0470_),
    .A2(_0474_));
 sg13g2_a22oi_1 _1740_ (.Y(_0410_),
    .B1(_0409_),
    .B2(_0491_),
    .A2(_0408_),
    .A1(_0406_));
 sg13g2_a21oi_1 _1741_ (.A1(net220),
    .A2(_0410_),
    .Y(_0357_),
    .B1(_0405_));
 sg13g2_nand3_1 _1742_ (.B(_0457_),
    .C(_0461_),
    .A(net945),
    .Y(_0411_));
 sg13g2_a21oi_1 _1743_ (.A1(_0495_),
    .A2(_0411_),
    .Y(_0358_),
    .B1(net251));
 sg13g2_nand3_1 _1744_ (.B(_0457_),
    .C(_0461_),
    .A(net941),
    .Y(_0412_));
 sg13g2_a21oi_1 _1745_ (.A1(_0479_),
    .A2(_0412_),
    .Y(_0359_),
    .B1(net251));
 sg13g2_nand3_1 _1746_ (.B(_0457_),
    .C(_0461_),
    .A(net922),
    .Y(_0413_));
 sg13g2_a21oi_1 _1747_ (.A1(_0486_),
    .A2(_0413_),
    .Y(_0360_),
    .B1(net251));
 sg13g2_nand4_1 _1748_ (.B(\hvsync_gen.vpos[2] ),
    .C(\hvsync_gen.vpos[3] ),
    .A(\hvsync_gen.vpos[9] ),
    .Y(_0414_),
    .D(_0458_));
 sg13g2_o21ai_1 _1749_ (.B1(net254),
    .Y(_0415_),
    .A1(_0515_),
    .A2(_0414_));
 sg13g2_or4_1 _1750_ (.A(_0434_),
    .B(_0373_),
    .C(_0375_),
    .D(_0415_),
    .X(_0416_));
 sg13g2_o21ai_1 _1751_ (.B1(net918),
    .Y(_0361_),
    .A1(_0438_),
    .A2(net221));
 sg13g2_nor3_1 _1752_ (.A(net251),
    .B(_0455_),
    .C(_0458_),
    .Y(_0417_));
 sg13g2_mux2_1 _1753_ (.A0(net845),
    .A1(_0417_),
    .S(net221),
    .X(_0362_));
 sg13g2_nand3_1 _1754_ (.B(_0455_),
    .C(net221),
    .A(net916),
    .Y(_0418_));
 sg13g2_and2_2 _1755_ (.A(net221),
    .B(_0415_),
    .X(_0419_));
 sg13g2_a21oi_1 _1756_ (.A1(_0455_),
    .A2(net221),
    .Y(_0420_),
    .B1(net916));
 sg13g2_nor2_1 _1757_ (.A(_0419_),
    .B(_0420_),
    .Y(_0421_));
 sg13g2_and2_1 _1758_ (.A(_0418_),
    .B(_0421_),
    .X(_0363_));
 sg13g2_nor2b_1 _1759_ (.A(net953),
    .B_N(_0418_),
    .Y(_0422_));
 sg13g2_and4_2 _1760_ (.A(\hvsync_gen.vpos[2] ),
    .B(net953),
    .C(_0455_),
    .D(net221),
    .X(_0423_));
 sg13g2_nor3_1 _1761_ (.A(_0419_),
    .B(_0422_),
    .C(_0423_),
    .Y(_0364_));
 sg13g2_xnor2_1 _1762_ (.Y(_0424_),
    .A(net960),
    .B(_0423_));
 sg13g2_nor2_1 _1763_ (.A(_0419_),
    .B(net961),
    .Y(_0365_));
 sg13g2_a21oi_1 _1764_ (.A1(\hvsync_gen.vpos[4] ),
    .A2(_0423_),
    .Y(_0425_),
    .B1(net920));
 sg13g2_and3_1 _1765_ (.X(_0426_),
    .A(net920),
    .B(net974),
    .C(_0423_));
 sg13g2_nor3_1 _1766_ (.A(_0419_),
    .B(net921),
    .C(_0426_),
    .Y(_0366_));
 sg13g2_xnor2_1 _1767_ (.Y(_0427_),
    .A(net954),
    .B(_0426_));
 sg13g2_nor2_1 _1768_ (.A(_0419_),
    .B(_0427_),
    .Y(_0367_));
 sg13g2_a21oi_1 _1769_ (.A1(\hvsync_gen.vpos[6] ),
    .A2(_0426_),
    .Y(_0428_),
    .B1(net926));
 sg13g2_and3_1 _1770_ (.X(_0429_),
    .A(net926),
    .B(\hvsync_gen.vpos[6] ),
    .C(_0426_));
 sg13g2_nor3_1 _1771_ (.A(_0419_),
    .B(net927),
    .C(_0429_),
    .Y(_0368_));
 sg13g2_a21oi_1 _1772_ (.A1(net947),
    .A2(_0429_),
    .Y(_0430_),
    .B1(_0419_));
 sg13g2_o21ai_1 _1773_ (.B1(_0430_),
    .Y(_0431_),
    .A1(net947),
    .A2(_0429_));
 sg13g2_inv_1 _1774_ (.Y(_0369_),
    .A(_0431_));
 sg13g2_nand2_1 _1775_ (.Y(_0432_),
    .A(\hvsync_gen.vpos[9] ),
    .B(_0430_));
 sg13g2_nand3_1 _1776_ (.B(net254),
    .C(_0429_),
    .A(net947),
    .Y(_0433_));
 sg13g2_o21ai_1 _1777_ (.B1(_0432_),
    .Y(_0370_),
    .A1(\hvsync_gen.vpos[9] ),
    .A2(net948));
 sg13g2_dfrbp_1 _1778_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net421),
    .D(_0018_),
    .Q_N(_0877_),
    .Q(\rule[7] ));
 sg13g2_dfrbp_1 _1779_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net99),
    .D(net944),
    .Q_N(_0876_),
    .Q(left));
 sg13g2_dfrbp_1 _1780_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net98),
    .D(_0020_),
    .Q_N(_0875_),
    .Q(\cellsbuf_[0].A ));
 sg13g2_dfrbp_1 _1781_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net96),
    .D(_0021_),
    .Q_N(_0874_),
    .Q(\next_cellsbuf_[1].A ));
 sg13g2_dfrbp_1 _1782_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net95),
    .D(net602),
    .Q_N(_0873_),
    .Q(\next_cellsbuf_[2].A ));
 sg13g2_dfrbp_1 _1783_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net94),
    .D(net619),
    .Q_N(_0872_),
    .Q(\next_cellsbuf_[3].A ));
 sg13g2_dfrbp_1 _1784_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net93),
    .D(_0024_),
    .Q_N(_0871_),
    .Q(\next_cellsbuf_[4].A ));
 sg13g2_dfrbp_1 _1785_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net92),
    .D(net635),
    .Q_N(_0870_),
    .Q(\next_cellsbuf_[5].A ));
 sg13g2_dfrbp_1 _1786_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net91),
    .D(_0026_),
    .Q_N(_0869_),
    .Q(\next_cellsbuf_[6].A ));
 sg13g2_dfrbp_1 _1787_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net90),
    .D(net526),
    .Q_N(_0868_),
    .Q(\next_cellsbuf_[7].A ));
 sg13g2_dfrbp_1 _1788_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net89),
    .D(net789),
    .Q_N(_0867_),
    .Q(\next_cellsbuf_[8].A ));
 sg13g2_dfrbp_1 _1789_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net88),
    .D(_0029_),
    .Q_N(_0866_),
    .Q(\next_cellsbuf_[9].A ));
 sg13g2_dfrbp_1 _1790_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net87),
    .D(net775),
    .Q_N(_0865_),
    .Q(\next_cellsbuf_[10].A ));
 sg13g2_dfrbp_1 _1791_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net86),
    .D(net604),
    .Q_N(_0864_),
    .Q(\next_cellsbuf_[11].A ));
 sg13g2_dfrbp_1 _1792_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net85),
    .D(_0032_),
    .Q_N(_0863_),
    .Q(\next_cellsbuf_[12].A ));
 sg13g2_dfrbp_1 _1793_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net84),
    .D(_0033_),
    .Q_N(_0862_),
    .Q(\next_cellsbuf_[13].A ));
 sg13g2_dfrbp_1 _1794_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net83),
    .D(_0034_),
    .Q_N(_0861_),
    .Q(\next_cellsbuf_[14].A ));
 sg13g2_dfrbp_1 _1795_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net82),
    .D(net886),
    .Q_N(_0860_),
    .Q(\next_cellsbuf_[15].A ));
 sg13g2_dfrbp_1 _1796_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net81),
    .D(net855),
    .Q_N(_0859_),
    .Q(\next_cellsbuf_[16].A ));
 sg13g2_dfrbp_1 _1797_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net80),
    .D(_0037_),
    .Q_N(_0858_),
    .Q(\next_cellsbuf_[17].A ));
 sg13g2_dfrbp_1 _1798_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net79),
    .D(net721),
    .Q_N(_0857_),
    .Q(\next_cellsbuf_[18].A ));
 sg13g2_dfrbp_1 _1799_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net78),
    .D(net615),
    .Q_N(_0856_),
    .Q(\next_cellsbuf_[19].A ));
 sg13g2_dfrbp_1 _1800_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net77),
    .D(net509),
    .Q_N(_0855_),
    .Q(\next_cellsbuf_[20].A ));
 sg13g2_dfrbp_1 _1801_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net76),
    .D(_0041_),
    .Q_N(_0854_),
    .Q(\next_cellsbuf_[21].A ));
 sg13g2_dfrbp_1 _1802_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net75),
    .D(net705),
    .Q_N(_0853_),
    .Q(\next_cellsbuf_[22].A ));
 sg13g2_dfrbp_1 _1803_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net74),
    .D(_0043_),
    .Q_N(_0852_),
    .Q(\next_cellsbuf_[23].A ));
 sg13g2_dfrbp_1 _1804_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net73),
    .D(net488),
    .Q_N(_0851_),
    .Q(\next_cellsbuf_[24].A ));
 sg13g2_dfrbp_1 _1805_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net72),
    .D(_0045_),
    .Q_N(_0850_),
    .Q(\next_cellsbuf_[25].A ));
 sg13g2_dfrbp_1 _1806_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net71),
    .D(_0046_),
    .Q_N(_0849_),
    .Q(\next_cellsbuf_[26].A ));
 sg13g2_dfrbp_1 _1807_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net70),
    .D(net592),
    .Q_N(_0848_),
    .Q(\next_cellsbuf_[27].A ));
 sg13g2_dfrbp_1 _1808_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net69),
    .D(_0048_),
    .Q_N(_0847_),
    .Q(\next_cellsbuf_[28].A ));
 sg13g2_dfrbp_1 _1809_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net68),
    .D(net596),
    .Q_N(_0846_),
    .Q(\next_cellsbuf_[29].A ));
 sg13g2_dfrbp_1 _1810_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net67),
    .D(_0050_),
    .Q_N(_0845_),
    .Q(\next_cellsbuf_[30].A ));
 sg13g2_dfrbp_1 _1811_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net66),
    .D(net588),
    .Q_N(_0844_),
    .Q(\next_cellsbuf_[31].A ));
 sg13g2_dfrbp_1 _1812_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net65),
    .D(_0052_),
    .Q_N(_0843_),
    .Q(\next_cellsbuf_[32].A ));
 sg13g2_dfrbp_1 _1813_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net64),
    .D(_0053_),
    .Q_N(_0842_),
    .Q(\next_cellsbuf_[33].A ));
 sg13g2_dfrbp_1 _1814_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net63),
    .D(net568),
    .Q_N(_0841_),
    .Q(\next_cellsbuf_[34].A ));
 sg13g2_dfrbp_1 _1815_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net62),
    .D(_0055_),
    .Q_N(_0840_),
    .Q(\next_cellsbuf_[35].A ));
 sg13g2_dfrbp_1 _1816_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net61),
    .D(net814),
    .Q_N(_0839_),
    .Q(\next_cellsbuf_[36].A ));
 sg13g2_dfrbp_1 _1817_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net60),
    .D(net809),
    .Q_N(_0838_),
    .Q(\next_cellsbuf_[37].A ));
 sg13g2_dfrbp_1 _1818_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net59),
    .D(net566),
    .Q_N(_0837_),
    .Q(\next_cellsbuf_[38].A ));
 sg13g2_dfrbp_1 _1819_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net58),
    .D(_0059_),
    .Q_N(_0836_),
    .Q(\next_cellsbuf_[39].A ));
 sg13g2_dfrbp_1 _1820_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net57),
    .D(net500),
    .Q_N(_0835_),
    .Q(\next_cellsbuf_[40].A ));
 sg13g2_dfrbp_1 _1821_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net56),
    .D(_0061_),
    .Q_N(_0834_),
    .Q(\next_cellsbuf_[41].A ));
 sg13g2_dfrbp_1 _1822_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net55),
    .D(_0062_),
    .Q_N(_0833_),
    .Q(\next_cellsbuf_[42].A ));
 sg13g2_dfrbp_1 _1823_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net54),
    .D(_0063_),
    .Q_N(_0832_),
    .Q(\next_cellsbuf_[43].A ));
 sg13g2_dfrbp_1 _1824_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net53),
    .D(net539),
    .Q_N(_0831_),
    .Q(\next_cellsbuf_[44].A ));
 sg13g2_dfrbp_1 _1825_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net52),
    .D(net858),
    .Q_N(_0830_),
    .Q(\next_cellsbuf_[45].A ));
 sg13g2_dfrbp_1 _1826_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net51),
    .D(net818),
    .Q_N(_0829_),
    .Q(\next_cellsbuf_[46].A ));
 sg13g2_dfrbp_1 _1827_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net50),
    .D(net710),
    .Q_N(_0828_),
    .Q(\next_cellsbuf_[47].A ));
 sg13g2_dfrbp_1 _1828_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net49),
    .D(_0068_),
    .Q_N(_0827_),
    .Q(\next_cellsbuf_[48].A ));
 sg13g2_dfrbp_1 _1829_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net48),
    .D(net641),
    .Q_N(_0826_),
    .Q(\next_cellsbuf_[49].A ));
 sg13g2_dfrbp_1 _1830_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net47),
    .D(_0070_),
    .Q_N(_0825_),
    .Q(\next_cellsbuf_[50].A ));
 sg13g2_dfrbp_1 _1831_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net46),
    .D(_0071_),
    .Q_N(_0824_),
    .Q(\next_cellsbuf_[51].A ));
 sg13g2_dfrbp_1 _1832_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net45),
    .D(net650),
    .Q_N(_0823_),
    .Q(\next_cellsbuf_[52].A ));
 sg13g2_dfrbp_1 _1833_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net44),
    .D(_0073_),
    .Q_N(_0822_),
    .Q(\next_cellsbuf_[53].A ));
 sg13g2_dfrbp_1 _1834_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net43),
    .D(net729),
    .Q_N(_0821_),
    .Q(\next_cellsbuf_[54].A ));
 sg13g2_dfrbp_1 _1835_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net42),
    .D(_0075_),
    .Q_N(_0820_),
    .Q(\next_cellsbuf_[55].A ));
 sg13g2_dfrbp_1 _1836_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net41),
    .D(net656),
    .Q_N(_0819_),
    .Q(\next_cellsbuf_[56].A ));
 sg13g2_dfrbp_1 _1837_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net40),
    .D(_0077_),
    .Q_N(_0818_),
    .Q(\next_cellsbuf_[57].A ));
 sg13g2_dfrbp_1 _1838_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net39),
    .D(_0078_),
    .Q_N(_0817_),
    .Q(\next_cellsbuf_[58].A ));
 sg13g2_dfrbp_1 _1839_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net38),
    .D(_0079_),
    .Q_N(_0816_),
    .Q(\next_cellsbuf_[59].A ));
 sg13g2_dfrbp_1 _1840_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net37),
    .D(net745),
    .Q_N(_0815_),
    .Q(\next_cellsbuf_[60].A ));
 sg13g2_dfrbp_1 _1841_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net36),
    .D(net703),
    .Q_N(_0814_),
    .Q(\next_cellsbuf_[61].A ));
 sg13g2_dfrbp_1 _1842_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net35),
    .D(_0082_),
    .Q_N(_0813_),
    .Q(\next_cellsbuf_[62].A ));
 sg13g2_dfrbp_1 _1843_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net34),
    .D(net658),
    .Q_N(_0812_),
    .Q(\next_cellsbuf_[63].A ));
 sg13g2_dfrbp_1 _1844_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net33),
    .D(_0084_),
    .Q_N(_0811_),
    .Q(\next_cellsbuf_[64].A ));
 sg13g2_dfrbp_1 _1845_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net32),
    .D(_0085_),
    .Q_N(_0810_),
    .Q(\next_cellsbuf_[65].A ));
 sg13g2_dfrbp_1 _1846_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net31),
    .D(net460),
    .Q_N(_0809_),
    .Q(\next_cellsbuf_[66].A ));
 sg13g2_dfrbp_1 _1847_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net30),
    .D(net529),
    .Q_N(_0808_),
    .Q(\next_cellsbuf_[67].A ));
 sg13g2_dfrbp_1 _1848_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net29),
    .D(_0088_),
    .Q_N(_0807_),
    .Q(\next_cellsbuf_[68].A ));
 sg13g2_dfrbp_1 _1849_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net28),
    .D(net834),
    .Q_N(_0806_),
    .Q(\next_cellsbuf_[69].A ));
 sg13g2_dfrbp_1 _1850_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net27),
    .D(net718),
    .Q_N(_0805_),
    .Q(\next_cellsbuf_[70].A ));
 sg13g2_dfrbp_1 _1851_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net26),
    .D(_0091_),
    .Q_N(_0804_),
    .Q(\next_cellsbuf_[71].A ));
 sg13g2_dfrbp_1 _1852_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net25),
    .D(_0092_),
    .Q_N(_0803_),
    .Q(\next_cellsbuf_[72].A ));
 sg13g2_dfrbp_1 _1853_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net24),
    .D(net757),
    .Q_N(_0802_),
    .Q(\next_cellsbuf_[73].A ));
 sg13g2_dfrbp_1 _1854_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net23),
    .D(net550),
    .Q_N(_0801_),
    .Q(\next_cellsbuf_[74].A ));
 sg13g2_dfrbp_1 _1855_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net22),
    .D(_0095_),
    .Q_N(_0800_),
    .Q(\next_cellsbuf_[75].A ));
 sg13g2_dfrbp_1 _1856_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net21),
    .D(net582),
    .Q_N(_0799_),
    .Q(\next_cellsbuf_[76].A ));
 sg13g2_dfrbp_1 _1857_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net20),
    .D(net532),
    .Q_N(_0798_),
    .Q(\next_cellsbuf_[77].A ));
 sg13g2_dfrbp_1 _1858_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net19),
    .D(_0098_),
    .Q_N(_0797_),
    .Q(\next_cellsbuf_[78].A ));
 sg13g2_dfrbp_1 _1859_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net18),
    .D(net676),
    .Q_N(_0796_),
    .Q(\next_cellsbuf_[79].A ));
 sg13g2_dfrbp_1 _1860_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net17),
    .D(_0100_),
    .Q_N(_0795_),
    .Q(\next_cellsbuf_[80].A ));
 sg13g2_dfrbp_1 _1861_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net438),
    .D(net684),
    .Q_N(_0794_),
    .Q(\next_cellsbuf_[81].A ));
 sg13g2_dfrbp_1 _1862_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net437),
    .D(_0102_),
    .Q_N(_0793_),
    .Q(\next_cellsbuf_[82].A ));
 sg13g2_dfrbp_1 _1863_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net436),
    .D(net648),
    .Q_N(_0792_),
    .Q(\next_cellsbuf_[83].A ));
 sg13g2_dfrbp_1 _1864_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net435),
    .D(_0104_),
    .Q_N(_0791_),
    .Q(\next_cellsbuf_[84].A ));
 sg13g2_dfrbp_1 _1865_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net434),
    .D(net696),
    .Q_N(_0790_),
    .Q(\next_cellsbuf_[85].A ));
 sg13g2_dfrbp_1 _1866_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net433),
    .D(net672),
    .Q_N(_0789_),
    .Q(\next_cellsbuf_[86].A ));
 sg13g2_dfrbp_1 _1867_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net432),
    .D(_0107_),
    .Q_N(_0788_),
    .Q(\next_cellsbuf_[87].A ));
 sg13g2_dfrbp_1 _1868_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net431),
    .D(_0108_),
    .Q_N(_0787_),
    .Q(\next_cellsbuf_[88].A ));
 sg13g2_dfrbp_1 _1869_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net430),
    .D(_0109_),
    .Q_N(_0786_),
    .Q(\next_cellsbuf_[89].A ));
 sg13g2_dfrbp_1 _1870_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net429),
    .D(_0110_),
    .Q_N(_0785_),
    .Q(\next_cellsbuf_[90].A ));
 sg13g2_dfrbp_1 _1871_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net420),
    .D(net759),
    .Q_N(_0784_),
    .Q(\next_cellsbuf_[91].A ));
 sg13g2_dfrbp_1 _1872_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net419),
    .D(_0112_),
    .Q_N(_0783_),
    .Q(\next_cellsbuf_[92].A ));
 sg13g2_dfrbp_1 _1873_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net418),
    .D(_0113_),
    .Q_N(_0782_),
    .Q(\next_cellsbuf_[93].A ));
 sg13g2_dfrbp_1 _1874_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net417),
    .D(net643),
    .Q_N(_0781_),
    .Q(\next_cellsbuf_[94].A ));
 sg13g2_dfrbp_1 _1875_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net416),
    .D(_0115_),
    .Q_N(_0780_),
    .Q(\next_cellsbuf_[95].A ));
 sg13g2_dfrbp_1 _1876_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net415),
    .D(_0116_),
    .Q_N(_0779_),
    .Q(\next_cellsbuf_[96].A ));
 sg13g2_dfrbp_1 _1877_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net414),
    .D(net825),
    .Q_N(_0778_),
    .Q(\next_cellsbuf_[97].A ));
 sg13g2_dfrbp_1 _1878_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net413),
    .D(_0118_),
    .Q_N(_0777_),
    .Q(\next_cellsbuf_[98].A ));
 sg13g2_dfrbp_1 _1879_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net412),
    .D(net726),
    .Q_N(_0776_),
    .Q(\next_cellsbuf_[99].A ));
 sg13g2_dfrbp_1 _1880_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net411),
    .D(net560),
    .Q_N(_0775_),
    .Q(\next_cellsbuf_[100].A ));
 sg13g2_dfrbp_1 _1881_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net410),
    .D(_0121_),
    .Q_N(_0774_),
    .Q(\next_cellsbuf_[101].A ));
 sg13g2_dfrbp_1 _1882_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net409),
    .D(net574),
    .Q_N(_0773_),
    .Q(\next_cellsbuf_[102].A ));
 sg13g2_dfrbp_1 _1883_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net408),
    .D(net511),
    .Q_N(_0772_),
    .Q(\next_cellsbuf_[103].A ));
 sg13g2_dfrbp_1 _1884_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net407),
    .D(_0124_),
    .Q_N(_0771_),
    .Q(\next_cellsbuf_[104].A ));
 sg13g2_dfrbp_1 _1885_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net406),
    .D(_0125_),
    .Q_N(_0770_),
    .Q(\next_cellsbuf_[105].A ));
 sg13g2_dfrbp_1 _1886_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net405),
    .D(net778),
    .Q_N(_0769_),
    .Q(\next_cellsbuf_[106].A ));
 sg13g2_dfrbp_1 _1887_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net404),
    .D(net669),
    .Q_N(_0768_),
    .Q(\next_cellsbuf_[107].A ));
 sg13g2_dfrbp_1 _1888_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net403),
    .D(net516),
    .Q_N(_0767_),
    .Q(\next_cellsbuf_[108].A ));
 sg13g2_dfrbp_1 _1889_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net402),
    .D(_0129_),
    .Q_N(_0766_),
    .Q(\next_cellsbuf_[109].A ));
 sg13g2_dfrbp_1 _1890_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net401),
    .D(_0130_),
    .Q_N(_0765_),
    .Q(\next_cellsbuf_[110].A ));
 sg13g2_dfrbp_1 _1891_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net400),
    .D(net454),
    .Q_N(_0764_),
    .Q(\next_cellsbuf_[111].A ));
 sg13g2_dfrbp_1 _1892_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net399),
    .D(net692),
    .Q_N(_0763_),
    .Q(\next_cellsbuf_[112].A ));
 sg13g2_dfrbp_1 _1893_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net398),
    .D(net486),
    .Q_N(_0762_),
    .Q(\next_cellsbuf_[113].A ));
 sg13g2_dfrbp_1 _1894_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net397),
    .D(_0134_),
    .Q_N(_0761_),
    .Q(\next_cellsbuf_[114].A ));
 sg13g2_dfrbp_1 _1895_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net396),
    .D(net507),
    .Q_N(_0760_),
    .Q(\next_cellsbuf_[115].A ));
 sg13g2_dfrbp_1 _1896_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net395),
    .D(_0136_),
    .Q_N(_0759_),
    .Q(\next_cellsbuf_[116].A ));
 sg13g2_dfrbp_1 _1897_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net394),
    .D(_0137_),
    .Q_N(_0758_),
    .Q(\next_cellsbuf_[117].A ));
 sg13g2_dfrbp_1 _1898_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net393),
    .D(_0138_),
    .Q_N(_0757_),
    .Q(\next_cellsbuf_[118].A ));
 sg13g2_dfrbp_1 _1899_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net392),
    .D(net608),
    .Q_N(_0756_),
    .Q(\next_cellsbuf_[119].A ));
 sg13g2_dfrbp_1 _1900_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net391),
    .D(_0140_),
    .Q_N(_0755_),
    .Q(\next_cellsbuf_[120].A ));
 sg13g2_dfrbp_1 _1901_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net390),
    .D(_0141_),
    .Q_N(_0754_),
    .Q(\next_cellsbuf_[121].A ));
 sg13g2_dfrbp_1 _1902_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net389),
    .D(net633),
    .Q_N(_0753_),
    .Q(\next_cellsbuf_[122].A ));
 sg13g2_dfrbp_1 _1903_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net388),
    .D(_0143_),
    .Q_N(_0752_),
    .Q(\next_cellsbuf_[123].A ));
 sg13g2_dfrbp_1 _1904_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net387),
    .D(net518),
    .Q_N(_0751_),
    .Q(\next_cellsbuf_[124].A ));
 sg13g2_dfrbp_1 _1905_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net386),
    .D(_0145_),
    .Q_N(_0750_),
    .Q(\next_cellsbuf_[125].A ));
 sg13g2_dfrbp_1 _1906_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net385),
    .D(_0146_),
    .Q_N(_0749_),
    .Q(\next_cellsbuf_[126].A ));
 sg13g2_dfrbp_1 _1907_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net384),
    .D(net464),
    .Q_N(_0748_),
    .Q(\next_cellsbuf_[127].A ));
 sg13g2_dfrbp_1 _1908_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net383),
    .D(net623),
    .Q_N(_0747_),
    .Q(\next_cellsbuf_[128].A ));
 sg13g2_dfrbp_1 _1909_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net382),
    .D(_0149_),
    .Q_N(_0746_),
    .Q(\next_cellsbuf_[129].A ));
 sg13g2_dfrbp_1 _1910_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net381),
    .D(net698),
    .Q_N(_0745_),
    .Q(\next_cellsbuf_[130].A ));
 sg13g2_dfrbp_1 _1911_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net380),
    .D(net652),
    .Q_N(_0744_),
    .Q(\next_cellsbuf_[131].A ));
 sg13g2_dfrbp_1 _1912_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net379),
    .D(net625),
    .Q_N(_0743_),
    .Q(\next_cellsbuf_[132].A ));
 sg13g2_dfrbp_1 _1913_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net378),
    .D(net621),
    .Q_N(_0742_),
    .Q(\next_cellsbuf_[133].A ));
 sg13g2_dfrbp_1 _1914_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net377),
    .D(net599),
    .Q_N(_0741_),
    .Q(\next_cellsbuf_[134].A ));
 sg13g2_dfrbp_1 _1915_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net376),
    .D(_0155_),
    .Q_N(_0740_),
    .Q(\next_cellsbuf_[135].A ));
 sg13g2_dfrbp_1 _1916_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net375),
    .D(_0156_),
    .Q_N(_0739_),
    .Q(\next_cellsbuf_[136].A ));
 sg13g2_dfrbp_1 _1917_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net374),
    .D(net504),
    .Q_N(_0738_),
    .Q(\next_cellsbuf_[137].A ));
 sg13g2_dfrbp_1 _1918_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net373),
    .D(net502),
    .Q_N(_0737_),
    .Q(\next_cellsbuf_[138].A ));
 sg13g2_dfrbp_1 _1919_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net372),
    .D(_0159_),
    .Q_N(_0736_),
    .Q(\next_cellsbuf_[139].A ));
 sg13g2_dfrbp_1 _1920_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net371),
    .D(_0160_),
    .Q_N(_0735_),
    .Q(\next_cellsbuf_[140].A ));
 sg13g2_dfrbp_1 _1921_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net370),
    .D(net570),
    .Q_N(_0734_),
    .Q(\next_cellsbuf_[141].A ));
 sg13g2_dfrbp_1 _1922_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net369),
    .D(net812),
    .Q_N(_0733_),
    .Q(\next_cellsbuf_[142].A ));
 sg13g2_dfrbp_1 _1923_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net368),
    .D(net663),
    .Q_N(_0732_),
    .Q(\next_cellsbuf_[143].A ));
 sg13g2_dfrbp_1 _1924_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net367),
    .D(_0164_),
    .Q_N(_0731_),
    .Q(\next_cellsbuf_[144].A ));
 sg13g2_dfrbp_1 _1925_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net366),
    .D(_0165_),
    .Q_N(_0730_),
    .Q(\next_cellsbuf_[145].A ));
 sg13g2_dfrbp_1 _1926_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net365),
    .D(_0166_),
    .Q_N(_0729_),
    .Q(\next_cellsbuf_[146].A ));
 sg13g2_dfrbp_1 _1927_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net364),
    .D(net780),
    .Q_N(_0728_),
    .Q(\next_cellsbuf_[147].A ));
 sg13g2_dfrbp_1 _1928_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net363),
    .D(net585),
    .Q_N(_0727_),
    .Q(\next_cellsbuf_[148].A ));
 sg13g2_dfrbp_1 _1929_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net362),
    .D(_0169_),
    .Q_N(_0726_),
    .Q(\next_cellsbuf_[149].A ));
 sg13g2_dfrbp_1 _1930_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net361),
    .D(net752),
    .Q_N(_0725_),
    .Q(\next_cellsbuf_[150].A ));
 sg13g2_dfrbp_1 _1931_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net360),
    .D(_0171_),
    .Q_N(_0724_),
    .Q(\next_cellsbuf_[151].A ));
 sg13g2_dfrbp_1 _1932_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net359),
    .D(net755),
    .Q_N(_0723_),
    .Q(\next_cellsbuf_[152].A ));
 sg13g2_dfrbp_1 _1933_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net358),
    .D(net714),
    .Q_N(_0722_),
    .Q(\next_cellsbuf_[153].A ));
 sg13g2_dfrbp_1 _1934_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net357),
    .D(net686),
    .Q_N(_0721_),
    .Q(\next_cellsbuf_[154].A ));
 sg13g2_dfrbp_1 _1935_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net356),
    .D(net617),
    .Q_N(_0720_),
    .Q(\next_cellsbuf_[155].A ));
 sg13g2_dfrbp_1 _1936_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net355),
    .D(net590),
    .Q_N(_0719_),
    .Q(\next_cellsbuf_[156].A ));
 sg13g2_dfrbp_1 _1937_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net354),
    .D(net513),
    .Q_N(_0718_),
    .Q(\next_cellsbuf_[157].A ));
 sg13g2_dfrbp_1 _1938_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net353),
    .D(_0178_),
    .Q_N(_0717_),
    .Q(\next_cellsbuf_[158].A ));
 sg13g2_dfrbp_1 _1939_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net352),
    .D(net735),
    .Q_N(_0716_),
    .Q(\next_cellsbuf_[159].A ));
 sg13g2_dfrbp_1 _1940_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net351),
    .D(_0180_),
    .Q_N(_0017_),
    .Q(\fract_x[0] ));
 sg13g2_dfrbp_1 _1941_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net350),
    .D(net971),
    .Q_N(_0715_),
    .Q(\fract_x[1] ));
 sg13g2_dfrbp_1 _1942_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net349),
    .D(_0182_),
    .Q_N(_0714_),
    .Q(\cell_x[0] ));
 sg13g2_dfrbp_1 _1943_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net348),
    .D(_0183_),
    .Q_N(_0713_),
    .Q(\cell_x[1] ));
 sg13g2_dfrbp_1 _1944_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net347),
    .D(net968),
    .Q_N(_0712_),
    .Q(\cell_x[2] ));
 sg13g2_dfrbp_1 _1945_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net346),
    .D(net940),
    .Q_N(_0711_),
    .Q(\cell_x[3] ));
 sg13g2_dfrbp_1 _1946_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net345),
    .D(_0186_),
    .Q_N(_0710_),
    .Q(\cell_x[4] ));
 sg13g2_dfrbp_1 _1947_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net344),
    .D(_0187_),
    .Q_N(_0709_),
    .Q(\cell_x[5] ));
 sg13g2_dfrbp_1 _1948_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net343),
    .D(_0188_),
    .Q_N(_0708_),
    .Q(\cell_x[6] ));
 sg13g2_dfrbp_1 _1949_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net342),
    .D(_0189_),
    .Q_N(_0707_),
    .Q(\cell_x[7] ));
 sg13g2_dfrbp_1 _1950_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net341),
    .D(_0190_),
    .Q_N(_0706_),
    .Q(\cellsbuf_[1].A ));
 sg13g2_dfrbp_1 _1951_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net340),
    .D(net466),
    .Q_N(_0705_),
    .Q(\cellsbuf_[2].A ));
 sg13g2_dfrbp_1 _1952_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net339),
    .D(_0192_),
    .Q_N(_0704_),
    .Q(\cellsbuf_[3].A ));
 sg13g2_dfrbp_1 _1953_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net338),
    .D(_0193_),
    .Q_N(_0703_),
    .Q(\cellsbuf_[4].A ));
 sg13g2_dfrbp_1 _1954_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net337),
    .D(_0194_),
    .Q_N(_0702_),
    .Q(\cellsbuf_[5].A ));
 sg13g2_dfrbp_1 _1955_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net336),
    .D(net645),
    .Q_N(_0701_),
    .Q(\cellsbuf_[6].A ));
 sg13g2_dfrbp_1 _1956_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net335),
    .D(net690),
    .Q_N(_0700_),
    .Q(\cellsbuf_[7].A ));
 sg13g2_dfrbp_1 _1957_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net334),
    .D(_0197_),
    .Q_N(_0699_),
    .Q(\cellsbuf_[8].A ));
 sg13g2_dfrbp_1 _1958_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net333),
    .D(net580),
    .Q_N(_0698_),
    .Q(\cellsbuf_[9].A ));
 sg13g2_dfrbp_1 _1959_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net332),
    .D(_0199_),
    .Q_N(_0697_),
    .Q(\cellsbuf_[10].A ));
 sg13g2_dfrbp_1 _1960_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net331),
    .D(_0200_),
    .Q_N(_0696_),
    .Q(\cellsbuf_[11].A ));
 sg13g2_dfrbp_1 _1961_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net330),
    .D(net490),
    .Q_N(_0695_),
    .Q(\cellsbuf_[12].A ));
 sg13g2_dfrbp_1 _1962_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net329),
    .D(_0202_),
    .Q_N(_0694_),
    .Q(\cellsbuf_[13].A ));
 sg13g2_dfrbp_1 _1963_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net328),
    .D(_0203_),
    .Q_N(_0693_),
    .Q(\cellsbuf_[14].A ));
 sg13g2_dfrbp_1 _1964_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net327),
    .D(net450),
    .Q_N(_0692_),
    .Q(\cellsbuf_[15].A ));
 sg13g2_dfrbp_1 _1965_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net326),
    .D(net852),
    .Q_N(_0691_),
    .Q(\cellsbuf_[16].A ));
 sg13g2_dfrbp_1 _1966_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net325),
    .D(_0206_),
    .Q_N(_0690_),
    .Q(\cellsbuf_[17].A ));
 sg13g2_dfrbp_1 _1967_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net324),
    .D(net474),
    .Q_N(_0689_),
    .Q(\cellsbuf_[18].A ));
 sg13g2_dfrbp_1 _1968_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net323),
    .D(net548),
    .Q_N(_0688_),
    .Q(\cellsbuf_[19].A ));
 sg13g2_dfrbp_1 _1969_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net322),
    .D(net901),
    .Q_N(_0687_),
    .Q(\cellsbuf_[20].A ));
 sg13g2_dfrbp_1 _1970_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net321),
    .D(_0210_),
    .Q_N(_0686_),
    .Q(\cellsbuf_[21].A ));
 sg13g2_dfrbp_1 _1971_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net320),
    .D(net750),
    .Q_N(_0685_),
    .Q(\cellsbuf_[22].A ));
 sg13g2_dfrbp_1 _1972_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net319),
    .D(_0212_),
    .Q_N(_0684_),
    .Q(\cellsbuf_[23].A ));
 sg13g2_dfrbp_1 _1973_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net318),
    .D(net871),
    .Q_N(_0683_),
    .Q(\cellsbuf_[24].A ));
 sg13g2_dfrbp_1 _1974_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net317),
    .D(_0214_),
    .Q_N(_0682_),
    .Q(\cellsbuf_[25].A ));
 sg13g2_dfrbp_1 _1975_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net316),
    .D(net631),
    .Q_N(_0681_),
    .Q(\cellsbuf_[26].A ));
 sg13g2_dfrbp_1 _1976_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net315),
    .D(_0216_),
    .Q_N(_0680_),
    .Q(\cellsbuf_[27].A ));
 sg13g2_dfrbp_1 _1977_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net314),
    .D(net553),
    .Q_N(_0679_),
    .Q(\cellsbuf_[28].A ));
 sg13g2_dfrbp_1 _1978_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net313),
    .D(_0218_),
    .Q_N(_0678_),
    .Q(\cellsbuf_[29].A ));
 sg13g2_dfrbp_1 _1979_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net312),
    .D(_0219_),
    .Q_N(_0677_),
    .Q(\cellsbuf_[30].A ));
 sg13g2_dfrbp_1 _1980_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net311),
    .D(net712),
    .Q_N(_0676_),
    .Q(\cellsbuf_[31].A ));
 sg13g2_dfrbp_1 _1981_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net310),
    .D(_0221_),
    .Q_N(_0675_),
    .Q(\cellsbuf_[32].A ));
 sg13g2_dfrbp_1 _1982_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net309),
    .D(net524),
    .Q_N(_0674_),
    .Q(\cellsbuf_[33].A ));
 sg13g2_dfrbp_1 _1983_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net308),
    .D(net562),
    .Q_N(_0673_),
    .Q(\cellsbuf_[34].A ));
 sg13g2_dfrbp_1 _1984_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net307),
    .D(net732),
    .Q_N(_0672_),
    .Q(\cellsbuf_[35].A ));
 sg13g2_dfrbp_1 _1985_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net306),
    .D(_0225_),
    .Q_N(_0671_),
    .Q(\cellsbuf_[36].A ));
 sg13g2_dfrbp_1 _1986_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net305),
    .D(net494),
    .Q_N(_0670_),
    .Q(\cellsbuf_[37].A ));
 sg13g2_dfrbp_1 _1987_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net304),
    .D(_0227_),
    .Q_N(_0669_),
    .Q(\cellsbuf_[38].A ));
 sg13g2_dfrbp_1 _1988_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net303),
    .D(net456),
    .Q_N(_0668_),
    .Q(\cellsbuf_[39].A ));
 sg13g2_dfrbp_1 _1989_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net302),
    .D(_0229_),
    .Q_N(_0667_),
    .Q(\cellsbuf_[40].A ));
 sg13g2_dfrbp_1 _1990_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net301),
    .D(net861),
    .Q_N(_0666_),
    .Q(\cellsbuf_[41].A ));
 sg13g2_dfrbp_1 _1991_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net300),
    .D(_0231_),
    .Q_N(_0665_),
    .Q(\cellsbuf_[42].A ));
 sg13g2_dfrbp_1 _1992_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net299),
    .D(_0232_),
    .Q_N(_0664_),
    .Q(\cellsbuf_[43].A ));
 sg13g2_dfrbp_1 _1993_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net298),
    .D(net468),
    .Q_N(_0663_),
    .Q(\cellsbuf_[44].A ));
 sg13g2_dfrbp_1 _1994_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net297),
    .D(_0234_),
    .Q_N(_0662_),
    .Q(\cellsbuf_[45].A ));
 sg13g2_dfrbp_1 _1995_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net296),
    .D(_0235_),
    .Q_N(_0661_),
    .Q(\cellsbuf_[46].A ));
 sg13g2_dfrbp_1 _1996_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net295),
    .D(net556),
    .Q_N(_0660_),
    .Q(\cellsbuf_[47].A ));
 sg13g2_dfrbp_1 _1997_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net294),
    .D(_0237_),
    .Q_N(_0659_),
    .Q(\cellsbuf_[48].A ));
 sg13g2_dfrbp_1 _1998_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net293),
    .D(_0238_),
    .Q_N(_0658_),
    .Q(\cellsbuf_[49].A ));
 sg13g2_dfrbp_1 _1999_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net292),
    .D(net498),
    .Q_N(_0657_),
    .Q(\cellsbuf_[50].A ));
 sg13g2_dfrbp_1 _2000_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net291),
    .D(net783),
    .Q_N(_0656_),
    .Q(\cellsbuf_[51].A ));
 sg13g2_dfrbp_1 _2001_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net290),
    .D(_0241_),
    .Q_N(_0655_),
    .Q(\cellsbuf_[52].A ));
 sg13g2_dfrbp_1 _2002_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net289),
    .D(net610),
    .Q_N(_0654_),
    .Q(\cellsbuf_[53].A ));
 sg13g2_dfrbp_1 _2003_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net288),
    .D(_0243_),
    .Q_N(_0653_),
    .Q(\cellsbuf_[54].A ));
 sg13g2_dfrbp_1 _2004_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net287),
    .D(_0244_),
    .Q_N(_0652_),
    .Q(\cellsbuf_[55].A ));
 sg13g2_dfrbp_1 _2005_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net286),
    .D(_0245_),
    .Q_N(_0651_),
    .Q(\cellsbuf_[56].A ));
 sg13g2_dfrbp_1 _2006_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net285),
    .D(net462),
    .Q_N(_0650_),
    .Q(\cellsbuf_[57].A ));
 sg13g2_dfrbp_1 _2007_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net284),
    .D(_0247_),
    .Q_N(_0649_),
    .Q(\cellsbuf_[58].A ));
 sg13g2_dfrbp_1 _2008_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net283),
    .D(net482),
    .Q_N(_0648_),
    .Q(\cellsbuf_[59].A ));
 sg13g2_dfrbp_1 _2009_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net282),
    .D(_0249_),
    .Q_N(_0647_),
    .Q(\cellsbuf_[60].A ));
 sg13g2_dfrbp_1 _2010_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net281),
    .D(net627),
    .Q_N(_0646_),
    .Q(\cellsbuf_[61].A ));
 sg13g2_dfrbp_1 _2011_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net280),
    .D(net661),
    .Q_N(_0645_),
    .Q(\cellsbuf_[62].A ));
 sg13g2_dfrbp_1 _2012_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net279),
    .D(net868),
    .Q_N(_0644_),
    .Q(\cellsbuf_[63].A ));
 sg13g2_dfrbp_1 _2013_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net278),
    .D(net737),
    .Q_N(_0643_),
    .Q(\cellsbuf_[64].A ));
 sg13g2_dfrbp_1 _2014_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net277),
    .D(_0254_),
    .Q_N(_0642_),
    .Q(\cellsbuf_[65].A ));
 sg13g2_dfrbp_1 _2015_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net276),
    .D(_0255_),
    .Q_N(_0641_),
    .Q(\cellsbuf_[66].A ));
 sg13g2_dfrbp_1 _2016_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net275),
    .D(_0256_),
    .Q_N(_0640_),
    .Q(\cellsbuf_[67].A ));
 sg13g2_dfrbp_1 _2017_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net274),
    .D(net458),
    .Q_N(_0639_),
    .Q(\cellsbuf_[68].A ));
 sg13g2_dfrbp_1 _2018_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net273),
    .D(net786),
    .Q_N(_0638_),
    .Q(\cellsbuf_[69].A ));
 sg13g2_dfrbp_1 _2019_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net272),
    .D(_0259_),
    .Q_N(_0637_),
    .Q(\cellsbuf_[70].A ));
 sg13g2_dfrbp_1 _2020_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net271),
    .D(net558),
    .Q_N(_0636_),
    .Q(\cellsbuf_[71].A ));
 sg13g2_dfrbp_1 _2021_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net270),
    .D(net594),
    .Q_N(_0635_),
    .Q(\cellsbuf_[72].A ));
 sg13g2_dfrbp_1 _2022_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net269),
    .D(_0262_),
    .Q_N(_0634_),
    .Q(\cellsbuf_[73].A ));
 sg13g2_dfrbp_1 _2023_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net268),
    .D(net541),
    .Q_N(_0633_),
    .Q(\cellsbuf_[74].A ));
 sg13g2_dfrbp_1 _2024_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net267),
    .D(net612),
    .Q_N(_0632_),
    .Q(\cellsbuf_[75].A ));
 sg13g2_dfrbp_1 _2025_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net266),
    .D(net821),
    .Q_N(_0631_),
    .Q(\cellsbuf_[76].A ));
 sg13g2_dfrbp_1 _2026_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net265),
    .D(net838),
    .Q_N(_0630_),
    .Q(\cellsbuf_[77].A ));
 sg13g2_dfrbp_1 _2027_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net264),
    .D(_0267_),
    .Q_N(_0629_),
    .Q(\cellsbuf_[78].A ));
 sg13g2_dfrbp_1 _2028_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net263),
    .D(_0268_),
    .Q_N(_0628_),
    .Q(\cellsbuf_[79].A ));
 sg13g2_dfrbp_1 _2029_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net262),
    .D(_0269_),
    .Q_N(_0627_),
    .Q(\cellsbuf_[80].A ));
 sg13g2_dfrbp_1 _2030_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net261),
    .D(net448),
    .Q_N(_0626_),
    .Q(\cellsbuf_[81].A ));
 sg13g2_dfrbp_1 _2031_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net260),
    .D(_0271_),
    .Q_N(_0625_),
    .Q(\cellsbuf_[82].A ));
 sg13g2_dfrbp_1 _2032_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net259),
    .D(net452),
    .Q_N(_0624_),
    .Q(\cellsbuf_[83].A ));
 sg13g2_dfrbp_1 _2033_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net258),
    .D(_0273_),
    .Q_N(_0623_),
    .Q(\cellsbuf_[84].A ));
 sg13g2_dfrbp_1 _2034_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net257),
    .D(_0274_),
    .Q_N(_0622_),
    .Q(\cellsbuf_[85].A ));
 sg13g2_dfrbp_1 _2035_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net256),
    .D(_0275_),
    .Q_N(_0621_),
    .Q(\cellsbuf_[86].A ));
 sg13g2_dfrbp_1 _2036_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net255),
    .D(net520),
    .Q_N(_0620_),
    .Q(\cellsbuf_[87].A ));
 sg13g2_dfrbp_1 _2037_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net193),
    .D(net694),
    .Q_N(_0619_),
    .Q(\cellsbuf_[88].A ));
 sg13g2_dfrbp_1 _2038_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net192),
    .D(_0278_),
    .Q_N(_0618_),
    .Q(\cellsbuf_[89].A ));
 sg13g2_dfrbp_1 _2039_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net191),
    .D(net480),
    .Q_N(_0617_),
    .Q(\cellsbuf_[90].A ));
 sg13g2_dfrbp_1 _2040_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net190),
    .D(_0280_),
    .Q_N(_0616_),
    .Q(\cellsbuf_[91].A ));
 sg13g2_dfrbp_1 _2041_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net189),
    .D(_0281_),
    .Q_N(_0615_),
    .Q(\cellsbuf_[92].A ));
 sg13g2_dfrbp_1 _2042_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net188),
    .D(net578),
    .Q_N(_0614_),
    .Q(\cellsbuf_[93].A ));
 sg13g2_dfrbp_1 _2043_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net187),
    .D(_0283_),
    .Q_N(_0613_),
    .Q(\cellsbuf_[94].A ));
 sg13g2_dfrbp_1 _2044_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net186),
    .D(net534),
    .Q_N(_0612_),
    .Q(\cellsbuf_[95].A ));
 sg13g2_dfrbp_1 _2045_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net185),
    .D(_0285_),
    .Q_N(_0611_),
    .Q(\cellsbuf_[96].A ));
 sg13g2_dfrbp_1 _2046_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net184),
    .D(net772),
    .Q_N(_0610_),
    .Q(\cellsbuf_[97].A ));
 sg13g2_dfrbp_1 _2047_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net183),
    .D(_0287_),
    .Q_N(_0609_),
    .Q(\cellsbuf_[98].A ));
 sg13g2_dfrbp_1 _2048_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net182),
    .D(net496),
    .Q_N(_0608_),
    .Q(\cellsbuf_[99].A ));
 sg13g2_dfrbp_1 _2049_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net181),
    .D(net674),
    .Q_N(_0607_),
    .Q(\cellsbuf_[100].A ));
 sg13g2_dfrbp_1 _2050_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net180),
    .D(_0290_),
    .Q_N(_0606_),
    .Q(\cellsbuf_[101].A ));
 sg13g2_dfrbp_1 _2051_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net179),
    .D(net492),
    .Q_N(_0605_),
    .Q(\cellsbuf_[102].A ));
 sg13g2_dfrbp_1 _2052_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net178),
    .D(_0292_),
    .Q_N(_0604_),
    .Q(\cellsbuf_[103].A ));
 sg13g2_dfrbp_1 _2053_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net177),
    .D(net476),
    .Q_N(_0603_),
    .Q(\cellsbuf_[104].A ));
 sg13g2_dfrbp_1 _2054_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net176),
    .D(_0294_),
    .Q_N(_0602_),
    .Q(\cellsbuf_[105].A ));
 sg13g2_dfrbp_1 _2055_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net175),
    .D(_0295_),
    .Q_N(_0601_),
    .Q(\cellsbuf_[106].A ));
 sg13g2_dfrbp_1 _2056_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net174),
    .D(_0296_),
    .Q_N(_0600_),
    .Q(\cellsbuf_[107].A ));
 sg13g2_dfrbp_1 _2057_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net173),
    .D(_0297_),
    .Q_N(_0599_),
    .Q(\cellsbuf_[108].A ));
 sg13g2_dfrbp_1 _2058_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net172),
    .D(net478),
    .Q_N(_0598_),
    .Q(\cellsbuf_[109].A ));
 sg13g2_dfrbp_1 _2059_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net171),
    .D(net794),
    .Q_N(_0597_),
    .Q(\cellsbuf_[110].A ));
 sg13g2_dfrbp_1 _2060_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net170),
    .D(_0300_),
    .Q_N(_0596_),
    .Q(\cellsbuf_[111].A ));
 sg13g2_dfrbp_1 _2061_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net169),
    .D(_0301_),
    .Q_N(_0595_),
    .Q(\cellsbuf_[112].A ));
 sg13g2_dfrbp_1 _2062_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net168),
    .D(_0302_),
    .Q_N(_0594_),
    .Q(\cellsbuf_[113].A ));
 sg13g2_dfrbp_1 _2063_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net167),
    .D(net472),
    .Q_N(_0593_),
    .Q(\cellsbuf_[114].A ));
 sg13g2_dfrbp_1 _2064_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net166),
    .D(net708),
    .Q_N(_0592_),
    .Q(\cellsbuf_[115].A ));
 sg13g2_dfrbp_1 _2065_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net165),
    .D(_0305_),
    .Q_N(_0591_),
    .Q(\cellsbuf_[116].A ));
 sg13g2_dfrbp_1 _2066_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net164),
    .D(_0306_),
    .Q_N(_0590_),
    .Q(\cellsbuf_[117].A ));
 sg13g2_dfrbp_1 _2067_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net163),
    .D(_0307_),
    .Q_N(_0589_),
    .Q(\cellsbuf_[118].A ));
 sg13g2_dfrbp_1 _2068_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net162),
    .D(net536),
    .Q_N(_0588_),
    .Q(\cellsbuf_[119].A ));
 sg13g2_dfrbp_1 _2069_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net161),
    .D(_0309_),
    .Q_N(_0587_),
    .Q(\cellsbuf_[120].A ));
 sg13g2_dfrbp_1 _2070_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net160),
    .D(_0310_),
    .Q_N(_0586_),
    .Q(\cellsbuf_[121].A ));
 sg13g2_dfrbp_1 _2071_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net159),
    .D(net546),
    .Q_N(_0585_),
    .Q(\cellsbuf_[122].A ));
 sg13g2_dfrbp_1 _2072_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net158),
    .D(net606),
    .Q_N(_0584_),
    .Q(\cellsbuf_[123].A ));
 sg13g2_dfrbp_1 _2073_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net157),
    .D(_0313_),
    .Q_N(_0583_),
    .Q(\cellsbuf_[124].A ));
 sg13g2_dfrbp_1 _2074_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net156),
    .D(_0314_),
    .Q_N(_0582_),
    .Q(\cellsbuf_[125].A ));
 sg13g2_dfrbp_1 _2075_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net155),
    .D(net629),
    .Q_N(_0581_),
    .Q(\cellsbuf_[126].A ));
 sg13g2_dfrbp_1 _2076_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net154),
    .D(net724),
    .Q_N(_0580_),
    .Q(\cellsbuf_[127].A ));
 sg13g2_dfrbp_1 _2077_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net153),
    .D(_0317_),
    .Q_N(_0579_),
    .Q(\cellsbuf_[128].A ));
 sg13g2_dfrbp_1 _2078_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net152),
    .D(_0318_),
    .Q_N(_0578_),
    .Q(\cellsbuf_[129].A ));
 sg13g2_dfrbp_1 _2079_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net151),
    .D(_0319_),
    .Q_N(_0577_),
    .Q(\cellsbuf_[130].A ));
 sg13g2_dfrbp_1 _2080_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net150),
    .D(net522),
    .Q_N(_0576_),
    .Q(\cellsbuf_[131].A ));
 sg13g2_dfrbp_1 _2081_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net149),
    .D(_0321_),
    .Q_N(_0575_),
    .Q(\cellsbuf_[132].A ));
 sg13g2_dfrbp_1 _2082_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net148),
    .D(net444),
    .Q_N(_0574_),
    .Q(\cellsbuf_[133].A ));
 sg13g2_dfrbp_1 _2083_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net147),
    .D(_0323_),
    .Q_N(_0573_),
    .Q(\cellsbuf_[134].A ));
 sg13g2_dfrbp_1 _2084_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net146),
    .D(_0324_),
    .Q_N(_0572_),
    .Q(\cellsbuf_[135].A ));
 sg13g2_dfrbp_1 _2085_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net145),
    .D(net484),
    .Q_N(_0571_),
    .Q(\cellsbuf_[136].A ));
 sg13g2_dfrbp_1 _2086_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net144),
    .D(_0326_),
    .Q_N(_0570_),
    .Q(\cellsbuf_[137].A ));
 sg13g2_dfrbp_1 _2087_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net143),
    .D(_0327_),
    .Q_N(_0569_),
    .Q(\cellsbuf_[138].A ));
 sg13g2_dfrbp_1 _2088_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net142),
    .D(_0328_),
    .Q_N(_0568_),
    .Q(\cellsbuf_[139].A ));
 sg13g2_dfrbp_1 _2089_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net141),
    .D(net679),
    .Q_N(_0567_),
    .Q(\cellsbuf_[140].A ));
 sg13g2_dfrbp_1 _2090_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net140),
    .D(_0330_),
    .Q_N(_0566_),
    .Q(\cellsbuf_[141].A ));
 sg13g2_dfrbp_1 _2091_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net139),
    .D(net572),
    .Q_N(_0565_),
    .Q(\cellsbuf_[142].A ));
 sg13g2_dfrbp_1 _2092_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net138),
    .D(_0332_),
    .Q_N(_0564_),
    .Q(\cellsbuf_[143].A ));
 sg13g2_dfrbp_1 _2093_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net137),
    .D(net742),
    .Q_N(_0563_),
    .Q(\cellsbuf_[144].A ));
 sg13g2_dfrbp_1 _2094_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net136),
    .D(_0334_),
    .Q_N(_0562_),
    .Q(\cellsbuf_[145].A ));
 sg13g2_dfrbp_1 _2095_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net135),
    .D(net544),
    .Q_N(_0561_),
    .Q(\cellsbuf_[146].A ));
 sg13g2_dfrbp_1 _2096_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net134),
    .D(_0336_),
    .Q_N(_0560_),
    .Q(\cellsbuf_[147].A ));
 sg13g2_dfrbp_1 _2097_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net133),
    .D(_0337_),
    .Q_N(_0559_),
    .Q(\cellsbuf_[148].A ));
 sg13g2_dfrbp_1 _2098_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net132),
    .D(net800),
    .Q_N(_0558_),
    .Q(\cellsbuf_[149].A ));
 sg13g2_dfrbp_1 _2099_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net131),
    .D(_0339_),
    .Q_N(_0557_),
    .Q(\cellsbuf_[150].A ));
 sg13g2_dfrbp_1 _2100_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net130),
    .D(_0340_),
    .Q_N(_0556_),
    .Q(\cellsbuf_[151].A ));
 sg13g2_dfrbp_1 _2101_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net129),
    .D(net470),
    .Q_N(_0555_),
    .Q(\cellsbuf_[152].A ));
 sg13g2_dfrbp_1 _2102_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net128),
    .D(_0342_),
    .Q_N(_0554_),
    .Q(\cellsbuf_[153].A ));
 sg13g2_dfrbp_1 _2103_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net127),
    .D(_0343_),
    .Q_N(_0553_),
    .Q(\cellsbuf_[154].A ));
 sg13g2_dfrbp_1 _2104_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net126),
    .D(net654),
    .Q_N(_0552_),
    .Q(\cellsbuf_[155].A ));
 sg13g2_dfrbp_1 _2105_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net125),
    .D(net865),
    .Q_N(_0551_),
    .Q(\cellsbuf_[156].A ));
 sg13g2_dfrbp_1 _2106_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net124),
    .D(net904),
    .Q_N(_0550_),
    .Q(\cellsbuf_[157].A ));
 sg13g2_dfrbp_1 _2107_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net123),
    .D(net934),
    .Q_N(_0549_),
    .Q(\cellsbuf_[158].A ));
 sg13g2_dfrbp_1 _2108_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net122),
    .D(_0348_),
    .Q_N(_0548_),
    .Q(\cellsbuf_[159].A ));
 sg13g2_dfrbp_1 _2109_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net121),
    .D(_0349_),
    .Q_N(_0547_),
    .Q(\next_cellsbuf_[0].A ));
 sg13g2_dfrbp_1 _2110_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net120),
    .D(net442),
    .Q_N(_0016_),
    .Q(\row_count[0] ));
 sg13g2_dfrbp_1 _2111_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net118),
    .D(net937),
    .Q_N(_0546_),
    .Q(\row_count[1] ));
 sg13g2_dfrbp_1 _2112_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net116),
    .D(net932),
    .Q_N(_0545_),
    .Q(\row_count[2] ));
 sg13g2_dfrbp_1 _2113_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net114),
    .D(net966),
    .Q_N(_0011_),
    .Q(\row_count[3] ));
 sg13g2_dfrbp_1 _2114_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net112),
    .D(net911),
    .Q_N(_0014_),
    .Q(\row_count[4] ));
 sg13g2_dfrbp_1 _2115_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net110),
    .D(_0355_),
    .Q_N(_0544_),
    .Q(\row_count[5] ));
 sg13g2_dfrbp_1 _2116_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net108),
    .D(net925),
    .Q_N(_0543_),
    .Q(\row_count[6] ));
 sg13g2_dfrbp_1 _2117_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net106),
    .D(net964),
    .Q_N(_0010_),
    .Q(\row_count[7] ));
 sg13g2_dfrbp_1 _2118_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net104),
    .D(net946),
    .Q_N(_0012_),
    .Q(\i[0] ));
 sg13g2_dfrbp_1 _2119_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net102),
    .D(net942),
    .Q_N(_0009_),
    .Q(\i[1] ));
 sg13g2_dfrbp_1 _2120_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net422),
    .D(net923),
    .Q_N(_0013_),
    .Q(\i[2] ));
 sg13g2_dfrbp_1 _2121_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net423),
    .D(_0000_),
    .Q_N(_0878_),
    .Q(\rule[0] ));
 sg13g2_dfrbp_1 _2122_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net424),
    .D(_0001_),
    .Q_N(_0879_),
    .Q(\rule[1] ));
 sg13g2_dfrbp_1 _2123_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net425),
    .D(_0002_),
    .Q_N(_0880_),
    .Q(\rule[2] ));
 sg13g2_dfrbp_1 _2124_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net426),
    .D(_0003_),
    .Q_N(_0881_),
    .Q(\rule[3] ));
 sg13g2_dfrbp_1 _2125_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net427),
    .D(_0004_),
    .Q_N(_0882_),
    .Q(\rule[4] ));
 sg13g2_dfrbp_1 _2126_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net428),
    .D(_0005_),
    .Q_N(_0883_),
    .Q(\rule[5] ));
 sg13g2_dfrbp_1 _2127_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net439),
    .D(_0006_),
    .Q_N(_0884_),
    .Q(\rule[6] ));
 sg13g2_dfrbp_1 _2128_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net100),
    .D(_0007_),
    .Q_N(_0542_),
    .Q(hsync));
 sg13g2_dfrbp_1 _2129_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net119),
    .D(net919),
    .Q_N(_0015_),
    .Q(\fract_y[0] ));
 sg13g2_dfrbp_1 _2130_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net115),
    .D(_0362_),
    .Q_N(_0541_),
    .Q(\fract_y[1] ));
 sg13g2_dfrbp_1 _2131_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net111),
    .D(_0363_),
    .Q_N(_0540_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _2132_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net107),
    .D(_0364_),
    .Q_N(_0539_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _2133_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net103),
    .D(_0365_),
    .Q_N(_0538_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _2134_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net97),
    .D(_0366_),
    .Q_N(_0537_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _2135_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net113),
    .D(_0367_),
    .Q_N(_0536_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _2136_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net105),
    .D(net928),
    .Q_N(_0535_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _2137_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net117),
    .D(_0369_),
    .Q_N(_0534_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _2138_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net109),
    .D(net949),
    .Q_N(_0885_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _2139_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net101),
    .D(net846),
    .Q_N(_0533_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_tiehi _1859__18 (.L_HI(net18));
 sg13g2_tiehi _1858__19 (.L_HI(net19));
 sg13g2_tiehi _1857__20 (.L_HI(net20));
 sg13g2_tiehi _1856__21 (.L_HI(net21));
 sg13g2_tiehi _1855__22 (.L_HI(net22));
 sg13g2_tiehi _1854__23 (.L_HI(net23));
 sg13g2_tiehi _1853__24 (.L_HI(net24));
 sg13g2_tiehi _1852__25 (.L_HI(net25));
 sg13g2_tiehi _1851__26 (.L_HI(net26));
 sg13g2_tiehi _1850__27 (.L_HI(net27));
 sg13g2_tiehi _1849__28 (.L_HI(net28));
 sg13g2_tiehi _1848__29 (.L_HI(net29));
 sg13g2_tiehi _1847__30 (.L_HI(net30));
 sg13g2_tiehi _1846__31 (.L_HI(net31));
 sg13g2_tiehi _1845__32 (.L_HI(net32));
 sg13g2_tiehi _1844__33 (.L_HI(net33));
 sg13g2_tiehi _1843__34 (.L_HI(net34));
 sg13g2_tiehi _1842__35 (.L_HI(net35));
 sg13g2_tiehi _1841__36 (.L_HI(net36));
 sg13g2_tiehi _1840__37 (.L_HI(net37));
 sg13g2_tiehi _1839__38 (.L_HI(net38));
 sg13g2_tiehi _1838__39 (.L_HI(net39));
 sg13g2_tiehi _1837__40 (.L_HI(net40));
 sg13g2_tiehi _1836__41 (.L_HI(net41));
 sg13g2_tiehi _1835__42 (.L_HI(net42));
 sg13g2_tiehi _1834__43 (.L_HI(net43));
 sg13g2_tiehi _1833__44 (.L_HI(net44));
 sg13g2_tiehi _1832__45 (.L_HI(net45));
 sg13g2_tiehi _1831__46 (.L_HI(net46));
 sg13g2_tiehi _1830__47 (.L_HI(net47));
 sg13g2_tiehi _1829__48 (.L_HI(net48));
 sg13g2_tiehi _1828__49 (.L_HI(net49));
 sg13g2_tiehi _1827__50 (.L_HI(net50));
 sg13g2_tiehi _1826__51 (.L_HI(net51));
 sg13g2_tiehi _1825__52 (.L_HI(net52));
 sg13g2_tiehi _1824__53 (.L_HI(net53));
 sg13g2_tiehi _1823__54 (.L_HI(net54));
 sg13g2_tiehi _1822__55 (.L_HI(net55));
 sg13g2_tiehi _1821__56 (.L_HI(net56));
 sg13g2_tiehi _1820__57 (.L_HI(net57));
 sg13g2_tiehi _1819__58 (.L_HI(net58));
 sg13g2_tiehi _1818__59 (.L_HI(net59));
 sg13g2_tiehi _1817__60 (.L_HI(net60));
 sg13g2_tiehi _1816__61 (.L_HI(net61));
 sg13g2_tiehi _1815__62 (.L_HI(net62));
 sg13g2_tiehi _1814__63 (.L_HI(net63));
 sg13g2_tiehi _1813__64 (.L_HI(net64));
 sg13g2_tiehi _1812__65 (.L_HI(net65));
 sg13g2_tiehi _1811__66 (.L_HI(net66));
 sg13g2_tiehi _1810__67 (.L_HI(net67));
 sg13g2_tiehi _1809__68 (.L_HI(net68));
 sg13g2_tiehi _1808__69 (.L_HI(net69));
 sg13g2_tiehi _1807__70 (.L_HI(net70));
 sg13g2_tiehi _1806__71 (.L_HI(net71));
 sg13g2_tiehi _1805__72 (.L_HI(net72));
 sg13g2_tiehi _1804__73 (.L_HI(net73));
 sg13g2_tiehi _1803__74 (.L_HI(net74));
 sg13g2_tiehi _1802__75 (.L_HI(net75));
 sg13g2_tiehi _1801__76 (.L_HI(net76));
 sg13g2_tiehi _1800__77 (.L_HI(net77));
 sg13g2_tiehi _1799__78 (.L_HI(net78));
 sg13g2_tiehi _1798__79 (.L_HI(net79));
 sg13g2_tiehi _1797__80 (.L_HI(net80));
 sg13g2_tiehi _1796__81 (.L_HI(net81));
 sg13g2_tiehi _1795__82 (.L_HI(net82));
 sg13g2_tiehi _1794__83 (.L_HI(net83));
 sg13g2_tiehi _1793__84 (.L_HI(net84));
 sg13g2_tiehi _1792__85 (.L_HI(net85));
 sg13g2_tiehi _1791__86 (.L_HI(net86));
 sg13g2_tiehi _1790__87 (.L_HI(net87));
 sg13g2_tiehi _1789__88 (.L_HI(net88));
 sg13g2_tiehi _1788__89 (.L_HI(net89));
 sg13g2_tiehi _1787__90 (.L_HI(net90));
 sg13g2_tiehi _1786__91 (.L_HI(net91));
 sg13g2_tiehi _1785__92 (.L_HI(net92));
 sg13g2_tiehi _1784__93 (.L_HI(net93));
 sg13g2_tiehi _1783__94 (.L_HI(net94));
 sg13g2_tiehi _1782__95 (.L_HI(net95));
 sg13g2_tiehi _1781__96 (.L_HI(net96));
 sg13g2_tiehi _2134__97 (.L_HI(net97));
 sg13g2_tiehi _1780__98 (.L_HI(net98));
 sg13g2_tiehi _1779__99 (.L_HI(net99));
 sg13g2_tiehi _2128__100 (.L_HI(net100));
 sg13g2_tiehi _2139__101 (.L_HI(net101));
 sg13g2_tiehi _2119__102 (.L_HI(net102));
 sg13g2_tiehi _2133__103 (.L_HI(net103));
 sg13g2_tiehi _2118__104 (.L_HI(net104));
 sg13g2_tiehi _2136__105 (.L_HI(net105));
 sg13g2_tiehi _2117__106 (.L_HI(net106));
 sg13g2_tiehi _2132__107 (.L_HI(net107));
 sg13g2_tiehi _2116__108 (.L_HI(net108));
 sg13g2_tiehi _2138__109 (.L_HI(net109));
 sg13g2_tiehi _2115__110 (.L_HI(net110));
 sg13g2_tiehi _2131__111 (.L_HI(net111));
 sg13g2_tiehi _2114__112 (.L_HI(net112));
 sg13g2_tiehi _2135__113 (.L_HI(net113));
 sg13g2_tiehi _2113__114 (.L_HI(net114));
 sg13g2_tiehi _2130__115 (.L_HI(net115));
 sg13g2_tiehi _2112__116 (.L_HI(net116));
 sg13g2_tiehi _2137__117 (.L_HI(net117));
 sg13g2_tiehi _2111__118 (.L_HI(net118));
 sg13g2_tiehi _2129__119 (.L_HI(net119));
 sg13g2_tiehi _2110__120 (.L_HI(net120));
 sg13g2_tiehi _2109__121 (.L_HI(net121));
 sg13g2_tiehi _2108__122 (.L_HI(net122));
 sg13g2_tiehi _2107__123 (.L_HI(net123));
 sg13g2_tiehi _2106__124 (.L_HI(net124));
 sg13g2_tiehi _2105__125 (.L_HI(net125));
 sg13g2_tiehi _2104__126 (.L_HI(net126));
 sg13g2_tiehi _2103__127 (.L_HI(net127));
 sg13g2_tiehi _2102__128 (.L_HI(net128));
 sg13g2_tiehi _2101__129 (.L_HI(net129));
 sg13g2_tiehi _2100__130 (.L_HI(net130));
 sg13g2_tiehi _2099__131 (.L_HI(net131));
 sg13g2_tiehi _2098__132 (.L_HI(net132));
 sg13g2_tiehi _2097__133 (.L_HI(net133));
 sg13g2_tiehi _2096__134 (.L_HI(net134));
 sg13g2_tiehi _2095__135 (.L_HI(net135));
 sg13g2_tiehi _2094__136 (.L_HI(net136));
 sg13g2_tiehi _2093__137 (.L_HI(net137));
 sg13g2_tiehi _2092__138 (.L_HI(net138));
 sg13g2_tiehi _2091__139 (.L_HI(net139));
 sg13g2_tiehi _2090__140 (.L_HI(net140));
 sg13g2_tiehi _2089__141 (.L_HI(net141));
 sg13g2_tiehi _2088__142 (.L_HI(net142));
 sg13g2_tiehi _2087__143 (.L_HI(net143));
 sg13g2_tiehi _2086__144 (.L_HI(net144));
 sg13g2_tiehi _2085__145 (.L_HI(net145));
 sg13g2_tiehi _2084__146 (.L_HI(net146));
 sg13g2_tiehi _2083__147 (.L_HI(net147));
 sg13g2_tiehi _2082__148 (.L_HI(net148));
 sg13g2_tiehi _2081__149 (.L_HI(net149));
 sg13g2_tiehi _2080__150 (.L_HI(net150));
 sg13g2_tiehi _2079__151 (.L_HI(net151));
 sg13g2_tiehi _2078__152 (.L_HI(net152));
 sg13g2_tiehi _2077__153 (.L_HI(net153));
 sg13g2_tiehi _2076__154 (.L_HI(net154));
 sg13g2_tiehi _2075__155 (.L_HI(net155));
 sg13g2_tiehi _2074__156 (.L_HI(net156));
 sg13g2_tiehi _2073__157 (.L_HI(net157));
 sg13g2_tiehi _2072__158 (.L_HI(net158));
 sg13g2_tiehi _2071__159 (.L_HI(net159));
 sg13g2_tiehi _2070__160 (.L_HI(net160));
 sg13g2_tiehi _2069__161 (.L_HI(net161));
 sg13g2_tiehi _2068__162 (.L_HI(net162));
 sg13g2_tiehi _2067__163 (.L_HI(net163));
 sg13g2_tiehi _2066__164 (.L_HI(net164));
 sg13g2_tiehi _2065__165 (.L_HI(net165));
 sg13g2_tiehi _2064__166 (.L_HI(net166));
 sg13g2_tiehi _2063__167 (.L_HI(net167));
 sg13g2_tiehi _2062__168 (.L_HI(net168));
 sg13g2_tiehi _2061__169 (.L_HI(net169));
 sg13g2_tiehi _2060__170 (.L_HI(net170));
 sg13g2_tiehi _2059__171 (.L_HI(net171));
 sg13g2_tiehi _2058__172 (.L_HI(net172));
 sg13g2_tiehi _2057__173 (.L_HI(net173));
 sg13g2_tiehi _2056__174 (.L_HI(net174));
 sg13g2_tiehi _2055__175 (.L_HI(net175));
 sg13g2_tiehi _2054__176 (.L_HI(net176));
 sg13g2_tiehi _2053__177 (.L_HI(net177));
 sg13g2_tiehi _2052__178 (.L_HI(net178));
 sg13g2_tiehi _2051__179 (.L_HI(net179));
 sg13g2_tiehi _2050__180 (.L_HI(net180));
 sg13g2_tiehi _2049__181 (.L_HI(net181));
 sg13g2_tiehi _2048__182 (.L_HI(net182));
 sg13g2_tiehi _2047__183 (.L_HI(net183));
 sg13g2_tiehi _2046__184 (.L_HI(net184));
 sg13g2_tiehi _2045__185 (.L_HI(net185));
 sg13g2_tiehi _2044__186 (.L_HI(net186));
 sg13g2_tiehi _2043__187 (.L_HI(net187));
 sg13g2_tiehi _2042__188 (.L_HI(net188));
 sg13g2_tiehi _2041__189 (.L_HI(net189));
 sg13g2_tiehi _2040__190 (.L_HI(net190));
 sg13g2_tiehi _2039__191 (.L_HI(net191));
 sg13g2_tiehi _2038__192 (.L_HI(net192));
 sg13g2_tiehi _2037__193 (.L_HI(net193));
 sg13g2_tiehi _2036__194 (.L_HI(net255));
 sg13g2_tiehi _2035__195 (.L_HI(net256));
 sg13g2_tiehi _2034__196 (.L_HI(net257));
 sg13g2_tiehi _2033__197 (.L_HI(net258));
 sg13g2_tiehi _2032__198 (.L_HI(net259));
 sg13g2_tiehi _2031__199 (.L_HI(net260));
 sg13g2_tiehi _2030__200 (.L_HI(net261));
 sg13g2_tiehi _2029__201 (.L_HI(net262));
 sg13g2_tiehi _2028__202 (.L_HI(net263));
 sg13g2_tiehi _2027__203 (.L_HI(net264));
 sg13g2_tiehi _2026__204 (.L_HI(net265));
 sg13g2_tiehi _2025__205 (.L_HI(net266));
 sg13g2_tiehi _2024__206 (.L_HI(net267));
 sg13g2_tiehi _2023__207 (.L_HI(net268));
 sg13g2_tiehi _2022__208 (.L_HI(net269));
 sg13g2_tiehi _2021__209 (.L_HI(net270));
 sg13g2_tiehi _2020__210 (.L_HI(net271));
 sg13g2_tiehi _2019__211 (.L_HI(net272));
 sg13g2_tiehi _2018__212 (.L_HI(net273));
 sg13g2_tiehi _2017__213 (.L_HI(net274));
 sg13g2_tiehi _2016__214 (.L_HI(net275));
 sg13g2_tiehi _2015__215 (.L_HI(net276));
 sg13g2_tiehi _2014__216 (.L_HI(net277));
 sg13g2_tiehi _2013__217 (.L_HI(net278));
 sg13g2_tiehi _2012__218 (.L_HI(net279));
 sg13g2_tiehi _2011__219 (.L_HI(net280));
 sg13g2_tiehi _2010__220 (.L_HI(net281));
 sg13g2_tiehi _2009__221 (.L_HI(net282));
 sg13g2_tiehi _2008__222 (.L_HI(net283));
 sg13g2_tiehi _2007__223 (.L_HI(net284));
 sg13g2_tiehi _2006__224 (.L_HI(net285));
 sg13g2_tiehi _2005__225 (.L_HI(net286));
 sg13g2_tiehi _2004__226 (.L_HI(net287));
 sg13g2_tiehi _2003__227 (.L_HI(net288));
 sg13g2_tiehi _2002__228 (.L_HI(net289));
 sg13g2_tiehi _2001__229 (.L_HI(net290));
 sg13g2_tiehi _2000__230 (.L_HI(net291));
 sg13g2_tiehi _1999__231 (.L_HI(net292));
 sg13g2_tiehi _1998__232 (.L_HI(net293));
 sg13g2_tiehi _1997__233 (.L_HI(net294));
 sg13g2_tiehi _1996__234 (.L_HI(net295));
 sg13g2_tiehi _1995__235 (.L_HI(net296));
 sg13g2_tiehi _1994__236 (.L_HI(net297));
 sg13g2_tiehi _1993__237 (.L_HI(net298));
 sg13g2_tiehi _1992__238 (.L_HI(net299));
 sg13g2_tiehi _1991__239 (.L_HI(net300));
 sg13g2_tiehi _1990__240 (.L_HI(net301));
 sg13g2_tiehi _1989__241 (.L_HI(net302));
 sg13g2_tiehi _1988__242 (.L_HI(net303));
 sg13g2_tiehi _1987__243 (.L_HI(net304));
 sg13g2_tiehi _1986__244 (.L_HI(net305));
 sg13g2_tiehi _1985__245 (.L_HI(net306));
 sg13g2_tiehi _1984__246 (.L_HI(net307));
 sg13g2_tiehi _1983__247 (.L_HI(net308));
 sg13g2_tiehi _1982__248 (.L_HI(net309));
 sg13g2_tiehi _1981__249 (.L_HI(net310));
 sg13g2_tiehi _1980__250 (.L_HI(net311));
 sg13g2_tiehi _1979__251 (.L_HI(net312));
 sg13g2_tiehi _1978__252 (.L_HI(net313));
 sg13g2_tiehi _1977__253 (.L_HI(net314));
 sg13g2_tiehi _1976__254 (.L_HI(net315));
 sg13g2_tiehi _1975__255 (.L_HI(net316));
 sg13g2_tiehi _1974__256 (.L_HI(net317));
 sg13g2_tiehi _1973__257 (.L_HI(net318));
 sg13g2_tiehi _1972__258 (.L_HI(net319));
 sg13g2_tiehi _1971__259 (.L_HI(net320));
 sg13g2_tiehi _1970__260 (.L_HI(net321));
 sg13g2_tiehi _1969__261 (.L_HI(net322));
 sg13g2_tiehi _1968__262 (.L_HI(net323));
 sg13g2_tiehi _1967__263 (.L_HI(net324));
 sg13g2_tiehi _1966__264 (.L_HI(net325));
 sg13g2_tiehi _1965__265 (.L_HI(net326));
 sg13g2_tiehi _1964__266 (.L_HI(net327));
 sg13g2_tiehi _1963__267 (.L_HI(net328));
 sg13g2_tiehi _1962__268 (.L_HI(net329));
 sg13g2_tiehi _1961__269 (.L_HI(net330));
 sg13g2_tiehi _1960__270 (.L_HI(net331));
 sg13g2_tiehi _1959__271 (.L_HI(net332));
 sg13g2_tiehi _1958__272 (.L_HI(net333));
 sg13g2_tiehi _1957__273 (.L_HI(net334));
 sg13g2_tiehi _1956__274 (.L_HI(net335));
 sg13g2_tiehi _1955__275 (.L_HI(net336));
 sg13g2_tiehi _1954__276 (.L_HI(net337));
 sg13g2_tiehi _1953__277 (.L_HI(net338));
 sg13g2_tiehi _1952__278 (.L_HI(net339));
 sg13g2_tiehi _1951__279 (.L_HI(net340));
 sg13g2_tiehi _1950__280 (.L_HI(net341));
 sg13g2_tiehi _1949__281 (.L_HI(net342));
 sg13g2_tiehi _1948__282 (.L_HI(net343));
 sg13g2_tiehi _1947__283 (.L_HI(net344));
 sg13g2_tiehi _1946__284 (.L_HI(net345));
 sg13g2_tiehi _1945__285 (.L_HI(net346));
 sg13g2_tiehi _1944__286 (.L_HI(net347));
 sg13g2_tiehi _1943__287 (.L_HI(net348));
 sg13g2_tiehi _1942__288 (.L_HI(net349));
 sg13g2_tiehi _1941__289 (.L_HI(net350));
 sg13g2_tiehi _1940__290 (.L_HI(net351));
 sg13g2_tiehi _1939__291 (.L_HI(net352));
 sg13g2_tiehi _1938__292 (.L_HI(net353));
 sg13g2_tiehi _1937__293 (.L_HI(net354));
 sg13g2_tiehi _1936__294 (.L_HI(net355));
 sg13g2_tiehi _1935__295 (.L_HI(net356));
 sg13g2_tiehi _1934__296 (.L_HI(net357));
 sg13g2_tiehi _1933__297 (.L_HI(net358));
 sg13g2_tiehi _1932__298 (.L_HI(net359));
 sg13g2_tiehi _1931__299 (.L_HI(net360));
 sg13g2_tiehi _1930__300 (.L_HI(net361));
 sg13g2_tiehi _1929__301 (.L_HI(net362));
 sg13g2_tiehi _1928__302 (.L_HI(net363));
 sg13g2_tiehi _1927__303 (.L_HI(net364));
 sg13g2_tiehi _1926__304 (.L_HI(net365));
 sg13g2_tiehi _1925__305 (.L_HI(net366));
 sg13g2_tiehi _1924__306 (.L_HI(net367));
 sg13g2_tiehi _1923__307 (.L_HI(net368));
 sg13g2_tiehi _1922__308 (.L_HI(net369));
 sg13g2_tiehi _1921__309 (.L_HI(net370));
 sg13g2_tiehi _1920__310 (.L_HI(net371));
 sg13g2_tiehi _1919__311 (.L_HI(net372));
 sg13g2_tiehi _1918__312 (.L_HI(net373));
 sg13g2_tiehi _1917__313 (.L_HI(net374));
 sg13g2_tiehi _1916__314 (.L_HI(net375));
 sg13g2_tiehi _1915__315 (.L_HI(net376));
 sg13g2_tiehi _1914__316 (.L_HI(net377));
 sg13g2_tiehi _1913__317 (.L_HI(net378));
 sg13g2_tiehi _1912__318 (.L_HI(net379));
 sg13g2_tiehi _1911__319 (.L_HI(net380));
 sg13g2_tiehi _1910__320 (.L_HI(net381));
 sg13g2_tiehi _1909__321 (.L_HI(net382));
 sg13g2_tiehi _1908__322 (.L_HI(net383));
 sg13g2_tiehi _1907__323 (.L_HI(net384));
 sg13g2_tiehi _1906__324 (.L_HI(net385));
 sg13g2_tiehi _1905__325 (.L_HI(net386));
 sg13g2_tiehi _1904__326 (.L_HI(net387));
 sg13g2_tiehi _1903__327 (.L_HI(net388));
 sg13g2_tiehi _1902__328 (.L_HI(net389));
 sg13g2_tiehi _1901__329 (.L_HI(net390));
 sg13g2_tiehi _1900__330 (.L_HI(net391));
 sg13g2_tiehi _1899__331 (.L_HI(net392));
 sg13g2_tiehi _1898__332 (.L_HI(net393));
 sg13g2_tiehi _1897__333 (.L_HI(net394));
 sg13g2_tiehi _1896__334 (.L_HI(net395));
 sg13g2_tiehi _1895__335 (.L_HI(net396));
 sg13g2_tiehi _1894__336 (.L_HI(net397));
 sg13g2_tiehi _1893__337 (.L_HI(net398));
 sg13g2_tiehi _1892__338 (.L_HI(net399));
 sg13g2_tiehi _1891__339 (.L_HI(net400));
 sg13g2_tiehi _1890__340 (.L_HI(net401));
 sg13g2_tiehi _1889__341 (.L_HI(net402));
 sg13g2_tiehi _1888__342 (.L_HI(net403));
 sg13g2_tiehi _1887__343 (.L_HI(net404));
 sg13g2_tiehi _1886__344 (.L_HI(net405));
 sg13g2_tiehi _1885__345 (.L_HI(net406));
 sg13g2_tiehi _1884__346 (.L_HI(net407));
 sg13g2_tiehi _1883__347 (.L_HI(net408));
 sg13g2_tiehi _1882__348 (.L_HI(net409));
 sg13g2_tiehi _1881__349 (.L_HI(net410));
 sg13g2_tiehi _1880__350 (.L_HI(net411));
 sg13g2_tiehi _1879__351 (.L_HI(net412));
 sg13g2_tiehi _1878__352 (.L_HI(net413));
 sg13g2_tiehi _1877__353 (.L_HI(net414));
 sg13g2_tiehi _1876__354 (.L_HI(net415));
 sg13g2_tiehi _1875__355 (.L_HI(net416));
 sg13g2_tiehi _1874__356 (.L_HI(net417));
 sg13g2_tiehi _1873__357 (.L_HI(net418));
 sg13g2_tiehi _1872__358 (.L_HI(net419));
 sg13g2_tiehi _1871__359 (.L_HI(net420));
 sg13g2_tiehi _1778__360 (.L_HI(net421));
 sg13g2_tiehi _2120__361 (.L_HI(net422));
 sg13g2_tiehi _2121__362 (.L_HI(net423));
 sg13g2_tiehi _2122__363 (.L_HI(net424));
 sg13g2_tiehi _2123__364 (.L_HI(net425));
 sg13g2_tiehi _2124__365 (.L_HI(net426));
 sg13g2_tiehi _2125__366 (.L_HI(net427));
 sg13g2_tiehi _2126__367 (.L_HI(net428));
 sg13g2_tiehi _1870__368 (.L_HI(net429));
 sg13g2_tiehi _1869__369 (.L_HI(net430));
 sg13g2_tiehi _1868__370 (.L_HI(net431));
 sg13g2_tiehi _1867__371 (.L_HI(net432));
 sg13g2_tiehi _1866__372 (.L_HI(net433));
 sg13g2_tiehi _1865__373 (.L_HI(net434));
 sg13g2_tiehi _1864__374 (.L_HI(net435));
 sg13g2_tiehi _1863__375 (.L_HI(net436));
 sg13g2_tiehi _1862__376 (.L_HI(net437));
 sg13g2_tiehi _1861__377 (.L_HI(net438));
 sg13g2_tiehi _2127__378 (.L_HI(net439));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_znah_vga_ca_2 (.L_LO(net2));
 sg13g2_tielo tt_um_znah_vga_ca_3 (.L_LO(net3));
 sg13g2_tielo tt_um_znah_vga_ca_4 (.L_LO(net4));
 sg13g2_tielo tt_um_znah_vga_ca_5 (.L_LO(net5));
 sg13g2_tielo tt_um_znah_vga_ca_6 (.L_LO(net6));
 sg13g2_tielo tt_um_znah_vga_ca_7 (.L_LO(net7));
 sg13g2_tielo tt_um_znah_vga_ca_8 (.L_LO(net8));
 sg13g2_tielo tt_um_znah_vga_ca_9 (.L_LO(net9));
 sg13g2_tielo tt_um_znah_vga_ca_10 (.L_LO(net10));
 sg13g2_tielo tt_um_znah_vga_ca_11 (.L_LO(net11));
 sg13g2_tielo tt_um_znah_vga_ca_12 (.L_LO(net12));
 sg13g2_tielo tt_um_znah_vga_ca_13 (.L_LO(net13));
 sg13g2_tielo tt_um_znah_vga_ca_14 (.L_LO(net14));
 sg13g2_tielo tt_um_znah_vga_ca_15 (.L_LO(net15));
 sg13g2_tielo tt_um_znah_vga_ca_16 (.L_LO(net16));
 sg13g2_tiehi _1860__17 (.L_HI(net17));
 sg13g2_buf_2 _2518_ (.A(\hvsync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _2519_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout194 (.X(net194),
    .A(net197));
 sg13g2_buf_2 fanout195 (.A(net197),
    .X(net195));
 sg13g2_buf_4 fanout196 (.X(net196),
    .A(net197));
 sg13g2_buf_2 fanout197 (.A(net219),
    .X(net197));
 sg13g2_buf_4 fanout198 (.X(net198),
    .A(net200));
 sg13g2_buf_4 fanout199 (.X(net199),
    .A(net200));
 sg13g2_buf_2 fanout200 (.A(net219),
    .X(net200));
 sg13g2_buf_4 fanout201 (.X(net201),
    .A(net203));
 sg13g2_buf_4 fanout202 (.X(net202),
    .A(net203));
 sg13g2_buf_4 fanout203 (.X(net203),
    .A(net207));
 sg13g2_buf_4 fanout204 (.X(net204),
    .A(net207));
 sg13g2_buf_2 fanout205 (.A(net207),
    .X(net205));
 sg13g2_buf_4 fanout206 (.X(net206),
    .A(net207));
 sg13g2_buf_2 fanout207 (.A(net219),
    .X(net207));
 sg13g2_buf_4 fanout208 (.X(net208),
    .A(net210));
 sg13g2_buf_2 fanout209 (.A(net210),
    .X(net209));
 sg13g2_buf_4 fanout210 (.X(net210),
    .A(net213));
 sg13g2_buf_4 fanout211 (.X(net211),
    .A(net212));
 sg13g2_buf_4 fanout212 (.X(net212),
    .A(net213));
 sg13g2_buf_2 fanout213 (.A(net219),
    .X(net213));
 sg13g2_buf_4 fanout214 (.X(net214),
    .A(net217));
 sg13g2_buf_4 fanout215 (.X(net215),
    .A(net216));
 sg13g2_buf_4 fanout216 (.X(net216),
    .A(net217));
 sg13g2_buf_2 fanout217 (.A(net218),
    .X(net217));
 sg13g2_buf_4 fanout218 (.X(net218),
    .A(net219));
 sg13g2_buf_4 fanout219 (.X(net219),
    .A(_0532_));
 sg13g2_buf_2 fanout220 (.A(_0465_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_0376_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_0376_),
    .X(net222));
 sg13g2_buf_4 fanout223 (.X(net223),
    .A(net226));
 sg13g2_buf_4 fanout224 (.X(net224),
    .A(net226));
 sg13g2_buf_4 fanout225 (.X(net225),
    .A(net226));
 sg13g2_buf_2 fanout226 (.A(net238),
    .X(net226));
 sg13g2_buf_4 fanout227 (.X(net227),
    .A(net230));
 sg13g2_buf_4 fanout228 (.X(net228),
    .A(net230));
 sg13g2_buf_4 fanout229 (.X(net229),
    .A(net230));
 sg13g2_buf_2 fanout230 (.A(net238),
    .X(net230));
 sg13g2_buf_4 fanout231 (.X(net231),
    .A(net234));
 sg13g2_buf_4 fanout232 (.X(net232),
    .A(net234));
 sg13g2_buf_2 fanout233 (.A(net234),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(net238),
    .X(net234));
 sg13g2_buf_4 fanout235 (.X(net235),
    .A(net237));
 sg13g2_buf_4 fanout236 (.X(net236),
    .A(net237));
 sg13g2_buf_4 fanout237 (.X(net237),
    .A(net238));
 sg13g2_buf_2 fanout238 (.A(_0507_),
    .X(net238));
 sg13g2_buf_4 fanout239 (.X(net239),
    .A(net245));
 sg13g2_buf_4 fanout240 (.X(net240),
    .A(net244));
 sg13g2_buf_2 fanout241 (.A(net244),
    .X(net241));
 sg13g2_buf_4 fanout242 (.X(net242),
    .A(net244));
 sg13g2_buf_2 fanout243 (.A(net244),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(net245),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_0507_),
    .X(net245));
 sg13g2_buf_4 fanout246 (.X(net246),
    .A(net249));
 sg13g2_buf_4 fanout247 (.X(net247),
    .A(net248));
 sg13g2_buf_4 fanout248 (.X(net248),
    .A(net249));
 sg13g2_buf_2 fanout249 (.A(net250),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_0507_),
    .X(net250));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(_0441_));
 sg13g2_buf_2 fanout252 (.A(net253),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(net254),
    .X(net253));
 sg13g2_buf_4 fanout254 (.X(net254),
    .A(rst_n));
 sg13g2_tielo tt_um_znah_vga_ca_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload0 (.A(clknet_leaf_44_clk));
 sg13g2_inv_4 clkload1 (.A(clknet_leaf_47_clk));
 sg13g2_inv_4 clkload2 (.A(clknet_leaf_35_clk));
 sg13g2_inv_2 clkload3 (.A(clknet_leaf_37_clk));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_31_clk));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_15_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_26_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_20_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0017_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0016_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0350_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold4 (.A(\cellsbuf_[132].A ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0322_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold6 (.A(\cell_x[1] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0378_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold8 (.A(\cellsbuf_[80].A ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0270_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold10 (.A(\cellsbuf_[14].A ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0204_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold12 (.A(\cellsbuf_[82].A ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0272_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold14 (.A(\next_cellsbuf_[110].A ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0131_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold16 (.A(\cellsbuf_[38].A ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0228_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold18 (.A(\cellsbuf_[67].A ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0257_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold20 (.A(\next_cellsbuf_[65].A ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0086_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold22 (.A(\cellsbuf_[56].A ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0246_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold24 (.A(\next_cellsbuf_[126].A ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0147_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold26 (.A(\cellsbuf_[1].A ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0191_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold28 (.A(\cellsbuf_[43].A ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0233_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold30 (.A(\cellsbuf_[151].A ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0341_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold32 (.A(\cellsbuf_[113].A ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0303_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold34 (.A(\cellsbuf_[17].A ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0207_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold36 (.A(\cellsbuf_[103].A ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0293_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold38 (.A(\cellsbuf_[108].A ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0298_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold40 (.A(\cellsbuf_[89].A ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0279_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold42 (.A(\cellsbuf_[58].A ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0248_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold44 (.A(\cellsbuf_[135].A ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0325_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold46 (.A(\next_cellsbuf_[113].A ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0133_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold48 (.A(\next_cellsbuf_[24].A ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0044_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold50 (.A(\cellsbuf_[11].A ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0201_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold52 (.A(\cellsbuf_[101].A ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0291_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold54 (.A(\cellsbuf_[36].A ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0226_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold56 (.A(\cellsbuf_[98].A ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0288_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold58 (.A(\cellsbuf_[49].A ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0239_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold60 (.A(\next_cellsbuf_[40].A ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0060_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold62 (.A(\next_cellsbuf_[138].A ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0158_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold64 (.A(\next_cellsbuf_[137].A ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0157_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold66 (.A(\next_cellsbuf_[109].A ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold67 (.A(\next_cellsbuf_[115].A ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0135_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold69 (.A(\next_cellsbuf_[20].A ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0040_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold71 (.A(\next_cellsbuf_[103].A ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0123_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold73 (.A(\next_cellsbuf_[157].A ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0177_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold75 (.A(\next_cellsbuf_[114].A ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold76 (.A(\next_cellsbuf_[108].A ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0128_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold78 (.A(\next_cellsbuf_[124].A ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0144_),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold80 (.A(\cellsbuf_[86].A ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0276_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold82 (.A(\cellsbuf_[130].A ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0320_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold84 (.A(\cellsbuf_[32].A ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0222_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold86 (.A(\next_cellsbuf_[6].A ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0027_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold88 (.A(\next_cellsbuf_[64].A ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold89 (.A(\next_cellsbuf_[67].A ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0087_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold91 (.A(\cellsbuf_[85].A ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold92 (.A(\next_cellsbuf_[77].A ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0097_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold94 (.A(\cellsbuf_[94].A ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0284_),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold96 (.A(\cellsbuf_[118].A ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0308_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold98 (.A(\next_cellsbuf_[104].A ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold99 (.A(\next_cellsbuf_[43].A ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0064_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold101 (.A(\cellsbuf_[73].A ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0263_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold103 (.A(\cellsbuf_[55].A ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold104 (.A(\cellsbuf_[145].A ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0335_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold106 (.A(\cellsbuf_[121].A ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0311_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold108 (.A(\cellsbuf_[18].A ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0208_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold110 (.A(\next_cellsbuf_[74].A ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0094_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold112 (.A(\cellsbuf_[107].A ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold113 (.A(\cellsbuf_[27].A ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0217_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold115 (.A(\cellsbuf_[48].A ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold116 (.A(\cellsbuf_[46].A ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0236_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold118 (.A(\cellsbuf_[70].A ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0260_),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold120 (.A(\next_cellsbuf_[100].A ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0120_),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold122 (.A(\cellsbuf_[33].A ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0223_),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold124 (.A(\cellsbuf_[84].A ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold125 (.A(\cellsbuf_[45].A ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold126 (.A(\next_cellsbuf_[38].A ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0058_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold128 (.A(\next_cellsbuf_[34].A ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0054_),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold130 (.A(\next_cellsbuf_[140].A ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0161_),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold132 (.A(\cellsbuf_[141].A ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0331_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold134 (.A(\next_cellsbuf_[102].A ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0122_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold136 (.A(\next_cellsbuf_[116].A ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold137 (.A(\next_cellsbuf_[42].A ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold138 (.A(\cellsbuf_[92].A ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0282_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold140 (.A(\cellsbuf_[8].A ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0198_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold142 (.A(\next_cellsbuf_[76].A ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0096_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold144 (.A(\cellsbuf_[42].A ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold145 (.A(\next_cellsbuf_[148].A ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0168_),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold147 (.A(\cellsbuf_[10].A ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold148 (.A(\next_cellsbuf_[31].A ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0051_),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold150 (.A(\next_cellsbuf_[156].A ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0176_),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold152 (.A(\next_cellsbuf_[27].A ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0047_),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold154 (.A(\cellsbuf_[71].A ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0261_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold156 (.A(\next_cellsbuf_[29].A ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0049_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold158 (.A(\cellsbuf_[112].A ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold159 (.A(\next_cellsbuf_[134].A ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0154_),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold161 (.A(\cellsbuf_[129].A ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold162 (.A(\next_cellsbuf_[1].A ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0022_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold164 (.A(\next_cellsbuf_[11].A ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0031_),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold166 (.A(\cellsbuf_[122].A ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0312_),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold168 (.A(\next_cellsbuf_[119].A ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0139_),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold170 (.A(\cellsbuf_[52].A ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0242_),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold172 (.A(\cellsbuf_[74].A ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0264_),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold174 (.A(\cellsbuf_[111].A ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold175 (.A(\next_cellsbuf_[19].A ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0039_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold177 (.A(\next_cellsbuf_[155].A ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0175_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold179 (.A(\next_cellsbuf_[3].A ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0023_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold181 (.A(\next_cellsbuf_[133].A ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0153_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold183 (.A(\next_cellsbuf_[128].A ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0148_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold185 (.A(\next_cellsbuf_[132].A ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0152_),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold187 (.A(\cellsbuf_[60].A ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0250_),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold189 (.A(\cellsbuf_[125].A ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0315_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold191 (.A(\cellsbuf_[25].A ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0215_),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold193 (.A(\next_cellsbuf_[122].A ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0142_),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold195 (.A(\next_cellsbuf_[5].A ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0025_),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold197 (.A(\next_cellsbuf_[4].A ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold198 (.A(\next_cellsbuf_[25].A ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold199 (.A(\cellsbuf_[128].A ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold200 (.A(\cellsbuf_[13].A ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold201 (.A(\next_cellsbuf_[49].A ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0069_),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold203 (.A(\next_cellsbuf_[94].A ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0114_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold205 (.A(\cellsbuf_[5].A ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0195_),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold207 (.A(\next_cellsbuf_[95].A ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold208 (.A(\next_cellsbuf_[83].A ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0103_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold210 (.A(\next_cellsbuf_[52].A ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0072_),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold212 (.A(\next_cellsbuf_[131].A ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0151_),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold214 (.A(\cellsbuf_[154].A ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0344_),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold216 (.A(\next_cellsbuf_[56].A ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0076_),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold218 (.A(\next_cellsbuf_[63].A ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0083_),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold220 (.A(\next_cellsbuf_[41].A ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold221 (.A(\cellsbuf_[61].A ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0251_),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold223 (.A(\next_cellsbuf_[143].A ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0163_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold225 (.A(\cellsbuf_[37].A ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold226 (.A(\next_cellsbuf_[50].A ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold227 (.A(\next_cellsbuf_[28].A ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold228 (.A(\next_cellsbuf_[75].A ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold229 (.A(\next_cellsbuf_[107].A ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0127_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold231 (.A(\next_cellsbuf_[144].A ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold232 (.A(\next_cellsbuf_[86].A ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0106_),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold234 (.A(\cellsbuf_[99].A ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0289_),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold236 (.A(\next_cellsbuf_[79].A ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0099_),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold238 (.A(\cellsbuf_[120].A ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold239 (.A(\cellsbuf_[139].A ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0329_),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold241 (.A(\cellsbuf_[91].A ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold242 (.A(\next_cellsbuf_[125].A ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold243 (.A(\next_cellsbuf_[87].A ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold244 (.A(\next_cellsbuf_[81].A ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0101_),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold246 (.A(\next_cellsbuf_[154].A ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0174_),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold248 (.A(\next_cellsbuf_[139].A ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold249 (.A(\cellsbuf_[47].A ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold250 (.A(\cellsbuf_[6].A ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0196_),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold252 (.A(\next_cellsbuf_[112].A ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0132_),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold254 (.A(\cellsbuf_[87].A ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0277_),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold256 (.A(\next_cellsbuf_[85].A ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0105_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold258 (.A(\next_cellsbuf_[130].A ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0150_),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold260 (.A(\cellsbuf_[93].A ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold261 (.A(\next_cellsbuf_[78].A ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold262 (.A(\cellsbuf_[150].A ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold263 (.A(\next_cellsbuf_[61].A ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0081_),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold265 (.A(\next_cellsbuf_[22].A ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0042_),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold267 (.A(\next_cellsbuf_[57].A ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold268 (.A(\cellsbuf_[114].A ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0304_),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold270 (.A(\next_cellsbuf_[47].A ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0067_),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold272 (.A(\cellsbuf_[30].A ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0220_),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold274 (.A(\next_cellsbuf_[153].A ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0173_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold276 (.A(\cellsbuf_[29].A ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold277 (.A(\next_cellsbuf_[135].A ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold278 (.A(\next_cellsbuf_[70].A ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0090_),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold280 (.A(\next_cellsbuf_[84].A ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold281 (.A(\next_cellsbuf_[18].A ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0038_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold283 (.A(\cellsbuf_[4].A ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold284 (.A(\cellsbuf_[126].A ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0316_),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold286 (.A(\next_cellsbuf_[99].A ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0119_),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold288 (.A(\cellsbuf_[88].A ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold289 (.A(\next_cellsbuf_[54].A ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0074_),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold291 (.A(\cellsbuf_[44].A ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold292 (.A(\cellsbuf_[34].A ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0224_),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold294 (.A(\cellsbuf_[131].A ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold295 (.A(\next_cellsbuf_[158].A ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0179_),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold297 (.A(\cellsbuf_[64].A ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0253_),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold299 (.A(\next_cellsbuf_[136].A ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold300 (.A(\next_cellsbuf_[39].A ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold301 (.A(\cellsbuf_[134].A ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold302 (.A(\cellsbuf_[143].A ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0333_),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold304 (.A(\cellsbuf_[117].A ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold305 (.A(\next_cellsbuf_[60].A ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0080_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold307 (.A(\cellsbuf_[102].A ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold308 (.A(\cellsbuf_[35].A ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold309 (.A(\cellsbuf_[59].A ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold310 (.A(\cellsbuf_[21].A ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0211_),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold312 (.A(\next_cellsbuf_[150].A ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0170_),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold314 (.A(\next_cellsbuf_[149].A ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold315 (.A(\next_cellsbuf_[152].A ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0172_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold317 (.A(\next_cellsbuf_[73].A ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold318 (.A(_0093_),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold319 (.A(\next_cellsbuf_[91].A ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0111_),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold321 (.A(\cellsbuf_[106].A ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold322 (.A(\next_cellsbuf_[30].A ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold323 (.A(\next_cellsbuf_[62].A ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold324 (.A(\next_cellsbuf_[123].A ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold325 (.A(\next_cellsbuf_[23].A ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold326 (.A(\next_cellsbuf_[55].A ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold327 (.A(\next_cellsbuf_[151].A ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold328 (.A(\cellsbuf_[138].A ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold329 (.A(\cellsbuf_[72].A ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold330 (.A(\cellsbuf_[54].A ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold331 (.A(\cellsbuf_[100].A ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold332 (.A(\cellsbuf_[96].A ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0286_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold334 (.A(\next_cellsbuf_[88].A ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold335 (.A(\next_cellsbuf_[10].A ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0030_),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold337 (.A(\cellsbuf_[97].A ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold338 (.A(\next_cellsbuf_[106].A ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0126_),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold340 (.A(\next_cellsbuf_[147].A ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0167_),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold342 (.A(\cellsbuf_[137].A ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold343 (.A(\cellsbuf_[50].A ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0240_),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold345 (.A(\cellsbuf_[83].A ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold346 (.A(\cellsbuf_[69].A ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold347 (.A(_0258_),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold348 (.A(\next_cellsbuf_[80].A ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold349 (.A(\next_cellsbuf_[8].A ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold350 (.A(_0028_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold351 (.A(\cellsbuf_[53].A ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold352 (.A(\next_cellsbuf_[129].A ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold353 (.A(\next_cellsbuf_[92].A ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold354 (.A(\cellsbuf_[109].A ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0299_),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold356 (.A(\next_cellsbuf_[58].A ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold357 (.A(\cellsbuf_[116].A ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold358 (.A(\cellsbuf_[26].A ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold359 (.A(\next_cellsbuf_[0].A ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold360 (.A(\cellsbuf_[148].A ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold361 (.A(_0338_),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold362 (.A(\next_cellsbuf_[120].A ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold363 (.A(\next_cellsbuf_[59].A ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold364 (.A(\cellsbuf_[153].A ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold365 (.A(\next_cellsbuf_[48].A ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold366 (.A(\next_cellsbuf_[12].A ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold367 (.A(\next_cellsbuf_[145].A ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold368 (.A(\next_cellsbuf_[82].A ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold369 (.A(\next_cellsbuf_[37].A ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0057_),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold371 (.A(\next_cellsbuf_[13].A ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold372 (.A(\next_cellsbuf_[142].A ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0162_),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold374 (.A(\next_cellsbuf_[36].A ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0056_),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold376 (.A(\next_cellsbuf_[93].A ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold377 (.A(\cellsbuf_[105].A ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold378 (.A(\next_cellsbuf_[46].A ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0066_),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold380 (.A(\cellsbuf_[124].A ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold381 (.A(\cellsbuf_[75].A ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0265_),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold383 (.A(\next_cellsbuf_[51].A ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold384 (.A(\cellsbuf_[66].A ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold385 (.A(\next_cellsbuf_[97].A ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0117_),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold387 (.A(\cellsbuf_[95].A ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold388 (.A(\next_cellsbuf_[89].A ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold389 (.A(\cellsbuf_[31].A ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold390 (.A(\cellsbuf_[65].A ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold391 (.A(\cellsbuf_[3].A ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold392 (.A(\next_cellsbuf_[117].A ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold393 (.A(\cellsbuf_[81].A ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold394 (.A(\next_cellsbuf_[69].A ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0089_),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold396 (.A(\cellsbuf_[110].A ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold397 (.A(\cellsbuf_[152].A ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold398 (.A(\cellsbuf_[76].A ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0266_),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold400 (.A(\next_cellsbuf_[121].A ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold401 (.A(\next_cellsbuf_[21].A ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold402 (.A(\next_cellsbuf_[32].A ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold403 (.A(\next_cellsbuf_[90].A ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold404 (.A(\cellsbuf_[136].A ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold405 (.A(\next_cellsbuf_[53].A ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold406 (.A(\fract_y[1] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0008_),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold408 (.A(\cellsbuf_[115].A ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold409 (.A(\next_cellsbuf_[35].A ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold410 (.A(\next_cellsbuf_[68].A ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold411 (.A(\next_cellsbuf_[105].A ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold412 (.A(\cellsbuf_[15].A ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0205_),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold414 (.A(\cellsbuf_[12].A ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold415 (.A(\next_cellsbuf_[16].A ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold416 (.A(_0036_),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold417 (.A(\next_cellsbuf_[26].A ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold418 (.A(\next_cellsbuf_[45].A ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold419 (.A(_0065_),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold420 (.A(\cellsbuf_[119].A ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold421 (.A(\cellsbuf_[40].A ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold422 (.A(_0230_),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold423 (.A(\cellsbuf_[79].A ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold424 (.A(\cellsbuf_[28].A ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold425 (.A(\cellsbuf_[155].A ),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold426 (.A(_0345_),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold427 (.A(\cellsbuf_[41].A ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold428 (.A(\cellsbuf_[62].A ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold429 (.A(_0252_),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold430 (.A(\next_cellsbuf_[98].A ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold431 (.A(\cellsbuf_[23].A ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold432 (.A(_0213_),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold433 (.A(\cellsbuf_[104].A ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold434 (.A(\cellsbuf_[9].A ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold435 (.A(\cellsbuf_[78].A ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold436 (.A(\cellsbuf_[51].A ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold437 (.A(\cellsbuf_[0].A ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold438 (.A(\cellsbuf_[133].A ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold439 (.A(\cellsbuf_[24].A ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold440 (.A(\cellsbuf_[7].A ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold441 (.A(\next_cellsbuf_[33].A ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold442 (.A(\cellsbuf_[39].A ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold443 (.A(\cellsbuf_[16].A ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold444 (.A(\cellsbuf_[77].A ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold445 (.A(\next_cellsbuf_[146].A ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold446 (.A(\next_cellsbuf_[15].A ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold447 (.A(_0035_),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold448 (.A(\next_cellsbuf_[14].A ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold449 (.A(\cellsbuf_[140].A ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold450 (.A(\next_cellsbuf_[71].A ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold451 (.A(\next_cellsbuf_[72].A ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold452 (.A(\next_cellsbuf_[9].A ),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold453 (.A(\cellsbuf_[127].A ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold454 (.A(\cellsbuf_[57].A ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold455 (.A(\next_cellsbuf_[118].A ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold456 (.A(\cellsbuf_[149].A ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold457 (.A(\cellsbuf_[144].A ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold458 (.A(\cellsbuf_[147].A ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold459 (.A(\next_cellsbuf_[101].A ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold460 (.A(\cellsbuf_[123].A ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold461 (.A(\cellsbuf_[19].A ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold462 (.A(_0209_),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold463 (.A(\cellsbuf_[90].A ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold464 (.A(\cellsbuf_[156].A ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold465 (.A(_0346_),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold466 (.A(\next_cellsbuf_[96].A ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold467 (.A(\cellsbuf_[146].A ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold468 (.A(\cellsbuf_[22].A ),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold469 (.A(\cellsbuf_[20].A ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold470 (.A(\cellsbuf_[142].A ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold471 (.A(_0014_),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold472 (.A(_0354_),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold473 (.A(\cellsbuf_[2].A ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold474 (.A(\cell_x[6] ),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold475 (.A(_0385_),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold476 (.A(\next_cellsbuf_[17].A ),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold477 (.A(\hvsync_gen.vpos[2] ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold478 (.A(_0015_),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold479 (.A(_0416_),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold480 (.A(_0361_),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold481 (.A(\hvsync_gen.vpos[5] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold482 (.A(_0425_),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold483 (.A(\i[2] ),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold484 (.A(_0360_),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold485 (.A(\row_count[6] ),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold486 (.A(_0356_),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold487 (.A(\hvsync_gen.vpos[7] ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold488 (.A(_0428_),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold489 (.A(_0368_),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold490 (.A(\row_count[5] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold491 (.A(_0402_),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold492 (.A(\row_count[2] ),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold493 (.A(_0352_),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold494 (.A(\cellsbuf_[157].A ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold495 (.A(_0347_),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold496 (.A(\row_count[1] ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold497 (.A(_0391_),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold498 (.A(_0351_),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold499 (.A(\cell_x[3] ),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold500 (.A(_0381_),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold501 (.A(_0185_),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold502 (.A(\i[1] ),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold503 (.A(_0359_),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold504 (.A(\cellsbuf_[159].A ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold505 (.A(_0019_),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold506 (.A(\i[0] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold507 (.A(_0358_),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold508 (.A(\hvsync_gen.vpos[8] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold509 (.A(_0433_),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold510 (.A(_0370_),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold511 (.A(\cellsbuf_[158].A ),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold512 (.A(\cell_x[0] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold513 (.A(_0377_),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold514 (.A(\hvsync_gen.vpos[3] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold515 (.A(\hvsync_gen.vpos[6] ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold516 (.A(\cell_x[4] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold517 (.A(_0383_),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold518 (.A(\cell_x[7] ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold519 (.A(_0388_),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold520 (.A(\cell_x[5] ),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold521 (.A(\hvsync_gen.vpos[4] ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold522 (.A(_0424_),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold523 (.A(\cell_x[2] ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold524 (.A(\row_count[7] ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold525 (.A(_0357_),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold526 (.A(\row_count[3] ),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold527 (.A(_0353_),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold528 (.A(\cell_x[2] ),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold529 (.A(_0184_),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold530 (.A(\fract_x[1] ),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold531 (.A(_0452_),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold532 (.A(_0181_),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold533 (.A(\fract_x[1] ),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold534 (.A(\cell_x[5] ),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold535 (.A(\hvsync_gen.vpos[4] ),
    .X(net974));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_4 FILLER_13_56 ();
 sg13g2_fill_1 FILLER_13_60 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_4 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_74 ();
 sg13g2_decap_8 FILLER_14_81 ();
 sg13g2_decap_8 FILLER_14_88 ();
 sg13g2_decap_8 FILLER_14_95 ();
 sg13g2_decap_8 FILLER_14_102 ();
 sg13g2_decap_8 FILLER_14_109 ();
 sg13g2_decap_8 FILLER_14_116 ();
 sg13g2_decap_8 FILLER_14_123 ();
 sg13g2_decap_8 FILLER_14_130 ();
 sg13g2_decap_8 FILLER_14_137 ();
 sg13g2_decap_8 FILLER_14_144 ();
 sg13g2_decap_8 FILLER_14_151 ();
 sg13g2_decap_8 FILLER_14_158 ();
 sg13g2_decap_8 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_decap_8 FILLER_14_179 ();
 sg13g2_decap_8 FILLER_14_186 ();
 sg13g2_decap_8 FILLER_14_193 ();
 sg13g2_decap_8 FILLER_14_200 ();
 sg13g2_decap_8 FILLER_14_207 ();
 sg13g2_decap_8 FILLER_14_214 ();
 sg13g2_decap_8 FILLER_14_221 ();
 sg13g2_decap_8 FILLER_14_228 ();
 sg13g2_decap_8 FILLER_14_235 ();
 sg13g2_decap_8 FILLER_14_242 ();
 sg13g2_decap_8 FILLER_14_249 ();
 sg13g2_decap_8 FILLER_14_256 ();
 sg13g2_decap_8 FILLER_14_263 ();
 sg13g2_decap_8 FILLER_14_270 ();
 sg13g2_decap_8 FILLER_14_277 ();
 sg13g2_decap_8 FILLER_14_284 ();
 sg13g2_decap_8 FILLER_14_291 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_fill_2 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_318 ();
 sg13g2_decap_4 FILLER_14_325 ();
 sg13g2_decap_8 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_4 FILLER_15_35 ();
 sg13g2_fill_1 FILLER_15_85 ();
 sg13g2_decap_8 FILLER_15_99 ();
 sg13g2_decap_8 FILLER_15_106 ();
 sg13g2_decap_8 FILLER_15_113 ();
 sg13g2_decap_8 FILLER_15_120 ();
 sg13g2_decap_8 FILLER_15_127 ();
 sg13g2_decap_8 FILLER_15_134 ();
 sg13g2_decap_8 FILLER_15_141 ();
 sg13g2_decap_8 FILLER_15_148 ();
 sg13g2_decap_8 FILLER_15_155 ();
 sg13g2_decap_8 FILLER_15_162 ();
 sg13g2_decap_8 FILLER_15_169 ();
 sg13g2_decap_8 FILLER_15_176 ();
 sg13g2_decap_8 FILLER_15_183 ();
 sg13g2_decap_8 FILLER_15_190 ();
 sg13g2_decap_8 FILLER_15_197 ();
 sg13g2_decap_8 FILLER_15_204 ();
 sg13g2_decap_8 FILLER_15_211 ();
 sg13g2_decap_8 FILLER_15_218 ();
 sg13g2_decap_8 FILLER_15_225 ();
 sg13g2_decap_8 FILLER_15_232 ();
 sg13g2_decap_8 FILLER_15_239 ();
 sg13g2_decap_8 FILLER_15_246 ();
 sg13g2_decap_8 FILLER_15_253 ();
 sg13g2_decap_4 FILLER_15_260 ();
 sg13g2_fill_2 FILLER_15_264 ();
 sg13g2_decap_8 FILLER_15_270 ();
 sg13g2_decap_8 FILLER_15_277 ();
 sg13g2_decap_4 FILLER_15_284 ();
 sg13g2_decap_4 FILLER_15_298 ();
 sg13g2_fill_1 FILLER_15_302 ();
 sg13g2_decap_8 FILLER_15_347 ();
 sg13g2_decap_8 FILLER_15_354 ();
 sg13g2_decap_8 FILLER_15_361 ();
 sg13g2_decap_8 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_4 FILLER_15_403 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_fill_1 FILLER_16_61 ();
 sg13g2_decap_8 FILLER_16_102 ();
 sg13g2_decap_8 FILLER_16_109 ();
 sg13g2_decap_8 FILLER_16_116 ();
 sg13g2_decap_8 FILLER_16_123 ();
 sg13g2_decap_8 FILLER_16_130 ();
 sg13g2_decap_8 FILLER_16_137 ();
 sg13g2_decap_8 FILLER_16_144 ();
 sg13g2_decap_8 FILLER_16_151 ();
 sg13g2_decap_8 FILLER_16_158 ();
 sg13g2_decap_8 FILLER_16_165 ();
 sg13g2_decap_8 FILLER_16_172 ();
 sg13g2_decap_8 FILLER_16_179 ();
 sg13g2_decap_8 FILLER_16_186 ();
 sg13g2_decap_8 FILLER_16_193 ();
 sg13g2_decap_8 FILLER_16_200 ();
 sg13g2_decap_8 FILLER_16_207 ();
 sg13g2_decap_8 FILLER_16_214 ();
 sg13g2_decap_8 FILLER_16_221 ();
 sg13g2_decap_8 FILLER_16_228 ();
 sg13g2_decap_8 FILLER_16_235 ();
 sg13g2_fill_1 FILLER_16_242 ();
 sg13g2_decap_4 FILLER_16_253 ();
 sg13g2_fill_1 FILLER_16_257 ();
 sg13g2_decap_4 FILLER_16_285 ();
 sg13g2_decap_8 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_fill_2 FILLER_17_35 ();
 sg13g2_fill_1 FILLER_17_37 ();
 sg13g2_fill_2 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_fill_2 FILLER_17_264 ();
 sg13g2_decap_8 FILLER_17_276 ();
 sg13g2_fill_1 FILLER_17_283 ();
 sg13g2_fill_2 FILLER_17_314 ();
 sg13g2_fill_1 FILLER_17_316 ();
 sg13g2_decap_8 FILLER_17_369 ();
 sg13g2_decap_8 FILLER_17_376 ();
 sg13g2_decap_8 FILLER_17_383 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_fill_1 FILLER_18_54 ();
 sg13g2_decap_8 FILLER_18_115 ();
 sg13g2_decap_8 FILLER_18_122 ();
 sg13g2_decap_8 FILLER_18_129 ();
 sg13g2_decap_8 FILLER_18_136 ();
 sg13g2_decap_8 FILLER_18_143 ();
 sg13g2_decap_8 FILLER_18_150 ();
 sg13g2_decap_8 FILLER_18_157 ();
 sg13g2_decap_8 FILLER_18_164 ();
 sg13g2_decap_8 FILLER_18_171 ();
 sg13g2_decap_8 FILLER_18_178 ();
 sg13g2_decap_8 FILLER_18_185 ();
 sg13g2_decap_8 FILLER_18_192 ();
 sg13g2_decap_8 FILLER_18_199 ();
 sg13g2_decap_8 FILLER_18_206 ();
 sg13g2_fill_2 FILLER_18_213 ();
 sg13g2_fill_2 FILLER_18_330 ();
 sg13g2_decap_8 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_375 ();
 sg13g2_decap_8 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_18_389 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_fill_1 FILLER_19_21 ();
 sg13g2_fill_1 FILLER_19_83 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_4 FILLER_19_203 ();
 sg13g2_fill_2 FILLER_19_207 ();
 sg13g2_fill_1 FILLER_19_255 ();
 sg13g2_fill_2 FILLER_19_329 ();
 sg13g2_fill_1 FILLER_19_331 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_fill_2 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_30 ();
 sg13g2_decap_8 FILLER_20_137 ();
 sg13g2_decap_8 FILLER_20_144 ();
 sg13g2_decap_8 FILLER_20_151 ();
 sg13g2_decap_8 FILLER_20_158 ();
 sg13g2_decap_8 FILLER_20_165 ();
 sg13g2_decap_8 FILLER_20_172 ();
 sg13g2_decap_8 FILLER_20_179 ();
 sg13g2_decap_8 FILLER_20_186 ();
 sg13g2_decap_8 FILLER_20_193 ();
 sg13g2_decap_8 FILLER_20_200 ();
 sg13g2_decap_4 FILLER_20_207 ();
 sg13g2_fill_1 FILLER_20_265 ();
 sg13g2_fill_1 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_37 ();
 sg13g2_fill_2 FILLER_21_58 ();
 sg13g2_fill_1 FILLER_21_128 ();
 sg13g2_decap_8 FILLER_21_155 ();
 sg13g2_decap_8 FILLER_21_162 ();
 sg13g2_decap_8 FILLER_21_169 ();
 sg13g2_decap_8 FILLER_21_176 ();
 sg13g2_decap_8 FILLER_21_183 ();
 sg13g2_decap_8 FILLER_21_190 ();
 sg13g2_decap_8 FILLER_21_197 ();
 sg13g2_decap_8 FILLER_21_204 ();
 sg13g2_decap_8 FILLER_21_211 ();
 sg13g2_fill_1 FILLER_21_218 ();
 sg13g2_decap_4 FILLER_21_228 ();
 sg13g2_fill_1 FILLER_21_232 ();
 sg13g2_fill_1 FILLER_21_320 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_fill_2 FILLER_22_28 ();
 sg13g2_decap_4 FILLER_22_63 ();
 sg13g2_fill_1 FILLER_22_67 ();
 sg13g2_fill_2 FILLER_22_77 ();
 sg13g2_fill_1 FILLER_22_83 ();
 sg13g2_decap_8 FILLER_22_162 ();
 sg13g2_decap_8 FILLER_22_169 ();
 sg13g2_decap_8 FILLER_22_176 ();
 sg13g2_decap_8 FILLER_22_183 ();
 sg13g2_decap_8 FILLER_22_190 ();
 sg13g2_decap_8 FILLER_22_197 ();
 sg13g2_decap_8 FILLER_22_204 ();
 sg13g2_fill_2 FILLER_22_211 ();
 sg13g2_fill_1 FILLER_22_213 ();
 sg13g2_decap_8 FILLER_22_233 ();
 sg13g2_fill_1 FILLER_22_250 ();
 sg13g2_fill_2 FILLER_22_264 ();
 sg13g2_fill_1 FILLER_22_266 ();
 sg13g2_fill_1 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_4 FILLER_23_28 ();
 sg13g2_decap_4 FILLER_23_58 ();
 sg13g2_fill_2 FILLER_23_62 ();
 sg13g2_fill_2 FILLER_23_74 ();
 sg13g2_fill_1 FILLER_23_76 ();
 sg13g2_decap_8 FILLER_23_164 ();
 sg13g2_decap_8 FILLER_23_171 ();
 sg13g2_decap_8 FILLER_23_178 ();
 sg13g2_decap_8 FILLER_23_185 ();
 sg13g2_decap_8 FILLER_23_192 ();
 sg13g2_decap_8 FILLER_23_199 ();
 sg13g2_fill_1 FILLER_23_206 ();
 sg13g2_decap_4 FILLER_23_233 ();
 sg13g2_fill_1 FILLER_23_263 ();
 sg13g2_fill_1 FILLER_23_305 ();
 sg13g2_fill_2 FILLER_23_325 ();
 sg13g2_fill_2 FILLER_23_345 ();
 sg13g2_fill_1 FILLER_23_347 ();
 sg13g2_fill_2 FILLER_23_362 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_fill_2 FILLER_24_28 ();
 sg13g2_fill_1 FILLER_24_56 ();
 sg13g2_fill_2 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_142 ();
 sg13g2_decap_8 FILLER_24_156 ();
 sg13g2_fill_1 FILLER_24_163 ();
 sg13g2_decap_8 FILLER_24_169 ();
 sg13g2_decap_8 FILLER_24_176 ();
 sg13g2_decap_8 FILLER_24_183 ();
 sg13g2_decap_8 FILLER_24_190 ();
 sg13g2_decap_8 FILLER_24_197 ();
 sg13g2_decap_4 FILLER_24_204 ();
 sg13g2_fill_2 FILLER_24_208 ();
 sg13g2_fill_2 FILLER_24_293 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_fill_1 FILLER_24_322 ();
 sg13g2_fill_2 FILLER_24_332 ();
 sg13g2_fill_1 FILLER_24_334 ();
 sg13g2_fill_2 FILLER_24_365 ();
 sg13g2_fill_1 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_14 ();
 sg13g2_fill_2 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_56 ();
 sg13g2_decap_4 FILLER_25_131 ();
 sg13g2_decap_8 FILLER_25_177 ();
 sg13g2_decap_8 FILLER_25_184 ();
 sg13g2_decap_8 FILLER_25_191 ();
 sg13g2_decap_8 FILLER_25_198 ();
 sg13g2_decap_8 FILLER_25_205 ();
 sg13g2_fill_2 FILLER_25_212 ();
 sg13g2_fill_1 FILLER_25_214 ();
 sg13g2_fill_2 FILLER_25_305 ();
 sg13g2_fill_2 FILLER_25_327 ();
 sg13g2_fill_1 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_21 ();
 sg13g2_fill_2 FILLER_26_34 ();
 sg13g2_fill_2 FILLER_26_80 ();
 sg13g2_fill_2 FILLER_26_100 ();
 sg13g2_fill_1 FILLER_26_102 ();
 sg13g2_fill_2 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_180 ();
 sg13g2_decap_8 FILLER_26_187 ();
 sg13g2_decap_8 FILLER_26_194 ();
 sg13g2_decap_8 FILLER_26_201 ();
 sg13g2_fill_2 FILLER_26_208 ();
 sg13g2_fill_1 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_fill_2 FILLER_26_231 ();
 sg13g2_fill_1 FILLER_26_233 ();
 sg13g2_decap_4 FILLER_26_243 ();
 sg13g2_fill_1 FILLER_26_247 ();
 sg13g2_fill_1 FILLER_26_252 ();
 sg13g2_fill_1 FILLER_26_328 ();
 sg13g2_fill_1 FILLER_26_363 ();
 sg13g2_decap_8 FILLER_26_390 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_4 ();
 sg13g2_fill_2 FILLER_27_40 ();
 sg13g2_decap_4 FILLER_27_96 ();
 sg13g2_fill_2 FILLER_27_130 ();
 sg13g2_decap_8 FILLER_27_171 ();
 sg13g2_decap_8 FILLER_27_178 ();
 sg13g2_decap_8 FILLER_27_185 ();
 sg13g2_decap_4 FILLER_27_192 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_fill_2 FILLER_27_238 ();
 sg13g2_fill_1 FILLER_27_240 ();
 sg13g2_decap_4 FILLER_27_245 ();
 sg13g2_fill_2 FILLER_27_249 ();
 sg13g2_fill_2 FILLER_27_256 ();
 sg13g2_fill_2 FILLER_27_288 ();
 sg13g2_fill_1 FILLER_27_290 ();
 sg13g2_fill_1 FILLER_27_317 ();
 sg13g2_fill_1 FILLER_27_359 ();
 sg13g2_decap_8 FILLER_27_383 ();
 sg13g2_decap_8 FILLER_27_390 ();
 sg13g2_decap_8 FILLER_27_397 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_2 ();
 sg13g2_fill_1 FILLER_28_52 ();
 sg13g2_fill_1 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_169 ();
 sg13g2_decap_8 FILLER_28_176 ();
 sg13g2_fill_1 FILLER_28_183 ();
 sg13g2_fill_2 FILLER_28_239 ();
 sg13g2_fill_1 FILLER_28_241 ();
 sg13g2_fill_1 FILLER_28_273 ();
 sg13g2_decap_4 FILLER_28_296 ();
 sg13g2_fill_2 FILLER_28_300 ();
 sg13g2_fill_2 FILLER_28_350 ();
 sg13g2_fill_1 FILLER_28_352 ();
 sg13g2_decap_8 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_2 FILLER_29_26 ();
 sg13g2_fill_2 FILLER_29_80 ();
 sg13g2_fill_1 FILLER_29_82 ();
 sg13g2_decap_8 FILLER_29_123 ();
 sg13g2_decap_8 FILLER_29_162 ();
 sg13g2_decap_8 FILLER_29_169 ();
 sg13g2_decap_4 FILLER_29_176 ();
 sg13g2_fill_1 FILLER_29_180 ();
 sg13g2_fill_2 FILLER_29_246 ();
 sg13g2_fill_2 FILLER_29_258 ();
 sg13g2_fill_1 FILLER_29_260 ();
 sg13g2_decap_4 FILLER_29_302 ();
 sg13g2_fill_2 FILLER_29_306 ();
 sg13g2_fill_1 FILLER_29_336 ();
 sg13g2_fill_1 FILLER_29_351 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_fill_2 FILLER_30_66 ();
 sg13g2_fill_1 FILLER_30_68 ();
 sg13g2_fill_1 FILLER_30_111 ();
 sg13g2_decap_8 FILLER_30_164 ();
 sg13g2_decap_8 FILLER_30_171 ();
 sg13g2_fill_2 FILLER_30_178 ();
 sg13g2_fill_1 FILLER_30_233 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_decap_8 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_fill_2 FILLER_31_26 ();
 sg13g2_fill_1 FILLER_31_28 ();
 sg13g2_fill_2 FILLER_31_42 ();
 sg13g2_fill_1 FILLER_31_44 ();
 sg13g2_fill_2 FILLER_31_63 ();
 sg13g2_fill_2 FILLER_31_111 ();
 sg13g2_fill_1 FILLER_31_113 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_decap_8 FILLER_31_165 ();
 sg13g2_decap_8 FILLER_31_172 ();
 sg13g2_fill_2 FILLER_31_179 ();
 sg13g2_decap_8 FILLER_31_204 ();
 sg13g2_fill_1 FILLER_31_211 ();
 sg13g2_fill_1 FILLER_31_240 ();
 sg13g2_fill_1 FILLER_31_255 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_fill_2 FILLER_31_352 ();
 sg13g2_decap_8 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_15 ();
 sg13g2_fill_2 FILLER_32_35 ();
 sg13g2_fill_1 FILLER_32_37 ();
 sg13g2_decap_8 FILLER_32_104 ();
 sg13g2_fill_1 FILLER_32_111 ();
 sg13g2_decap_8 FILLER_32_165 ();
 sg13g2_decap_8 FILLER_32_172 ();
 sg13g2_decap_4 FILLER_32_179 ();
 sg13g2_fill_1 FILLER_32_183 ();
 sg13g2_fill_2 FILLER_32_203 ();
 sg13g2_fill_1 FILLER_32_205 ();
 sg13g2_fill_2 FILLER_32_225 ();
 sg13g2_fill_2 FILLER_32_231 ();
 sg13g2_fill_2 FILLER_32_334 ();
 sg13g2_decap_8 FILLER_32_384 ();
 sg13g2_decap_8 FILLER_32_391 ();
 sg13g2_decap_8 FILLER_32_398 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_104 ();
 sg13g2_fill_2 FILLER_33_125 ();
 sg13g2_fill_1 FILLER_33_127 ();
 sg13g2_decap_8 FILLER_33_155 ();
 sg13g2_decap_8 FILLER_33_162 ();
 sg13g2_decap_8 FILLER_33_169 ();
 sg13g2_fill_2 FILLER_33_176 ();
 sg13g2_fill_1 FILLER_33_178 ();
 sg13g2_decap_4 FILLER_33_205 ();
 sg13g2_fill_1 FILLER_33_209 ();
 sg13g2_fill_2 FILLER_33_280 ();
 sg13g2_fill_2 FILLER_33_327 ();
 sg13g2_fill_1 FILLER_33_338 ();
 sg13g2_decap_8 FILLER_33_375 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_fill_2 FILLER_34_26 ();
 sg13g2_fill_1 FILLER_34_28 ();
 sg13g2_fill_1 FILLER_34_138 ();
 sg13g2_decap_8 FILLER_34_158 ();
 sg13g2_decap_8 FILLER_34_165 ();
 sg13g2_decap_8 FILLER_34_172 ();
 sg13g2_fill_2 FILLER_34_236 ();
 sg13g2_fill_1 FILLER_34_306 ();
 sg13g2_decap_8 FILLER_34_372 ();
 sg13g2_decap_8 FILLER_34_379 ();
 sg13g2_decap_8 FILLER_34_386 ();
 sg13g2_decap_8 FILLER_34_393 ();
 sg13g2_decap_8 FILLER_34_400 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_42 ();
 sg13g2_fill_2 FILLER_35_62 ();
 sg13g2_fill_1 FILLER_35_64 ();
 sg13g2_fill_1 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_104 ();
 sg13g2_decap_8 FILLER_35_128 ();
 sg13g2_fill_2 FILLER_35_135 ();
 sg13g2_decap_8 FILLER_35_172 ();
 sg13g2_decap_4 FILLER_35_209 ();
 sg13g2_fill_2 FILLER_35_213 ();
 sg13g2_fill_2 FILLER_35_225 ();
 sg13g2_fill_1 FILLER_35_240 ();
 sg13g2_fill_2 FILLER_35_264 ();
 sg13g2_fill_1 FILLER_35_266 ();
 sg13g2_fill_2 FILLER_35_302 ();
 sg13g2_fill_1 FILLER_35_304 ();
 sg13g2_fill_2 FILLER_35_344 ();
 sg13g2_decap_8 FILLER_35_372 ();
 sg13g2_decap_8 FILLER_35_379 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_fill_2 FILLER_36_49 ();
 sg13g2_fill_2 FILLER_36_60 ();
 sg13g2_fill_1 FILLER_36_62 ();
 sg13g2_fill_1 FILLER_36_80 ();
 sg13g2_fill_2 FILLER_36_103 ();
 sg13g2_fill_1 FILLER_36_105 ();
 sg13g2_decap_4 FILLER_36_132 ();
 sg13g2_fill_1 FILLER_36_136 ();
 sg13g2_decap_8 FILLER_36_163 ();
 sg13g2_decap_8 FILLER_36_170 ();
 sg13g2_decap_8 FILLER_36_177 ();
 sg13g2_decap_4 FILLER_36_184 ();
 sg13g2_fill_2 FILLER_36_188 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_fill_1 FILLER_36_224 ();
 sg13g2_decap_4 FILLER_36_230 ();
 sg13g2_fill_2 FILLER_36_234 ();
 sg13g2_fill_2 FILLER_36_240 ();
 sg13g2_fill_2 FILLER_36_283 ();
 sg13g2_fill_2 FILLER_36_338 ();
 sg13g2_decap_8 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_fill_2 FILLER_37_19 ();
 sg13g2_fill_1 FILLER_37_21 ();
 sg13g2_decap_4 FILLER_37_52 ();
 sg13g2_fill_2 FILLER_37_86 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_fill_2 FILLER_37_105 ();
 sg13g2_decap_4 FILLER_37_129 ();
 sg13g2_fill_2 FILLER_37_137 ();
 sg13g2_fill_2 FILLER_37_149 ();
 sg13g2_decap_4 FILLER_37_173 ();
 sg13g2_decap_4 FILLER_37_216 ();
 sg13g2_fill_1 FILLER_37_220 ();
 sg13g2_fill_1 FILLER_37_240 ();
 sg13g2_fill_1 FILLER_37_303 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_fill_1 FILLER_38_19 ();
 sg13g2_fill_1 FILLER_38_85 ();
 sg13g2_decap_8 FILLER_38_158 ();
 sg13g2_decap_4 FILLER_38_165 ();
 sg13g2_fill_2 FILLER_38_205 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_368 ();
 sg13g2_decap_8 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_382 ();
 sg13g2_decap_8 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_fill_1 FILLER_39_35 ();
 sg13g2_fill_2 FILLER_39_46 ();
 sg13g2_fill_1 FILLER_39_48 ();
 sg13g2_fill_1 FILLER_39_87 ();
 sg13g2_fill_2 FILLER_39_114 ();
 sg13g2_fill_1 FILLER_39_121 ();
 sg13g2_decap_8 FILLER_39_148 ();
 sg13g2_decap_8 FILLER_39_155 ();
 sg13g2_fill_1 FILLER_39_162 ();
 sg13g2_fill_1 FILLER_39_199 ();
 sg13g2_fill_1 FILLER_39_274 ();
 sg13g2_fill_2 FILLER_39_311 ();
 sg13g2_fill_1 FILLER_39_313 ();
 sg13g2_decap_8 FILLER_39_355 ();
 sg13g2_decap_8 FILLER_39_362 ();
 sg13g2_decap_8 FILLER_39_369 ();
 sg13g2_decap_8 FILLER_39_376 ();
 sg13g2_decap_8 FILLER_39_383 ();
 sg13g2_decap_8 FILLER_39_390 ();
 sg13g2_decap_8 FILLER_39_397 ();
 sg13g2_decap_4 FILLER_39_404 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_fill_2 FILLER_40_36 ();
 sg13g2_fill_1 FILLER_40_52 ();
 sg13g2_fill_2 FILLER_40_57 ();
 sg13g2_fill_1 FILLER_40_59 ();
 sg13g2_fill_1 FILLER_40_105 ();
 sg13g2_decap_4 FILLER_40_168 ();
 sg13g2_fill_1 FILLER_40_172 ();
 sg13g2_fill_2 FILLER_40_186 ();
 sg13g2_fill_1 FILLER_40_188 ();
 sg13g2_fill_1 FILLER_40_216 ();
 sg13g2_fill_2 FILLER_40_237 ();
 sg13g2_fill_2 FILLER_40_265 ();
 sg13g2_fill_1 FILLER_40_267 ();
 sg13g2_decap_8 FILLER_40_355 ();
 sg13g2_decap_8 FILLER_40_362 ();
 sg13g2_decap_8 FILLER_40_369 ();
 sg13g2_decap_8 FILLER_40_376 ();
 sg13g2_decap_8 FILLER_40_383 ();
 sg13g2_decap_8 FILLER_40_390 ();
 sg13g2_decap_8 FILLER_40_397 ();
 sg13g2_decap_4 FILLER_40_404 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_41 ();
 sg13g2_fill_1 FILLER_41_68 ();
 sg13g2_fill_1 FILLER_41_84 ();
 sg13g2_decap_4 FILLER_41_174 ();
 sg13g2_fill_2 FILLER_41_188 ();
 sg13g2_fill_1 FILLER_41_190 ();
 sg13g2_fill_1 FILLER_41_200 ();
 sg13g2_decap_4 FILLER_41_246 ();
 sg13g2_fill_2 FILLER_41_254 ();
 sg13g2_fill_1 FILLER_41_256 ();
 sg13g2_fill_1 FILLER_41_287 ();
 sg13g2_fill_2 FILLER_41_321 ();
 sg13g2_decap_8 FILLER_41_359 ();
 sg13g2_decap_8 FILLER_41_366 ();
 sg13g2_decap_8 FILLER_41_373 ();
 sg13g2_decap_8 FILLER_41_380 ();
 sg13g2_decap_8 FILLER_41_387 ();
 sg13g2_decap_8 FILLER_41_394 ();
 sg13g2_decap_8 FILLER_41_401 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_11 ();
 sg13g2_fill_2 FILLER_42_32 ();
 sg13g2_fill_1 FILLER_42_61 ();
 sg13g2_fill_1 FILLER_42_119 ();
 sg13g2_decap_4 FILLER_42_129 ();
 sg13g2_decap_4 FILLER_42_187 ();
 sg13g2_decap_8 FILLER_42_235 ();
 sg13g2_decap_8 FILLER_42_242 ();
 sg13g2_fill_1 FILLER_42_249 ();
 sg13g2_decap_4 FILLER_42_259 ();
 sg13g2_fill_1 FILLER_42_295 ();
 sg13g2_fill_2 FILLER_42_305 ();
 sg13g2_fill_2 FILLER_42_316 ();
 sg13g2_fill_1 FILLER_42_326 ();
 sg13g2_decap_8 FILLER_42_367 ();
 sg13g2_decap_8 FILLER_42_374 ();
 sg13g2_decap_8 FILLER_42_381 ();
 sg13g2_decap_8 FILLER_42_388 ();
 sg13g2_decap_8 FILLER_42_395 ();
 sg13g2_decap_8 FILLER_42_402 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_16 ();
 sg13g2_fill_1 FILLER_43_32 ();
 sg13g2_decap_4 FILLER_43_86 ();
 sg13g2_fill_1 FILLER_43_90 ();
 sg13g2_fill_2 FILLER_43_108 ();
 sg13g2_fill_1 FILLER_43_110 ();
 sg13g2_decap_8 FILLER_43_128 ();
 sg13g2_fill_2 FILLER_43_139 ();
 sg13g2_fill_1 FILLER_43_190 ();
 sg13g2_fill_2 FILLER_43_230 ();
 sg13g2_fill_1 FILLER_43_232 ();
 sg13g2_decap_8 FILLER_43_360 ();
 sg13g2_decap_8 FILLER_43_367 ();
 sg13g2_decap_8 FILLER_43_374 ();
 sg13g2_decap_8 FILLER_43_381 ();
 sg13g2_decap_8 FILLER_43_388 ();
 sg13g2_decap_8 FILLER_43_395 ();
 sg13g2_decap_8 FILLER_43_402 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_2 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_fill_2 FILLER_44_103 ();
 sg13g2_fill_1 FILLER_44_105 ();
 sg13g2_fill_2 FILLER_44_159 ();
 sg13g2_decap_8 FILLER_44_210 ();
 sg13g2_decap_4 FILLER_44_217 ();
 sg13g2_fill_1 FILLER_44_221 ();
 sg13g2_fill_2 FILLER_44_303 ();
 sg13g2_fill_1 FILLER_44_315 ();
 sg13g2_fill_1 FILLER_44_325 ();
 sg13g2_decap_8 FILLER_44_361 ();
 sg13g2_decap_8 FILLER_44_368 ();
 sg13g2_decap_8 FILLER_44_375 ();
 sg13g2_decap_8 FILLER_44_382 ();
 sg13g2_decap_8 FILLER_44_389 ();
 sg13g2_decap_8 FILLER_44_396 ();
 sg13g2_decap_4 FILLER_44_403 ();
 sg13g2_fill_2 FILLER_44_407 ();
 sg13g2_fill_2 FILLER_45_26 ();
 sg13g2_fill_2 FILLER_45_93 ();
 sg13g2_fill_1 FILLER_45_95 ();
 sg13g2_fill_2 FILLER_45_105 ();
 sg13g2_fill_1 FILLER_45_107 ();
 sg13g2_fill_1 FILLER_45_183 ();
 sg13g2_fill_2 FILLER_45_203 ();
 sg13g2_fill_2 FILLER_45_265 ();
 sg13g2_fill_1 FILLER_45_267 ();
 sg13g2_decap_8 FILLER_45_359 ();
 sg13g2_decap_8 FILLER_45_366 ();
 sg13g2_decap_8 FILLER_45_373 ();
 sg13g2_decap_8 FILLER_45_380 ();
 sg13g2_decap_8 FILLER_45_387 ();
 sg13g2_decap_8 FILLER_45_394 ();
 sg13g2_decap_8 FILLER_45_401 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_2 ();
 sg13g2_fill_1 FILLER_46_22 ();
 sg13g2_decap_4 FILLER_46_84 ();
 sg13g2_decap_4 FILLER_46_92 ();
 sg13g2_fill_1 FILLER_46_96 ();
 sg13g2_fill_2 FILLER_46_143 ();
 sg13g2_decap_4 FILLER_46_163 ();
 sg13g2_fill_2 FILLER_46_179 ();
 sg13g2_fill_2 FILLER_46_191 ();
 sg13g2_fill_1 FILLER_46_193 ();
 sg13g2_decap_4 FILLER_46_211 ();
 sg13g2_fill_2 FILLER_46_272 ();
 sg13g2_decap_8 FILLER_46_353 ();
 sg13g2_decap_8 FILLER_46_360 ();
 sg13g2_decap_8 FILLER_46_367 ();
 sg13g2_decap_8 FILLER_46_374 ();
 sg13g2_decap_8 FILLER_46_381 ();
 sg13g2_decap_8 FILLER_46_388 ();
 sg13g2_decap_8 FILLER_46_395 ();
 sg13g2_decap_8 FILLER_46_402 ();
 sg13g2_fill_2 FILLER_47_26 ();
 sg13g2_fill_1 FILLER_47_63 ();
 sg13g2_decap_4 FILLER_47_130 ();
 sg13g2_fill_1 FILLER_47_147 ();
 sg13g2_fill_2 FILLER_47_153 ();
 sg13g2_fill_1 FILLER_47_163 ();
 sg13g2_fill_2 FILLER_47_216 ();
 sg13g2_fill_2 FILLER_47_241 ();
 sg13g2_fill_1 FILLER_47_243 ();
 sg13g2_fill_1 FILLER_47_249 ();
 sg13g2_fill_2 FILLER_47_277 ();
 sg13g2_fill_1 FILLER_47_279 ();
 sg13g2_fill_2 FILLER_47_303 ();
 sg13g2_fill_1 FILLER_47_324 ();
 sg13g2_decap_8 FILLER_47_339 ();
 sg13g2_decap_8 FILLER_47_346 ();
 sg13g2_decap_8 FILLER_47_353 ();
 sg13g2_decap_8 FILLER_47_360 ();
 sg13g2_decap_8 FILLER_47_367 ();
 sg13g2_decap_8 FILLER_47_374 ();
 sg13g2_decap_8 FILLER_47_381 ();
 sg13g2_decap_8 FILLER_47_388 ();
 sg13g2_decap_8 FILLER_47_395 ();
 sg13g2_decap_8 FILLER_47_402 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_2 ();
 sg13g2_fill_1 FILLER_48_22 ();
 sg13g2_fill_2 FILLER_48_32 ();
 sg13g2_fill_2 FILLER_48_92 ();
 sg13g2_fill_1 FILLER_48_94 ();
 sg13g2_decap_4 FILLER_48_121 ();
 sg13g2_decap_4 FILLER_48_144 ();
 sg13g2_fill_1 FILLER_48_240 ();
 sg13g2_fill_2 FILLER_48_246 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_fill_1 FILLER_48_312 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_fill_2 FILLER_48_406 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_fill_2 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_28 ();
 sg13g2_fill_1 FILLER_49_62 ();
 sg13g2_fill_2 FILLER_49_177 ();
 sg13g2_fill_2 FILLER_49_205 ();
 sg13g2_fill_1 FILLER_49_226 ();
 sg13g2_fill_1 FILLER_49_253 ();
 sg13g2_fill_2 FILLER_49_280 ();
 sg13g2_fill_1 FILLER_49_282 ();
 sg13g2_decap_4 FILLER_49_313 ();
 sg13g2_fill_1 FILLER_49_317 ();
 sg13g2_decap_8 FILLER_49_344 ();
 sg13g2_decap_8 FILLER_49_351 ();
 sg13g2_decap_8 FILLER_49_358 ();
 sg13g2_decap_8 FILLER_49_365 ();
 sg13g2_decap_8 FILLER_49_372 ();
 sg13g2_decap_8 FILLER_49_379 ();
 sg13g2_decap_8 FILLER_49_386 ();
 sg13g2_decap_8 FILLER_49_393 ();
 sg13g2_decap_8 FILLER_49_400 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_fill_1 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_58 ();
 sg13g2_fill_2 FILLER_50_83 ();
 sg13g2_decap_8 FILLER_50_120 ();
 sg13g2_fill_1 FILLER_50_127 ();
 sg13g2_fill_2 FILLER_50_154 ();
 sg13g2_fill_2 FILLER_50_197 ();
 sg13g2_fill_2 FILLER_50_225 ();
 sg13g2_fill_1 FILLER_50_227 ();
 sg13g2_fill_2 FILLER_50_242 ();
 sg13g2_fill_1 FILLER_50_244 ();
 sg13g2_fill_1 FILLER_50_277 ();
 sg13g2_decap_8 FILLER_50_339 ();
 sg13g2_decap_8 FILLER_50_346 ();
 sg13g2_decap_8 FILLER_50_353 ();
 sg13g2_decap_8 FILLER_50_360 ();
 sg13g2_decap_8 FILLER_50_367 ();
 sg13g2_decap_8 FILLER_50_374 ();
 sg13g2_decap_8 FILLER_50_381 ();
 sg13g2_decap_8 FILLER_50_388 ();
 sg13g2_decap_8 FILLER_50_395 ();
 sg13g2_decap_8 FILLER_50_402 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_2 ();
 sg13g2_decap_8 FILLER_51_67 ();
 sg13g2_fill_1 FILLER_51_74 ();
 sg13g2_fill_1 FILLER_51_136 ();
 sg13g2_fill_2 FILLER_51_173 ();
 sg13g2_fill_1 FILLER_51_175 ();
 sg13g2_fill_1 FILLER_51_201 ();
 sg13g2_fill_2 FILLER_51_216 ();
 sg13g2_fill_2 FILLER_51_244 ();
 sg13g2_fill_2 FILLER_51_268 ();
 sg13g2_fill_2 FILLER_51_307 ();
 sg13g2_fill_1 FILLER_51_309 ();
 sg13g2_decap_8 FILLER_51_347 ();
 sg13g2_decap_8 FILLER_51_354 ();
 sg13g2_decap_8 FILLER_51_361 ();
 sg13g2_decap_8 FILLER_51_368 ();
 sg13g2_decap_8 FILLER_51_375 ();
 sg13g2_decap_8 FILLER_51_382 ();
 sg13g2_decap_8 FILLER_51_389 ();
 sg13g2_decap_8 FILLER_51_396 ();
 sg13g2_decap_4 FILLER_51_403 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_7 ();
 sg13g2_decap_4 FILLER_52_12 ();
 sg13g2_fill_2 FILLER_52_16 ();
 sg13g2_fill_2 FILLER_52_45 ();
 sg13g2_fill_1 FILLER_52_56 ();
 sg13g2_fill_2 FILLER_52_83 ();
 sg13g2_fill_2 FILLER_52_201 ();
 sg13g2_fill_1 FILLER_52_203 ();
 sg13g2_fill_1 FILLER_52_225 ();
 sg13g2_fill_1 FILLER_52_240 ();
 sg13g2_fill_1 FILLER_52_255 ();
 sg13g2_fill_1 FILLER_52_304 ();
 sg13g2_decap_8 FILLER_52_357 ();
 sg13g2_decap_8 FILLER_52_364 ();
 sg13g2_decap_8 FILLER_52_371 ();
 sg13g2_decap_8 FILLER_52_378 ();
 sg13g2_decap_8 FILLER_52_385 ();
 sg13g2_decap_8 FILLER_52_392 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_fill_2 FILLER_52_406 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_2 ();
 sg13g2_fill_2 FILLER_53_59 ();
 sg13g2_fill_1 FILLER_53_61 ();
 sg13g2_fill_2 FILLER_53_88 ();
 sg13g2_fill_1 FILLER_53_90 ();
 sg13g2_fill_1 FILLER_53_105 ();
 sg13g2_decap_4 FILLER_53_189 ();
 sg13g2_fill_1 FILLER_53_193 ();
 sg13g2_fill_2 FILLER_53_220 ();
 sg13g2_fill_1 FILLER_53_222 ();
 sg13g2_fill_2 FILLER_53_244 ();
 sg13g2_fill_2 FILLER_53_277 ();
 sg13g2_fill_1 FILLER_53_279 ();
 sg13g2_fill_2 FILLER_53_308 ();
 sg13g2_fill_1 FILLER_53_310 ();
 sg13g2_fill_2 FILLER_53_320 ();
 sg13g2_decap_8 FILLER_53_363 ();
 sg13g2_decap_8 FILLER_53_370 ();
 sg13g2_decap_8 FILLER_53_377 ();
 sg13g2_decap_8 FILLER_53_384 ();
 sg13g2_decap_8 FILLER_53_391 ();
 sg13g2_decap_8 FILLER_53_398 ();
 sg13g2_decap_4 FILLER_53_405 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_21 ();
 sg13g2_fill_1 FILLER_54_57 ();
 sg13g2_fill_2 FILLER_54_111 ();
 sg13g2_fill_1 FILLER_54_151 ();
 sg13g2_fill_1 FILLER_54_183 ();
 sg13g2_fill_2 FILLER_54_227 ();
 sg13g2_decap_4 FILLER_54_268 ();
 sg13g2_fill_1 FILLER_54_272 ();
 sg13g2_fill_2 FILLER_54_281 ();
 sg13g2_fill_1 FILLER_54_283 ();
 sg13g2_fill_2 FILLER_54_308 ();
 sg13g2_decap_8 FILLER_54_359 ();
 sg13g2_decap_8 FILLER_54_366 ();
 sg13g2_decap_8 FILLER_54_373 ();
 sg13g2_decap_8 FILLER_54_380 ();
 sg13g2_decap_8 FILLER_54_387 ();
 sg13g2_decap_8 FILLER_54_394 ();
 sg13g2_decap_8 FILLER_54_401 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_fill_2 FILLER_55_26 ();
 sg13g2_fill_2 FILLER_55_47 ();
 sg13g2_fill_1 FILLER_55_84 ();
 sg13g2_fill_2 FILLER_55_100 ();
 sg13g2_fill_1 FILLER_55_120 ();
 sg13g2_fill_2 FILLER_55_157 ();
 sg13g2_fill_1 FILLER_55_159 ();
 sg13g2_fill_1 FILLER_55_164 ();
 sg13g2_fill_1 FILLER_55_196 ();
 sg13g2_fill_2 FILLER_55_206 ();
 sg13g2_fill_2 FILLER_55_221 ();
 sg13g2_fill_2 FILLER_55_232 ();
 sg13g2_decap_4 FILLER_55_265 ();
 sg13g2_fill_1 FILLER_55_279 ();
 sg13g2_fill_2 FILLER_55_325 ();
 sg13g2_fill_1 FILLER_55_327 ();
 sg13g2_decap_8 FILLER_55_368 ();
 sg13g2_decap_8 FILLER_55_375 ();
 sg13g2_decap_8 FILLER_55_382 ();
 sg13g2_decap_8 FILLER_55_389 ();
 sg13g2_decap_8 FILLER_55_396 ();
 sg13g2_decap_4 FILLER_55_403 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_21 ();
 sg13g2_fill_1 FILLER_56_23 ();
 sg13g2_fill_1 FILLER_56_52 ();
 sg13g2_fill_2 FILLER_56_67 ();
 sg13g2_fill_1 FILLER_56_69 ();
 sg13g2_fill_1 FILLER_56_113 ();
 sg13g2_fill_2 FILLER_56_155 ();
 sg13g2_decap_8 FILLER_56_175 ();
 sg13g2_fill_2 FILLER_56_182 ();
 sg13g2_fill_2 FILLER_56_208 ();
 sg13g2_fill_1 FILLER_56_210 ();
 sg13g2_decap_8 FILLER_56_372 ();
 sg13g2_decap_8 FILLER_56_379 ();
 sg13g2_decap_8 FILLER_56_386 ();
 sg13g2_decap_8 FILLER_56_393 ();
 sg13g2_decap_8 FILLER_56_400 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_fill_1 FILLER_57_56 ();
 sg13g2_fill_1 FILLER_57_83 ();
 sg13g2_fill_1 FILLER_57_119 ();
 sg13g2_fill_2 FILLER_57_138 ();
 sg13g2_fill_1 FILLER_57_140 ();
 sg13g2_fill_1 FILLER_57_150 ();
 sg13g2_decap_4 FILLER_57_181 ();
 sg13g2_fill_2 FILLER_57_185 ();
 sg13g2_fill_2 FILLER_57_197 ();
 sg13g2_fill_1 FILLER_57_199 ();
 sg13g2_fill_2 FILLER_57_215 ();
 sg13g2_fill_1 FILLER_57_217 ();
 sg13g2_fill_1 FILLER_57_244 ();
 sg13g2_fill_2 FILLER_57_280 ();
 sg13g2_fill_1 FILLER_57_282 ();
 sg13g2_decap_8 FILLER_57_371 ();
 sg13g2_decap_8 FILLER_57_378 ();
 sg13g2_decap_8 FILLER_57_385 ();
 sg13g2_decap_8 FILLER_57_392 ();
 sg13g2_decap_8 FILLER_57_399 ();
 sg13g2_fill_2 FILLER_57_406 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_fill_2 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_2 ();
 sg13g2_fill_2 FILLER_58_50 ();
 sg13g2_fill_1 FILLER_58_52 ();
 sg13g2_fill_2 FILLER_58_151 ();
 sg13g2_fill_1 FILLER_58_172 ();
 sg13g2_fill_2 FILLER_58_220 ();
 sg13g2_fill_1 FILLER_58_245 ();
 sg13g2_fill_1 FILLER_58_263 ();
 sg13g2_decap_8 FILLER_58_287 ();
 sg13g2_decap_8 FILLER_58_294 ();
 sg13g2_decap_4 FILLER_58_301 ();
 sg13g2_fill_2 FILLER_58_305 ();
 sg13g2_fill_1 FILLER_58_317 ();
 sg13g2_fill_2 FILLER_58_342 ();
 sg13g2_fill_1 FILLER_58_344 ();
 sg13g2_decap_8 FILLER_58_371 ();
 sg13g2_decap_8 FILLER_58_378 ();
 sg13g2_decap_8 FILLER_58_385 ();
 sg13g2_decap_8 FILLER_58_392 ();
 sg13g2_decap_8 FILLER_58_399 ();
 sg13g2_fill_2 FILLER_58_406 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_21 ();
 sg13g2_fill_2 FILLER_59_56 ();
 sg13g2_fill_2 FILLER_59_68 ();
 sg13g2_fill_1 FILLER_59_98 ();
 sg13g2_fill_2 FILLER_59_109 ();
 sg13g2_fill_1 FILLER_59_111 ();
 sg13g2_fill_2 FILLER_59_138 ();
 sg13g2_fill_1 FILLER_59_166 ();
 sg13g2_decap_4 FILLER_59_187 ();
 sg13g2_fill_1 FILLER_59_202 ();
 sg13g2_fill_1 FILLER_59_213 ();
 sg13g2_fill_1 FILLER_59_220 ();
 sg13g2_decap_4 FILLER_59_235 ();
 sg13g2_fill_2 FILLER_59_239 ();
 sg13g2_decap_8 FILLER_59_294 ();
 sg13g2_decap_8 FILLER_59_301 ();
 sg13g2_decap_4 FILLER_59_308 ();
 sg13g2_decap_8 FILLER_59_373 ();
 sg13g2_decap_8 FILLER_59_380 ();
 sg13g2_decap_8 FILLER_59_387 ();
 sg13g2_decap_8 FILLER_59_394 ();
 sg13g2_decap_8 FILLER_59_401 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_fill_2 FILLER_60_40 ();
 sg13g2_fill_2 FILLER_60_69 ();
 sg13g2_fill_1 FILLER_60_71 ();
 sg13g2_fill_2 FILLER_60_81 ();
 sg13g2_fill_1 FILLER_60_83 ();
 sg13g2_fill_1 FILLER_60_111 ();
 sg13g2_fill_2 FILLER_60_122 ();
 sg13g2_fill_1 FILLER_60_124 ();
 sg13g2_fill_2 FILLER_60_158 ();
 sg13g2_fill_1 FILLER_60_160 ();
 sg13g2_decap_8 FILLER_60_187 ();
 sg13g2_decap_4 FILLER_60_194 ();
 sg13g2_fill_2 FILLER_60_198 ();
 sg13g2_decap_8 FILLER_60_214 ();
 sg13g2_decap_4 FILLER_60_221 ();
 sg13g2_fill_2 FILLER_60_225 ();
 sg13g2_decap_8 FILLER_60_232 ();
 sg13g2_decap_8 FILLER_60_239 ();
 sg13g2_fill_1 FILLER_60_246 ();
 sg13g2_fill_2 FILLER_60_262 ();
 sg13g2_fill_1 FILLER_60_355 ();
 sg13g2_decap_8 FILLER_60_369 ();
 sg13g2_decap_8 FILLER_60_376 ();
 sg13g2_decap_8 FILLER_60_383 ();
 sg13g2_decap_8 FILLER_60_390 ();
 sg13g2_decap_8 FILLER_60_397 ();
 sg13g2_decap_4 FILLER_60_404 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_fill_2 FILLER_61_111 ();
 sg13g2_fill_1 FILLER_61_113 ();
 sg13g2_fill_1 FILLER_61_123 ();
 sg13g2_fill_1 FILLER_61_142 ();
 sg13g2_fill_2 FILLER_61_156 ();
 sg13g2_fill_1 FILLER_61_158 ();
 sg13g2_fill_2 FILLER_61_163 ();
 sg13g2_fill_1 FILLER_61_165 ();
 sg13g2_fill_2 FILLER_61_171 ();
 sg13g2_fill_1 FILLER_61_173 ();
 sg13g2_decap_8 FILLER_61_183 ();
 sg13g2_decap_8 FILLER_61_190 ();
 sg13g2_fill_2 FILLER_61_201 ();
 sg13g2_decap_4 FILLER_61_212 ();
 sg13g2_fill_1 FILLER_61_221 ();
 sg13g2_fill_1 FILLER_61_235 ();
 sg13g2_decap_4 FILLER_61_362 ();
 sg13g2_fill_1 FILLER_61_366 ();
 sg13g2_decap_8 FILLER_61_376 ();
 sg13g2_decap_8 FILLER_61_383 ();
 sg13g2_decap_8 FILLER_61_390 ();
 sg13g2_decap_8 FILLER_61_397 ();
 sg13g2_decap_4 FILLER_61_404 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_fill_1 FILLER_62_112 ();
 sg13g2_fill_1 FILLER_62_122 ();
 sg13g2_fill_2 FILLER_62_132 ();
 sg13g2_fill_1 FILLER_62_134 ();
 sg13g2_fill_1 FILLER_62_171 ();
 sg13g2_decap_4 FILLER_62_176 ();
 sg13g2_fill_1 FILLER_62_199 ();
 sg13g2_fill_1 FILLER_62_282 ();
 sg13g2_fill_2 FILLER_62_293 ();
 sg13g2_decap_8 FILLER_62_367 ();
 sg13g2_decap_8 FILLER_62_374 ();
 sg13g2_decap_8 FILLER_62_381 ();
 sg13g2_decap_8 FILLER_62_388 ();
 sg13g2_decap_8 FILLER_62_395 ();
 sg13g2_decap_8 FILLER_62_402 ();
 sg13g2_fill_1 FILLER_63_26 ();
 sg13g2_fill_1 FILLER_63_50 ();
 sg13g2_fill_2 FILLER_63_77 ();
 sg13g2_fill_2 FILLER_63_114 ();
 sg13g2_fill_2 FILLER_63_124 ();
 sg13g2_fill_1 FILLER_63_126 ();
 sg13g2_fill_2 FILLER_63_205 ();
 sg13g2_fill_1 FILLER_63_243 ();
 sg13g2_fill_2 FILLER_63_291 ();
 sg13g2_fill_1 FILLER_63_306 ();
 sg13g2_decap_8 FILLER_63_382 ();
 sg13g2_decap_8 FILLER_63_389 ();
 sg13g2_decap_8 FILLER_63_396 ();
 sg13g2_decap_4 FILLER_63_403 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_fill_1 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_147 ();
 sg13g2_fill_1 FILLER_64_159 ();
 sg13g2_decap_4 FILLER_64_174 ();
 sg13g2_fill_1 FILLER_64_178 ();
 sg13g2_fill_1 FILLER_64_218 ();
 sg13g2_fill_1 FILLER_64_244 ();
 sg13g2_fill_1 FILLER_64_302 ();
 sg13g2_fill_2 FILLER_64_316 ();
 sg13g2_fill_1 FILLER_64_336 ();
 sg13g2_fill_2 FILLER_64_351 ();
 sg13g2_fill_1 FILLER_64_353 ();
 sg13g2_decap_8 FILLER_64_389 ();
 sg13g2_decap_8 FILLER_64_396 ();
 sg13g2_decap_4 FILLER_64_403 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_fill_2 FILLER_65_30 ();
 sg13g2_fill_1 FILLER_65_32 ();
 sg13g2_fill_2 FILLER_65_78 ();
 sg13g2_fill_1 FILLER_65_90 ();
 sg13g2_fill_1 FILLER_65_104 ();
 sg13g2_fill_2 FILLER_65_142 ();
 sg13g2_fill_1 FILLER_65_153 ();
 sg13g2_decap_8 FILLER_65_167 ();
 sg13g2_decap_8 FILLER_65_174 ();
 sg13g2_decap_4 FILLER_65_181 ();
 sg13g2_decap_8 FILLER_65_204 ();
 sg13g2_fill_2 FILLER_65_272 ();
 sg13g2_fill_1 FILLER_65_274 ();
 sg13g2_decap_8 FILLER_65_305 ();
 sg13g2_decap_4 FILLER_65_312 ();
 sg13g2_fill_1 FILLER_65_316 ();
 sg13g2_fill_1 FILLER_65_358 ();
 sg13g2_decap_8 FILLER_65_385 ();
 sg13g2_decap_8 FILLER_65_392 ();
 sg13g2_decap_8 FILLER_65_399 ();
 sg13g2_fill_2 FILLER_65_406 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_4 FILLER_66_7 ();
 sg13g2_fill_2 FILLER_66_43 ();
 sg13g2_fill_1 FILLER_66_45 ();
 sg13g2_fill_1 FILLER_66_99 ();
 sg13g2_fill_2 FILLER_66_126 ();
 sg13g2_decap_4 FILLER_66_155 ();
 sg13g2_fill_2 FILLER_66_159 ();
 sg13g2_fill_1 FILLER_66_187 ();
 sg13g2_fill_2 FILLER_66_193 ();
 sg13g2_fill_1 FILLER_66_195 ();
 sg13g2_fill_2 FILLER_66_247 ();
 sg13g2_fill_1 FILLER_66_285 ();
 sg13g2_decap_8 FILLER_66_389 ();
 sg13g2_decap_8 FILLER_66_396 ();
 sg13g2_decap_4 FILLER_66_403 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_fill_1 FILLER_67_14 ();
 sg13g2_fill_2 FILLER_67_19 ();
 sg13g2_fill_1 FILLER_67_21 ();
 sg13g2_fill_2 FILLER_67_45 ();
 sg13g2_fill_1 FILLER_67_47 ();
 sg13g2_fill_1 FILLER_67_75 ();
 sg13g2_decap_8 FILLER_67_148 ();
 sg13g2_decap_4 FILLER_67_155 ();
 sg13g2_fill_2 FILLER_67_159 ();
 sg13g2_fill_1 FILLER_67_196 ();
 sg13g2_fill_2 FILLER_67_250 ();
 sg13g2_fill_1 FILLER_67_290 ();
 sg13g2_fill_1 FILLER_67_301 ();
 sg13g2_fill_2 FILLER_67_333 ();
 sg13g2_decap_8 FILLER_67_387 ();
 sg13g2_decap_8 FILLER_67_394 ();
 sg13g2_decap_8 FILLER_67_401 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_fill_1 FILLER_68_14 ();
 sg13g2_fill_2 FILLER_68_80 ();
 sg13g2_fill_1 FILLER_68_82 ();
 sg13g2_fill_1 FILLER_68_114 ();
 sg13g2_decap_8 FILLER_68_141 ();
 sg13g2_fill_2 FILLER_68_148 ();
 sg13g2_fill_1 FILLER_68_206 ();
 sg13g2_fill_1 FILLER_68_305 ();
 sg13g2_fill_2 FILLER_68_315 ();
 sg13g2_fill_1 FILLER_68_317 ();
 sg13g2_fill_1 FILLER_68_373 ();
 sg13g2_decap_8 FILLER_68_387 ();
 sg13g2_decap_8 FILLER_68_394 ();
 sg13g2_decap_8 FILLER_68_401 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_fill_2 FILLER_69_21 ();
 sg13g2_fill_1 FILLER_69_23 ();
 sg13g2_decap_4 FILLER_69_50 ();
 sg13g2_fill_2 FILLER_69_67 ();
 sg13g2_decap_8 FILLER_69_132 ();
 sg13g2_decap_8 FILLER_69_139 ();
 sg13g2_decap_4 FILLER_69_146 ();
 sg13g2_fill_1 FILLER_69_176 ();
 sg13g2_fill_2 FILLER_69_186 ();
 sg13g2_fill_1 FILLER_69_219 ();
 sg13g2_fill_1 FILLER_69_236 ();
 sg13g2_fill_1 FILLER_69_242 ();
 sg13g2_fill_2 FILLER_69_269 ();
 sg13g2_fill_1 FILLER_69_325 ();
 sg13g2_fill_1 FILLER_69_358 ();
 sg13g2_decap_8 FILLER_69_385 ();
 sg13g2_decap_8 FILLER_69_392 ();
 sg13g2_decap_8 FILLER_69_399 ();
 sg13g2_fill_2 FILLER_69_406 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_4 FILLER_70_21 ();
 sg13g2_fill_1 FILLER_70_25 ();
 sg13g2_fill_2 FILLER_70_36 ();
 sg13g2_decap_4 FILLER_70_55 ();
 sg13g2_fill_2 FILLER_70_69 ();
 sg13g2_fill_1 FILLER_70_109 ();
 sg13g2_fill_2 FILLER_70_146 ();
 sg13g2_fill_1 FILLER_70_193 ();
 sg13g2_fill_2 FILLER_70_208 ();
 sg13g2_fill_1 FILLER_70_210 ();
 sg13g2_fill_2 FILLER_70_268 ();
 sg13g2_fill_2 FILLER_70_275 ();
 sg13g2_fill_2 FILLER_70_297 ();
 sg13g2_fill_1 FILLER_70_299 ();
 sg13g2_fill_1 FILLER_70_347 ();
 sg13g2_fill_2 FILLER_70_367 ();
 sg13g2_fill_1 FILLER_70_369 ();
 sg13g2_decap_8 FILLER_70_383 ();
 sg13g2_decap_8 FILLER_70_390 ();
 sg13g2_decap_8 FILLER_70_397 ();
 sg13g2_decap_4 FILLER_70_404 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_fill_1 FILLER_71_14 ();
 sg13g2_fill_1 FILLER_71_46 ();
 sg13g2_fill_2 FILLER_71_73 ();
 sg13g2_fill_2 FILLER_71_89 ();
 sg13g2_fill_1 FILLER_71_91 ();
 sg13g2_fill_2 FILLER_71_118 ();
 sg13g2_decap_4 FILLER_71_147 ();
 sg13g2_fill_2 FILLER_71_151 ();
 sg13g2_fill_2 FILLER_71_221 ();
 sg13g2_fill_1 FILLER_71_223 ();
 sg13g2_fill_2 FILLER_71_256 ();
 sg13g2_fill_2 FILLER_71_284 ();
 sg13g2_fill_1 FILLER_71_286 ();
 sg13g2_fill_2 FILLER_71_317 ();
 sg13g2_decap_8 FILLER_71_386 ();
 sg13g2_decap_8 FILLER_71_393 ();
 sg13g2_decap_8 FILLER_71_400 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_fill_1 FILLER_72_7 ();
 sg13g2_fill_2 FILLER_72_44 ();
 sg13g2_fill_1 FILLER_72_46 ();
 sg13g2_fill_1 FILLER_72_66 ();
 sg13g2_fill_1 FILLER_72_108 ();
 sg13g2_decap_8 FILLER_72_145 ();
 sg13g2_decap_4 FILLER_72_152 ();
 sg13g2_fill_2 FILLER_72_156 ();
 sg13g2_decap_8 FILLER_72_223 ();
 sg13g2_fill_2 FILLER_72_230 ();
 sg13g2_fill_1 FILLER_72_243 ();
 sg13g2_decap_4 FILLER_72_275 ();
 sg13g2_fill_1 FILLER_72_315 ();
 sg13g2_fill_2 FILLER_72_342 ();
 sg13g2_fill_1 FILLER_72_344 ();
 sg13g2_decap_8 FILLER_72_381 ();
 sg13g2_decap_8 FILLER_72_388 ();
 sg13g2_decap_8 FILLER_72_395 ();
 sg13g2_decap_8 FILLER_72_402 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_4 FILLER_73_7 ();
 sg13g2_fill_2 FILLER_73_41 ();
 sg13g2_fill_1 FILLER_73_43 ();
 sg13g2_fill_2 FILLER_73_70 ();
 sg13g2_fill_1 FILLER_73_154 ();
 sg13g2_fill_2 FILLER_73_185 ();
 sg13g2_fill_1 FILLER_73_187 ();
 sg13g2_decap_8 FILLER_73_227 ();
 sg13g2_fill_2 FILLER_73_234 ();
 sg13g2_fill_1 FILLER_73_236 ();
 sg13g2_decap_8 FILLER_73_242 ();
 sg13g2_decap_4 FILLER_73_249 ();
 sg13g2_fill_1 FILLER_73_253 ();
 sg13g2_decap_4 FILLER_73_262 ();
 sg13g2_fill_2 FILLER_73_266 ();
 sg13g2_decap_8 FILLER_73_273 ();
 sg13g2_decap_8 FILLER_73_280 ();
 sg13g2_fill_2 FILLER_73_287 ();
 sg13g2_fill_1 FILLER_73_289 ();
 sg13g2_fill_1 FILLER_73_294 ();
 sg13g2_fill_2 FILLER_73_318 ();
 sg13g2_decap_8 FILLER_73_381 ();
 sg13g2_decap_8 FILLER_73_388 ();
 sg13g2_decap_8 FILLER_73_395 ();
 sg13g2_decap_8 FILLER_73_402 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_4 FILLER_74_7 ();
 sg13g2_fill_2 FILLER_74_11 ();
 sg13g2_fill_2 FILLER_74_112 ();
 sg13g2_fill_1 FILLER_74_124 ();
 sg13g2_decap_8 FILLER_74_142 ();
 sg13g2_fill_2 FILLER_74_149 ();
 sg13g2_fill_1 FILLER_74_151 ();
 sg13g2_fill_2 FILLER_74_224 ();
 sg13g2_decap_8 FILLER_74_247 ();
 sg13g2_decap_8 FILLER_74_280 ();
 sg13g2_decap_8 FILLER_74_287 ();
 sg13g2_fill_2 FILLER_74_336 ();
 sg13g2_fill_1 FILLER_74_338 ();
 sg13g2_fill_2 FILLER_74_349 ();
 sg13g2_fill_1 FILLER_74_351 ();
 sg13g2_decap_8 FILLER_74_378 ();
 sg13g2_decap_8 FILLER_74_385 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_decap_8 FILLER_74_399 ();
 sg13g2_fill_2 FILLER_74_406 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_4 FILLER_75_14 ();
 sg13g2_fill_2 FILLER_75_18 ();
 sg13g2_decap_8 FILLER_75_128 ();
 sg13g2_decap_8 FILLER_75_135 ();
 sg13g2_decap_8 FILLER_75_142 ();
 sg13g2_decap_4 FILLER_75_149 ();
 sg13g2_fill_2 FILLER_75_153 ();
 sg13g2_decap_8 FILLER_75_225 ();
 sg13g2_decap_8 FILLER_75_239 ();
 sg13g2_fill_2 FILLER_75_246 ();
 sg13g2_fill_1 FILLER_75_248 ();
 sg13g2_fill_2 FILLER_75_253 ();
 sg13g2_fill_1 FILLER_75_255 ();
 sg13g2_decap_8 FILLER_75_274 ();
 sg13g2_decap_8 FILLER_75_281 ();
 sg13g2_fill_2 FILLER_75_288 ();
 sg13g2_decap_4 FILLER_75_321 ();
 sg13g2_fill_2 FILLER_75_325 ();
 sg13g2_fill_1 FILLER_75_335 ();
 sg13g2_fill_2 FILLER_75_350 ();
 sg13g2_decap_8 FILLER_75_383 ();
 sg13g2_decap_8 FILLER_75_390 ();
 sg13g2_decap_8 FILLER_75_397 ();
 sg13g2_decap_4 FILLER_75_404 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_4 FILLER_76_21 ();
 sg13g2_fill_2 FILLER_76_44 ();
 sg13g2_fill_2 FILLER_76_83 ();
 sg13g2_fill_1 FILLER_76_85 ();
 sg13g2_decap_8 FILLER_76_131 ();
 sg13g2_decap_8 FILLER_76_138 ();
 sg13g2_decap_8 FILLER_76_145 ();
 sg13g2_decap_8 FILLER_76_152 ();
 sg13g2_decap_4 FILLER_76_159 ();
 sg13g2_fill_1 FILLER_76_163 ();
 sg13g2_fill_1 FILLER_76_191 ();
 sg13g2_decap_8 FILLER_76_218 ();
 sg13g2_fill_2 FILLER_76_241 ();
 sg13g2_decap_8 FILLER_76_383 ();
 sg13g2_decap_8 FILLER_76_390 ();
 sg13g2_decap_8 FILLER_76_397 ();
 sg13g2_decap_4 FILLER_76_404 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_7 ();
 sg13g2_fill_2 FILLER_77_49 ();
 sg13g2_fill_1 FILLER_77_51 ();
 sg13g2_fill_2 FILLER_77_62 ();
 sg13g2_fill_1 FILLER_77_64 ();
 sg13g2_fill_1 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_fill_2 FILLER_77_168 ();
 sg13g2_fill_1 FILLER_77_170 ();
 sg13g2_decap_8 FILLER_77_215 ();
 sg13g2_decap_8 FILLER_77_222 ();
 sg13g2_fill_2 FILLER_77_229 ();
 sg13g2_fill_2 FILLER_77_261 ();
 sg13g2_fill_1 FILLER_77_263 ();
 sg13g2_fill_2 FILLER_77_279 ();
 sg13g2_fill_2 FILLER_77_343 ();
 sg13g2_fill_1 FILLER_77_345 ();
 sg13g2_decap_8 FILLER_77_381 ();
 sg13g2_decap_8 FILLER_77_388 ();
 sg13g2_decap_8 FILLER_77_395 ();
 sg13g2_decap_8 FILLER_77_402 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_4 FILLER_78_14 ();
 sg13g2_fill_2 FILLER_78_18 ();
 sg13g2_decap_8 FILLER_78_124 ();
 sg13g2_decap_8 FILLER_78_131 ();
 sg13g2_decap_8 FILLER_78_138 ();
 sg13g2_decap_8 FILLER_78_145 ();
 sg13g2_decap_8 FILLER_78_152 ();
 sg13g2_decap_8 FILLER_78_159 ();
 sg13g2_decap_8 FILLER_78_166 ();
 sg13g2_fill_2 FILLER_78_173 ();
 sg13g2_fill_1 FILLER_78_175 ();
 sg13g2_fill_2 FILLER_78_189 ();
 sg13g2_fill_1 FILLER_78_191 ();
 sg13g2_decap_8 FILLER_78_222 ();
 sg13g2_decap_8 FILLER_78_229 ();
 sg13g2_fill_2 FILLER_78_236 ();
 sg13g2_decap_8 FILLER_78_269 ();
 sg13g2_decap_8 FILLER_78_276 ();
 sg13g2_fill_2 FILLER_78_283 ();
 sg13g2_fill_1 FILLER_78_285 ();
 sg13g2_decap_8 FILLER_78_385 ();
 sg13g2_decap_8 FILLER_78_392 ();
 sg13g2_decap_8 FILLER_78_399 ();
 sg13g2_fill_2 FILLER_78_406 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_9 ();
 sg13g2_fill_2 FILLER_79_72 ();
 sg13g2_fill_1 FILLER_79_74 ();
 sg13g2_fill_2 FILLER_79_85 ();
 sg13g2_fill_1 FILLER_79_87 ();
 sg13g2_fill_2 FILLER_79_97 ();
 sg13g2_fill_1 FILLER_79_108 ();
 sg13g2_decap_8 FILLER_79_113 ();
 sg13g2_decap_8 FILLER_79_120 ();
 sg13g2_decap_8 FILLER_79_127 ();
 sg13g2_decap_8 FILLER_79_134 ();
 sg13g2_decap_8 FILLER_79_141 ();
 sg13g2_decap_8 FILLER_79_148 ();
 sg13g2_decap_8 FILLER_79_155 ();
 sg13g2_decap_8 FILLER_79_162 ();
 sg13g2_decap_8 FILLER_79_169 ();
 sg13g2_decap_4 FILLER_79_176 ();
 sg13g2_decap_8 FILLER_79_219 ();
 sg13g2_decap_8 FILLER_79_226 ();
 sg13g2_decap_8 FILLER_79_233 ();
 sg13g2_decap_8 FILLER_79_266 ();
 sg13g2_decap_8 FILLER_79_273 ();
 sg13g2_decap_8 FILLER_79_280 ();
 sg13g2_fill_2 FILLER_79_300 ();
 sg13g2_fill_2 FILLER_79_321 ();
 sg13g2_fill_1 FILLER_79_323 ();
 sg13g2_decap_8 FILLER_79_378 ();
 sg13g2_decap_8 FILLER_79_385 ();
 sg13g2_decap_8 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_fill_2 FILLER_79_406 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_4 FILLER_80_7 ();
 sg13g2_fill_2 FILLER_80_58 ();
 sg13g2_fill_1 FILLER_80_60 ();
 sg13g2_fill_2 FILLER_80_83 ();
 sg13g2_fill_2 FILLER_80_102 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_4 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_195 ();
 sg13g2_decap_8 FILLER_80_202 ();
 sg13g2_decap_8 FILLER_80_209 ();
 sg13g2_decap_8 FILLER_80_216 ();
 sg13g2_decap_8 FILLER_80_223 ();
 sg13g2_decap_8 FILLER_80_230 ();
 sg13g2_decap_8 FILLER_80_237 ();
 sg13g2_decap_8 FILLER_80_244 ();
 sg13g2_decap_8 FILLER_80_255 ();
 sg13g2_decap_8 FILLER_80_262 ();
 sg13g2_decap_8 FILLER_80_269 ();
 sg13g2_decap_8 FILLER_80_276 ();
 sg13g2_decap_8 FILLER_80_283 ();
 sg13g2_decap_8 FILLER_80_290 ();
 sg13g2_fill_2 FILLER_80_319 ();
 sg13g2_fill_1 FILLER_80_321 ();
 sg13g2_decap_8 FILLER_80_368 ();
 sg13g2_decap_8 FILLER_80_375 ();
 sg13g2_decap_8 FILLER_80_382 ();
 sg13g2_decap_8 FILLER_80_389 ();
 sg13g2_decap_8 FILLER_80_396 ();
 sg13g2_decap_4 FILLER_80_403 ();
 sg13g2_fill_2 FILLER_80_407 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net8;
 assign uio_out[0] = net9;
 assign uio_out[1] = net10;
 assign uio_out[2] = net11;
 assign uio_out[3] = net12;
 assign uio_out[4] = net13;
 assign uio_out[5] = net14;
 assign uio_out[6] = net15;
 assign uio_out[7] = net16;
endmodule

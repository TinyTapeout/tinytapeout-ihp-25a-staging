module tt_um_rejunity_decoder (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net1;
 wire net2;
 wire net3;

 sg13g2_inv_1 _0510_ (.Y(_0129_),
    .A(net262));
 sg13g2_inv_1 _0511_ (.Y(_0139_),
    .A(net275));
 sg13g2_inv_1 _0512_ (.Y(_0150_),
    .A(net286));
 sg13g2_inv_1 _0513_ (.Y(_0161_),
    .A(net292));
 sg13g2_inv_2 _0514_ (.Y(_0172_),
    .A(net303));
 sg13g2_inv_1 _0515_ (.Y(_0182_),
    .A(net264));
 sg13g2_inv_1 _0516_ (.Y(_0193_),
    .A(net259));
 sg13g2_inv_2 _0517_ (.Y(_0204_),
    .A(net307));
 sg13g2_nor2_2 _0518_ (.A(_0204_),
    .B(net2),
    .Y(_0215_));
 sg13g2_nand2b_2 _0519_ (.Y(_0226_),
    .B(net307),
    .A_N(net2));
 sg13g2_nor2_2 _0520_ (.A(net278),
    .B(net288),
    .Y(_0237_));
 sg13g2_nand2_2 _0521_ (.Y(_0248_),
    .A(net255),
    .B(net249));
 sg13g2_and2_2 _0522_ (.A(net305),
    .B(net299),
    .X(_0258_));
 sg13g2_nand2_1 _0523_ (.Y(_0269_),
    .A(net303),
    .B(net297));
 sg13g2_nor2_2 _0524_ (.A(net292),
    .B(net298),
    .Y(_0280_));
 sg13g2_or2_2 _0525_ (.X(_0291_),
    .B(net299),
    .A(net293));
 sg13g2_nor2_2 _0526_ (.A(net291),
    .B(net302),
    .Y(_0301_));
 sg13g2_a21oi_2 _0527_ (.B1(net295),
    .Y(_0311_),
    .A2(net301),
    .A1(net306));
 sg13g2_a21o_2 _0528_ (.A2(net298),
    .A1(net302),
    .B1(net291),
    .X(_0322_));
 sg13g2_nor2_1 _0529_ (.A(net287),
    .B(net294),
    .Y(_0333_));
 sg13g2_or2_2 _0530_ (.X(_0343_),
    .B(net294),
    .A(net287));
 sg13g2_nor2_1 _0531_ (.A(_0258_),
    .B(net241),
    .Y(_0354_));
 sg13g2_nand2_1 _0532_ (.Y(_0365_),
    .A(_0269_),
    .B(net242));
 sg13g2_nand2_1 _0533_ (.Y(_0376_),
    .A(_0237_),
    .B(_0311_));
 sg13g2_nand2_1 _0534_ (.Y(_0387_),
    .A(net266),
    .B(_0376_));
 sg13g2_nor2_2 _0535_ (.A(net261),
    .B(net258),
    .Y(_0398_));
 sg13g2_nand2_2 _0536_ (.Y(_0407_),
    .A(net257),
    .B(net243));
 sg13g2_a21oi_2 _0537_ (.B1(_0226_),
    .Y(_0418_),
    .A2(net240),
    .A1(_0387_));
 sg13g2_and2_1 _0538_ (.A(net290),
    .B(net297),
    .X(_0428_));
 sg13g2_nand2_2 _0539_ (.Y(_0439_),
    .A(net293),
    .B(net299));
 sg13g2_and3_2 _0540_ (.X(_0450_),
    .A(net294),
    .B(net1),
    .C(net300));
 sg13g2_nand4_1 _0541_ (.B(net296),
    .C(net304),
    .A(net285),
    .Y(_0461_),
    .D(net301));
 sg13g2_and2_1 _0542_ (.A(net253),
    .B(_0461_),
    .X(_0466_));
 sg13g2_nor2_2 _0543_ (.A(net279),
    .B(net248),
    .Y(_0467_));
 sg13g2_nand2_2 _0544_ (.Y(_0468_),
    .A(net256),
    .B(net272));
 sg13g2_nand2_1 _0545_ (.Y(_0469_),
    .A(net267),
    .B(_0466_));
 sg13g2_and2_1 _0546_ (.A(net285),
    .B(net290),
    .X(_0470_));
 sg13g2_nand2_2 _0547_ (.Y(_0471_),
    .A(net284),
    .B(net291));
 sg13g2_nor2_2 _0548_ (.A(net276),
    .B(_0470_),
    .Y(_0472_));
 sg13g2_nor2_1 _0549_ (.A(net267),
    .B(_0472_),
    .Y(_0473_));
 sg13g2_o21ai_1 _0550_ (.B1(net245),
    .Y(_0474_),
    .A1(net276),
    .A2(net239));
 sg13g2_a21oi_1 _0551_ (.A1(net295),
    .A2(net301),
    .Y(_0475_),
    .B1(net289));
 sg13g2_nand2_2 _0552_ (.Y(_0476_),
    .A(net250),
    .B(_0439_));
 sg13g2_nor2_2 _0553_ (.A(net279),
    .B(net271),
    .Y(_0477_));
 sg13g2_nand2_1 _0554_ (.Y(_0478_),
    .A(net255),
    .B(net238));
 sg13g2_nand2_1 _0555_ (.Y(_0479_),
    .A(net238),
    .B(net237));
 sg13g2_nand3_1 _0556_ (.B(_0469_),
    .C(_0474_),
    .A(net259),
    .Y(_0480_));
 sg13g2_o21ai_1 _0557_ (.B1(net261),
    .Y(_0481_),
    .A1(net260),
    .A2(_0479_));
 sg13g2_nor2_1 _0558_ (.A(net257),
    .B(net243),
    .Y(_0482_));
 sg13g2_nand2_2 _0559_ (.Y(_0483_),
    .A(net262),
    .B(net259));
 sg13g2_nand3_1 _0560_ (.B(_0480_),
    .C(_0481_),
    .A(_0418_),
    .Y(_0484_));
 sg13g2_nand2_1 _0561_ (.Y(_0485_),
    .A(_0237_),
    .B(_0280_));
 sg13g2_a21oi_1 _0562_ (.A1(_0237_),
    .A2(_0280_),
    .Y(_0486_),
    .B1(net246));
 sg13g2_a21o_1 _0563_ (.A2(_0486_),
    .A1(net258),
    .B1(net231),
    .X(_0487_));
 sg13g2_o21ai_1 _0564_ (.B1(net279),
    .Y(_0488_),
    .A1(_0258_),
    .A2(net241));
 sg13g2_nand2_2 _0565_ (.Y(_0489_),
    .A(net262),
    .B(net268));
 sg13g2_nor2_2 _0566_ (.A(net256),
    .B(net248),
    .Y(_0490_));
 sg13g2_nand2_2 _0567_ (.Y(_0491_),
    .A(net279),
    .B(net271));
 sg13g2_nor2_2 _0568_ (.A(net247),
    .B(_0488_),
    .Y(_0492_));
 sg13g2_nand2_1 _0569_ (.Y(_0493_),
    .A(net261),
    .B(_0492_));
 sg13g2_and2_2 _0570_ (.A(net307),
    .B(net2),
    .X(_0494_));
 sg13g2_nand2_2 _0571_ (.Y(_0495_),
    .A(net307),
    .B(net2));
 sg13g2_nand3_1 _0572_ (.B(_0493_),
    .C(_0494_),
    .A(_0487_),
    .Y(_0496_));
 sg13g2_nor2_2 _0573_ (.A(net261),
    .B(net244),
    .Y(_0497_));
 sg13g2_nand2_2 _0574_ (.Y(_0498_),
    .A(net257),
    .B(net258));
 sg13g2_a21oi_1 _0575_ (.A1(net267),
    .A2(_0248_),
    .Y(_0499_),
    .B1(_0498_));
 sg13g2_and2_2 _0576_ (.A(net278),
    .B(net288),
    .X(_0500_));
 sg13g2_nand2_2 _0577_ (.Y(_0501_),
    .A(net280),
    .B(net289));
 sg13g2_nand2_1 _0578_ (.Y(_0502_),
    .A(net276),
    .B(net239));
 sg13g2_nor2_2 _0579_ (.A(_0439_),
    .B(_0501_),
    .Y(_0503_));
 sg13g2_nand2_2 _0580_ (.Y(_0504_),
    .A(net261),
    .B(net244));
 sg13g2_nor2_1 _0581_ (.A(net258),
    .B(_0489_),
    .Y(_0505_));
 sg13g2_nand2b_2 _0582_ (.Y(_0506_),
    .B(net243),
    .A_N(_0489_));
 sg13g2_and2_1 _0583_ (.A(_0503_),
    .B(_0505_),
    .X(_0507_));
 sg13g2_nand2_1 _0584_ (.Y(_0508_),
    .A(_0503_),
    .B(_0505_));
 sg13g2_o21ai_1 _0585_ (.B1(_0204_),
    .Y(_0509_),
    .A1(_0499_),
    .A2(_0507_));
 sg13g2_nand3_1 _0586_ (.B(_0496_),
    .C(_0509_),
    .A(_0484_),
    .Y(uo_out[0]));
 sg13g2_nor2_1 _0587_ (.A(net284),
    .B(_0450_),
    .Y(_0000_));
 sg13g2_or2_1 _0588_ (.X(_0001_),
    .B(_0450_),
    .A(net284));
 sg13g2_nand2_1 _0589_ (.Y(_0002_),
    .A(_0471_),
    .B(_0001_));
 sg13g2_nand3_1 _0590_ (.B(_0471_),
    .C(_0001_),
    .A(net278),
    .Y(_0003_));
 sg13g2_nor2_1 _0591_ (.A(net277),
    .B(net249),
    .Y(_0004_));
 sg13g2_nand2_1 _0592_ (.Y(_0005_),
    .A(net255),
    .B(net288));
 sg13g2_nor2_1 _0593_ (.A(net306),
    .B(net300),
    .Y(_0006_));
 sg13g2_or2_2 _0594_ (.X(_0007_),
    .B(net300),
    .A(net306));
 sg13g2_nand2_2 _0595_ (.Y(_0008_),
    .A(net295),
    .B(_0007_));
 sg13g2_inv_1 _0596_ (.Y(_0009_),
    .A(_0008_));
 sg13g2_o21ai_1 _0597_ (.B1(_0003_),
    .Y(_0010_),
    .A1(_0005_),
    .A2(_0009_));
 sg13g2_nor2_2 _0598_ (.A(net251),
    .B(_0280_),
    .Y(_0011_));
 sg13g2_nand2_2 _0599_ (.Y(_0012_),
    .A(net288),
    .B(_0291_));
 sg13g2_nor3_2 _0600_ (.A(net295),
    .B(net306),
    .C(net300),
    .Y(_0013_));
 sg13g2_or3_2 _0601_ (.A(net293),
    .B(net306),
    .C(net299),
    .X(_0014_));
 sg13g2_nand2_2 _0602_ (.Y(_0015_),
    .A(net289),
    .B(_0014_));
 sg13g2_nor2_2 _0603_ (.A(net256),
    .B(net271),
    .Y(_0016_));
 sg13g2_nand2_2 _0604_ (.Y(_0017_),
    .A(net275),
    .B(net245));
 sg13g2_nor2_1 _0605_ (.A(net242),
    .B(_0017_),
    .Y(_0018_));
 sg13g2_a21oi_2 _0606_ (.B1(net289),
    .Y(_0019_),
    .A2(_0007_),
    .A1(net295));
 sg13g2_nor4_1 _0607_ (.A(net280),
    .B(net269),
    .C(_0011_),
    .D(_0019_),
    .Y(_0020_));
 sg13g2_a221oi_1 _0608_ (.B2(_0018_),
    .C1(_0020_),
    .B1(_0015_),
    .A1(net269),
    .Y(_0021_),
    .A2(_0010_));
 sg13g2_nor2_1 _0609_ (.A(_0439_),
    .B(_0005_),
    .Y(_0022_));
 sg13g2_nor2_1 _0610_ (.A(_0450_),
    .B(_0012_),
    .Y(_0023_));
 sg13g2_a22oi_1 _0611_ (.Y(_0024_),
    .B1(_0023_),
    .B2(_0016_),
    .A2(_0022_),
    .A1(net271));
 sg13g2_nor2_2 _0612_ (.A(net250),
    .B(_0311_),
    .Y(_0025_));
 sg13g2_inv_1 _0613_ (.Y(_0026_),
    .A(_0025_));
 sg13g2_o21ai_1 _0614_ (.B1(_0365_),
    .Y(_0027_),
    .A1(net250),
    .A2(_0008_));
 sg13g2_a22oi_1 _0615_ (.Y(_0028_),
    .B1(_0027_),
    .B2(_0490_),
    .A2(_0025_),
    .A1(net236));
 sg13g2_a21oi_1 _0616_ (.A1(_0024_),
    .A2(_0028_),
    .Y(_0029_),
    .B1(_0504_));
 sg13g2_nor2_1 _0617_ (.A(_0248_),
    .B(_0311_),
    .Y(_0030_));
 sg13g2_nor2_1 _0618_ (.A(net269),
    .B(_0030_),
    .Y(_0031_));
 sg13g2_nor3_1 _0619_ (.A(net278),
    .B(net238),
    .C(_0025_),
    .Y(_0032_));
 sg13g2_o21ai_1 _0620_ (.B1(net232),
    .Y(_0033_),
    .A1(net247),
    .A2(_0032_));
 sg13g2_a21oi_1 _0621_ (.A1(_0003_),
    .A2(_0031_),
    .Y(_0034_),
    .B1(_0033_));
 sg13g2_nand3_1 _0622_ (.B(_0490_),
    .C(_0015_),
    .A(_0343_),
    .Y(_0035_));
 sg13g2_nor2_1 _0623_ (.A(_0476_),
    .B(_0013_),
    .Y(_0036_));
 sg13g2_nor3_1 _0624_ (.A(_0476_),
    .B(_0013_),
    .C(_0017_),
    .Y(_0037_));
 sg13g2_nor2_2 _0625_ (.A(net300),
    .B(net241),
    .Y(_0038_));
 sg13g2_a221oi_1 _0626_ (.B2(net236),
    .C1(_0037_),
    .B1(_0038_),
    .A1(_0467_),
    .Y(_0039_),
    .A2(_0019_));
 sg13g2_a21oi_1 _0627_ (.A1(_0035_),
    .A2(_0039_),
    .Y(_0040_),
    .B1(_0498_));
 sg13g2_nor3_1 _0628_ (.A(_0029_),
    .B(_0034_),
    .C(_0040_),
    .Y(_0041_));
 sg13g2_o21ai_1 _0629_ (.B1(_0041_),
    .Y(_0042_),
    .A1(_0407_),
    .A2(_0021_));
 sg13g2_nand2_1 _0630_ (.Y(_0043_),
    .A(_0475_),
    .B(_0490_));
 sg13g2_nor2_1 _0631_ (.A(net249),
    .B(_0428_),
    .Y(_0044_));
 sg13g2_a22oi_1 _0632_ (.Y(_0045_),
    .B1(_0500_),
    .B2(_0439_),
    .A2(_0476_),
    .A1(_0472_));
 sg13g2_nor2b_2 _0633_ (.A(net288),
    .B_N(net278),
    .Y(_0046_));
 sg13g2_nand2_1 _0634_ (.Y(_0047_),
    .A(net278),
    .B(net250));
 sg13g2_o21ai_1 _0635_ (.B1(_0043_),
    .Y(_0048_),
    .A1(net272),
    .A2(_0045_));
 sg13g2_nand2_1 _0636_ (.Y(_0049_),
    .A(net253),
    .B(_0012_));
 sg13g2_nand3_1 _0637_ (.B(_0343_),
    .C(_0012_),
    .A(net255),
    .Y(_0050_));
 sg13g2_nor2_2 _0638_ (.A(net254),
    .B(net238),
    .Y(_0051_));
 sg13g2_nand2_1 _0639_ (.Y(_0052_),
    .A(_0471_),
    .B(_0051_));
 sg13g2_nand2_1 _0640_ (.Y(_0053_),
    .A(_0050_),
    .B(_0052_));
 sg13g2_a21oi_1 _0641_ (.A1(net281),
    .A2(net242),
    .Y(_0054_),
    .B1(_0022_));
 sg13g2_nand2_2 _0642_ (.Y(_0055_),
    .A(net272),
    .B(net230));
 sg13g2_nor2_2 _0643_ (.A(net257),
    .B(net264),
    .Y(_0056_));
 sg13g2_nand2_2 _0644_ (.Y(_0057_),
    .A(net243),
    .B(_0056_));
 sg13g2_inv_1 _0645_ (.Y(_0058_),
    .A(_0057_));
 sg13g2_a21oi_1 _0646_ (.A1(_0248_),
    .A2(_0501_),
    .Y(_0059_),
    .B1(_0280_));
 sg13g2_a22oi_1 _0647_ (.Y(_0060_),
    .B1(_0011_),
    .B2(net233),
    .A2(net236),
    .A1(net238));
 sg13g2_nor2_2 _0648_ (.A(net255),
    .B(_0038_),
    .Y(_0061_));
 sg13g2_nor3_1 _0649_ (.A(_0472_),
    .B(_0506_),
    .C(_0061_),
    .Y(_0062_));
 sg13g2_nand3_1 _0650_ (.B(_0439_),
    .C(net235),
    .A(net247),
    .Y(_0063_));
 sg13g2_nand2_1 _0651_ (.Y(_0064_),
    .A(_0060_),
    .B(_0063_));
 sg13g2_nand2_1 _0652_ (.Y(_0065_),
    .A(net272),
    .B(_0054_));
 sg13g2_o21ai_1 _0653_ (.B1(_0065_),
    .Y(_0066_),
    .A1(net272),
    .A2(_0053_));
 sg13g2_a221oi_1 _0654_ (.B2(_0059_),
    .C1(_0062_),
    .B1(_0058_),
    .A1(_0398_),
    .Y(_0067_),
    .A2(_0048_));
 sg13g2_o21ai_1 _0655_ (.B1(_0067_),
    .Y(_0068_),
    .A1(_0498_),
    .A2(_0066_));
 sg13g2_a21oi_1 _0656_ (.A1(net232),
    .A2(_0064_),
    .Y(_0069_),
    .B1(_0068_));
 sg13g2_nor2_1 _0657_ (.A(net238),
    .B(_0491_),
    .Y(_0070_));
 sg13g2_nor2_1 _0658_ (.A(net263),
    .B(_0070_),
    .Y(_0071_));
 sg13g2_nor2_1 _0659_ (.A(net266),
    .B(net258),
    .Y(_0072_));
 sg13g2_o21ai_1 _0660_ (.B1(net278),
    .Y(_0073_),
    .A1(net305),
    .A2(net298));
 sg13g2_o21ai_1 _0661_ (.B1(net277),
    .Y(_0074_),
    .A1(net241),
    .A2(_0007_));
 sg13g2_a21oi_1 _0662_ (.A1(_0072_),
    .A2(_0074_),
    .Y(_0075_),
    .B1(net240));
 sg13g2_a21oi_1 _0663_ (.A1(net237),
    .A2(_0000_),
    .Y(_0076_),
    .B1(_0486_));
 sg13g2_a22oi_1 _0664_ (.Y(_0077_),
    .B1(_0016_),
    .B2(net286),
    .A2(_0488_),
    .A1(net271));
 sg13g2_nor2_1 _0665_ (.A(_0483_),
    .B(_0077_),
    .Y(_0078_));
 sg13g2_a21oi_1 _0666_ (.A1(_0497_),
    .A2(_0076_),
    .Y(_0079_),
    .B1(_0078_));
 sg13g2_o21ai_1 _0667_ (.B1(_0079_),
    .Y(_0080_),
    .A1(_0071_),
    .A2(_0075_));
 sg13g2_a22oi_1 _0668_ (.Y(_0081_),
    .B1(_0080_),
    .B2(_0494_),
    .A2(_0042_),
    .A1(_0215_));
 sg13g2_o21ai_1 _0669_ (.B1(_0081_),
    .Y(uo_out[1]),
    .A1(net308),
    .A2(_0069_));
 sg13g2_nor2b_2 _0670_ (.A(net300),
    .B_N(net286),
    .Y(_0082_));
 sg13g2_nor2b_2 _0671_ (.A(net293),
    .B_N(net299),
    .Y(_0083_));
 sg13g2_nor2b_2 _0672_ (.A(net286),
    .B_N(net299),
    .Y(_0084_));
 sg13g2_nand2_1 _0673_ (.Y(_0085_),
    .A(net250),
    .B(net300));
 sg13g2_nor2b_2 _0674_ (.A(net297),
    .B_N(net290),
    .Y(_0086_));
 sg13g2_or4_2 _0675_ (.A(net242),
    .B(net239),
    .C(_0082_),
    .D(_0084_),
    .X(_0087_));
 sg13g2_xnor2_1 _0676_ (.Y(_0088_),
    .A(net292),
    .B(net298));
 sg13g2_nand2_1 _0677_ (.Y(_0089_),
    .A(net249),
    .B(_0088_));
 sg13g2_nand2_1 _0678_ (.Y(_0090_),
    .A(_0046_),
    .B(_0088_));
 sg13g2_o21ai_1 _0679_ (.B1(_0090_),
    .Y(_0091_),
    .A1(net275),
    .A2(_0087_));
 sg13g2_nand3_1 _0680_ (.B(net231),
    .C(_0091_),
    .A(net265),
    .Y(_0092_));
 sg13g2_a22oi_1 _0681_ (.Y(_0093_),
    .B1(_0088_),
    .B2(net283),
    .A2(_0084_),
    .A1(_0161_));
 sg13g2_nor2_1 _0682_ (.A(net252),
    .B(_0093_),
    .Y(_0094_));
 sg13g2_nand2_1 _0683_ (.Y(_0095_),
    .A(net291),
    .B(_0082_));
 sg13g2_a21oi_1 _0684_ (.A1(_0089_),
    .A2(_0095_),
    .Y(_0096_),
    .B1(net275));
 sg13g2_xor2_1 _0685_ (.B(net258),
    .A(net264),
    .X(_0097_));
 sg13g2_nand2_1 _0686_ (.Y(_0098_),
    .A(net262),
    .B(_0097_));
 sg13g2_o21ai_1 _0687_ (.B1(_0098_),
    .Y(_0099_),
    .A1(net264),
    .A2(_0407_));
 sg13g2_o21ai_1 _0688_ (.B1(_0099_),
    .Y(_0100_),
    .A1(_0094_),
    .A2(_0096_));
 sg13g2_nand2_2 _0689_ (.Y(_0101_),
    .A(_0055_),
    .B(_0057_));
 sg13g2_nor2_1 _0690_ (.A(net252),
    .B(_0087_),
    .Y(_0102_));
 sg13g2_mux2_2 _0691_ (.A0(_0087_),
    .A1(_0093_),
    .S(net252),
    .X(_0103_));
 sg13g2_inv_1 _0692_ (.Y(_0104_),
    .A(_0103_));
 sg13g2_a21o_1 _0693_ (.A2(_0086_),
    .A1(net235),
    .B1(_0091_),
    .X(_0105_));
 sg13g2_and2_1 _0694_ (.A(net257),
    .B(_0097_),
    .X(_0106_));
 sg13g2_a22oi_1 _0695_ (.Y(_0107_),
    .B1(_0105_),
    .B2(_0106_),
    .A2(_0104_),
    .A1(_0101_));
 sg13g2_nand3_1 _0696_ (.B(_0100_),
    .C(_0107_),
    .A(_0092_),
    .Y(_0108_));
 sg13g2_nand2_1 _0697_ (.Y(_0109_),
    .A(net304),
    .B(_0108_));
 sg13g2_a21oi_2 _0698_ (.B1(net277),
    .Y(_0110_),
    .A2(_0014_),
    .A1(net285));
 sg13g2_inv_1 _0699_ (.Y(_0111_),
    .A(_0110_));
 sg13g2_a221oi_1 _0700_ (.B2(_0002_),
    .C1(net267),
    .B1(_0110_),
    .A1(net235),
    .Y(_0112_),
    .A2(_0014_));
 sg13g2_nor2_2 _0701_ (.A(_0501_),
    .B(_0008_),
    .Y(_0113_));
 sg13g2_a22oi_1 _0702_ (.Y(_0114_),
    .B1(net241),
    .B2(net276),
    .A2(_0280_),
    .A1(_0237_));
 sg13g2_o21ai_1 _0703_ (.B1(net267),
    .Y(_0115_),
    .A1(_0113_),
    .A2(_0114_));
 sg13g2_nand2b_1 _0704_ (.Y(_0116_),
    .B(_0115_),
    .A_N(_0112_));
 sg13g2_nor2_1 _0705_ (.A(_0472_),
    .B(_0503_),
    .Y(_0117_));
 sg13g2_nor2_1 _0706_ (.A(net267),
    .B(_0237_),
    .Y(_0118_));
 sg13g2_a21oi_1 _0707_ (.A1(_0074_),
    .A2(_0118_),
    .Y(_0119_),
    .B1(_0504_));
 sg13g2_o21ai_1 _0708_ (.B1(_0119_),
    .Y(_0120_),
    .A1(_0387_),
    .A2(_0117_));
 sg13g2_o21ai_1 _0709_ (.B1(net255),
    .Y(_0121_),
    .A1(_0471_),
    .A2(net234));
 sg13g2_a22oi_1 _0710_ (.Y(_0122_),
    .B1(_0121_),
    .B2(net270),
    .A2(_0061_),
    .A1(_0026_));
 sg13g2_o21ai_1 _0711_ (.B1(net240),
    .Y(_0123_),
    .A1(_0070_),
    .A2(_0122_));
 sg13g2_nand2_1 _0712_ (.Y(_0124_),
    .A(_0461_),
    .B(net237));
 sg13g2_a22oi_1 _0713_ (.Y(_0125_),
    .B1(_0012_),
    .B2(net233),
    .A2(net235),
    .A1(net245));
 sg13g2_a21oi_1 _0714_ (.A1(net246),
    .A2(net235),
    .Y(_0126_),
    .B1(_0492_));
 sg13g2_nand3b_1 _0715_ (.B(_0124_),
    .C(_0125_),
    .Y(_0127_),
    .A_N(_0492_));
 sg13g2_a22oi_1 _0716_ (.Y(_0128_),
    .B1(_0127_),
    .B2(net231),
    .A2(_0116_),
    .A1(net230));
 sg13g2_nand4_1 _0717_ (.B(_0120_),
    .C(_0123_),
    .A(_0494_),
    .Y(_0130_),
    .D(_0128_));
 sg13g2_o21ai_1 _0718_ (.B1(_0130_),
    .Y(uo_out[2]),
    .A1(net307),
    .A2(_0109_));
 sg13g2_nor2_1 _0719_ (.A(_0017_),
    .B(_0038_),
    .Y(_0131_));
 sg13g2_nor2_2 _0720_ (.A(net254),
    .B(_0019_),
    .Y(_0132_));
 sg13g2_nor2_2 _0721_ (.A(net246),
    .B(_0132_),
    .Y(_0133_));
 sg13g2_o21ai_1 _0722_ (.B1(net232),
    .Y(_0134_),
    .A1(_0131_),
    .A2(_0133_));
 sg13g2_nor4_1 _0723_ (.A(net276),
    .B(net268),
    .C(net239),
    .D(_0498_),
    .Y(_0135_));
 sg13g2_o21ai_1 _0724_ (.B1(_0215_),
    .Y(_0136_),
    .A1(_0506_),
    .A2(_0110_));
 sg13g2_nor2_1 _0725_ (.A(_0135_),
    .B(_0136_),
    .Y(_0137_));
 sg13g2_a21oi_1 _0726_ (.A1(net296),
    .A2(net235),
    .Y(_0138_),
    .B1(net247));
 sg13g2_nand2_2 _0727_ (.Y(_0140_),
    .A(net266),
    .B(_0502_));
 sg13g2_nand3b_1 _0728_ (.B(_0140_),
    .C(net260),
    .Y(_0141_),
    .A_N(_0131_));
 sg13g2_o21ai_1 _0729_ (.B1(net269),
    .Y(_0142_),
    .A1(_0439_),
    .A2(_0501_));
 sg13g2_nor2_1 _0730_ (.A(net260),
    .B(_0018_),
    .Y(_0143_));
 sg13g2_nand2_1 _0731_ (.Y(_0144_),
    .A(_0142_),
    .B(_0143_));
 sg13g2_nand4_1 _0732_ (.B(_0495_),
    .C(_0141_),
    .A(net263),
    .Y(_0145_),
    .D(_0144_));
 sg13g2_nor2_1 _0733_ (.A(_0008_),
    .B(_0082_),
    .Y(_0146_));
 sg13g2_nor3_1 _0734_ (.A(net289),
    .B(_0450_),
    .C(_0013_),
    .Y(_0147_));
 sg13g2_nor3_1 _0735_ (.A(_0011_),
    .B(_0017_),
    .C(_0147_),
    .Y(_0148_));
 sg13g2_a22oi_1 _0736_ (.Y(_0149_),
    .B1(_0025_),
    .B2(_0439_),
    .A2(_0019_),
    .A1(_0291_));
 sg13g2_a22oi_1 _0737_ (.Y(_0151_),
    .B1(_0084_),
    .B2(net306),
    .A2(net234),
    .A1(net287));
 sg13g2_a221oi_1 _0738_ (.B2(net305),
    .C1(net294),
    .B1(_0084_),
    .A1(net287),
    .Y(_0152_),
    .A2(_0006_));
 sg13g2_nor2_1 _0739_ (.A(net279),
    .B(_0152_),
    .Y(_0153_));
 sg13g2_a21oi_1 _0740_ (.A1(net281),
    .A2(_0149_),
    .Y(_0154_),
    .B1(_0153_));
 sg13g2_a221oi_1 _0741_ (.B2(net273),
    .C1(_0148_),
    .B1(_0154_),
    .A1(net236),
    .Y(_0155_),
    .A2(_0146_));
 sg13g2_nor2_1 _0742_ (.A(_0504_),
    .B(_0155_),
    .Y(_0156_));
 sg13g2_a21oi_1 _0743_ (.A1(_0476_),
    .A2(_0015_),
    .Y(_0157_),
    .B1(_0450_));
 sg13g2_nand2b_1 _0744_ (.Y(_0158_),
    .B(net236),
    .A_N(_0157_));
 sg13g2_a22oi_1 _0745_ (.Y(_0159_),
    .B1(_0008_),
    .B2(_0011_),
    .A2(_0007_),
    .A1(net242));
 sg13g2_nand3_1 _0746_ (.B(_0016_),
    .C(_0085_),
    .A(_0311_),
    .Y(_0160_));
 sg13g2_o21ai_1 _0747_ (.B1(_0160_),
    .Y(_0162_),
    .A1(_0468_),
    .A2(_0159_));
 sg13g2_nand2b_1 _0748_ (.Y(_0163_),
    .B(_0158_),
    .A_N(_0162_));
 sg13g2_a22oi_1 _0749_ (.Y(_0164_),
    .B1(net238),
    .B2(_0322_),
    .A2(net239),
    .A1(_0269_));
 sg13g2_nor2_1 _0750_ (.A(_0491_),
    .B(_0164_),
    .Y(_0165_));
 sg13g2_o21ai_1 _0751_ (.B1(net240),
    .Y(_0166_),
    .A1(_0163_),
    .A2(_0165_));
 sg13g2_nand2_1 _0752_ (.Y(_0167_),
    .A(net294),
    .B(_0151_));
 sg13g2_mux2_1 _0753_ (.A0(_0157_),
    .A1(_0167_),
    .S(net255),
    .X(_0168_));
 sg13g2_or3_1 _0754_ (.A(net272),
    .B(_0498_),
    .C(_0168_),
    .X(_0169_));
 sg13g2_o21ai_1 _0755_ (.B1(net255),
    .Y(_0170_),
    .A1(_0011_),
    .A2(_0147_));
 sg13g2_nand3_1 _0756_ (.B(_0488_),
    .C(_0170_),
    .A(net271),
    .Y(_0171_));
 sg13g2_nor2_1 _0757_ (.A(net281),
    .B(_0164_),
    .Y(_0173_));
 sg13g2_a21oi_1 _0758_ (.A1(net280),
    .A2(_0146_),
    .Y(_0174_),
    .B1(_0173_));
 sg13g2_o21ai_1 _0759_ (.B1(_0171_),
    .Y(_0175_),
    .A1(net273),
    .A2(_0174_));
 sg13g2_a21oi_1 _0760_ (.A1(_0311_),
    .A2(_0085_),
    .Y(_0176_),
    .B1(net281));
 sg13g2_a21o_1 _0761_ (.A2(_0159_),
    .A1(net280),
    .B1(_0176_),
    .X(_0177_));
 sg13g2_o21ai_1 _0762_ (.B1(net2),
    .Y(_0178_),
    .A1(_0055_),
    .A2(_0177_));
 sg13g2_a21oi_1 _0763_ (.A1(net232),
    .A2(_0175_),
    .Y(_0179_),
    .B1(_0178_));
 sg13g2_nand3_1 _0764_ (.B(_0169_),
    .C(_0179_),
    .A(_0166_),
    .Y(_0180_));
 sg13g2_o21ai_1 _0765_ (.B1(net308),
    .Y(_0181_),
    .A1(_0156_),
    .A2(_0180_));
 sg13g2_a22oi_1 _0766_ (.Y(uo_out[3]),
    .B1(_0145_),
    .B2(_0181_),
    .A2(_0137_),
    .A1(_0134_));
 sg13g2_a21oi_2 _0767_ (.B1(net269),
    .Y(_0183_),
    .A2(_0046_),
    .A1(_0291_));
 sg13g2_a21oi_1 _0768_ (.A1(_0050_),
    .A2(_0138_),
    .Y(_0184_),
    .B1(_0183_));
 sg13g2_and2_1 _0769_ (.A(net240),
    .B(_0184_),
    .X(_0185_));
 sg13g2_nand3_1 _0770_ (.B(net232),
    .C(_0053_),
    .A(net272),
    .Y(_0186_));
 sg13g2_nor2_1 _0771_ (.A(_0506_),
    .B(_0045_),
    .Y(_0187_));
 sg13g2_nand2b_1 _0772_ (.Y(_0188_),
    .B(_0059_),
    .A_N(_0055_));
 sg13g2_nand4_1 _0773_ (.B(net247),
    .C(net238),
    .A(net281),
    .Y(_0189_),
    .D(net230));
 sg13g2_a21oi_1 _0774_ (.A1(_0485_),
    .A2(_0054_),
    .Y(_0190_),
    .B1(_0057_));
 sg13g2_nor4_1 _0775_ (.A(net269),
    .B(_0472_),
    .C(_0483_),
    .D(_0061_),
    .Y(_0191_));
 sg13g2_nor4_1 _0776_ (.A(net308),
    .B(_0187_),
    .C(_0190_),
    .D(_0191_),
    .Y(_0192_));
 sg13g2_nand4_1 _0777_ (.B(_0188_),
    .C(_0189_),
    .A(_0186_),
    .Y(_0194_),
    .D(_0192_));
 sg13g2_o21ai_1 _0778_ (.B1(_0495_),
    .Y(_0195_),
    .A1(_0185_),
    .A2(_0194_));
 sg13g2_xor2_1 _0779_ (.B(net299),
    .A(net305),
    .X(_0196_));
 sg13g2_xnor2_1 _0780_ (.Y(_0197_),
    .A(net302),
    .B(net297));
 sg13g2_a22oi_1 _0781_ (.Y(_0198_),
    .B1(_0197_),
    .B2(net290),
    .A2(_0280_),
    .A1(net302));
 sg13g2_nand2_1 _0782_ (.Y(_0199_),
    .A(net297),
    .B(_0301_));
 sg13g2_nand3b_1 _0783_ (.B(net306),
    .C(net293),
    .Y(_0200_),
    .A_N(net299));
 sg13g2_a22oi_1 _0784_ (.Y(_0201_),
    .B1(_0086_),
    .B2(net302),
    .A2(_0301_),
    .A1(net297));
 sg13g2_a221oi_1 _0785_ (.B2(net302),
    .C1(net249),
    .B1(_0086_),
    .A1(net297),
    .Y(_0202_),
    .A2(_0301_));
 sg13g2_a221oi_1 _0786_ (.B2(net290),
    .C1(net284),
    .B1(_0197_),
    .A1(net302),
    .Y(_0203_),
    .A2(_0280_));
 sg13g2_or2_1 _0787_ (.X(_0205_),
    .B(_0203_),
    .A(_0202_));
 sg13g2_a221oi_1 _0788_ (.B2(_0161_),
    .C1(net249),
    .B1(_0197_),
    .A1(_0172_),
    .Y(_0206_),
    .A2(_0428_));
 sg13g2_a21o_1 _0789_ (.A2(_0201_),
    .A1(net249),
    .B1(_0206_),
    .X(_0207_));
 sg13g2_mux2_1 _0790_ (.A0(_0205_),
    .A1(_0207_),
    .S(net253),
    .X(_0208_));
 sg13g2_a221oi_1 _0791_ (.B2(_0161_),
    .C1(net283),
    .B1(_0197_),
    .A1(_0172_),
    .Y(_0209_),
    .A2(_0428_));
 sg13g2_a21o_1 _0792_ (.A2(_0198_),
    .A1(net283),
    .B1(_0209_),
    .X(_0210_));
 sg13g2_a21oi_1 _0793_ (.A1(net283),
    .A2(_0198_),
    .Y(_0211_),
    .B1(_0209_));
 sg13g2_o21ai_1 _0794_ (.B1(net237),
    .Y(_0212_),
    .A1(_0202_),
    .A2(_0203_));
 sg13g2_o21ai_1 _0795_ (.B1(_0212_),
    .Y(_0213_),
    .A1(_0017_),
    .A2(_0211_));
 sg13g2_a21o_1 _0796_ (.A2(_0208_),
    .A1(net265),
    .B1(_0213_),
    .X(_0214_));
 sg13g2_mux2_1 _0797_ (.A0(_0207_),
    .A1(_0210_),
    .S(net252),
    .X(_0216_));
 sg13g2_mux2_1 _0798_ (.A0(_0208_),
    .A1(_0216_),
    .S(net265),
    .X(_0217_));
 sg13g2_mux2_1 _0799_ (.A0(_0214_),
    .A1(_0217_),
    .S(net257),
    .X(_0218_));
 sg13g2_nor2_1 _0800_ (.A(net244),
    .B(_0218_),
    .Y(_0219_));
 sg13g2_o21ai_1 _0801_ (.B1(net243),
    .Y(_0220_),
    .A1(net262),
    .A2(_0217_));
 sg13g2_and2_1 _0802_ (.A(net244),
    .B(_0218_),
    .X(_0221_));
 sg13g2_nand2_1 _0803_ (.Y(_0222_),
    .A(net257),
    .B(_0214_));
 sg13g2_nand2_1 _0804_ (.Y(_0223_),
    .A(net254),
    .B(_0205_));
 sg13g2_a221oi_1 _0805_ (.B2(_0223_),
    .C1(_0489_),
    .B1(_0073_),
    .A1(net277),
    .Y(_0224_),
    .A2(_0365_));
 sg13g2_nand2b_1 _0806_ (.Y(_0225_),
    .B(net258),
    .A_N(_0224_));
 sg13g2_a221oi_1 _0807_ (.B2(_0056_),
    .C1(_0225_),
    .B1(_0216_),
    .A1(_0129_),
    .Y(_0227_),
    .A2(_0214_));
 sg13g2_or4_1 _0808_ (.A(_0495_),
    .B(_0219_),
    .C(_0221_),
    .D(_0227_),
    .X(_0228_));
 sg13g2_a21oi_1 _0809_ (.A1(net276),
    .A2(net241),
    .Y(_0229_),
    .B1(_0466_));
 sg13g2_nor3_1 _0810_ (.A(net268),
    .B(_0503_),
    .C(_0229_),
    .Y(_0230_));
 sg13g2_nor3_2 _0811_ (.A(_0280_),
    .B(_0450_),
    .C(_0047_),
    .Y(_0231_));
 sg13g2_nand2_1 _0812_ (.Y(_0232_),
    .A(_0398_),
    .B(_0231_));
 sg13g2_a22oi_1 _0813_ (.Y(_0233_),
    .B1(_0232_),
    .B2(_0418_),
    .A2(_0230_),
    .A1(_0215_));
 sg13g2_a21oi_2 _0814_ (.B1(net268),
    .Y(_0234_),
    .A2(net235),
    .A1(_0322_));
 sg13g2_o21ai_1 _0815_ (.B1(_0234_),
    .Y(_0235_),
    .A1(net276),
    .A2(_0002_));
 sg13g2_nor3_1 _0816_ (.A(net280),
    .B(_0450_),
    .C(_0012_),
    .Y(_0236_));
 sg13g2_o21ai_1 _0817_ (.B1(net230),
    .Y(_0238_),
    .A1(_0142_),
    .A2(_0236_));
 sg13g2_nor2b_1 _0818_ (.A(_0238_),
    .B_N(_0235_),
    .Y(_0239_));
 sg13g2_nor2_1 _0819_ (.A(net270),
    .B(_0061_),
    .Y(_0240_));
 sg13g2_o21ai_1 _0820_ (.B1(_0240_),
    .Y(_0241_),
    .A1(net280),
    .A2(_0027_));
 sg13g2_o21ai_1 _0821_ (.B1(_0133_),
    .Y(_0242_),
    .A1(net280),
    .A2(_0036_));
 sg13g2_a21oi_1 _0822_ (.A1(_0241_),
    .A2(_0242_),
    .Y(_0243_),
    .B1(_0483_));
 sg13g2_nand3_1 _0823_ (.B(net233),
    .C(_0015_),
    .A(net241),
    .Y(_0244_));
 sg13g2_a22oi_1 _0824_ (.Y(_0245_),
    .B1(_0012_),
    .B2(_0016_),
    .A2(_0008_),
    .A1(_0490_));
 sg13g2_nor2_1 _0825_ (.A(_0019_),
    .B(_0245_),
    .Y(_0246_));
 sg13g2_a21oi_1 _0826_ (.A1(net236),
    .A2(_0036_),
    .Y(_0247_),
    .B1(_0246_));
 sg13g2_a21oi_1 _0827_ (.A1(_0244_),
    .A2(_0247_),
    .Y(_0249_),
    .B1(_0504_));
 sg13g2_nor4_2 _0828_ (.A(_0233_),
    .B(_0239_),
    .C(_0243_),
    .Y(_0250_),
    .D(_0249_));
 sg13g2_a21oi_1 _0829_ (.A1(_0195_),
    .A2(_0228_),
    .Y(uo_out[4]),
    .B1(_0250_));
 sg13g2_a21o_1 _0830_ (.A2(_0088_),
    .A1(net249),
    .B1(_0172_),
    .X(_0251_));
 sg13g2_o21ai_1 _0831_ (.B1(_0466_),
    .Y(_0252_),
    .A1(net239),
    .A2(_0251_));
 sg13g2_a21o_1 _0832_ (.A2(_0093_),
    .A1(net303),
    .B1(net253),
    .X(_0253_));
 sg13g2_nand3_1 _0833_ (.B(_0252_),
    .C(_0253_),
    .A(net245),
    .Y(_0254_));
 sg13g2_nand2_1 _0834_ (.Y(_0255_),
    .A(net304),
    .B(_0103_));
 sg13g2_o21ai_1 _0835_ (.B1(net257),
    .Y(_0256_),
    .A1(_0254_),
    .A2(_0255_));
 sg13g2_a21oi_1 _0836_ (.A1(_0254_),
    .A2(_0255_),
    .Y(_0257_),
    .B1(_0256_));
 sg13g2_nand4_1 _0837_ (.B(net243),
    .C(_0252_),
    .A(net265),
    .Y(_0259_),
    .D(_0253_));
 sg13g2_nand3_1 _0838_ (.B(_0072_),
    .C(_0103_),
    .A(net304),
    .Y(_0260_));
 sg13g2_nand2_1 _0839_ (.Y(_0261_),
    .A(_0259_),
    .B(_0260_));
 sg13g2_nand4_1 _0840_ (.B(_0471_),
    .C(_0490_),
    .A(net304),
    .Y(_0262_),
    .D(_0089_));
 sg13g2_nand3_1 _0841_ (.B(net233),
    .C(_0087_),
    .A(net303),
    .Y(_0263_));
 sg13g2_nand3_1 _0842_ (.B(_0262_),
    .C(_0263_),
    .A(_0254_),
    .Y(_0264_));
 sg13g2_a21oi_1 _0843_ (.A1(net231),
    .A2(_0264_),
    .Y(_0265_),
    .B1(_0261_));
 sg13g2_nand2b_1 _0844_ (.Y(_0266_),
    .B(_0265_),
    .A_N(_0257_));
 sg13g2_a21oi_1 _0845_ (.A1(_0257_),
    .A2(_0261_),
    .Y(_0267_),
    .B1(net307));
 sg13g2_a22oi_1 _0846_ (.Y(_0268_),
    .B1(_0197_),
    .B2(net290),
    .A2(_0301_),
    .A1(net297));
 sg13g2_o21ai_1 _0847_ (.B1(_0200_),
    .Y(_0270_),
    .A1(net293),
    .A2(_0196_));
 sg13g2_o21ai_1 _0848_ (.B1(_0073_),
    .Y(_0271_),
    .A1(net250),
    .A2(_0083_));
 sg13g2_xor2_1 _0849_ (.B(net305),
    .A(net293),
    .X(_0272_));
 sg13g2_xnor2_1 _0850_ (.Y(_0273_),
    .A(net293),
    .B(net305));
 sg13g2_nor2_1 _0851_ (.A(_0500_),
    .B(_0273_),
    .Y(_0274_));
 sg13g2_a22oi_1 _0852_ (.Y(_0275_),
    .B1(_0271_),
    .B2(_0274_),
    .A2(_0270_),
    .A1(_0500_));
 sg13g2_o21ai_1 _0853_ (.B1(_0275_),
    .Y(_0276_),
    .A1(_0248_),
    .A2(_0268_));
 sg13g2_nand2_1 _0854_ (.Y(_0277_),
    .A(net250),
    .B(_0270_));
 sg13g2_o21ai_1 _0855_ (.B1(_0277_),
    .Y(_0278_),
    .A1(net250),
    .A2(_0272_));
 sg13g2_a221oi_1 _0856_ (.B2(_0161_),
    .C1(_0273_),
    .B1(_0084_),
    .A1(net288),
    .Y(_0279_),
    .A2(_0006_));
 sg13g2_and2_1 _0857_ (.A(net236),
    .B(_0279_),
    .X(_0281_));
 sg13g2_a221oi_1 _0858_ (.B2(_0016_),
    .C1(_0281_),
    .B1(_0278_),
    .A1(net271),
    .Y(_0282_),
    .A2(_0276_));
 sg13g2_a22oi_1 _0859_ (.Y(_0283_),
    .B1(_0279_),
    .B2(net278),
    .A2(_0273_),
    .A1(_0237_));
 sg13g2_o21ai_1 _0860_ (.B1(_0283_),
    .Y(_0284_),
    .A1(_0005_),
    .A2(_0268_));
 sg13g2_mux2_1 _0861_ (.A0(_0276_),
    .A1(_0284_),
    .S(net269),
    .X(_0285_));
 sg13g2_a21oi_1 _0862_ (.A1(net263),
    .A2(_0282_),
    .Y(_0286_),
    .B1(_0285_));
 sg13g2_a21oi_1 _0863_ (.A1(net263),
    .A2(_0285_),
    .Y(_0287_),
    .B1(net260));
 sg13g2_nor2b_1 _0864_ (.A(_0286_),
    .B_N(_0287_),
    .Y(_0288_));
 sg13g2_nand2b_1 _0865_ (.Y(_0289_),
    .B(_0497_),
    .A_N(_0282_));
 sg13g2_nor4_1 _0866_ (.A(net305),
    .B(net247),
    .C(_0047_),
    .D(_0088_),
    .Y(_0290_));
 sg13g2_a221oi_1 _0867_ (.B2(net247),
    .C1(_0290_),
    .B1(_0284_),
    .A1(_0467_),
    .Y(_0292_),
    .A2(_0278_));
 sg13g2_o21ai_1 _0868_ (.B1(_0289_),
    .Y(_0293_),
    .A1(_0483_),
    .A2(_0292_));
 sg13g2_o21ai_1 _0869_ (.B1(_0215_),
    .Y(_0294_),
    .A1(_0288_),
    .A2(_0293_));
 sg13g2_o21ai_1 _0870_ (.B1(_0075_),
    .Y(_0295_),
    .A1(net243),
    .A2(_0493_));
 sg13g2_a22oi_1 _0871_ (.Y(_0296_),
    .B1(_0295_),
    .B2(_0494_),
    .A2(_0267_),
    .A1(_0266_));
 sg13g2_nand2_2 _0872_ (.Y(uo_out[5]),
    .A(_0294_),
    .B(_0296_));
 sg13g2_o21ai_1 _0873_ (.B1(_0474_),
    .Y(_0297_),
    .A1(_0468_),
    .A2(net239));
 sg13g2_o21ai_1 _0874_ (.B1(_0493_),
    .Y(_0298_),
    .A1(net261),
    .A2(_0113_));
 sg13g2_a22oi_1 _0875_ (.Y(_0299_),
    .B1(_0298_),
    .B2(_0487_),
    .A2(_0234_),
    .A1(net240));
 sg13g2_a21oi_1 _0876_ (.A1(_0119_),
    .A2(_0297_),
    .Y(_0300_),
    .B1(_0495_));
 sg13g2_or2_1 _0877_ (.X(_0302_),
    .B(_0502_),
    .A(_0489_));
 sg13g2_a21oi_1 _0878_ (.A1(net259),
    .A2(_0302_),
    .Y(_0303_),
    .B1(_0494_));
 sg13g2_nand2_1 _0879_ (.Y(_0304_),
    .A(_0471_),
    .B(net237));
 sg13g2_a22oi_1 _0880_ (.Y(_0305_),
    .B1(_0132_),
    .B2(net261),
    .A2(_0472_),
    .A1(net245));
 sg13g2_nor3_1 _0881_ (.A(_0226_),
    .B(_0056_),
    .C(_0305_),
    .Y(_0306_));
 sg13g2_a221oi_1 _0882_ (.B2(_0508_),
    .C1(_0306_),
    .B1(_0303_),
    .A1(_0299_),
    .Y(uo_out[6]),
    .A2(_0300_));
 sg13g2_a22oi_1 _0883_ (.Y(_0307_),
    .B1(_0461_),
    .B2(_0051_),
    .A2(net242),
    .A1(net254));
 sg13g2_a221oi_1 _0884_ (.B2(net267),
    .C1(net261),
    .B1(_0307_),
    .A1(_0111_),
    .Y(_0308_),
    .A2(_0234_));
 sg13g2_o21ai_1 _0885_ (.B1(net263),
    .Y(_0309_),
    .A1(net241),
    .A2(_0007_));
 sg13g2_nor3_1 _0886_ (.A(_0011_),
    .B(_0017_),
    .C(_0309_),
    .Y(_0310_));
 sg13g2_nor3_1 _0887_ (.A(_0472_),
    .B(_0489_),
    .C(_0132_),
    .Y(_0312_));
 sg13g2_nor3_1 _0888_ (.A(_0308_),
    .B(_0310_),
    .C(_0312_),
    .Y(_0313_));
 sg13g2_nand3_1 _0889_ (.B(net233),
    .C(net234),
    .A(net242),
    .Y(_0314_));
 sg13g2_nand3_1 _0890_ (.B(_0126_),
    .C(_0314_),
    .A(_0479_),
    .Y(_0315_));
 sg13g2_nor3_1 _0891_ (.A(_0468_),
    .B(_0025_),
    .C(_0038_),
    .Y(_0316_));
 sg13g2_a221oi_1 _0892_ (.B2(net270),
    .C1(_0316_),
    .B1(_0113_),
    .A1(net237),
    .Y(_0317_),
    .A2(_0001_));
 sg13g2_nor2_1 _0893_ (.A(_0498_),
    .B(_0317_),
    .Y(_0318_));
 sg13g2_a21oi_1 _0894_ (.A1(net231),
    .A2(_0315_),
    .Y(_0319_),
    .B1(_0318_));
 sg13g2_o21ai_1 _0895_ (.B1(_0319_),
    .Y(_0320_),
    .A1(net260),
    .A2(_0313_));
 sg13g2_mux2_1 _0896_ (.A0(_0237_),
    .A1(_0051_),
    .S(net246),
    .X(_0321_));
 sg13g2_nor3_1 _0897_ (.A(_0483_),
    .B(_0184_),
    .C(_0321_),
    .Y(_0323_));
 sg13g2_nor3_1 _0898_ (.A(_0472_),
    .B(_0503_),
    .C(_0506_),
    .Y(_0324_));
 sg13g2_nor2b_1 _0899_ (.A(_0057_),
    .B_N(_0114_),
    .Y(_0325_));
 sg13g2_o21ai_1 _0900_ (.B1(_0499_),
    .Y(_0326_),
    .A1(net267),
    .A2(_0051_));
 sg13g2_o21ai_1 _0901_ (.B1(_0326_),
    .Y(_0327_),
    .A1(_0407_),
    .A2(_0125_));
 sg13g2_nor4_1 _0902_ (.A(_0323_),
    .B(_0324_),
    .C(_0325_),
    .D(_0327_),
    .Y(_0328_));
 sg13g2_a22oi_1 _0903_ (.Y(_0329_),
    .B1(_0240_),
    .B2(_0376_),
    .A2(_0133_),
    .A1(_0478_));
 sg13g2_nand2_1 _0904_ (.Y(_0330_),
    .A(net276),
    .B(_0011_));
 sg13g2_a21oi_1 _0905_ (.A1(_0478_),
    .A2(_0330_),
    .Y(_0331_),
    .B1(_0057_));
 sg13g2_o21ai_1 _0906_ (.B1(_0505_),
    .Y(_0332_),
    .A1(_0110_),
    .A2(_0113_));
 sg13g2_a221oi_1 _0907_ (.B2(_0001_),
    .C1(_0018_),
    .B1(_0490_),
    .A1(_0354_),
    .Y(_0334_),
    .A2(net233));
 sg13g2_a21oi_1 _0908_ (.A1(_0469_),
    .A2(_0304_),
    .Y(_0335_),
    .B1(_0498_));
 sg13g2_o21ai_1 _0909_ (.B1(_0332_),
    .Y(_0336_),
    .A1(_0407_),
    .A2(_0334_));
 sg13g2_nor3_1 _0910_ (.A(_0331_),
    .B(_0335_),
    .C(_0336_),
    .Y(_0337_));
 sg13g2_o21ai_1 _0911_ (.B1(_0337_),
    .Y(_0338_),
    .A1(_0483_),
    .A2(_0329_));
 sg13g2_a22oi_1 _0912_ (.Y(_0339_),
    .B1(_0338_),
    .B2(_0215_),
    .A2(_0320_),
    .A1(_0494_));
 sg13g2_o21ai_1 _0913_ (.B1(_0339_),
    .Y(uo_out[7]),
    .A1(net307),
    .A2(_0328_));
 sg13g2_and3_1 _0914_ (.X(_0340_),
    .A(net284),
    .B(net302),
    .C(_0083_));
 sg13g2_nand3_1 _0915_ (.B(net305),
    .C(_0083_),
    .A(net286),
    .Y(_0341_));
 sg13g2_nand2_1 _0916_ (.Y(_0342_),
    .A(net290),
    .B(net234));
 sg13g2_nand2_1 _0917_ (.Y(_0344_),
    .A(net284),
    .B(_0342_));
 sg13g2_o21ai_1 _0918_ (.B1(_0439_),
    .Y(_0345_),
    .A1(_0322_),
    .A2(net234));
 sg13g2_a221oi_1 _0919_ (.B2(net251),
    .C1(_0340_),
    .B1(_0345_),
    .A1(net239),
    .Y(_0346_),
    .A2(net234));
 sg13g2_a21oi_1 _0920_ (.A1(net290),
    .A2(_0197_),
    .Y(_0347_),
    .B1(_0083_));
 sg13g2_or2_1 _0921_ (.X(_0348_),
    .B(_0083_),
    .A(_0258_));
 sg13g2_a22oi_1 _0922_ (.Y(_0349_),
    .B1(_0348_),
    .B2(net235),
    .A2(_0347_),
    .A1(_0046_));
 sg13g2_o21ai_1 _0923_ (.B1(_0349_),
    .Y(_0350_),
    .A1(net275),
    .A2(_0346_));
 sg13g2_nand2_1 _0924_ (.Y(_0351_),
    .A(net264),
    .B(_0350_));
 sg13g2_nand2_1 _0925_ (.Y(_0352_),
    .A(_0322_),
    .B(_0019_));
 sg13g2_a21oi_1 _0926_ (.A1(net283),
    .A2(_0347_),
    .Y(_0353_),
    .B1(net277));
 sg13g2_or3_2 _0927_ (.A(_0258_),
    .B(_0301_),
    .C(_0086_),
    .X(_0355_));
 sg13g2_or2_1 _0928_ (.X(_0356_),
    .B(_0086_),
    .A(net234));
 sg13g2_o21ai_1 _0929_ (.B1(_0355_),
    .Y(_0357_),
    .A1(_0082_),
    .A2(_0084_));
 sg13g2_a22oi_1 _0930_ (.Y(_0358_),
    .B1(_0357_),
    .B2(net275),
    .A2(_0353_),
    .A1(_0352_));
 sg13g2_a21oi_1 _0931_ (.A1(net245),
    .A2(_0358_),
    .Y(_0359_),
    .B1(net262));
 sg13g2_nand2_1 _0932_ (.Y(_0360_),
    .A(_0351_),
    .B(_0359_));
 sg13g2_mux2_1 _0933_ (.A0(_0346_),
    .A1(_0357_),
    .S(net252),
    .X(_0361_));
 sg13g2_inv_1 _0934_ (.Y(_0362_),
    .A(_0361_));
 sg13g2_nor3_1 _0935_ (.A(net264),
    .B(_0350_),
    .C(_0362_),
    .Y(_0363_));
 sg13g2_o21ai_1 _0936_ (.B1(net262),
    .Y(_0364_),
    .A1(net245),
    .A2(_0361_));
 sg13g2_o21ai_1 _0937_ (.B1(_0360_),
    .Y(_0366_),
    .A1(_0363_),
    .A2(_0364_));
 sg13g2_a21oi_1 _0938_ (.A1(net245),
    .A2(_0361_),
    .Y(_0367_),
    .B1(_0358_));
 sg13g2_nand2b_1 _0939_ (.Y(_0368_),
    .B(_0359_),
    .A_N(_0367_));
 sg13g2_nor2_1 _0940_ (.A(net254),
    .B(_0352_),
    .Y(_0369_));
 sg13g2_a221oi_1 _0941_ (.B2(_0237_),
    .C1(_0369_),
    .B1(_0356_),
    .A1(_0004_),
    .Y(_0370_),
    .A2(_0345_));
 sg13g2_o21ai_1 _0942_ (.B1(net258),
    .Y(_0371_),
    .A1(_0489_),
    .A2(_0370_));
 sg13g2_a21oi_1 _0943_ (.A1(_0056_),
    .A2(_0350_),
    .Y(_0372_),
    .B1(_0371_));
 sg13g2_a221oi_1 _0944_ (.B2(_0372_),
    .C1(_0226_),
    .B1(_0368_),
    .A1(net243),
    .Y(_0373_),
    .A2(_0366_));
 sg13g2_nor2_1 _0945_ (.A(_0506_),
    .B(_0174_),
    .Y(_0374_));
 sg13g2_nor2_1 _0946_ (.A(_0057_),
    .B(_0177_),
    .Y(_0375_));
 sg13g2_nor2_1 _0947_ (.A(_0374_),
    .B(_0375_),
    .Y(_0377_));
 sg13g2_a21oi_1 _0948_ (.A1(net273),
    .A2(_0168_),
    .Y(_0378_),
    .B1(_0407_));
 sg13g2_o21ai_1 _0949_ (.B1(_0378_),
    .Y(_0379_),
    .A1(net272),
    .A2(_0154_));
 sg13g2_and2_1 _0950_ (.A(net247),
    .B(_0152_),
    .X(_0380_));
 sg13g2_o21ai_1 _0951_ (.B1(_0170_),
    .Y(_0381_),
    .A1(_0477_),
    .A2(_0380_));
 sg13g2_nor2_1 _0952_ (.A(_0468_),
    .B(_0149_),
    .Y(_0382_));
 sg13g2_o21ai_1 _0953_ (.B1(_0381_),
    .Y(_0383_),
    .A1(_0491_),
    .A2(_0167_));
 sg13g2_o21ai_1 _0954_ (.B1(net230),
    .Y(_0384_),
    .A1(_0382_),
    .A2(_0383_));
 sg13g2_o21ai_1 _0955_ (.B1(net231),
    .Y(_0385_),
    .A1(_0492_),
    .A2(_0163_));
 sg13g2_nand4_1 _0956_ (.B(_0379_),
    .C(_0384_),
    .A(_0377_),
    .Y(_0386_),
    .D(_0385_));
 sg13g2_nand2_1 _0957_ (.Y(_0388_),
    .A(_0494_),
    .B(_0386_));
 sg13g2_or2_1 _0958_ (.X(_0389_),
    .B(_0103_),
    .A(net265));
 sg13g2_nand2_1 _0959_ (.Y(_0390_),
    .A(net264),
    .B(_0103_));
 sg13g2_o21ai_1 _0960_ (.B1(_0389_),
    .Y(_0391_),
    .A1(_0105_),
    .A2(_0390_));
 sg13g2_and2_1 _0961_ (.A(net230),
    .B(_0391_),
    .X(_0392_));
 sg13g2_o21ai_1 _0962_ (.B1(_0390_),
    .Y(_0393_),
    .A1(net264),
    .A2(_0105_));
 sg13g2_or2_1 _0963_ (.X(_0394_),
    .B(_0391_),
    .A(_0504_));
 sg13g2_nor3_1 _0964_ (.A(net240),
    .B(net231),
    .C(_0393_),
    .Y(_0395_));
 sg13g2_a21oi_1 _0965_ (.A1(_0393_),
    .A2(_0394_),
    .Y(_0396_),
    .B1(_0395_));
 sg13g2_o21ai_1 _0966_ (.B1(_0204_),
    .Y(_0397_),
    .A1(_0392_),
    .A2(_0396_));
 sg13g2_nand3b_1 _0967_ (.B(_0388_),
    .C(_0397_),
    .Y(uio_out[0]),
    .A_N(_0373_));
 sg13g2_nand3_1 _0968_ (.B(net231),
    .C(_0132_),
    .A(net266),
    .Y(_0399_));
 sg13g2_a21oi_1 _0969_ (.A1(_0217_),
    .A2(_0222_),
    .Y(_0400_),
    .B1(_0220_));
 sg13g2_o21ai_1 _0970_ (.B1(_0494_),
    .Y(_0401_),
    .A1(_0227_),
    .A2(_0400_));
 sg13g2_nand3_1 _0971_ (.B(net244),
    .C(_0049_),
    .A(net266),
    .Y(_0402_));
 sg13g2_nand3_1 _0972_ (.B(_0303_),
    .C(_0402_),
    .A(_0504_),
    .Y(_0403_));
 sg13g2_and2_1 _0973_ (.A(_0226_),
    .B(_0403_),
    .X(_0404_));
 sg13g2_a22oi_1 _0974_ (.Y(uio_out[1]),
    .B1(_0401_),
    .B2(_0404_),
    .A2(_0399_),
    .A1(_0418_));
 sg13g2_a22oi_1 _0975_ (.Y(_0405_),
    .B1(_0030_),
    .B2(net269),
    .A2(_0019_),
    .A1(net237));
 sg13g2_nor2_1 _0976_ (.A(net263),
    .B(_0405_),
    .Y(_0406_));
 sg13g2_nor3_1 _0977_ (.A(net277),
    .B(_0489_),
    .C(_0013_),
    .Y(_0408_));
 sg13g2_a221oi_1 _0978_ (.B2(_0044_),
    .C1(_0406_),
    .B1(_0408_),
    .A1(_0032_),
    .Y(_0409_),
    .A2(_0056_));
 sg13g2_a22oi_1 _0979_ (.Y(_0410_),
    .B1(_0229_),
    .B2(net268),
    .A2(_0074_),
    .A1(_0473_));
 sg13g2_nor2_1 _0980_ (.A(_0498_),
    .B(_0410_),
    .Y(_0411_));
 sg13g2_nor2_1 _0981_ (.A(_0483_),
    .B(_0133_),
    .Y(_0412_));
 sg13g2_o21ai_1 _0982_ (.B1(_0412_),
    .Y(_0413_),
    .A1(net270),
    .A2(_0231_));
 sg13g2_o21ai_1 _0983_ (.B1(_0413_),
    .Y(_0414_),
    .A1(net260),
    .A2(_0409_));
 sg13g2_o21ai_1 _0984_ (.B1(_0215_),
    .Y(_0415_),
    .A1(_0411_),
    .A2(_0414_));
 sg13g2_nand3_1 _0985_ (.B(_0343_),
    .C(_0012_),
    .A(net280),
    .Y(_0416_));
 sg13g2_o21ai_1 _0986_ (.B1(_0204_),
    .Y(_0417_),
    .A1(_0503_),
    .A2(_0506_));
 sg13g2_nand2_1 _0987_ (.Y(_0419_),
    .A(net240),
    .B(_0060_));
 sg13g2_o21ai_1 _0988_ (.B1(net232),
    .Y(_0420_),
    .A1(_0138_),
    .A2(_0183_));
 sg13g2_a22oi_1 _0989_ (.Y(_0421_),
    .B1(_0044_),
    .B2(net233),
    .A2(net237),
    .A1(net242));
 sg13g2_a221oi_1 _0990_ (.B2(net230),
    .C1(_0417_),
    .B1(_0421_),
    .A1(_0058_),
    .Y(_0422_),
    .A2(_0416_));
 sg13g2_nand3_1 _0991_ (.B(_0420_),
    .C(_0422_),
    .A(_0419_),
    .Y(_0423_));
 sg13g2_nand2_2 _0992_ (.Y(uio_out[2]),
    .A(_0415_),
    .B(_0423_));
 sg13g2_and2_1 _0993_ (.A(_0172_),
    .B(_0088_),
    .X(_0424_));
 sg13g2_o21ai_1 _0994_ (.B1(_0344_),
    .Y(_0425_),
    .A1(net283),
    .A2(_0424_));
 sg13g2_nand2b_1 _0995_ (.Y(_0426_),
    .B(net252),
    .A_N(_0425_));
 sg13g2_nand2_1 _0996_ (.Y(_0427_),
    .A(net283),
    .B(_0424_));
 sg13g2_o21ai_1 _0997_ (.B1(_0427_),
    .Y(_0429_),
    .A1(net283),
    .A2(_0199_));
 sg13g2_nand2_1 _0998_ (.Y(_0430_),
    .A(net275),
    .B(_0429_));
 sg13g2_nand3_1 _0999_ (.B(_0426_),
    .C(_0430_),
    .A(_0099_),
    .Y(_0431_));
 sg13g2_nand2_1 _1000_ (.Y(_0432_),
    .A(_0172_),
    .B(_0091_));
 sg13g2_nor2_1 _1001_ (.A(_0483_),
    .B(_0140_),
    .Y(_0433_));
 sg13g2_a21oi_1 _1002_ (.A1(_0432_),
    .A2(_0433_),
    .Y(_0434_),
    .B1(net307));
 sg13g2_a22oi_1 _1003_ (.Y(_0435_),
    .B1(_0429_),
    .B2(net252),
    .A2(_0102_),
    .A1(_0172_));
 sg13g2_nand2_1 _1004_ (.Y(_0436_),
    .A(_0101_),
    .B(_0435_));
 sg13g2_nor3_1 _1005_ (.A(net275),
    .B(net303),
    .C(_0087_),
    .Y(_0437_));
 sg13g2_nor2b_1 _1006_ (.A(_0437_),
    .B_N(_0106_),
    .Y(_0438_));
 sg13g2_o21ai_1 _1007_ (.B1(_0438_),
    .Y(_0440_),
    .A1(net252),
    .A2(_0425_));
 sg13g2_nand4_1 _1008_ (.B(_0434_),
    .C(_0436_),
    .A(_0431_),
    .Y(_0441_),
    .D(_0440_));
 sg13g2_nor3_1 _1009_ (.A(_0082_),
    .B(_0084_),
    .C(_0272_),
    .Y(_0442_));
 sg13g2_a21oi_1 _1010_ (.A1(net294),
    .A2(net234),
    .Y(_0443_),
    .B1(net286));
 sg13g2_a21oi_1 _1011_ (.A1(net286),
    .A2(_0355_),
    .Y(_0444_),
    .B1(_0443_));
 sg13g2_mux2_1 _1012_ (.A0(_0442_),
    .A1(_0444_),
    .S(net279),
    .X(_0445_));
 sg13g2_nand2_1 _1013_ (.Y(_0446_),
    .A(net271),
    .B(_0445_));
 sg13g2_a22oi_1 _1014_ (.Y(_0447_),
    .B1(_0342_),
    .B2(net284),
    .A2(_0199_),
    .A1(_0000_));
 sg13g2_o21ai_1 _1015_ (.B1(_0341_),
    .Y(_0448_),
    .A1(net286),
    .A2(_0355_));
 sg13g2_a22oi_1 _1016_ (.Y(_0449_),
    .B1(_0448_),
    .B2(_0016_),
    .A2(_0447_),
    .A1(net236));
 sg13g2_nand2_1 _1017_ (.Y(_0451_),
    .A(_0446_),
    .B(_0449_));
 sg13g2_a22oi_1 _1018_ (.Y(_0452_),
    .B1(_0082_),
    .B2(_0273_),
    .A2(_0333_),
    .A1(_0258_));
 sg13g2_nor2_1 _1019_ (.A(net279),
    .B(_0452_),
    .Y(_0453_));
 sg13g2_a21oi_1 _1020_ (.A1(net279),
    .A2(_0447_),
    .Y(_0454_),
    .B1(_0453_));
 sg13g2_nand2_1 _1021_ (.Y(_0455_),
    .A(_0014_),
    .B(_0019_));
 sg13g2_a22oi_1 _1022_ (.Y(_0456_),
    .B1(_0455_),
    .B2(_0490_),
    .A2(_0448_),
    .A1(net233));
 sg13g2_o21ai_1 _1023_ (.B1(_0456_),
    .Y(_0457_),
    .A1(net273),
    .A2(_0454_));
 sg13g2_a21oi_1 _1024_ (.A1(net273),
    .A2(_0454_),
    .Y(_0458_),
    .B1(_0407_));
 sg13g2_o21ai_1 _1025_ (.B1(_0458_),
    .Y(_0459_),
    .A1(net273),
    .A2(_0445_));
 sg13g2_nand2_1 _1026_ (.Y(_0460_),
    .A(_0016_),
    .B(_0442_));
 sg13g2_o21ai_1 _1027_ (.B1(_0460_),
    .Y(_0462_),
    .A1(_0491_),
    .A2(_0452_));
 sg13g2_a221oi_1 _1028_ (.B2(_0477_),
    .C1(_0462_),
    .B1(_0448_),
    .A1(_0467_),
    .Y(_0463_),
    .A2(_0444_));
 sg13g2_o21ai_1 _1029_ (.B1(_0459_),
    .Y(_0464_),
    .A1(_0504_),
    .A2(_0463_));
 sg13g2_a221oi_1 _1030_ (.B2(net232),
    .C1(_0464_),
    .B1(_0457_),
    .A1(net230),
    .Y(_0465_),
    .A2(_0451_));
 sg13g2_o21ai_1 _1031_ (.B1(_0441_),
    .Y(uio_out[3]),
    .A1(_0226_),
    .A2(_0465_));
 sg13g2_tiehi tt_um_rejunity_decoder_9 (.L_HI(net9));
 sg13g2_tiehi tt_um_rejunity_decoder_10 (.L_HI(net10));
 sg13g2_tiehi tt_um_rejunity_decoder_11 (.L_HI(net11));
 sg13g2_tiehi tt_um_rejunity_decoder_12 (.L_HI(net12));
 sg13g2_tiehi tt_um_rejunity_decoder_13 (.L_HI(net13));
 sg13g2_tiehi tt_um_rejunity_decoder_14 (.L_HI(net14));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_tielo tt_um_rejunity_decoder_4 (.L_LO(net4));
 sg13g2_tielo tt_um_rejunity_decoder_5 (.L_LO(net5));
 sg13g2_tielo tt_um_rejunity_decoder_6 (.L_LO(net6));
 sg13g2_tielo tt_um_rejunity_decoder_7 (.L_LO(net7));
 sg13g2_tiehi tt_um_rejunity_decoder_8 (.L_HI(net8));
 sg13g2_buf_4 fanout230 (.X(net230),
    .A(_0497_));
 sg13g2_buf_4 fanout231 (.X(net231),
    .A(_0482_));
 sg13g2_buf_4 fanout232 (.X(net232),
    .A(_0482_));
 sg13g2_buf_4 fanout233 (.X(net233),
    .A(_0467_));
 sg13g2_buf_4 fanout234 (.X(net234),
    .A(_0006_));
 sg13g2_buf_4 fanout235 (.X(net235),
    .A(_0500_));
 sg13g2_buf_2 fanout236 (.A(_0477_),
    .X(net236));
 sg13g2_buf_4 fanout237 (.X(net237),
    .A(_0477_));
 sg13g2_buf_4 fanout238 (.X(net238),
    .A(_0475_));
 sg13g2_buf_4 fanout239 (.X(net239),
    .A(_0470_));
 sg13g2_buf_4 fanout240 (.X(net240),
    .A(_0398_));
 sg13g2_buf_4 fanout241 (.X(net241),
    .A(_0343_));
 sg13g2_buf_4 fanout242 (.X(net242),
    .A(_0333_));
 sg13g2_buf_4 fanout243 (.X(net243),
    .A(_0193_));
 sg13g2_buf_2 fanout244 (.A(_0193_),
    .X(net244));
 sg13g2_buf_4 fanout245 (.X(net245),
    .A(net248));
 sg13g2_buf_2 fanout246 (.A(net248),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(net248),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_0182_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(net251),
    .X(net249));
 sg13g2_buf_4 fanout250 (.X(net250),
    .A(net251));
 sg13g2_buf_2 fanout251 (.A(_0150_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(net253),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(net254),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(net256),
    .X(net254));
 sg13g2_buf_4 fanout255 (.X(net255),
    .A(net256));
 sg13g2_buf_2 fanout256 (.A(_0139_),
    .X(net256));
 sg13g2_buf_4 fanout257 (.X(net257),
    .A(_0129_));
 sg13g2_buf_4 fanout258 (.X(net258),
    .A(net260));
 sg13g2_buf_2 fanout259 (.A(net260),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(ui_in[7]),
    .X(net260));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(net262));
 sg13g2_buf_4 fanout262 (.X(net262),
    .A(net263));
 sg13g2_buf_2 fanout263 (.A(ui_in[6]),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(net265),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(net266),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(net274),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(net268),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(net274),
    .X(net268));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(net274));
 sg13g2_buf_1 fanout270 (.A(net274),
    .X(net270));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(net273));
 sg13g2_buf_2 fanout272 (.A(net273),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(net274),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(ui_in[5]),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(net277),
    .X(net275));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(net277));
 sg13g2_buf_2 fanout277 (.A(ui_in[4]),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(net282),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(net282),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(net282),
    .X(net280));
 sg13g2_buf_1 fanout281 (.A(net282),
    .X(net281));
 sg13g2_buf_1 fanout282 (.A(ui_in[4]),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(net284),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(net285),
    .X(net284));
 sg13g2_buf_1 fanout285 (.A(ui_in[3]),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(net288),
    .X(net286));
 sg13g2_buf_1 fanout287 (.A(net288),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(net289),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(ui_in[3]),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(net291),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(net292),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(net296),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(net295),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(net295),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(net296),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(ui_in[2]),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(net301),
    .X(net297));
 sg13g2_buf_1 fanout298 (.A(net301),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(net300),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(net301),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(ui_in[1]),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(net303),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(net304),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(net1),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(net306),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(net1),
    .X(net306));
 sg13g2_buf_4 fanout307 (.X(net307),
    .A(net308));
 sg13g2_buf_2 fanout308 (.A(ena),
    .X(net308));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(uio_in[7]),
    .X(net2));
 sg13g2_tielo tt_um_rejunity_decoder_3 (.L_LO(net3));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_fill_2 FILLER_19_231 ();
 sg13g2_fill_1 FILLER_19_233 ();
 sg13g2_decap_8 FILLER_19_240 ();
 sg13g2_decap_8 FILLER_19_247 ();
 sg13g2_decap_8 FILLER_19_254 ();
 sg13g2_fill_2 FILLER_19_261 ();
 sg13g2_decap_8 FILLER_19_268 ();
 sg13g2_decap_8 FILLER_19_275 ();
 sg13g2_decap_8 FILLER_19_292 ();
 sg13g2_decap_8 FILLER_19_299 ();
 sg13g2_decap_8 FILLER_19_306 ();
 sg13g2_decap_8 FILLER_19_313 ();
 sg13g2_decap_8 FILLER_19_320 ();
 sg13g2_decap_8 FILLER_19_327 ();
 sg13g2_fill_2 FILLER_19_334 ();
 sg13g2_decap_8 FILLER_19_346 ();
 sg13g2_fill_2 FILLER_19_353 ();
 sg13g2_fill_1 FILLER_19_355 ();
 sg13g2_decap_8 FILLER_19_361 ();
 sg13g2_decap_8 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_4 FILLER_20_210 ();
 sg13g2_fill_2 FILLER_20_214 ();
 sg13g2_decap_4 FILLER_20_223 ();
 sg13g2_fill_1 FILLER_20_227 ();
 sg13g2_decap_4 FILLER_20_249 ();
 sg13g2_fill_1 FILLER_20_253 ();
 sg13g2_decap_4 FILLER_20_275 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_313 ();
 sg13g2_decap_8 FILLER_20_320 ();
 sg13g2_fill_2 FILLER_20_327 ();
 sg13g2_fill_1 FILLER_20_329 ();
 sg13g2_fill_2 FILLER_20_350 ();
 sg13g2_fill_1 FILLER_20_352 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_fill_1 FILLER_21_189 ();
 sg13g2_decap_4 FILLER_21_194 ();
 sg13g2_decap_4 FILLER_21_203 ();
 sg13g2_fill_2 FILLER_21_207 ();
 sg13g2_decap_4 FILLER_21_232 ();
 sg13g2_decap_4 FILLER_21_260 ();
 sg13g2_fill_1 FILLER_21_264 ();
 sg13g2_fill_2 FILLER_21_269 ();
 sg13g2_fill_1 FILLER_21_271 ();
 sg13g2_decap_4 FILLER_21_285 ();
 sg13g2_decap_4 FILLER_21_293 ();
 sg13g2_fill_1 FILLER_21_302 ();
 sg13g2_fill_2 FILLER_21_313 ();
 sg13g2_fill_2 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_decap_4 FILLER_21_359 ();
 sg13g2_decap_8 FILLER_21_384 ();
 sg13g2_decap_8 FILLER_21_391 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_fill_2 FILLER_22_185 ();
 sg13g2_fill_2 FILLER_22_191 ();
 sg13g2_decap_8 FILLER_22_223 ();
 sg13g2_fill_2 FILLER_22_230 ();
 sg13g2_decap_4 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_277 ();
 sg13g2_decap_4 FILLER_22_284 ();
 sg13g2_decap_4 FILLER_22_294 ();
 sg13g2_fill_2 FILLER_22_298 ();
 sg13g2_fill_1 FILLER_22_308 ();
 sg13g2_fill_2 FILLER_22_312 ();
 sg13g2_fill_1 FILLER_22_314 ();
 sg13g2_fill_2 FILLER_22_347 ();
 sg13g2_fill_1 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_fill_1 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_4 FILLER_23_159 ();
 sg13g2_fill_1 FILLER_23_163 ();
 sg13g2_fill_1 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_206 ();
 sg13g2_fill_2 FILLER_23_227 ();
 sg13g2_fill_1 FILLER_23_229 ();
 sg13g2_fill_2 FILLER_23_241 ();
 sg13g2_decap_4 FILLER_23_249 ();
 sg13g2_fill_1 FILLER_23_253 ();
 sg13g2_decap_4 FILLER_23_269 ();
 sg13g2_decap_4 FILLER_23_295 ();
 sg13g2_fill_1 FILLER_23_310 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_fill_2 FILLER_23_336 ();
 sg13g2_fill_1 FILLER_23_342 ();
 sg13g2_fill_2 FILLER_23_354 ();
 sg13g2_fill_1 FILLER_23_356 ();
 sg13g2_fill_1 FILLER_23_371 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_166 ();
 sg13g2_fill_1 FILLER_24_173 ();
 sg13g2_fill_1 FILLER_24_192 ();
 sg13g2_decap_8 FILLER_24_213 ();
 sg13g2_fill_1 FILLER_24_220 ();
 sg13g2_decap_4 FILLER_24_227 ();
 sg13g2_fill_1 FILLER_24_231 ();
 sg13g2_decap_4 FILLER_24_254 ();
 sg13g2_decap_8 FILLER_24_275 ();
 sg13g2_decap_8 FILLER_24_282 ();
 sg13g2_decap_4 FILLER_24_289 ();
 sg13g2_fill_1 FILLER_24_293 ();
 sg13g2_decap_8 FILLER_24_330 ();
 sg13g2_fill_2 FILLER_24_337 ();
 sg13g2_fill_1 FILLER_24_339 ();
 sg13g2_fill_1 FILLER_24_371 ();
 sg13g2_fill_2 FILLER_24_382 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_4 FILLER_25_147 ();
 sg13g2_fill_2 FILLER_25_174 ();
 sg13g2_fill_1 FILLER_25_176 ();
 sg13g2_fill_2 FILLER_25_198 ();
 sg13g2_fill_1 FILLER_25_200 ();
 sg13g2_decap_8 FILLER_25_212 ();
 sg13g2_fill_1 FILLER_25_219 ();
 sg13g2_fill_2 FILLER_25_232 ();
 sg13g2_fill_2 FILLER_25_239 ();
 sg13g2_fill_1 FILLER_25_241 ();
 sg13g2_fill_1 FILLER_25_255 ();
 sg13g2_fill_1 FILLER_25_278 ();
 sg13g2_decap_8 FILLER_25_293 ();
 sg13g2_decap_8 FILLER_25_300 ();
 sg13g2_fill_2 FILLER_25_317 ();
 sg13g2_fill_1 FILLER_25_319 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_fill_2 FILLER_25_347 ();
 sg13g2_fill_2 FILLER_25_366 ();
 sg13g2_fill_1 FILLER_25_368 ();
 sg13g2_fill_1 FILLER_25_383 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_4 FILLER_26_147 ();
 sg13g2_fill_1 FILLER_26_151 ();
 sg13g2_decap_4 FILLER_26_178 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_fill_1 FILLER_26_200 ();
 sg13g2_fill_2 FILLER_26_205 ();
 sg13g2_fill_2 FILLER_26_218 ();
 sg13g2_fill_1 FILLER_26_220 ();
 sg13g2_fill_1 FILLER_26_231 ();
 sg13g2_fill_1 FILLER_26_237 ();
 sg13g2_decap_8 FILLER_26_251 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_fill_2 FILLER_26_263 ();
 sg13g2_decap_4 FILLER_26_277 ();
 sg13g2_fill_2 FILLER_26_281 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_fill_1 FILLER_26_303 ();
 sg13g2_fill_1 FILLER_26_323 ();
 sg13g2_fill_2 FILLER_26_330 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_363 ();
 sg13g2_decap_8 FILLER_26_370 ();
 sg13g2_fill_2 FILLER_26_377 ();
 sg13g2_fill_1 FILLER_26_379 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_4 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_fill_2 FILLER_27_176 ();
 sg13g2_fill_1 FILLER_27_178 ();
 sg13g2_fill_1 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_fill_2 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_233 ();
 sg13g2_decap_8 FILLER_27_239 ();
 sg13g2_decap_4 FILLER_27_251 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_fill_1 FILLER_27_296 ();
 sg13g2_fill_1 FILLER_27_306 ();
 sg13g2_fill_2 FILLER_27_330 ();
 sg13g2_decap_4 FILLER_27_342 ();
 sg13g2_fill_1 FILLER_27_346 ();
 sg13g2_fill_2 FILLER_27_368 ();
 sg13g2_fill_1 FILLER_27_374 ();
 sg13g2_decap_4 FILLER_27_380 ();
 sg13g2_fill_2 FILLER_27_389 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_4 FILLER_28_140 ();
 sg13g2_fill_1 FILLER_28_162 ();
 sg13g2_fill_2 FILLER_28_168 ();
 sg13g2_decap_4 FILLER_28_180 ();
 sg13g2_fill_1 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_197 ();
 sg13g2_fill_1 FILLER_28_204 ();
 sg13g2_fill_1 FILLER_28_209 ();
 sg13g2_fill_2 FILLER_28_214 ();
 sg13g2_fill_1 FILLER_28_226 ();
 sg13g2_decap_4 FILLER_28_233 ();
 sg13g2_decap_4 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_276 ();
 sg13g2_fill_2 FILLER_28_303 ();
 sg13g2_fill_1 FILLER_28_305 ();
 sg13g2_decap_4 FILLER_28_312 ();
 sg13g2_fill_2 FILLER_28_316 ();
 sg13g2_decap_8 FILLER_28_344 ();
 sg13g2_fill_1 FILLER_28_355 ();
 sg13g2_fill_2 FILLER_28_362 ();
 sg13g2_fill_1 FILLER_28_364 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_fill_2 FILLER_29_147 ();
 sg13g2_fill_1 FILLER_29_149 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_fill_2 FILLER_29_175 ();
 sg13g2_decap_4 FILLER_29_195 ();
 sg13g2_fill_2 FILLER_29_208 ();
 sg13g2_fill_2 FILLER_29_225 ();
 sg13g2_fill_1 FILLER_29_227 ();
 sg13g2_decap_8 FILLER_29_235 ();
 sg13g2_fill_2 FILLER_29_242 ();
 sg13g2_decap_4 FILLER_29_254 ();
 sg13g2_fill_1 FILLER_29_258 ();
 sg13g2_decap_8 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_271 ();
 sg13g2_fill_2 FILLER_29_284 ();
 sg13g2_fill_2 FILLER_29_296 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_4 FILLER_29_328 ();
 sg13g2_fill_1 FILLER_29_332 ();
 sg13g2_fill_2 FILLER_29_358 ();
 sg13g2_fill_1 FILLER_29_360 ();
 sg13g2_decap_4 FILLER_29_370 ();
 sg13g2_fill_1 FILLER_29_374 ();
 sg13g2_decap_4 FILLER_29_384 ();
 sg13g2_fill_1 FILLER_29_393 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_4 FILLER_30_154 ();
 sg13g2_fill_2 FILLER_30_158 ();
 sg13g2_fill_2 FILLER_30_167 ();
 sg13g2_decap_8 FILLER_30_174 ();
 sg13g2_fill_2 FILLER_30_200 ();
 sg13g2_fill_1 FILLER_30_202 ();
 sg13g2_decap_8 FILLER_30_225 ();
 sg13g2_fill_1 FILLER_30_232 ();
 sg13g2_decap_4 FILLER_30_237 ();
 sg13g2_decap_8 FILLER_30_279 ();
 sg13g2_fill_1 FILLER_30_286 ();
 sg13g2_decap_8 FILLER_30_305 ();
 sg13g2_fill_1 FILLER_30_312 ();
 sg13g2_fill_1 FILLER_30_323 ();
 sg13g2_fill_1 FILLER_30_329 ();
 sg13g2_fill_2 FILLER_30_340 ();
 sg13g2_fill_2 FILLER_30_357 ();
 sg13g2_fill_1 FILLER_30_359 ();
 sg13g2_fill_2 FILLER_30_371 ();
 sg13g2_fill_1 FILLER_30_373 ();
 sg13g2_fill_2 FILLER_30_380 ();
 sg13g2_fill_1 FILLER_30_382 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_4 FILLER_31_176 ();
 sg13g2_fill_1 FILLER_31_180 ();
 sg13g2_decap_4 FILLER_31_195 ();
 sg13g2_fill_1 FILLER_31_199 ();
 sg13g2_decap_8 FILLER_31_209 ();
 sg13g2_decap_4 FILLER_31_239 ();
 sg13g2_fill_1 FILLER_31_248 ();
 sg13g2_fill_1 FILLER_31_260 ();
 sg13g2_decap_4 FILLER_31_266 ();
 sg13g2_fill_2 FILLER_31_306 ();
 sg13g2_fill_1 FILLER_31_308 ();
 sg13g2_fill_1 FILLER_31_327 ();
 sg13g2_fill_2 FILLER_31_343 ();
 sg13g2_fill_1 FILLER_31_356 ();
 sg13g2_fill_1 FILLER_31_361 ();
 sg13g2_fill_2 FILLER_31_377 ();
 sg13g2_decap_4 FILLER_31_383 ();
 sg13g2_fill_1 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_fill_1 FILLER_32_165 ();
 sg13g2_fill_2 FILLER_32_180 ();
 sg13g2_fill_2 FILLER_32_186 ();
 sg13g2_fill_1 FILLER_32_188 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_fill_2 FILLER_32_217 ();
 sg13g2_fill_1 FILLER_32_219 ();
 sg13g2_decap_8 FILLER_32_236 ();
 sg13g2_fill_2 FILLER_32_257 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_decap_4 FILLER_32_287 ();
 sg13g2_fill_2 FILLER_32_300 ();
 sg13g2_fill_1 FILLER_32_307 ();
 sg13g2_decap_8 FILLER_32_313 ();
 sg13g2_fill_2 FILLER_32_320 ();
 sg13g2_fill_1 FILLER_32_322 ();
 sg13g2_decap_4 FILLER_32_328 ();
 sg13g2_fill_1 FILLER_32_332 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_decap_8 FILLER_32_346 ();
 sg13g2_fill_2 FILLER_32_359 ();
 sg13g2_fill_2 FILLER_32_366 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_fill_2 FILLER_33_168 ();
 sg13g2_fill_1 FILLER_33_181 ();
 sg13g2_fill_2 FILLER_33_200 ();
 sg13g2_decap_8 FILLER_33_213 ();
 sg13g2_fill_2 FILLER_33_220 ();
 sg13g2_fill_2 FILLER_33_237 ();
 sg13g2_decap_4 FILLER_33_248 ();
 sg13g2_fill_1 FILLER_33_252 ();
 sg13g2_decap_4 FILLER_33_259 ();
 sg13g2_fill_1 FILLER_33_285 ();
 sg13g2_fill_1 FILLER_33_290 ();
 sg13g2_decap_4 FILLER_33_328 ();
 sg13g2_fill_1 FILLER_33_342 ();
 sg13g2_decap_4 FILLER_33_357 ();
 sg13g2_fill_1 FILLER_33_361 ();
 sg13g2_decap_8 FILLER_33_369 ();
 sg13g2_decap_4 FILLER_33_385 ();
 sg13g2_fill_1 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_395 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_4 FILLER_34_161 ();
 sg13g2_fill_1 FILLER_34_165 ();
 sg13g2_decap_4 FILLER_34_177 ();
 sg13g2_fill_1 FILLER_34_181 ();
 sg13g2_fill_2 FILLER_34_188 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_fill_1 FILLER_34_203 ();
 sg13g2_fill_2 FILLER_34_241 ();
 sg13g2_decap_4 FILLER_34_257 ();
 sg13g2_fill_2 FILLER_34_261 ();
 sg13g2_fill_1 FILLER_34_268 ();
 sg13g2_decap_4 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_289 ();
 sg13g2_fill_1 FILLER_34_291 ();
 sg13g2_fill_1 FILLER_34_304 ();
 sg13g2_fill_2 FILLER_34_311 ();
 sg13g2_fill_1 FILLER_34_313 ();
 sg13g2_decap_4 FILLER_34_318 ();
 sg13g2_fill_2 FILLER_34_322 ();
 sg13g2_fill_1 FILLER_34_351 ();
 sg13g2_decap_4 FILLER_34_360 ();
 sg13g2_decap_4 FILLER_34_368 ();
 sg13g2_fill_2 FILLER_34_372 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_fill_2 FILLER_35_168 ();
 sg13g2_fill_2 FILLER_35_178 ();
 sg13g2_fill_2 FILLER_35_188 ();
 sg13g2_fill_1 FILLER_35_190 ();
 sg13g2_decap_8 FILLER_35_205 ();
 sg13g2_fill_2 FILLER_35_220 ();
 sg13g2_fill_2 FILLER_35_232 ();
 sg13g2_decap_8 FILLER_35_265 ();
 sg13g2_decap_8 FILLER_35_283 ();
 sg13g2_fill_2 FILLER_35_290 ();
 sg13g2_fill_1 FILLER_35_318 ();
 sg13g2_fill_2 FILLER_35_324 ();
 sg13g2_fill_1 FILLER_35_339 ();
 sg13g2_fill_2 FILLER_35_361 ();
 sg13g2_fill_1 FILLER_35_363 ();
 sg13g2_fill_1 FILLER_35_375 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_4 FILLER_36_175 ();
 sg13g2_fill_1 FILLER_36_179 ();
 sg13g2_fill_1 FILLER_36_184 ();
 sg13g2_fill_1 FILLER_36_191 ();
 sg13g2_fill_2 FILLER_36_206 ();
 sg13g2_fill_1 FILLER_36_208 ();
 sg13g2_fill_1 FILLER_36_214 ();
 sg13g2_fill_2 FILLER_36_220 ();
 sg13g2_fill_1 FILLER_36_238 ();
 sg13g2_fill_2 FILLER_36_255 ();
 sg13g2_fill_1 FILLER_36_261 ();
 sg13g2_fill_2 FILLER_36_267 ();
 sg13g2_decap_4 FILLER_36_279 ();
 sg13g2_fill_1 FILLER_36_283 ();
 sg13g2_decap_8 FILLER_36_305 ();
 sg13g2_decap_4 FILLER_36_312 ();
 sg13g2_fill_2 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_333 ();
 sg13g2_fill_1 FILLER_36_335 ();
 sg13g2_fill_1 FILLER_36_346 ();
 sg13g2_decap_8 FILLER_36_366 ();
 sg13g2_fill_1 FILLER_36_373 ();
 sg13g2_decap_4 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_decap_8 FILLER_36_395 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_fill_1 FILLER_37_217 ();
 sg13g2_fill_1 FILLER_37_240 ();
 sg13g2_fill_2 FILLER_37_250 ();
 sg13g2_fill_1 FILLER_37_252 ();
 sg13g2_fill_1 FILLER_37_271 ();
 sg13g2_decap_8 FILLER_37_276 ();
 sg13g2_fill_2 FILLER_37_283 ();
 sg13g2_decap_8 FILLER_37_312 ();
 sg13g2_fill_1 FILLER_37_319 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_fill_1 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_380 ();
 sg13g2_decap_8 FILLER_37_387 ();
 sg13g2_decap_8 FILLER_37_394 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_148 ();
 sg13g2_decap_8 FILLER_38_155 ();
 sg13g2_decap_8 FILLER_38_162 ();
 sg13g2_decap_8 FILLER_38_169 ();
 sg13g2_decap_8 FILLER_38_176 ();
 sg13g2_decap_8 FILLER_38_183 ();
 sg13g2_decap_8 FILLER_38_190 ();
 sg13g2_decap_8 FILLER_38_197 ();
 sg13g2_decap_8 FILLER_38_204 ();
 sg13g2_decap_8 FILLER_38_211 ();
 sg13g2_decap_8 FILLER_38_218 ();
 sg13g2_decap_8 FILLER_38_225 ();
 sg13g2_fill_2 FILLER_38_232 ();
 sg13g2_fill_1 FILLER_38_234 ();
 sg13g2_decap_4 FILLER_38_243 ();
 sg13g2_decap_4 FILLER_38_262 ();
 sg13g2_decap_8 FILLER_38_274 ();
 sg13g2_decap_4 FILLER_38_291 ();
 sg13g2_decap_8 FILLER_38_304 ();
 sg13g2_decap_8 FILLER_38_311 ();
 sg13g2_decap_8 FILLER_38_318 ();
 sg13g2_decap_8 FILLER_38_331 ();
 sg13g2_decap_8 FILLER_38_338 ();
 sg13g2_decap_8 FILLER_38_345 ();
 sg13g2_decap_8 FILLER_38_352 ();
 sg13g2_decap_8 FILLER_38_359 ();
 sg13g2_fill_2 FILLER_38_366 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net8;
 assign uio_oe[1] = net9;
 assign uio_oe[2] = net10;
 assign uio_oe[3] = net11;
 assign uio_oe[4] = net12;
 assign uio_oe[5] = net13;
 assign uio_oe[6] = net14;
 assign uio_oe[7] = net3;
 assign uio_out[4] = net4;
 assign uio_out[5] = net5;
 assign uio_out[6] = net6;
 assign uio_out[7] = net7;
endmodule

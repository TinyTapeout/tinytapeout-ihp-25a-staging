module tt_um_wokwi_group_1 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire \proj_10.net4 ;
 wire \proj_10.net5 ;
 wire \proj_10.net7 ;
 wire \proj_10.net8 ;
 wire \proj_10.net9 ;
 wire \proj_11.net10 ;
 wire \proj_11.net16 ;
 wire \proj_11.net18 ;
 wire \proj_11.net19 ;
 wire \proj_11.net20 ;
 wire \proj_11.net21 ;
 wire \proj_11.net22 ;
 wire \proj_11.net23 ;
 wire \proj_11.net24 ;
 wire \proj_11.net25 ;
 wire \proj_11.net3 ;
 wire \proj_11.net4 ;
 wire \proj_11.net5 ;
 wire \proj_11.net6 ;
 wire \proj_11.net7 ;
 wire \proj_11.net8 ;
 wire \proj_11.net9 ;
 wire \proj_12.net10 ;
 wire \proj_12.net11 ;
 wire \proj_12.net12 ;
 wire \proj_12.net13 ;
 wire \proj_12.net14 ;
 wire \proj_12.net15 ;
 wire \proj_12.net16 ;
 wire \proj_12.net22 ;
 wire \proj_12.net23 ;
 wire \proj_12.net24 ;
 wire \proj_12.net25 ;
 wire \proj_12.net26 ;
 wire \proj_12.net27 ;
 wire \proj_12.net28 ;
 wire \proj_12.net29 ;
 wire \proj_12.net30 ;
 wire \proj_12.net31 ;
 wire \proj_12.net32 ;
 wire \proj_12.net33 ;
 wire \proj_12.net34 ;
 wire \proj_12.net35 ;
 wire \proj_12.net36 ;
 wire \proj_12.net37 ;
 wire \proj_12.net38 ;
 wire \proj_12.net39 ;
 wire \proj_12.net40 ;
 wire \proj_12.net41 ;
 wire \proj_12.net42 ;
 wire \proj_12.net43 ;
 wire \proj_12.net44 ;
 wire \proj_12.net45 ;
 wire \proj_12.net46 ;
 wire \proj_12.net47 ;
 wire \proj_12.net48 ;
 wire \proj_12.net49 ;
 wire \proj_12.net50 ;
 wire \proj_12.net9 ;
 wire \proj_14.net15 ;
 wire \proj_14.net16 ;
 wire \proj_14.net17 ;
 wire \proj_14.net18 ;
 wire \proj_14.net19 ;
 wire \proj_14.net20 ;
 wire \proj_14.net9 ;
 wire \proj__0.net10 ;
 wire \proj__0.net11 ;
 wire \proj__0.net9 ;
 wire \proj__1.net13 ;
 wire \proj__1.net14 ;
 wire \proj__1.net7 ;
 wire \proj__2.net11 ;
 wire \proj__2.net12 ;
 wire \proj__2.net13 ;
 wire \proj__2.net4 ;
 wire \proj__2.net5 ;
 wire \proj__3.net10 ;
 wire \proj__3.net11 ;
 wire \proj__3.net12 ;
 wire \proj__3.net13 ;
 wire \proj__3.net14 ;
 wire \proj__3.net9 ;
 wire \proj__4.net10 ;
 wire clk_regs;
 wire \proj__4.net12 ;
 wire \proj__4.net13 ;
 wire \proj__5.net10 ;
 wire \proj__5.net9 ;
 wire \proj__6.net10 ;
 wire \proj__6.net11 ;
 wire \proj__6.net12 ;
 wire \proj__6.net17 ;
 wire \proj__6.net18 ;
 wire \proj__6.net19 ;
 wire \proj__6.net20 ;
 wire \proj__6.net21 ;
 wire \proj__6.net22 ;
 wire \proj__6.net23 ;
 wire \proj__6.net24 ;
 wire \proj__6.net25 ;
 wire \proj__7.net10 ;
 wire \proj__7.net8 ;
 wire \proj__7.net9 ;
 wire \proj__8.net10 ;
 wire \proj__8.net100 ;
 wire \proj__8.net101 ;
 wire \proj__8.net102 ;
 wire \proj__8.net103 ;
 wire \proj__8.net104 ;
 wire \proj__8.net105 ;
 wire \proj__8.net106 ;
 wire \proj__8.net107 ;
 wire \proj__8.net108 ;
 wire \proj__8.net109 ;
 wire \proj__8.net11 ;
 wire \proj__8.net110 ;
 wire \proj__8.net111 ;
 wire \proj__8.net112 ;
 wire \proj__8.net113 ;
 wire \proj__8.net114 ;
 wire \proj__8.net115 ;
 wire \proj__8.net116 ;
 wire \proj__8.net117 ;
 wire \proj__8.net118 ;
 wire \proj__8.net119 ;
 wire \proj__8.net120 ;
 wire \proj__8.net121 ;
 wire \proj__8.net122 ;
 wire \proj__8.net123 ;
 wire \proj__8.net124 ;
 wire \proj__8.net125 ;
 wire \proj__8.net126 ;
 wire \proj__8.net127 ;
 wire \proj__8.net128 ;
 wire \proj__8.net129 ;
 wire \proj__8.net130 ;
 wire \proj__8.net131 ;
 wire \proj__8.net132 ;
 wire \proj__8.net133 ;
 wire \proj__8.net134 ;
 wire \proj__8.net135 ;
 wire \proj__8.net136 ;
 wire \proj__8.net137 ;
 wire \proj__8.net138 ;
 wire \proj__8.net139 ;
 wire \proj__8.net140 ;
 wire \proj__8.net141 ;
 wire \proj__8.net142 ;
 wire \proj__8.net143 ;
 wire \proj__8.net144 ;
 wire \proj__8.net145 ;
 wire \proj__8.net146 ;
 wire \proj__8.net147 ;
 wire \proj__8.net148 ;
 wire \proj__8.net149 ;
 wire \proj__8.net150 ;
 wire \proj__8.net151 ;
 wire \proj__8.net152 ;
 wire \proj__8.net153 ;
 wire \proj__8.net154 ;
 wire \proj__8.net155 ;
 wire \proj__8.net156 ;
 wire \proj__8.net157 ;
 wire \proj__8.net158 ;
 wire \proj__8.net159 ;
 wire \proj__8.net160 ;
 wire \proj__8.net161 ;
 wire \proj__8.net162 ;
 wire \proj__8.net163 ;
 wire \proj__8.net164 ;
 wire \proj__8.net165 ;
 wire \proj__8.net166 ;
 wire \proj__8.net167 ;
 wire \proj__8.net168 ;
 wire \proj__8.net169 ;
 wire \proj__8.net17 ;
 wire \proj__8.net170 ;
 wire \proj__8.net171 ;
 wire \proj__8.net172 ;
 wire \proj__8.net173 ;
 wire \proj__8.net174 ;
 wire \proj__8.net175 ;
 wire \proj__8.net176 ;
 wire \proj__8.net177 ;
 wire \proj__8.net178 ;
 wire \proj__8.net179 ;
 wire \proj__8.net18 ;
 wire \proj__8.net180 ;
 wire \proj__8.net181 ;
 wire \proj__8.net182 ;
 wire \proj__8.net183 ;
 wire \proj__8.net184 ;
 wire \proj__8.net185 ;
 wire \proj__8.net186 ;
 wire \proj__8.net187 ;
 wire \proj__8.net188 ;
 wire \proj__8.net189 ;
 wire \proj__8.net19 ;
 wire \proj__8.net190 ;
 wire \proj__8.net191 ;
 wire \proj__8.net192 ;
 wire \proj__8.net193 ;
 wire \proj__8.net194 ;
 wire \proj__8.net195 ;
 wire \proj__8.net196 ;
 wire \proj__8.net197 ;
 wire \proj__8.net198 ;
 wire \proj__8.net199 ;
 wire \proj__8.net20 ;
 wire \proj__8.net200 ;
 wire \proj__8.net201 ;
 wire \proj__8.net202 ;
 wire \proj__8.net203 ;
 wire \proj__8.net204 ;
 wire \proj__8.net205 ;
 wire \proj__8.net206 ;
 wire \proj__8.net207 ;
 wire \proj__8.net208 ;
 wire \proj__8.net209 ;
 wire \proj__8.net21 ;
 wire \proj__8.net210 ;
 wire \proj__8.net211 ;
 wire \proj__8.net212 ;
 wire \proj__8.net213 ;
 wire \proj__8.net214 ;
 wire \proj__8.net215 ;
 wire \proj__8.net216 ;
 wire \proj__8.net217 ;
 wire \proj__8.net218 ;
 wire \proj__8.net219 ;
 wire \proj__8.net22 ;
 wire \proj__8.net220 ;
 wire \proj__8.net221 ;
 wire \proj__8.net222 ;
 wire \proj__8.net223 ;
 wire \proj__8.net224 ;
 wire \proj__8.net225 ;
 wire \proj__8.net226 ;
 wire \proj__8.net227 ;
 wire \proj__8.net228 ;
 wire \proj__8.net229 ;
 wire \proj__8.net23 ;
 wire \proj__8.net230 ;
 wire \proj__8.net231 ;
 wire \proj__8.net232 ;
 wire \proj__8.net233 ;
 wire \proj__8.net234 ;
 wire \proj__8.net235 ;
 wire \proj__8.net236 ;
 wire \proj__8.net237 ;
 wire \proj__8.net238 ;
 wire \proj__8.net239 ;
 wire \proj__8.net24 ;
 wire \proj__8.net240 ;
 wire \proj__8.net241 ;
 wire \proj__8.net242 ;
 wire \proj__8.net243 ;
 wire \proj__8.net244 ;
 wire \proj__8.net245 ;
 wire \proj__8.net246 ;
 wire \proj__8.net247 ;
 wire \proj__8.net248 ;
 wire \proj__8.net249 ;
 wire \proj__8.net25 ;
 wire \proj__8.net250 ;
 wire \proj__8.net251 ;
 wire \proj__8.net252 ;
 wire \proj__8.net253 ;
 wire \proj__8.net254 ;
 wire \proj__8.net255 ;
 wire \proj__8.net256 ;
 wire \proj__8.net257 ;
 wire \proj__8.net258 ;
 wire \proj__8.net259 ;
 wire \proj__8.net26 ;
 wire \proj__8.net260 ;
 wire \proj__8.net261 ;
 wire \proj__8.net262 ;
 wire \proj__8.net263 ;
 wire \proj__8.net264 ;
 wire \proj__8.net265 ;
 wire \proj__8.net266 ;
 wire \proj__8.net267 ;
 wire \proj__8.net268 ;
 wire \proj__8.net269 ;
 wire \proj__8.net27 ;
 wire \proj__8.net270 ;
 wire \proj__8.net271 ;
 wire \proj__8.net272 ;
 wire \proj__8.net273 ;
 wire \proj__8.net274 ;
 wire \proj__8.net275 ;
 wire \proj__8.net276 ;
 wire \proj__8.net277 ;
 wire \proj__8.net278 ;
 wire \proj__8.net279 ;
 wire \proj__8.net28 ;
 wire \proj__8.net280 ;
 wire \proj__8.net281 ;
 wire \proj__8.net282 ;
 wire \proj__8.net283 ;
 wire \proj__8.net284 ;
 wire \proj__8.net285 ;
 wire \proj__8.net286 ;
 wire \proj__8.net287 ;
 wire \proj__8.net288 ;
 wire \proj__8.net289 ;
 wire \proj__8.net29 ;
 wire \proj__8.net290 ;
 wire \proj__8.net291 ;
 wire \proj__8.net292 ;
 wire \proj__8.net293 ;
 wire \proj__8.net294 ;
 wire \proj__8.net295 ;
 wire \proj__8.net296 ;
 wire \proj__8.net297 ;
 wire \proj__8.net298 ;
 wire \proj__8.net299 ;
 wire \proj__8.net3 ;
 wire \proj__8.net30 ;
 wire \proj__8.net300 ;
 wire \proj__8.net301 ;
 wire \proj__8.net302 ;
 wire \proj__8.net303 ;
 wire \proj__8.net304 ;
 wire \proj__8.net305 ;
 wire \proj__8.net306 ;
 wire \proj__8.net307 ;
 wire \proj__8.net308 ;
 wire \proj__8.net309 ;
 wire \proj__8.net31 ;
 wire \proj__8.net310 ;
 wire \proj__8.net311 ;
 wire \proj__8.net312 ;
 wire \proj__8.net313 ;
 wire \proj__8.net314 ;
 wire \proj__8.net315 ;
 wire \proj__8.net316 ;
 wire \proj__8.net317 ;
 wire \proj__8.net318 ;
 wire \proj__8.net319 ;
 wire \proj__8.net32 ;
 wire \proj__8.net320 ;
 wire \proj__8.net321 ;
 wire \proj__8.net322 ;
 wire \proj__8.net323 ;
 wire \proj__8.net324 ;
 wire \proj__8.net325 ;
 wire \proj__8.net326 ;
 wire \proj__8.net327 ;
 wire \proj__8.net328 ;
 wire \proj__8.net329 ;
 wire \proj__8.net33 ;
 wire \proj__8.net330 ;
 wire \proj__8.net331 ;
 wire \proj__8.net332 ;
 wire \proj__8.net333 ;
 wire \proj__8.net334 ;
 wire \proj__8.net335 ;
 wire \proj__8.net336 ;
 wire \proj__8.net337 ;
 wire \proj__8.net338 ;
 wire \proj__8.net339 ;
 wire \proj__8.net34 ;
 wire \proj__8.net340 ;
 wire \proj__8.net341 ;
 wire \proj__8.net342 ;
 wire \proj__8.net343 ;
 wire \proj__8.net344 ;
 wire \proj__8.net345 ;
 wire \proj__8.net346 ;
 wire \proj__8.net347 ;
 wire \proj__8.net348 ;
 wire \proj__8.net349 ;
 wire \proj__8.net35 ;
 wire \proj__8.net350 ;
 wire \proj__8.net351 ;
 wire \proj__8.net352 ;
 wire \proj__8.net353 ;
 wire \proj__8.net354 ;
 wire \proj__8.net355 ;
 wire \proj__8.net356 ;
 wire \proj__8.net357 ;
 wire \proj__8.net358 ;
 wire \proj__8.net359 ;
 wire \proj__8.net36 ;
 wire \proj__8.net360 ;
 wire \proj__8.net361 ;
 wire \proj__8.net362 ;
 wire \proj__8.net363 ;
 wire \proj__8.net364 ;
 wire \proj__8.net365 ;
 wire \proj__8.net366 ;
 wire \proj__8.net367 ;
 wire \proj__8.net368 ;
 wire \proj__8.net369 ;
 wire \proj__8.net37 ;
 wire \proj__8.net370 ;
 wire \proj__8.net371 ;
 wire \proj__8.net372 ;
 wire \proj__8.net373 ;
 wire \proj__8.net374 ;
 wire \proj__8.net375 ;
 wire \proj__8.net376 ;
 wire \proj__8.net377 ;
 wire \proj__8.net378 ;
 wire \proj__8.net379 ;
 wire \proj__8.net38 ;
 wire \proj__8.net380 ;
 wire \proj__8.net381 ;
 wire \proj__8.net382 ;
 wire \proj__8.net383 ;
 wire \proj__8.net384 ;
 wire \proj__8.net385 ;
 wire \proj__8.net386 ;
 wire \proj__8.net387 ;
 wire \proj__8.net388 ;
 wire \proj__8.net389 ;
 wire \proj__8.net39 ;
 wire \proj__8.net390 ;
 wire \proj__8.net391 ;
 wire \proj__8.net392 ;
 wire \proj__8.net393 ;
 wire \proj__8.net394 ;
 wire \proj__8.net395 ;
 wire \proj__8.net396 ;
 wire \proj__8.net397 ;
 wire \proj__8.net398 ;
 wire \proj__8.net399 ;
 wire \proj__8.net4 ;
 wire \proj__8.net40 ;
 wire \proj__8.net400 ;
 wire \proj__8.net401 ;
 wire \proj__8.net402 ;
 wire \proj__8.net403 ;
 wire \proj__8.net404 ;
 wire \proj__8.net405 ;
 wire \proj__8.net406 ;
 wire \proj__8.net407 ;
 wire \proj__8.net408 ;
 wire \proj__8.net409 ;
 wire \proj__8.net41 ;
 wire \proj__8.net410 ;
 wire \proj__8.net411 ;
 wire \proj__8.net412 ;
 wire \proj__8.net413 ;
 wire \proj__8.net414 ;
 wire \proj__8.net415 ;
 wire \proj__8.net416 ;
 wire \proj__8.net417 ;
 wire \proj__8.net418 ;
 wire \proj__8.net419 ;
 wire \proj__8.net42 ;
 wire \proj__8.net420 ;
 wire \proj__8.net421 ;
 wire \proj__8.net422 ;
 wire \proj__8.net423 ;
 wire \proj__8.net424 ;
 wire \proj__8.net425 ;
 wire \proj__8.net426 ;
 wire \proj__8.net427 ;
 wire \proj__8.net428 ;
 wire \proj__8.net429 ;
 wire \proj__8.net43 ;
 wire \proj__8.net430 ;
 wire \proj__8.net431 ;
 wire \proj__8.net432 ;
 wire \proj__8.net433 ;
 wire \proj__8.net434 ;
 wire \proj__8.net435 ;
 wire \proj__8.net436 ;
 wire \proj__8.net437 ;
 wire \proj__8.net438 ;
 wire \proj__8.net439 ;
 wire \proj__8.net44 ;
 wire \proj__8.net440 ;
 wire \proj__8.net441 ;
 wire \proj__8.net442 ;
 wire \proj__8.net443 ;
 wire \proj__8.net444 ;
 wire \proj__8.net445 ;
 wire \proj__8.net446 ;
 wire \proj__8.net447 ;
 wire \proj__8.net448 ;
 wire \proj__8.net449 ;
 wire \proj__8.net45 ;
 wire \proj__8.net450 ;
 wire \proj__8.net451 ;
 wire \proj__8.net452 ;
 wire \proj__8.net453 ;
 wire \proj__8.net454 ;
 wire \proj__8.net455 ;
 wire \proj__8.net456 ;
 wire \proj__8.net457 ;
 wire \proj__8.net458 ;
 wire \proj__8.net459 ;
 wire \proj__8.net46 ;
 wire \proj__8.net460 ;
 wire \proj__8.net461 ;
 wire \proj__8.net462 ;
 wire \proj__8.net463 ;
 wire \proj__8.net464 ;
 wire \proj__8.net465 ;
 wire \proj__8.net466 ;
 wire \proj__8.net467 ;
 wire \proj__8.net468 ;
 wire \proj__8.net469 ;
 wire \proj__8.net47 ;
 wire \proj__8.net470 ;
 wire \proj__8.net471 ;
 wire \proj__8.net472 ;
 wire \proj__8.net473 ;
 wire \proj__8.net474 ;
 wire \proj__8.net475 ;
 wire \proj__8.net476 ;
 wire \proj__8.net477 ;
 wire \proj__8.net478 ;
 wire \proj__8.net479 ;
 wire \proj__8.net48 ;
 wire \proj__8.net480 ;
 wire \proj__8.net49 ;
 wire \proj__8.net50 ;
 wire \proj__8.net51 ;
 wire \proj__8.net52 ;
 wire \proj__8.net53 ;
 wire \proj__8.net54 ;
 wire \proj__8.net55 ;
 wire \proj__8.net56 ;
 wire \proj__8.net57 ;
 wire \proj__8.net58 ;
 wire \proj__8.net59 ;
 wire \proj__8.net60 ;
 wire \proj__8.net61 ;
 wire \proj__8.net62 ;
 wire \proj__8.net63 ;
 wire \proj__8.net64 ;
 wire \proj__8.net65 ;
 wire \proj__8.net66 ;
 wire \proj__8.net67 ;
 wire \proj__8.net68 ;
 wire \proj__8.net69 ;
 wire \proj__8.net70 ;
 wire \proj__8.net71 ;
 wire \proj__8.net72 ;
 wire \proj__8.net73 ;
 wire \proj__8.net74 ;
 wire \proj__8.net75 ;
 wire \proj__8.net76 ;
 wire \proj__8.net77 ;
 wire \proj__8.net78 ;
 wire \proj__8.net79 ;
 wire \proj__8.net80 ;
 wire \proj__8.net81 ;
 wire \proj__8.net82 ;
 wire \proj__8.net83 ;
 wire \proj__8.net84 ;
 wire \proj__8.net85 ;
 wire \proj__8.net86 ;
 wire \proj__8.net87 ;
 wire \proj__8.net88 ;
 wire \proj__8.net89 ;
 wire \proj__8.net90 ;
 wire \proj__8.net91 ;
 wire \proj__8.net92 ;
 wire \proj__8.net93 ;
 wire \proj__8.net94 ;
 wire \proj__8.net95 ;
 wire \proj__8.net96 ;
 wire \proj__8.net97 ;
 wire \proj__8.net98 ;
 wire \proj__8.net99 ;
 wire \proj__9.net10 ;
 wire \proj__9.net11 ;
 wire \proj__9.net12 ;
 wire \proj__9.net17 ;
 wire \proj__9.net18 ;
 wire \proj__9.net19 ;
 wire \proj__9.net20 ;
 wire \proj__9.net21 ;
 wire \proj__9.net22 ;
 wire \proj__9.net23 ;
 wire \proj__9.net24 ;
 wire \proj__9.net25 ;
 wire \proj__9.net26 ;
 wire \proj__9.net27 ;
 wire \proj__9.net28 ;
 wire \proj__9.net7 ;
 wire \proj__9.net8 ;
 wire \proj__9.net9 ;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire \proj_11.flop1/_0_ ;
 wire \proj_11.flop1/_1_ ;
 wire net34;
 wire net35;
 wire \proj_11.flop2/_0_ ;
 wire \proj_11.flop2/_1_ ;
 wire net36;
 wire net37;
 wire \proj_11.flop3/_0_ ;
 wire \proj_11.flop3/_1_ ;
 wire net38;
 wire net39;
 wire \proj_11.flop4/_0_ ;
 wire \proj_11.flop4/_1_ ;
 wire net40;
 wire net41;
 wire \proj_11.flop5/_0_ ;
 wire \proj_11.flop5/_1_ ;
 wire net42;
 wire net43;
 wire \proj_11.flop6/_0_ ;
 wire \proj_11.flop6/_1_ ;
 wire net44;
 wire net45;
 wire \proj_11.flop7/_0_ ;
 wire \proj_11.flop7/_1_ ;
 wire net46;
 wire net47;
 wire \proj_11.flop8/_0_ ;
 wire \proj_11.flop8/_1_ ;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire \proj__8.flop10/notq ;
 wire net52;
 wire \proj__8.flop11/notq ;
 wire net53;
 wire net54;
 wire \proj__8.flop13/notq ;
 wire net55;
 wire \proj__8.flop14/notq ;
 wire net56;
 wire \proj__8.flop15/notq ;
 wire net57;
 wire net58;
 wire \proj__8.flop17/notq ;
 wire net59;
 wire \proj__8.flop18/notq ;
 wire net60;
 wire \proj__8.flop19/notq ;
 wire net82;
 wire net83;
 wire \proj__8.flop21/notq ;
 wire net84;
 wire \proj__8.flop22/notq ;
 wire net85;
 wire \proj__8.flop23/notq ;
 wire net86;
 wire net87;
 wire \proj__8.flop25/notq ;
 wire net88;
 wire \proj__8.flop26/notq ;
 wire net89;
 wire \proj__8.flop27/notq ;
 wire net90;
 wire net91;
 wire \proj__8.flop29/notq ;
 wire net92;
 wire \proj__8.flop30/notq ;
 wire net93;
 wire \proj__8.flop31/notq ;
 wire net94;
 wire net95;
 wire \proj__8.flop33/notq ;
 wire net96;
 wire \proj__8.flop34/notq ;
 wire net97;
 wire \proj__8.flop35/notq ;
 wire net98;
 wire net99;
 wire \proj__8.flop37/notq ;
 wire net100;
 wire \proj__8.flop38/notq ;
 wire net101;
 wire \proj__8.flop39/notq ;
 wire net102;
 wire net103;
 wire \proj__8.flop41/notq ;
 wire net104;
 wire \proj__8.flop6/notq ;
 wire net105;
 wire \proj__8.flop7/notq ;
 wire net106;
 wire net107;
 wire \proj__8.flop9/notq ;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net108;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_1_0__leaf_clk_regs;
 wire clknet_1_1__leaf_clk_regs;
 wire net109;
 wire net110;

 sg13g2_inv_1 _076_ (.Y(_039_),
    .A(net6));
 sg13g2_inv_1 _077_ (.Y(_040_),
    .A(\proj__0.net9 ));
 sg13g2_inv_1 _078_ (.Y(_041_),
    .A(\proj__0.net10 ));
 sg13g2_inv_1 _079_ (.Y(_042_),
    .A(\proj__0.net11 ));
 sg13g2_nor2_1 _080_ (.A(net8),
    .B(net7),
    .Y(_043_));
 sg13g2_nor2_2 _081_ (.A(net5),
    .B(net6),
    .Y(_044_));
 sg13g2_nor4_2 _082_ (.A(net5),
    .B(net6),
    .C(net8),
    .Y(_045_),
    .D(net7));
 sg13g2_nor2b_2 _083_ (.A(net8),
    .B_N(net7),
    .Y(_046_));
 sg13g2_nor2b_2 _084_ (.A(net5),
    .B_N(net6),
    .Y(_047_));
 sg13g2_and2_2 _085_ (.A(_046_),
    .B(_047_),
    .X(_048_));
 sg13g2_and3_2 _086_ (.X(_049_),
    .A(net8),
    .B(net7),
    .C(_044_));
 sg13g2_nor2b_2 _087_ (.A(net7),
    .B_N(net8),
    .Y(_050_));
 sg13g2_nor2b_1 _088_ (.A(net6),
    .B_N(net5),
    .Y(_051_));
 sg13g2_and2_2 _089_ (.A(_050_),
    .B(_051_),
    .X(_052_));
 sg13g2_and2_1 _090_ (.A(_046_),
    .B(_051_),
    .X(_053_));
 sg13g2_nand4_1 _091_ (.B(net7),
    .C(\proj_14.net9 ),
    .A(net8),
    .Y(_054_),
    .D(_047_));
 sg13g2_and2_1 _092_ (.A(net5),
    .B(net6),
    .X(_055_));
 sg13g2_and2_2 _093_ (.A(_050_),
    .B(_055_),
    .X(_056_));
 sg13g2_and2_1 _094_ (.A(_044_),
    .B(_046_),
    .X(_057_));
 sg13g2_nand3_1 _095_ (.B(_047_),
    .C(_050_),
    .A(\proj_10.net4 ),
    .Y(_058_));
 sg13g2_and2_1 _096_ (.A(_046_),
    .B(_055_),
    .X(_059_));
 sg13g2_a21oi_1 _097_ (.A1(\proj__7.net8 ),
    .A2(_059_),
    .Y(_060_),
    .B1(_045_));
 sg13g2_and2_2 _098_ (.A(_043_),
    .B(_055_),
    .X(_061_));
 sg13g2_and2_1 _099_ (.A(_043_),
    .B(_047_),
    .X(_062_));
 sg13g2_nand2_1 _100_ (.Y(_063_),
    .A(_054_),
    .B(_058_));
 sg13g2_a221oi_1 _101_ (.B2(\proj__3.net9 ),
    .C1(_063_),
    .B1(_061_),
    .A1(\proj__4.net10 ),
    .Y(_064_),
    .A2(_057_));
 sg13g2_a22oi_1 _102_ (.Y(_065_),
    .B1(_056_),
    .B2(\proj_11.net3 ),
    .A2(_048_),
    .A1(\proj__6.net10 ));
 sg13g2_a22oi_1 _103_ (.Y(_066_),
    .B1(_062_),
    .B2(\proj__2.net4 ),
    .A2(_052_),
    .A1(\proj__9.net7 ));
 sg13g2_a22oi_1 _104_ (.Y(_067_),
    .B1(_053_),
    .B2(\proj__5.net9 ),
    .A2(_049_),
    .A1(\proj_12.net9 ));
 sg13g2_and4_1 _105_ (.A(_060_),
    .B(_065_),
    .C(_066_),
    .D(_067_),
    .X(_000_));
 sg13g2_a22oi_1 _106_ (.Y(uo_out[0]),
    .B1(_064_),
    .B2(_000_),
    .A2(_045_),
    .A1(_040_));
 sg13g2_a22oi_1 _107_ (.Y(_001_),
    .B1(_061_),
    .B2(\proj__3.net10 ),
    .A2(_053_),
    .A1(\proj__5.net10 ));
 sg13g2_nand3_1 _108_ (.B(_044_),
    .C(_050_),
    .A(\proj__8.net3 ),
    .Y(_002_));
 sg13g2_nand3_1 _109_ (.B(_047_),
    .C(_050_),
    .A(\proj_10.net5 ),
    .Y(_003_));
 sg13g2_and4_1 _110_ (.A(net8),
    .B(net7),
    .C(net3),
    .D(_055_),
    .X(_004_));
 sg13g2_a22oi_1 _111_ (.Y(_005_),
    .B1(_062_),
    .B2(\proj__2.net5 ),
    .A2(_052_),
    .A1(\proj__9.net8 ));
 sg13g2_and3_1 _112_ (.X(_006_),
    .A(_060_),
    .B(_001_),
    .C(_005_));
 sg13g2_a221oi_1 _113_ (.B2(\proj_11.net4 ),
    .C1(_004_),
    .B1(_056_),
    .A1(\proj_12.net10 ),
    .Y(_007_),
    .A2(_049_));
 sg13g2_a22oi_1 _114_ (.Y(_008_),
    .B1(_057_),
    .B2(net108),
    .A2(_048_),
    .A1(\proj__6.net11 ));
 sg13g2_and4_1 _115_ (.A(_002_),
    .B(_003_),
    .C(_007_),
    .D(_008_),
    .X(_009_));
 sg13g2_a22oi_1 _116_ (.Y(uo_out[1]),
    .B1(_006_),
    .B2(_009_),
    .A2(_045_),
    .A1(_041_));
 sg13g2_nand2_1 _117_ (.Y(_010_),
    .A(\proj__4.net12 ),
    .B(_057_));
 sg13g2_nand2_1 _118_ (.Y(_011_),
    .A(\proj__9.net9 ),
    .B(_052_));
 sg13g2_nand2_1 _119_ (.Y(_012_),
    .A(\proj__6.net12 ),
    .B(_048_));
 sg13g2_a22oi_1 _120_ (.Y(_013_),
    .B1(_061_),
    .B2(\proj__3.net11 ),
    .A2(_056_),
    .A1(\proj_11.net5 ));
 sg13g2_and3_1 _121_ (.X(_014_),
    .A(_010_),
    .B(_012_),
    .C(_013_));
 sg13g2_a22oi_1 _122_ (.Y(_015_),
    .B1(_053_),
    .B2(net72),
    .A2(_049_),
    .A1(\proj_12.net11 ));
 sg13g2_and4_1 _123_ (.A(_060_),
    .B(_002_),
    .C(_011_),
    .D(_015_),
    .X(_016_));
 sg13g2_a22oi_1 _124_ (.Y(uo_out[2]),
    .B1(_014_),
    .B2(_016_),
    .A2(_045_),
    .A1(_042_));
 sg13g2_a22oi_1 _125_ (.Y(_017_),
    .B1(_061_),
    .B2(\proj__3.net12 ),
    .A2(_053_),
    .A1(net70));
 sg13g2_a22oi_1 _126_ (.Y(_018_),
    .B1(_057_),
    .B2(\proj__4.net13 ),
    .A2(_048_),
    .A1(net62));
 sg13g2_nand3_1 _127_ (.B(_043_),
    .C(_051_),
    .A(\proj__1.net7 ),
    .Y(_019_));
 sg13g2_a22oi_1 _128_ (.Y(_020_),
    .B1(_059_),
    .B2(\proj__7.net9 ),
    .A2(_056_),
    .A1(\proj_11.net6 ));
 sg13g2_a22oi_1 _129_ (.Y(_021_),
    .B1(_052_),
    .B2(\proj__9.net10 ),
    .A2(_049_),
    .A1(\proj_12.net12 ));
 sg13g2_and4_1 _130_ (.A(_002_),
    .B(_019_),
    .C(_020_),
    .D(_021_),
    .X(_022_));
 sg13g2_nand3_1 _131_ (.B(_018_),
    .C(_022_),
    .A(_017_),
    .Y(uo_out[3]));
 sg13g2_a21o_1 _132_ (.A2(_046_),
    .A1(_039_),
    .B1(_045_),
    .X(_023_));
 sg13g2_o21ai_1 _133_ (.B1(net67),
    .Y(_024_),
    .A1(_059_),
    .A2(_023_));
 sg13g2_nand2_1 _134_ (.Y(_025_),
    .A(\proj__9.net11 ),
    .B(_052_));
 sg13g2_a22oi_1 _135_ (.Y(_026_),
    .B1(_049_),
    .B2(\proj_12.net13 ),
    .A2(_048_),
    .A1(clknet_1_0__leaf_clk));
 sg13g2_a22oi_1 _136_ (.Y(_027_),
    .B1(_061_),
    .B2(\proj__3.net13 ),
    .A2(_056_),
    .A1(\proj_11.net7 ));
 sg13g2_nand4_1 _137_ (.B(_025_),
    .C(_026_),
    .A(_002_),
    .Y(_028_),
    .D(_027_));
 sg13g2_nand2b_1 _138_ (.Y(uo_out[4]),
    .B(_024_),
    .A_N(_028_));
 sg13g2_nand2_1 _139_ (.Y(_029_),
    .A(\proj__7.net10 ),
    .B(_059_));
 sg13g2_a22oi_1 _140_ (.Y(_030_),
    .B1(_052_),
    .B2(\proj__9.net12 ),
    .A2(_049_),
    .A1(\proj_12.net14 ));
 sg13g2_a22oi_1 _141_ (.Y(_031_),
    .B1(_061_),
    .B2(\proj__3.net14 ),
    .A2(_056_),
    .A1(\proj_11.net8 ));
 sg13g2_nand4_1 _142_ (.B(_029_),
    .C(_030_),
    .A(_002_),
    .Y(_032_),
    .D(_031_));
 sg13g2_a21o_1 _143_ (.A2(_023_),
    .A1(net64),
    .B1(_032_),
    .X(uo_out[5]));
 sg13g2_or2_1 _144_ (.X(_033_),
    .B(_023_),
    .A(_061_));
 sg13g2_nand2_1 _145_ (.Y(_034_),
    .A(net63),
    .B(_033_));
 sg13g2_a22oi_1 _146_ (.Y(_035_),
    .B1(_056_),
    .B2(\proj_11.net9 ),
    .A2(_049_),
    .A1(\proj_12.net15 ));
 sg13g2_nand3_1 _147_ (.B(_034_),
    .C(_035_),
    .A(_029_),
    .Y(uo_out[6]));
 sg13g2_nand2_1 _148_ (.Y(_036_),
    .A(net61),
    .B(_033_));
 sg13g2_nand3_1 _149_ (.B(_044_),
    .C(_050_),
    .A(\proj__8.net4 ),
    .Y(_037_));
 sg13g2_a22oi_1 _150_ (.Y(_038_),
    .B1(_056_),
    .B2(\proj_11.net10 ),
    .A2(_049_),
    .A1(\proj_12.net16 ));
 sg13g2_nand4_1 _151_ (.B(_036_),
    .C(_037_),
    .A(_029_),
    .Y(uo_out[7]),
    .D(_038_));
 sg13g2_tielo \proj_11.flop2/_5__10  (.L_LO(net10));
 sg13g2_tielo \proj_11.flop3/_5__11  (.L_LO(net11));
 sg13g2_tielo \proj_11.flop4/_5__12  (.L_LO(net12));
 sg13g2_tielo \proj_11.flop5/_5__13  (.L_LO(net13));
 sg13g2_tielo \proj_11.flop6/_5__14  (.L_LO(net14));
 sg13g2_tielo \proj_11.flop7/_5__15  (.L_LO(net15));
 sg13g2_tielo \proj_11.flop8/_5__16  (.L_LO(net16));
 sg13g2_tielo tt_um_wokwi_group_1_17 (.L_LO(net17));
 sg13g2_tielo tt_um_wokwi_group_1_18 (.L_LO(net18));
 sg13g2_tielo tt_um_wokwi_group_1_19 (.L_LO(net19));
 sg13g2_tielo tt_um_wokwi_group_1_20 (.L_LO(net20));
 sg13g2_tielo tt_um_wokwi_group_1_21 (.L_LO(net21));
 sg13g2_tielo tt_um_wokwi_group_1_22 (.L_LO(net22));
 sg13g2_tielo tt_um_wokwi_group_1_23 (.L_LO(net23));
 sg13g2_tielo tt_um_wokwi_group_1_24 (.L_LO(net24));
 sg13g2_tielo tt_um_wokwi_group_1_25 (.L_LO(net25));
 sg13g2_tielo tt_um_wokwi_group_1_26 (.L_LO(net26));
 sg13g2_tielo tt_um_wokwi_group_1_27 (.L_LO(net27));
 sg13g2_tielo tt_um_wokwi_group_1_28 (.L_LO(net28));
 sg13g2_tielo tt_um_wokwi_group_1_29 (.L_LO(net29));
 sg13g2_tielo tt_um_wokwi_group_1_30 (.L_LO(net30));
 sg13g2_tielo tt_um_wokwi_group_1_31 (.L_LO(net31));
 sg13g2_tielo tt_um_wokwi_group_1_32 (.L_LO(net32));
 sg13g2_tielo \proj_11.flop1/dffsr_33  (.L_LO(net33));
 sg13g2_and2_1 \proj_10.and1/_0_  (.A(net73),
    .B(\proj_10.net7 ),
    .X(\proj_10.net8 ));
 sg13g2_and2_1 \proj_10.and2/_0_  (.A(net75),
    .B(net80),
    .X(\proj_10.net9 ));
 sg13g2_or2_1 \proj_10.or1/_0_  (.X(\proj_10.net5 ),
    .B(\proj_10.net8 ),
    .A(\proj_10.net9 ));
 sg13g2_xor2_1 \proj_10.xor1/_0_  (.B(net80),
    .A(net75),
    .X(\proj_10.net7 ));
 sg13g2_xor2_1 \proj_10.xor2/_0_  (.B(\proj_10.net7 ),
    .A(net73),
    .X(\proj_10.net4 ));
 sg13g2_inv_1 \proj_11.flop1/_4_  (.Y(\proj_11.flop1/_0_ ),
    .A(\proj_11.net18 ));
 sg13g2_inv_1 \proj_11.flop1/_5_  (.Y(\proj_11.flop1/_1_ ),
    .A(net9));
 sg13g2_tielo \proj_11.flop1/dffsr_34  (.L_LO(net34));
 sg13g2_tielo \proj_11.flop2/dffsr_35  (.L_LO(net35));
 sg13g2_sdfbbp_1 \proj_11.flop1/dffsr  (.Q(\proj_11.net4 ),
    .Q_N(\proj_11.net19 ),
    .RESET_B(\proj_11.flop1/_0_ ),
    .SET_B(\proj_11.flop1/_1_ ),
    .D(\proj_11.net19 ),
    .SCE(net34),
    .SCD(net33),
    .CLK(\proj_11.net3 ));
 sg13g2_inv_1 \proj_11.flop2/_4_  (.Y(\proj_11.flop2/_0_ ),
    .A(\proj_11.net18 ));
 sg13g2_inv_1 \proj_11.flop2/_5_  (.Y(\proj_11.flop2/_1_ ),
    .A(net10));
 sg13g2_tielo \proj_11.flop2/dffsr_36  (.L_LO(net36));
 sg13g2_tielo \proj_11.flop3/dffsr_37  (.L_LO(net37));
 sg13g2_sdfbbp_1 \proj_11.flop2/dffsr  (.Q(\proj_11.net5 ),
    .Q_N(\proj_11.net20 ),
    .RESET_B(\proj_11.flop2/_0_ ),
    .SET_B(\proj_11.flop2/_1_ ),
    .D(\proj_11.net20 ),
    .SCE(net36),
    .SCD(net35),
    .CLK(\proj_11.net4 ));
 sg13g2_inv_1 \proj_11.flop3/_4_  (.Y(\proj_11.flop3/_0_ ),
    .A(\proj_11.net18 ));
 sg13g2_inv_1 \proj_11.flop3/_5_  (.Y(\proj_11.flop3/_1_ ),
    .A(net11));
 sg13g2_tielo \proj_11.flop3/dffsr_38  (.L_LO(net38));
 sg13g2_tielo \proj_11.flop4/dffsr_39  (.L_LO(net39));
 sg13g2_sdfbbp_1 \proj_11.flop3/dffsr  (.Q(\proj_11.net6 ),
    .Q_N(\proj_11.net21 ),
    .RESET_B(\proj_11.flop3/_0_ ),
    .SET_B(\proj_11.flop3/_1_ ),
    .D(\proj_11.net21 ),
    .SCE(net38),
    .SCD(net37),
    .CLK(\proj_11.net5 ));
 sg13g2_inv_1 \proj_11.flop4/_4_  (.Y(\proj_11.flop4/_0_ ),
    .A(\proj_11.net18 ));
 sg13g2_inv_1 \proj_11.flop4/_5_  (.Y(\proj_11.flop4/_1_ ),
    .A(net12));
 sg13g2_tielo \proj_11.flop4/dffsr_40  (.L_LO(net40));
 sg13g2_tielo \proj_11.flop5/dffsr_41  (.L_LO(net41));
 sg13g2_sdfbbp_1 \proj_11.flop4/dffsr  (.Q(\proj_11.net3 ),
    .Q_N(\proj_11.net16 ),
    .RESET_B(\proj_11.flop4/_0_ ),
    .SET_B(\proj_11.flop4/_1_ ),
    .D(net110),
    .SCE(net40),
    .SCD(net39),
    .CLK(clknet_1_1__leaf_clk_regs));
 sg13g2_inv_1 \proj_11.flop5/_4_  (.Y(\proj_11.flop5/_0_ ),
    .A(\proj_11.net18 ));
 sg13g2_inv_1 \proj_11.flop5/_5_  (.Y(\proj_11.flop5/_1_ ),
    .A(net13));
 sg13g2_tielo \proj_11.flop5/dffsr_42  (.L_LO(net42));
 sg13g2_tielo \proj_11.flop6/dffsr_43  (.L_LO(net43));
 sg13g2_sdfbbp_1 \proj_11.flop5/dffsr  (.Q(\proj_11.net7 ),
    .Q_N(\proj_11.net22 ),
    .RESET_B(\proj_11.flop5/_0_ ),
    .SET_B(\proj_11.flop5/_1_ ),
    .D(\proj_11.net22 ),
    .SCE(net42),
    .SCD(net41),
    .CLK(\proj_11.net6 ));
 sg13g2_inv_1 \proj_11.flop6/_4_  (.Y(\proj_11.flop6/_0_ ),
    .A(\proj_11.net18 ));
 sg13g2_inv_1 \proj_11.flop6/_5_  (.Y(\proj_11.flop6/_1_ ),
    .A(net14));
 sg13g2_tielo \proj_11.flop6/dffsr_44  (.L_LO(net44));
 sg13g2_tielo \proj_11.flop7/dffsr_45  (.L_LO(net45));
 sg13g2_sdfbbp_1 \proj_11.flop6/dffsr  (.Q(\proj_11.net9 ),
    .Q_N(\proj_11.net23 ),
    .RESET_B(\proj_11.flop6/_0_ ),
    .SET_B(\proj_11.flop6/_1_ ),
    .D(\proj_11.net23 ),
    .SCE(net44),
    .SCD(net43),
    .CLK(\proj_11.net8 ));
 sg13g2_inv_1 \proj_11.flop7/_4_  (.Y(\proj_11.flop7/_0_ ),
    .A(\proj_11.net18 ));
 sg13g2_inv_1 \proj_11.flop7/_5_  (.Y(\proj_11.flop7/_1_ ),
    .A(net15));
 sg13g2_tielo \proj_11.flop7/dffsr_46  (.L_LO(net46));
 sg13g2_tielo \proj_11.flop8/dffsr_47  (.L_LO(net47));
 sg13g2_sdfbbp_1 \proj_11.flop7/dffsr  (.Q(\proj_11.net8 ),
    .Q_N(\proj_11.net24 ),
    .RESET_B(\proj_11.flop7/_0_ ),
    .SET_B(\proj_11.flop7/_1_ ),
    .D(\proj_11.net24 ),
    .SCE(net46),
    .SCD(net45),
    .CLK(\proj_11.net7 ));
 sg13g2_inv_1 \proj_11.flop8/_4_  (.Y(\proj_11.flop8/_0_ ),
    .A(\proj_11.net18 ));
 sg13g2_inv_1 \proj_11.flop8/_5_  (.Y(\proj_11.flop8/_1_ ),
    .A(net16));
 sg13g2_tielo \proj_11.flop8/dffsr_48  (.L_LO(net48));
 sg13g2_tiehi \proj__8.flop1/_1__49  (.L_HI(net49));
 sg13g2_sdfbbp_1 \proj_11.flop8/dffsr  (.Q(\proj_11.net10 ),
    .Q_N(\proj_11.net25 ),
    .RESET_B(\proj_11.flop8/_0_ ),
    .SET_B(\proj_11.flop8/_1_ ),
    .D(\proj_11.net25 ),
    .SCE(net48),
    .SCD(net47),
    .CLK(\proj_11.net9 ));
 sg13g2_inv_2 \proj_11.not1/_0_  (.Y(\proj_11.net18 ),
    .A(net1));
 sg13g2_and2_1 \proj_12.and1/_0_  (.A(net63),
    .B(net61),
    .X(\proj_12.net45 ));
 sg13g2_and2_1 \proj_12.and2/_0_  (.A(\proj_12.net47 ),
    .B(\proj_12.net46 ),
    .X(\proj_12.net16 ));
 sg13g2_and2_1 \proj_12.and3/_0_  (.A(net71),
    .B(net69),
    .X(\proj_12.net48 ));
 sg13g2_and2_1 \proj_12.and4/_0_  (.A(\proj_12.net49 ),
    .B(\proj_12.net48 ),
    .X(\proj_12.net47 ));
 sg13g2_and2_1 \proj_12.and5/_0_  (.A(\proj_12.net50 ),
    .B(\proj_12.net45 ),
    .X(\proj_12.net46 ));
 sg13g2_and2_1 \proj_12.and6/_0_  (.A(net81),
    .B(net74),
    .X(\proj_12.net49 ));
 sg13g2_and2_1 \proj_12.and7/_0_  (.A(net67),
    .B(net64),
    .X(\proj_12.net50 ));
 sg13g2_or2_1 \proj_12.or1/_0_  (.X(\proj_12.net11 ),
    .B(\proj_12.net22 ),
    .A(\proj_12.net23 ));
 sg13g2_or2_1 \proj_12.or10/_0_  (.X(\proj_12.net22 ),
    .B(\proj_12.net30 ),
    .A(\proj_12.net31 ));
 sg13g2_or2_1 \proj_12.or11/_0_  (.X(\proj_12.net32 ),
    .B(net66),
    .A(net63));
 sg13g2_or2_1 \proj_12.or12/_0_  (.X(\proj_12.net30 ),
    .B(net78),
    .A(net72));
 sg13g2_or2_1 \proj_12.or13/_0_  (.X(\proj_12.net23 ),
    .B(\proj_12.net32 ),
    .A(net62));
 sg13g2_or2_1 \proj_12.or14/_0_  (.X(\proj_12.net31 ),
    .B(net70),
    .A(net68));
 sg13g2_or2_1 \proj_12.or15/_0_  (.X(\proj_12.net35 ),
    .B(\proj_12.net33 ),
    .A(\proj_12.net34 ));
 sg13g2_or2_1 \proj_12.or16/_0_  (.X(\proj_12.net10 ),
    .B(\proj_12.net35 ),
    .A(\proj_12.net36 ));
 sg13g2_or2_1 \proj_12.or17/_0_  (.X(\proj_12.net36 ),
    .B(net63),
    .A(net62));
 sg13g2_or2_1 \proj_12.or18/_0_  (.X(\proj_12.net34 ),
    .B(net73),
    .A(net70));
 sg13g2_or2_1 \proj_12.or19/_0_  (.X(\proj_12.net33 ),
    .B(net77),
    .A(net81));
 sg13g2_or2_1 \proj_12.or2/_0_  (.X(\proj_12.net26 ),
    .B(\proj_12.net24 ),
    .A(\proj_12.net25 ));
 sg13g2_or2_1 \proj_12.or20/_0_  (.X(\proj_12.net39 ),
    .B(\proj_12.net37 ),
    .A(\proj_12.net38 ));
 sg13g2_or2_1 \proj_12.or21/_0_  (.X(\proj_12.net12 ),
    .B(\proj_12.net39 ),
    .A(net61));
 sg13g2_or2_1 \proj_12.or22/_0_  (.X(\proj_12.net38 ),
    .B(net68),
    .A(net64));
 sg13g2_or2_1 \proj_12.or23/_0_  (.X(\proj_12.net37 ),
    .B(net74),
    .A(net71));
 sg13g2_or2_1 \proj_12.or24/_0_  (.X(\proj_12.net40 ),
    .B(net65),
    .A(net61));
 sg13g2_or2_1 \proj_12.or25/_0_  (.X(\proj_12.net14 ),
    .B(\proj_12.net29 ),
    .A(\proj_12.net40 ));
 sg13g2_or2_1 \proj_12.or26/_0_  (.X(\proj_12.net43 ),
    .B(\proj_12.net41 ),
    .A(\proj_12.net42 ));
 sg13g2_or2_1 \proj_12.or27/_0_  (.X(\proj_12.net15 ),
    .B(\proj_12.net43 ),
    .A(\proj_12.net44 ));
 sg13g2_or2_1 \proj_12.or28/_0_  (.X(\proj_12.net44 ),
    .B(net64),
    .A(net61));
 sg13g2_or2_1 \proj_12.or29/_0_  (.X(\proj_12.net42 ),
    .B(net69),
    .A(net67));
 sg13g2_or2_1 \proj_12.or3/_0_  (.X(\proj_12.net9 ),
    .B(\proj_12.net26 ),
    .A(\proj_12.net27 ));
 sg13g2_or2_1 \proj_12.or30/_0_  (.X(\proj_12.net41 ),
    .B(net74),
    .A(net71));
 sg13g2_or2_1 \proj_12.or4/_0_  (.X(\proj_12.net13 ),
    .B(\proj_12.net28 ),
    .A(net61));
 sg13g2_or2_1 \proj_12.or5/_0_  (.X(\proj_12.net28 ),
    .B(net74),
    .A(net66));
 sg13g2_or2_1 \proj_12.or6/_0_  (.X(\proj_12.net27 ),
    .B(net63),
    .A(net62));
 sg13g2_or2_1 \proj_12.or7/_0_  (.X(\proj_12.net25 ),
    .B(net68),
    .A(net66));
 sg13g2_or2_1 \proj_12.or8/_0_  (.X(\proj_12.net24 ),
    .B(net74),
    .A(net72));
 sg13g2_or2_1 \proj_12.or9/_0_  (.X(\proj_12.net29 ),
    .B(net69),
    .A(net67));
 sg13g2_xor2_1 \proj_14.xor1/_0_  (.B(net80),
    .A(net75),
    .X(\proj_14.net15 ));
 sg13g2_xor2_1 \proj_14.xor2/_0_  (.B(net73),
    .A(net70),
    .X(\proj_14.net16 ));
 sg13g2_xor2_1 \proj_14.xor3/_0_  (.B(net68),
    .A(net66),
    .X(\proj_14.net17 ));
 sg13g2_xor2_1 \proj_14.xor4/_0_  (.B(net63),
    .A(net62),
    .X(\proj_14.net18 ));
 sg13g2_xor2_1 \proj_14.xor5/_0_  (.B(\proj_14.net15 ),
    .A(\proj_14.net16 ),
    .X(\proj_14.net19 ));
 sg13g2_xor2_1 \proj_14.xor6/_0_  (.B(\proj_14.net17 ),
    .A(\proj_14.net18 ),
    .X(\proj_14.net20 ));
 sg13g2_xor2_1 \proj_14.xor7/_0_  (.B(\proj_14.net19 ),
    .A(\proj_14.net20 ),
    .X(\proj_14.net9 ));
 sg13g2_and2_1 \proj__0.and2/_0_  (.A(net76),
    .B(net78),
    .X(\proj__0.net9 ));
 sg13g2_and2_1 \proj__0.and3/_0_  (.A(net70),
    .B(net72),
    .X(\proj__0.net10 ));
 sg13g2_or2_1 \proj__0.or1/_0_  (.X(\proj__0.net11 ),
    .B(\proj__0.net9 ),
    .A(\proj__0.net10 ));
 sg13g2_mux2_1 \proj__1.mux1/_0_  (.A0(net81),
    .A1(net74),
    .S(net66),
    .X(\proj__1.net13 ));
 sg13g2_mux2_1 \proj__1.mux3/_0_  (.A0(\proj__1.net13 ),
    .A1(\proj__1.net14 ),
    .S(net68),
    .X(\proj__1.net7 ));
 sg13g2_mux2_1 \proj__1.mux4/_0_  (.A0(net71),
    .A1(net69),
    .S(net65),
    .X(\proj__1.net14 ));
 sg13g2_and2_1 \proj__2.and3/_0_  (.A(\proj__2.net11 ),
    .B(net72),
    .X(\proj__2.net12 ));
 sg13g2_and2_1 \proj__2.and4/_0_  (.A(net79),
    .B(net75),
    .X(\proj__2.net13 ));
 sg13g2_or2_1 \proj__2.or1/_0_  (.X(\proj__2.net5 ),
    .B(\proj__2.net12 ),
    .A(\proj__2.net13 ));
 sg13g2_xor2_1 \proj__2.xor1/_0_  (.B(net79),
    .A(net75),
    .X(\proj__2.net11 ));
 sg13g2_xor2_1 \proj__2.xor2/_0_  (.B(\proj__2.net11 ),
    .A(net72),
    .X(\proj__2.net4 ));
 sg13g2_inv_1 \proj__3.not1/_0_  (.Y(\proj__3.net12 ),
    .A(net69));
 sg13g2_inv_1 \proj__3.not2/_0_  (.Y(\proj__3.net11 ),
    .A(net71));
 sg13g2_inv_1 \proj__3.not3/_0_  (.Y(\proj__3.net13 ),
    .A(net67));
 sg13g2_inv_1 \proj__3.not4/_0_  (.Y(\proj__3.net9 ),
    .A(net78));
 sg13g2_inv_1 \proj__3.not5/_0_  (.Y(\proj__3.net10 ),
    .A(net76));
 sg13g2_inv_1 \proj__3.not6/_0_  (.Y(\proj__3.net14 ),
    .A(net64));
 sg13g2_and2_1 \proj__4.and1/_0_  (.A(net78),
    .B(clknet_1_1__leaf_clk),
    .X(\proj__4.net10 ));
 sg13g2_nand2_1 \proj__4.nand1/_0_  (.Y(\proj__4.net13 ),
    .A(net71),
    .B(net74));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_or2_1 \proj__4.or1/_0_  (.X(\proj__4.net12 ),
    .B(net107),
    .A(net70));
 sg13g2_nand2_1 \proj__5.nand1/_0_  (.Y(\proj__5.net9 ),
    .A(net76),
    .B(net78));
 sg13g2_or2_1 \proj__5.or1/_0_  (.X(\proj__5.net10 ),
    .B(net78),
    .A(net76));
 sg13g2_or2_1 \proj__6.or1/_0_  (.X(\proj__6.net17 ),
    .B(net81),
    .A(net73));
 sg13g2_or2_1 \proj__6.or2/_0_  (.X(\proj__6.net18 ),
    .B(net68),
    .A(net4));
 sg13g2_or2_1 \proj__6.or3/_0_  (.X(\proj__6.net19 ),
    .B(net74),
    .A(net71));
 sg13g2_or2_1 \proj__6.or4/_0_  (.X(\proj__6.net20 ),
    .B(net66),
    .A(net4));
 sg13g2_or2_1 \proj__6.or5/_0_  (.X(\proj__6.net21 ),
    .B(net69),
    .A(net68));
 sg13g2_or2_1 \proj__6.or6/_0_  (.X(\proj__6.net22 ),
    .B(net64),
    .A(net63));
 sg13g2_or2_1 \proj__6.or7/_0_  (.X(\proj__6.net23 ),
    .B(\proj__6.net17 ),
    .A(\proj__6.net18 ));
 sg13g2_or2_1 \proj__6.or8/_0_  (.X(\proj__6.net24 ),
    .B(\proj__6.net19 ),
    .A(\proj__6.net20 ));
 sg13g2_or2_1 \proj__6.or9/_0_  (.X(\proj__6.net25 ),
    .B(\proj__6.net21 ),
    .A(\proj__6.net22 ));
 sg13g2_xor2_1 \proj__6.xor1/_0_  (.B(\proj__6.net23 ),
    .A(net62),
    .X(\proj__6.net10 ));
 sg13g2_xor2_1 \proj__6.xor2/_0_  (.B(\proj__6.net24 ),
    .A(net62),
    .X(\proj__6.net11 ));
 sg13g2_xor2_1 \proj__6.xor3/_0_  (.B(\proj__6.net25 ),
    .A(net61),
    .X(\proj__6.net12 ));
 sg13g2_and2_1 \proj__7.and1/_0_  (.A(net73),
    .B(net77),
    .X(\proj__7.net8 ));
 sg13g2_mux2_1 \proj__7.mux1/_0_  (.A0(net65),
    .A1(net63),
    .S(net61),
    .X(\proj__7.net10 ));
 sg13g2_inv_1 \proj__7.not1/_0_  (.Y(\proj__7.net9 ),
    .A(net69));
 sg13g2_dfrbp_1 \proj__8.flop1/_1_  (.CLK(\proj__8.net10 ),
    .RESET_B(net49),
    .D(net81),
    .Q_N(\proj__8.net11 ),
    .Q(\proj__8.net3 ));
 sg13g2_tiehi \proj__8.flop10/_1__50  (.L_HI(net50));
 sg13g2_dfrbp_1 \proj__8.flop10/_1_  (.CLK(\proj__8.net25 ),
    .RESET_B(net50),
    .D(\proj__8.net26 ),
    .Q_N(\proj__8.flop10/notq ),
    .Q(\proj__8.net27 ));
 sg13g2_tiehi \proj__8.flop11/_1__51  (.L_HI(net51));
 sg13g2_dfrbp_1 \proj__8.flop11/_1_  (.CLK(\proj__8.net29 ),
    .RESET_B(net51),
    .D(\proj__8.net28 ),
    .Q_N(\proj__8.flop11/notq ),
    .Q(\proj__8.net30 ));
 sg13g2_tiehi \proj__8.flop12/_1__52  (.L_HI(net52));
 sg13g2_dfrbp_1 \proj__8.flop12/_1_  (.CLK(\proj__8.net27 ),
    .RESET_B(net52),
    .D(\proj__8.net31 ),
    .Q_N(\proj__8.net29 ),
    .Q(\proj__8.net32 ));
 sg13g2_tiehi \proj__8.flop13/_1__53  (.L_HI(net53));
 sg13g2_dfrbp_1 \proj__8.flop13/_1_  (.CLK(\proj__8.net30 ),
    .RESET_B(net53),
    .D(\proj__8.net33 ),
    .Q_N(\proj__8.flop13/notq ),
    .Q(\proj__8.net34 ));
 sg13g2_tiehi \proj__8.flop14/_1__54  (.L_HI(net54));
 sg13g2_dfrbp_1 \proj__8.flop14/_1_  (.CLK(\proj__8.net34 ),
    .RESET_B(net54),
    .D(\proj__8.net35 ),
    .Q_N(\proj__8.flop14/notq ),
    .Q(\proj__8.net36 ));
 sg13g2_tiehi \proj__8.flop15/_1__55  (.L_HI(net55));
 sg13g2_dfrbp_1 \proj__8.flop15/_1_  (.CLK(\proj__8.net38 ),
    .RESET_B(net55),
    .D(\proj__8.net37 ),
    .Q_N(\proj__8.flop15/notq ),
    .Q(\proj__8.net39 ));
 sg13g2_tiehi \proj__8.flop16/_1__56  (.L_HI(net56));
 sg13g2_dfrbp_1 \proj__8.flop16/_1_  (.CLK(\proj__8.net36 ),
    .RESET_B(net56),
    .D(\proj__8.net40 ),
    .Q_N(\proj__8.net38 ),
    .Q(\proj__8.net41 ));
 sg13g2_tiehi \proj__8.flop17/_1__57  (.L_HI(net57));
 sg13g2_dfrbp_1 \proj__8.flop17/_1_  (.CLK(\proj__8.net39 ),
    .RESET_B(net57),
    .D(\proj__8.net42 ),
    .Q_N(\proj__8.flop17/notq ),
    .Q(\proj__8.net43 ));
 sg13g2_tiehi \proj__8.flop18/_1__58  (.L_HI(net58));
 sg13g2_dfrbp_1 \proj__8.flop18/_1_  (.CLK(\proj__8.net43 ),
    .RESET_B(net58),
    .D(\proj__8.net44 ),
    .Q_N(\proj__8.flop18/notq ),
    .Q(\proj__8.net45 ));
 sg13g2_tiehi \proj__8.flop19/_1__59  (.L_HI(net59));
 sg13g2_dfrbp_1 \proj__8.flop19/_1_  (.CLK(\proj__8.net47 ),
    .RESET_B(net59),
    .D(\proj__8.net46 ),
    .Q_N(\proj__8.flop19/notq ),
    .Q(\proj__8.net48 ));
 sg13g2_tiehi \proj__8.flop20/_1__60  (.L_HI(net60));
 sg13g2_dfrbp_1 \proj__8.flop20/_1_  (.CLK(\proj__8.net45 ),
    .RESET_B(net60),
    .D(\proj__8.net49 ),
    .Q_N(\proj__8.net47 ),
    .Q(\proj__8.net50 ));
 sg13g2_tiehi \proj__8.flop21/_1__61  (.L_HI(net82));
 sg13g2_dfrbp_1 \proj__8.flop21/_1_  (.CLK(\proj__8.net48 ),
    .RESET_B(net82),
    .D(\proj__8.net51 ),
    .Q_N(\proj__8.flop21/notq ),
    .Q(\proj__8.net52 ));
 sg13g2_tiehi \proj__8.flop22/_1__62  (.L_HI(net83));
 sg13g2_dfrbp_1 \proj__8.flop22/_1_  (.CLK(\proj__8.net52 ),
    .RESET_B(net83),
    .D(\proj__8.net53 ),
    .Q_N(\proj__8.flop22/notq ),
    .Q(\proj__8.net54 ));
 sg13g2_tiehi \proj__8.flop23/_1__63  (.L_HI(net84));
 sg13g2_dfrbp_1 \proj__8.flop23/_1_  (.CLK(\proj__8.net56 ),
    .RESET_B(net84),
    .D(\proj__8.net55 ),
    .Q_N(\proj__8.flop23/notq ),
    .Q(\proj__8.net57 ));
 sg13g2_tiehi \proj__8.flop24/_1__64  (.L_HI(net85));
 sg13g2_dfrbp_1 \proj__8.flop24/_1_  (.CLK(\proj__8.net54 ),
    .RESET_B(net85),
    .D(\proj__8.net58 ),
    .Q_N(\proj__8.net56 ),
    .Q(\proj__8.net59 ));
 sg13g2_tiehi \proj__8.flop25/_1__65  (.L_HI(net86));
 sg13g2_dfrbp_1 \proj__8.flop25/_1_  (.CLK(\proj__8.net57 ),
    .RESET_B(net86),
    .D(\proj__8.net60 ),
    .Q_N(\proj__8.flop25/notq ),
    .Q(\proj__8.net61 ));
 sg13g2_tiehi \proj__8.flop26/_1__66  (.L_HI(net87));
 sg13g2_dfrbp_1 \proj__8.flop26/_1_  (.CLK(\proj__8.net61 ),
    .RESET_B(net87),
    .D(\proj__8.net62 ),
    .Q_N(\proj__8.flop26/notq ),
    .Q(\proj__8.net63 ));
 sg13g2_tiehi \proj__8.flop27/_1__67  (.L_HI(net88));
 sg13g2_dfrbp_1 \proj__8.flop27/_1_  (.CLK(\proj__8.net65 ),
    .RESET_B(net88),
    .D(\proj__8.net64 ),
    .Q_N(\proj__8.flop27/notq ),
    .Q(\proj__8.net66 ));
 sg13g2_tiehi \proj__8.flop28/_1__68  (.L_HI(net89));
 sg13g2_dfrbp_1 \proj__8.flop28/_1_  (.CLK(\proj__8.net63 ),
    .RESET_B(net89),
    .D(\proj__8.net67 ),
    .Q_N(\proj__8.net65 ),
    .Q(\proj__8.net68 ));
 sg13g2_tiehi \proj__8.flop29/_1__69  (.L_HI(net90));
 sg13g2_dfrbp_1 \proj__8.flop29/_1_  (.CLK(\proj__8.net66 ),
    .RESET_B(net90),
    .D(\proj__8.net69 ),
    .Q_N(\proj__8.flop29/notq ),
    .Q(\proj__8.net70 ));
 sg13g2_tiehi \proj__8.flop30/_1__70  (.L_HI(net91));
 sg13g2_dfrbp_1 \proj__8.flop30/_1_  (.CLK(\proj__8.net70 ),
    .RESET_B(net91),
    .D(\proj__8.net71 ),
    .Q_N(\proj__8.flop30/notq ),
    .Q(\proj__8.net72 ));
 sg13g2_tiehi \proj__8.flop31/_1__71  (.L_HI(net92));
 sg13g2_dfrbp_1 \proj__8.flop31/_1_  (.CLK(\proj__8.net74 ),
    .RESET_B(net92),
    .D(\proj__8.net73 ),
    .Q_N(\proj__8.flop31/notq ),
    .Q(\proj__8.net75 ));
 sg13g2_tiehi \proj__8.flop32/_1__72  (.L_HI(net93));
 sg13g2_dfrbp_1 \proj__8.flop32/_1_  (.CLK(\proj__8.net72 ),
    .RESET_B(net93),
    .D(\proj__8.net76 ),
    .Q_N(\proj__8.net74 ),
    .Q(\proj__8.net77 ));
 sg13g2_tiehi \proj__8.flop33/_1__73  (.L_HI(net94));
 sg13g2_dfrbp_1 \proj__8.flop33/_1_  (.CLK(\proj__8.net75 ),
    .RESET_B(net94),
    .D(\proj__8.net78 ),
    .Q_N(\proj__8.flop33/notq ),
    .Q(\proj__8.net79 ));
 sg13g2_tiehi \proj__8.flop34/_1__74  (.L_HI(net95));
 sg13g2_dfrbp_1 \proj__8.flop34/_1_  (.CLK(\proj__8.net79 ),
    .RESET_B(net95),
    .D(\proj__8.net80 ),
    .Q_N(\proj__8.flop34/notq ),
    .Q(\proj__8.net81 ));
 sg13g2_tiehi \proj__8.flop35/_1__75  (.L_HI(net96));
 sg13g2_dfrbp_1 \proj__8.flop35/_1_  (.CLK(\proj__8.net83 ),
    .RESET_B(net96),
    .D(\proj__8.net82 ),
    .Q_N(\proj__8.flop35/notq ),
    .Q(\proj__8.net84 ));
 sg13g2_tiehi \proj__8.flop36/_1__76  (.L_HI(net97));
 sg13g2_dfrbp_1 \proj__8.flop36/_1_  (.CLK(\proj__8.net81 ),
    .RESET_B(net97),
    .D(\proj__8.net85 ),
    .Q_N(\proj__8.net83 ),
    .Q(\proj__8.net86 ));
 sg13g2_tiehi \proj__8.flop37/_1__77  (.L_HI(net98));
 sg13g2_dfrbp_1 \proj__8.flop37/_1_  (.CLK(\proj__8.net84 ),
    .RESET_B(net98),
    .D(\proj__8.net87 ),
    .Q_N(\proj__8.flop37/notq ),
    .Q(\proj__8.net88 ));
 sg13g2_tiehi \proj__8.flop38/_1__78  (.L_HI(net99));
 sg13g2_dfrbp_1 \proj__8.flop38/_1_  (.CLK(\proj__8.net88 ),
    .RESET_B(net99),
    .D(\proj__8.net89 ),
    .Q_N(\proj__8.flop38/notq ),
    .Q(\proj__8.net90 ));
 sg13g2_tiehi \proj__8.flop39/_1__79  (.L_HI(net100));
 sg13g2_dfrbp_1 \proj__8.flop39/_1_  (.CLK(\proj__8.net92 ),
    .RESET_B(net100),
    .D(\proj__8.net91 ),
    .Q_N(\proj__8.flop39/notq ),
    .Q(\proj__8.net93 ));
 sg13g2_tiehi \proj__8.flop40/_1__80  (.L_HI(net101));
 sg13g2_dfrbp_1 \proj__8.flop40/_1_  (.CLK(\proj__8.net90 ),
    .RESET_B(net101),
    .D(\proj__8.net94 ),
    .Q_N(\proj__8.net92 ),
    .Q(\proj__8.net95 ));
 sg13g2_tiehi \proj__8.flop41/_1__81  (.L_HI(net102));
 sg13g2_dfrbp_1 \proj__8.flop41/_1_  (.CLK(\proj__8.net93 ),
    .RESET_B(net102),
    .D(\proj__8.net96 ),
    .Q_N(\proj__8.flop41/notq ),
    .Q(\proj__8.net10 ));
 sg13g2_tiehi \proj__8.flop6/_1__82  (.L_HI(net103));
 sg13g2_dfrbp_1 \proj__8.flop6/_1_  (.CLK(clknet_1_0__leaf_clk_regs),
    .RESET_B(net103),
    .D(\proj__8.net17 ),
    .Q_N(\proj__8.flop6/notq ),
    .Q(\proj__8.net18 ));
 sg13g2_tiehi \proj__8.flop7/_1__83  (.L_HI(net104));
 sg13g2_dfrbp_1 \proj__8.flop7/_1_  (.CLK(\proj__8.net20 ),
    .RESET_B(net104),
    .D(\proj__8.net19 ),
    .Q_N(\proj__8.flop7/notq ),
    .Q(\proj__8.net21 ));
 sg13g2_tiehi \proj__8.flop8/_1__84  (.L_HI(net105));
 sg13g2_dfrbp_1 \proj__8.flop8/_1_  (.CLK(\proj__8.net18 ),
    .RESET_B(net105),
    .D(\proj__8.net22 ),
    .Q_N(\proj__8.net20 ),
    .Q(\proj__8.net23 ));
 sg13g2_tiehi \proj__8.flop9/_1__85  (.L_HI(net106));
 sg13g2_dfrbp_1 \proj__8.flop9/_1_  (.CLK(\proj__8.net21 ),
    .RESET_B(net106),
    .D(\proj__8.net24 ),
    .Q_N(\proj__8.flop9/notq ),
    .Q(\proj__8.net25 ));
 sg13g2_inv_1 \proj__4.not1/_0__1  (.Y(net107),
    .A(clknet_1_1__leaf_clk));
 sg13g2_inv_1 \proj__8.not1/_0_  (.Y(\proj__8.net17 ),
    .A(net109));
 sg13g2_inv_1 \proj__8.not10/_0_  (.Y(\proj__8.net40 ),
    .A(\proj__8.net41 ));
 sg13g2_inv_1 \proj__8.not100/_0_  (.Y(\proj__8.net160 ),
    .A(\proj__8.net159 ));
 sg13g2_inv_1 \proj__8.not101/_0_  (.Y(\proj__8.net154 ),
    .A(\proj__8.net160 ));
 sg13g2_inv_1 \proj__8.not102/_0_  (.Y(\proj__8.net162 ),
    .A(\proj__8.net161 ));
 sg13g2_inv_1 \proj__8.not103/_0_  (.Y(\proj__8.net163 ),
    .A(\proj__8.net162 ));
 sg13g2_inv_1 \proj__8.not104/_0_  (.Y(\proj__8.net164 ),
    .A(\proj__8.net163 ));
 sg13g2_inv_1 \proj__8.not105/_0_  (.Y(\proj__8.net165 ),
    .A(\proj__8.net164 ));
 sg13g2_inv_1 \proj__8.not106/_0_  (.Y(\proj__8.net167 ),
    .A(\proj__8.net166 ));
 sg13g2_inv_1 \proj__8.not107/_0_  (.Y(\proj__8.net168 ),
    .A(\proj__8.net167 ));
 sg13g2_inv_1 \proj__8.not108/_0_  (.Y(\proj__8.net169 ),
    .A(\proj__8.net168 ));
 sg13g2_inv_1 \proj__8.not109/_0_  (.Y(\proj__8.net161 ),
    .A(\proj__8.net169 ));
 sg13g2_inv_1 \proj__8.not11/_0_  (.Y(\proj__8.net37 ),
    .A(\proj__8.net39 ));
 sg13g2_inv_1 \proj__8.not110/_0_  (.Y(\proj__8.net171 ),
    .A(\proj__8.net170 ));
 sg13g2_inv_1 \proj__8.not111/_0_  (.Y(\proj__8.net172 ),
    .A(\proj__8.net171 ));
 sg13g2_inv_1 \proj__8.not112/_0_  (.Y(\proj__8.net173 ),
    .A(\proj__8.net172 ));
 sg13g2_inv_1 \proj__8.not113/_0_  (.Y(\proj__8.net174 ),
    .A(\proj__8.net173 ));
 sg13g2_inv_1 \proj__8.not114/_0_  (.Y(\proj__8.net175 ),
    .A(\proj__8.net165 ));
 sg13g2_inv_1 \proj__8.not115/_0_  (.Y(\proj__8.net176 ),
    .A(\proj__8.net175 ));
 sg13g2_inv_1 \proj__8.not116/_0_  (.Y(\proj__8.net177 ),
    .A(\proj__8.net176 ));
 sg13g2_inv_1 \proj__8.not117/_0_  (.Y(\proj__8.net170 ),
    .A(\proj__8.net177 ));
 sg13g2_inv_1 \proj__8.not118/_0_  (.Y(\proj__8.net179 ),
    .A(\proj__8.net178 ));
 sg13g2_inv_1 \proj__8.not119/_0_  (.Y(\proj__8.net180 ),
    .A(\proj__8.net179 ));
 sg13g2_inv_1 \proj__8.not12/_0_  (.Y(\proj__8.net42 ),
    .A(\proj__8.net43 ));
 sg13g2_inv_1 \proj__8.not120/_0_  (.Y(\proj__8.net181 ),
    .A(\proj__8.net180 ));
 sg13g2_inv_1 \proj__8.not121/_0_  (.Y(\proj__8.net182 ),
    .A(\proj__8.net181 ));
 sg13g2_inv_1 \proj__8.not122/_0_  (.Y(\proj__8.net183 ),
    .A(\proj__8.net174 ));
 sg13g2_inv_1 \proj__8.not123/_0_  (.Y(\proj__8.net184 ),
    .A(\proj__8.net183 ));
 sg13g2_inv_1 \proj__8.not124/_0_  (.Y(\proj__8.net185 ),
    .A(\proj__8.net184 ));
 sg13g2_inv_1 \proj__8.not125/_0_  (.Y(\proj__8.net178 ),
    .A(\proj__8.net185 ));
 sg13g2_inv_1 \proj__8.not126/_0_  (.Y(\proj__8.net187 ),
    .A(\proj__8.net186 ));
 sg13g2_inv_1 \proj__8.not127/_0_  (.Y(\proj__8.net188 ),
    .A(\proj__8.net187 ));
 sg13g2_inv_1 \proj__8.not128/_0_  (.Y(\proj__8.net189 ),
    .A(\proj__8.net188 ));
 sg13g2_inv_1 \proj__8.not129/_0_  (.Y(\proj__8.net190 ),
    .A(\proj__8.net189 ));
 sg13g2_inv_1 \proj__8.not13/_0_  (.Y(\proj__8.net44 ),
    .A(\proj__8.net45 ));
 sg13g2_inv_1 \proj__8.not130/_0_  (.Y(\proj__8.net191 ),
    .A(\proj__8.net182 ));
 sg13g2_inv_1 \proj__8.not131/_0_  (.Y(\proj__8.net192 ),
    .A(\proj__8.net191 ));
 sg13g2_inv_1 \proj__8.not132/_0_  (.Y(\proj__8.net193 ),
    .A(\proj__8.net192 ));
 sg13g2_inv_1 \proj__8.not133/_0_  (.Y(\proj__8.net186 ),
    .A(\proj__8.net193 ));
 sg13g2_inv_1 \proj__8.not134/_0_  (.Y(\proj__8.net195 ),
    .A(\proj__8.net194 ));
 sg13g2_inv_1 \proj__8.not135/_0_  (.Y(\proj__8.net196 ),
    .A(\proj__8.net195 ));
 sg13g2_inv_1 \proj__8.not136/_0_  (.Y(\proj__8.net197 ),
    .A(\proj__8.net196 ));
 sg13g2_inv_1 \proj__8.not137/_0_  (.Y(\proj__8.net198 ),
    .A(\proj__8.net197 ));
 sg13g2_inv_1 \proj__8.not138/_0_  (.Y(\proj__8.net199 ),
    .A(\proj__8.net126 ));
 sg13g2_inv_1 \proj__8.not139/_0_  (.Y(\proj__8.net200 ),
    .A(\proj__8.net199 ));
 sg13g2_inv_1 \proj__8.not14/_0_  (.Y(\proj__8.net49 ),
    .A(\proj__8.net50 ));
 sg13g2_inv_1 \proj__8.not140/_0_  (.Y(\proj__8.net201 ),
    .A(\proj__8.net200 ));
 sg13g2_inv_1 \proj__8.not141/_0_  (.Y(\proj__8.net194 ),
    .A(\proj__8.net201 ));
 sg13g2_inv_1 \proj__8.not142/_0_  (.Y(\proj__8.net203 ),
    .A(\proj__8.net202 ));
 sg13g2_inv_1 \proj__8.not143/_0_  (.Y(\proj__8.net204 ),
    .A(\proj__8.net203 ));
 sg13g2_inv_1 \proj__8.not144/_0_  (.Y(\proj__8.net205 ),
    .A(\proj__8.net204 ));
 sg13g2_inv_1 \proj__8.not145/_0_  (.Y(\proj__8.net206 ),
    .A(\proj__8.net205 ));
 sg13g2_inv_1 \proj__8.not146/_0_  (.Y(\proj__8.net207 ),
    .A(\proj__8.net198 ));
 sg13g2_inv_1 \proj__8.not147/_0_  (.Y(\proj__8.net208 ),
    .A(\proj__8.net207 ));
 sg13g2_inv_1 \proj__8.not148/_0_  (.Y(\proj__8.net209 ),
    .A(\proj__8.net208 ));
 sg13g2_inv_1 \proj__8.not149/_0_  (.Y(\proj__8.net202 ),
    .A(\proj__8.net209 ));
 sg13g2_inv_1 \proj__8.not15/_0_  (.Y(\proj__8.net46 ),
    .A(\proj__8.net48 ));
 sg13g2_inv_1 \proj__8.not150/_0_  (.Y(\proj__8.net211 ),
    .A(\proj__8.net210 ));
 sg13g2_inv_1 \proj__8.not151/_0_  (.Y(\proj__8.net212 ),
    .A(\proj__8.net211 ));
 sg13g2_inv_1 \proj__8.not152/_0_  (.Y(\proj__8.net213 ),
    .A(\proj__8.net212 ));
 sg13g2_inv_1 \proj__8.not153/_0_  (.Y(\proj__8.net214 ),
    .A(\proj__8.net213 ));
 sg13g2_inv_1 \proj__8.not154/_0_  (.Y(\proj__8.net215 ),
    .A(\proj__8.net206 ));
 sg13g2_inv_1 \proj__8.not155/_0_  (.Y(\proj__8.net216 ),
    .A(\proj__8.net215 ));
 sg13g2_inv_1 \proj__8.not156/_0_  (.Y(\proj__8.net217 ),
    .A(\proj__8.net216 ));
 sg13g2_inv_1 \proj__8.not157/_0_  (.Y(\proj__8.net210 ),
    .A(\proj__8.net217 ));
 sg13g2_inv_1 \proj__8.not158/_0_  (.Y(\proj__8.net219 ),
    .A(\proj__8.net218 ));
 sg13g2_inv_1 \proj__8.not159/_0_  (.Y(\proj__8.net220 ),
    .A(\proj__8.net219 ));
 sg13g2_inv_1 \proj__8.not16/_0_  (.Y(\proj__8.net51 ),
    .A(\proj__8.net52 ));
 sg13g2_inv_1 \proj__8.not160/_0_  (.Y(\proj__8.net221 ),
    .A(\proj__8.net220 ));
 sg13g2_inv_1 \proj__8.not161/_0_  (.Y(\proj__8.net166 ),
    .A(\proj__8.net221 ));
 sg13g2_inv_1 \proj__8.not162/_0_  (.Y(\proj__8.net222 ),
    .A(\proj__8.net214 ));
 sg13g2_inv_1 \proj__8.not163/_0_  (.Y(\proj__8.net223 ),
    .A(\proj__8.net222 ));
 sg13g2_inv_1 \proj__8.not164/_0_  (.Y(\proj__8.net224 ),
    .A(\proj__8.net223 ));
 sg13g2_inv_1 \proj__8.not165/_0_  (.Y(\proj__8.net218 ),
    .A(\proj__8.net224 ));
 sg13g2_inv_1 \proj__8.not166/_0_  (.Y(\proj__8.net226 ),
    .A(\proj__8.net225 ));
 sg13g2_inv_1 \proj__8.not167/_0_  (.Y(\proj__8.net227 ),
    .A(\proj__8.net226 ));
 sg13g2_inv_1 \proj__8.not168/_0_  (.Y(\proj__8.net228 ),
    .A(\proj__8.net227 ));
 sg13g2_inv_1 \proj__8.not169/_0_  (.Y(\proj__8.net229 ),
    .A(\proj__8.net228 ));
 sg13g2_inv_1 \proj__8.not17/_0_  (.Y(\proj__8.net53 ),
    .A(\proj__8.net54 ));
 sg13g2_inv_1 \proj__8.not170/_0_  (.Y(\proj__8.net231 ),
    .A(\proj__8.net230 ));
 sg13g2_inv_1 \proj__8.not171/_0_  (.Y(\proj__8.net232 ),
    .A(\proj__8.net231 ));
 sg13g2_inv_1 \proj__8.not172/_0_  (.Y(\proj__8.net233 ),
    .A(\proj__8.net232 ));
 sg13g2_inv_1 \proj__8.not173/_0_  (.Y(\proj__8.net225 ),
    .A(\proj__8.net233 ));
 sg13g2_inv_1 \proj__8.not174/_0_  (.Y(\proj__8.net235 ),
    .A(\proj__8.net234 ));
 sg13g2_inv_1 \proj__8.not175/_0_  (.Y(\proj__8.net236 ),
    .A(\proj__8.net235 ));
 sg13g2_inv_1 \proj__8.not176/_0_  (.Y(\proj__8.net237 ),
    .A(\proj__8.net236 ));
 sg13g2_inv_1 \proj__8.not177/_0_  (.Y(\proj__8.net238 ),
    .A(\proj__8.net237 ));
 sg13g2_inv_1 \proj__8.not178/_0_  (.Y(\proj__8.net239 ),
    .A(\proj__8.net229 ));
 sg13g2_inv_1 \proj__8.not179/_0_  (.Y(\proj__8.net240 ),
    .A(\proj__8.net239 ));
 sg13g2_inv_1 \proj__8.not18/_0_  (.Y(\proj__8.net58 ),
    .A(\proj__8.net59 ));
 sg13g2_inv_1 \proj__8.not180/_0_  (.Y(\proj__8.net241 ),
    .A(\proj__8.net240 ));
 sg13g2_inv_1 \proj__8.not181/_0_  (.Y(\proj__8.net234 ),
    .A(\proj__8.net241 ));
 sg13g2_inv_1 \proj__8.not182/_0_  (.Y(\proj__8.net243 ),
    .A(\proj__8.net242 ));
 sg13g2_inv_1 \proj__8.not183/_0_  (.Y(\proj__8.net244 ),
    .A(\proj__8.net243 ));
 sg13g2_inv_1 \proj__8.not184/_0_  (.Y(\proj__8.net245 ),
    .A(\proj__8.net244 ));
 sg13g2_inv_1 \proj__8.not185/_0_  (.Y(\proj__8.net246 ),
    .A(\proj__8.net245 ));
 sg13g2_inv_1 \proj__8.not186/_0_  (.Y(\proj__8.net247 ),
    .A(\proj__8.net238 ));
 sg13g2_inv_1 \proj__8.not187/_0_  (.Y(\proj__8.net248 ),
    .A(\proj__8.net247 ));
 sg13g2_inv_1 \proj__8.not188/_0_  (.Y(\proj__8.net249 ),
    .A(\proj__8.net248 ));
 sg13g2_inv_1 \proj__8.not189/_0_  (.Y(\proj__8.net242 ),
    .A(\proj__8.net249 ));
 sg13g2_inv_1 \proj__8.not19/_0_  (.Y(\proj__8.net55 ),
    .A(\proj__8.net57 ));
 sg13g2_inv_1 \proj__8.not190/_0_  (.Y(\proj__8.net251 ),
    .A(\proj__8.net250 ));
 sg13g2_inv_1 \proj__8.not191/_0_  (.Y(\proj__8.net252 ),
    .A(\proj__8.net251 ));
 sg13g2_inv_1 \proj__8.not192/_0_  (.Y(\proj__8.net253 ),
    .A(\proj__8.net252 ));
 sg13g2_inv_1 \proj__8.not193/_0_  (.Y(\proj__8.net254 ),
    .A(\proj__8.net253 ));
 sg13g2_inv_1 \proj__8.not194/_0_  (.Y(\proj__8.net255 ),
    .A(\proj__8.net246 ));
 sg13g2_inv_1 \proj__8.not195/_0_  (.Y(\proj__8.net256 ),
    .A(\proj__8.net255 ));
 sg13g2_inv_1 \proj__8.not196/_0_  (.Y(\proj__8.net257 ),
    .A(\proj__8.net256 ));
 sg13g2_inv_1 \proj__8.not197/_0_  (.Y(\proj__8.net250 ),
    .A(\proj__8.net257 ));
 sg13g2_inv_1 \proj__8.not198/_0_  (.Y(\proj__8.net259 ),
    .A(\proj__8.net258 ));
 sg13g2_inv_1 \proj__8.not199/_0_  (.Y(\proj__8.net260 ),
    .A(\proj__8.net259 ));
 sg13g2_inv_1 \proj__8.not2/_0_  (.Y(\proj__8.net22 ),
    .A(\proj__8.net23 ));
 sg13g2_inv_1 \proj__8.not20/_0_  (.Y(\proj__8.net60 ),
    .A(\proj__8.net61 ));
 sg13g2_inv_1 \proj__8.not200/_0_  (.Y(\proj__8.net261 ),
    .A(\proj__8.net260 ));
 sg13g2_inv_1 \proj__8.not201/_0_  (.Y(\proj__8.net262 ),
    .A(\proj__8.net261 ));
 sg13g2_inv_1 \proj__8.not202/_0_  (.Y(\proj__8.net263 ),
    .A(\proj__8.net190 ));
 sg13g2_inv_1 \proj__8.not203/_0_  (.Y(\proj__8.net264 ),
    .A(\proj__8.net263 ));
 sg13g2_inv_1 \proj__8.not204/_0_  (.Y(\proj__8.net265 ),
    .A(\proj__8.net264 ));
 sg13g2_inv_1 \proj__8.not205/_0_  (.Y(\proj__8.net258 ),
    .A(\proj__8.net265 ));
 sg13g2_inv_1 \proj__8.not206/_0_  (.Y(\proj__8.net267 ),
    .A(\proj__8.net266 ));
 sg13g2_inv_1 \proj__8.not207/_0_  (.Y(\proj__8.net268 ),
    .A(\proj__8.net267 ));
 sg13g2_inv_1 \proj__8.not208/_0_  (.Y(\proj__8.net269 ),
    .A(\proj__8.net268 ));
 sg13g2_inv_1 \proj__8.not209/_0_  (.Y(\proj__8.net270 ),
    .A(\proj__8.net269 ));
 sg13g2_inv_1 \proj__8.not21/_0_  (.Y(\proj__8.net62 ),
    .A(\proj__8.net63 ));
 sg13g2_inv_1 \proj__8.not210/_0_  (.Y(\proj__8.net271 ),
    .A(\proj__8.net262 ));
 sg13g2_inv_1 \proj__8.not211/_0_  (.Y(\proj__8.net272 ),
    .A(\proj__8.net271 ));
 sg13g2_inv_1 \proj__8.not212/_0_  (.Y(\proj__8.net273 ),
    .A(\proj__8.net272 ));
 sg13g2_inv_1 \proj__8.not213/_0_  (.Y(\proj__8.net266 ),
    .A(\proj__8.net273 ));
 sg13g2_inv_1 \proj__8.not214/_0_  (.Y(\proj__8.net275 ),
    .A(\proj__8.net274 ));
 sg13g2_inv_1 \proj__8.not215/_0_  (.Y(\proj__8.net276 ),
    .A(\proj__8.net275 ));
 sg13g2_inv_1 \proj__8.not216/_0_  (.Y(\proj__8.net277 ),
    .A(\proj__8.net276 ));
 sg13g2_inv_1 \proj__8.not217/_0_  (.Y(\proj__8.net278 ),
    .A(\proj__8.net277 ));
 sg13g2_inv_1 \proj__8.not218/_0_  (.Y(\proj__8.net279 ),
    .A(\proj__8.net270 ));
 sg13g2_inv_1 \proj__8.not219/_0_  (.Y(\proj__8.net280 ),
    .A(\proj__8.net279 ));
 sg13g2_inv_1 \proj__8.not22/_0_  (.Y(\proj__8.net67 ),
    .A(\proj__8.net68 ));
 sg13g2_inv_1 \proj__8.not220/_0_  (.Y(\proj__8.net281 ),
    .A(\proj__8.net280 ));
 sg13g2_inv_1 \proj__8.not221/_0_  (.Y(\proj__8.net274 ),
    .A(\proj__8.net281 ));
 sg13g2_inv_1 \proj__8.not222/_0_  (.Y(\proj__8.net283 ),
    .A(\proj__8.net282 ));
 sg13g2_inv_1 \proj__8.not223/_0_  (.Y(\proj__8.net284 ),
    .A(\proj__8.net283 ));
 sg13g2_inv_1 \proj__8.not224/_0_  (.Y(\proj__8.net285 ),
    .A(\proj__8.net284 ));
 sg13g2_inv_1 \proj__8.not225/_0_  (.Y(\proj__8.net230 ),
    .A(\proj__8.net285 ));
 sg13g2_inv_1 \proj__8.not226/_0_  (.Y(\proj__8.net286 ),
    .A(\proj__8.net278 ));
 sg13g2_inv_1 \proj__8.not227/_0_  (.Y(\proj__8.net287 ),
    .A(\proj__8.net286 ));
 sg13g2_inv_1 \proj__8.not228/_0_  (.Y(\proj__8.net288 ),
    .A(\proj__8.net287 ));
 sg13g2_inv_1 \proj__8.not229/_0_  (.Y(\proj__8.net282 ),
    .A(\proj__8.net288 ));
 sg13g2_inv_1 \proj__8.not23/_0_  (.Y(\proj__8.net64 ),
    .A(\proj__8.net66 ));
 sg13g2_inv_1 \proj__8.not230/_0_  (.Y(\proj__8.net290 ),
    .A(\proj__8.net289 ));
 sg13g2_inv_1 \proj__8.not231/_0_  (.Y(\proj__8.net291 ),
    .A(\proj__8.net290 ));
 sg13g2_inv_1 \proj__8.not232/_0_  (.Y(\proj__8.net292 ),
    .A(\proj__8.net291 ));
 sg13g2_inv_1 \proj__8.not233/_0_  (.Y(\proj__8.net293 ),
    .A(\proj__8.net292 ));
 sg13g2_inv_1 \proj__8.not234/_0_  (.Y(\proj__8.net295 ),
    .A(\proj__8.net294 ));
 sg13g2_inv_1 \proj__8.not235/_0_  (.Y(\proj__8.net296 ),
    .A(\proj__8.net295 ));
 sg13g2_inv_1 \proj__8.not236/_0_  (.Y(\proj__8.net297 ),
    .A(\proj__8.net296 ));
 sg13g2_inv_1 \proj__8.not237/_0_  (.Y(\proj__8.net289 ),
    .A(\proj__8.net297 ));
 sg13g2_inv_1 \proj__8.not238/_0_  (.Y(\proj__8.net299 ),
    .A(\proj__8.net298 ));
 sg13g2_inv_1 \proj__8.not239/_0_  (.Y(\proj__8.net300 ),
    .A(\proj__8.net299 ));
 sg13g2_inv_1 \proj__8.not24/_0_  (.Y(\proj__8.net69 ),
    .A(\proj__8.net70 ));
 sg13g2_inv_1 \proj__8.not240/_0_  (.Y(\proj__8.net301 ),
    .A(\proj__8.net300 ));
 sg13g2_inv_1 \proj__8.not241/_0_  (.Y(\proj__8.net302 ),
    .A(\proj__8.net301 ));
 sg13g2_inv_1 \proj__8.not242/_0_  (.Y(\proj__8.net303 ),
    .A(\proj__8.net293 ));
 sg13g2_inv_1 \proj__8.not243/_0_  (.Y(\proj__8.net304 ),
    .A(\proj__8.net303 ));
 sg13g2_inv_1 \proj__8.not244/_0_  (.Y(\proj__8.net305 ),
    .A(\proj__8.net304 ));
 sg13g2_inv_1 \proj__8.not245/_0_  (.Y(\proj__8.net298 ),
    .A(\proj__8.net305 ));
 sg13g2_inv_1 \proj__8.not246/_0_  (.Y(\proj__8.net307 ),
    .A(\proj__8.net306 ));
 sg13g2_inv_1 \proj__8.not247/_0_  (.Y(\proj__8.net308 ),
    .A(\proj__8.net307 ));
 sg13g2_inv_1 \proj__8.not248/_0_  (.Y(\proj__8.net309 ),
    .A(\proj__8.net308 ));
 sg13g2_inv_1 \proj__8.not249/_0_  (.Y(\proj__8.net310 ),
    .A(\proj__8.net309 ));
 sg13g2_inv_1 \proj__8.not25/_0_  (.Y(\proj__8.net71 ),
    .A(\proj__8.net72 ));
 sg13g2_inv_1 \proj__8.not250/_0_  (.Y(\proj__8.net311 ),
    .A(\proj__8.net302 ));
 sg13g2_inv_1 \proj__8.not251/_0_  (.Y(\proj__8.net312 ),
    .A(\proj__8.net311 ));
 sg13g2_inv_1 \proj__8.not252/_0_  (.Y(\proj__8.net313 ),
    .A(\proj__8.net312 ));
 sg13g2_inv_1 \proj__8.not253/_0_  (.Y(\proj__8.net306 ),
    .A(\proj__8.net313 ));
 sg13g2_inv_1 \proj__8.not254/_0_  (.Y(\proj__8.net315 ),
    .A(\proj__8.net314 ));
 sg13g2_inv_1 \proj__8.not255/_0_  (.Y(\proj__8.net316 ),
    .A(\proj__8.net315 ));
 sg13g2_inv_1 \proj__8.not256/_0_  (.Y(\proj__8.net317 ),
    .A(\proj__8.net316 ));
 sg13g2_inv_1 \proj__8.not257/_0_  (.Y(\proj__8.net318 ),
    .A(\proj__8.net317 ));
 sg13g2_inv_1 \proj__8.not258/_0_  (.Y(\proj__8.net319 ),
    .A(\proj__8.net310 ));
 sg13g2_inv_1 \proj__8.not259/_0_  (.Y(\proj__8.net320 ),
    .A(\proj__8.net319 ));
 sg13g2_inv_1 \proj__8.not26/_0_  (.Y(\proj__8.net76 ),
    .A(\proj__8.net77 ));
 sg13g2_inv_1 \proj__8.not260/_0_  (.Y(\proj__8.net321 ),
    .A(\proj__8.net320 ));
 sg13g2_inv_1 \proj__8.not261/_0_  (.Y(\proj__8.net314 ),
    .A(\proj__8.net321 ));
 sg13g2_inv_1 \proj__8.not262/_0_  (.Y(\proj__8.net323 ),
    .A(\proj__8.net322 ));
 sg13g2_inv_1 \proj__8.not263/_0_  (.Y(\proj__8.net324 ),
    .A(\proj__8.net323 ));
 sg13g2_inv_1 \proj__8.not264/_0_  (.Y(\proj__8.net325 ),
    .A(\proj__8.net324 ));
 sg13g2_inv_1 \proj__8.not265/_0_  (.Y(\proj__8.net326 ),
    .A(\proj__8.net325 ));
 sg13g2_inv_1 \proj__8.not266/_0_  (.Y(\proj__8.net327 ),
    .A(\proj__8.net254 ));
 sg13g2_inv_1 \proj__8.not267/_0_  (.Y(\proj__8.net328 ),
    .A(\proj__8.net327 ));
 sg13g2_inv_1 \proj__8.not268/_0_  (.Y(\proj__8.net329 ),
    .A(\proj__8.net328 ));
 sg13g2_inv_1 \proj__8.not269/_0_  (.Y(\proj__8.net322 ),
    .A(\proj__8.net329 ));
 sg13g2_inv_1 \proj__8.not27/_0_  (.Y(\proj__8.net73 ),
    .A(\proj__8.net75 ));
 sg13g2_inv_1 \proj__8.not270/_0_  (.Y(\proj__8.net331 ),
    .A(\proj__8.net330 ));
 sg13g2_inv_1 \proj__8.not271/_0_  (.Y(\proj__8.net332 ),
    .A(\proj__8.net331 ));
 sg13g2_inv_1 \proj__8.not272/_0_  (.Y(\proj__8.net333 ),
    .A(\proj__8.net332 ));
 sg13g2_inv_1 \proj__8.not273/_0_  (.Y(\proj__8.net334 ),
    .A(\proj__8.net333 ));
 sg13g2_inv_1 \proj__8.not274/_0_  (.Y(\proj__8.net335 ),
    .A(\proj__8.net326 ));
 sg13g2_inv_1 \proj__8.not275/_0_  (.Y(\proj__8.net336 ),
    .A(\proj__8.net335 ));
 sg13g2_inv_1 \proj__8.not276/_0_  (.Y(\proj__8.net337 ),
    .A(\proj__8.net336 ));
 sg13g2_inv_1 \proj__8.not277/_0_  (.Y(\proj__8.net330 ),
    .A(\proj__8.net337 ));
 sg13g2_inv_1 \proj__8.not278/_0_  (.Y(\proj__8.net339 ),
    .A(\proj__8.net338 ));
 sg13g2_inv_1 \proj__8.not279/_0_  (.Y(\proj__8.net340 ),
    .A(\proj__8.net339 ));
 sg13g2_inv_1 \proj__8.not28/_0_  (.Y(\proj__8.net78 ),
    .A(\proj__8.net79 ));
 sg13g2_inv_1 \proj__8.not280/_0_  (.Y(\proj__8.net341 ),
    .A(\proj__8.net340 ));
 sg13g2_inv_1 \proj__8.not281/_0_  (.Y(\proj__8.net342 ),
    .A(\proj__8.net341 ));
 sg13g2_inv_1 \proj__8.not282/_0_  (.Y(\proj__8.net343 ),
    .A(\proj__8.net334 ));
 sg13g2_inv_1 \proj__8.not283/_0_  (.Y(\proj__8.net344 ),
    .A(\proj__8.net343 ));
 sg13g2_inv_1 \proj__8.not284/_0_  (.Y(\proj__8.net345 ),
    .A(\proj__8.net344 ));
 sg13g2_inv_1 \proj__8.not285/_0_  (.Y(\proj__8.net338 ),
    .A(\proj__8.net345 ));
 sg13g2_inv_1 \proj__8.not286/_0_  (.Y(\proj__8.net347 ),
    .A(\proj__8.net346 ));
 sg13g2_inv_1 \proj__8.not287/_0_  (.Y(\proj__8.net348 ),
    .A(\proj__8.net347 ));
 sg13g2_inv_1 \proj__8.not288/_0_  (.Y(\proj__8.net349 ),
    .A(\proj__8.net348 ));
 sg13g2_inv_1 \proj__8.not289/_0_  (.Y(\proj__8.net294 ),
    .A(\proj__8.net349 ));
 sg13g2_inv_1 \proj__8.not29/_0_  (.Y(\proj__8.net80 ),
    .A(\proj__8.net81 ));
 sg13g2_inv_1 \proj__8.not290/_0_  (.Y(\proj__8.net350 ),
    .A(\proj__8.net342 ));
 sg13g2_inv_1 \proj__8.not291/_0_  (.Y(\proj__8.net351 ),
    .A(\proj__8.net350 ));
 sg13g2_inv_1 \proj__8.not292/_0_  (.Y(\proj__8.net352 ),
    .A(\proj__8.net351 ));
 sg13g2_inv_1 \proj__8.not293/_0_  (.Y(\proj__8.net346 ),
    .A(\proj__8.net352 ));
 sg13g2_inv_1 \proj__8.not294/_0_  (.Y(\proj__8.net354 ),
    .A(\proj__8.net353 ));
 sg13g2_inv_1 \proj__8.not295/_0_  (.Y(\proj__8.net355 ),
    .A(\proj__8.net354 ));
 sg13g2_inv_1 \proj__8.not296/_0_  (.Y(\proj__8.net356 ),
    .A(\proj__8.net355 ));
 sg13g2_inv_1 \proj__8.not297/_0_  (.Y(\proj__8.net357 ),
    .A(\proj__8.net356 ));
 sg13g2_inv_1 \proj__8.not298/_0_  (.Y(\proj__8.net359 ),
    .A(\proj__8.net358 ));
 sg13g2_inv_1 \proj__8.not299/_0_  (.Y(\proj__8.net360 ),
    .A(\proj__8.net359 ));
 sg13g2_inv_1 \proj__8.not3/_0_  (.Y(\proj__8.net19 ),
    .A(\proj__8.net21 ));
 sg13g2_inv_1 \proj__8.not30/_0_  (.Y(\proj__8.net85 ),
    .A(\proj__8.net86 ));
 sg13g2_inv_1 \proj__8.not300/_0_  (.Y(\proj__8.net361 ),
    .A(\proj__8.net360 ));
 sg13g2_inv_1 \proj__8.not301/_0_  (.Y(\proj__8.net353 ),
    .A(\proj__8.net361 ));
 sg13g2_inv_1 \proj__8.not302/_0_  (.Y(\proj__8.net363 ),
    .A(\proj__8.net362 ));
 sg13g2_inv_1 \proj__8.not303/_0_  (.Y(\proj__8.net364 ),
    .A(\proj__8.net363 ));
 sg13g2_inv_1 \proj__8.not304/_0_  (.Y(\proj__8.net365 ),
    .A(\proj__8.net364 ));
 sg13g2_inv_1 \proj__8.not305/_0_  (.Y(\proj__8.net366 ),
    .A(\proj__8.net365 ));
 sg13g2_inv_1 \proj__8.not306/_0_  (.Y(\proj__8.net367 ),
    .A(\proj__8.net357 ));
 sg13g2_inv_1 \proj__8.not307/_0_  (.Y(\proj__8.net368 ),
    .A(\proj__8.net367 ));
 sg13g2_inv_1 \proj__8.not308/_0_  (.Y(\proj__8.net369 ),
    .A(\proj__8.net368 ));
 sg13g2_inv_1 \proj__8.not309/_0_  (.Y(\proj__8.net362 ),
    .A(\proj__8.net369 ));
 sg13g2_inv_1 \proj__8.not31/_0_  (.Y(\proj__8.net82 ),
    .A(\proj__8.net84 ));
 sg13g2_inv_1 \proj__8.not310/_0_  (.Y(\proj__8.net371 ),
    .A(\proj__8.net370 ));
 sg13g2_inv_1 \proj__8.not311/_0_  (.Y(\proj__8.net372 ),
    .A(\proj__8.net371 ));
 sg13g2_inv_1 \proj__8.not312/_0_  (.Y(\proj__8.net373 ),
    .A(\proj__8.net372 ));
 sg13g2_inv_1 \proj__8.not313/_0_  (.Y(\proj__8.net374 ),
    .A(\proj__8.net373 ));
 sg13g2_inv_1 \proj__8.not314/_0_  (.Y(\proj__8.net375 ),
    .A(\proj__8.net366 ));
 sg13g2_inv_1 \proj__8.not315/_0_  (.Y(\proj__8.net376 ),
    .A(\proj__8.net375 ));
 sg13g2_inv_1 \proj__8.not316/_0_  (.Y(\proj__8.net377 ),
    .A(\proj__8.net376 ));
 sg13g2_inv_1 \proj__8.not317/_0_  (.Y(\proj__8.net370 ),
    .A(\proj__8.net377 ));
 sg13g2_inv_1 \proj__8.not318/_0_  (.Y(\proj__8.net379 ),
    .A(\proj__8.net378 ));
 sg13g2_inv_1 \proj__8.not319/_0_  (.Y(\proj__8.net380 ),
    .A(\proj__8.net379 ));
 sg13g2_inv_1 \proj__8.not32/_0_  (.Y(\proj__8.net87 ),
    .A(\proj__8.net88 ));
 sg13g2_inv_1 \proj__8.not320/_0_  (.Y(\proj__8.net381 ),
    .A(\proj__8.net380 ));
 sg13g2_inv_1 \proj__8.not321/_0_  (.Y(\proj__8.net382 ),
    .A(\proj__8.net381 ));
 sg13g2_inv_1 \proj__8.not322/_0_  (.Y(\proj__8.net383 ),
    .A(\proj__8.net374 ));
 sg13g2_inv_1 \proj__8.not323/_0_  (.Y(\proj__8.net384 ),
    .A(\proj__8.net383 ));
 sg13g2_inv_1 \proj__8.not324/_0_  (.Y(\proj__8.net385 ),
    .A(\proj__8.net384 ));
 sg13g2_inv_1 \proj__8.not325/_0_  (.Y(\proj__8.net378 ),
    .A(\proj__8.net385 ));
 sg13g2_inv_1 \proj__8.not326/_0_  (.Y(\proj__8.net387 ),
    .A(\proj__8.net386 ));
 sg13g2_inv_1 \proj__8.not327/_0_  (.Y(\proj__8.net388 ),
    .A(\proj__8.net387 ));
 sg13g2_inv_1 \proj__8.not328/_0_  (.Y(\proj__8.net389 ),
    .A(\proj__8.net388 ));
 sg13g2_inv_1 \proj__8.not329/_0_  (.Y(\proj__8.net390 ),
    .A(\proj__8.net389 ));
 sg13g2_inv_1 \proj__8.not33/_0_  (.Y(\proj__8.net89 ),
    .A(\proj__8.net90 ));
 sg13g2_inv_1 \proj__8.not330/_0_  (.Y(\proj__8.net391 ),
    .A(\proj__8.net318 ));
 sg13g2_inv_1 \proj__8.not331/_0_  (.Y(\proj__8.net392 ),
    .A(\proj__8.net391 ));
 sg13g2_inv_1 \proj__8.not332/_0_  (.Y(\proj__8.net393 ),
    .A(\proj__8.net392 ));
 sg13g2_inv_1 \proj__8.not333/_0_  (.Y(\proj__8.net386 ),
    .A(\proj__8.net393 ));
 sg13g2_inv_1 \proj__8.not334/_0_  (.Y(\proj__8.net395 ),
    .A(\proj__8.net394 ));
 sg13g2_inv_1 \proj__8.not335/_0_  (.Y(\proj__8.net396 ),
    .A(\proj__8.net395 ));
 sg13g2_inv_1 \proj__8.not336/_0_  (.Y(\proj__8.net397 ),
    .A(\proj__8.net396 ));
 sg13g2_inv_1 \proj__8.not337/_0_  (.Y(\proj__8.net398 ),
    .A(\proj__8.net397 ));
 sg13g2_inv_1 \proj__8.not338/_0_  (.Y(\proj__8.net399 ),
    .A(\proj__8.net390 ));
 sg13g2_inv_1 \proj__8.not339/_0_  (.Y(\proj__8.net400 ),
    .A(\proj__8.net399 ));
 sg13g2_inv_1 \proj__8.not34/_0_  (.Y(\proj__8.net94 ),
    .A(\proj__8.net95 ));
 sg13g2_inv_1 \proj__8.not340/_0_  (.Y(\proj__8.net401 ),
    .A(\proj__8.net400 ));
 sg13g2_inv_1 \proj__8.not341/_0_  (.Y(\proj__8.net394 ),
    .A(\proj__8.net401 ));
 sg13g2_inv_1 \proj__8.not342/_0_  (.Y(\proj__8.net403 ),
    .A(\proj__8.net402 ));
 sg13g2_inv_1 \proj__8.not343/_0_  (.Y(\proj__8.net404 ),
    .A(\proj__8.net403 ));
 sg13g2_inv_1 \proj__8.not344/_0_  (.Y(\proj__8.net405 ),
    .A(\proj__8.net404 ));
 sg13g2_inv_1 \proj__8.not345/_0_  (.Y(\proj__8.net406 ),
    .A(\proj__8.net405 ));
 sg13g2_inv_1 \proj__8.not346/_0_  (.Y(\proj__8.net407 ),
    .A(\proj__8.net398 ));
 sg13g2_inv_1 \proj__8.not347/_0_  (.Y(\proj__8.net408 ),
    .A(\proj__8.net407 ));
 sg13g2_inv_1 \proj__8.not348/_0_  (.Y(\proj__8.net409 ),
    .A(\proj__8.net408 ));
 sg13g2_inv_1 \proj__8.not349/_0_  (.Y(\proj__8.net402 ),
    .A(\proj__8.net409 ));
 sg13g2_inv_1 \proj__8.not35/_0_  (.Y(\proj__8.net91 ),
    .A(\proj__8.net93 ));
 sg13g2_inv_1 \proj__8.not350/_0_  (.Y(\proj__8.net411 ),
    .A(\proj__8.net410 ));
 sg13g2_inv_1 \proj__8.not351/_0_  (.Y(\proj__8.net412 ),
    .A(\proj__8.net411 ));
 sg13g2_inv_1 \proj__8.not352/_0_  (.Y(\proj__8.net413 ),
    .A(\proj__8.net412 ));
 sg13g2_inv_1 \proj__8.not353/_0_  (.Y(\proj__8.net358 ),
    .A(\proj__8.net413 ));
 sg13g2_inv_1 \proj__8.not354/_0_  (.Y(\proj__8.net414 ),
    .A(\proj__8.net406 ));
 sg13g2_inv_1 \proj__8.not355/_0_  (.Y(\proj__8.net415 ),
    .A(\proj__8.net414 ));
 sg13g2_inv_1 \proj__8.not356/_0_  (.Y(\proj__8.net416 ),
    .A(\proj__8.net415 ));
 sg13g2_inv_1 \proj__8.not357/_0_  (.Y(\proj__8.net410 ),
    .A(\proj__8.net416 ));
 sg13g2_inv_1 \proj__8.not358/_0_  (.Y(\proj__8.net418 ),
    .A(\proj__8.net417 ));
 sg13g2_inv_1 \proj__8.not359/_0_  (.Y(\proj__8.net419 ),
    .A(\proj__8.net418 ));
 sg13g2_inv_1 \proj__8.not36/_0_  (.Y(\proj__8.net96 ),
    .A(\proj__8.net10 ));
 sg13g2_inv_1 \proj__8.not360/_0_  (.Y(\proj__8.net420 ),
    .A(\proj__8.net419 ));
 sg13g2_inv_1 \proj__8.not361/_0_  (.Y(\proj__8.net421 ),
    .A(\proj__8.net420 ));
 sg13g2_inv_1 \proj__8.not362/_0_  (.Y(\proj__8.net423 ),
    .A(\proj__8.net422 ));
 sg13g2_inv_1 \proj__8.not363/_0_  (.Y(\proj__8.net424 ),
    .A(\proj__8.net423 ));
 sg13g2_inv_1 \proj__8.not364/_0_  (.Y(\proj__8.net425 ),
    .A(\proj__8.net424 ));
 sg13g2_inv_1 \proj__8.not365/_0_  (.Y(\proj__8.net417 ),
    .A(\proj__8.net425 ));
 sg13g2_inv_1 \proj__8.not366/_0_  (.Y(\proj__8.net427 ),
    .A(\proj__8.net426 ));
 sg13g2_inv_1 \proj__8.not367/_0_  (.Y(\proj__8.net428 ),
    .A(\proj__8.net427 ));
 sg13g2_inv_1 \proj__8.not368/_0_  (.Y(\proj__8.net429 ),
    .A(\proj__8.net428 ));
 sg13g2_inv_1 \proj__8.not369/_0_  (.Y(\proj__8.net430 ),
    .A(\proj__8.net429 ));
 sg13g2_inv_1 \proj__8.not370/_0_  (.Y(\proj__8.net431 ),
    .A(\proj__8.net421 ));
 sg13g2_inv_1 \proj__8.not371/_0_  (.Y(\proj__8.net432 ),
    .A(\proj__8.net431 ));
 sg13g2_inv_1 \proj__8.not372/_0_  (.Y(\proj__8.net433 ),
    .A(\proj__8.net432 ));
 sg13g2_inv_1 \proj__8.not373/_0_  (.Y(\proj__8.net426 ),
    .A(\proj__8.net433 ));
 sg13g2_inv_1 \proj__8.not374/_0_  (.Y(\proj__8.net435 ),
    .A(\proj__8.net434 ));
 sg13g2_inv_1 \proj__8.not375/_0_  (.Y(\proj__8.net436 ),
    .A(\proj__8.net435 ));
 sg13g2_inv_1 \proj__8.not376/_0_  (.Y(\proj__8.net437 ),
    .A(\proj__8.net436 ));
 sg13g2_inv_1 \proj__8.not377/_0_  (.Y(\proj__8.net438 ),
    .A(\proj__8.net437 ));
 sg13g2_inv_1 \proj__8.not378/_0_  (.Y(\proj__8.net439 ),
    .A(\proj__8.net430 ));
 sg13g2_inv_1 \proj__8.not379/_0_  (.Y(\proj__8.net440 ),
    .A(\proj__8.net439 ));
 sg13g2_inv_1 \proj__8.not38/_0_  (.Y(\proj__8.net98 ),
    .A(\proj__8.net97 ));
 sg13g2_inv_1 \proj__8.not380/_0_  (.Y(\proj__8.net441 ),
    .A(\proj__8.net440 ));
 sg13g2_inv_1 \proj__8.not381/_0_  (.Y(\proj__8.net434 ),
    .A(\proj__8.net441 ));
 sg13g2_inv_1 \proj__8.not382/_0_  (.Y(\proj__8.net443 ),
    .A(\proj__8.net442 ));
 sg13g2_inv_1 \proj__8.not383/_0_  (.Y(\proj__8.net444 ),
    .A(\proj__8.net443 ));
 sg13g2_inv_1 \proj__8.not384/_0_  (.Y(\proj__8.net445 ),
    .A(\proj__8.net444 ));
 sg13g2_inv_1 \proj__8.not385/_0_  (.Y(\proj__8.net446 ),
    .A(\proj__8.net445 ));
 sg13g2_inv_1 \proj__8.not386/_0_  (.Y(\proj__8.net447 ),
    .A(\proj__8.net438 ));
 sg13g2_inv_1 \proj__8.not387/_0_  (.Y(\proj__8.net448 ),
    .A(\proj__8.net447 ));
 sg13g2_inv_1 \proj__8.not388/_0_  (.Y(\proj__8.net449 ),
    .A(\proj__8.net448 ));
 sg13g2_inv_1 \proj__8.not389/_0_  (.Y(\proj__8.net442 ),
    .A(\proj__8.net449 ));
 sg13g2_inv_1 \proj__8.not39/_0_  (.Y(\proj__8.net99 ),
    .A(\proj__8.net98 ));
 sg13g2_inv_1 \proj__8.not390/_0_  (.Y(\proj__8.net451 ),
    .A(\proj__8.net450 ));
 sg13g2_inv_1 \proj__8.not391/_0_  (.Y(\proj__8.net452 ),
    .A(\proj__8.net451 ));
 sg13g2_inv_1 \proj__8.not392/_0_  (.Y(\proj__8.net453 ),
    .A(\proj__8.net452 ));
 sg13g2_inv_1 \proj__8.not393/_0_  (.Y(\proj__8.net454 ),
    .A(\proj__8.net453 ));
 sg13g2_inv_1 \proj__8.not394/_0_  (.Y(\proj__8.net455 ),
    .A(\proj__8.net382 ));
 sg13g2_inv_1 \proj__8.not395/_0_  (.Y(\proj__8.net456 ),
    .A(\proj__8.net455 ));
 sg13g2_inv_1 \proj__8.not396/_0_  (.Y(\proj__8.net457 ),
    .A(\proj__8.net456 ));
 sg13g2_inv_1 \proj__8.not397/_0_  (.Y(\proj__8.net450 ),
    .A(\proj__8.net457 ));
 sg13g2_inv_1 \proj__8.not398/_0_  (.Y(\proj__8.net459 ),
    .A(\proj__8.net458 ));
 sg13g2_inv_1 \proj__8.not399/_0_  (.Y(\proj__8.net460 ),
    .A(\proj__8.net459 ));
 sg13g2_inv_1 \proj__8.not4/_0_  (.Y(\proj__8.net24 ),
    .A(\proj__8.net25 ));
 sg13g2_inv_1 \proj__8.not40/_0_  (.Y(\proj__8.net100 ),
    .A(\proj__8.net99 ));
 sg13g2_inv_1 \proj__8.not400/_0_  (.Y(\proj__8.net461 ),
    .A(\proj__8.net460 ));
 sg13g2_inv_1 \proj__8.not401/_0_  (.Y(\proj__8.net462 ),
    .A(\proj__8.net461 ));
 sg13g2_inv_1 \proj__8.not402/_0_  (.Y(\proj__8.net463 ),
    .A(\proj__8.net454 ));
 sg13g2_inv_1 \proj__8.not403/_0_  (.Y(\proj__8.net464 ),
    .A(\proj__8.net463 ));
 sg13g2_inv_1 \proj__8.not404/_0_  (.Y(\proj__8.net465 ),
    .A(\proj__8.net464 ));
 sg13g2_inv_1 \proj__8.not405/_0_  (.Y(\proj__8.net458 ),
    .A(\proj__8.net465 ));
 sg13g2_inv_1 \proj__8.not406/_0_  (.Y(\proj__8.net467 ),
    .A(\proj__8.net466 ));
 sg13g2_inv_1 \proj__8.not407/_0_  (.Y(\proj__8.net468 ),
    .A(\proj__8.net467 ));
 sg13g2_inv_1 \proj__8.not408/_0_  (.Y(\proj__8.net469 ),
    .A(\proj__8.net468 ));
 sg13g2_inv_1 \proj__8.not409/_0_  (.Y(\proj__8.net470 ),
    .A(\proj__8.net469 ));
 sg13g2_inv_1 \proj__8.not41/_0_  (.Y(\proj__8.net101 ),
    .A(\proj__8.net100 ));
 sg13g2_inv_1 \proj__8.not410/_0_  (.Y(\proj__8.net471 ),
    .A(\proj__8.net462 ));
 sg13g2_inv_1 \proj__8.not411/_0_  (.Y(\proj__8.net472 ),
    .A(\proj__8.net471 ));
 sg13g2_inv_1 \proj__8.not412/_0_  (.Y(\proj__8.net473 ),
    .A(\proj__8.net472 ));
 sg13g2_inv_1 \proj__8.not413/_0_  (.Y(\proj__8.net466 ),
    .A(\proj__8.net473 ));
 sg13g2_inv_1 \proj__8.not414/_0_  (.Y(\proj__8.net475 ),
    .A(\proj__8.net474 ));
 sg13g2_inv_1 \proj__8.not415/_0_  (.Y(\proj__8.net476 ),
    .A(\proj__8.net475 ));
 sg13g2_inv_1 \proj__8.not416/_0_  (.Y(\proj__8.net477 ),
    .A(\proj__8.net476 ));
 sg13g2_inv_1 \proj__8.not417/_0_  (.Y(\proj__8.net422 ),
    .A(\proj__8.net477 ));
 sg13g2_inv_1 \proj__8.not418/_0_  (.Y(\proj__8.net478 ),
    .A(\proj__8.net470 ));
 sg13g2_inv_1 \proj__8.not419/_0_  (.Y(\proj__8.net479 ),
    .A(\proj__8.net478 ));
 sg13g2_inv_1 \proj__8.not42/_0_  (.Y(\proj__8.net103 ),
    .A(\proj__8.net102 ));
 sg13g2_inv_1 \proj__8.not420/_0_  (.Y(\proj__8.net480 ),
    .A(\proj__8.net479 ));
 sg13g2_inv_1 \proj__8.not421/_0_  (.Y(\proj__8.net474 ),
    .A(\proj__8.net480 ));
 sg13g2_inv_1 \proj__8.not43/_0_  (.Y(\proj__8.net104 ),
    .A(\proj__8.net103 ));
 sg13g2_inv_1 \proj__8.not44/_0_  (.Y(\proj__8.net105 ),
    .A(\proj__8.net104 ));
 sg13g2_inv_1 \proj__8.not45/_0_  (.Y(\proj__8.net97 ),
    .A(\proj__8.net105 ));
 sg13g2_inv_1 \proj__8.not46/_0_  (.Y(\proj__8.net107 ),
    .A(\proj__8.net106 ));
 sg13g2_inv_1 \proj__8.not47/_0_  (.Y(\proj__8.net108 ),
    .A(\proj__8.net107 ));
 sg13g2_inv_1 \proj__8.not48/_0_  (.Y(\proj__8.net109 ),
    .A(\proj__8.net108 ));
 sg13g2_inv_1 \proj__8.not49/_0_  (.Y(\proj__8.net110 ),
    .A(\proj__8.net109 ));
 sg13g2_inv_1 \proj__8.not5/_0_  (.Y(\proj__8.net26 ),
    .A(\proj__8.net27 ));
 sg13g2_inv_1 \proj__8.not50/_0_  (.Y(\proj__8.net111 ),
    .A(\proj__8.net101 ));
 sg13g2_inv_1 \proj__8.not51/_0_  (.Y(\proj__8.net112 ),
    .A(\proj__8.net111 ));
 sg13g2_inv_1 \proj__8.not52/_0_  (.Y(\proj__8.net113 ),
    .A(\proj__8.net112 ));
 sg13g2_inv_1 \proj__8.not53/_0_  (.Y(\proj__8.net106 ),
    .A(\proj__8.net113 ));
 sg13g2_inv_1 \proj__8.not54/_0_  (.Y(\proj__8.net115 ),
    .A(\proj__8.net114 ));
 sg13g2_inv_1 \proj__8.not55/_0_  (.Y(\proj__8.net116 ),
    .A(\proj__8.net115 ));
 sg13g2_inv_1 \proj__8.not56/_0_  (.Y(\proj__8.net117 ),
    .A(\proj__8.net116 ));
 sg13g2_inv_1 \proj__8.not57/_0_  (.Y(\proj__8.net118 ),
    .A(\proj__8.net117 ));
 sg13g2_inv_1 \proj__8.not58/_0_  (.Y(\proj__8.net119 ),
    .A(\proj__8.net110 ));
 sg13g2_inv_1 \proj__8.not59/_0_  (.Y(\proj__8.net120 ),
    .A(\proj__8.net119 ));
 sg13g2_inv_1 \proj__8.not6/_0_  (.Y(\proj__8.net31 ),
    .A(\proj__8.net32 ));
 sg13g2_inv_1 \proj__8.not60/_0_  (.Y(\proj__8.net121 ),
    .A(\proj__8.net120 ));
 sg13g2_inv_1 \proj__8.not61/_0_  (.Y(\proj__8.net114 ),
    .A(\proj__8.net121 ));
 sg13g2_inv_1 \proj__8.not62/_0_  (.Y(\proj__8.net123 ),
    .A(\proj__8.net122 ));
 sg13g2_inv_1 \proj__8.not63/_0_  (.Y(\proj__8.net124 ),
    .A(\proj__8.net123 ));
 sg13g2_inv_1 \proj__8.not64/_0_  (.Y(\proj__8.net125 ),
    .A(\proj__8.net124 ));
 sg13g2_inv_1 \proj__8.not65/_0_  (.Y(\proj__8.net126 ),
    .A(\proj__8.net125 ));
 sg13g2_inv_1 \proj__8.not66/_0_  (.Y(\proj__8.net127 ),
    .A(\proj__8.net118 ));
 sg13g2_inv_1 \proj__8.not67/_0_  (.Y(\proj__8.net128 ),
    .A(\proj__8.net127 ));
 sg13g2_inv_1 \proj__8.not68/_0_  (.Y(\proj__8.net129 ),
    .A(\proj__8.net128 ));
 sg13g2_inv_1 \proj__8.not69/_0_  (.Y(\proj__8.net122 ),
    .A(\proj__8.net129 ));
 sg13g2_inv_1 \proj__8.not7/_0_  (.Y(\proj__8.net28 ),
    .A(\proj__8.net30 ));
 sg13g2_inv_1 \proj__8.not70/_0_  (.Y(\proj__8.net131 ),
    .A(\proj__8.net130 ));
 sg13g2_inv_1 \proj__8.not71/_0_  (.Y(\proj__8.net132 ),
    .A(\proj__8.net131 ));
 sg13g2_inv_1 \proj__8.not72/_0_  (.Y(\proj__8.net133 ),
    .A(\proj__8.net132 ));
 sg13g2_inv_1 \proj__8.not73/_0_  (.Y(\proj__8.net134 ),
    .A(\proj__8.net133 ));
 sg13g2_inv_1 \proj__8.not74/_0_  (.Y(\proj__8.net135 ),
    .A(\proj__8.net80 ));
 sg13g2_inv_1 \proj__8.not75/_0_  (.Y(\proj__8.net136 ),
    .A(\proj__8.net135 ));
 sg13g2_inv_1 \proj__8.not76/_0_  (.Y(\proj__8.net137 ),
    .A(\proj__8.net136 ));
 sg13g2_inv_1 \proj__8.not77/_0_  (.Y(\proj__8.net130 ),
    .A(\proj__8.net137 ));
 sg13g2_inv_1 \proj__8.not78/_0_  (.Y(\proj__8.net139 ),
    .A(\proj__8.net138 ));
 sg13g2_inv_1 \proj__8.not79/_0_  (.Y(\proj__8.net140 ),
    .A(\proj__8.net139 ));
 sg13g2_inv_1 \proj__8.not8/_0_  (.Y(\proj__8.net33 ),
    .A(\proj__8.net34 ));
 sg13g2_inv_1 \proj__8.not80/_0_  (.Y(\proj__8.net141 ),
    .A(\proj__8.net140 ));
 sg13g2_inv_1 \proj__8.not81/_0_  (.Y(\proj__8.net142 ),
    .A(\proj__8.net141 ));
 sg13g2_inv_1 \proj__8.not82/_0_  (.Y(\proj__8.net143 ),
    .A(\proj__8.net134 ));
 sg13g2_inv_1 \proj__8.not83/_0_  (.Y(\proj__8.net144 ),
    .A(\proj__8.net143 ));
 sg13g2_inv_1 \proj__8.not84/_0_  (.Y(\proj__8.net145 ),
    .A(\proj__8.net144 ));
 sg13g2_inv_1 \proj__8.not85/_0_  (.Y(\proj__8.net138 ),
    .A(\proj__8.net145 ));
 sg13g2_inv_1 \proj__8.not86/_0_  (.Y(\proj__8.net147 ),
    .A(\proj__8.net146 ));
 sg13g2_inv_1 \proj__8.not87/_0_  (.Y(\proj__8.net148 ),
    .A(\proj__8.net147 ));
 sg13g2_inv_1 \proj__8.not88/_0_  (.Y(\proj__8.net149 ),
    .A(\proj__8.net148 ));
 sg13g2_inv_1 \proj__8.not89/_0_  (.Y(\proj__8.net150 ),
    .A(\proj__8.net149 ));
 sg13g2_inv_1 \proj__8.not9/_0_  (.Y(\proj__8.net35 ),
    .A(\proj__8.net36 ));
 sg13g2_inv_1 \proj__8.not90/_0_  (.Y(\proj__8.net151 ),
    .A(\proj__8.net142 ));
 sg13g2_inv_1 \proj__8.not91/_0_  (.Y(\proj__8.net152 ),
    .A(\proj__8.net151 ));
 sg13g2_inv_1 \proj__8.not92/_0_  (.Y(\proj__8.net153 ),
    .A(\proj__8.net152 ));
 sg13g2_inv_1 \proj__8.not93/_0_  (.Y(\proj__8.net146 ),
    .A(\proj__8.net153 ));
 sg13g2_inv_1 \proj__8.not94/_0_  (.Y(\proj__8.net155 ),
    .A(\proj__8.net154 ));
 sg13g2_inv_1 \proj__8.not95/_0_  (.Y(\proj__8.net156 ),
    .A(\proj__8.net155 ));
 sg13g2_inv_1 \proj__8.not96/_0_  (.Y(\proj__8.net157 ),
    .A(\proj__8.net156 ));
 sg13g2_inv_1 \proj__8.not97/_0_  (.Y(\proj__8.net102 ),
    .A(\proj__8.net157 ));
 sg13g2_inv_1 \proj__8.not98/_0_  (.Y(\proj__8.net158 ),
    .A(\proj__8.net150 ));
 sg13g2_inv_1 \proj__8.not99/_0_  (.Y(\proj__8.net159 ),
    .A(\proj__8.net158 ));
 sg13g2_or2_1 \proj__8.or1/_0_  (.X(\proj__8.net4 ),
    .B(\proj__8.net11 ),
    .A(\proj__8.net446 ));
 sg13g2_and2_1 \proj__9.and1/_0_  (.A(\proj__9.net18 ),
    .B(\proj__9.net18 ),
    .X(\proj__9.net20 ));
 sg13g2_nand2_1 \proj__9.nand1/_0_  (.Y(\proj__9.net17 ),
    .A(net75),
    .B(net75));
 sg13g2_nand2_1 \proj__9.nand10/_0_  (.Y(\proj__9.net25 ),
    .A(net67),
    .B(net67));
 sg13g2_nand2_1 \proj__9.nand11/_0_  (.Y(\proj__9.net26 ),
    .A(net64),
    .B(net64));
 sg13g2_nand2_1 \proj__9.nand12/_0_  (.Y(\proj__9.net27 ),
    .A(\proj__9.net26 ),
    .B(\proj__9.net25 ));
 sg13g2_nand2_1 \proj__9.nand13/_0_  (.Y(\proj__9.net11 ),
    .A(\proj__9.net27 ),
    .B(\proj__9.net27 ));
 sg13g2_nand2_1 \proj__9.nand2/_0_  (.Y(\proj__9.net18 ),
    .A(net75),
    .B(net78));
 sg13g2_nand2_1 \proj__9.nand3/_0_  (.Y(\proj__9.net19 ),
    .A(net78),
    .B(net79));
 sg13g2_nand2_1 \proj__9.nand4/_0_  (.Y(\proj__9.net22 ),
    .A(\proj__9.net21 ),
    .B(\proj__9.net20 ));
 sg13g2_nand2_1 \proj__9.nand5/_0_  (.Y(\proj__9.net7 ),
    .A(\proj__9.net22 ),
    .B(\proj__9.net22 ));
 sg13g2_nand2_1 \proj__9.nand6/_0_  (.Y(\proj__9.net21 ),
    .A(\proj__9.net17 ),
    .B(\proj__9.net19 ));
 sg13g2_nand2_1 \proj__9.nand7/_0_  (.Y(\proj__9.net23 ),
    .A(net72),
    .B(net72));
 sg13g2_nand2_1 \proj__9.nand8/_0_  (.Y(\proj__9.net24 ),
    .A(net70),
    .B(net2));
 sg13g2_nand2_1 \proj__9.nand9/_0_  (.Y(\proj__9.net9 ),
    .A(\proj__9.net24 ),
    .B(\proj__9.net23 ));
 sg13g2_inv_1 \proj__9.not1/_0_  (.Y(\proj__9.net12 ),
    .A(\proj__9.net28 ));
 sg13g2_or2_1 \proj__9.or1/_0_  (.X(\proj__9.net10 ),
    .B(net71),
    .A(net69));
 sg13g2_or2_1 \proj__9.or2/_0_  (.X(\proj__9.net28 ),
    .B(net67),
    .A(net65));
 sg13g2_xor2_1 \proj__9.xor1/_0_  (.B(net79),
    .A(net76),
    .X(\proj__9.net8 ));
 sg13g2_buf_2 fanout61 (.A(ui_in[7]),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(ui_in[7]),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(net4),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(net66),
    .X(net64));
 sg13g2_buf_1 fanout65 (.A(net66),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(ui_in[5]),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(net68),
    .X(net67));
 sg13g2_buf_4 fanout68 (.X(net68),
    .A(net3));
 sg13g2_buf_2 fanout69 (.A(net70),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(net2),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(net73),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(net73),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(ui_in[2]),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(net77),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(net76),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(net77),
    .X(net76));
 sg13g2_buf_1 fanout77 (.A(ui_in[1]),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(net80),
    .X(net78));
 sg13g2_buf_1 fanout79 (.A(net80),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(net81),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(ui_in[0]),
    .X(net81));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[3]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[6]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(uio_in[0]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(uio_in[1]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(uio_in[2]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[3]),
    .X(net8));
 sg13g2_tielo \proj_11.flop1/_5__9  (.L_LO(net9));
 sg13g2_inv_1 \proj__4.not1/_0__2  (.Y(net108),
    .A(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_1_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_1_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_1_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_1_1__leaf_clk_regs));
 sg13g2_buf_1 clkload1 (.A(clknet_1_0__leaf_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(\proj__8.net18 ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold2 (.A(\proj_11.net16 ),
    .X(net110));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_fill_1 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_153 ();
 sg13g2_decap_8 FILLER_13_160 ();
 sg13g2_decap_8 FILLER_13_167 ();
 sg13g2_decap_8 FILLER_13_174 ();
 sg13g2_decap_8 FILLER_13_181 ();
 sg13g2_decap_8 FILLER_13_188 ();
 sg13g2_decap_8 FILLER_13_195 ();
 sg13g2_decap_8 FILLER_13_202 ();
 sg13g2_decap_8 FILLER_13_209 ();
 sg13g2_decap_8 FILLER_13_216 ();
 sg13g2_decap_8 FILLER_13_223 ();
 sg13g2_decap_8 FILLER_13_230 ();
 sg13g2_decap_8 FILLER_13_237 ();
 sg13g2_decap_8 FILLER_13_244 ();
 sg13g2_decap_8 FILLER_13_251 ();
 sg13g2_decap_8 FILLER_13_258 ();
 sg13g2_decap_8 FILLER_13_265 ();
 sg13g2_decap_8 FILLER_13_272 ();
 sg13g2_decap_8 FILLER_13_279 ();
 sg13g2_decap_8 FILLER_13_286 ();
 sg13g2_decap_8 FILLER_13_293 ();
 sg13g2_decap_8 FILLER_13_300 ();
 sg13g2_decap_8 FILLER_13_307 ();
 sg13g2_decap_8 FILLER_13_314 ();
 sg13g2_decap_8 FILLER_13_321 ();
 sg13g2_decap_8 FILLER_13_328 ();
 sg13g2_decap_8 FILLER_13_335 ();
 sg13g2_decap_8 FILLER_13_342 ();
 sg13g2_decap_8 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_356 ();
 sg13g2_decap_8 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_370 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_4 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_155 ();
 sg13g2_fill_1 FILLER_15_162 ();
 sg13g2_decap_8 FILLER_15_166 ();
 sg13g2_fill_2 FILLER_15_173 ();
 sg13g2_decap_8 FILLER_15_179 ();
 sg13g2_fill_2 FILLER_15_212 ();
 sg13g2_decap_8 FILLER_15_218 ();
 sg13g2_decap_8 FILLER_15_225 ();
 sg13g2_decap_8 FILLER_15_232 ();
 sg13g2_decap_8 FILLER_15_239 ();
 sg13g2_decap_8 FILLER_15_246 ();
 sg13g2_decap_8 FILLER_15_253 ();
 sg13g2_decap_8 FILLER_15_260 ();
 sg13g2_decap_8 FILLER_15_267 ();
 sg13g2_decap_8 FILLER_15_274 ();
 sg13g2_decap_8 FILLER_15_281 ();
 sg13g2_decap_8 FILLER_15_288 ();
 sg13g2_decap_8 FILLER_15_295 ();
 sg13g2_decap_8 FILLER_15_302 ();
 sg13g2_decap_8 FILLER_15_309 ();
 sg13g2_decap_8 FILLER_15_316 ();
 sg13g2_decap_8 FILLER_15_323 ();
 sg13g2_decap_8 FILLER_15_330 ();
 sg13g2_decap_8 FILLER_15_337 ();
 sg13g2_decap_8 FILLER_15_344 ();
 sg13g2_decap_8 FILLER_15_351 ();
 sg13g2_decap_8 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_fill_2 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_193 ();
 sg13g2_decap_8 FILLER_16_229 ();
 sg13g2_decap_8 FILLER_16_236 ();
 sg13g2_decap_8 FILLER_16_243 ();
 sg13g2_decap_8 FILLER_16_250 ();
 sg13g2_decap_8 FILLER_16_257 ();
 sg13g2_decap_8 FILLER_16_264 ();
 sg13g2_decap_8 FILLER_16_271 ();
 sg13g2_decap_8 FILLER_16_278 ();
 sg13g2_decap_8 FILLER_16_285 ();
 sg13g2_decap_8 FILLER_16_292 ();
 sg13g2_decap_8 FILLER_16_299 ();
 sg13g2_decap_8 FILLER_16_306 ();
 sg13g2_decap_8 FILLER_16_313 ();
 sg13g2_decap_8 FILLER_16_320 ();
 sg13g2_decap_8 FILLER_16_327 ();
 sg13g2_decap_8 FILLER_16_334 ();
 sg13g2_decap_8 FILLER_16_341 ();
 sg13g2_decap_8 FILLER_16_348 ();
 sg13g2_decap_8 FILLER_16_355 ();
 sg13g2_decap_8 FILLER_16_362 ();
 sg13g2_decap_8 FILLER_16_369 ();
 sg13g2_decap_8 FILLER_16_376 ();
 sg13g2_decap_8 FILLER_16_383 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_decap_8 FILLER_16_397 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_4 FILLER_17_162 ();
 sg13g2_decap_8 FILLER_17_170 ();
 sg13g2_decap_8 FILLER_17_177 ();
 sg13g2_fill_2 FILLER_17_184 ();
 sg13g2_decap_4 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_201 ();
 sg13g2_decap_8 FILLER_17_211 ();
 sg13g2_fill_1 FILLER_17_218 ();
 sg13g2_decap_8 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_230 ();
 sg13g2_decap_8 FILLER_17_237 ();
 sg13g2_decap_8 FILLER_17_244 ();
 sg13g2_decap_8 FILLER_17_251 ();
 sg13g2_decap_8 FILLER_17_258 ();
 sg13g2_decap_8 FILLER_17_265 ();
 sg13g2_decap_8 FILLER_17_272 ();
 sg13g2_decap_8 FILLER_17_279 ();
 sg13g2_decap_8 FILLER_17_286 ();
 sg13g2_decap_8 FILLER_17_293 ();
 sg13g2_decap_8 FILLER_17_300 ();
 sg13g2_decap_8 FILLER_17_307 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_decap_8 FILLER_17_328 ();
 sg13g2_fill_2 FILLER_17_335 ();
 sg13g2_fill_1 FILLER_17_337 ();
 sg13g2_fill_1 FILLER_17_341 ();
 sg13g2_fill_2 FILLER_17_345 ();
 sg13g2_fill_1 FILLER_17_347 ();
 sg13g2_decap_8 FILLER_17_354 ();
 sg13g2_decap_8 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_fill_2 FILLER_18_151 ();
 sg13g2_decap_8 FILLER_18_234 ();
 sg13g2_decap_8 FILLER_18_241 ();
 sg13g2_decap_8 FILLER_18_248 ();
 sg13g2_decap_8 FILLER_18_255 ();
 sg13g2_fill_2 FILLER_18_262 ();
 sg13g2_fill_1 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_271 ();
 sg13g2_fill_1 FILLER_18_275 ();
 sg13g2_decap_4 FILLER_18_279 ();
 sg13g2_fill_1 FILLER_18_283 ();
 sg13g2_fill_1 FILLER_18_287 ();
 sg13g2_decap_4 FILLER_18_291 ();
 sg13g2_fill_1 FILLER_18_295 ();
 sg13g2_fill_1 FILLER_18_299 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_fill_1 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_fill_2 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_327 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_4 FILLER_18_371 ();
 sg13g2_fill_1 FILLER_18_375 ();
 sg13g2_fill_1 FILLER_18_379 ();
 sg13g2_fill_1 FILLER_18_383 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_fill_2 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_167 ();
 sg13g2_decap_8 FILLER_19_174 ();
 sg13g2_decap_4 FILLER_19_181 ();
 sg13g2_fill_2 FILLER_19_185 ();
 sg13g2_decap_4 FILLER_19_190 ();
 sg13g2_decap_8 FILLER_19_198 ();
 sg13g2_fill_2 FILLER_19_205 ();
 sg13g2_fill_1 FILLER_19_207 ();
 sg13g2_fill_2 FILLER_19_211 ();
 sg13g2_fill_1 FILLER_19_213 ();
 sg13g2_decap_8 FILLER_19_218 ();
 sg13g2_decap_8 FILLER_19_225 ();
 sg13g2_decap_8 FILLER_19_232 ();
 sg13g2_decap_4 FILLER_19_239 ();
 sg13g2_fill_1 FILLER_19_246 ();
 sg13g2_decap_8 FILLER_19_334 ();
 sg13g2_decap_8 FILLER_19_341 ();
 sg13g2_fill_2 FILLER_19_348 ();
 sg13g2_fill_1 FILLER_19_389 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_4 FILLER_20_105 ();
 sg13g2_fill_2 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_137 ();
 sg13g2_decap_4 FILLER_20_144 ();
 sg13g2_fill_1 FILLER_20_229 ();
 sg13g2_fill_1 FILLER_20_233 ();
 sg13g2_decap_8 FILLER_20_258 ();
 sg13g2_decap_8 FILLER_20_265 ();
 sg13g2_decap_8 FILLER_20_272 ();
 sg13g2_decap_8 FILLER_20_279 ();
 sg13g2_decap_8 FILLER_20_286 ();
 sg13g2_decap_8 FILLER_20_293 ();
 sg13g2_fill_2 FILLER_20_300 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_decap_4 FILLER_20_354 ();
 sg13g2_fill_2 FILLER_20_358 ();
 sg13g2_decap_8 FILLER_20_375 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_fill_2 FILLER_20_389 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_fill_1 FILLER_21_84 ();
 sg13g2_fill_2 FILLER_21_114 ();
 sg13g2_fill_1 FILLER_21_116 ();
 sg13g2_fill_2 FILLER_21_120 ();
 sg13g2_fill_1 FILLER_21_177 ();
 sg13g2_decap_8 FILLER_21_207 ();
 sg13g2_fill_2 FILLER_21_214 ();
 sg13g2_fill_1 FILLER_21_216 ();
 sg13g2_fill_2 FILLER_21_223 ();
 sg13g2_fill_1 FILLER_21_228 ();
 sg13g2_decap_8 FILLER_21_232 ();
 sg13g2_decap_4 FILLER_21_239 ();
 sg13g2_fill_2 FILLER_21_243 ();
 sg13g2_fill_2 FILLER_21_248 ();
 sg13g2_fill_1 FILLER_21_250 ();
 sg13g2_fill_1 FILLER_21_255 ();
 sg13g2_decap_8 FILLER_21_282 ();
 sg13g2_fill_1 FILLER_21_289 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_fill_1 FILLER_21_346 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_4 FILLER_21_383 ();
 sg13g2_fill_1 FILLER_21_387 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_4 FILLER_22_63 ();
 sg13g2_fill_2 FILLER_22_96 ();
 sg13g2_fill_1 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_103 ();
 sg13g2_decap_8 FILLER_22_110 ();
 sg13g2_decap_4 FILLER_22_117 ();
 sg13g2_fill_1 FILLER_22_121 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_4 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_141 ();
 sg13g2_fill_2 FILLER_22_148 ();
 sg13g2_decap_4 FILLER_22_156 ();
 sg13g2_fill_2 FILLER_22_160 ();
 sg13g2_decap_8 FILLER_22_166 ();
 sg13g2_decap_8 FILLER_22_173 ();
 sg13g2_decap_4 FILLER_22_180 ();
 sg13g2_fill_2 FILLER_22_184 ();
 sg13g2_fill_2 FILLER_22_189 ();
 sg13g2_fill_1 FILLER_22_191 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_fill_1 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_312 ();
 sg13g2_decap_4 FILLER_22_319 ();
 sg13g2_fill_1 FILLER_22_323 ();
 sg13g2_fill_1 FILLER_22_330 ();
 sg13g2_fill_1 FILLER_22_334 ();
 sg13g2_decap_4 FILLER_22_353 ();
 sg13g2_fill_2 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_77 ();
 sg13g2_fill_1 FILLER_23_79 ();
 sg13g2_fill_1 FILLER_23_110 ();
 sg13g2_fill_2 FILLER_23_114 ();
 sg13g2_decap_8 FILLER_23_120 ();
 sg13g2_decap_4 FILLER_23_127 ();
 sg13g2_fill_2 FILLER_23_131 ();
 sg13g2_fill_2 FILLER_23_202 ();
 sg13g2_fill_1 FILLER_23_210 ();
 sg13g2_fill_1 FILLER_23_223 ();
 sg13g2_fill_1 FILLER_23_227 ();
 sg13g2_decap_8 FILLER_23_232 ();
 sg13g2_decap_8 FILLER_23_239 ();
 sg13g2_decap_8 FILLER_23_246 ();
 sg13g2_fill_1 FILLER_23_253 ();
 sg13g2_fill_1 FILLER_23_283 ();
 sg13g2_decap_8 FILLER_23_288 ();
 sg13g2_decap_8 FILLER_23_295 ();
 sg13g2_decap_8 FILLER_23_302 ();
 sg13g2_decap_8 FILLER_23_309 ();
 sg13g2_fill_2 FILLER_23_325 ();
 sg13g2_decap_8 FILLER_23_339 ();
 sg13g2_decap_4 FILLER_23_346 ();
 sg13g2_decap_4 FILLER_23_353 ();
 sg13g2_fill_1 FILLER_23_360 ();
 sg13g2_fill_1 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_4 FILLER_24_84 ();
 sg13g2_decap_4 FILLER_24_91 ();
 sg13g2_decap_4 FILLER_24_99 ();
 sg13g2_fill_2 FILLER_24_103 ();
 sg13g2_decap_8 FILLER_24_131 ();
 sg13g2_fill_2 FILLER_24_138 ();
 sg13g2_decap_4 FILLER_24_146 ();
 sg13g2_fill_2 FILLER_24_150 ();
 sg13g2_decap_4 FILLER_24_156 ();
 sg13g2_fill_2 FILLER_24_160 ();
 sg13g2_decap_8 FILLER_24_188 ();
 sg13g2_fill_2 FILLER_24_195 ();
 sg13g2_fill_2 FILLER_24_223 ();
 sg13g2_fill_1 FILLER_24_225 ();
 sg13g2_decap_4 FILLER_24_230 ();
 sg13g2_fill_1 FILLER_24_234 ();
 sg13g2_decap_4 FILLER_24_267 ();
 sg13g2_fill_2 FILLER_24_271 ();
 sg13g2_decap_8 FILLER_24_332 ();
 sg13g2_decap_4 FILLER_24_339 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_4 FILLER_25_105 ();
 sg13g2_fill_2 FILLER_25_109 ();
 sg13g2_fill_1 FILLER_25_140 ();
 sg13g2_fill_2 FILLER_25_167 ();
 sg13g2_decap_8 FILLER_25_172 ();
 sg13g2_fill_2 FILLER_25_205 ();
 sg13g2_fill_1 FILLER_25_207 ();
 sg13g2_decap_8 FILLER_25_241 ();
 sg13g2_fill_1 FILLER_25_248 ();
 sg13g2_decap_8 FILLER_25_253 ();
 sg13g2_decap_4 FILLER_25_260 ();
 sg13g2_decap_8 FILLER_25_277 ();
 sg13g2_fill_2 FILLER_25_284 ();
 sg13g2_fill_1 FILLER_25_286 ();
 sg13g2_fill_1 FILLER_25_290 ();
 sg13g2_decap_8 FILLER_25_300 ();
 sg13g2_fill_1 FILLER_25_307 ();
 sg13g2_fill_2 FILLER_25_320 ();
 sg13g2_fill_1 FILLER_25_326 ();
 sg13g2_decap_4 FILLER_25_335 ();
 sg13g2_fill_2 FILLER_25_339 ();
 sg13g2_decap_4 FILLER_25_354 ();
 sg13g2_fill_2 FILLER_25_358 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_4 FILLER_26_119 ();
 sg13g2_fill_2 FILLER_26_123 ();
 sg13g2_decap_8 FILLER_26_129 ();
 sg13g2_fill_2 FILLER_26_151 ();
 sg13g2_fill_1 FILLER_26_159 ();
 sg13g2_decap_4 FILLER_26_169 ();
 sg13g2_decap_8 FILLER_26_177 ();
 sg13g2_decap_4 FILLER_26_184 ();
 sg13g2_fill_2 FILLER_26_188 ();
 sg13g2_fill_1 FILLER_26_194 ();
 sg13g2_decap_8 FILLER_26_198 ();
 sg13g2_decap_8 FILLER_26_205 ();
 sg13g2_fill_2 FILLER_26_212 ();
 sg13g2_fill_1 FILLER_26_214 ();
 sg13g2_decap_8 FILLER_26_222 ();
 sg13g2_decap_4 FILLER_26_229 ();
 sg13g2_decap_8 FILLER_26_236 ();
 sg13g2_decap_8 FILLER_26_243 ();
 sg13g2_decap_4 FILLER_26_361 ();
 sg13g2_fill_2 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_4 FILLER_27_133 ();
 sg13g2_decap_4 FILLER_27_152 ();
 sg13g2_fill_2 FILLER_27_156 ();
 sg13g2_decap_8 FILLER_27_167 ();
 sg13g2_decap_8 FILLER_27_174 ();
 sg13g2_decap_8 FILLER_27_181 ();
 sg13g2_decap_8 FILLER_27_188 ();
 sg13g2_decap_8 FILLER_27_195 ();
 sg13g2_fill_2 FILLER_27_202 ();
 sg13g2_fill_1 FILLER_27_267 ();
 sg13g2_decap_8 FILLER_27_272 ();
 sg13g2_decap_8 FILLER_27_279 ();
 sg13g2_decap_8 FILLER_27_300 ();
 sg13g2_fill_2 FILLER_27_307 ();
 sg13g2_fill_1 FILLER_27_313 ();
 sg13g2_decap_4 FILLER_27_319 ();
 sg13g2_decap_8 FILLER_27_327 ();
 sg13g2_fill_2 FILLER_27_334 ();
 sg13g2_fill_1 FILLER_27_336 ();
 sg13g2_decap_4 FILLER_27_345 ();
 sg13g2_decap_8 FILLER_27_359 ();
 sg13g2_decap_8 FILLER_27_366 ();
 sg13g2_decap_8 FILLER_27_376 ();
 sg13g2_fill_2 FILLER_27_383 ();
 sg13g2_fill_1 FILLER_27_397 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_105 ();
 sg13g2_fill_1 FILLER_28_118 ();
 sg13g2_decap_8 FILLER_28_128 ();
 sg13g2_fill_2 FILLER_28_135 ();
 sg13g2_decap_8 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_156 ();
 sg13g2_decap_8 FILLER_28_172 ();
 sg13g2_decap_8 FILLER_28_179 ();
 sg13g2_decap_8 FILLER_28_186 ();
 sg13g2_decap_8 FILLER_28_193 ();
 sg13g2_decap_8 FILLER_28_200 ();
 sg13g2_decap_8 FILLER_28_207 ();
 sg13g2_decap_8 FILLER_28_214 ();
 sg13g2_decap_8 FILLER_28_221 ();
 sg13g2_decap_8 FILLER_28_228 ();
 sg13g2_fill_2 FILLER_28_235 ();
 sg13g2_fill_1 FILLER_28_244 ();
 sg13g2_decap_4 FILLER_28_271 ();
 sg13g2_fill_2 FILLER_28_275 ();
 sg13g2_decap_4 FILLER_28_281 ();
 sg13g2_fill_2 FILLER_28_285 ();
 sg13g2_decap_4 FILLER_28_295 ();
 sg13g2_fill_1 FILLER_28_299 ();
 sg13g2_fill_1 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_324 ();
 sg13g2_fill_2 FILLER_28_331 ();
 sg13g2_fill_1 FILLER_28_367 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_fill_2 FILLER_29_98 ();
 sg13g2_fill_1 FILLER_29_100 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_132 ();
 sg13g2_fill_1 FILLER_29_136 ();
 sg13g2_decap_8 FILLER_29_149 ();
 sg13g2_decap_4 FILLER_29_156 ();
 sg13g2_decap_8 FILLER_29_169 ();
 sg13g2_decap_8 FILLER_29_176 ();
 sg13g2_decap_8 FILLER_29_183 ();
 sg13g2_decap_8 FILLER_29_190 ();
 sg13g2_decap_8 FILLER_29_197 ();
 sg13g2_decap_8 FILLER_29_204 ();
 sg13g2_decap_8 FILLER_29_211 ();
 sg13g2_fill_2 FILLER_29_218 ();
 sg13g2_fill_1 FILLER_29_220 ();
 sg13g2_fill_1 FILLER_29_265 ();
 sg13g2_decap_8 FILLER_29_292 ();
 sg13g2_fill_2 FILLER_29_299 ();
 sg13g2_fill_1 FILLER_29_301 ();
 sg13g2_fill_1 FILLER_29_324 ();
 sg13g2_decap_8 FILLER_29_331 ();
 sg13g2_fill_2 FILLER_29_338 ();
 sg13g2_fill_1 FILLER_29_340 ();
 sg13g2_fill_2 FILLER_29_349 ();
 sg13g2_decap_8 FILLER_29_359 ();
 sg13g2_fill_2 FILLER_29_366 ();
 sg13g2_fill_1 FILLER_29_368 ();
 sg13g2_fill_2 FILLER_29_383 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_4 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_97 ();
 sg13g2_decap_8 FILLER_30_108 ();
 sg13g2_decap_4 FILLER_30_115 ();
 sg13g2_fill_1 FILLER_30_158 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_fill_2 FILLER_30_210 ();
 sg13g2_fill_1 FILLER_30_212 ();
 sg13g2_decap_4 FILLER_30_217 ();
 sg13g2_fill_2 FILLER_30_221 ();
 sg13g2_decap_4 FILLER_30_234 ();
 sg13g2_fill_2 FILLER_30_238 ();
 sg13g2_decap_4 FILLER_30_244 ();
 sg13g2_decap_8 FILLER_30_251 ();
 sg13g2_decap_4 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_262 ();
 sg13g2_decap_8 FILLER_30_279 ();
 sg13g2_fill_2 FILLER_30_286 ();
 sg13g2_fill_1 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_299 ();
 sg13g2_fill_2 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_decap_4 FILLER_30_334 ();
 sg13g2_fill_1 FILLER_30_359 ();
 sg13g2_fill_1 FILLER_30_368 ();
 sg13g2_fill_1 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_fill_2 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_80 ();
 sg13g2_decap_8 FILLER_31_87 ();
 sg13g2_decap_8 FILLER_31_94 ();
 sg13g2_fill_2 FILLER_31_101 ();
 sg13g2_fill_1 FILLER_31_103 ();
 sg13g2_fill_2 FILLER_31_122 ();
 sg13g2_decap_8 FILLER_31_130 ();
 sg13g2_decap_8 FILLER_31_137 ();
 sg13g2_decap_8 FILLER_31_144 ();
 sg13g2_decap_8 FILLER_31_151 ();
 sg13g2_decap_8 FILLER_31_158 ();
 sg13g2_decap_8 FILLER_31_165 ();
 sg13g2_decap_8 FILLER_31_172 ();
 sg13g2_decap_8 FILLER_31_179 ();
 sg13g2_decap_8 FILLER_31_186 ();
 sg13g2_decap_8 FILLER_31_193 ();
 sg13g2_decap_8 FILLER_31_200 ();
 sg13g2_decap_4 FILLER_31_249 ();
 sg13g2_fill_2 FILLER_31_253 ();
 sg13g2_decap_8 FILLER_31_272 ();
 sg13g2_fill_1 FILLER_31_279 ();
 sg13g2_decap_8 FILLER_31_300 ();
 sg13g2_decap_8 FILLER_31_351 ();
 sg13g2_decap_8 FILLER_31_383 ();
 sg13g2_fill_2 FILLER_31_390 ();
 sg13g2_fill_1 FILLER_31_392 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_4 FILLER_32_56 ();
 sg13g2_fill_2 FILLER_32_60 ();
 sg13g2_fill_2 FILLER_32_71 ();
 sg13g2_fill_1 FILLER_32_76 ();
 sg13g2_decap_8 FILLER_32_83 ();
 sg13g2_fill_1 FILLER_32_90 ();
 sg13g2_fill_1 FILLER_32_103 ();
 sg13g2_fill_1 FILLER_32_107 ();
 sg13g2_decap_8 FILLER_32_114 ();
 sg13g2_decap_8 FILLER_32_121 ();
 sg13g2_decap_8 FILLER_32_128 ();
 sg13g2_decap_8 FILLER_32_135 ();
 sg13g2_decap_8 FILLER_32_142 ();
 sg13g2_decap_8 FILLER_32_149 ();
 sg13g2_decap_8 FILLER_32_156 ();
 sg13g2_decap_8 FILLER_32_163 ();
 sg13g2_decap_8 FILLER_32_170 ();
 sg13g2_decap_8 FILLER_32_177 ();
 sg13g2_decap_8 FILLER_32_184 ();
 sg13g2_decap_8 FILLER_32_191 ();
 sg13g2_decap_8 FILLER_32_198 ();
 sg13g2_decap_4 FILLER_32_205 ();
 sg13g2_fill_2 FILLER_32_209 ();
 sg13g2_decap_8 FILLER_32_215 ();
 sg13g2_fill_2 FILLER_32_222 ();
 sg13g2_fill_1 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_232 ();
 sg13g2_decap_8 FILLER_32_239 ();
 sg13g2_fill_2 FILLER_32_246 ();
 sg13g2_fill_1 FILLER_32_248 ();
 sg13g2_fill_2 FILLER_32_262 ();
 sg13g2_fill_1 FILLER_32_270 ();
 sg13g2_decap_4 FILLER_32_276 ();
 sg13g2_fill_1 FILLER_32_280 ();
 sg13g2_fill_1 FILLER_32_306 ();
 sg13g2_fill_2 FILLER_32_320 ();
 sg13g2_fill_1 FILLER_32_322 ();
 sg13g2_fill_2 FILLER_32_335 ();
 sg13g2_decap_8 FILLER_32_376 ();
 sg13g2_decap_4 FILLER_32_383 ();
 sg13g2_fill_1 FILLER_32_387 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_4 FILLER_33_63 ();
 sg13g2_fill_1 FILLER_33_67 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_fill_2 FILLER_33_203 ();
 sg13g2_fill_1 FILLER_33_259 ();
 sg13g2_decap_4 FILLER_33_295 ();
 sg13g2_fill_1 FILLER_33_309 ();
 sg13g2_fill_2 FILLER_33_316 ();
 sg13g2_decap_8 FILLER_33_326 ();
 sg13g2_fill_1 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_360 ();
 sg13g2_decap_8 FILLER_33_367 ();
 sg13g2_fill_2 FILLER_33_374 ();
 sg13g2_decap_4 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_4 FILLER_34_210 ();
 sg13g2_fill_2 FILLER_34_214 ();
 sg13g2_decap_4 FILLER_34_220 ();
 sg13g2_fill_2 FILLER_34_224 ();
 sg13g2_fill_2 FILLER_34_230 ();
 sg13g2_decap_8 FILLER_34_236 ();
 sg13g2_decap_8 FILLER_34_243 ();
 sg13g2_decap_8 FILLER_34_250 ();
 sg13g2_decap_4 FILLER_34_257 ();
 sg13g2_decap_8 FILLER_34_275 ();
 sg13g2_fill_2 FILLER_34_282 ();
 sg13g2_fill_1 FILLER_34_284 ();
 sg13g2_fill_1 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_300 ();
 sg13g2_decap_8 FILLER_34_307 ();
 sg13g2_decap_4 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_335 ();
 sg13g2_fill_2 FILLER_34_342 ();
 sg13g2_fill_1 FILLER_34_344 ();
 sg13g2_fill_2 FILLER_34_355 ();
 sg13g2_fill_1 FILLER_34_357 ();
 sg13g2_fill_2 FILLER_34_362 ();
 sg13g2_fill_1 FILLER_34_364 ();
 sg13g2_fill_2 FILLER_34_379 ();
 sg13g2_fill_1 FILLER_34_381 ();
 sg13g2_decap_4 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_4 FILLER_35_203 ();
 sg13g2_fill_2 FILLER_35_207 ();
 sg13g2_fill_2 FILLER_35_260 ();
 sg13g2_fill_1 FILLER_35_310 ();
 sg13g2_decap_4 FILLER_35_332 ();
 sg13g2_fill_2 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_347 ();
 sg13g2_fill_2 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_234 ();
 sg13g2_decap_8 FILLER_36_241 ();
 sg13g2_decap_4 FILLER_36_248 ();
 sg13g2_fill_2 FILLER_36_252 ();
 sg13g2_fill_1 FILLER_36_259 ();
 sg13g2_fill_1 FILLER_36_275 ();
 sg13g2_decap_4 FILLER_36_296 ();
 sg13g2_fill_1 FILLER_36_300 ();
 sg13g2_decap_4 FILLER_36_312 ();
 sg13g2_decap_8 FILLER_36_326 ();
 sg13g2_fill_2 FILLER_36_338 ();
 sg13g2_fill_1 FILLER_36_345 ();
 sg13g2_decap_4 FILLER_36_362 ();
 sg13g2_fill_1 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_382 ();
 sg13g2_fill_2 FILLER_36_389 ();
 sg13g2_fill_1 FILLER_36_391 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_4 FILLER_37_231 ();
 sg13g2_fill_2 FILLER_37_235 ();
 sg13g2_decap_4 FILLER_37_279 ();
 sg13g2_fill_1 FILLER_37_283 ();
 sg13g2_fill_2 FILLER_37_293 ();
 sg13g2_fill_1 FILLER_37_295 ();
 sg13g2_fill_2 FILLER_37_309 ();
 sg13g2_decap_4 FILLER_37_319 ();
 sg13g2_fill_2 FILLER_37_323 ();
 sg13g2_fill_1 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_380 ();
 sg13g2_decap_8 FILLER_37_387 ();
 sg13g2_decap_8 FILLER_37_394 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_4 FILLER_38_236 ();
 sg13g2_fill_2 FILLER_38_240 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_fill_2 FILLER_38_257 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_fill_1 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_333 ();
 sg13g2_fill_2 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_354 ();
 sg13g2_fill_2 FILLER_38_374 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net17;
 assign uio_oe[1] = net18;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_oe[4] = net21;
 assign uio_oe[5] = net22;
 assign uio_oe[6] = net23;
 assign uio_oe[7] = net24;
 assign uio_out[0] = net25;
 assign uio_out[1] = net26;
 assign uio_out[2] = net27;
 assign uio_out[3] = net28;
 assign uio_out[4] = net29;
 assign uio_out[5] = net30;
 assign uio_out[6] = net31;
 assign uio_out[7] = net32;
endmodule

module tt_um_devinatkin_basys3_uart (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \Led_Cycle_inst.buttons[0] ;
 wire \Led_Cycle_inst.buttons[1] ;
 wire \Led_Cycle_inst.buttons[2] ;
 wire \Led_Cycle_inst.buttons[3] ;
 wire \Led_Cycle_inst.buttons[4] ;
 wire \Led_Cycle_inst.clk_reduced ;
 wire \Led_Cycle_inst.clk_reducer.counter[0] ;
 wire \Led_Cycle_inst.clk_reducer.counter[10] ;
 wire \Led_Cycle_inst.clk_reducer.counter[11] ;
 wire \Led_Cycle_inst.clk_reducer.counter[12] ;
 wire \Led_Cycle_inst.clk_reducer.counter[13] ;
 wire \Led_Cycle_inst.clk_reducer.counter[14] ;
 wire \Led_Cycle_inst.clk_reducer.counter[15] ;
 wire \Led_Cycle_inst.clk_reducer.counter[16] ;
 wire \Led_Cycle_inst.clk_reducer.counter[17] ;
 wire \Led_Cycle_inst.clk_reducer.counter[18] ;
 wire \Led_Cycle_inst.clk_reducer.counter[19] ;
 wire \Led_Cycle_inst.clk_reducer.counter[1] ;
 wire \Led_Cycle_inst.clk_reducer.counter[20] ;
 wire \Led_Cycle_inst.clk_reducer.counter[21] ;
 wire \Led_Cycle_inst.clk_reducer.counter[22] ;
 wire \Led_Cycle_inst.clk_reducer.counter[23] ;
 wire \Led_Cycle_inst.clk_reducer.counter[24] ;
 wire \Led_Cycle_inst.clk_reducer.counter[25] ;
 wire \Led_Cycle_inst.clk_reducer.counter[26] ;
 wire \Led_Cycle_inst.clk_reducer.counter[27] ;
 wire \Led_Cycle_inst.clk_reducer.counter[28] ;
 wire \Led_Cycle_inst.clk_reducer.counter[29] ;
 wire \Led_Cycle_inst.clk_reducer.counter[2] ;
 wire \Led_Cycle_inst.clk_reducer.counter[30] ;
 wire \Led_Cycle_inst.clk_reducer.counter[31] ;
 wire \Led_Cycle_inst.clk_reducer.counter[3] ;
 wire \Led_Cycle_inst.clk_reducer.counter[4] ;
 wire \Led_Cycle_inst.clk_reducer.counter[5] ;
 wire \Led_Cycle_inst.clk_reducer.counter[6] ;
 wire \Led_Cycle_inst.clk_reducer.counter[7] ;
 wire \Led_Cycle_inst.clk_reducer.counter[8] ;
 wire \Led_Cycle_inst.clk_reducer.counter[9] ;
 wire \Led_Cycle_inst.csr.read_ptr[0] ;
 wire \Led_Cycle_inst.csr.read_ptr[1] ;
 wire \Led_Cycle_inst.csr.read_ptr[2] ;
 wire \Led_Cycle_inst.csr.read_ptr[3] ;
 wire \Led_Cycle_inst.genblk1[0].pwm_unit.counter[0] ;
 wire \Led_Cycle_inst.genblk1[0].pwm_unit.counter[1] ;
 wire \Led_Cycle_inst.genblk1[0].pwm_unit.counter[2] ;
 wire \Led_Cycle_inst.genblk1[0].pwm_unit.counter[3] ;
 wire \Led_Cycle_inst.genblk1[0].pwm_unit.counter[4] ;
 wire \Led_Cycle_inst.genblk1[0].pwm_unit.counter[5] ;
 wire \Led_Cycle_inst.genblk1[0].pwm_unit.pwm_out ;
 wire \Led_Cycle_inst.genblk1[10].pwm_unit.counter[0] ;
 wire \Led_Cycle_inst.genblk1[10].pwm_unit.counter[1] ;
 wire \Led_Cycle_inst.genblk1[10].pwm_unit.counter[2] ;
 wire \Led_Cycle_inst.genblk1[10].pwm_unit.counter[3] ;
 wire \Led_Cycle_inst.genblk1[10].pwm_unit.counter[4] ;
 wire \Led_Cycle_inst.genblk1[10].pwm_unit.counter[5] ;
 wire \Led_Cycle_inst.genblk1[10].pwm_unit.pwm_out ;
 wire \Led_Cycle_inst.genblk1[11].pwm_unit.counter[0] ;
 wire \Led_Cycle_inst.genblk1[11].pwm_unit.counter[1] ;
 wire \Led_Cycle_inst.genblk1[11].pwm_unit.counter[2] ;
 wire \Led_Cycle_inst.genblk1[11].pwm_unit.counter[3] ;
 wire \Led_Cycle_inst.genblk1[11].pwm_unit.counter[4] ;
 wire \Led_Cycle_inst.genblk1[11].pwm_unit.counter[5] ;
 wire \Led_Cycle_inst.genblk1[11].pwm_unit.pwm_out ;
 wire \Led_Cycle_inst.genblk1[12].pwm_unit.counter[0] ;
 wire \Led_Cycle_inst.genblk1[12].pwm_unit.counter[1] ;
 wire \Led_Cycle_inst.genblk1[12].pwm_unit.counter[2] ;
 wire \Led_Cycle_inst.genblk1[12].pwm_unit.counter[3] ;
 wire \Led_Cycle_inst.genblk1[12].pwm_unit.counter[4] ;
 wire \Led_Cycle_inst.genblk1[12].pwm_unit.counter[5] ;
 wire \Led_Cycle_inst.genblk1[12].pwm_unit.pwm_out ;
 wire \Led_Cycle_inst.genblk1[13].pwm_unit.counter[0] ;
 wire \Led_Cycle_inst.genblk1[13].pwm_unit.counter[1] ;
 wire \Led_Cycle_inst.genblk1[13].pwm_unit.counter[2] ;
 wire \Led_Cycle_inst.genblk1[13].pwm_unit.counter[3] ;
 wire \Led_Cycle_inst.genblk1[13].pwm_unit.counter[4] ;
 wire \Led_Cycle_inst.genblk1[13].pwm_unit.counter[5] ;
 wire \Led_Cycle_inst.genblk1[13].pwm_unit.pwm_out ;
 wire \Led_Cycle_inst.genblk1[14].pwm_unit.counter[0] ;
 wire \Led_Cycle_inst.genblk1[14].pwm_unit.counter[1] ;
 wire \Led_Cycle_inst.genblk1[14].pwm_unit.counter[2] ;
 wire \Led_Cycle_inst.genblk1[14].pwm_unit.counter[3] ;
 wire \Led_Cycle_inst.genblk1[14].pwm_unit.counter[4] ;
 wire \Led_Cycle_inst.genblk1[14].pwm_unit.counter[5] ;
 wire \Led_Cycle_inst.genblk1[14].pwm_unit.pwm_out ;
 wire \Led_Cycle_inst.genblk1[15].pwm_unit.counter[0] ;
 wire \Led_Cycle_inst.genblk1[15].pwm_unit.counter[1] ;
 wire \Led_Cycle_inst.genblk1[15].pwm_unit.counter[2] ;
 wire \Led_Cycle_inst.genblk1[15].pwm_unit.counter[3] ;
 wire \Led_Cycle_inst.genblk1[15].pwm_unit.counter[4] ;
 wire \Led_Cycle_inst.genblk1[15].pwm_unit.counter[5] ;
 wire \Led_Cycle_inst.genblk1[15].pwm_unit.pwm_out ;
 wire \Led_Cycle_inst.genblk1[1].pwm_unit.counter[0] ;
 wire \Led_Cycle_inst.genblk1[1].pwm_unit.counter[1] ;
 wire \Led_Cycle_inst.genblk1[1].pwm_unit.counter[2] ;
 wire \Led_Cycle_inst.genblk1[1].pwm_unit.counter[3] ;
 wire \Led_Cycle_inst.genblk1[1].pwm_unit.counter[4] ;
 wire \Led_Cycle_inst.genblk1[1].pwm_unit.counter[5] ;
 wire \Led_Cycle_inst.genblk1[1].pwm_unit.pwm_out ;
 wire \Led_Cycle_inst.genblk1[2].pwm_unit.counter[0] ;
 wire \Led_Cycle_inst.genblk1[2].pwm_unit.counter[1] ;
 wire \Led_Cycle_inst.genblk1[2].pwm_unit.counter[2] ;
 wire \Led_Cycle_inst.genblk1[2].pwm_unit.counter[3] ;
 wire \Led_Cycle_inst.genblk1[2].pwm_unit.counter[4] ;
 wire \Led_Cycle_inst.genblk1[2].pwm_unit.counter[5] ;
 wire \Led_Cycle_inst.genblk1[2].pwm_unit.pwm_out ;
 wire \Led_Cycle_inst.genblk1[3].pwm_unit.counter[0] ;
 wire \Led_Cycle_inst.genblk1[3].pwm_unit.counter[1] ;
 wire \Led_Cycle_inst.genblk1[3].pwm_unit.counter[2] ;
 wire \Led_Cycle_inst.genblk1[3].pwm_unit.counter[3] ;
 wire \Led_Cycle_inst.genblk1[3].pwm_unit.counter[4] ;
 wire \Led_Cycle_inst.genblk1[3].pwm_unit.counter[5] ;
 wire \Led_Cycle_inst.genblk1[3].pwm_unit.pwm_out ;
 wire \Led_Cycle_inst.genblk1[4].pwm_unit.counter[0] ;
 wire \Led_Cycle_inst.genblk1[4].pwm_unit.counter[1] ;
 wire \Led_Cycle_inst.genblk1[4].pwm_unit.counter[2] ;
 wire \Led_Cycle_inst.genblk1[4].pwm_unit.counter[3] ;
 wire \Led_Cycle_inst.genblk1[4].pwm_unit.counter[4] ;
 wire \Led_Cycle_inst.genblk1[4].pwm_unit.counter[5] ;
 wire \Led_Cycle_inst.genblk1[4].pwm_unit.pwm_out ;
 wire \Led_Cycle_inst.genblk1[5].pwm_unit.counter[0] ;
 wire \Led_Cycle_inst.genblk1[5].pwm_unit.counter[1] ;
 wire \Led_Cycle_inst.genblk1[5].pwm_unit.counter[2] ;
 wire \Led_Cycle_inst.genblk1[5].pwm_unit.counter[3] ;
 wire \Led_Cycle_inst.genblk1[5].pwm_unit.counter[4] ;
 wire \Led_Cycle_inst.genblk1[5].pwm_unit.counter[5] ;
 wire \Led_Cycle_inst.genblk1[5].pwm_unit.pwm_out ;
 wire \Led_Cycle_inst.genblk1[6].pwm_unit.counter[0] ;
 wire \Led_Cycle_inst.genblk1[6].pwm_unit.counter[1] ;
 wire \Led_Cycle_inst.genblk1[6].pwm_unit.counter[2] ;
 wire \Led_Cycle_inst.genblk1[6].pwm_unit.counter[3] ;
 wire \Led_Cycle_inst.genblk1[6].pwm_unit.counter[4] ;
 wire \Led_Cycle_inst.genblk1[6].pwm_unit.counter[5] ;
 wire \Led_Cycle_inst.genblk1[6].pwm_unit.pwm_out ;
 wire \Led_Cycle_inst.genblk1[7].pwm_unit.counter[0] ;
 wire \Led_Cycle_inst.genblk1[7].pwm_unit.counter[1] ;
 wire \Led_Cycle_inst.genblk1[7].pwm_unit.counter[2] ;
 wire \Led_Cycle_inst.genblk1[7].pwm_unit.counter[3] ;
 wire \Led_Cycle_inst.genblk1[7].pwm_unit.counter[4] ;
 wire \Led_Cycle_inst.genblk1[7].pwm_unit.counter[5] ;
 wire \Led_Cycle_inst.genblk1[7].pwm_unit.pwm_out ;
 wire \Led_Cycle_inst.genblk1[8].pwm_unit.counter[0] ;
 wire \Led_Cycle_inst.genblk1[8].pwm_unit.counter[1] ;
 wire \Led_Cycle_inst.genblk1[8].pwm_unit.counter[2] ;
 wire \Led_Cycle_inst.genblk1[8].pwm_unit.counter[3] ;
 wire \Led_Cycle_inst.genblk1[8].pwm_unit.counter[4] ;
 wire \Led_Cycle_inst.genblk1[8].pwm_unit.counter[5] ;
 wire \Led_Cycle_inst.genblk1[8].pwm_unit.pwm_out ;
 wire \Led_Cycle_inst.genblk1[9].pwm_unit.counter[0] ;
 wire \Led_Cycle_inst.genblk1[9].pwm_unit.counter[1] ;
 wire \Led_Cycle_inst.genblk1[9].pwm_unit.counter[2] ;
 wire \Led_Cycle_inst.genblk1[9].pwm_unit.counter[3] ;
 wire \Led_Cycle_inst.genblk1[9].pwm_unit.counter[4] ;
 wire \Led_Cycle_inst.genblk1[9].pwm_unit.counter[5] ;
 wire \Led_Cycle_inst.genblk1[9].pwm_unit.pwm_out ;
 wire \SegmentDisplay.an[0] ;
 wire \SegmentDisplay.an[1] ;
 wire \SegmentDisplay.an[2] ;
 wire \SegmentDisplay.an[3] ;
 wire \SegmentDisplay.bcd2[0] ;
 wire \SegmentDisplay.bcd2[1] ;
 wire \SegmentDisplay.bcd2[2] ;
 wire \SegmentDisplay.bcd2[3] ;
 wire \SegmentDisplay.bcd3[0] ;
 wire \SegmentDisplay.bcd3[1] ;
 wire \SegmentDisplay.bcd3[2] ;
 wire \SegmentDisplay.bcd3[3] ;
 wire \SegmentDisplay.digit0[0] ;
 wire \SegmentDisplay.digit0[1] ;
 wire \SegmentDisplay.digit0[2] ;
 wire \SegmentDisplay.digit0[3] ;
 wire \SegmentDisplay.digit0[4] ;
 wire \SegmentDisplay.digit0[5] ;
 wire \SegmentDisplay.digit0[6] ;
 wire \SegmentDisplay.digit1[0] ;
 wire \SegmentDisplay.digit1[1] ;
 wire \SegmentDisplay.digit1[2] ;
 wire \SegmentDisplay.digit1[3] ;
 wire \SegmentDisplay.digit1[4] ;
 wire \SegmentDisplay.digit1[5] ;
 wire \SegmentDisplay.digit1[6] ;
 wire \SegmentDisplay.digit2[0] ;
 wire \SegmentDisplay.digit2[1] ;
 wire \SegmentDisplay.digit2[2] ;
 wire \SegmentDisplay.digit2[3] ;
 wire \SegmentDisplay.digit2[4] ;
 wire \SegmentDisplay.digit2[5] ;
 wire \SegmentDisplay.digit2[6] ;
 wire \SegmentDisplay.digit3[0] ;
 wire \SegmentDisplay.digit3[1] ;
 wire \SegmentDisplay.digit3[2] ;
 wire \SegmentDisplay.digit3[3] ;
 wire \SegmentDisplay.digit3[4] ;
 wire \SegmentDisplay.digit3[5] ;
 wire \SegmentDisplay.digit3[6] ;
 wire \SegmentDisplay.out_sel[0] ;
 wire \SegmentDisplay.out_sel[1] ;
 wire \SegmentDisplay.out_sel[2] ;
 wire \SegmentDisplay.out_sel[3] ;
 wire \SegmentDisplay.seg_driver.clk_reduced ;
 wire \SegmentDisplay.seg_driver.clk_reducer.counter[0] ;
 wire \SegmentDisplay.seg_driver.clk_reducer.counter[10] ;
 wire \SegmentDisplay.seg_driver.clk_reducer.counter[11] ;
 wire \SegmentDisplay.seg_driver.clk_reducer.counter[12] ;
 wire \SegmentDisplay.seg_driver.clk_reducer.counter[1] ;
 wire \SegmentDisplay.seg_driver.clk_reducer.counter[2] ;
 wire \SegmentDisplay.seg_driver.clk_reducer.counter[3] ;
 wire \SegmentDisplay.seg_driver.clk_reducer.counter[4] ;
 wire \SegmentDisplay.seg_driver.clk_reducer.counter[5] ;
 wire \SegmentDisplay.seg_driver.clk_reducer.counter[6] ;
 wire \SegmentDisplay.seg_driver.clk_reducer.counter[7] ;
 wire \SegmentDisplay.seg_driver.clk_reducer.counter[8] ;
 wire \SegmentDisplay.seg_driver.clk_reducer.counter[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire \input_value_check_inst.character_buff[0][0] ;
 wire \input_value_check_inst.character_buff[0][1] ;
 wire \input_value_check_inst.character_buff[0][2] ;
 wire \input_value_check_inst.character_buff[0][3] ;
 wire \input_value_check_inst.character_buff[0][4] ;
 wire \input_value_check_inst.character_buff[0][5] ;
 wire \input_value_check_inst.character_buff[0][6] ;
 wire \input_value_check_inst.character_buff[0][7] ;
 wire \input_value_check_inst.character_buff[1][0] ;
 wire \input_value_check_inst.character_buff[1][1] ;
 wire \input_value_check_inst.character_buff[1][2] ;
 wire \input_value_check_inst.character_buff[1][3] ;
 wire \input_value_check_inst.character_buff[1][4] ;
 wire \input_value_check_inst.character_buff[1][5] ;
 wire \input_value_check_inst.character_buff[1][6] ;
 wire \input_value_check_inst.character_buff[1][7] ;
 wire \input_value_check_inst.character_buff[2][0] ;
 wire \input_value_check_inst.character_buff[2][1] ;
 wire \input_value_check_inst.character_buff[2][2] ;
 wire \input_value_check_inst.character_buff[2][3] ;
 wire \input_value_check_inst.character_buff[2][4] ;
 wire \input_value_check_inst.character_buff[2][5] ;
 wire \input_value_check_inst.character_buff[2][6] ;
 wire \input_value_check_inst.character_buff[2][7] ;
 wire \input_value_check_inst.character_buff[3][0] ;
 wire \input_value_check_inst.character_buff[3][1] ;
 wire \input_value_check_inst.character_buff[3][2] ;
 wire \input_value_check_inst.character_buff[3][3] ;
 wire \input_value_check_inst.character_buff[3][4] ;
 wire \input_value_check_inst.character_buff[3][5] ;
 wire \input_value_check_inst.character_buff[3][6] ;
 wire \input_value_check_inst.character_buff[3][7] ;
 wire \input_value_check_inst.character_buff[4][0] ;
 wire \input_value_check_inst.character_buff[4][1] ;
 wire \input_value_check_inst.character_buff[4][2] ;
 wire \input_value_check_inst.character_buff[4][3] ;
 wire \input_value_check_inst.character_buff[4][4] ;
 wire \input_value_check_inst.character_buff[4][5] ;
 wire \input_value_check_inst.character_buff[4][6] ;
 wire \input_value_check_inst.character_buff[4][7] ;
 wire \input_value_check_inst.character_buff[5][0] ;
 wire \input_value_check_inst.character_buff[5][1] ;
 wire \input_value_check_inst.character_buff[5][2] ;
 wire \input_value_check_inst.character_buff[5][3] ;
 wire \input_value_check_inst.character_buff[5][4] ;
 wire \input_value_check_inst.character_buff[5][5] ;
 wire \input_value_check_inst.character_buff[5][6] ;
 wire \input_value_check_inst.character_buff[5][7] ;
 wire \input_value_check_inst.character_buff[6][0] ;
 wire \input_value_check_inst.character_buff[6][1] ;
 wire \input_value_check_inst.character_buff[6][2] ;
 wire \input_value_check_inst.character_buff[6][3] ;
 wire \input_value_check_inst.character_buff[6][4] ;
 wire \input_value_check_inst.character_buff[6][5] ;
 wire \input_value_check_inst.character_buff[6][6] ;
 wire \input_value_check_inst.character_buff[6][7] ;
 wire \input_value_check_inst.character_buff[7][0] ;
 wire \input_value_check_inst.character_buff[7][1] ;
 wire \input_value_check_inst.character_buff[7][2] ;
 wire \input_value_check_inst.character_buff[7][3] ;
 wire \input_value_check_inst.character_buff[7][4] ;
 wire \input_value_check_inst.character_buff[7][5] ;
 wire \input_value_check_inst.character_buff[7][6] ;
 wire \input_value_check_inst.character_buff[7][7] ;
 wire \input_value_check_inst.character_buff[8][0] ;
 wire \input_value_check_inst.character_buff[8][1] ;
 wire \input_value_check_inst.character_buff[8][2] ;
 wire \input_value_check_inst.character_buff[8][3] ;
 wire \input_value_check_inst.character_buff[8][4] ;
 wire \input_value_check_inst.character_buff[8][5] ;
 wire \input_value_check_inst.character_buff[8][6] ;
 wire \input_value_check_inst.character_buff[8][7] ;
 wire \input_value_check_inst.character_buff[9][0] ;
 wire \input_value_check_inst.character_buff[9][1] ;
 wire \input_value_check_inst.character_buff[9][2] ;
 wire \input_value_check_inst.character_buff[9][3] ;
 wire \input_value_check_inst.character_buff[9][4] ;
 wire \input_value_check_inst.character_buff[9][5] ;
 wire \input_value_check_inst.character_buff[9][6] ;
 wire \input_value_check_inst.character_buff[9][7] ;
 wire \output_value_inst.character_buff[0][0] ;
 wire \output_value_inst.character_buff[0][1] ;
 wire \output_value_inst.character_buff[0][2] ;
 wire \output_value_inst.character_buff[0][3] ;
 wire \output_value_inst.character_buff[0][4] ;
 wire \output_value_inst.character_buff[0][5] ;
 wire \output_value_inst.character_buff[0][6] ;
 wire \output_value_inst.character_buff[1][0] ;
 wire \output_value_inst.character_buff[1][1] ;
 wire \output_value_inst.character_buff[1][2] ;
 wire \output_value_inst.character_buff[1][3] ;
 wire \output_value_inst.character_buff[1][4] ;
 wire \output_value_inst.character_buff[1][5] ;
 wire \output_value_inst.character_buff[1][6] ;
 wire \output_value_inst.character_buff[2][0] ;
 wire \output_value_inst.character_buff[2][1] ;
 wire \output_value_inst.character_buff[2][2] ;
 wire \output_value_inst.character_buff[2][3] ;
 wire \output_value_inst.character_buff[2][4] ;
 wire \output_value_inst.character_buff[2][5] ;
 wire \output_value_inst.character_buff[2][6] ;
 wire \output_value_inst.character_buff[3][0] ;
 wire \output_value_inst.character_buff[3][1] ;
 wire \output_value_inst.character_buff[3][2] ;
 wire \output_value_inst.character_buff[3][3] ;
 wire \output_value_inst.character_buff[3][4] ;
 wire \output_value_inst.character_buff[3][5] ;
 wire \output_value_inst.character_buff[3][6] ;
 wire \output_value_inst.character_buff[4][0] ;
 wire \output_value_inst.character_buff[4][1] ;
 wire \output_value_inst.character_buff[4][2] ;
 wire \output_value_inst.character_buff[4][3] ;
 wire \output_value_inst.character_buff[4][4] ;
 wire \output_value_inst.character_buff[4][6] ;
 wire \output_value_inst.character_buff[5][0] ;
 wire \output_value_inst.character_buff[5][1] ;
 wire \output_value_inst.character_buff[5][2] ;
 wire \output_value_inst.character_buff[5][3] ;
 wire \output_value_inst.character_buff[5][4] ;
 wire \output_value_inst.character_buff[5][6] ;
 wire \output_value_inst.character_buff[6][0] ;
 wire \output_value_inst.character_buff[6][1] ;
 wire \output_value_inst.character_buff[6][2] ;
 wire \output_value_inst.character_buff[6][3] ;
 wire \output_value_inst.character_buff[6][4] ;
 wire \output_value_inst.character_buff[6][6] ;
 wire \output_value_inst.character_buff[7][0] ;
 wire \output_value_inst.character_buff[7][1] ;
 wire \output_value_inst.character_buff[7][2] ;
 wire \output_value_inst.character_buff[7][3] ;
 wire \output_value_inst.character_buff[7][4] ;
 wire \output_value_inst.character_buff[7][6] ;
 wire \output_value_inst.character_buff[8][0] ;
 wire \output_value_inst.character_buff[8][1] ;
 wire \output_value_inst.character_buff[8][2] ;
 wire \output_value_inst.character_buff[8][3] ;
 wire \output_value_inst.character_buff[8][4] ;
 wire \output_value_inst.character_buff[8][6] ;
 wire \output_value_inst.character_buff[9][0] ;
 wire \output_value_inst.character_buff[9][1] ;
 wire \output_value_inst.character_buff[9][2] ;
 wire \output_value_inst.character_buff[9][3] ;
 wire \output_value_inst.character_buff[9][4] ;
 wire \output_value_inst.character_buff[9][6] ;
 wire \output_value_inst.element_data_reg[0] ;
 wire \output_value_inst.element_data_reg[10] ;
 wire \output_value_inst.element_data_reg[11] ;
 wire \output_value_inst.element_data_reg[1] ;
 wire \output_value_inst.element_data_reg[2] ;
 wire \output_value_inst.element_data_reg[3] ;
 wire \output_value_inst.element_data_reg[4] ;
 wire \output_value_inst.element_data_reg[5] ;
 wire \output_value_inst.element_data_reg[6] ;
 wire \output_value_inst.element_data_reg[7] ;
 wire \output_value_inst.element_data_reg[8] ;
 wire \output_value_inst.element_data_reg[9] ;
 wire \output_value_inst.led_data_reg[0] ;
 wire \output_value_inst.led_data_reg[10] ;
 wire \output_value_inst.led_data_reg[11] ;
 wire \output_value_inst.led_data_reg[12] ;
 wire \output_value_inst.led_data_reg[13] ;
 wire \output_value_inst.led_data_reg[14] ;
 wire \output_value_inst.led_data_reg[15] ;
 wire \output_value_inst.led_data_reg[1] ;
 wire \output_value_inst.led_data_reg[2] ;
 wire \output_value_inst.led_data_reg[3] ;
 wire \output_value_inst.led_data_reg[4] ;
 wire \output_value_inst.led_data_reg[5] ;
 wire \output_value_inst.led_data_reg[6] ;
 wire \output_value_inst.led_data_reg[7] ;
 wire \output_value_inst.led_data_reg[8] ;
 wire \output_value_inst.led_data_reg[9] ;
 wire \output_value_inst.output_data[0] ;
 wire \output_value_inst.output_data[1] ;
 wire \output_value_inst.output_data[2] ;
 wire \output_value_inst.output_data[3] ;
 wire \output_value_inst.output_data[4] ;
 wire \output_value_inst.output_data[5] ;
 wire \output_value_inst.output_data[6] ;
 wire \output_value_inst.output_valid ;
 wire \output_value_inst.ready_to_send ;
 wire \output_value_inst.send_element_data ;
 wire \output_value_inst.send_led_data ;
 wire \output_value_inst.tx_ready ;
 wire \rx_data[0] ;
 wire \rx_data[1] ;
 wire \rx_data[2] ;
 wire \rx_data[3] ;
 wire \rx_data[4] ;
 wire \rx_data[5] ;
 wire \rx_data[6] ;
 wire \rx_data[7] ;
 wire rx_valid;
 wire \tx_data[0] ;
 wire \tx_data[1] ;
 wire \tx_data[2] ;
 wire \tx_data[3] ;
 wire tx_signal;
 wire tx_valid;
 wire \uart_inst.tx_data[4] ;
 wire \uart_inst.tx_data[5] ;
 wire \uart_inst.tx_data[6] ;
 wire \uart_inst.uart_rx_inst.CLK_CNT[0] ;
 wire \uart_inst.uart_rx_inst.CLK_CNT[1] ;
 wire \uart_inst.uart_rx_inst.CLK_CNT[2] ;
 wire \uart_inst.uart_rx_inst.CLK_CNT[3] ;
 wire \uart_inst.uart_rx_inst.CLK_CNT[4] ;
 wire \uart_inst.uart_rx_inst.CLK_CNT[5] ;
 wire \uart_inst.uart_rx_inst.CLK_CNT[6] ;
 wire \uart_inst.uart_rx_inst.CLK_CNT[7] ;
 wire \uart_inst.uart_rx_inst.CLK_CNT[8] ;
 wire \uart_inst.uart_rx_inst.CLK_CNT[9] ;
 wire \uart_inst.uart_rx_inst.DATA_CNT[0] ;
 wire \uart_inst.uart_rx_inst.DATA_CNT[1] ;
 wire \uart_inst.uart_rx_inst.DATA_CNT[2] ;
 wire \uart_inst.uart_rx_inst.DATA_CNT[3] ;
 wire \uart_inst.uart_rx_inst.DATA_TEMP_REG[0] ;
 wire \uart_inst.uart_rx_inst.DATA_TEMP_REG[1] ;
 wire \uart_inst.uart_rx_inst.DATA_TEMP_REG[2] ;
 wire \uart_inst.uart_rx_inst.DATA_TEMP_REG[3] ;
 wire \uart_inst.uart_rx_inst.DATA_TEMP_REG[4] ;
 wire \uart_inst.uart_rx_inst.DATA_TEMP_REG[5] ;
 wire \uart_inst.uart_rx_inst.DATA_TEMP_REG[6] ;
 wire \uart_inst.uart_rx_inst.DATA_TEMP_REG[7] ;
 wire \uart_inst.uart_rx_inst.SAMPLING_COUNT[0] ;
 wire \uart_inst.uart_rx_inst.SAMPLING_COUNT[1] ;
 wire \uart_inst.uart_rx_inst.SIGNAL_Q[0] ;
 wire \uart_inst.uart_rx_inst.SIGNAL_Q[1] ;
 wire \uart_inst.uart_rx_inst.SIGNAL_Q[2] ;
 wire \uart_inst.uart_rx_inst.SIGNAL_Q[3] ;
 wire \uart_inst.uart_rx_inst.SIGNAL_Q[4] ;
 wire \uart_inst.uart_rx_inst.SIGNAL_R ;
 wire \uart_inst.uart_rx_inst.state[0] ;
 wire \uart_inst.uart_rx_inst.state[1] ;
 wire \uart_inst.uart_rx_inst.state[2] ;
 wire \uart_inst.uart_tx_inst.CLK_CNT[0] ;
 wire \uart_inst.uart_tx_inst.CLK_CNT[1] ;
 wire \uart_inst.uart_tx_inst.CLK_CNT[2] ;
 wire \uart_inst.uart_tx_inst.CLK_CNT[3] ;
 wire \uart_inst.uart_tx_inst.CLK_CNT[4] ;
 wire \uart_inst.uart_tx_inst.CLK_CNT[5] ;
 wire \uart_inst.uart_tx_inst.CLK_CNT[6] ;
 wire \uart_inst.uart_tx_inst.CLK_CNT[7] ;
 wire \uart_inst.uart_tx_inst.CLK_CNT[8] ;
 wire \uart_inst.uart_tx_inst.CLK_CNT[9] ;
 wire \uart_inst.uart_tx_inst.DATA_CNT[0] ;
 wire \uart_inst.uart_tx_inst.DATA_CNT[1] ;
 wire \uart_inst.uart_tx_inst.DATA_CNT[2] ;
 wire \uart_inst.uart_tx_inst.DATA_REG[0] ;
 wire \uart_inst.uart_tx_inst.DATA_REG[1] ;
 wire \uart_inst.uart_tx_inst.DATA_REG[2] ;
 wire \uart_inst.uart_tx_inst.DATA_REG[3] ;
 wire \uart_inst.uart_tx_inst.DATA_REG[4] ;
 wire \uart_inst.uart_tx_inst.DATA_REG[5] ;
 wire \uart_inst.uart_tx_inst.DATA_REG[6] ;
 wire \uart_inst.uart_tx_inst.state[0] ;
 wire \uart_inst.uart_tx_inst.state[1] ;
 wire \uart_inst.uart_tx_inst.state[2] ;
 wire \uart_tx_fifo_inst.fifo[0][0] ;
 wire \uart_tx_fifo_inst.fifo[0][1] ;
 wire \uart_tx_fifo_inst.fifo[0][2] ;
 wire \uart_tx_fifo_inst.fifo[0][3] ;
 wire \uart_tx_fifo_inst.fifo[0][4] ;
 wire \uart_tx_fifo_inst.fifo[0][5] ;
 wire \uart_tx_fifo_inst.fifo[0][6] ;
 wire \uart_tx_fifo_inst.fifo[1][0] ;
 wire \uart_tx_fifo_inst.fifo[1][1] ;
 wire \uart_tx_fifo_inst.fifo[1][2] ;
 wire \uart_tx_fifo_inst.fifo[1][3] ;
 wire \uart_tx_fifo_inst.fifo[1][4] ;
 wire \uart_tx_fifo_inst.fifo[1][5] ;
 wire \uart_tx_fifo_inst.fifo[1][6] ;
 wire \uart_tx_fifo_inst.fifo[2][0] ;
 wire \uart_tx_fifo_inst.fifo[2][1] ;
 wire \uart_tx_fifo_inst.fifo[2][2] ;
 wire \uart_tx_fifo_inst.fifo[2][3] ;
 wire \uart_tx_fifo_inst.fifo[2][4] ;
 wire \uart_tx_fifo_inst.fifo[2][5] ;
 wire \uart_tx_fifo_inst.fifo[2][6] ;
 wire \uart_tx_fifo_inst.fifo[3][0] ;
 wire \uart_tx_fifo_inst.fifo[3][1] ;
 wire \uart_tx_fifo_inst.fifo[3][2] ;
 wire \uart_tx_fifo_inst.fifo[3][3] ;
 wire \uart_tx_fifo_inst.fifo[3][4] ;
 wire \uart_tx_fifo_inst.fifo[3][5] ;
 wire \uart_tx_fifo_inst.fifo[3][6] ;
 wire \uart_tx_fifo_inst.fifo[4][0] ;
 wire \uart_tx_fifo_inst.fifo[4][1] ;
 wire \uart_tx_fifo_inst.fifo[4][2] ;
 wire \uart_tx_fifo_inst.fifo[4][3] ;
 wire \uart_tx_fifo_inst.fifo[4][4] ;
 wire \uart_tx_fifo_inst.fifo[4][5] ;
 wire \uart_tx_fifo_inst.fifo[4][6] ;
 wire \uart_tx_fifo_inst.fifo[5][0] ;
 wire \uart_tx_fifo_inst.fifo[5][1] ;
 wire \uart_tx_fifo_inst.fifo[5][2] ;
 wire \uart_tx_fifo_inst.fifo[5][3] ;
 wire \uart_tx_fifo_inst.fifo[5][4] ;
 wire \uart_tx_fifo_inst.fifo[5][5] ;
 wire \uart_tx_fifo_inst.fifo[5][6] ;
 wire \uart_tx_fifo_inst.fifo[6][0] ;
 wire \uart_tx_fifo_inst.fifo[6][1] ;
 wire \uart_tx_fifo_inst.fifo[6][2] ;
 wire \uart_tx_fifo_inst.fifo[6][3] ;
 wire \uart_tx_fifo_inst.fifo[6][4] ;
 wire \uart_tx_fifo_inst.fifo[6][5] ;
 wire \uart_tx_fifo_inst.fifo[6][6] ;
 wire \uart_tx_fifo_inst.fifo[7][0] ;
 wire \uart_tx_fifo_inst.fifo[7][1] ;
 wire \uart_tx_fifo_inst.fifo[7][2] ;
 wire \uart_tx_fifo_inst.fifo[7][3] ;
 wire \uart_tx_fifo_inst.fifo[7][4] ;
 wire \uart_tx_fifo_inst.fifo[7][5] ;
 wire \uart_tx_fifo_inst.fifo[7][6] ;
 wire \uart_tx_fifo_inst.fifo[8][0] ;
 wire \uart_tx_fifo_inst.fifo[8][1] ;
 wire \uart_tx_fifo_inst.fifo[8][2] ;
 wire \uart_tx_fifo_inst.fifo[8][3] ;
 wire \uart_tx_fifo_inst.fifo[8][4] ;
 wire \uart_tx_fifo_inst.fifo[8][5] ;
 wire \uart_tx_fifo_inst.fifo[8][6] ;
 wire \uart_tx_fifo_inst.fifo[9][0] ;
 wire \uart_tx_fifo_inst.fifo[9][1] ;
 wire \uart_tx_fifo_inst.fifo[9][2] ;
 wire \uart_tx_fifo_inst.fifo[9][3] ;
 wire \uart_tx_fifo_inst.fifo[9][4] ;
 wire \uart_tx_fifo_inst.fifo[9][5] ;
 wire \uart_tx_fifo_inst.fifo[9][6] ;
 wire \uart_tx_fifo_inst.fifo_valid[0] ;
 wire \uart_tx_fifo_inst.fifo_valid[1] ;
 wire \uart_tx_fifo_inst.fifo_valid[2] ;
 wire \uart_tx_fifo_inst.fifo_valid[3] ;
 wire \uart_tx_fifo_inst.fifo_valid[4] ;
 wire \uart_tx_fifo_inst.fifo_valid[5] ;
 wire \uart_tx_fifo_inst.fifo_valid[6] ;
 wire \uart_tx_fifo_inst.fifo_valid[7] ;
 wire \uart_tx_fifo_inst.fifo_valid[8] ;
 wire \uart_tx_fifo_inst.fifo_valid[9] ;
 wire net604;
 wire net4;
 wire net605;
 wire net606;
 wire clknet_leaf_0_clk;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;

 sg13g2_inv_1 _3686_ (.Y(_0762_),
    .A(net1198));
 sg13g2_inv_1 _3687_ (.Y(_0763_),
    .A(net1119));
 sg13g2_inv_1 _3688_ (.Y(_0764_),
    .A(net1323));
 sg13g2_inv_1 _3689_ (.Y(_0765_),
    .A(net1227));
 sg13g2_inv_1 _3690_ (.Y(_0766_),
    .A(net1407));
 sg13g2_inv_1 _3691_ (.Y(_0767_),
    .A(net1314));
 sg13g2_inv_1 _3692_ (.Y(_0768_),
    .A(net1307));
 sg13g2_inv_1 _3693_ (.Y(_0769_),
    .A(net1320));
 sg13g2_inv_1 _3694_ (.Y(_0770_),
    .A(net1350));
 sg13g2_inv_2 _3695_ (.Y(_0771_),
    .A(net879));
 sg13g2_inv_1 _3696_ (.Y(_0772_),
    .A(net1272));
 sg13g2_inv_1 _3697_ (.Y(_0773_),
    .A(\Led_Cycle_inst.genblk1[15].pwm_unit.pwm_out ));
 sg13g2_inv_1 _3698_ (.Y(_0774_),
    .A(net1687));
 sg13g2_inv_1 _3699_ (.Y(_0775_),
    .A(net1182));
 sg13g2_inv_1 _3700_ (.Y(_0776_),
    .A(net1109));
 sg13g2_inv_1 _3701_ (.Y(_0777_),
    .A(net1753));
 sg13g2_inv_1 _3702_ (.Y(_0778_),
    .A(net1121));
 sg13g2_inv_1 _3703_ (.Y(_0779_),
    .A(net1064));
 sg13g2_inv_1 _3704_ (.Y(_0780_),
    .A(net1748));
 sg13g2_inv_1 _3705_ (.Y(_0781_),
    .A(net1164));
 sg13g2_inv_1 _3706_ (.Y(_0782_),
    .A(net1088));
 sg13g2_inv_1 _3707_ (.Y(_0783_),
    .A(net1681));
 sg13g2_inv_1 _3708_ (.Y(_0784_),
    .A(\Led_Cycle_inst.genblk1[2].pwm_unit.pwm_out ));
 sg13g2_inv_1 _3709_ (.Y(_0785_),
    .A(\output_value_inst.led_data_reg[1] ));
 sg13g2_inv_1 _3710_ (.Y(_0786_),
    .A(\Led_Cycle_inst.genblk1[1].pwm_unit.pwm_out ));
 sg13g2_inv_1 _3711_ (.Y(_0787_),
    .A(net1155));
 sg13g2_inv_1 _3712_ (.Y(_0788_),
    .A(uo_out[7]));
 sg13g2_inv_1 _3713_ (.Y(_0789_),
    .A(\SegmentDisplay.an[3] ));
 sg13g2_inv_1 _3714_ (.Y(_0790_),
    .A(\SegmentDisplay.an[1] ));
 sg13g2_inv_1 _3715_ (.Y(_0791_),
    .A(\SegmentDisplay.an[0] ));
 sg13g2_inv_1 _3716_ (.Y(_0792_),
    .A(net1649));
 sg13g2_inv_1 _3717_ (.Y(_0793_),
    .A(net883));
 sg13g2_inv_1 _3718_ (.Y(_0794_),
    .A(net964));
 sg13g2_inv_1 _3719_ (.Y(_0795_),
    .A(net885));
 sg13g2_inv_1 _3720_ (.Y(_0796_),
    .A(net707));
 sg13g2_inv_1 _3721_ (.Y(_0797_),
    .A(net722));
 sg13g2_inv_1 _3722_ (.Y(_0798_),
    .A(net688));
 sg13g2_inv_1 _3723_ (.Y(_0799_),
    .A(net716));
 sg13g2_inv_1 _3724_ (.Y(_0800_),
    .A(net972));
 sg13g2_inv_1 _3725_ (.Y(_0801_),
    .A(net713));
 sg13g2_inv_1 _3726_ (.Y(_0802_),
    .A(net1026));
 sg13g2_inv_1 _3727_ (.Y(_0803_),
    .A(net1145));
 sg13g2_inv_1 _3728_ (.Y(_0804_),
    .A(net1220));
 sg13g2_inv_1 _3729_ (.Y(_0805_),
    .A(net1225));
 sg13g2_inv_1 _3730_ (.Y(_0806_),
    .A(net1081));
 sg13g2_inv_1 _3731_ (.Y(_0807_),
    .A(net1262));
 sg13g2_inv_1 _3732_ (.Y(_0808_),
    .A(net987));
 sg13g2_inv_1 _3733_ (.Y(_0809_),
    .A(net1266));
 sg13g2_inv_1 _3734_ (.Y(_0810_),
    .A(net1472));
 sg13g2_inv_1 _3735_ (.Y(_0811_),
    .A(net1187));
 sg13g2_inv_1 _3736_ (.Y(_0812_),
    .A(net1282));
 sg13g2_inv_1 _3737_ (.Y(_0813_),
    .A(net1296));
 sg13g2_inv_1 _3738_ (.Y(_0814_),
    .A(uo_out[6]));
 sg13g2_inv_1 _3739_ (.Y(_0815_),
    .A(net1420));
 sg13g2_inv_1 _3740_ (.Y(_0816_),
    .A(net1578));
 sg13g2_inv_1 _3741_ (.Y(_0817_),
    .A(net1582));
 sg13g2_inv_1 _3742_ (.Y(_0818_),
    .A(net1339));
 sg13g2_inv_1 _3743_ (.Y(_0819_),
    .A(\uart_tx_fifo_inst.fifo_valid[3] ));
 sg13g2_inv_1 _3744_ (.Y(_0820_),
    .A(net1473));
 sg13g2_inv_1 _3745_ (.Y(_0821_),
    .A(net1507));
 sg13g2_inv_1 _3746_ (.Y(_0822_),
    .A(net1029));
 sg13g2_inv_1 _3747_ (.Y(_0823_),
    .A(net1205));
 sg13g2_inv_1 _3748_ (.Y(_0824_),
    .A(net1066));
 sg13g2_inv_1 _3749_ (.Y(_0825_),
    .A(net1083));
 sg13g2_inv_1 _3750_ (.Y(_0826_),
    .A(net1002));
 sg13g2_inv_1 _3751_ (.Y(_0827_),
    .A(net1041));
 sg13g2_inv_1 _3752_ (.Y(_0828_),
    .A(net1022));
 sg13g2_inv_1 _3753_ (.Y(_0829_),
    .A(net989));
 sg13g2_inv_1 _3754_ (.Y(_0830_),
    .A(net979));
 sg13g2_inv_1 _3755_ (.Y(_0831_),
    .A(net997));
 sg13g2_inv_1 _3756_ (.Y(_0832_),
    .A(net995));
 sg13g2_inv_1 _3757_ (.Y(_0833_),
    .A(net1368));
 sg13g2_inv_1 _3758_ (.Y(_0834_),
    .A(net1300));
 sg13g2_inv_1 _3759_ (.Y(_0835_),
    .A(net1149));
 sg13g2_inv_1 _3760_ (.Y(_0836_),
    .A(net1505));
 sg13g2_inv_1 _3761_ (.Y(_0837_),
    .A(net1447));
 sg13g2_inv_1 _3762_ (.Y(_0838_),
    .A(net1493));
 sg13g2_inv_1 _3763_ (.Y(_0839_),
    .A(net1460));
 sg13g2_inv_1 _3764_ (.Y(_0840_),
    .A(net1645));
 sg13g2_inv_2 _3765_ (.Y(_0841_),
    .A(net1650));
 sg13g2_inv_1 _3766_ (.Y(_0842_),
    .A(net1289));
 sg13g2_inv_1 _3767_ (.Y(_0843_),
    .A(net1325));
 sg13g2_inv_1 _3768_ (.Y(_0844_),
    .A(net1426));
 sg13g2_inv_1 _3769_ (.Y(_0845_),
    .A(net1436));
 sg13g2_inv_1 _3770_ (.Y(_0846_),
    .A(\input_value_check_inst.character_buff[3][0] ));
 sg13g2_inv_1 _3771_ (.Y(_0847_),
    .A(net1348));
 sg13g2_inv_1 _3772_ (.Y(_0848_),
    .A(net1206));
 sg13g2_inv_1 _3773_ (.Y(_0849_),
    .A(net1241));
 sg13g2_inv_1 _3774_ (.Y(_0850_),
    .A(net1284));
 sg13g2_inv_1 _3775_ (.Y(_0851_),
    .A(net1249));
 sg13g2_inv_1 _3776_ (.Y(_0852_),
    .A(net1142));
 sg13g2_inv_1 _3777_ (.Y(_0853_),
    .A(net1171));
 sg13g2_inv_1 _3778_ (.Y(_0854_),
    .A(net1363));
 sg13g2_inv_1 _3779_ (.Y(_0855_),
    .A(net1233));
 sg13g2_inv_1 _3780_ (.Y(_0856_),
    .A(net1268));
 sg13g2_inv_1 _3781_ (.Y(_0857_),
    .A(net1211));
 sg13g2_inv_1 _3782_ (.Y(_0858_),
    .A(net1330));
 sg13g2_inv_1 _3783_ (.Y(_0859_),
    .A(net1168));
 sg13g2_inv_1 _3784_ (.Y(_0860_),
    .A(net1305));
 sg13g2_inv_1 _3785_ (.Y(_0861_),
    .A(net1130));
 sg13g2_inv_1 _3786_ (.Y(_0862_),
    .A(net1322));
 sg13g2_inv_1 _3787_ (.Y(_0863_),
    .A(net1270));
 sg13g2_inv_1 _3788_ (.Y(_0864_),
    .A(net1366));
 sg13g2_inv_1 _3789_ (.Y(_0865_),
    .A(net1295));
 sg13g2_inv_1 _3790_ (.Y(_0866_),
    .A(net1215));
 sg13g2_inv_1 _3791_ (.Y(_0867_),
    .A(net1134));
 sg13g2_inv_1 _3792_ (.Y(_0868_),
    .A(net1252));
 sg13g2_inv_1 _3793_ (.Y(_0869_),
    .A(net1246));
 sg13g2_inv_1 _3794_ (.Y(_0870_),
    .A(net1341));
 sg13g2_inv_1 _3795_ (.Y(_0871_),
    .A(net1153));
 sg13g2_inv_1 _3796_ (.Y(_0872_),
    .A(net1248));
 sg13g2_inv_1 _3797_ (.Y(_0873_),
    .A(net1390));
 sg13g2_inv_1 _3798_ (.Y(_0874_),
    .A(net1044));
 sg13g2_inv_1 _3799_ (.Y(_0875_),
    .A(net1151));
 sg13g2_inv_2 _3800_ (.Y(_0876_),
    .A(net889));
 sg13g2_inv_1 _3801_ (.Y(_0877_),
    .A(net1552));
 sg13g2_inv_1 _3802_ (.Y(_0878_),
    .A(net1562));
 sg13g2_inv_1 _3803_ (.Y(_0879_),
    .A(net1494));
 sg13g2_inv_1 _3804_ (.Y(_0880_),
    .A(net1383));
 sg13g2_inv_1 _3805_ (.Y(_0881_),
    .A(net1385));
 sg13g2_inv_1 _3806_ (.Y(_0882_),
    .A(net1103));
 sg13g2_inv_1 _3807_ (.Y(_0883_),
    .A(net1571));
 sg13g2_inv_1 _3808_ (.Y(_0884_),
    .A(net1072));
 sg13g2_inv_1 _3809_ (.Y(_0885_),
    .A(net1092));
 sg13g2_inv_1 _3810_ (.Y(_0886_),
    .A(net1138));
 sg13g2_inv_1 _3811_ (.Y(_0887_),
    .A(net1038));
 sg13g2_inv_1 _3812_ (.Y(_0888_),
    .A(net1224));
 sg13g2_inv_1 _3813_ (.Y(_0889_),
    .A(net1179));
 sg13g2_inv_1 _3814_ (.Y(_0890_),
    .A(net709));
 sg13g2_inv_1 _3815_ (.Y(_0891_),
    .A(\uart_tx_fifo_inst.fifo[8][6] ));
 sg13g2_inv_1 _3816_ (.Y(_0892_),
    .A(net1419));
 sg13g2_inv_1 _3817_ (.Y(_0893_),
    .A(net1357));
 sg13g2_inv_1 _3818_ (.Y(_0894_),
    .A(\uart_tx_fifo_inst.fifo[8][1] ));
 sg13g2_inv_1 _3819_ (.Y(_0895_),
    .A(\uart_tx_fifo_inst.fifo[8][0] ));
 sg13g2_inv_2 _3820_ (.Y(_0896_),
    .A(net836));
 sg13g2_inv_2 _3821_ (.Y(_0897_),
    .A(net840));
 sg13g2_inv_1 _3822_ (.Y(_0898_),
    .A(net835));
 sg13g2_inv_1 _3823_ (.Y(_0899_),
    .A(net833));
 sg13g2_inv_2 _3824_ (.Y(_0900_),
    .A(net918));
 sg13g2_inv_1 _3825_ (.Y(_0901_),
    .A(net990));
 sg13g2_inv_1 _3826_ (.Y(_0902_),
    .A(net1048));
 sg13g2_inv_1 _3827_ (.Y(_0903_),
    .A(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[4] ));
 sg13g2_inv_1 _3828_ (.Y(_0904_),
    .A(net1068));
 sg13g2_inv_1 _3829_ (.Y(_0905_),
    .A(net1079));
 sg13g2_inv_1 _3830_ (.Y(_0906_),
    .A(net828));
 sg13g2_inv_1 _3831_ (.Y(_0907_),
    .A(net1020));
 sg13g2_inv_1 _3832_ (.Y(_0908_),
    .A(net1034));
 sg13g2_inv_1 _3833_ (.Y(_0909_),
    .A(net1100));
 sg13g2_inv_1 _3834_ (.Y(_0910_),
    .A(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[4] ));
 sg13g2_inv_1 _3835_ (.Y(_0911_),
    .A(net1060));
 sg13g2_inv_1 _3836_ (.Y(_0912_),
    .A(_0103_));
 sg13g2_inv_1 _3837_ (.Y(_0913_),
    .A(net2));
 sg13g2_inv_1 _3838_ (.Y(_0914_),
    .A(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[4] ));
 sg13g2_inv_1 _3839_ (.Y(_0915_),
    .A(net1024));
 sg13g2_inv_1 _3840_ (.Y(_0916_),
    .A(net1095));
 sg13g2_inv_1 _3841_ (.Y(_0917_),
    .A(net1077));
 sg13g2_inv_1 _3842_ (.Y(_0918_),
    .A(net1004));
 sg13g2_inv_1 _3843_ (.Y(_0919_),
    .A(net1042));
 sg13g2_inv_1 _3844_ (.Y(_0920_),
    .A(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[2] ));
 sg13g2_inv_1 _3845_ (.Y(_0921_),
    .A(net1085));
 sg13g2_inv_1 _3846_ (.Y(_0922_),
    .A(net1036));
 sg13g2_inv_1 _3847_ (.Y(_0923_),
    .A(\Led_Cycle_inst.clk_reducer.counter[10] ));
 sg13g2_inv_1 _3848_ (.Y(_0924_),
    .A(net1070));
 sg13g2_inv_1 _3849_ (.Y(_0925_),
    .A(net1761));
 sg13g2_inv_1 _3850_ (.Y(_0926_),
    .A(_0123_));
 sg13g2_inv_1 _3851_ (.Y(_0927_),
    .A(_0128_));
 sg13g2_inv_1 _3852_ (.Y(_0928_),
    .A(_0131_));
 sg13g2_inv_1 _3853_ (.Y(_0929_),
    .A(_0133_));
 sg13g2_inv_1 _3854_ (.Y(_0930_),
    .A(net1756));
 sg13g2_inv_1 _3855_ (.Y(_0931_),
    .A(net1663));
 sg13g2_inv_1 _3856_ (.Y(_0932_),
    .A(_0146_));
 sg13g2_inv_1 _3857_ (.Y(_0933_),
    .A(_0150_));
 sg13g2_inv_1 _3858_ (.Y(_0934_),
    .A(net1770));
 sg13g2_inv_1 _3859_ (.Y(_0935_),
    .A(_0153_));
 sg13g2_inv_1 _3860_ (.Y(_0936_),
    .A(net1751));
 sg13g2_inv_1 _3861_ (.Y(_0937_),
    .A(_0157_));
 sg13g2_inv_1 _3862_ (.Y(_0938_),
    .A(_0158_));
 sg13g2_inv_1 _3863_ (.Y(_0939_),
    .A(net1740));
 sg13g2_inv_2 _3864_ (.Y(_0940_),
    .A(net831));
 sg13g2_inv_1 _3865_ (.Y(_0941_),
    .A(_0168_));
 sg13g2_inv_1 _3866_ (.Y(_0942_),
    .A(net638));
 sg13g2_inv_1 _3867_ (.Y(_0943_),
    .A(_0170_));
 sg13g2_inv_1 _3868_ (.Y(_0944_),
    .A(net642));
 sg13g2_inv_1 _3869_ (.Y(_0945_),
    .A(net659));
 sg13g2_inv_1 _3870_ (.Y(_0946_),
    .A(net669));
 sg13g2_inv_1 _3871_ (.Y(_0947_),
    .A(net644));
 sg13g2_inv_1 _3872_ (.Y(_0948_),
    .A(net667));
 sg13g2_inv_1 _3873_ (.Y(_0949_),
    .A(_0187_));
 sg13g2_inv_1 _3874_ (.Y(_0950_),
    .A(_0188_));
 sg13g2_inv_1 _3875_ (.Y(_0951_),
    .A(net685));
 sg13g2_inv_1 _3876_ (.Y(_0952_),
    .A(net661));
 sg13g2_inv_1 _3877_ (.Y(_0953_),
    .A(net651));
 sg13g2_inv_1 _3878_ (.Y(_0954_),
    .A(net687));
 sg13g2_inv_1 _3879_ (.Y(_0955_),
    .A(_0202_));
 sg13g2_inv_1 _3880_ (.Y(_0956_),
    .A(net624));
 sg13g2_inv_1 _3881_ (.Y(_0957_),
    .A(net631));
 sg13g2_inv_1 _3882_ (.Y(_0958_),
    .A(net614));
 sg13g2_inv_1 _3883_ (.Y(_0959_),
    .A(net616));
 sg13g2_inv_1 _3884_ (.Y(_0960_),
    .A(net622));
 sg13g2_inv_1 _3885_ (.Y(_0961_),
    .A(net620));
 sg13g2_and2_2 _3886_ (.A(\Led_Cycle_inst.csr.read_ptr[1] ),
    .B(net841),
    .X(_0962_));
 sg13g2_nand2_2 _3887_ (.Y(_0963_),
    .A(net839),
    .B(net841));
 sg13g2_nor2_2 _3888_ (.A(net834),
    .B(_0963_),
    .Y(_0964_));
 sg13g2_nor2_1 _3889_ (.A(net833),
    .B(_0964_),
    .Y(_0965_));
 sg13g2_xnor2_1 _3890_ (.Y(_0205_),
    .A(net826),
    .B(_0964_));
 sg13g2_nand2_1 _3891_ (.Y(_0966_),
    .A(_0896_),
    .B(net838));
 sg13g2_xnor2_1 _3892_ (.Y(_0967_),
    .A(net836),
    .B(_0962_));
 sg13g2_inv_1 _3893_ (.Y(_0204_),
    .A(_0967_));
 sg13g2_nor2b_2 _3894_ (.A(net840),
    .B_N(net838),
    .Y(_0968_));
 sg13g2_nand2_2 _3895_ (.Y(_0969_),
    .A(net838),
    .B(_0897_));
 sg13g2_nor2_2 _3896_ (.A(net838),
    .B(_0897_),
    .Y(_0970_));
 sg13g2_nand2b_2 _3897_ (.Y(_0971_),
    .B(net840),
    .A_N(net839));
 sg13g2_nand2_1 _3898_ (.Y(_0203_),
    .A(_0969_),
    .B(_0971_));
 sg13g2_nand2_1 _3899_ (.Y(_0972_),
    .A(net941),
    .B(net890));
 sg13g2_nor2_1 _3900_ (.A(net1331),
    .B(\uart_inst.uart_rx_inst.CLK_CNT[0] ),
    .Y(_0973_));
 sg13g2_or4_2 _3901_ (.A(\uart_inst.uart_rx_inst.CLK_CNT[3] ),
    .B(\uart_inst.uart_rx_inst.CLK_CNT[2] ),
    .C(\uart_inst.uart_rx_inst.CLK_CNT[1] ),
    .D(\uart_inst.uart_rx_inst.CLK_CNT[0] ),
    .X(_0974_));
 sg13g2_nor3_1 _3902_ (.A(\uart_inst.uart_rx_inst.CLK_CNT[5] ),
    .B(net1783),
    .C(_0974_),
    .Y(_0975_));
 sg13g2_or4_1 _3903_ (.A(\uart_inst.uart_rx_inst.CLK_CNT[6] ),
    .B(\uart_inst.uart_rx_inst.CLK_CNT[5] ),
    .C(\uart_inst.uart_rx_inst.CLK_CNT[4] ),
    .D(_0974_),
    .X(_0976_));
 sg13g2_nor4_2 _3904_ (.A(net1430),
    .B(\uart_inst.uart_rx_inst.CLK_CNT[8] ),
    .C(\uart_inst.uart_rx_inst.CLK_CNT[7] ),
    .Y(_0977_),
    .D(_0976_));
 sg13g2_or4_2 _3905_ (.A(\uart_inst.uart_rx_inst.CLK_CNT[9] ),
    .B(\uart_inst.uart_rx_inst.CLK_CNT[8] ),
    .C(\uart_inst.uart_rx_inst.CLK_CNT[7] ),
    .D(_0976_),
    .X(_0978_));
 sg13g2_nor2_1 _3906_ (.A(net913),
    .B(_0978_),
    .Y(_0979_));
 sg13g2_nand3_1 _3907_ (.B(net1387),
    .C(net1280),
    .A(net1500),
    .Y(_0980_));
 sg13g2_nor2_1 _3908_ (.A(net680),
    .B(_0980_),
    .Y(_0981_));
 sg13g2_nand2_1 _3909_ (.Y(_0982_),
    .A(_0979_),
    .B(_0981_));
 sg13g2_nand2b_1 _3910_ (.Y(_0983_),
    .B(_0982_),
    .A_N(_0972_));
 sg13g2_nor2_2 _3911_ (.A(net914),
    .B(net908),
    .Y(_0984_));
 sg13g2_nand2_2 _3912_ (.Y(_0985_),
    .A(net962),
    .B(net954));
 sg13g2_nand2b_1 _3913_ (.Y(_0986_),
    .B(net1529),
    .A_N(net1356));
 sg13g2_o21ai_1 _3914_ (.B1(_0983_),
    .Y(_0050_),
    .A1(_0985_),
    .A2(_0986_));
 sg13g2_a21oi_1 _3915_ (.A1(\uart_inst.uart_rx_inst.state[2] ),
    .A2(_0977_),
    .Y(_0987_),
    .B1(\uart_inst.uart_rx_inst.state[0] ));
 sg13g2_nor3_1 _3916_ (.A(net704),
    .B(_0985_),
    .C(_0987_),
    .Y(_0988_));
 sg13g2_a21oi_1 _3917_ (.A1(net913),
    .A2(\uart_inst.uart_rx_inst.state[0] ),
    .Y(_0989_),
    .B1(net705));
 sg13g2_nand2_1 _3918_ (.Y(_0049_),
    .A(net940),
    .B(net706));
 sg13g2_nor2_1 _3919_ (.A(net1361),
    .B(\uart_inst.uart_tx_inst.CLK_CNT[0] ),
    .Y(_0990_));
 sg13g2_nor4_2 _3920_ (.A(net1651),
    .B(\uart_inst.uart_tx_inst.CLK_CNT[2] ),
    .C(\uart_inst.uart_tx_inst.CLK_CNT[1] ),
    .Y(_0991_),
    .D(\uart_inst.uart_tx_inst.CLK_CNT[0] ));
 sg13g2_or4_2 _3921_ (.A(\uart_inst.uart_tx_inst.CLK_CNT[9] ),
    .B(\uart_inst.uart_tx_inst.CLK_CNT[8] ),
    .C(\uart_inst.uart_tx_inst.CLK_CNT[7] ),
    .D(\uart_inst.uart_tx_inst.CLK_CNT[6] ),
    .X(_0992_));
 sg13g2_nor2_1 _3922_ (.A(\uart_inst.uart_tx_inst.CLK_CNT[5] ),
    .B(\uart_inst.uart_tx_inst.CLK_CNT[4] ),
    .Y(_0993_));
 sg13g2_nand2_2 _3923_ (.Y(_0994_),
    .A(_0991_),
    .B(_0993_));
 sg13g2_nor2_2 _3924_ (.A(_0992_),
    .B(_0994_),
    .Y(_0995_));
 sg13g2_nor3_1 _3925_ (.A(net914),
    .B(_0992_),
    .C(_0994_),
    .Y(_0996_));
 sg13g2_nand2_1 _3926_ (.Y(_0997_),
    .A(\uart_inst.uart_tx_inst.DATA_CNT[1] ),
    .B(\uart_inst.uart_tx_inst.DATA_CNT[0] ));
 sg13g2_nor2_1 _3927_ (.A(_0108_),
    .B(_0997_),
    .Y(_0998_));
 sg13g2_nand2_1 _3928_ (.Y(_0999_),
    .A(net808),
    .B(_0998_));
 sg13g2_nand4_1 _3929_ (.B(\uart_inst.uart_tx_inst.state[1] ),
    .C(net808),
    .A(net952),
    .Y(_1000_),
    .D(_0998_));
 sg13g2_nand2_1 _3930_ (.Y(_1001_),
    .A(net954),
    .B(net1546));
 sg13g2_o21ai_1 _3931_ (.B1(_1000_),
    .Y(_0054_),
    .A1(net808),
    .A2(_1001_));
 sg13g2_nand2_1 _3932_ (.Y(_1002_),
    .A(net1546),
    .B(net808));
 sg13g2_nand2b_1 _3933_ (.Y(_1003_),
    .B(net1678),
    .A_N(net808));
 sg13g2_nor2b_1 _3934_ (.A(tx_valid),
    .B_N(\uart_inst.uart_tx_inst.state[0] ),
    .Y(_1004_));
 sg13g2_nand2_1 _3935_ (.Y(_1005_),
    .A(_0107_),
    .B(\uart_inst.uart_tx_inst.state[0] ));
 sg13g2_nor2b_1 _3936_ (.A(_1004_),
    .B_N(_1005_),
    .Y(_1006_));
 sg13g2_nand4_1 _3937_ (.B(_1002_),
    .C(_1003_),
    .A(net952),
    .Y(_0052_),
    .D(_1006_));
 sg13g2_nand3_1 _3938_ (.B(net1575),
    .C(_0999_),
    .A(net952),
    .Y(_1007_));
 sg13g2_nand3_1 _3939_ (.B(\uart_inst.uart_tx_inst.state[0] ),
    .C(net808),
    .A(net1213),
    .Y(_1008_));
 sg13g2_nand2b_1 _3940_ (.Y(_1009_),
    .B(net952),
    .A_N(_0107_));
 sg13g2_o21ai_1 _3941_ (.B1(net1576),
    .Y(_0053_),
    .A1(_1008_),
    .A2(_1009_));
 sg13g2_and2_1 _3942_ (.A(net1356),
    .B(_0979_),
    .X(_1010_));
 sg13g2_nand3b_1 _3943_ (.B(net1598),
    .C(net941),
    .Y(_1011_),
    .A_N(_1010_));
 sg13g2_o21ai_1 _3944_ (.B1(_1011_),
    .Y(_0051_),
    .A1(_0972_),
    .A2(_0982_));
 sg13g2_and3_1 _3945_ (.X(_1012_),
    .A(\input_value_check_inst.character_buff[9][4] ),
    .B(\input_value_check_inst.character_buff[9][1] ),
    .C(\input_value_check_inst.character_buff[9][0] ));
 sg13g2_nor2_1 _3946_ (.A(net913),
    .B(\input_value_check_inst.character_buff[9][5] ),
    .Y(_1013_));
 sg13g2_nand4_1 _3947_ (.B(\input_value_check_inst.character_buff[8][0] ),
    .C(_1012_),
    .A(\input_value_check_inst.character_buff[8][1] ),
    .Y(_1014_),
    .D(_1013_));
 sg13g2_nor4_1 _3948_ (.A(\input_value_check_inst.character_buff[9][7] ),
    .B(_0874_),
    .C(\input_value_check_inst.character_buff[9][3] ),
    .D(\input_value_check_inst.character_buff[9][2] ),
    .Y(_1015_));
 sg13g2_nor4_1 _3949_ (.A(\input_value_check_inst.character_buff[8][5] ),
    .B(_0870_),
    .C(\input_value_check_inst.character_buff[8][3] ),
    .D(_0872_),
    .Y(_1016_));
 sg13g2_nor4_1 _3950_ (.A(\input_value_check_inst.character_buff[6][3] ),
    .B(\input_value_check_inst.character_buff[6][2] ),
    .C(\input_value_check_inst.character_buff[6][1] ),
    .D(\input_value_check_inst.character_buff[6][0] ),
    .Y(_1017_));
 sg13g2_nor4_2 _3951_ (.A(\input_value_check_inst.character_buff[6][7] ),
    .B(\input_value_check_inst.character_buff[6][6] ),
    .C(_0858_),
    .Y(_1018_),
    .D(\input_value_check_inst.character_buff[6][4] ));
 sg13g2_nor4_1 _3952_ (.A(\input_value_check_inst.character_buff[5][3] ),
    .B(\input_value_check_inst.character_buff[5][2] ),
    .C(\input_value_check_inst.character_buff[5][1] ),
    .D(\input_value_check_inst.character_buff[5][0] ),
    .Y(_1019_));
 sg13g2_nor4_1 _3953_ (.A(_0850_),
    .B(\input_value_check_inst.character_buff[4][2] ),
    .C(\input_value_check_inst.character_buff[4][1] ),
    .D(\input_value_check_inst.character_buff[4][0] ),
    .Y(_1020_));
 sg13g2_nor4_1 _3954_ (.A(\input_value_check_inst.character_buff[4][7] ),
    .B(_0847_),
    .C(_0848_),
    .D(_0849_),
    .Y(_1021_));
 sg13g2_nor4_1 _3955_ (.A(_0865_),
    .B(\input_value_check_inst.character_buff[7][2] ),
    .C(_0866_),
    .D(\input_value_check_inst.character_buff[7][0] ),
    .Y(_1022_));
 sg13g2_and4_1 _3956_ (.A(_0863_),
    .B(_0864_),
    .C(\input_value_check_inst.character_buff[7][5] ),
    .D(\input_value_check_inst.character_buff[7][4] ),
    .X(_1023_));
 sg13g2_nand4_1 _3957_ (.B(_1018_),
    .C(_1022_),
    .A(_1017_),
    .Y(_1024_),
    .D(_1023_));
 sg13g2_nor4_1 _3958_ (.A(\input_value_check_inst.character_buff[5][7] ),
    .B(\input_value_check_inst.character_buff[5][6] ),
    .C(_0854_),
    .D(_0855_),
    .Y(_1025_));
 sg13g2_nand4_1 _3959_ (.B(_1020_),
    .C(_1021_),
    .A(_1019_),
    .Y(_1026_),
    .D(_1025_));
 sg13g2_nand4_1 _3960_ (.B(\input_value_check_inst.character_buff[8][6] ),
    .C(_1015_),
    .A(_0868_),
    .Y(_1027_),
    .D(_1016_));
 sg13g2_nor4_2 _3961_ (.A(_1014_),
    .B(_1024_),
    .C(_1026_),
    .Y(_1028_),
    .D(_1027_));
 sg13g2_inv_1 _3962_ (.Y(_1029_),
    .A(net798));
 sg13g2_o21ai_1 _3963_ (.B1(\input_value_check_inst.character_buff[1][3] ),
    .Y(_1030_),
    .A1(\input_value_check_inst.character_buff[1][2] ),
    .A2(\input_value_check_inst.character_buff[1][1] ));
 sg13g2_nor2_1 _3964_ (.A(\input_value_check_inst.character_buff[1][7] ),
    .B(\input_value_check_inst.character_buff[1][6] ),
    .Y(_1031_));
 sg13g2_and4_2 _3965_ (.A(\input_value_check_inst.character_buff[1][5] ),
    .B(\input_value_check_inst.character_buff[1][4] ),
    .C(_1030_),
    .D(_1031_),
    .X(_1032_));
 sg13g2_nand2_1 _3966_ (.Y(_1033_),
    .A(\input_value_check_inst.character_buff[1][1] ),
    .B(\input_value_check_inst.character_buff[1][0] ));
 sg13g2_nand3_1 _3967_ (.B(\input_value_check_inst.character_buff[1][1] ),
    .C(\input_value_check_inst.character_buff[1][0] ),
    .A(\input_value_check_inst.character_buff[1][2] ),
    .Y(_1034_));
 sg13g2_nand2b_1 _3968_ (.Y(_1035_),
    .B(\input_value_check_inst.character_buff[1][6] ),
    .A_N(\input_value_check_inst.character_buff[1][7] ));
 sg13g2_nor3_1 _3969_ (.A(\input_value_check_inst.character_buff[1][4] ),
    .B(\input_value_check_inst.character_buff[1][3] ),
    .C(_1035_),
    .Y(_1036_));
 sg13g2_nor3_1 _3970_ (.A(\input_value_check_inst.character_buff[1][2] ),
    .B(\input_value_check_inst.character_buff[1][1] ),
    .C(\input_value_check_inst.character_buff[1][0] ),
    .Y(_1037_));
 sg13g2_nor4_1 _3971_ (.A(\input_value_check_inst.character_buff[1][4] ),
    .B(\input_value_check_inst.character_buff[1][3] ),
    .C(_1035_),
    .D(_1037_),
    .Y(_1038_));
 sg13g2_a21oi_1 _3972_ (.A1(_1034_),
    .A2(_1038_),
    .Y(_1039_),
    .B1(_1032_));
 sg13g2_nor3_1 _3973_ (.A(_0116_),
    .B(_1032_),
    .C(_1033_),
    .Y(_1040_));
 sg13g2_nor2_1 _3974_ (.A(_1039_),
    .B(_1040_),
    .Y(_1041_));
 sg13g2_nand2_1 _3975_ (.Y(_1042_),
    .A(net1569),
    .B(_1032_));
 sg13g2_nand3_1 _3976_ (.B(_1041_),
    .C(_1042_),
    .A(net798),
    .Y(_1043_));
 sg13g2_o21ai_1 _3977_ (.B1(_1043_),
    .Y(_1044_),
    .A1(net1779),
    .A2(net798));
 sg13g2_nand2_2 _3978_ (.Y(_1045_),
    .A(net940),
    .B(_1044_));
 sg13g2_inv_1 _3979_ (.Y(_1046_),
    .A(_1045_));
 sg13g2_o21ai_1 _3980_ (.B1(_0116_),
    .Y(_1047_),
    .A1(_1032_),
    .A2(_1033_));
 sg13g2_nand3_1 _3981_ (.B(_1041_),
    .C(_1047_),
    .A(net798),
    .Y(_1048_));
 sg13g2_o21ai_1 _3982_ (.B1(_1048_),
    .Y(_1049_),
    .A1(_0814_),
    .A2(net798));
 sg13g2_xor2_1 _3983_ (.B(\input_value_check_inst.character_buff[1][0] ),
    .A(\input_value_check_inst.character_buff[1][1] ),
    .X(_1050_));
 sg13g2_a22oi_1 _3984_ (.Y(_1051_),
    .B1(_1036_),
    .B2(_1050_),
    .A2(_1032_),
    .A1(_0925_));
 sg13g2_o21ai_1 _3985_ (.B1(net940),
    .Y(_1052_),
    .A1(uo_out[5]),
    .A2(net796));
 sg13g2_a21o_1 _3986_ (.A2(_1051_),
    .A1(net798),
    .B1(_1052_),
    .X(_1053_));
 sg13g2_inv_1 _3987_ (.Y(_0605_),
    .A(_1053_));
 sg13g2_or3_2 _3988_ (.A(_1045_),
    .B(_1049_),
    .C(_0605_),
    .X(_1054_));
 sg13g2_mux2_1 _3989_ (.A0(\input_value_check_inst.character_buff[1][0] ),
    .A1(_0117_),
    .S(_1032_),
    .X(_1055_));
 sg13g2_or2_2 _3990_ (.X(_1056_),
    .B(_1055_),
    .A(_1039_));
 sg13g2_o21ai_1 _3991_ (.B1(net940),
    .Y(_1057_),
    .A1(net1769),
    .A2(net796));
 sg13g2_a21o_1 _3992_ (.A2(_1056_),
    .A1(net796),
    .B1(_1057_),
    .X(_1058_));
 sg13g2_inv_1 _3993_ (.Y(_0604_),
    .A(_1058_));
 sg13g2_and2_1 _3994_ (.A(_1053_),
    .B(_1058_),
    .X(_1059_));
 sg13g2_nor2_1 _3995_ (.A(_1053_),
    .B(_1058_),
    .Y(_1060_));
 sg13g2_nand2_2 _3996_ (.Y(_1061_),
    .A(net940),
    .B(_1049_));
 sg13g2_inv_1 _3997_ (.Y(_0606_),
    .A(_1061_));
 sg13g2_nor2_1 _3998_ (.A(_1060_),
    .B(_1061_),
    .Y(_1062_));
 sg13g2_nor2_1 _3999_ (.A(_1059_),
    .B(_1061_),
    .Y(_1063_));
 sg13g2_nor3_1 _4000_ (.A(_1059_),
    .B(_1060_),
    .C(_1061_),
    .Y(_1064_));
 sg13g2_o21ai_1 _4001_ (.B1(_1054_),
    .Y(_0008_),
    .A1(_1046_),
    .A2(_1064_));
 sg13g2_nor2_1 _4002_ (.A(_1053_),
    .B(_0604_),
    .Y(_1065_));
 sg13g2_and2_1 _4003_ (.A(_1061_),
    .B(_1065_),
    .X(_1066_));
 sg13g2_o21ai_1 _4004_ (.B1(_1054_),
    .Y(_0009_),
    .A1(_1046_),
    .A2(_1066_));
 sg13g2_nor2_1 _4005_ (.A(_1049_),
    .B(_1053_),
    .Y(_1067_));
 sg13g2_a21o_1 _4006_ (.A2(_1061_),
    .A1(_1058_),
    .B1(_1067_),
    .X(_1068_));
 sg13g2_o21ai_1 _4007_ (.B1(_1045_),
    .Y(_1069_),
    .A1(_1064_),
    .A2(_1068_));
 sg13g2_nand2_1 _4008_ (.Y(_0010_),
    .A(_1054_),
    .B(_1069_));
 sg13g2_a22oi_1 _4009_ (.Y(_1070_),
    .B1(_1065_),
    .B2(_1045_),
    .A2(_1061_),
    .A1(_1059_));
 sg13g2_inv_1 _4010_ (.Y(_0011_),
    .A(_1070_));
 sg13g2_o21ai_1 _4011_ (.B1(_1045_),
    .Y(_1071_),
    .A1(_1059_),
    .A2(_1062_));
 sg13g2_nand2_1 _4012_ (.Y(_0012_),
    .A(_1054_),
    .B(_1071_));
 sg13g2_o21ai_1 _4013_ (.B1(_1045_),
    .Y(_1072_),
    .A1(_1062_),
    .A2(_1067_));
 sg13g2_nand2_1 _4014_ (.Y(_0013_),
    .A(_1054_),
    .B(_1072_));
 sg13g2_xnor2_1 _4015_ (.Y(_1073_),
    .A(\output_value_inst.led_data_reg[7] ),
    .B(\Led_Cycle_inst.genblk1[7].pwm_unit.pwm_out ));
 sg13g2_xor2_1 _4016_ (.B(\Led_Cycle_inst.genblk1[5].pwm_unit.pwm_out ),
    .A(\output_value_inst.led_data_reg[5] ),
    .X(_1074_));
 sg13g2_xor2_1 _4017_ (.B(\Led_Cycle_inst.genblk1[8].pwm_unit.pwm_out ),
    .A(\output_value_inst.led_data_reg[8] ),
    .X(_1075_));
 sg13g2_xor2_1 _4018_ (.B(\Led_Cycle_inst.genblk1[4].pwm_unit.pwm_out ),
    .A(\output_value_inst.led_data_reg[4] ),
    .X(_1076_));
 sg13g2_xor2_1 _4019_ (.B(\Led_Cycle_inst.genblk1[14].pwm_unit.pwm_out ),
    .A(\output_value_inst.led_data_reg[14] ),
    .X(_1077_));
 sg13g2_a22oi_1 _4020_ (.Y(_1078_),
    .B1(\output_value_inst.led_data_reg[1] ),
    .B2(_0786_),
    .A2(\Led_Cycle_inst.genblk1[15].pwm_unit.pwm_out ),
    .A1(_0772_));
 sg13g2_xor2_1 _4021_ (.B(\Led_Cycle_inst.genblk1[3].pwm_unit.pwm_out ),
    .A(\output_value_inst.led_data_reg[3] ),
    .X(_1079_));
 sg13g2_xor2_1 _4022_ (.B(\Led_Cycle_inst.genblk1[11].pwm_unit.pwm_out ),
    .A(\output_value_inst.led_data_reg[11] ),
    .X(_1080_));
 sg13g2_xor2_1 _4023_ (.B(\Led_Cycle_inst.genblk1[6].pwm_unit.pwm_out ),
    .A(\output_value_inst.led_data_reg[6] ),
    .X(_1081_));
 sg13g2_xor2_1 _4024_ (.B(\Led_Cycle_inst.genblk1[10].pwm_unit.pwm_out ),
    .A(\output_value_inst.led_data_reg[10] ),
    .X(_1082_));
 sg13g2_xor2_1 _4025_ (.B(\Led_Cycle_inst.genblk1[13].pwm_unit.pwm_out ),
    .A(\output_value_inst.led_data_reg[13] ),
    .X(_1083_));
 sg13g2_xor2_1 _4026_ (.B(\Led_Cycle_inst.genblk1[12].pwm_unit.pwm_out ),
    .A(\output_value_inst.led_data_reg[12] ),
    .X(_1084_));
 sg13g2_xor2_1 _4027_ (.B(\Led_Cycle_inst.genblk1[9].pwm_unit.pwm_out ),
    .A(\output_value_inst.led_data_reg[9] ),
    .X(_1085_));
 sg13g2_xor2_1 _4028_ (.B(\Led_Cycle_inst.genblk1[0].pwm_unit.pwm_out ),
    .A(\output_value_inst.led_data_reg[0] ),
    .X(_1086_));
 sg13g2_nor4_2 _4029_ (.A(_1074_),
    .B(_1076_),
    .C(_1081_),
    .Y(_1087_),
    .D(_1083_));
 sg13g2_a221oi_1 _4030_ (.B2(\Led_Cycle_inst.genblk1[2].pwm_unit.pwm_out ),
    .C1(_1080_),
    .B1(_0783_),
    .A1(\output_value_inst.led_data_reg[15] ),
    .Y(_1088_),
    .A2(_0773_));
 sg13g2_a22oi_1 _4031_ (.Y(_1089_),
    .B1(_0785_),
    .B2(\Led_Cycle_inst.genblk1[1].pwm_unit.pwm_out ),
    .A2(_0784_),
    .A1(\output_value_inst.led_data_reg[2] ));
 sg13g2_nand4_1 _4032_ (.B(_1087_),
    .C(_1088_),
    .A(_1078_),
    .Y(_1090_),
    .D(_1089_));
 sg13g2_nor3_1 _4033_ (.A(_1079_),
    .B(_1084_),
    .C(_1085_),
    .Y(_1091_));
 sg13g2_nor4_1 _4034_ (.A(_1075_),
    .B(_1077_),
    .C(_1082_),
    .D(_1086_),
    .Y(_1092_));
 sg13g2_nand3_1 _4035_ (.B(_1091_),
    .C(_1092_),
    .A(_1073_),
    .Y(_1093_));
 sg13g2_o21ai_1 _4036_ (.B1(net963),
    .Y(_1094_),
    .A1(_1090_),
    .A2(_1093_));
 sg13g2_a21oi_1 _4037_ (.A1(net1656),
    .A2(net792),
    .Y(_1095_),
    .B1(net901));
 sg13g2_o21ai_1 _4038_ (.B1(_1095_),
    .Y(_1096_),
    .A1(_0926_),
    .A2(net792));
 sg13g2_mux2_1 _4039_ (.A0(net1759),
    .A1(\output_value_inst.led_data_reg[1] ),
    .S(net793),
    .X(_1097_));
 sg13g2_nand2_1 _4040_ (.Y(_1098_),
    .A(net949),
    .B(net1760));
 sg13g2_inv_1 _4041_ (.Y(_0696_),
    .A(_1098_));
 sg13g2_a21oi_1 _4042_ (.A1(_0783_),
    .A2(net792),
    .Y(_1099_),
    .B1(net901));
 sg13g2_o21ai_1 _4043_ (.B1(_1099_),
    .Y(_1100_),
    .A1(\Led_Cycle_inst.genblk1[2].pwm_unit.pwm_out ),
    .A2(net792));
 sg13g2_inv_1 _4044_ (.Y(_0697_),
    .A(net1682));
 sg13g2_a21oi_1 _4045_ (.A1(_1098_),
    .A2(_1100_),
    .Y(_0720_),
    .B1(net1657));
 sg13g2_inv_1 _4046_ (.Y(_0378_),
    .A(_0720_));
 sg13g2_nand2b_1 _4047_ (.Y(_1101_),
    .B(net793),
    .A_N(net1734));
 sg13g2_o21ai_1 _4048_ (.B1(_1101_),
    .Y(_1102_),
    .A1(net1697),
    .A2(net793));
 sg13g2_nand3b_1 _4049_ (.B(net1698),
    .C(net949),
    .Y(_1103_),
    .A_N(_0720_));
 sg13g2_o21ai_1 _4050_ (.B1(_1103_),
    .Y(_0028_),
    .A1(_0378_),
    .A2(net1698));
 sg13g2_nor3_1 _4051_ (.A(_1096_),
    .B(_1097_),
    .C(_1102_),
    .Y(_1104_));
 sg13g2_nand2_1 _4052_ (.Y(_1105_),
    .A(_1097_),
    .B(net1698));
 sg13g2_a22oi_1 _4053_ (.Y(_1106_),
    .B1(_0697_),
    .B2(_1104_),
    .A2(_0696_),
    .A1(net1657));
 sg13g2_o21ai_1 _4054_ (.B1(_1106_),
    .Y(_0029_),
    .A1(net1657),
    .A2(net1699));
 sg13g2_nor2_1 _4055_ (.A(net1682),
    .B(net1735),
    .Y(_0030_));
 sg13g2_nor2_1 _4056_ (.A(\input_value_check_inst.character_buff[2][7] ),
    .B(\input_value_check_inst.character_buff[2][6] ),
    .Y(_1107_));
 sg13g2_nand2_1 _4057_ (.Y(_1108_),
    .A(\input_value_check_inst.character_buff[2][5] ),
    .B(\input_value_check_inst.character_buff[2][4] ));
 sg13g2_nor2b_1 _4058_ (.A(\input_value_check_inst.character_buff[2][6] ),
    .B_N(_0129_),
    .Y(_1109_));
 sg13g2_nor2_1 _4059_ (.A(\input_value_check_inst.character_buff[2][2] ),
    .B(\input_value_check_inst.character_buff[2][1] ),
    .Y(_1110_));
 sg13g2_nand3_1 _4060_ (.B(\input_value_check_inst.character_buff[2][4] ),
    .C(\input_value_check_inst.character_buff[2][3] ),
    .A(\input_value_check_inst.character_buff[2][5] ),
    .Y(_1111_));
 sg13g2_o21ai_1 _4061_ (.B1(_1109_),
    .Y(_1112_),
    .A1(_1110_),
    .A2(_1111_));
 sg13g2_nor2b_1 _4062_ (.A(\input_value_check_inst.character_buff[2][1] ),
    .B_N(\input_value_check_inst.character_buff[2][0] ),
    .Y(_1113_));
 sg13g2_nand4_1 _4063_ (.B(_0839_),
    .C(_1107_),
    .A(\input_value_check_inst.character_buff[2][3] ),
    .Y(_1114_),
    .D(_1113_));
 sg13g2_a22oi_1 _4064_ (.Y(_1115_),
    .B1(_1112_),
    .B2(_1114_),
    .A2(_1108_),
    .A1(_1107_));
 sg13g2_a21oi_1 _4065_ (.A1(\input_value_check_inst.character_buff[2][6] ),
    .A2(\input_value_check_inst.character_buff[2][5] ),
    .Y(_1116_),
    .B1(_0129_));
 sg13g2_nand2_1 _4066_ (.Y(_1117_),
    .A(\input_value_check_inst.character_buff[2][1] ),
    .B(\input_value_check_inst.character_buff[2][0] ));
 sg13g2_nand3_1 _4067_ (.B(\input_value_check_inst.character_buff[2][1] ),
    .C(\input_value_check_inst.character_buff[2][0] ),
    .A(\input_value_check_inst.character_buff[2][2] ),
    .Y(_1118_));
 sg13g2_nor2_1 _4068_ (.A(\input_value_check_inst.character_buff[2][4] ),
    .B(\input_value_check_inst.character_buff[2][3] ),
    .Y(_1119_));
 sg13g2_a21oi_1 _4069_ (.A1(_1118_),
    .A2(_1119_),
    .Y(_1120_),
    .B1(_1116_));
 sg13g2_and3_1 _4070_ (.X(_1121_),
    .A(_0841_),
    .B(_0129_),
    .C(_1110_));
 sg13g2_nor4_1 _4071_ (.A(\input_value_check_inst.character_buff[2][7] ),
    .B(_1109_),
    .C(_1120_),
    .D(_1121_),
    .Y(_1122_));
 sg13g2_nor2b_1 _4072_ (.A(_1115_),
    .B_N(_1122_),
    .Y(_1123_));
 sg13g2_xor2_1 _4073_ (.B(\input_value_check_inst.character_buff[2][0] ),
    .A(\input_value_check_inst.character_buff[2][1] ),
    .X(_1124_));
 sg13g2_a22oi_1 _4074_ (.Y(_1125_),
    .B1(_1123_),
    .B2(_1124_),
    .A2(_1115_),
    .A1(_0927_));
 sg13g2_nor2_1 _4075_ (.A(net782),
    .B(_1125_),
    .Y(_1126_));
 sg13g2_mux2_1 _4076_ (.A0(net1744),
    .A1(_1125_),
    .S(net795),
    .X(_1127_));
 sg13g2_nand2b_1 _4077_ (.Y(_1128_),
    .B(net1764),
    .A_N(net795));
 sg13g2_o21ai_1 _4078_ (.B1(_0132_),
    .Y(_1129_),
    .A1(_1115_),
    .A2(_1117_));
 sg13g2_nor2_1 _4079_ (.A(_0132_),
    .B(_1117_),
    .Y(_1130_));
 sg13g2_nor2b_1 _4080_ (.A(_1130_),
    .B_N(_1122_),
    .Y(_1131_));
 sg13g2_o21ai_1 _4081_ (.B1(_1129_),
    .Y(_1132_),
    .A1(_1115_),
    .A2(_1131_));
 sg13g2_o21ai_1 _4082_ (.B1(_1128_),
    .Y(_1133_),
    .A1(net783),
    .A2(_1132_));
 sg13g2_inv_1 _4083_ (.Y(_1134_),
    .A(_1133_));
 sg13g2_nor2_1 _4084_ (.A(net1746),
    .B(_1028_),
    .Y(_1135_));
 sg13g2_xnor2_1 _4085_ (.Y(_1136_),
    .A(\input_value_check_inst.character_buff[2][3] ),
    .B(_1130_));
 sg13g2_nand2_1 _4086_ (.Y(_1137_),
    .A(_1123_),
    .B(_1136_));
 sg13g2_a21oi_1 _4087_ (.A1(_0929_),
    .A2(_1115_),
    .Y(_1138_),
    .B1(net782));
 sg13g2_a21oi_1 _4088_ (.A1(_1137_),
    .A2(_1138_),
    .Y(_1139_),
    .B1(_1135_));
 sg13g2_and2_2 _4089_ (.A(net930),
    .B(net1747),
    .X(_0611_));
 sg13g2_nand3_1 _4090_ (.B(_1134_),
    .C(_0611_),
    .A(_1127_),
    .Y(_1140_));
 sg13g2_and2_1 _4091_ (.A(net930),
    .B(_1133_),
    .X(_0610_));
 sg13g2_a22oi_1 _4092_ (.Y(_1141_),
    .B1(_1123_),
    .B2(_0841_),
    .A2(_1115_),
    .A1(_0928_));
 sg13g2_nor2_1 _4093_ (.A(net782),
    .B(_1141_),
    .Y(_1142_));
 sg13g2_mux2_2 _4094_ (.A0(net1667),
    .A1(_1141_),
    .S(net795),
    .X(_1143_));
 sg13g2_nor2_1 _4095_ (.A(net894),
    .B(_1143_),
    .Y(_1144_));
 sg13g2_a21oi_1 _4096_ (.A1(_1127_),
    .A2(_1144_),
    .Y(_1145_),
    .B1(_0610_));
 sg13g2_nand2b_1 _4097_ (.Y(_1146_),
    .B(net930),
    .A_N(_1127_));
 sg13g2_a21oi_1 _4098_ (.A1(_1127_),
    .A2(_1143_),
    .Y(_1147_),
    .B1(net894));
 sg13g2_a21oi_1 _4099_ (.A1(_1133_),
    .A2(_1147_),
    .Y(_1148_),
    .B1(_1145_));
 sg13g2_o21ai_1 _4100_ (.B1(_1140_),
    .Y(_0014_),
    .A1(_0611_),
    .A2(_1148_));
 sg13g2_or2_1 _4101_ (.X(_1149_),
    .B(_1143_),
    .A(_1127_));
 sg13g2_nand2_1 _4102_ (.Y(_1150_),
    .A(_0610_),
    .B(_1149_));
 sg13g2_nand3_1 _4103_ (.B(_1147_),
    .C(_1149_),
    .A(_0610_),
    .Y(_1151_));
 sg13g2_nand2b_1 _4104_ (.Y(_1152_),
    .B(_1151_),
    .A_N(_0611_));
 sg13g2_nand2_1 _4105_ (.Y(_0015_),
    .A(_1140_),
    .B(_1152_));
 sg13g2_nor2_1 _4106_ (.A(_1133_),
    .B(_1146_),
    .Y(_1153_));
 sg13g2_and2_1 _4107_ (.A(_1143_),
    .B(_1153_),
    .X(_1154_));
 sg13g2_o21ai_1 _4108_ (.B1(_1140_),
    .Y(_0016_),
    .A1(_0611_),
    .A2(_1154_));
 sg13g2_nor2b_1 _4109_ (.A(_1145_),
    .B_N(_1151_),
    .Y(_1155_));
 sg13g2_o21ai_1 _4110_ (.B1(_1140_),
    .Y(_0017_),
    .A1(_0611_),
    .A2(_1155_));
 sg13g2_or2_1 _4111_ (.X(_1156_),
    .B(_1147_),
    .A(_0610_));
 sg13g2_nand2b_1 _4112_ (.Y(_1157_),
    .B(_1143_),
    .A_N(_1139_));
 sg13g2_o21ai_1 _4113_ (.B1(_1156_),
    .Y(_0018_),
    .A1(_1146_),
    .A2(net1668));
 sg13g2_and2_1 _4114_ (.A(_1150_),
    .B(_1156_),
    .X(_1158_));
 sg13g2_o21ai_1 _4115_ (.B1(_1140_),
    .Y(_0019_),
    .A1(_0611_),
    .A2(_1158_));
 sg13g2_a21oi_1 _4116_ (.A1(_0610_),
    .A2(_1149_),
    .Y(_1159_),
    .B1(_1153_));
 sg13g2_o21ai_1 _4117_ (.B1(_1140_),
    .Y(_0020_),
    .A1(_0611_),
    .A2(_1159_));
 sg13g2_a21oi_1 _4118_ (.A1(net1646),
    .A2(net792),
    .Y(_1160_),
    .B1(net901));
 sg13g2_o21ai_1 _4119_ (.B1(_1160_),
    .Y(_1161_),
    .A1(_0930_),
    .A2(net792));
 sg13g2_mux2_2 _4120_ (.A0(net1762),
    .A1(\output_value_inst.led_data_reg[13] ),
    .S(net790),
    .X(_1162_));
 sg13g2_nand2_1 _4121_ (.Y(_1163_),
    .A(net945),
    .B(net1763));
 sg13g2_inv_1 _4122_ (.Y(_0708_),
    .A(_1163_));
 sg13g2_a21oi_1 _4123_ (.A1(_0774_),
    .A2(net794),
    .Y(_1164_),
    .B1(net901));
 sg13g2_o21ai_1 _4124_ (.B1(_1164_),
    .Y(_1165_),
    .A1(\Led_Cycle_inst.genblk1[14].pwm_unit.pwm_out ),
    .A2(net794));
 sg13g2_inv_1 _4125_ (.Y(_0709_),
    .A(net1688));
 sg13g2_a21oi_1 _4126_ (.A1(_1163_),
    .A2(_1165_),
    .Y(_0533_),
    .B1(net1647));
 sg13g2_inv_1 _4127_ (.Y(_0379_),
    .A(_0533_));
 sg13g2_nand2b_1 _4128_ (.Y(_1166_),
    .B(net790),
    .A_N(_0141_));
 sg13g2_o21ai_1 _4129_ (.B1(_1166_),
    .Y(_1167_),
    .A1(net1719),
    .A2(net790));
 sg13g2_nand3b_1 _4130_ (.B(net1720),
    .C(net946),
    .Y(_1168_),
    .A_N(_0533_));
 sg13g2_o21ai_1 _4131_ (.B1(_1168_),
    .Y(_0037_),
    .A1(_0379_),
    .A2(net1720));
 sg13g2_or3_1 _4132_ (.A(_1162_),
    .B(_1165_),
    .C(_1167_),
    .X(_1169_));
 sg13g2_a21oi_1 _4133_ (.A1(_1162_),
    .A2(_1167_),
    .Y(_1170_),
    .B1(net1647));
 sg13g2_a22oi_1 _4134_ (.Y(_0038_),
    .B1(_1169_),
    .B2(net1721),
    .A2(_1163_),
    .A1(net1647));
 sg13g2_nor3_1 _4135_ (.A(_1161_),
    .B(_1162_),
    .C(_1167_),
    .Y(_1171_));
 sg13g2_nor2_1 _4136_ (.A(net1688),
    .B(net1757),
    .Y(_0039_));
 sg13g2_o21ai_1 _4137_ (.B1(\input_value_check_inst.character_buff[3][3] ),
    .Y(_1172_),
    .A1(\input_value_check_inst.character_buff[3][2] ),
    .A2(\input_value_check_inst.character_buff[3][1] ));
 sg13g2_nor2_1 _4138_ (.A(\input_value_check_inst.character_buff[3][7] ),
    .B(\input_value_check_inst.character_buff[3][6] ),
    .Y(_1173_));
 sg13g2_and4_1 _4139_ (.A(\input_value_check_inst.character_buff[3][5] ),
    .B(\input_value_check_inst.character_buff[3][4] ),
    .C(_1172_),
    .D(_1173_),
    .X(_1174_));
 sg13g2_nand4_1 _4140_ (.B(\input_value_check_inst.character_buff[3][4] ),
    .C(_1172_),
    .A(\input_value_check_inst.character_buff[3][5] ),
    .Y(_1175_),
    .D(_1173_));
 sg13g2_nand2b_1 _4141_ (.Y(_1176_),
    .B(\input_value_check_inst.character_buff[3][6] ),
    .A_N(\input_value_check_inst.character_buff[3][7] ));
 sg13g2_nor3_1 _4142_ (.A(\input_value_check_inst.character_buff[3][2] ),
    .B(\input_value_check_inst.character_buff[3][1] ),
    .C(\input_value_check_inst.character_buff[3][0] ),
    .Y(_1177_));
 sg13g2_nor4_1 _4143_ (.A(\input_value_check_inst.character_buff[3][4] ),
    .B(\input_value_check_inst.character_buff[3][3] ),
    .C(_1176_),
    .D(_1177_),
    .Y(_1178_));
 sg13g2_nand2b_1 _4144_ (.Y(_1179_),
    .B(_0137_),
    .A_N(\input_value_check_inst.character_buff[3][2] ));
 sg13g2_nand3_1 _4145_ (.B(\input_value_check_inst.character_buff[3][0] ),
    .C(_1175_),
    .A(\input_value_check_inst.character_buff[3][1] ),
    .Y(_1180_));
 sg13g2_nand3_1 _4146_ (.B(\input_value_check_inst.character_buff[3][0] ),
    .C(_1179_),
    .A(\input_value_check_inst.character_buff[3][1] ),
    .Y(_1181_));
 sg13g2_a21oi_1 _4147_ (.A1(_1178_),
    .A2(_1181_),
    .Y(_1182_),
    .B1(_1174_));
 sg13g2_and2_1 _4148_ (.A(_0138_),
    .B(_1174_),
    .X(_1183_));
 sg13g2_nor3_1 _4149_ (.A(net782),
    .B(_1182_),
    .C(_1183_),
    .Y(_1184_));
 sg13g2_a21oi_2 _4150_ (.B1(_1184_),
    .Y(_1185_),
    .A2(net783),
    .A1(net1618));
 sg13g2_nor2_2 _4151_ (.A(net894),
    .B(net1619),
    .Y(_0615_));
 sg13g2_a21oi_1 _4152_ (.A1(_0137_),
    .A2(_1180_),
    .Y(_1186_),
    .B1(_1182_));
 sg13g2_mux2_2 _4153_ (.A0(net1736),
    .A1(_1186_),
    .S(net795),
    .X(_1187_));
 sg13g2_nor2_1 _4154_ (.A(_0136_),
    .B(_1175_),
    .Y(_1188_));
 sg13g2_xnor2_1 _4155_ (.Y(_1189_),
    .A(\input_value_check_inst.character_buff[3][1] ),
    .B(\input_value_check_inst.character_buff[3][0] ));
 sg13g2_nor4_1 _4156_ (.A(\input_value_check_inst.character_buff[3][4] ),
    .B(\input_value_check_inst.character_buff[3][3] ),
    .C(_1176_),
    .D(_1189_),
    .Y(_1190_));
 sg13g2_o21ai_1 _4157_ (.B1(net795),
    .Y(_1191_),
    .A1(_1188_),
    .A2(_1190_));
 sg13g2_o21ai_1 _4158_ (.B1(_1191_),
    .Y(_1192_),
    .A1(_0143_),
    .A2(net795));
 sg13g2_or4_2 _4159_ (.A(net894),
    .B(_1185_),
    .C(_1187_),
    .D(_1192_),
    .X(_1193_));
 sg13g2_nand2_2 _4160_ (.Y(_1194_),
    .A(net938),
    .B(_1187_));
 sg13g2_inv_1 _4161_ (.Y(_0614_),
    .A(_1194_));
 sg13g2_nand2_1 _4162_ (.Y(_1195_),
    .A(_0846_),
    .B(_1178_));
 sg13g2_o21ai_1 _4163_ (.B1(_1195_),
    .Y(_1196_),
    .A1(_0135_),
    .A2(_1175_));
 sg13g2_nand2_1 _4164_ (.Y(_1197_),
    .A(net795),
    .B(_1196_));
 sg13g2_mux2_2 _4165_ (.A0(_0931_),
    .A1(_1196_),
    .S(net795),
    .X(_1198_));
 sg13g2_inv_1 _4166_ (.Y(_1199_),
    .A(_1198_));
 sg13g2_nand2_1 _4167_ (.Y(_1200_),
    .A(net938),
    .B(_1198_));
 sg13g2_or2_1 _4168_ (.X(_1201_),
    .B(_1200_),
    .A(_1192_));
 sg13g2_o21ai_1 _4169_ (.B1(_1194_),
    .Y(_1202_),
    .A1(_1192_),
    .A2(_1200_));
 sg13g2_nand2_1 _4170_ (.Y(_1203_),
    .A(net938),
    .B(_1192_));
 sg13g2_o21ai_1 _4171_ (.B1(net938),
    .Y(_1204_),
    .A1(_1192_),
    .A2(_1198_));
 sg13g2_inv_1 _4172_ (.Y(_1205_),
    .A(_1204_));
 sg13g2_a22oi_1 _4173_ (.Y(_1206_),
    .B1(_1205_),
    .B2(_1187_),
    .A2(_1201_),
    .A1(_1194_));
 sg13g2_o21ai_1 _4174_ (.B1(_1193_),
    .Y(_0021_),
    .A1(_0615_),
    .A2(_1206_));
 sg13g2_a21o_1 _4175_ (.A2(_1198_),
    .A1(_1192_),
    .B1(_1194_),
    .X(_1207_));
 sg13g2_nor2_1 _4176_ (.A(_1204_),
    .B(_1207_),
    .Y(_1208_));
 sg13g2_o21ai_1 _4177_ (.B1(_1193_),
    .Y(_0022_),
    .A1(_0615_),
    .A2(_1208_));
 sg13g2_nor3_1 _4178_ (.A(_1187_),
    .B(_1198_),
    .C(_1203_),
    .Y(_1209_));
 sg13g2_o21ai_1 _4179_ (.B1(_1193_),
    .Y(_0023_),
    .A1(_0615_),
    .A2(_1209_));
 sg13g2_o21ai_1 _4180_ (.B1(_1202_),
    .Y(_1210_),
    .A1(_1204_),
    .A2(_1207_));
 sg13g2_inv_1 _4181_ (.Y(_1211_),
    .A(_1210_));
 sg13g2_o21ai_1 _4182_ (.B1(_1193_),
    .Y(_0024_),
    .A1(_0615_),
    .A2(_1211_));
 sg13g2_nand2_1 _4183_ (.Y(_1212_),
    .A(_1194_),
    .B(_1204_));
 sg13g2_nand2_1 _4184_ (.Y(_1213_),
    .A(_1185_),
    .B(_1199_));
 sg13g2_o21ai_1 _4185_ (.B1(_1212_),
    .Y(_0025_),
    .A1(_1203_),
    .A2(_1213_));
 sg13g2_and2_1 _4186_ (.A(_1207_),
    .B(_1212_),
    .X(_1214_));
 sg13g2_o21ai_1 _4187_ (.B1(_1193_),
    .Y(_0026_),
    .A1(_0615_),
    .A2(_1214_));
 sg13g2_o21ai_1 _4188_ (.B1(_1207_),
    .Y(_1215_),
    .A1(_1187_),
    .A2(_1203_));
 sg13g2_inv_1 _4189_ (.Y(_1216_),
    .A(_1215_));
 sg13g2_o21ai_1 _4190_ (.B1(_1193_),
    .Y(_0027_),
    .A1(_0615_),
    .A2(_1216_));
 sg13g2_a21oi_1 _4191_ (.A1(net1690),
    .A2(net788),
    .Y(_1217_),
    .B1(net899));
 sg13g2_o21ai_1 _4192_ (.B1(_1217_),
    .Y(_1218_),
    .A1(_0932_),
    .A2(net788));
 sg13g2_mux2_1 _4193_ (.A0(\Led_Cycle_inst.genblk1[9].pwm_unit.pwm_out ),
    .A1(\output_value_inst.led_data_reg[9] ),
    .S(net789),
    .X(_1219_));
 sg13g2_nand2_1 _4194_ (.Y(_1220_),
    .A(net922),
    .B(net1755));
 sg13g2_inv_1 _4195_ (.Y(_0704_),
    .A(_1220_));
 sg13g2_a21oi_1 _4196_ (.A1(_0777_),
    .A2(net791),
    .Y(_1221_),
    .B1(net892));
 sg13g2_o21ai_1 _4197_ (.B1(_1221_),
    .Y(_1222_),
    .A1(net1782),
    .A2(net791));
 sg13g2_inv_1 _4198_ (.Y(_0705_),
    .A(net1754));
 sg13g2_a21oi_1 _4199_ (.A1(_1220_),
    .A2(_1222_),
    .Y(_0422_),
    .B1(_1218_));
 sg13g2_inv_1 _4200_ (.Y(_0376_),
    .A(_0422_));
 sg13g2_nand2b_1 _4201_ (.Y(_1223_),
    .B(net788),
    .A_N(net1741));
 sg13g2_o21ai_1 _4202_ (.B1(_1223_),
    .Y(_1224_),
    .A1(net1752),
    .A2(net788));
 sg13g2_nand3b_1 _4203_ (.B(net1742),
    .C(net922),
    .Y(_1225_),
    .A_N(_0422_));
 sg13g2_o21ai_1 _4204_ (.B1(_1225_),
    .Y(_0034_),
    .A1(_0376_),
    .A2(net1742));
 sg13g2_or3_1 _4205_ (.A(_1219_),
    .B(_1222_),
    .C(_1224_),
    .X(_1226_));
 sg13g2_a21oi_1 _4206_ (.A1(_1219_),
    .A2(_1224_),
    .Y(_1227_),
    .B1(_1218_));
 sg13g2_a22oi_1 _4207_ (.Y(_0035_),
    .B1(_1226_),
    .B2(_1227_),
    .A2(_1220_),
    .A1(_1218_));
 sg13g2_nor3_1 _4208_ (.A(_1218_),
    .B(_1219_),
    .C(net1742),
    .Y(_1228_));
 sg13g2_nor2_1 _4209_ (.A(net1754),
    .B(_1228_),
    .Y(_0036_));
 sg13g2_nor2_2 _4210_ (.A(\SegmentDisplay.out_sel[3] ),
    .B(net830),
    .Y(_1229_));
 sg13g2_nor3_2 _4211_ (.A(\SegmentDisplay.out_sel[3] ),
    .B(\SegmentDisplay.out_sel[0] ),
    .C(net830),
    .Y(_1230_));
 sg13g2_nand3_1 _4212_ (.B(\SegmentDisplay.digit1[3] ),
    .C(_1230_),
    .A(net828),
    .Y(_1231_));
 sg13g2_nor2_2 _4213_ (.A(\SegmentDisplay.out_sel[0] ),
    .B(net827),
    .Y(_1232_));
 sg13g2_nor2b_2 _4214_ (.A(net829),
    .B_N(\SegmentDisplay.out_sel[3] ),
    .Y(_1233_));
 sg13g2_nand3_1 _4215_ (.B(_1232_),
    .C(_1233_),
    .A(\SegmentDisplay.digit3[3] ),
    .Y(_1234_));
 sg13g2_nor3_2 _4216_ (.A(\SegmentDisplay.out_sel[3] ),
    .B(\SegmentDisplay.out_sel[0] ),
    .C(net827),
    .Y(_1235_));
 sg13g2_nand3_1 _4217_ (.B(\SegmentDisplay.digit2[3] ),
    .C(_1235_),
    .A(net830),
    .Y(_1236_));
 sg13g2_nor2b_2 _4218_ (.A(net828),
    .B_N(\SegmentDisplay.out_sel[0] ),
    .Y(_1237_));
 sg13g2_nand3_1 _4219_ (.B(_1229_),
    .C(_1237_),
    .A(\SegmentDisplay.digit0[3] ),
    .Y(_1238_));
 sg13g2_nand4_1 _4220_ (.B(_1234_),
    .C(_1236_),
    .A(_1231_),
    .Y(_1239_),
    .D(_1238_));
 sg13g2_nand3_1 _4221_ (.B(\SegmentDisplay.digit2[6] ),
    .C(_1235_),
    .A(net829),
    .Y(_1240_));
 sg13g2_nand3_1 _4222_ (.B(\SegmentDisplay.digit1[6] ),
    .C(_1230_),
    .A(net828),
    .Y(_1241_));
 sg13g2_nand3_1 _4223_ (.B(_1229_),
    .C(_1237_),
    .A(\SegmentDisplay.digit0[6] ),
    .Y(_1242_));
 sg13g2_nand3_1 _4224_ (.B(_1232_),
    .C(_1233_),
    .A(\SegmentDisplay.digit3[6] ),
    .Y(_1243_));
 sg13g2_nand4_1 _4225_ (.B(_1241_),
    .C(_1242_),
    .A(_1240_),
    .Y(_1244_),
    .D(_1243_));
 sg13g2_nand3_1 _4226_ (.B(\SegmentDisplay.digit1[2] ),
    .C(_1230_),
    .A(net827),
    .Y(_1245_));
 sg13g2_nand3_1 _4227_ (.B(_1229_),
    .C(_1237_),
    .A(\SegmentDisplay.digit0[2] ),
    .Y(_1246_));
 sg13g2_nand3_1 _4228_ (.B(\SegmentDisplay.digit2[2] ),
    .C(_1235_),
    .A(net829),
    .Y(_1247_));
 sg13g2_nand3_1 _4229_ (.B(_1232_),
    .C(_1233_),
    .A(\SegmentDisplay.digit3[2] ),
    .Y(_1248_));
 sg13g2_nand4_1 _4230_ (.B(_1246_),
    .C(_1247_),
    .A(_1245_),
    .Y(_1249_),
    .D(_1248_));
 sg13g2_nand3_1 _4231_ (.B(_1229_),
    .C(_1237_),
    .A(\SegmentDisplay.digit0[1] ),
    .Y(_1250_));
 sg13g2_nand3_1 _4232_ (.B(_1232_),
    .C(_1233_),
    .A(\SegmentDisplay.digit3[1] ),
    .Y(_1251_));
 sg13g2_nand3_1 _4233_ (.B(\SegmentDisplay.digit1[1] ),
    .C(_1230_),
    .A(net827),
    .Y(_1252_));
 sg13g2_nand3_1 _4234_ (.B(\SegmentDisplay.digit2[1] ),
    .C(_1235_),
    .A(net829),
    .Y(_1253_));
 sg13g2_nand4_1 _4235_ (.B(_1251_),
    .C(_1252_),
    .A(_1250_),
    .Y(_1254_),
    .D(_1253_));
 sg13g2_xnor2_1 _4236_ (.Y(_1255_),
    .A(_0100_),
    .B(_1254_));
 sg13g2_nand3_1 _4237_ (.B(_1232_),
    .C(_1233_),
    .A(\SegmentDisplay.digit3[0] ),
    .Y(_1256_));
 sg13g2_nand3_1 _4238_ (.B(\SegmentDisplay.digit1[0] ),
    .C(_1230_),
    .A(net827),
    .Y(_1257_));
 sg13g2_nand3_1 _4239_ (.B(\SegmentDisplay.digit2[0] ),
    .C(_1235_),
    .A(net829),
    .Y(_1258_));
 sg13g2_nand3_1 _4240_ (.B(_1229_),
    .C(_1237_),
    .A(\SegmentDisplay.digit0[0] ),
    .Y(_1259_));
 sg13g2_nand4_1 _4241_ (.B(_1257_),
    .C(_1258_),
    .A(_1256_),
    .Y(_1260_),
    .D(_1259_));
 sg13g2_nor2_1 _4242_ (.A(\output_value_inst.element_data_reg[10] ),
    .B(\SegmentDisplay.out_sel[3] ),
    .Y(_1261_));
 sg13g2_xnor2_1 _4243_ (.Y(_1262_),
    .A(uo_out[7]),
    .B(\output_value_inst.element_data_reg[11] ));
 sg13g2_nor2_1 _4244_ (.A(\output_value_inst.element_data_reg[7] ),
    .B(\SegmentDisplay.out_sel[0] ),
    .Y(_1263_));
 sg13g2_xnor2_1 _4245_ (.Y(_1264_),
    .A(\output_value_inst.element_data_reg[9] ),
    .B(net830));
 sg13g2_xor2_1 _4246_ (.B(net828),
    .A(\output_value_inst.element_data_reg[8] ),
    .X(_1265_));
 sg13g2_a22oi_1 _4247_ (.Y(_1266_),
    .B1(\SegmentDisplay.out_sel[0] ),
    .B2(\output_value_inst.element_data_reg[7] ),
    .A2(\SegmentDisplay.out_sel[3] ),
    .A1(\output_value_inst.element_data_reg[10] ));
 sg13g2_nor3_1 _4248_ (.A(_1261_),
    .B(_1263_),
    .C(_1264_),
    .Y(_1267_));
 sg13g2_nand4_1 _4249_ (.B(_1265_),
    .C(_1266_),
    .A(_1262_),
    .Y(_1268_),
    .D(_1267_));
 sg13g2_nand3_1 _4250_ (.B(\SegmentDisplay.digit1[5] ),
    .C(_1230_),
    .A(net827),
    .Y(_1269_));
 sg13g2_nand3_1 _4251_ (.B(_1229_),
    .C(_1237_),
    .A(\SegmentDisplay.digit0[5] ),
    .Y(_1270_));
 sg13g2_nand3_1 _4252_ (.B(\SegmentDisplay.digit2[5] ),
    .C(_1235_),
    .A(net829),
    .Y(_1271_));
 sg13g2_nand3_1 _4253_ (.B(_1232_),
    .C(_1233_),
    .A(\SegmentDisplay.digit3[5] ),
    .Y(_1272_));
 sg13g2_nand4_1 _4254_ (.B(_1270_),
    .C(_1271_),
    .A(_1269_),
    .Y(_1273_),
    .D(_1272_));
 sg13g2_nand3_1 _4255_ (.B(\SegmentDisplay.digit1[4] ),
    .C(_1230_),
    .A(net827),
    .Y(_1274_));
 sg13g2_nand3_1 _4256_ (.B(_1229_),
    .C(_1237_),
    .A(\SegmentDisplay.digit0[4] ),
    .Y(_1275_));
 sg13g2_nand3_1 _4257_ (.B(_1232_),
    .C(_1233_),
    .A(\SegmentDisplay.digit3[4] ),
    .Y(_1276_));
 sg13g2_nand3_1 _4258_ (.B(\SegmentDisplay.digit2[4] ),
    .C(_1235_),
    .A(net829),
    .Y(_1277_));
 sg13g2_nand4_1 _4259_ (.B(_1275_),
    .C(_1276_),
    .A(_1274_),
    .Y(_1278_),
    .D(_1277_));
 sg13g2_nor2_1 _4260_ (.A(_0912_),
    .B(_1278_),
    .Y(_1279_));
 sg13g2_xnor2_1 _4261_ (.Y(_1280_),
    .A(_0101_),
    .B(_1249_));
 sg13g2_xnor2_1 _4262_ (.Y(_1281_),
    .A(_0792_),
    .B(_1260_));
 sg13g2_a21oi_1 _4263_ (.A1(_0912_),
    .A2(_1278_),
    .Y(_1282_),
    .B1(_1268_));
 sg13g2_xor2_1 _4264_ (.B(_1239_),
    .A(_0102_),
    .X(_1283_));
 sg13g2_xor2_1 _4265_ (.B(_1244_),
    .A(_0105_),
    .X(_1284_));
 sg13g2_xor2_1 _4266_ (.B(_1273_),
    .A(_0104_),
    .X(_1285_));
 sg13g2_and4_1 _4267_ (.A(_1255_),
    .B(_1280_),
    .C(_1281_),
    .D(_1282_),
    .X(_1286_));
 sg13g2_nor4_1 _4268_ (.A(_1279_),
    .B(_1283_),
    .C(_1284_),
    .D(_1285_),
    .Y(_1287_));
 sg13g2_a21oi_1 _4269_ (.A1(_1286_),
    .A2(_1287_),
    .Y(_1288_),
    .B1(net914));
 sg13g2_nand2b_1 _4270_ (.Y(_1289_),
    .B(net1242),
    .A_N(net732));
 sg13g2_nand2_1 _4271_ (.Y(_1290_),
    .A(\SegmentDisplay.out_sel[0] ),
    .B(net730));
 sg13g2_and3_1 _4272_ (.X(_1291_),
    .A(net951),
    .B(_1289_),
    .C(_1290_));
 sg13g2_nand3_1 _4273_ (.B(_1289_),
    .C(_1290_),
    .A(net951),
    .Y(_1292_));
 sg13g2_nand2b_1 _4274_ (.Y(_1293_),
    .B(net733),
    .A_N(_1273_));
 sg13g2_mux2_1 _4275_ (.A0(_0104_),
    .A1(_1273_),
    .S(net732),
    .X(_1294_));
 sg13g2_nor2_1 _4276_ (.A(net895),
    .B(_1294_),
    .Y(_1295_));
 sg13g2_nand2b_1 _4277_ (.Y(_1296_),
    .B(net732),
    .A_N(_1244_));
 sg13g2_or2_1 _4278_ (.X(_1297_),
    .B(net732),
    .A(net1712));
 sg13g2_a21oi_2 _4279_ (.B1(net895),
    .Y(_1298_),
    .A2(_1297_),
    .A1(_1296_));
 sg13g2_o21ai_1 _4280_ (.B1(_1291_),
    .Y(_0375_),
    .A1(_1295_),
    .A2(_1298_));
 sg13g2_inv_1 _4281_ (.Y(_0544_),
    .A(_0375_));
 sg13g2_nand2b_1 _4282_ (.Y(_1299_),
    .B(net732),
    .A_N(_1278_));
 sg13g2_mux2_1 _4283_ (.A0(net1743),
    .A1(_1278_),
    .S(net732),
    .X(_1300_));
 sg13g2_nor2_1 _4284_ (.A(net895),
    .B(_1300_),
    .Y(_1301_));
 sg13g2_mux2_1 _4285_ (.A0(_1300_),
    .A1(_1301_),
    .S(_0375_),
    .X(_0043_));
 sg13g2_and3_1 _4286_ (.X(_1302_),
    .A(_1291_),
    .B(_1294_),
    .C(_1300_));
 sg13g2_nor2_1 _4287_ (.A(_1294_),
    .B(_1300_),
    .Y(_1303_));
 sg13g2_mux2_1 _4288_ (.A0(_1295_),
    .A1(_1303_),
    .S(_1291_),
    .X(_1304_));
 sg13g2_a21o_1 _4289_ (.A2(_1302_),
    .A1(_1298_),
    .B1(_1304_),
    .X(_0044_));
 sg13g2_nor2b_1 _4290_ (.A(_1302_),
    .B_N(_1298_),
    .Y(_0045_));
 sg13g2_a21oi_1 _4291_ (.A1(net1765),
    .A2(net731),
    .Y(_1305_),
    .B1(net897));
 sg13g2_o21ai_1 _4292_ (.B1(_1305_),
    .Y(_1306_),
    .A1(_0933_),
    .A2(net731));
 sg13g2_mux2_1 _4293_ (.A0(net1758),
    .A1(\SegmentDisplay.an[2] ),
    .S(net730),
    .X(_1307_));
 sg13g2_nand2_2 _4294_ (.Y(_1308_),
    .A(net939),
    .B(_1307_));
 sg13g2_inv_1 _4295_ (.Y(_0692_),
    .A(_1308_));
 sg13g2_a21oi_1 _4296_ (.A1(_0789_),
    .A2(net730),
    .Y(_1309_),
    .B1(net895));
 sg13g2_o21ai_1 _4297_ (.B1(_1309_),
    .Y(_1310_),
    .A1(net1767),
    .A2(net730));
 sg13g2_inv_1 _4298_ (.Y(_0693_),
    .A(_1310_));
 sg13g2_a21oi_2 _4299_ (.B1(_1306_),
    .Y(_0535_),
    .A2(_1310_),
    .A1(_1308_));
 sg13g2_inv_1 _4300_ (.Y(_0373_),
    .A(_0535_));
 sg13g2_mux2_2 _4301_ (.A0(_0934_),
    .A1(_0906_),
    .S(net730),
    .X(_1311_));
 sg13g2_inv_1 _4302_ (.Y(_1312_),
    .A(_1311_));
 sg13g2_nor2_1 _4303_ (.A(_1306_),
    .B(_1311_),
    .Y(_1313_));
 sg13g2_nor2_1 _4304_ (.A(net895),
    .B(_1312_),
    .Y(_1314_));
 sg13g2_mux2_1 _4305_ (.A0(_1314_),
    .A1(_1312_),
    .S(_0535_),
    .X(_0046_));
 sg13g2_or3_1 _4306_ (.A(_1307_),
    .B(_1310_),
    .C(_1311_),
    .X(_1315_));
 sg13g2_a21oi_1 _4307_ (.A1(_1307_),
    .A2(_1311_),
    .Y(_1316_),
    .B1(_1306_));
 sg13g2_a22oi_1 _4308_ (.Y(_0047_),
    .B1(_1315_),
    .B2(_1316_),
    .A2(_1308_),
    .A1(_1306_));
 sg13g2_a21oi_1 _4309_ (.A1(_1308_),
    .A2(_1313_),
    .Y(_0048_),
    .B1(_1310_));
 sg13g2_o21ai_1 _4310_ (.B1(net941),
    .Y(_1317_),
    .A1(uo_out[3]),
    .A2(net796));
 sg13g2_o21ai_1 _4311_ (.B1(\input_value_check_inst.character_buff[0][3] ),
    .Y(_1318_),
    .A1(\input_value_check_inst.character_buff[0][2] ),
    .A2(\input_value_check_inst.character_buff[0][1] ));
 sg13g2_nor2_1 _4312_ (.A(\input_value_check_inst.character_buff[0][7] ),
    .B(\input_value_check_inst.character_buff[0][6] ),
    .Y(_1319_));
 sg13g2_nand4_1 _4313_ (.B(\input_value_check_inst.character_buff[0][4] ),
    .C(_1318_),
    .A(\input_value_check_inst.character_buff[0][5] ),
    .Y(_1320_),
    .D(_1319_));
 sg13g2_nand2_1 _4314_ (.Y(_1321_),
    .A(\input_value_check_inst.character_buff[0][1] ),
    .B(\input_value_check_inst.character_buff[0][0] ));
 sg13g2_nand3_1 _4315_ (.B(\input_value_check_inst.character_buff[0][1] ),
    .C(\input_value_check_inst.character_buff[0][0] ),
    .A(\input_value_check_inst.character_buff[0][2] ),
    .Y(_1322_));
 sg13g2_nor2b_1 _4316_ (.A(\input_value_check_inst.character_buff[0][7] ),
    .B_N(\input_value_check_inst.character_buff[0][6] ),
    .Y(_1323_));
 sg13g2_nor2_1 _4317_ (.A(\input_value_check_inst.character_buff[0][4] ),
    .B(\input_value_check_inst.character_buff[0][3] ),
    .Y(_1324_));
 sg13g2_nand2_1 _4318_ (.Y(_1325_),
    .A(_0829_),
    .B(_0831_));
 sg13g2_or3_1 _4319_ (.A(\input_value_check_inst.character_buff[0][2] ),
    .B(\input_value_check_inst.character_buff[0][1] ),
    .C(\input_value_check_inst.character_buff[0][0] ),
    .X(_1326_));
 sg13g2_nand4_1 _4320_ (.B(_1323_),
    .C(_1324_),
    .A(_1322_),
    .Y(_1327_),
    .D(_1326_));
 sg13g2_nor2b_1 _4321_ (.A(_1321_),
    .B_N(_1320_),
    .Y(_1328_));
 sg13g2_a22oi_1 _4322_ (.Y(_1329_),
    .B1(_1328_),
    .B2(_0937_),
    .A2(_1327_),
    .A1(_1320_));
 sg13g2_o21ai_1 _4323_ (.B1(_1329_),
    .Y(_1330_),
    .A1(_0938_),
    .A2(_1320_));
 sg13g2_a21oi_1 _4324_ (.A1(net796),
    .A2(_1330_),
    .Y(_0603_),
    .B1(_1317_));
 sg13g2_o21ai_1 _4325_ (.B1(_1329_),
    .Y(_1331_),
    .A1(_0937_),
    .A2(_1328_));
 sg13g2_o21ai_1 _4326_ (.B1(net940),
    .Y(_1332_),
    .A1(net1737),
    .A2(net796));
 sg13g2_a21oi_2 _4327_ (.B1(_1332_),
    .Y(_0602_),
    .A2(_1331_),
    .A1(net797));
 sg13g2_inv_1 _4328_ (.Y(_1333_),
    .A(_0602_));
 sg13g2_nand4_1 _4329_ (.B(_1323_),
    .C(_1324_),
    .A(_1321_),
    .Y(_1334_),
    .D(_1325_));
 sg13g2_o21ai_1 _4330_ (.B1(_1334_),
    .Y(_1335_),
    .A1(_0154_),
    .A2(_1320_));
 sg13g2_nand2_1 _4331_ (.Y(_1336_),
    .A(net797),
    .B(_1335_));
 sg13g2_mux2_1 _4332_ (.A0(_0935_),
    .A1(_1335_),
    .S(net796),
    .X(_1337_));
 sg13g2_nand2_2 _4333_ (.Y(_1338_),
    .A(net942),
    .B(_1337_));
 sg13g2_nand3_1 _4334_ (.B(_1333_),
    .C(_1338_),
    .A(_0603_),
    .Y(_1339_));
 sg13g2_nand2b_1 _4335_ (.Y(_1340_),
    .B(_0831_),
    .A_N(_1327_));
 sg13g2_o21ai_1 _4336_ (.B1(_1340_),
    .Y(_1341_),
    .A1(_0156_),
    .A2(_1320_));
 sg13g2_nand2_1 _4337_ (.Y(_1342_),
    .A(net797),
    .B(_1341_));
 sg13g2_mux2_1 _4338_ (.A0(_0936_),
    .A1(_1341_),
    .S(net796),
    .X(_1343_));
 sg13g2_nand2_1 _4339_ (.Y(_1344_),
    .A(net941),
    .B(_1343_));
 sg13g2_o21ai_1 _4340_ (.B1(_1333_),
    .Y(_1345_),
    .A1(_1337_),
    .A2(_1344_));
 sg13g2_nand2_1 _4341_ (.Y(_1346_),
    .A(_1338_),
    .B(_1344_));
 sg13g2_nand2_1 _4342_ (.Y(_1347_),
    .A(_0602_),
    .B(_1346_));
 sg13g2_and2_1 _4343_ (.A(_1345_),
    .B(_1347_),
    .X(_1348_));
 sg13g2_o21ai_1 _4344_ (.B1(_1339_),
    .Y(_0000_),
    .A1(net755),
    .A2(_1348_));
 sg13g2_nand3_1 _4345_ (.B(_1337_),
    .C(_1343_),
    .A(net940),
    .Y(_1349_));
 sg13g2_and2_1 _4346_ (.A(_0602_),
    .B(_1349_),
    .X(_1350_));
 sg13g2_and2_1 _4347_ (.A(_1346_),
    .B(_1350_),
    .X(_1351_));
 sg13g2_nand2_1 _4348_ (.Y(_1352_),
    .A(_1346_),
    .B(_1350_));
 sg13g2_o21ai_1 _4349_ (.B1(_1339_),
    .Y(_0001_),
    .A1(net755),
    .A2(_1351_));
 sg13g2_nor2_1 _4350_ (.A(_0602_),
    .B(_1338_),
    .Y(_1353_));
 sg13g2_nor3_1 _4351_ (.A(_0602_),
    .B(_1338_),
    .C(_1343_),
    .Y(_1354_));
 sg13g2_o21ai_1 _4352_ (.B1(_1339_),
    .Y(_0002_),
    .A1(net755),
    .A2(_1354_));
 sg13g2_and2_1 _4353_ (.A(_1345_),
    .B(_1352_),
    .X(_1355_));
 sg13g2_o21ai_1 _4354_ (.B1(_1339_),
    .Y(_0003_),
    .A1(net755),
    .A2(_1355_));
 sg13g2_or3_1 _4355_ (.A(net755),
    .B(_1338_),
    .C(_1343_),
    .X(_1356_));
 sg13g2_o21ai_1 _4356_ (.B1(_1356_),
    .Y(_0004_),
    .A1(_0602_),
    .A2(_1346_));
 sg13g2_a21oi_1 _4357_ (.A1(_1338_),
    .A2(_1344_),
    .Y(_1357_),
    .B1(_1350_));
 sg13g2_o21ai_1 _4358_ (.B1(_1339_),
    .Y(_0005_),
    .A1(net755),
    .A2(_1357_));
 sg13g2_nor2_1 _4359_ (.A(_1350_),
    .B(_1353_),
    .Y(_1358_));
 sg13g2_o21ai_1 _4360_ (.B1(_1339_),
    .Y(_0006_),
    .A1(net755),
    .A2(_1358_));
 sg13g2_a21oi_1 _4361_ (.A1(net1707),
    .A2(net789),
    .Y(_1359_),
    .B1(net892));
 sg13g2_o21ai_1 _4362_ (.B1(_1359_),
    .Y(_1360_),
    .A1(_0939_),
    .A2(net789));
 sg13g2_mux2_2 _4363_ (.A0(\Led_Cycle_inst.genblk1[5].pwm_unit.pwm_out ),
    .A1(net1675),
    .S(net790),
    .X(_1361_));
 sg13g2_nand2_1 _4364_ (.Y(_1362_),
    .A(net946),
    .B(net1676));
 sg13g2_inv_1 _4365_ (.Y(_0700_),
    .A(_1362_));
 sg13g2_a21oi_1 _4366_ (.A1(_0780_),
    .A2(net790),
    .Y(_1363_),
    .B1(net900));
 sg13g2_o21ai_1 _4367_ (.B1(_1363_),
    .Y(_1364_),
    .A1(\Led_Cycle_inst.genblk1[6].pwm_unit.pwm_out ),
    .A2(net791));
 sg13g2_inv_1 _4368_ (.Y(_0701_),
    .A(net1749));
 sg13g2_a21oi_1 _4369_ (.A1(_1362_),
    .A2(_1364_),
    .Y(_0372_),
    .B1(_1360_));
 sg13g2_inv_1 _4370_ (.Y(_0377_),
    .A(net1709));
 sg13g2_nand2b_1 _4371_ (.Y(_1365_),
    .B(net791),
    .A_N(_0162_));
 sg13g2_o21ai_1 _4372_ (.B1(_1365_),
    .Y(_1366_),
    .A1(net1728),
    .A2(net790));
 sg13g2_nand3b_1 _4373_ (.B(net1729),
    .C(net951),
    .Y(_1367_),
    .A_N(_0372_));
 sg13g2_o21ai_1 _4374_ (.B1(_1367_),
    .Y(_0031_),
    .A1(_0377_),
    .A2(net1729));
 sg13g2_or3_1 _4375_ (.A(_1361_),
    .B(_1364_),
    .C(_1366_),
    .X(_1368_));
 sg13g2_a21oi_1 _4376_ (.A1(_1361_),
    .A2(_1366_),
    .Y(_1369_),
    .B1(net1708));
 sg13g2_a22oi_1 _4377_ (.Y(_0032_),
    .B1(_1368_),
    .B2(net1730),
    .A2(_1362_),
    .A1(net1708));
 sg13g2_nor3_1 _4378_ (.A(_1360_),
    .B(_1361_),
    .C(_1366_),
    .Y(_1370_));
 sg13g2_nor2_1 _4379_ (.A(net1749),
    .B(_1370_),
    .Y(_0033_));
 sg13g2_nand2b_1 _4380_ (.Y(_1371_),
    .B(net734),
    .A_N(_1239_));
 sg13g2_mux2_1 _4381_ (.A0(net1733),
    .A1(_1239_),
    .S(net734),
    .X(_1372_));
 sg13g2_o21ai_1 _4382_ (.B1(_1371_),
    .Y(_1373_),
    .A1(net1733),
    .A2(net734));
 sg13g2_nand2b_1 _4383_ (.Y(_1374_),
    .B(net735),
    .A_N(_1254_));
 sg13g2_mux2_1 _4384_ (.A0(_0100_),
    .A1(_1254_),
    .S(net734),
    .X(_1375_));
 sg13g2_nand2b_1 _4385_ (.Y(_1376_),
    .B(net951),
    .A_N(_1375_));
 sg13g2_nand2b_1 _4386_ (.Y(_1377_),
    .B(net735),
    .A_N(_1249_));
 sg13g2_or2_1 _4387_ (.X(_1378_),
    .B(net735),
    .A(net1738));
 sg13g2_a21o_1 _4388_ (.A2(_1378_),
    .A1(_1377_),
    .B1(net906),
    .X(_1379_));
 sg13g2_a21o_1 _4389_ (.A2(_1379_),
    .A1(_1376_),
    .B1(_1372_),
    .X(_0374_));
 sg13g2_inv_1 _4390_ (.Y(_0519_),
    .A(_0374_));
 sg13g2_mux2_1 _4391_ (.A0(net1686),
    .A1(_1260_),
    .S(net734),
    .X(_1380_));
 sg13g2_nor2_1 _4392_ (.A(net906),
    .B(_1380_),
    .Y(_1381_));
 sg13g2_mux2_1 _4393_ (.A0(_1380_),
    .A1(_1381_),
    .S(_0374_),
    .X(_0040_));
 sg13g2_nor2_1 _4394_ (.A(net906),
    .B(_1372_),
    .Y(_1382_));
 sg13g2_nand2_1 _4395_ (.Y(_1383_),
    .A(_1375_),
    .B(_1380_));
 sg13g2_or2_1 _4396_ (.X(_1384_),
    .B(_1380_),
    .A(_1375_));
 sg13g2_o21ai_1 _4397_ (.B1(_1384_),
    .Y(_1385_),
    .A1(_1379_),
    .A2(_1383_));
 sg13g2_nor2_1 _4398_ (.A(_1373_),
    .B(_1376_),
    .Y(_1386_));
 sg13g2_a21o_1 _4399_ (.A2(_1385_),
    .A1(_1382_),
    .B1(_1386_),
    .X(_0041_));
 sg13g2_nor2_1 _4400_ (.A(_1372_),
    .B(_1383_),
    .Y(_1387_));
 sg13g2_nor2_1 _4401_ (.A(_1379_),
    .B(_1387_),
    .Y(_0042_));
 sg13g2_o21ai_1 _4402_ (.B1(_1045_),
    .Y(_1388_),
    .A1(_1063_),
    .A2(_1068_));
 sg13g2_nand2_1 _4403_ (.Y(_0007_),
    .A(_1054_),
    .B(_1388_));
 sg13g2_nor2_1 _4404_ (.A(\uart_tx_fifo_inst.fifo_valid[3] ),
    .B(\uart_tx_fifo_inst.fifo_valid[2] ),
    .Y(_1389_));
 sg13g2_nor2_2 _4405_ (.A(\uart_tx_fifo_inst.fifo_valid[1] ),
    .B(\uart_tx_fifo_inst.fifo_valid[0] ),
    .Y(_1390_));
 sg13g2_nand2_1 _4406_ (.Y(_1391_),
    .A(_1389_),
    .B(_1390_));
 sg13g2_nor2_1 _4407_ (.A(\uart_tx_fifo_inst.fifo_valid[7] ),
    .B(\uart_tx_fifo_inst.fifo_valid[6] ),
    .Y(_1392_));
 sg13g2_nor3_1 _4408_ (.A(\uart_tx_fifo_inst.fifo_valid[7] ),
    .B(\uart_tx_fifo_inst.fifo_valid[6] ),
    .C(\uart_tx_fifo_inst.fifo_valid[5] ),
    .Y(_1393_));
 sg13g2_nand4_1 _4409_ (.B(_1389_),
    .C(_1390_),
    .A(_0818_),
    .Y(_1394_),
    .D(_1393_));
 sg13g2_nor2_1 _4410_ (.A(\uart_tx_fifo_inst.fifo_valid[9] ),
    .B(\uart_tx_fifo_inst.fifo_valid[8] ),
    .Y(_1395_));
 sg13g2_nand2b_1 _4411_ (.Y(_1396_),
    .B(_1395_),
    .A_N(_1394_));
 sg13g2_nand2_2 _4412_ (.Y(_1397_),
    .A(net962),
    .B(_1396_));
 sg13g2_nor2_1 _4413_ (.A(_0159_),
    .B(_1397_),
    .Y(_1398_));
 sg13g2_nor2_1 _4414_ (.A(net911),
    .B(_1398_),
    .Y(_1399_));
 sg13g2_nor3_1 _4415_ (.A(net911),
    .B(_0159_),
    .C(_1397_),
    .Y(_1400_));
 sg13g2_a22oi_1 _4416_ (.Y(_1401_),
    .B1(net779),
    .B2(net1287),
    .A2(net752),
    .A1(\uart_tx_fifo_inst.fifo[8][0] ));
 sg13g2_nand2b_1 _4417_ (.Y(_1402_),
    .B(\uart_tx_fifo_inst.fifo_valid[9] ),
    .A_N(\uart_tx_fifo_inst.fifo_valid[8] ));
 sg13g2_a21oi_1 _4418_ (.A1(_0816_),
    .A2(_1402_),
    .Y(_1403_),
    .B1(\uart_tx_fifo_inst.fifo_valid[6] ));
 sg13g2_o21ai_1 _4419_ (.B1(_0818_),
    .Y(_1404_),
    .A1(\uart_tx_fifo_inst.fifo_valid[5] ),
    .A2(_1403_));
 sg13g2_a21oi_2 _4420_ (.B1(\uart_tx_fifo_inst.fifo_valid[2] ),
    .Y(_1405_),
    .A2(_1404_),
    .A1(_0819_));
 sg13g2_nor2_1 _4421_ (.A(\uart_tx_fifo_inst.fifo_valid[1] ),
    .B(_1405_),
    .Y(_1406_));
 sg13g2_nor2_2 _4422_ (.A(\uart_tx_fifo_inst.fifo_valid[0] ),
    .B(_1406_),
    .Y(_1407_));
 sg13g2_o21ai_1 _4423_ (.B1(_0821_),
    .Y(_1408_),
    .A1(\uart_tx_fifo_inst.fifo_valid[1] ),
    .A2(_1405_));
 sg13g2_nand2_1 _4424_ (.Y(_1409_),
    .A(_0817_),
    .B(_0121_));
 sg13g2_o21ai_1 _4425_ (.B1(_1389_),
    .Y(_1410_),
    .A1(_1392_),
    .A2(_1409_));
 sg13g2_and2_1 _4426_ (.A(_1390_),
    .B(_1410_),
    .X(_1411_));
 sg13g2_nand2_1 _4427_ (.Y(_1412_),
    .A(_1390_),
    .B(_1410_));
 sg13g2_and2_1 _4428_ (.A(net770),
    .B(_1412_),
    .X(_1413_));
 sg13g2_nand2_2 _4429_ (.Y(_1414_),
    .A(net770),
    .B(_1412_));
 sg13g2_nor2_1 _4430_ (.A(net914),
    .B(_0876_),
    .Y(_1415_));
 sg13g2_nand2_1 _4431_ (.Y(_1416_),
    .A(net962),
    .B(net889));
 sg13g2_nor2_1 _4432_ (.A(_0876_),
    .B(_1397_),
    .Y(_1417_));
 sg13g2_nand2_1 _4433_ (.Y(_1418_),
    .A(net959),
    .B(_1417_));
 sg13g2_or2_1 _4434_ (.X(_1419_),
    .B(_1395_),
    .A(_1394_));
 sg13g2_a21oi_2 _4435_ (.B1(_1391_),
    .Y(_1420_),
    .A2(_1393_),
    .A1(_0121_));
 sg13g2_inv_1 _4436_ (.Y(_1421_),
    .A(_1420_));
 sg13g2_nor2_2 _4437_ (.A(_1419_),
    .B(_1420_),
    .Y(_1422_));
 sg13g2_nand3_1 _4438_ (.B(_1417_),
    .C(_1422_),
    .A(net959),
    .Y(_1423_));
 sg13g2_nor2_2 _4439_ (.A(_1414_),
    .B(_1423_),
    .Y(_1424_));
 sg13g2_nor2_1 _4440_ (.A(net1288),
    .B(_1424_),
    .Y(_0225_));
 sg13g2_a22oi_1 _4441_ (.Y(_1425_),
    .B1(net779),
    .B2(net1112),
    .A2(net752),
    .A1(\uart_tx_fifo_inst.fifo[8][1] ));
 sg13g2_nor2_1 _4442_ (.A(_1424_),
    .B(net1113),
    .Y(_0226_));
 sg13g2_a22oi_1 _4443_ (.Y(_1426_),
    .B1(net774),
    .B2(\uart_tx_fifo_inst.fifo[7][2] ),
    .A2(net747),
    .A1(net1357));
 sg13g2_nor2_1 _4444_ (.A(_1424_),
    .B(net1358),
    .Y(_0227_));
 sg13g2_a22oi_1 _4445_ (.Y(_1427_),
    .B1(net773),
    .B2(net695),
    .A2(net746),
    .A1(\uart_tx_fifo_inst.fifo[8][3] ));
 sg13g2_nor2_1 _4446_ (.A(_1424_),
    .B(net696),
    .Y(_0228_));
 sg13g2_a22oi_1 _4447_ (.Y(_1428_),
    .B1(net780),
    .B2(net1098),
    .A2(net753),
    .A1(\uart_tx_fifo_inst.fifo[8][4] ));
 sg13g2_nor2_1 _4448_ (.A(_1424_),
    .B(net1099),
    .Y(_0229_));
 sg13g2_a22oi_1 _4449_ (.Y(_1429_),
    .B1(net773),
    .B2(net1328),
    .A2(net746),
    .A1(\uart_tx_fifo_inst.fifo[8][5] ));
 sg13g2_nor2_1 _4450_ (.A(_1424_),
    .B(net1329),
    .Y(_0230_));
 sg13g2_a22oi_1 _4451_ (.Y(_1430_),
    .B1(net778),
    .B2(net1018),
    .A2(net751),
    .A1(\uart_tx_fifo_inst.fifo[8][6] ));
 sg13g2_nor2_1 _4452_ (.A(_1424_),
    .B(net1019),
    .Y(_0231_));
 sg13g2_and3_1 _4453_ (.X(_1431_),
    .A(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[0] ),
    .B(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[1] ),
    .C(net1161));
 sg13g2_and2_1 _4454_ (.A(net1491),
    .B(_1431_),
    .X(_1432_));
 sg13g2_nand2_1 _4455_ (.Y(_1433_),
    .A(net1715),
    .B(_1432_));
 sg13g2_o21ai_1 _4456_ (.B1(net946),
    .Y(_1434_),
    .A1(_0916_),
    .A2(_1433_));
 sg13g2_nor2_1 _4457_ (.A(_0953_),
    .B(_1434_),
    .Y(_0232_));
 sg13g2_xnor2_1 _4458_ (.Y(_1435_),
    .A(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[0] ),
    .B(net1557));
 sg13g2_nor2_1 _4459_ (.A(_1434_),
    .B(net1558),
    .Y(_0233_));
 sg13g2_a21oi_1 _4460_ (.A1(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[0] ),
    .A2(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[1] ),
    .Y(_1436_),
    .B1(net1161));
 sg13g2_nor3_1 _4461_ (.A(net900),
    .B(_1431_),
    .C(net1162),
    .Y(_0234_));
 sg13g2_o21ai_1 _4462_ (.B1(net945),
    .Y(_1437_),
    .A1(net1491),
    .A2(_1431_));
 sg13g2_nor2_1 _4463_ (.A(_1432_),
    .B(net1492),
    .Y(_0235_));
 sg13g2_or2_1 _4464_ (.X(_1438_),
    .B(_1432_),
    .A(net1715));
 sg13g2_and3_1 _4465_ (.X(_0236_),
    .A(net945),
    .B(_1433_),
    .C(_1438_));
 sg13g2_a21oi_1 _4466_ (.A1(_0916_),
    .A2(_1433_),
    .Y(_0237_),
    .B1(_1434_));
 sg13g2_nand2_1 _4467_ (.Y(_1439_),
    .A(net834),
    .B(_0963_));
 sg13g2_xnor2_1 _4468_ (.Y(_1440_),
    .A(_0940_),
    .B(_1439_));
 sg13g2_nor2_1 _4469_ (.A(_0967_),
    .B(_1440_),
    .Y(_1441_));
 sg13g2_and2_1 _4470_ (.A(_0967_),
    .B(_1440_),
    .X(_1442_));
 sg13g2_nor3_2 _4471_ (.A(_0966_),
    .B(_1441_),
    .C(_1442_),
    .Y(_1443_));
 sg13g2_nand2b_1 _4472_ (.Y(_1444_),
    .B(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[4] ),
    .A_N(_0200_));
 sg13g2_nor2_1 _4473_ (.A(_0896_),
    .B(net826),
    .Y(_1445_));
 sg13g2_nand2_1 _4474_ (.Y(_1446_),
    .A(net837),
    .B(net833));
 sg13g2_nor2_2 _4475_ (.A(net837),
    .B(net826),
    .Y(_1447_));
 sg13g2_nand2_1 _4476_ (.Y(_1448_),
    .A(_0896_),
    .B(net832));
 sg13g2_a21oi_1 _4477_ (.A1(net837),
    .A2(net840),
    .Y(_1449_),
    .B1(net826));
 sg13g2_o21ai_1 _4478_ (.B1(_1449_),
    .Y(_1450_),
    .A1(net840),
    .A2(_1448_));
 sg13g2_nor2_1 _4479_ (.A(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[2] ),
    .B(_1450_),
    .Y(_1451_));
 sg13g2_o21ai_1 _4480_ (.B1(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[1] ),
    .Y(_1452_),
    .A1(net609),
    .A2(_0210_));
 sg13g2_nor2_2 _4481_ (.A(net838),
    .B(net840),
    .Y(_1453_));
 sg13g2_or2_2 _4482_ (.X(_1454_),
    .B(net841),
    .A(net839));
 sg13g2_nand2_1 _4483_ (.Y(_1455_),
    .A(_0962_),
    .B(_1445_));
 sg13g2_o21ai_1 _4484_ (.B1(_1455_),
    .Y(_1456_),
    .A1(_1448_),
    .A2(_1454_));
 sg13g2_nand2_1 _4485_ (.Y(_1457_),
    .A(net836),
    .B(_1453_));
 sg13g2_nor2_2 _4486_ (.A(_1446_),
    .B(_1454_),
    .Y(_1458_));
 sg13g2_a21oi_2 _4487_ (.B1(_1458_),
    .Y(_1459_),
    .A2(_1447_),
    .A1(_0962_));
 sg13g2_inv_1 _4488_ (.Y(_1460_),
    .A(_1459_));
 sg13g2_nor3_1 _4489_ (.A(net609),
    .B(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[1] ),
    .C(_0210_),
    .Y(_1461_));
 sg13g2_o21ai_1 _4490_ (.B1(_1452_),
    .Y(_1462_),
    .A1(_1456_),
    .A2(_1461_));
 sg13g2_nand2_1 _4491_ (.Y(_1463_),
    .A(_1459_),
    .B(_1462_));
 sg13g2_nor2b_1 _4492_ (.A(_0210_),
    .B_N(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[1] ),
    .Y(_1464_));
 sg13g2_a22oi_1 _4493_ (.Y(_1465_),
    .B1(_1460_),
    .B2(_1464_),
    .A2(_1450_),
    .A1(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[2] ));
 sg13g2_a221oi_1 _4494_ (.B2(_1465_),
    .C1(_1451_),
    .B1(_1463_),
    .A1(_1443_),
    .Y(_1466_),
    .A2(_1444_));
 sg13g2_a21oi_1 _4495_ (.A1(_0914_),
    .A2(_0200_),
    .Y(_1467_),
    .B1(_1443_));
 sg13g2_nand2_1 _4496_ (.Y(_1468_),
    .A(net943),
    .B(net635));
 sg13g2_nor3_1 _4497_ (.A(_1466_),
    .B(_1467_),
    .C(_1468_),
    .Y(_0238_));
 sg13g2_and3_1 _4498_ (.X(_1469_),
    .A(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[0] ),
    .B(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[1] ),
    .C(net1277));
 sg13g2_and2_1 _4499_ (.A(net1483),
    .B(_1469_),
    .X(_1470_));
 sg13g2_nand2_1 _4500_ (.Y(_1471_),
    .A(net1710),
    .B(_1470_));
 sg13g2_o21ai_1 _4501_ (.B1(net919),
    .Y(_1472_),
    .A1(_0917_),
    .A2(_1471_));
 sg13g2_nor2_1 _4502_ (.A(_0956_),
    .B(_1472_),
    .Y(_0239_));
 sg13g2_xnor2_1 _4503_ (.Y(_1473_),
    .A(net1555),
    .B(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[1] ));
 sg13g2_nor2_1 _4504_ (.A(_1472_),
    .B(net1556),
    .Y(_0240_));
 sg13g2_a21oi_1 _4505_ (.A1(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[0] ),
    .A2(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[1] ),
    .Y(_1474_),
    .B1(net1277));
 sg13g2_nor3_1 _4506_ (.A(net892),
    .B(_1469_),
    .C(net1278),
    .Y(_0241_));
 sg13g2_o21ai_1 _4507_ (.B1(net920),
    .Y(_1475_),
    .A1(net1483),
    .A2(_1469_));
 sg13g2_nor2_1 _4508_ (.A(_1470_),
    .B(net1484),
    .Y(_0242_));
 sg13g2_or2_1 _4509_ (.X(_1476_),
    .B(_1470_),
    .A(net1710));
 sg13g2_and3_1 _4510_ (.X(_0243_),
    .A(net919),
    .B(_1471_),
    .C(_1476_));
 sg13g2_a21oi_1 _4511_ (.A1(_0917_),
    .A2(_1471_),
    .Y(_0244_),
    .B1(_1472_));
 sg13g2_nand2_2 _4512_ (.Y(_1477_),
    .A(net836),
    .B(_1454_));
 sg13g2_and2_1 _4513_ (.A(_0899_),
    .B(_1477_),
    .X(_1478_));
 sg13g2_xnor2_1 _4514_ (.Y(_1479_),
    .A(net832),
    .B(_1477_));
 sg13g2_inv_1 _4515_ (.Y(_1480_),
    .A(_1479_));
 sg13g2_xnor2_1 _4516_ (.Y(_1481_),
    .A(net835),
    .B(_1453_));
 sg13g2_nor2b_1 _4517_ (.A(_1479_),
    .B_N(_1481_),
    .Y(_1482_));
 sg13g2_nor2_1 _4518_ (.A(net837),
    .B(net839),
    .Y(_1483_));
 sg13g2_nor3_1 _4519_ (.A(net836),
    .B(_0167_),
    .C(_0971_),
    .Y(_1484_));
 sg13g2_a21oi_1 _4520_ (.A1(_1453_),
    .A2(_1482_),
    .Y(_1485_),
    .B1(_1484_));
 sg13g2_nor2_1 _4521_ (.A(_0167_),
    .B(_0969_),
    .Y(_1486_));
 sg13g2_a22oi_1 _4522_ (.Y(_1487_),
    .B1(_1486_),
    .B2(_0896_),
    .A2(_1480_),
    .A1(_0964_));
 sg13g2_nand2_1 _4523_ (.Y(_1488_),
    .A(_0968_),
    .B(_1482_));
 sg13g2_and2_1 _4524_ (.A(_0940_),
    .B(_1477_),
    .X(_1489_));
 sg13g2_xnor2_1 _4525_ (.Y(_1490_),
    .A(_0940_),
    .B(_1477_));
 sg13g2_nand2_1 _4526_ (.Y(_1491_),
    .A(_1481_),
    .B(_1490_));
 sg13g2_nor2_2 _4527_ (.A(net831),
    .B(_0963_),
    .Y(_1492_));
 sg13g2_nor2_2 _4528_ (.A(net836),
    .B(_1454_),
    .Y(_1493_));
 sg13g2_nand2_1 _4529_ (.Y(_1494_),
    .A(_0896_),
    .B(_1453_));
 sg13g2_a22oi_1 _4530_ (.Y(_1495_),
    .B1(_1494_),
    .B2(_1478_),
    .A2(_1492_),
    .A1(_0896_));
 sg13g2_and2_1 _4531_ (.A(_1491_),
    .B(_1495_),
    .X(_1496_));
 sg13g2_nand3_1 _4532_ (.B(_1488_),
    .C(_1496_),
    .A(_1485_),
    .Y(_1497_));
 sg13g2_nand4_1 _4533_ (.B(_1487_),
    .C(_1488_),
    .A(_1485_),
    .Y(_1498_),
    .D(_1496_));
 sg13g2_inv_1 _4534_ (.Y(_1499_),
    .A(_1498_));
 sg13g2_nand2_1 _4535_ (.Y(_1500_),
    .A(_1485_),
    .B(_1498_));
 sg13g2_a21oi_1 _4536_ (.A1(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[0] ),
    .A2(_0224_),
    .Y(_1501_),
    .B1(_1500_));
 sg13g2_and2_1 _4537_ (.A(_1487_),
    .B(_1497_),
    .X(_1502_));
 sg13g2_a22oi_1 _4538_ (.Y(_1503_),
    .B1(_1502_),
    .B2(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[1] ),
    .A2(_1500_),
    .A1(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[0] ));
 sg13g2_nand2b_1 _4539_ (.Y(_1504_),
    .B(_1503_),
    .A_N(_1501_));
 sg13g2_nand3b_1 _4540_ (.B(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[4] ),
    .C(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[2] ),
    .Y(_1505_),
    .A_N(_0198_));
 sg13g2_nor2_1 _4541_ (.A(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[1] ),
    .B(_1502_),
    .Y(_1506_));
 sg13g2_a21oi_1 _4542_ (.A1(_1460_),
    .A2(_1505_),
    .Y(_1507_),
    .B1(_1506_));
 sg13g2_nand2b_1 _4543_ (.Y(_1508_),
    .B(_0198_),
    .A_N(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[2] ));
 sg13g2_o21ai_1 _4544_ (.B1(_1459_),
    .Y(_1509_),
    .A1(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[4] ),
    .A2(_1508_));
 sg13g2_nand3_1 _4545_ (.B(net646),
    .C(_1509_),
    .A(net945),
    .Y(_1510_));
 sg13g2_a21oi_1 _4546_ (.A1(_1504_),
    .A2(_1507_),
    .Y(_0245_),
    .B1(net647));
 sg13g2_and3_1 _4547_ (.X(_1511_),
    .A(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[0] ),
    .B(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[1] ),
    .C(net1274));
 sg13g2_and2_1 _4548_ (.A(net1403),
    .B(_1511_),
    .X(_1512_));
 sg13g2_nand2_1 _4549_ (.Y(_1513_),
    .A(net1727),
    .B(_1512_));
 sg13g2_o21ai_1 _4550_ (.B1(net921),
    .Y(_1514_),
    .A1(_0918_),
    .A2(_1513_));
 sg13g2_nor2_1 _4551_ (.A(_0952_),
    .B(_1514_),
    .Y(_0246_));
 sg13g2_xnor2_1 _4552_ (.Y(_1515_),
    .A(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[0] ),
    .B(net1423));
 sg13g2_nor2_1 _4553_ (.A(_1514_),
    .B(net1424),
    .Y(_0247_));
 sg13g2_a21oi_1 _4554_ (.A1(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[0] ),
    .A2(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[1] ),
    .Y(_1516_),
    .B1(net1274));
 sg13g2_nor3_1 _4555_ (.A(net891),
    .B(_1511_),
    .C(net1275),
    .Y(_0248_));
 sg13g2_o21ai_1 _4556_ (.B1(net921),
    .Y(_1517_),
    .A1(net1403),
    .A2(_1511_));
 sg13g2_nor2_1 _4557_ (.A(_1512_),
    .B(net1404),
    .Y(_0249_));
 sg13g2_or2_1 _4558_ (.X(_1518_),
    .B(_1512_),
    .A(net1727));
 sg13g2_and3_1 _4559_ (.X(_0250_),
    .A(net921),
    .B(_1513_),
    .C(_1518_));
 sg13g2_a21oi_1 _4560_ (.A1(_0918_),
    .A2(_1513_),
    .Y(_0251_),
    .B1(_1514_));
 sg13g2_nand3_1 _4561_ (.B(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[2] ),
    .C(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[4] ),
    .A(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[1] ),
    .Y(_1519_));
 sg13g2_o21ai_1 _4562_ (.B1(_1499_),
    .Y(_1520_),
    .A1(_0196_),
    .A2(_1519_));
 sg13g2_nor2_1 _4563_ (.A(net833),
    .B(_0971_),
    .Y(_1521_));
 sg13g2_nor2_2 _4564_ (.A(net836),
    .B(net832),
    .Y(_1522_));
 sg13g2_nor2b_1 _4565_ (.A(_0971_),
    .B_N(_1522_),
    .Y(_1523_));
 sg13g2_nand2_1 _4566_ (.Y(_1524_),
    .A(_0970_),
    .B(_1522_));
 sg13g2_o21ai_1 _4567_ (.B1(_1524_),
    .Y(_1525_),
    .A1(_0969_),
    .A2(_1448_));
 sg13g2_xnor2_1 _4568_ (.Y(_1526_),
    .A(net833),
    .B(_1483_));
 sg13g2_nor2_1 _4569_ (.A(_0203_),
    .B(_1446_),
    .Y(_1527_));
 sg13g2_or4_1 _4570_ (.A(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[0] ),
    .B(_1525_),
    .C(_1526_),
    .D(_1527_),
    .X(_1528_));
 sg13g2_nor3_1 _4571_ (.A(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[1] ),
    .B(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[2] ),
    .C(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[4] ),
    .Y(_1529_));
 sg13g2_nand2_1 _4572_ (.Y(_1530_),
    .A(_0196_),
    .B(_1529_));
 sg13g2_nand2_1 _4573_ (.Y(_1531_),
    .A(net919),
    .B(net665));
 sg13g2_a221oi_1 _4574_ (.B2(_1498_),
    .C1(_1531_),
    .B1(_1530_),
    .A1(_1520_),
    .Y(_0252_),
    .A2(_1528_));
 sg13g2_and3_1 _4575_ (.X(_1532_),
    .A(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[0] ),
    .B(net1370),
    .C(net692));
 sg13g2_and2_1 _4576_ (.A(net1593),
    .B(_1532_),
    .X(_1533_));
 sg13g2_nand2_1 _4577_ (.Y(_1534_),
    .A(net1723),
    .B(_1533_));
 sg13g2_o21ai_1 _4578_ (.B1(net919),
    .Y(_1535_),
    .A1(_0919_),
    .A2(_1534_));
 sg13g2_nor2b_1 _4579_ (.A(_1535_),
    .B_N(net618),
    .Y(_0253_));
 sg13g2_xnor2_1 _4580_ (.Y(_1536_),
    .A(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[0] ),
    .B(net1370));
 sg13g2_nor2_1 _4581_ (.A(_1535_),
    .B(net1371),
    .Y(_0254_));
 sg13g2_a21oi_1 _4582_ (.A1(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[0] ),
    .A2(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[1] ),
    .Y(_1537_),
    .B1(net692));
 sg13g2_nor3_1 _4583_ (.A(net891),
    .B(_1532_),
    .C(net693),
    .Y(_0255_));
 sg13g2_o21ai_1 _4584_ (.B1(net919),
    .Y(_1538_),
    .A1(net1593),
    .A2(_1532_));
 sg13g2_nor2_1 _4585_ (.A(_1533_),
    .B(net1594),
    .Y(_0256_));
 sg13g2_or2_1 _4586_ (.X(_1539_),
    .B(_1533_),
    .A(net1723));
 sg13g2_and3_1 _4587_ (.X(_0257_),
    .A(net919),
    .B(_1534_),
    .C(_1539_));
 sg13g2_a21oi_1 _4588_ (.A1(_0919_),
    .A2(_1534_),
    .Y(_0258_),
    .B1(_1535_));
 sg13g2_nor2_1 _4589_ (.A(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[0] ),
    .B(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[2] ),
    .Y(_1540_));
 sg13g2_nand4_1 _4590_ (.B(_0194_),
    .C(_0952_),
    .A(_0193_),
    .Y(_1541_),
    .D(_1540_));
 sg13g2_nand2_1 _4591_ (.Y(_1542_),
    .A(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[4] ),
    .B(_1541_));
 sg13g2_nor2_1 _4592_ (.A(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[4] ),
    .B(_1541_),
    .Y(_1543_));
 sg13g2_a221oi_1 _4593_ (.B2(_1542_),
    .C1(_1543_),
    .B1(_1525_),
    .A1(_0203_),
    .Y(_1544_),
    .A2(_1445_));
 sg13g2_nor3_1 _4594_ (.A(_0193_),
    .B(_0194_),
    .C(_0222_),
    .Y(_1545_));
 sg13g2_nand3_1 _4595_ (.B(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[4] ),
    .C(_1545_),
    .A(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[2] ),
    .Y(_1546_));
 sg13g2_nand3_1 _4596_ (.B(net682),
    .C(_1546_),
    .A(net921),
    .Y(_1547_));
 sg13g2_nor2_1 _4597_ (.A(_1544_),
    .B(net683),
    .Y(_0259_));
 sg13g2_and3_1 _4598_ (.X(_1548_),
    .A(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[0] ),
    .B(net1352),
    .C(net1395));
 sg13g2_and2_1 _4599_ (.A(net1606),
    .B(_1548_),
    .X(_1549_));
 sg13g2_nand2_1 _4600_ (.Y(_1550_),
    .A(net1705),
    .B(_1549_));
 sg13g2_o21ai_1 _4601_ (.B1(net921),
    .Y(_1551_),
    .A1(_0921_),
    .A2(_1550_));
 sg13g2_nor2_1 _4602_ (.A(_0951_),
    .B(_1551_),
    .Y(_0260_));
 sg13g2_xnor2_1 _4603_ (.Y(_1552_),
    .A(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[0] ),
    .B(net1352));
 sg13g2_nor2_1 _4604_ (.A(_1551_),
    .B(net1353),
    .Y(_0261_));
 sg13g2_a21oi_1 _4605_ (.A1(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[0] ),
    .A2(net1352),
    .Y(_1553_),
    .B1(net1395));
 sg13g2_nor3_1 _4606_ (.A(net891),
    .B(_1548_),
    .C(net1396),
    .Y(_0262_));
 sg13g2_o21ai_1 _4607_ (.B1(net919),
    .Y(_1554_),
    .A1(net1606),
    .A2(_1548_));
 sg13g2_nor2_1 _4608_ (.A(_1549_),
    .B(net1607),
    .Y(_0263_));
 sg13g2_or2_1 _4609_ (.X(_1555_),
    .B(_1549_),
    .A(net1705));
 sg13g2_and3_1 _4610_ (.X(_0264_),
    .A(net921),
    .B(_1550_),
    .C(_1555_));
 sg13g2_a21oi_1 _4611_ (.A1(_0921_),
    .A2(_1550_),
    .Y(_0265_),
    .B1(_1551_));
 sg13g2_nor3_1 _4612_ (.A(net834),
    .B(net831),
    .C(_1454_),
    .Y(_1556_));
 sg13g2_nor2_1 _4613_ (.A(_1523_),
    .B(_1556_),
    .Y(_1557_));
 sg13g2_xnor2_1 _4614_ (.Y(_1558_),
    .A(net831),
    .B(_0964_));
 sg13g2_nor4_1 _4615_ (.A(net839),
    .B(_0897_),
    .C(net834),
    .D(net831),
    .Y(_1559_));
 sg13g2_nor3_1 _4616_ (.A(net837),
    .B(net841),
    .C(net833),
    .Y(_1560_));
 sg13g2_a21oi_1 _4617_ (.A1(net834),
    .A2(_1492_),
    .Y(_1561_),
    .B1(_1560_));
 sg13g2_a221oi_1 _4618_ (.B2(_0967_),
    .C1(_1559_),
    .B1(_1558_),
    .A1(_0965_),
    .Y(_1562_),
    .A2(_1439_));
 sg13g2_and2_1 _4619_ (.A(_0968_),
    .B(_1522_),
    .X(_1563_));
 sg13g2_a21oi_1 _4620_ (.A1(net834),
    .A2(_1492_),
    .Y(_1564_),
    .B1(_1563_));
 sg13g2_nand2_2 _4621_ (.Y(_1565_),
    .A(_1453_),
    .B(_1522_));
 sg13g2_nand2_1 _4622_ (.Y(_1566_),
    .A(_1561_),
    .B(_1562_));
 sg13g2_nand3_1 _4623_ (.B(_1561_),
    .C(_1562_),
    .A(_1557_),
    .Y(_1567_));
 sg13g2_nor2_1 _4624_ (.A(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[4] ),
    .B(_1557_),
    .Y(_1568_));
 sg13g2_nor2_1 _4625_ (.A(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[3] ),
    .B(_1564_),
    .Y(_1569_));
 sg13g2_nor2_1 _4626_ (.A(_1568_),
    .B(_1569_),
    .Y(_1570_));
 sg13g2_nand3_1 _4627_ (.B(_1557_),
    .C(_1566_),
    .A(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[4] ),
    .Y(_1571_));
 sg13g2_nand4_1 _4628_ (.B(net674),
    .C(_1534_),
    .A(net919),
    .Y(_1572_),
    .D(_1571_));
 sg13g2_a21oi_1 _4629_ (.A1(_1567_),
    .A2(_1570_),
    .Y(_0266_),
    .B1(net675));
 sg13g2_and3_1 _4630_ (.X(_1573_),
    .A(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[0] ),
    .B(net1364),
    .C(net1230));
 sg13g2_and2_1 _4631_ (.A(net1461),
    .B(_1573_),
    .X(_1574_));
 sg13g2_nand2_1 _4632_ (.Y(_1575_),
    .A(net1732),
    .B(_1574_));
 sg13g2_o21ai_1 _4633_ (.B1(net948),
    .Y(_1576_),
    .A1(_0922_),
    .A2(_1575_));
 sg13g2_nor2_1 _4634_ (.A(_0948_),
    .B(_1576_),
    .Y(_0267_));
 sg13g2_xnor2_1 _4635_ (.Y(_1577_),
    .A(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[0] ),
    .B(net1364));
 sg13g2_nor2_1 _4636_ (.A(_1576_),
    .B(net1365),
    .Y(_0268_));
 sg13g2_a21oi_1 _4637_ (.A1(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[0] ),
    .A2(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[1] ),
    .Y(_1578_),
    .B1(net1230));
 sg13g2_nor3_1 _4638_ (.A(net904),
    .B(_1573_),
    .C(net1231),
    .Y(_0269_));
 sg13g2_o21ai_1 _4639_ (.B1(net948),
    .Y(_1579_),
    .A1(net1461),
    .A2(_1573_));
 sg13g2_nor2_1 _4640_ (.A(_1574_),
    .B(net1462),
    .Y(_0270_));
 sg13g2_or2_1 _4641_ (.X(_1580_),
    .B(_1574_),
    .A(net1732));
 sg13g2_and3_1 _4642_ (.X(_0271_),
    .A(net948),
    .B(_1575_),
    .C(_1580_));
 sg13g2_a21oi_1 _4643_ (.A1(_0922_),
    .A2(_1575_),
    .Y(_0272_),
    .B1(_1576_));
 sg13g2_nor2_1 _4644_ (.A(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[4] ),
    .B(_1567_),
    .Y(_1581_));
 sg13g2_a21oi_1 _4645_ (.A1(net841),
    .A2(_1445_),
    .Y(_1582_),
    .B1(_1560_));
 sg13g2_or2_1 _4646_ (.X(_1583_),
    .B(_1582_),
    .A(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[3] ));
 sg13g2_nand2_2 _4647_ (.Y(_1584_),
    .A(_1455_),
    .B(_1565_));
 sg13g2_o21ai_1 _4648_ (.B1(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[2] ),
    .Y(_1585_),
    .A1(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[0] ),
    .A2(_0220_));
 sg13g2_and2_2 _4649_ (.A(_0962_),
    .B(_1522_),
    .X(_1586_));
 sg13g2_nor3_1 _4650_ (.A(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[0] ),
    .B(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[2] ),
    .C(_0220_),
    .Y(_1587_));
 sg13g2_o21ai_1 _4651_ (.B1(_1585_),
    .Y(_1588_),
    .A1(_1458_),
    .A2(_1586_));
 sg13g2_a21oi_1 _4652_ (.A1(_0190_),
    .A2(_1587_),
    .Y(_1589_),
    .B1(_1584_));
 sg13g2_nor3_1 _4653_ (.A(_0920_),
    .B(_0190_),
    .C(_0220_),
    .Y(_1590_));
 sg13g2_a221oi_1 _4654_ (.B2(_1589_),
    .C1(_1590_),
    .B1(_1588_),
    .A1(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[3] ),
    .Y(_1591_),
    .A2(_1582_));
 sg13g2_nor2_1 _4655_ (.A(_1581_),
    .B(_1591_),
    .Y(_1592_));
 sg13g2_nand2_1 _4656_ (.Y(_1593_),
    .A(net920),
    .B(net663));
 sg13g2_a221oi_1 _4657_ (.B2(_1592_),
    .C1(_1593_),
    .B1(_1583_),
    .A1(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[4] ),
    .Y(_0273_),
    .A2(_1567_));
 sg13g2_and3_1 _4658_ (.X(_1594_),
    .A(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[0] ),
    .B(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[1] ),
    .C(net1217));
 sg13g2_and2_1 _4659_ (.A(net1477),
    .B(_1594_),
    .X(_1595_));
 sg13g2_nand2_1 _4660_ (.Y(_1596_),
    .A(net1702),
    .B(_1595_));
 sg13g2_o21ai_1 _4661_ (.B1(net922),
    .Y(_1597_),
    .A1(_0909_),
    .A2(_1596_));
 sg13g2_nor2_1 _4662_ (.A(_0957_),
    .B(_1597_),
    .Y(_0274_));
 sg13g2_xnor2_1 _4663_ (.Y(_1598_),
    .A(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[0] ),
    .B(net1533));
 sg13g2_nor2_1 _4664_ (.A(_1597_),
    .B(net1534),
    .Y(_0275_));
 sg13g2_a21oi_1 _4665_ (.A1(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[0] ),
    .A2(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[1] ),
    .Y(_1599_),
    .B1(net1217));
 sg13g2_nor3_1 _4666_ (.A(net892),
    .B(_1594_),
    .C(net1218),
    .Y(_0276_));
 sg13g2_o21ai_1 _4667_ (.B1(net922),
    .Y(_1600_),
    .A1(net1477),
    .A2(_1594_));
 sg13g2_nor2_1 _4668_ (.A(_1595_),
    .B(net1478),
    .Y(_0277_));
 sg13g2_or2_1 _4669_ (.X(_1601_),
    .B(_1595_),
    .A(net1702));
 sg13g2_and3_1 _4670_ (.X(_0278_),
    .A(net922),
    .B(_1596_),
    .C(_1601_));
 sg13g2_a21oi_1 _4671_ (.A1(_0909_),
    .A2(_1596_),
    .Y(_0279_),
    .B1(_1597_));
 sg13g2_nor3_2 _4672_ (.A(net834),
    .B(net831),
    .C(_0969_),
    .Y(_1602_));
 sg13g2_nor2_2 _4673_ (.A(_0896_),
    .B(net832),
    .Y(_1603_));
 sg13g2_nor2_2 _4674_ (.A(net833),
    .B(_1457_),
    .Y(_1604_));
 sg13g2_nor2_1 _4675_ (.A(_1559_),
    .B(_1604_),
    .Y(_1605_));
 sg13g2_nand2_1 _4676_ (.Y(_1606_),
    .A(net832),
    .B(_1494_));
 sg13g2_nand3_1 _4677_ (.B(_1565_),
    .C(_1606_),
    .A(_1481_),
    .Y(_1607_));
 sg13g2_a221oi_1 _4678_ (.B2(_1494_),
    .C1(_1563_),
    .B1(_1489_),
    .A1(_0940_),
    .Y(_1608_),
    .A2(_0964_));
 sg13g2_nand3_1 _4679_ (.B(_1607_),
    .C(_1608_),
    .A(_1605_),
    .Y(_1609_));
 sg13g2_inv_1 _4680_ (.Y(_1610_),
    .A(_1609_));
 sg13g2_nor3_2 _4681_ (.A(_1586_),
    .B(_1602_),
    .C(_1609_),
    .Y(_1611_));
 sg13g2_nand2_1 _4682_ (.Y(_1612_),
    .A(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[0] ),
    .B(net1716));
 sg13g2_nand3_1 _4683_ (.B(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[1] ),
    .C(_1611_),
    .A(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[0] ),
    .Y(_1613_));
 sg13g2_nor3_1 _4684_ (.A(_1586_),
    .B(_1602_),
    .C(_1610_),
    .Y(_1614_));
 sg13g2_nand2_1 _4685_ (.Y(_1615_),
    .A(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[0] ),
    .B(_0206_));
 sg13g2_nand2_1 _4686_ (.Y(_1616_),
    .A(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[1] ),
    .B(_1615_));
 sg13g2_o21ai_1 _4687_ (.B1(_1605_),
    .Y(_1617_),
    .A1(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[1] ),
    .A2(_1615_));
 sg13g2_a21oi_1 _4688_ (.A1(_1616_),
    .A2(_1617_),
    .Y(_1618_),
    .B1(_1611_));
 sg13g2_a21oi_1 _4689_ (.A1(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[2] ),
    .A2(_1614_),
    .Y(_1619_),
    .B1(_1618_));
 sg13g2_o21ai_1 _4690_ (.B1(_1584_),
    .Y(_1620_),
    .A1(_0910_),
    .A2(_0177_));
 sg13g2_o21ai_1 _4691_ (.B1(_1620_),
    .Y(_1621_),
    .A1(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[2] ),
    .A2(_1614_));
 sg13g2_a21oi_1 _4692_ (.A1(_1613_),
    .A2(_1619_),
    .Y(_1622_),
    .B1(_1621_));
 sg13g2_a21oi_1 _4693_ (.A1(_0910_),
    .A2(_0177_),
    .Y(_1623_),
    .B1(_1584_));
 sg13g2_nand2_1 _4694_ (.Y(_1624_),
    .A(net920),
    .B(net655));
 sg13g2_nor3_1 _4695_ (.A(_1622_),
    .B(_1623_),
    .C(_1624_),
    .Y(_0280_));
 sg13g2_and3_1 _4696_ (.X(_1625_),
    .A(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[0] ),
    .B(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[1] ),
    .C(net1343));
 sg13g2_and2_1 _4697_ (.A(net1410),
    .B(_1625_),
    .X(_1626_));
 sg13g2_nand2_1 _4698_ (.Y(_1627_),
    .A(net1725),
    .B(_1626_));
 sg13g2_o21ai_1 _4699_ (.B1(net923),
    .Y(_1628_),
    .A1(_0908_),
    .A2(_1627_));
 sg13g2_nor2_1 _4700_ (.A(_0958_),
    .B(_1628_),
    .Y(_0281_));
 sg13g2_xnor2_1 _4701_ (.Y(_1629_),
    .A(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[0] ),
    .B(net1412));
 sg13g2_nor2_1 _4702_ (.A(_1628_),
    .B(net1413),
    .Y(_0282_));
 sg13g2_a21oi_1 _4703_ (.A1(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[0] ),
    .A2(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[1] ),
    .Y(_1630_),
    .B1(net1343));
 sg13g2_nor3_1 _4704_ (.A(net892),
    .B(_1625_),
    .C(net1344),
    .Y(_0283_));
 sg13g2_o21ai_1 _4705_ (.B1(net923),
    .Y(_1631_),
    .A1(net1410),
    .A2(_1625_));
 sg13g2_nor2_1 _4706_ (.A(_1626_),
    .B(net1411),
    .Y(_0284_));
 sg13g2_or2_1 _4707_ (.X(_1632_),
    .B(_1626_),
    .A(net1725));
 sg13g2_and3_1 _4708_ (.X(_0285_),
    .A(net923),
    .B(_1627_),
    .C(_1632_));
 sg13g2_a21oi_1 _4709_ (.A1(_0908_),
    .A2(_1627_),
    .Y(_0286_),
    .B1(_1628_));
 sg13g2_and2_1 _4710_ (.A(net837),
    .B(net839),
    .X(_1633_));
 sg13g2_a21oi_1 _4711_ (.A1(_0967_),
    .A2(_1492_),
    .Y(_1634_),
    .B1(_1604_));
 sg13g2_inv_1 _4712_ (.Y(_1635_),
    .A(_1634_));
 sg13g2_or3_1 _4713_ (.A(net831),
    .B(_1483_),
    .C(_1633_),
    .X(_1636_));
 sg13g2_a21oi_1 _4714_ (.A1(net831),
    .A2(_1493_),
    .Y(_1637_),
    .B1(_1586_));
 sg13g2_o21ai_1 _4715_ (.B1(net836),
    .Y(_1638_),
    .A1(_1486_),
    .A2(_1521_));
 sg13g2_o21ai_1 _4716_ (.B1(_1526_),
    .Y(_1639_),
    .A1(_1483_),
    .A2(_1633_));
 sg13g2_nand4_1 _4717_ (.B(_1637_),
    .C(_1638_),
    .A(_1636_),
    .Y(_1640_),
    .D(_1639_));
 sg13g2_nor2_2 _4718_ (.A(_1635_),
    .B(_1640_),
    .Y(_1641_));
 sg13g2_a21oi_1 _4719_ (.A1(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[1] ),
    .A2(_1634_),
    .Y(_1642_),
    .B1(_1638_));
 sg13g2_nor2_1 _4720_ (.A(_1641_),
    .B(_1642_),
    .Y(_1643_));
 sg13g2_nand3b_1 _4721_ (.B(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[4] ),
    .C(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[2] ),
    .Y(_1644_),
    .A_N(_0179_));
 sg13g2_a21oi_1 _4722_ (.A1(_1634_),
    .A2(_1640_),
    .Y(_1645_),
    .B1(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[1] ));
 sg13g2_a21oi_1 _4723_ (.A1(_1611_),
    .A2(_1644_),
    .Y(_1646_),
    .B1(_1645_));
 sg13g2_o21ai_1 _4724_ (.B1(_1646_),
    .Y(_1647_),
    .A1(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[0] ),
    .A2(_1643_));
 sg13g2_nor2_1 _4725_ (.A(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[2] ),
    .B(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[4] ),
    .Y(_1648_));
 sg13g2_a21o_1 _4726_ (.A2(_1648_),
    .A1(_0179_),
    .B1(_1611_),
    .X(_1649_));
 sg13g2_and4_1 _4727_ (.A(net922),
    .B(net649),
    .C(_1647_),
    .D(_1649_),
    .X(_0287_));
 sg13g2_and3_1 _4728_ (.X(_1650_),
    .A(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[0] ),
    .B(net1379),
    .C(net699));
 sg13g2_and2_1 _4729_ (.A(net1481),
    .B(_1650_),
    .X(_1651_));
 sg13g2_nand2_1 _4730_ (.Y(_1652_),
    .A(net1724),
    .B(_1651_));
 sg13g2_o21ai_1 _4731_ (.B1(net949),
    .Y(_1653_),
    .A1(_0907_),
    .A2(_1652_));
 sg13g2_nor2_1 _4732_ (.A(_0959_),
    .B(_1653_),
    .Y(_0288_));
 sg13g2_xnor2_1 _4733_ (.Y(_1654_),
    .A(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[0] ),
    .B(net1379));
 sg13g2_nor2_1 _4734_ (.A(_1653_),
    .B(net1380),
    .Y(_0289_));
 sg13g2_a21oi_1 _4735_ (.A1(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[0] ),
    .A2(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[1] ),
    .Y(_1655_),
    .B1(net699));
 sg13g2_nor3_1 _4736_ (.A(net902),
    .B(_1650_),
    .C(net700),
    .Y(_0290_));
 sg13g2_o21ai_1 _4737_ (.B1(net950),
    .Y(_1656_),
    .A1(net1481),
    .A2(_1650_));
 sg13g2_nor2_1 _4738_ (.A(_1651_),
    .B(net1482),
    .Y(_0291_));
 sg13g2_or2_1 _4739_ (.X(_1657_),
    .B(_1651_),
    .A(net1724));
 sg13g2_and3_1 _4740_ (.X(_0292_),
    .A(net949),
    .B(_1652_),
    .C(_1657_));
 sg13g2_a21oi_1 _4741_ (.A1(_0907_),
    .A2(_1652_),
    .Y(_0293_),
    .B1(_1653_));
 sg13g2_xnor2_1 _4742_ (.Y(_1658_),
    .A(net826),
    .B(_1439_));
 sg13g2_and2_1 _4743_ (.A(_0204_),
    .B(_1658_),
    .X(_1659_));
 sg13g2_a22oi_1 _4744_ (.Y(_1660_),
    .B1(_1659_),
    .B2(_0968_),
    .A2(_1492_),
    .A1(_0967_));
 sg13g2_a21oi_1 _4745_ (.A1(_0204_),
    .A2(_1440_),
    .Y(_1661_),
    .B1(_1658_));
 sg13g2_a21oi_1 _4746_ (.A1(_1441_),
    .A2(_1457_),
    .Y(_1662_),
    .B1(_1661_));
 sg13g2_a21oi_1 _4747_ (.A1(_0970_),
    .A2(_1442_),
    .Y(_1663_),
    .B1(_1662_));
 sg13g2_nand2_1 _4748_ (.Y(_1664_),
    .A(_1660_),
    .B(_1663_));
 sg13g2_a22oi_1 _4749_ (.Y(_1665_),
    .B1(_1659_),
    .B2(_0970_),
    .A2(_1493_),
    .A1(_1440_));
 sg13g2_a21oi_1 _4750_ (.A1(_1664_),
    .A2(_1665_),
    .Y(_1666_),
    .B1(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[0] ));
 sg13g2_nand4_1 _4751_ (.B(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[4] ),
    .C(_0949_),
    .A(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[2] ),
    .Y(_1667_),
    .D(_0950_));
 sg13g2_a21oi_1 _4752_ (.A1(_1641_),
    .A2(_1667_),
    .Y(_1668_),
    .B1(_1666_));
 sg13g2_nor3_1 _4753_ (.A(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[2] ),
    .B(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[4] ),
    .C(_0949_),
    .Y(_1669_));
 sg13g2_a21oi_1 _4754_ (.A1(_0188_),
    .A2(_1669_),
    .Y(_1670_),
    .B1(_1641_));
 sg13g2_nand2_1 _4755_ (.Y(_1671_),
    .A(net923),
    .B(net629));
 sg13g2_nor3_1 _4756_ (.A(_1668_),
    .B(_1670_),
    .C(_1671_),
    .Y(_0294_));
 sg13g2_and3_1 _4757_ (.X(_1672_),
    .A(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[0] ),
    .B(net1416),
    .C(net1234));
 sg13g2_and2_1 _4758_ (.A(net1634),
    .B(_1672_),
    .X(_1673_));
 sg13g2_nand2_1 _4759_ (.Y(_1674_),
    .A(net1726),
    .B(_1673_));
 sg13g2_o21ai_1 _4760_ (.B1(net944),
    .Y(_1675_),
    .A1(_0905_),
    .A2(_1674_));
 sg13g2_nor2_1 _4761_ (.A(_0946_),
    .B(_1675_),
    .Y(_0295_));
 sg13g2_xnor2_1 _4762_ (.Y(_1676_),
    .A(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[0] ),
    .B(net1416));
 sg13g2_nor2_1 _4763_ (.A(_1675_),
    .B(net1417),
    .Y(_0296_));
 sg13g2_a21oi_1 _4764_ (.A1(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[0] ),
    .A2(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[1] ),
    .Y(_1677_),
    .B1(net1234));
 sg13g2_nor3_1 _4765_ (.A(net899),
    .B(_1672_),
    .C(net1235),
    .Y(_0297_));
 sg13g2_o21ai_1 _4766_ (.B1(net944),
    .Y(_1678_),
    .A1(net1634),
    .A2(_1672_));
 sg13g2_nor2_1 _4767_ (.A(_1673_),
    .B(net1635),
    .Y(_0298_));
 sg13g2_or2_1 _4768_ (.X(_1679_),
    .B(_1673_),
    .A(net1726));
 sg13g2_and3_1 _4769_ (.X(_0299_),
    .A(net944),
    .B(_1674_),
    .C(_1679_));
 sg13g2_a21oi_1 _4770_ (.A1(_0905_),
    .A2(_1674_),
    .Y(_0300_),
    .B1(_1675_));
 sg13g2_nand3_1 _4771_ (.B(_1663_),
    .C(_1665_),
    .A(_1660_),
    .Y(_1680_));
 sg13g2_o21ai_1 _4772_ (.B1(_1680_),
    .Y(_1681_),
    .A1(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[4] ),
    .A2(_1660_));
 sg13g2_nand3b_1 _4773_ (.B(_1650_),
    .C(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[4] ),
    .Y(_1682_),
    .A_N(_0175_));
 sg13g2_and4_1 _4774_ (.A(net949),
    .B(net640),
    .C(_1681_),
    .D(_1682_),
    .X(_0301_));
 sg13g2_and3_1 _4775_ (.X(_1683_),
    .A(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[0] ),
    .B(net1337),
    .C(net1123));
 sg13g2_and2_1 _4776_ (.A(net1527),
    .B(_1683_),
    .X(_1684_));
 sg13g2_nand2_1 _4777_ (.Y(_1685_),
    .A(net1693),
    .B(_1684_));
 sg13g2_o21ai_1 _4778_ (.B1(net943),
    .Y(_1686_),
    .A1(_0904_),
    .A2(_1685_));
 sg13g2_nor2_1 _4779_ (.A(_0960_),
    .B(_1686_),
    .Y(_0302_));
 sg13g2_xnor2_1 _4780_ (.Y(_1687_),
    .A(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[0] ),
    .B(net1337));
 sg13g2_nor2_1 _4781_ (.A(_1686_),
    .B(net1338),
    .Y(_0303_));
 sg13g2_a21oi_1 _4782_ (.A1(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[0] ),
    .A2(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[1] ),
    .Y(_1688_),
    .B1(net1123));
 sg13g2_nor3_1 _4783_ (.A(net900),
    .B(_1683_),
    .C(net1124),
    .Y(_0304_));
 sg13g2_o21ai_1 _4784_ (.B1(net943),
    .Y(_1689_),
    .A1(net1527),
    .A2(_1683_));
 sg13g2_nor2_1 _4785_ (.A(_1684_),
    .B(net1528),
    .Y(_0305_));
 sg13g2_or2_1 _4786_ (.X(_1690_),
    .B(_1684_),
    .A(net1693));
 sg13g2_and3_1 _4787_ (.X(_0306_),
    .A(net944),
    .B(_1685_),
    .C(_1690_));
 sg13g2_a21oi_1 _4788_ (.A1(_0904_),
    .A2(_1685_),
    .Y(_0307_),
    .B1(_1686_));
 sg13g2_a21oi_1 _4789_ (.A1(_0968_),
    .A2(_1603_),
    .Y(_1691_),
    .B1(_1523_));
 sg13g2_nor2_1 _4790_ (.A(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[0] ),
    .B(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[2] ),
    .Y(_1692_));
 sg13g2_nand3_1 _4791_ (.B(_0946_),
    .C(_1692_),
    .A(_0173_),
    .Y(_1693_));
 sg13g2_o21ai_1 _4792_ (.B1(_1565_),
    .Y(_1694_),
    .A1(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[3] ),
    .A2(_1693_));
 sg13g2_a21oi_1 _4793_ (.A1(_0962_),
    .A2(_1603_),
    .Y(_1695_),
    .B1(_1694_));
 sg13g2_a221oi_1 _4794_ (.B2(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[3] ),
    .C1(_1695_),
    .B1(_1693_),
    .A1(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[4] ),
    .Y(_1696_),
    .A2(_1691_));
 sg13g2_or2_1 _4795_ (.X(_1697_),
    .B(_1604_),
    .A(_1586_));
 sg13g2_nand4_1 _4796_ (.B(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[2] ),
    .C(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[4] ),
    .A(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[3] ),
    .Y(_1698_),
    .D(_0946_));
 sg13g2_o21ai_1 _4797_ (.B1(_1697_),
    .Y(_1699_),
    .A1(_0173_),
    .A2(_1698_));
 sg13g2_o21ai_1 _4798_ (.B1(_1699_),
    .Y(_1700_),
    .A1(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[4] ),
    .A2(_1691_));
 sg13g2_nor2_1 _4799_ (.A(_1696_),
    .B(_1700_),
    .Y(_1701_));
 sg13g2_nor3_2 _4800_ (.A(net899),
    .B(_0945_),
    .C(_1701_),
    .Y(_0308_));
 sg13g2_nand2_1 _4801_ (.Y(_1702_),
    .A(net1694),
    .B(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[1] ));
 sg13g2_and3_1 _4802_ (.X(_1703_),
    .A(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[0] ),
    .B(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[1] ),
    .C(net1184));
 sg13g2_and2_1 _4803_ (.A(net1479),
    .B(_1703_),
    .X(_1704_));
 sg13g2_nand2_1 _4804_ (.Y(_1705_),
    .A(net1706),
    .B(_1704_));
 sg13g2_o21ai_1 _4805_ (.B1(net943),
    .Y(_1706_),
    .A1(_0902_),
    .A2(_1705_));
 sg13g2_nor2_1 _4806_ (.A(_0944_),
    .B(_1706_),
    .Y(_0309_));
 sg13g2_or2_1 _4807_ (.X(_1707_),
    .B(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[1] ),
    .A(net1694));
 sg13g2_and3_1 _4808_ (.X(_0310_),
    .A(net947),
    .B(net1695),
    .C(_1707_));
 sg13g2_a21oi_1 _4809_ (.A1(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[0] ),
    .A2(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[1] ),
    .Y(_1708_),
    .B1(net1184));
 sg13g2_nor3_1 _4810_ (.A(net900),
    .B(_1703_),
    .C(net1185),
    .Y(_0311_));
 sg13g2_o21ai_1 _4811_ (.B1(net943),
    .Y(_1709_),
    .A1(net1479),
    .A2(_1703_));
 sg13g2_nor2_1 _4812_ (.A(_1704_),
    .B(net1480),
    .Y(_0312_));
 sg13g2_or2_1 _4813_ (.X(_1710_),
    .B(_1704_),
    .A(net1706));
 sg13g2_and3_1 _4814_ (.X(_0313_),
    .A(net943),
    .B(_1705_),
    .C(_1710_));
 sg13g2_a21oi_1 _4815_ (.A1(_0902_),
    .A2(_1705_),
    .Y(_0314_),
    .B1(_1706_));
 sg13g2_o21ai_1 _4816_ (.B1(_1524_),
    .Y(_1711_),
    .A1(_1454_),
    .A2(_1491_));
 sg13g2_a21oi_1 _4817_ (.A1(_0964_),
    .A2(_1490_),
    .Y(_1712_),
    .B1(_1563_));
 sg13g2_nor2b_1 _4818_ (.A(_1711_),
    .B_N(_1712_),
    .Y(_1713_));
 sg13g2_nand2_1 _4819_ (.Y(_1714_),
    .A(_0969_),
    .B(_1481_));
 sg13g2_a21oi_1 _4820_ (.A1(_1490_),
    .A2(_1714_),
    .Y(_1715_),
    .B1(_1586_));
 sg13g2_nand3b_1 _4821_ (.B(_1713_),
    .C(_1715_),
    .Y(_1716_),
    .A_N(_1482_));
 sg13g2_o21ai_1 _4822_ (.B1(_1716_),
    .Y(_1717_),
    .A1(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[3] ),
    .A2(_1713_));
 sg13g2_nand3_1 _4823_ (.B(_1711_),
    .C(_1712_),
    .A(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[2] ),
    .Y(_1718_));
 sg13g2_nor2b_1 _4824_ (.A(_1684_),
    .B_N(_1718_),
    .Y(_1719_));
 sg13g2_a22oi_1 _4825_ (.Y(_1720_),
    .B1(_1717_),
    .B2(_1719_),
    .A2(_1697_),
    .A1(_0903_));
 sg13g2_and2_1 _4826_ (.A(net944),
    .B(net1485),
    .X(_1721_));
 sg13g2_o21ai_1 _4827_ (.B1(_1721_),
    .Y(_1722_),
    .A1(_0903_),
    .A2(_1697_));
 sg13g2_nor2_2 _4828_ (.A(_1720_),
    .B(net1486),
    .Y(_0315_));
 sg13g2_and3_1 _4829_ (.X(_1723_),
    .A(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[0] ),
    .B(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[1] ),
    .C(net1297));
 sg13g2_and2_1 _4830_ (.A(net1470),
    .B(_1723_),
    .X(_1724_));
 sg13g2_nand2_1 _4831_ (.Y(_1725_),
    .A(net1711),
    .B(_1724_));
 sg13g2_o21ai_1 _4832_ (.B1(net948),
    .Y(_1726_),
    .A1(_0901_),
    .A2(_1725_));
 sg13g2_nor2_1 _4833_ (.A(_0942_),
    .B(_1726_),
    .Y(_0316_));
 sg13g2_xnor2_1 _4834_ (.Y(_1727_),
    .A(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[0] ),
    .B(net1591));
 sg13g2_nor2_1 _4835_ (.A(_1726_),
    .B(net1592),
    .Y(_0317_));
 sg13g2_a21oi_1 _4836_ (.A1(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[0] ),
    .A2(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[1] ),
    .Y(_1728_),
    .B1(net1297));
 sg13g2_nor3_1 _4837_ (.A(net904),
    .B(_1723_),
    .C(net1298),
    .Y(_0318_));
 sg13g2_o21ai_1 _4838_ (.B1(net948),
    .Y(_1729_),
    .A1(net1470),
    .A2(_1723_));
 sg13g2_nor2_1 _4839_ (.A(_1724_),
    .B(net1471),
    .Y(_0319_));
 sg13g2_or2_1 _4840_ (.X(_1730_),
    .B(_1724_),
    .A(net1711));
 sg13g2_and3_1 _4841_ (.X(_0320_),
    .A(net949),
    .B(_1725_),
    .C(_1730_));
 sg13g2_a21oi_1 _4842_ (.A1(_0901_),
    .A2(_1725_),
    .Y(_0321_),
    .B1(_1726_));
 sg13g2_a21oi_1 _4843_ (.A1(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[4] ),
    .A2(_0943_),
    .Y(_1731_),
    .B1(_1716_));
 sg13g2_a21oi_1 _4844_ (.A1(net840),
    .A2(_0167_),
    .Y(_1732_),
    .B1(net832));
 sg13g2_nor2b_1 _4845_ (.A(_1732_),
    .B_N(net839),
    .Y(_1733_));
 sg13g2_o21ai_1 _4846_ (.B1(_0966_),
    .Y(_1734_),
    .A1(_1478_),
    .A2(_1733_));
 sg13g2_nor2_1 _4847_ (.A(_1484_),
    .B(_1563_),
    .Y(_1735_));
 sg13g2_nand3_1 _4848_ (.B(_1734_),
    .C(_1735_),
    .A(_1636_),
    .Y(_1736_));
 sg13g2_nand2b_1 _4849_ (.Y(_1737_),
    .B(_1702_),
    .A_N(_1736_));
 sg13g2_a21oi_2 _4850_ (.B1(_1586_),
    .Y(_1738_),
    .A2(_1493_),
    .A1(_0940_));
 sg13g2_nand3_1 _4851_ (.B(_1737_),
    .C(_1738_),
    .A(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[2] ),
    .Y(_1739_));
 sg13g2_nor2b_2 _4852_ (.A(_1736_),
    .B_N(_1738_),
    .Y(_1740_));
 sg13g2_nand2_1 _4853_ (.Y(_1741_),
    .A(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[0] ),
    .B(_0213_));
 sg13g2_nor2_1 _4854_ (.A(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[1] ),
    .B(_1741_),
    .Y(_1742_));
 sg13g2_a21oi_1 _4855_ (.A1(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[1] ),
    .A2(_1741_),
    .Y(_1743_),
    .B1(_1735_));
 sg13g2_nor3_1 _4856_ (.A(_1740_),
    .B(_1742_),
    .C(_1743_),
    .Y(_1744_));
 sg13g2_o21ai_1 _4857_ (.B1(_1744_),
    .Y(_1745_),
    .A1(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[2] ),
    .A2(_1738_));
 sg13g2_o21ai_1 _4858_ (.B1(_1716_),
    .Y(_1746_),
    .A1(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[4] ),
    .A2(_0943_));
 sg13g2_a21oi_1 _4859_ (.A1(_1739_),
    .A2(_1745_),
    .Y(_1747_),
    .B1(_1731_));
 sg13g2_nand3_1 _4860_ (.B(net671),
    .C(_1746_),
    .A(net943),
    .Y(_1748_));
 sg13g2_nor2_1 _4861_ (.A(_1747_),
    .B(net672),
    .Y(_0322_));
 sg13g2_and3_1 _4862_ (.X(_1749_),
    .A(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[0] ),
    .B(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[1] ),
    .C(net1237));
 sg13g2_and2_1 _4863_ (.A(net1405),
    .B(_1749_),
    .X(_1750_));
 sg13g2_nand2_1 _4864_ (.Y(_1751_),
    .A(net1714),
    .B(_1750_));
 sg13g2_o21ai_1 _4865_ (.B1(net950),
    .Y(_1752_),
    .A1(_0924_),
    .A2(_1751_));
 sg13g2_nor2_1 _4866_ (.A(_0961_),
    .B(_1752_),
    .Y(_0323_));
 sg13g2_xnor2_1 _4867_ (.Y(_1753_),
    .A(net1518),
    .B(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[1] ));
 sg13g2_nor2_1 _4868_ (.A(_1752_),
    .B(net1519),
    .Y(_0324_));
 sg13g2_a21oi_1 _4869_ (.A1(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[0] ),
    .A2(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[1] ),
    .Y(_1754_),
    .B1(net1237));
 sg13g2_nor3_1 _4870_ (.A(net904),
    .B(_1749_),
    .C(net1238),
    .Y(_0325_));
 sg13g2_o21ai_1 _4871_ (.B1(net950),
    .Y(_1755_),
    .A1(net1405),
    .A2(_1749_));
 sg13g2_nor2_1 _4872_ (.A(_1750_),
    .B(net1406),
    .Y(_0326_));
 sg13g2_or2_1 _4873_ (.X(_1756_),
    .B(_1750_),
    .A(net1714));
 sg13g2_and3_1 _4874_ (.X(_0327_),
    .A(net948),
    .B(_1751_),
    .C(_1756_));
 sg13g2_a21oi_1 _4875_ (.A1(_0924_),
    .A2(_1751_),
    .Y(_0328_),
    .B1(_1752_));
 sg13g2_nand4_1 _4876_ (.B(_0897_),
    .C(net835),
    .A(net838),
    .Y(_1757_),
    .D(net832));
 sg13g2_nand3_1 _4877_ (.B(net826),
    .C(_0962_),
    .A(net835),
    .Y(_1758_));
 sg13g2_nand2_1 _4878_ (.Y(_1759_),
    .A(_1757_),
    .B(_1758_));
 sg13g2_nor4_1 _4879_ (.A(net838),
    .B(net840),
    .C(_0898_),
    .D(net826),
    .Y(_1760_));
 sg13g2_a21oi_1 _4880_ (.A1(_0898_),
    .A2(_1521_),
    .Y(_1761_),
    .B1(_1760_));
 sg13g2_xnor2_1 _4881_ (.Y(_1762_),
    .A(_0205_),
    .B(_0967_));
 sg13g2_nand3b_1 _4882_ (.B(_1761_),
    .C(_1762_),
    .Y(_1763_),
    .A_N(_1759_));
 sg13g2_nor4_1 _4883_ (.A(net838),
    .B(_0897_),
    .C(_0898_),
    .D(net826),
    .Y(_1764_));
 sg13g2_nor3_1 _4884_ (.A(net834),
    .B(net832),
    .C(_1454_),
    .Y(_1765_));
 sg13g2_or2_1 _4885_ (.X(_1766_),
    .B(_1765_),
    .A(_1764_));
 sg13g2_nor2_2 _4886_ (.A(_1763_),
    .B(_1766_),
    .Y(_1767_));
 sg13g2_nor2_1 _4887_ (.A(_1759_),
    .B(_1767_),
    .Y(_1768_));
 sg13g2_nand2_1 _4888_ (.Y(_1769_),
    .A(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[0] ),
    .B(_0212_));
 sg13g2_o21ai_1 _4889_ (.B1(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[0] ),
    .Y(_1770_),
    .A1(_1759_),
    .A2(_1767_));
 sg13g2_nor2b_1 _4890_ (.A(_1766_),
    .B_N(_1763_),
    .Y(_1771_));
 sg13g2_a22oi_1 _4891_ (.Y(_1772_),
    .B1(_1771_),
    .B2(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[1] ),
    .A2(_1769_),
    .A1(_1768_));
 sg13g2_nand3_1 _4892_ (.B(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[4] ),
    .C(_0941_),
    .A(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[2] ),
    .Y(_1773_));
 sg13g2_nor2_1 _4893_ (.A(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[1] ),
    .B(_1771_),
    .Y(_1774_));
 sg13g2_a221oi_1 _4894_ (.B2(_1740_),
    .C1(_1774_),
    .B1(_1773_),
    .A1(_1770_),
    .Y(_1775_),
    .A2(_1772_));
 sg13g2_nor3_1 _4895_ (.A(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[2] ),
    .B(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[4] ),
    .C(_0941_),
    .Y(_1776_));
 sg13g2_o21ai_1 _4896_ (.B1(net626),
    .Y(_1777_),
    .A1(_1740_),
    .A2(_1776_));
 sg13g2_nor3_1 _4897_ (.A(net900),
    .B(_1775_),
    .C(net627),
    .Y(_0329_));
 sg13g2_and3_1 _4898_ (.X(_1778_),
    .A(net609),
    .B(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[1] ),
    .C(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[2] ));
 sg13g2_and2_1 _4899_ (.A(net1463),
    .B(_1778_),
    .X(_1779_));
 sg13g2_nand2_1 _4900_ (.Y(_1780_),
    .A(net1713),
    .B(_1779_));
 sg13g2_o21ai_1 _4901_ (.B1(net947),
    .Y(_1781_),
    .A1(_0915_),
    .A2(_1780_));
 sg13g2_nor2_1 _4902_ (.A(_0954_),
    .B(_1781_),
    .Y(_0330_));
 sg13g2_xnor2_1 _4903_ (.Y(_1782_),
    .A(net609),
    .B(net612));
 sg13g2_nor2_1 _4904_ (.A(_1781_),
    .B(_1782_),
    .Y(_0331_));
 sg13g2_a21oi_1 _4905_ (.A1(net609),
    .A2(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[1] ),
    .Y(_1783_),
    .B1(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[2] ));
 sg13g2_nor3_1 _4906_ (.A(net900),
    .B(_1778_),
    .C(net610),
    .Y(_0332_));
 sg13g2_o21ai_1 _4907_ (.B1(net943),
    .Y(_1784_),
    .A1(net1463),
    .A2(_1778_));
 sg13g2_nor2_1 _4908_ (.A(_1779_),
    .B(net1464),
    .Y(_0333_));
 sg13g2_or2_1 _4909_ (.X(_1785_),
    .B(_1779_),
    .A(net1713));
 sg13g2_and3_1 _4910_ (.X(_0334_),
    .A(net947),
    .B(_1780_),
    .C(_1785_));
 sg13g2_a21oi_1 _4911_ (.A1(_0915_),
    .A2(_1780_),
    .Y(_0335_),
    .B1(_1781_));
 sg13g2_nand4_1 _4912_ (.B(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[2] ),
    .C(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[4] ),
    .A(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[1] ),
    .Y(_1786_),
    .D(_0955_));
 sg13g2_a21oi_2 _4913_ (.B1(_1604_),
    .Y(_1787_),
    .A2(_1447_),
    .A1(_0962_));
 sg13g2_a22oi_1 _4914_ (.Y(_1788_),
    .B1(_1603_),
    .B2(_0969_),
    .A2(_1447_),
    .A1(_0971_));
 sg13g2_nor2_1 _4915_ (.A(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[0] ),
    .B(_1788_),
    .Y(_1789_));
 sg13g2_a22oi_1 _4916_ (.Y(_1790_),
    .B1(_1787_),
    .B2(_1789_),
    .A2(_1786_),
    .A1(_1767_));
 sg13g2_nor3_1 _4917_ (.A(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[1] ),
    .B(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[2] ),
    .C(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[4] ),
    .Y(_1791_));
 sg13g2_a21oi_1 _4918_ (.A1(_0202_),
    .A2(_1791_),
    .Y(_1792_),
    .B1(_1767_));
 sg13g2_nand2_1 _4919_ (.Y(_1793_),
    .A(net948),
    .B(net653));
 sg13g2_nor3_1 _4920_ (.A(_1790_),
    .B(_1792_),
    .C(_1793_),
    .Y(_0336_));
 sg13g2_nor2_1 _4921_ (.A(\Led_Cycle_inst.buttons[1] ),
    .B(\Led_Cycle_inst.buttons[0] ),
    .Y(_1794_));
 sg13g2_and2_1 _4922_ (.A(\Led_Cycle_inst.buttons[2] ),
    .B(_0111_),
    .X(_1795_));
 sg13g2_nor3_1 _4923_ (.A(\Led_Cycle_inst.buttons[3] ),
    .B(\Led_Cycle_inst.buttons[1] ),
    .C(\Led_Cycle_inst.buttons[0] ),
    .Y(_1796_));
 sg13g2_nor2_1 _4924_ (.A(\Led_Cycle_inst.buttons[3] ),
    .B(\Led_Cycle_inst.buttons[2] ),
    .Y(_1797_));
 sg13g2_and2_1 _4925_ (.A(\Led_Cycle_inst.buttons[1] ),
    .B(_0111_),
    .X(_1798_));
 sg13g2_nor3_1 _4926_ (.A(\Led_Cycle_inst.buttons[3] ),
    .B(\Led_Cycle_inst.buttons[2] ),
    .C(\Led_Cycle_inst.buttons[0] ),
    .Y(_1799_));
 sg13g2_and2_1 _4927_ (.A(_1798_),
    .B(_1799_),
    .X(_1800_));
 sg13g2_a22oi_1 _4928_ (.Y(_1801_),
    .B1(_1798_),
    .B2(_1799_),
    .A2(_1796_),
    .A1(_1795_));
 sg13g2_xor2_1 _4929_ (.B(\Led_Cycle_inst.buttons[3] ),
    .A(\Led_Cycle_inst.buttons[4] ),
    .X(_1802_));
 sg13g2_nand3b_1 _4930_ (.B(_1794_),
    .C(_1802_),
    .Y(_1803_),
    .A_N(\Led_Cycle_inst.buttons[2] ));
 sg13g2_nor3_1 _4931_ (.A(\Led_Cycle_inst.buttons[3] ),
    .B(\Led_Cycle_inst.buttons[2] ),
    .C(_0111_),
    .Y(_1804_));
 sg13g2_and2_1 _4932_ (.A(_1794_),
    .B(_1804_),
    .X(_1805_));
 sg13g2_nand2_1 _4933_ (.Y(_1806_),
    .A(_1794_),
    .B(_1804_));
 sg13g2_nand2_2 _4934_ (.Y(_1807_),
    .A(_1801_),
    .B(_1803_));
 sg13g2_inv_1 _4935_ (.Y(_1808_),
    .A(_1807_));
 sg13g2_o21ai_1 _4936_ (.B1(_1801_),
    .Y(_1809_),
    .A1(_1803_),
    .A2(_1806_));
 sg13g2_xnor2_1 _4937_ (.Y(_1810_),
    .A(\Led_Cycle_inst.clk_reducer.counter[16] ),
    .B(_1809_));
 sg13g2_xor2_1 _4938_ (.B(_1807_),
    .A(\Led_Cycle_inst.clk_reducer.counter[22] ),
    .X(_1811_));
 sg13g2_nor4_2 _4939_ (.A(net1585),
    .B(net1511),
    .C(net1428),
    .Y(_1812_),
    .D(net1208));
 sg13g2_nor4_2 _4940_ (.A(net1599),
    .B(net1468),
    .C(net1453),
    .Y(_1813_),
    .D(net1433));
 sg13g2_nor4_2 _4941_ (.A(\Led_Cycle_inst.clk_reducer.counter[1] ),
    .B(\Led_Cycle_inst.clk_reducer.counter[0] ),
    .C(\Led_Cycle_inst.clk_reducer.counter[3] ),
    .Y(_1814_),
    .D(\Led_Cycle_inst.clk_reducer.counter[2] ));
 sg13g2_nor2_1 _4942_ (.A(\Led_Cycle_inst.clk_reducer.counter[5] ),
    .B(\Led_Cycle_inst.clk_reducer.counter[4] ),
    .Y(_1815_));
 sg13g2_nand3_1 _4943_ (.B(\Led_Cycle_inst.clk_reducer.counter[18] ),
    .C(_1815_),
    .A(\Led_Cycle_inst.clk_reducer.counter[19] ),
    .Y(_1816_));
 sg13g2_nor4_1 _4944_ (.A(\Led_Cycle_inst.clk_reducer.counter[13] ),
    .B(\Led_Cycle_inst.clk_reducer.counter[12] ),
    .C(\Led_Cycle_inst.clk_reducer.counter[23] ),
    .D(_1816_),
    .Y(_1817_));
 sg13g2_and4_1 _4945_ (.A(_1812_),
    .B(_1813_),
    .C(_1814_),
    .D(_1817_),
    .X(_1818_));
 sg13g2_xor2_1 _4946_ (.B(_1803_),
    .A(\Led_Cycle_inst.clk_reducer.counter[17] ),
    .X(_1819_));
 sg13g2_xor2_1 _4947_ (.B(_1801_),
    .A(\Led_Cycle_inst.clk_reducer.counter[21] ),
    .X(_1820_));
 sg13g2_nand4_1 _4948_ (.B(_1818_),
    .C(_1819_),
    .A(_1811_),
    .Y(_1821_),
    .D(_1820_));
 sg13g2_a21oi_2 _4949_ (.B1(_1797_),
    .Y(_1822_),
    .A2(_1803_),
    .A1(_1801_));
 sg13g2_or4_1 _4950_ (.A(\Led_Cycle_inst.clk_reducer.counter[7] ),
    .B(\Led_Cycle_inst.clk_reducer.counter[10] ),
    .C(\Led_Cycle_inst.clk_reducer.counter[15] ),
    .D(_1822_),
    .X(_1823_));
 sg13g2_nand4_1 _4951_ (.B(\Led_Cycle_inst.clk_reducer.counter[10] ),
    .C(\Led_Cycle_inst.clk_reducer.counter[15] ),
    .A(\Led_Cycle_inst.clk_reducer.counter[7] ),
    .Y(_1824_),
    .D(_1822_));
 sg13g2_o21ai_1 _4952_ (.B1(_1807_),
    .Y(_1825_),
    .A1(\Led_Cycle_inst.buttons[3] ),
    .A2(_1800_));
 sg13g2_xnor2_1 _4953_ (.Y(_1826_),
    .A(\Led_Cycle_inst.clk_reducer.counter[20] ),
    .B(_1825_));
 sg13g2_a21oi_1 _4954_ (.A1(_1823_),
    .A2(_1824_),
    .Y(_1827_),
    .B1(_1826_));
 sg13g2_a221oi_1 _4955_ (.B2(_1803_),
    .C1(_1805_),
    .B1(_1801_),
    .A1(_1795_),
    .Y(_1828_),
    .A2(_1796_));
 sg13g2_nor4_1 _4956_ (.A(_0110_),
    .B(_0113_),
    .C(_0115_),
    .D(_1828_),
    .Y(_1829_));
 sg13g2_nand4_1 _4957_ (.B(_0113_),
    .C(_0115_),
    .A(_0110_),
    .Y(_1830_),
    .D(_1828_));
 sg13g2_nand2b_1 _4958_ (.Y(_1831_),
    .B(_1830_),
    .A_N(_1829_));
 sg13g2_a21oi_2 _4959_ (.B1(_1800_),
    .Y(_1832_),
    .A2(_1803_),
    .A1(_1801_));
 sg13g2_or3_1 _4960_ (.A(_0112_),
    .B(_0114_),
    .C(_1832_),
    .X(_1833_));
 sg13g2_nand3_1 _4961_ (.B(_0114_),
    .C(_1832_),
    .A(_0112_),
    .Y(_1834_));
 sg13g2_a21oi_1 _4962_ (.A1(_1833_),
    .A2(_1834_),
    .Y(_1835_),
    .B1(_1821_));
 sg13g2_nand4_1 _4963_ (.B(_1827_),
    .C(_1831_),
    .A(_1810_),
    .Y(_1836_),
    .D(_1835_));
 sg13g2_nand2_1 _4964_ (.Y(_1837_),
    .A(net916),
    .B(_1836_));
 sg13g2_and3_1 _4965_ (.X(_0337_),
    .A(net916),
    .B(net637),
    .C(_1836_));
 sg13g2_xnor2_1 _4966_ (.Y(_1838_),
    .A(net1600),
    .B(\Led_Cycle_inst.clk_reducer.counter[0] ));
 sg13g2_nor2_1 _4967_ (.A(net725),
    .B(net1601),
    .Y(_0338_));
 sg13g2_and3_1 _4968_ (.X(_1839_),
    .A(\Led_Cycle_inst.clk_reducer.counter[1] ),
    .B(\Led_Cycle_inst.clk_reducer.counter[0] ),
    .C(net1309));
 sg13g2_a21oi_1 _4969_ (.A1(\Led_Cycle_inst.clk_reducer.counter[1] ),
    .A2(\Led_Cycle_inst.clk_reducer.counter[0] ),
    .Y(_1840_),
    .B1(net1309));
 sg13g2_nor3_1 _4970_ (.A(net725),
    .B(_1839_),
    .C(net1310),
    .Y(_0339_));
 sg13g2_and4_1 _4971_ (.A(\Led_Cycle_inst.clk_reducer.counter[1] ),
    .B(\Led_Cycle_inst.clk_reducer.counter[0] ),
    .C(net1388),
    .D(net1309),
    .X(_1841_));
 sg13g2_nor2_1 _4972_ (.A(net1388),
    .B(_1839_),
    .Y(_1842_));
 sg13g2_nor3_1 _4973_ (.A(net725),
    .B(_1841_),
    .C(net1389),
    .Y(_0340_));
 sg13g2_and2_1 _4974_ (.A(net1536),
    .B(_1841_),
    .X(_1843_));
 sg13g2_nor2_1 _4975_ (.A(net1536),
    .B(_1841_),
    .Y(_1844_));
 sg13g2_nor3_1 _4976_ (.A(net725),
    .B(_1843_),
    .C(net1537),
    .Y(_0341_));
 sg13g2_nand2_1 _4977_ (.Y(_1845_),
    .A(net1596),
    .B(_1843_));
 sg13g2_xnor2_1 _4978_ (.Y(_1846_),
    .A(net1596),
    .B(_1843_));
 sg13g2_nor2_1 _4979_ (.A(net725),
    .B(_1846_),
    .Y(_0342_));
 sg13g2_xor2_1 _4980_ (.B(_1845_),
    .A(net1589),
    .X(_1847_));
 sg13g2_nor2_1 _4981_ (.A(net726),
    .B(net1590),
    .Y(_0343_));
 sg13g2_nor2_1 _4982_ (.A(net1632),
    .B(_1845_),
    .Y(_1848_));
 sg13g2_xnor2_1 _4983_ (.Y(_1849_),
    .A(\Led_Cycle_inst.clk_reducer.counter[7] ),
    .B(_1848_));
 sg13g2_nor2_1 _4984_ (.A(net726),
    .B(net1633),
    .Y(_0344_));
 sg13g2_and2_1 _4985_ (.A(\Led_Cycle_inst.clk_reducer.counter[6] ),
    .B(\Led_Cycle_inst.clk_reducer.counter[7] ),
    .X(_1850_));
 sg13g2_nand4_1 _4986_ (.B(\Led_Cycle_inst.clk_reducer.counter[4] ),
    .C(_1841_),
    .A(\Led_Cycle_inst.clk_reducer.counter[5] ),
    .Y(_1851_),
    .D(_1850_));
 sg13g2_xnor2_1 _4987_ (.Y(_1852_),
    .A(net1701),
    .B(_1851_));
 sg13g2_nor2b_1 _4988_ (.A(net726),
    .B_N(_1852_),
    .Y(_0345_));
 sg13g2_nor2_1 _4989_ (.A(_0112_),
    .B(_1851_),
    .Y(_1853_));
 sg13g2_xnor2_1 _4990_ (.Y(_1854_),
    .A(net1398),
    .B(_1853_));
 sg13g2_nor2_1 _4991_ (.A(net729),
    .B(net1399),
    .Y(_0346_));
 sg13g2_nand2_2 _4992_ (.Y(_1855_),
    .A(net1781),
    .B(net1398));
 sg13g2_nor2_1 _4993_ (.A(_1851_),
    .B(_1855_),
    .Y(_1856_));
 sg13g2_nor3_2 _4994_ (.A(_0923_),
    .B(_1851_),
    .C(_1855_),
    .Y(_1857_));
 sg13g2_nor2_1 _4995_ (.A(net1613),
    .B(_1856_),
    .Y(_1858_));
 sg13g2_nor3_1 _4996_ (.A(net726),
    .B(_1857_),
    .C(net1614),
    .Y(_0347_));
 sg13g2_xnor2_1 _4997_ (.Y(_1859_),
    .A(net1550),
    .B(_1857_));
 sg13g2_nor2_1 _4998_ (.A(net726),
    .B(net1551),
    .Y(_0348_));
 sg13g2_nand2_1 _4999_ (.Y(_1860_),
    .A(net1550),
    .B(net1400));
 sg13g2_nor4_2 _5000_ (.A(_0923_),
    .B(_1851_),
    .C(_1855_),
    .Y(_1861_),
    .D(_1860_));
 sg13g2_a21oi_1 _5001_ (.A1(\Led_Cycle_inst.clk_reducer.counter[11] ),
    .A2(_1857_),
    .Y(_1862_),
    .B1(net1400));
 sg13g2_nor3_1 _5002_ (.A(net729),
    .B(_1861_),
    .C(net1401),
    .Y(_0349_));
 sg13g2_and2_1 _5003_ (.A(net1640),
    .B(_1861_),
    .X(_1863_));
 sg13g2_nor2_1 _5004_ (.A(net1640),
    .B(_1861_),
    .Y(_1864_));
 sg13g2_nor3_1 _5005_ (.A(net728),
    .B(_1863_),
    .C(net1641),
    .Y(_0350_));
 sg13g2_xnor2_1 _5006_ (.Y(_1865_),
    .A(net1543),
    .B(_1863_));
 sg13g2_nor2_1 _5007_ (.A(net729),
    .B(net1544),
    .Y(_0351_));
 sg13g2_nor2b_1 _5008_ (.A(_0115_),
    .B_N(_1863_),
    .Y(_1866_));
 sg13g2_xnor2_1 _5009_ (.Y(_1867_),
    .A(net1503),
    .B(_1866_));
 sg13g2_nor2_1 _5010_ (.A(net726),
    .B(net1504),
    .Y(_0352_));
 sg13g2_and4_2 _5011_ (.A(\Led_Cycle_inst.clk_reducer.counter[13] ),
    .B(net1543),
    .C(net1503),
    .D(_1861_),
    .X(_1868_));
 sg13g2_nor2_1 _5012_ (.A(net1642),
    .B(_1868_),
    .Y(_1869_));
 sg13g2_and2_1 _5013_ (.A(net1642),
    .B(_1868_),
    .X(_1870_));
 sg13g2_nor3_1 _5014_ (.A(net728),
    .B(_1869_),
    .C(_1870_),
    .Y(_0353_));
 sg13g2_or2_1 _5015_ (.X(_1871_),
    .B(_1870_),
    .A(net1745));
 sg13g2_nand3_1 _5016_ (.B(\Led_Cycle_inst.clk_reducer.counter[17] ),
    .C(_1868_),
    .A(\Led_Cycle_inst.clk_reducer.counter[16] ),
    .Y(_1872_));
 sg13g2_and4_1 _5017_ (.A(net923),
    .B(_1836_),
    .C(_1871_),
    .D(_1872_),
    .X(_0354_));
 sg13g2_xnor2_1 _5018_ (.Y(_1873_),
    .A(net1665),
    .B(_1872_));
 sg13g2_nor2b_1 _5019_ (.A(net728),
    .B_N(net1666),
    .Y(_0355_));
 sg13g2_nor2_1 _5020_ (.A(net1244),
    .B(_1872_),
    .Y(_1874_));
 sg13g2_xnor2_1 _5021_ (.Y(_1875_),
    .A(\Led_Cycle_inst.clk_reducer.counter[19] ),
    .B(_1874_));
 sg13g2_nor2_1 _5022_ (.A(net728),
    .B(net1245),
    .Y(_0356_));
 sg13g2_and4_1 _5023_ (.A(\Led_Cycle_inst.clk_reducer.counter[16] ),
    .B(\Led_Cycle_inst.clk_reducer.counter[17] ),
    .C(\Led_Cycle_inst.clk_reducer.counter[19] ),
    .D(\Led_Cycle_inst.clk_reducer.counter[18] ),
    .X(_1876_));
 sg13g2_a21oi_1 _5024_ (.A1(_1868_),
    .A2(_1876_),
    .Y(_1877_),
    .B1(net1525));
 sg13g2_and3_1 _5025_ (.X(_1878_),
    .A(net1525),
    .B(_1868_),
    .C(_1876_));
 sg13g2_nor3_1 _5026_ (.A(net727),
    .B(net1526),
    .C(_1878_),
    .Y(_0357_));
 sg13g2_nor2_1 _5027_ (.A(net1631),
    .B(_1878_),
    .Y(_1879_));
 sg13g2_and4_2 _5028_ (.A(net1525),
    .B(\Led_Cycle_inst.clk_reducer.counter[21] ),
    .C(_1868_),
    .D(_1876_),
    .X(_1880_));
 sg13g2_nor3_1 _5029_ (.A(net727),
    .B(_1879_),
    .C(_1880_),
    .Y(_0358_));
 sg13g2_xnor2_1 _5030_ (.Y(_1881_),
    .A(net1692),
    .B(_1880_));
 sg13g2_nor2_1 _5031_ (.A(net727),
    .B(_1881_),
    .Y(_0359_));
 sg13g2_a21oi_1 _5032_ (.A1(net1692),
    .A2(_1880_),
    .Y(_1882_),
    .B1(net1680));
 sg13g2_nand3_1 _5033_ (.B(net1680),
    .C(_1880_),
    .A(net1692),
    .Y(_1883_));
 sg13g2_nor2_1 _5034_ (.A(net727),
    .B(_1882_),
    .Y(_1884_));
 sg13g2_and2_1 _5035_ (.A(_1883_),
    .B(_1884_),
    .X(_0360_));
 sg13g2_nor2b_1 _5036_ (.A(net1468),
    .B_N(_1883_),
    .Y(_1885_));
 sg13g2_and4_2 _5037_ (.A(net1777),
    .B(net1774),
    .C(net1468),
    .D(_1880_),
    .X(_1886_));
 sg13g2_nor3_1 _5038_ (.A(net727),
    .B(net1469),
    .C(_1886_),
    .Y(_0361_));
 sg13g2_xnor2_1 _5039_ (.Y(_1887_),
    .A(net1599),
    .B(net1775));
 sg13g2_nor2_1 _5040_ (.A(net727),
    .B(_1887_),
    .Y(_0362_));
 sg13g2_a21oi_1 _5041_ (.A1(\Led_Cycle_inst.clk_reducer.counter[25] ),
    .A2(_1886_),
    .Y(_1888_),
    .B1(net1433));
 sg13g2_and3_1 _5042_ (.X(_1889_),
    .A(\Led_Cycle_inst.clk_reducer.counter[25] ),
    .B(net1433),
    .C(_1886_));
 sg13g2_nor3_1 _5043_ (.A(net727),
    .B(net1434),
    .C(_1889_),
    .Y(_0363_));
 sg13g2_nor2_1 _5044_ (.A(net1453),
    .B(_1889_),
    .Y(_1890_));
 sg13g2_and4_1 _5045_ (.A(net1778),
    .B(net1453),
    .C(net1433),
    .D(_1886_),
    .X(_1891_));
 sg13g2_nor3_1 _5046_ (.A(net727),
    .B(net1454),
    .C(_1891_),
    .Y(_0364_));
 sg13g2_nor2_1 _5047_ (.A(net1511),
    .B(_1891_),
    .Y(_1892_));
 sg13g2_and2_1 _5048_ (.A(net1511),
    .B(_1891_),
    .X(_1893_));
 sg13g2_nor3_1 _5049_ (.A(net726),
    .B(net1512),
    .C(_1893_),
    .Y(_0365_));
 sg13g2_nor2_1 _5050_ (.A(net1585),
    .B(_1893_),
    .Y(_1894_));
 sg13g2_a21oi_1 _5051_ (.A1(net1585),
    .A2(_1893_),
    .Y(_1895_),
    .B1(net725));
 sg13g2_nor2b_1 _5052_ (.A(_1894_),
    .B_N(_1895_),
    .Y(_0366_));
 sg13g2_a21oi_1 _5053_ (.A1(\Led_Cycle_inst.clk_reducer.counter[29] ),
    .A2(_1893_),
    .Y(_1896_),
    .B1(net1208));
 sg13g2_and4_1 _5054_ (.A(\Led_Cycle_inst.clk_reducer.counter[29] ),
    .B(\Led_Cycle_inst.clk_reducer.counter[28] ),
    .C(net1208),
    .D(_1891_),
    .X(_1897_));
 sg13g2_nor3_1 _5055_ (.A(net725),
    .B(net1209),
    .C(_1897_),
    .Y(_0367_));
 sg13g2_xnor2_1 _5056_ (.Y(_1898_),
    .A(net1428),
    .B(_1897_));
 sg13g2_nor2_1 _5057_ (.A(net725),
    .B(net1429),
    .Y(_0368_));
 sg13g2_nor3_1 _5058_ (.A(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[0] ),
    .B(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[2] ),
    .C(net667),
    .Y(_1899_));
 sg13g2_nand3_1 _5059_ (.B(_0185_),
    .C(_1899_),
    .A(_0184_),
    .Y(_1900_));
 sg13g2_a21oi_1 _5060_ (.A1(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[4] ),
    .A2(_1900_),
    .Y(_1901_),
    .B1(_1787_));
 sg13g2_a22oi_1 _5061_ (.Y(_1902_),
    .B1(_1603_),
    .B2(_0962_),
    .A2(_1453_),
    .A1(_1447_));
 sg13g2_o21ai_1 _5062_ (.B1(_1902_),
    .Y(_1903_),
    .A1(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[4] ),
    .A2(_1900_));
 sg13g2_nor2_1 _5063_ (.A(_1901_),
    .B(_1903_),
    .Y(_1904_));
 sg13g2_nor3_1 _5064_ (.A(_0184_),
    .B(_0185_),
    .C(net667),
    .Y(_1905_));
 sg13g2_nand3_1 _5065_ (.B(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[4] ),
    .C(_1905_),
    .A(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[2] ),
    .Y(_1906_));
 sg13g2_nand3_1 _5066_ (.B(net677),
    .C(_1906_),
    .A(net948),
    .Y(_1907_));
 sg13g2_nor2_1 _5067_ (.A(_1904_),
    .B(net678),
    .Y(_0369_));
 sg13g2_nor2_1 _5068_ (.A(\Led_Cycle_inst.clk_reducer.counter[20] ),
    .B(_1801_),
    .Y(_1908_));
 sg13g2_nor3_1 _5069_ (.A(\Led_Cycle_inst.clk_reducer.counter[21] ),
    .B(net1777),
    .C(net1680),
    .Y(_1909_));
 sg13g2_o21ai_1 _5070_ (.B1(_1909_),
    .Y(_1910_),
    .A1(_1808_),
    .A2(_1908_));
 sg13g2_nand2_1 _5071_ (.Y(_1911_),
    .A(\Led_Cycle_inst.clk_reducer.counter[20] ),
    .B(_1801_));
 sg13g2_nor3_1 _5072_ (.A(\Led_Cycle_inst.clk_reducer.counter[22] ),
    .B(\Led_Cycle_inst.clk_reducer.counter[23] ),
    .C(_1908_),
    .Y(_1912_));
 sg13g2_xor2_1 _5073_ (.B(_1807_),
    .A(\Led_Cycle_inst.clk_reducer.counter[21] ),
    .X(_1913_));
 sg13g2_nand3_1 _5074_ (.B(_1912_),
    .C(_1913_),
    .A(_1911_),
    .Y(_1914_));
 sg13g2_inv_1 _5075_ (.Y(_1915_),
    .A(_1914_));
 sg13g2_xnor2_1 _5076_ (.Y(_1916_),
    .A(\Led_Cycle_inst.clk_reducer.counter[14] ),
    .B(_1822_));
 sg13g2_nor2_1 _5077_ (.A(_0181_),
    .B(_1809_),
    .Y(_1917_));
 sg13g2_xor2_1 _5078_ (.B(_1809_),
    .A(_0181_),
    .X(_1918_));
 sg13g2_nand2_1 _5079_ (.Y(_1919_),
    .A(\Led_Cycle_inst.clk_reducer.counter[19] ),
    .B(_1825_));
 sg13g2_nor2_1 _5080_ (.A(\Led_Cycle_inst.clk_reducer.counter[19] ),
    .B(_1825_),
    .Y(_1920_));
 sg13g2_nand3b_1 _5081_ (.B(\Led_Cycle_inst.clk_reducer.counter[18] ),
    .C(_1919_),
    .Y(_1921_),
    .A_N(_1920_));
 sg13g2_o21ai_1 _5082_ (.B1(\Led_Cycle_inst.clk_reducer.counter[17] ),
    .Y(_1922_),
    .A1(\Led_Cycle_inst.clk_reducer.counter[16] ),
    .A2(_1803_));
 sg13g2_a21o_1 _5083_ (.A2(_1803_),
    .A1(\Led_Cycle_inst.clk_reducer.counter[16] ),
    .B1(_1922_),
    .X(_1923_));
 sg13g2_nor2_1 _5084_ (.A(\Led_Cycle_inst.clk_reducer.counter[13] ),
    .B(_1828_),
    .Y(_1924_));
 sg13g2_xor2_1 _5085_ (.B(_1828_),
    .A(\Led_Cycle_inst.clk_reducer.counter[13] ),
    .X(_1925_));
 sg13g2_nand3_1 _5086_ (.B(_1918_),
    .C(_1925_),
    .A(_1916_),
    .Y(_1926_));
 sg13g2_nor4_1 _5087_ (.A(\Led_Cycle_inst.clk_reducer.counter[12] ),
    .B(_1921_),
    .C(_1923_),
    .D(_1926_),
    .Y(_1927_));
 sg13g2_o21ai_1 _5088_ (.B1(_0114_),
    .Y(_1928_),
    .A1(_0113_),
    .A2(_1822_));
 sg13g2_xnor2_1 _5089_ (.Y(_1929_),
    .A(\Led_Cycle_inst.clk_reducer.counter[10] ),
    .B(_1832_));
 sg13g2_nor2_1 _5090_ (.A(_1928_),
    .B(_1929_),
    .Y(_1930_));
 sg13g2_nor2_1 _5091_ (.A(\Led_Cycle_inst.clk_reducer.counter[8] ),
    .B(_1828_),
    .Y(_1931_));
 sg13g2_nand2_1 _5092_ (.Y(_1932_),
    .A(_0113_),
    .B(_1822_));
 sg13g2_nor2b_1 _5093_ (.A(_1931_),
    .B_N(_1932_),
    .Y(_1933_));
 sg13g2_nand2b_1 _5094_ (.Y(_1934_),
    .B(_1932_),
    .A_N(_1931_));
 sg13g2_nand2_1 _5095_ (.Y(_1935_),
    .A(\Led_Cycle_inst.clk_reducer.counter[8] ),
    .B(_1828_));
 sg13g2_nand3_1 _5096_ (.B(_1933_),
    .C(_1935_),
    .A(_1930_),
    .Y(_1936_));
 sg13g2_nor2b_1 _5097_ (.A(_1828_),
    .B_N(_0182_),
    .Y(_1937_));
 sg13g2_nand2_1 _5098_ (.Y(_1938_),
    .A(\Led_Cycle_inst.clk_reducer.counter[7] ),
    .B(_1832_));
 sg13g2_or2_1 _5099_ (.X(_1939_),
    .B(_1832_),
    .A(\Led_Cycle_inst.clk_reducer.counter[7] ));
 sg13g2_xnor2_1 _5100_ (.Y(_1940_),
    .A(\Led_Cycle_inst.clk_reducer.counter[6] ),
    .B(_1822_));
 sg13g2_and3_1 _5101_ (.X(_1941_),
    .A(_1938_),
    .B(_1939_),
    .C(_1940_));
 sg13g2_nand2_1 _5102_ (.Y(_1942_),
    .A(_0110_),
    .B(_1822_));
 sg13g2_nand2_1 _5103_ (.Y(_1943_),
    .A(_1939_),
    .B(_1942_));
 sg13g2_a22oi_1 _5104_ (.Y(_1944_),
    .B1(_1943_),
    .B2(_1938_),
    .A2(_1941_),
    .A1(_1937_));
 sg13g2_nor3_1 _5105_ (.A(\Led_Cycle_inst.clk_reducer.counter[10] ),
    .B(\Led_Cycle_inst.clk_reducer.counter[11] ),
    .C(_1832_),
    .Y(_1945_));
 sg13g2_a21oi_1 _5106_ (.A1(_1930_),
    .A2(_1934_),
    .Y(_1946_),
    .B1(_1945_));
 sg13g2_o21ai_1 _5107_ (.B1(_1946_),
    .Y(_1947_),
    .A1(_1936_),
    .A2(_1944_));
 sg13g2_and2_1 _5108_ (.A(_1927_),
    .B(_1947_),
    .X(_1948_));
 sg13g2_o21ai_1 _5109_ (.B1(_1919_),
    .Y(_1949_),
    .A1(_0180_),
    .A2(_1920_));
 sg13g2_nand3_1 _5110_ (.B(_1918_),
    .C(_1924_),
    .A(_1916_),
    .Y(_1950_));
 sg13g2_a22oi_1 _5111_ (.Y(_1951_),
    .B1(_1822_),
    .B2(_0115_),
    .A2(_1809_),
    .A1(_0181_));
 sg13g2_or2_1 _5112_ (.X(_1952_),
    .B(_1951_),
    .A(_1917_));
 sg13g2_a21oi_1 _5113_ (.A1(_1950_),
    .A2(_1952_),
    .Y(_1953_),
    .B1(_1923_));
 sg13g2_nor2_1 _5114_ (.A(_1922_),
    .B(_1953_),
    .Y(_1954_));
 sg13g2_o21ai_1 _5115_ (.B1(_1949_),
    .Y(_1955_),
    .A1(_1921_),
    .A2(_1954_));
 sg13g2_o21ai_1 _5116_ (.B1(_1915_),
    .Y(_1956_),
    .A1(_1948_),
    .A2(_1955_));
 sg13g2_nor2b_1 _5117_ (.A(_0182_),
    .B_N(_1828_),
    .Y(_1957_));
 sg13g2_nand2b_1 _5118_ (.Y(_1958_),
    .B(_1814_),
    .A_N(\Led_Cycle_inst.clk_reducer.counter[4] ));
 sg13g2_nor3_1 _5119_ (.A(_1937_),
    .B(_1957_),
    .C(_1958_),
    .Y(_1959_));
 sg13g2_nand3_1 _5120_ (.B(_1941_),
    .C(_1959_),
    .A(_1915_),
    .Y(_1960_));
 sg13g2_nor2_1 _5121_ (.A(_1936_),
    .B(_1960_),
    .Y(_1961_));
 sg13g2_nand3_1 _5122_ (.B(_1812_),
    .C(_1813_),
    .A(net918),
    .Y(_1962_));
 sg13g2_a221oi_1 _5123_ (.B2(_1927_),
    .C1(_1962_),
    .B1(_1961_),
    .A1(_1910_),
    .Y(_0370_),
    .A2(_1956_));
 sg13g2_nor3_1 _5124_ (.A(_1360_),
    .B(net1676),
    .C(_0701_),
    .Y(_0371_));
 sg13g2_and3_1 _5125_ (.X(_0380_),
    .A(net939),
    .B(net829),
    .C(_1235_));
 sg13g2_and3_1 _5126_ (.X(_0381_),
    .A(net939),
    .B(net827),
    .C(_1230_));
 sg13g2_and3_1 _5127_ (.X(_0382_),
    .A(net939),
    .B(_1229_),
    .C(_1237_));
 sg13g2_or4_1 _5128_ (.A(net913),
    .B(rx_valid),
    .C(net1144),
    .D(_0978_),
    .X(_1963_));
 sg13g2_o21ai_1 _5129_ (.B1(net936),
    .Y(_1964_),
    .A1(net709),
    .A2(net787));
 sg13g2_a21oi_1 _5130_ (.A1(_0832_),
    .A2(net787),
    .Y(_0383_),
    .B1(_1964_));
 sg13g2_o21ai_1 _5131_ (.B1(net936),
    .Y(_1965_),
    .A1(\uart_inst.uart_rx_inst.DATA_TEMP_REG[1] ),
    .A2(net787));
 sg13g2_a21oi_1 _5132_ (.A1(_0830_),
    .A2(net787),
    .Y(_0384_),
    .B1(_1965_));
 sg13g2_o21ai_1 _5133_ (.B1(net934),
    .Y(_1966_),
    .A1(\uart_inst.uart_rx_inst.DATA_TEMP_REG[2] ),
    .A2(net786));
 sg13g2_a21oi_1 _5134_ (.A1(_0828_),
    .A2(net786),
    .Y(_0385_),
    .B1(_1966_));
 sg13g2_o21ai_1 _5135_ (.B1(net935),
    .Y(_1967_),
    .A1(net1038),
    .A2(net786));
 sg13g2_a21oi_1 _5136_ (.A1(_0826_),
    .A2(net786),
    .Y(_0386_),
    .B1(_1967_));
 sg13g2_o21ai_1 _5137_ (.B1(net934),
    .Y(_1968_),
    .A1(net1138),
    .A2(net785));
 sg13g2_a21oi_1 _5138_ (.A1(_0825_),
    .A2(net785),
    .Y(_0387_),
    .B1(_1968_));
 sg13g2_o21ai_1 _5139_ (.B1(net934),
    .Y(_1969_),
    .A1(net1092),
    .A2(net785));
 sg13g2_a21oi_1 _5140_ (.A1(_0824_),
    .A2(net785),
    .Y(_0388_),
    .B1(_1969_));
 sg13g2_o21ai_1 _5141_ (.B1(net934),
    .Y(_1970_),
    .A1(net1072),
    .A2(net785));
 sg13g2_a21oi_1 _5142_ (.A1(_0823_),
    .A2(net785),
    .Y(_0389_),
    .B1(_1970_));
 sg13g2_o21ai_1 _5143_ (.B1(net933),
    .Y(_1971_),
    .A1(net1111),
    .A2(net785));
 sg13g2_a21oi_1 _5144_ (.A1(_0822_),
    .A2(net785),
    .Y(_0390_),
    .B1(_1971_));
 sg13g2_o21ai_1 _5145_ (.B1(net1301),
    .Y(_1972_),
    .A1(net913),
    .A2(_0913_));
 sg13g2_a21oi_1 _5146_ (.A1(net787),
    .A2(_1972_),
    .Y(_0391_),
    .B1(net893));
 sg13g2_nand2_1 _5147_ (.Y(_1973_),
    .A(net890),
    .B(_0979_));
 sg13g2_o21ai_1 _5148_ (.B1(net936),
    .Y(_1974_),
    .A1(\uart_inst.uart_rx_inst.DATA_TEMP_REG[1] ),
    .A2(net768));
 sg13g2_a21oi_1 _5149_ (.A1(_0890_),
    .A2(net768),
    .Y(_0392_),
    .B1(_1974_));
 sg13g2_o21ai_1 _5150_ (.B1(net934),
    .Y(_1975_),
    .A1(\uart_inst.uart_rx_inst.DATA_TEMP_REG[2] ),
    .A2(net767));
 sg13g2_a21oi_1 _5151_ (.A1(_0889_),
    .A2(net767),
    .Y(_0393_),
    .B1(_1975_));
 sg13g2_o21ai_1 _5152_ (.B1(net935),
    .Y(_1976_),
    .A1(net1038),
    .A2(net767));
 sg13g2_a21oi_1 _5153_ (.A1(_0888_),
    .A2(net767),
    .Y(_0394_),
    .B1(_1976_));
 sg13g2_o21ai_1 _5154_ (.B1(net933),
    .Y(_1977_),
    .A1(net1138),
    .A2(net766));
 sg13g2_a21oi_1 _5155_ (.A1(_0887_),
    .A2(net766),
    .Y(_0395_),
    .B1(_1977_));
 sg13g2_o21ai_1 _5156_ (.B1(net933),
    .Y(_1978_),
    .A1(net1092),
    .A2(net766));
 sg13g2_a21oi_1 _5157_ (.A1(_0886_),
    .A2(net766),
    .Y(_0396_),
    .B1(_1978_));
 sg13g2_o21ai_1 _5158_ (.B1(net933),
    .Y(_1979_),
    .A1(net1072),
    .A2(net766));
 sg13g2_a21oi_1 _5159_ (.A1(_0885_),
    .A2(net766),
    .Y(_0397_),
    .B1(_1979_));
 sg13g2_o21ai_1 _5160_ (.B1(net933),
    .Y(_1980_),
    .A1(\uart_inst.uart_rx_inst.DATA_TEMP_REG[7] ),
    .A2(net766));
 sg13g2_a21oi_1 _5161_ (.A1(_0884_),
    .A2(net766),
    .Y(_0398_),
    .B1(_1980_));
 sg13g2_a22oi_1 _5162_ (.Y(_1981_),
    .B1(net768),
    .B2(net1111),
    .A2(_1010_),
    .A1(net890));
 sg13g2_nor2_1 _5163_ (.A(net893),
    .B(_1981_),
    .Y(_0399_));
 sg13g2_a21oi_1 _5164_ (.A1(\uart_inst.uart_rx_inst.SIGNAL_R ),
    .A2(\uart_inst.uart_rx_inst.state[0] ),
    .Y(_1982_),
    .B1(net913));
 sg13g2_o21ai_1 _5165_ (.B1(_1982_),
    .Y(_1983_),
    .A1(net890),
    .A2(\uart_inst.uart_rx_inst.state[0] ));
 sg13g2_nor2_1 _5166_ (.A(net890),
    .B(_1983_),
    .Y(_1984_));
 sg13g2_nor3_1 _5167_ (.A(_0978_),
    .B(_0981_),
    .C(_1983_),
    .Y(_1985_));
 sg13g2_nor2_1 _5168_ (.A(_1984_),
    .B(_1985_),
    .Y(_1986_));
 sg13g2_nor2b_1 _5169_ (.A(_1986_),
    .B_N(net1280),
    .Y(_1987_));
 sg13g2_o21ai_1 _5170_ (.B1(net936),
    .Y(_1988_),
    .A1(net890),
    .A2(_1983_));
 sg13g2_nor2_1 _5171_ (.A(net1280),
    .B(_1985_),
    .Y(_1989_));
 sg13g2_nor3_1 _5172_ (.A(_1987_),
    .B(_1988_),
    .C(_1989_),
    .Y(_0400_));
 sg13g2_nor2_1 _5173_ (.A(net1387),
    .B(_1987_),
    .Y(_1990_));
 sg13g2_and2_1 _5174_ (.A(net1387),
    .B(_1987_),
    .X(_1991_));
 sg13g2_nor3_1 _5175_ (.A(_1988_),
    .B(_1990_),
    .C(_1991_),
    .Y(_0401_));
 sg13g2_a21oi_1 _5176_ (.A1(net1500),
    .A2(_1991_),
    .Y(_1992_),
    .B1(_1988_));
 sg13g2_o21ai_1 _5177_ (.B1(_1992_),
    .Y(_1993_),
    .A1(net1500),
    .A2(_1991_));
 sg13g2_inv_1 _5178_ (.Y(_0402_),
    .A(_1993_));
 sg13g2_and2_1 _5179_ (.A(net680),
    .B(_1992_),
    .X(_0403_));
 sg13g2_o21ai_1 _5180_ (.B1(_1982_),
    .Y(_1994_),
    .A1(net1144),
    .A2(_0978_));
 sg13g2_nor2_2 _5181_ (.A(net1173),
    .B(net1776),
    .Y(_1995_));
 sg13g2_nor2_1 _5182_ (.A(_1994_),
    .B(_1995_),
    .Y(_1996_));
 sg13g2_o21ai_1 _5183_ (.B1(_0883_),
    .Y(_1997_),
    .A1(\uart_inst.uart_rx_inst.state[2] ),
    .A2(_0978_));
 sg13g2_nand2b_1 _5184_ (.Y(_1998_),
    .B(_1995_),
    .A_N(\uart_inst.uart_rx_inst.state[0] ));
 sg13g2_nand2b_1 _5185_ (.Y(_1999_),
    .B(_1998_),
    .A_N(_1994_));
 sg13g2_inv_1 _5186_ (.Y(_2000_),
    .A(net765));
 sg13g2_a221oi_1 _5187_ (.B2(_0883_),
    .C1(net898),
    .B1(net765),
    .A1(_1996_),
    .Y(_0404_),
    .A2(_1997_));
 sg13g2_o21ai_1 _5188_ (.B1(net1331),
    .Y(_2001_),
    .A1(\uart_inst.uart_rx_inst.CLK_CNT[0] ),
    .A2(_1999_));
 sg13g2_o21ai_1 _5189_ (.B1(_2000_),
    .Y(_2002_),
    .A1(_0973_),
    .A2(_1995_));
 sg13g2_a21oi_1 _5190_ (.A1(net1332),
    .A2(_2002_),
    .Y(_0405_),
    .B1(net898));
 sg13g2_nand2_1 _5191_ (.Y(_2003_),
    .A(_0126_),
    .B(_0973_));
 sg13g2_xor2_1 _5192_ (.B(_0973_),
    .A(_0126_),
    .X(_2004_));
 sg13g2_nor2_1 _5193_ (.A(net1144),
    .B(_1995_),
    .Y(_2005_));
 sg13g2_or2_1 _5194_ (.X(_2006_),
    .B(_2005_),
    .A(net890));
 sg13g2_a21oi_1 _5195_ (.A1(net890),
    .A2(_0978_),
    .Y(_2007_),
    .B1(_2005_));
 sg13g2_o21ai_1 _5196_ (.B1(_2000_),
    .Y(_2008_),
    .A1(_2004_),
    .A2(_2007_));
 sg13g2_o21ai_1 _5197_ (.B1(net942),
    .Y(_2009_),
    .A1(net1501),
    .A2(_2000_));
 sg13g2_nor2b_1 _5198_ (.A(_2009_),
    .B_N(_2008_),
    .Y(_0406_));
 sg13g2_xnor2_1 _5199_ (.Y(_2010_),
    .A(net1620),
    .B(_2003_));
 sg13g2_o21ai_1 _5200_ (.B1(_2010_),
    .Y(_2011_),
    .A1(net1598),
    .A2(_0978_));
 sg13g2_o21ai_1 _5201_ (.B1(net940),
    .Y(_2012_),
    .A1(net1620),
    .A2(_2000_));
 sg13g2_a21oi_1 _5202_ (.A1(_1996_),
    .A2(_2011_),
    .Y(_0407_),
    .B1(_2012_));
 sg13g2_o21ai_1 _5203_ (.B1(net941),
    .Y(_2013_),
    .A1(net765),
    .A2(_2006_));
 sg13g2_nor3_1 _5204_ (.A(net1684),
    .B(_0974_),
    .C(net765),
    .Y(_2014_));
 sg13g2_o21ai_1 _5205_ (.B1(net1684),
    .Y(_2015_),
    .A1(_0974_),
    .A2(net765));
 sg13g2_nor2b_1 _5206_ (.A(_2014_),
    .B_N(_2015_),
    .Y(_2016_));
 sg13g2_nor2_1 _5207_ (.A(_2013_),
    .B(_2016_),
    .Y(_0408_));
 sg13g2_xnor2_1 _5208_ (.Y(_2017_),
    .A(net1449),
    .B(_2014_));
 sg13g2_nor2_1 _5209_ (.A(_2013_),
    .B(net1450),
    .Y(_0409_));
 sg13g2_or2_1 _5210_ (.X(_2018_),
    .B(net765),
    .A(_0976_));
 sg13g2_a21oi_1 _5211_ (.A1(net1103),
    .A2(net1784),
    .Y(_2019_),
    .B1(_2007_));
 sg13g2_o21ai_1 _5212_ (.B1(net941),
    .Y(_2020_),
    .A1(net765),
    .A2(_2019_));
 sg13g2_a21oi_1 _5213_ (.A1(_0882_),
    .A2(_2018_),
    .Y(_0410_),
    .B1(_2020_));
 sg13g2_or2_1 _5214_ (.X(_2021_),
    .B(_2018_),
    .A(net1584));
 sg13g2_a22oi_1 _5215_ (.Y(_2022_),
    .B1(_2018_),
    .B2(net1584),
    .A2(_2000_),
    .A1(_1995_));
 sg13g2_a21oi_1 _5216_ (.A1(_2021_),
    .A2(_2022_),
    .Y(_0411_),
    .B1(net893));
 sg13g2_xor2_1 _5217_ (.B(_2021_),
    .A(net1615),
    .X(_2023_));
 sg13g2_nor2_1 _5218_ (.A(_2013_),
    .B(_2023_),
    .Y(_0412_));
 sg13g2_o21ai_1 _5219_ (.B1(net1430),
    .Y(_2024_),
    .A1(\uart_inst.uart_rx_inst.CLK_CNT[8] ),
    .A2(_2021_));
 sg13g2_a21oi_1 _5220_ (.A1(\uart_inst.uart_rx_inst.state[2] ),
    .A2(_0977_),
    .Y(_2025_),
    .B1(_1995_));
 sg13g2_or2_1 _5221_ (.X(_2026_),
    .B(_2025_),
    .A(net765));
 sg13g2_a21oi_1 _5222_ (.A1(net1431),
    .A2(_2026_),
    .Y(_0413_),
    .B1(net893));
 sg13g2_nor2_1 _5223_ (.A(net962),
    .B(net908),
    .Y(_2027_));
 sg13g2_a22oi_1 _5224_ (.Y(_2028_),
    .B1(net872),
    .B2(\uart_inst.uart_rx_inst.SAMPLING_COUNT[0] ),
    .A2(_0984_),
    .A1(net657));
 sg13g2_inv_1 _5225_ (.Y(_0414_),
    .A(net658));
 sg13g2_a21oi_1 _5226_ (.A1(net962),
    .A2(\uart_inst.uart_rx_inst.SAMPLING_COUNT[0] ),
    .Y(_2029_),
    .B1(net1254));
 sg13g2_and3_1 _5227_ (.X(_2030_),
    .A(net962),
    .B(net1254),
    .C(\uart_inst.uart_rx_inst.SAMPLING_COUNT[0] ));
 sg13g2_nor3_1 _5228_ (.A(net896),
    .B(net1255),
    .C(_2030_),
    .Y(_0415_));
 sg13g2_nor3_2 _5229_ (.A(net914),
    .B(net1254),
    .C(\uart_inst.uart_rx_inst.SAMPLING_COUNT[0] ),
    .Y(_2031_));
 sg13g2_a21oi_1 _5230_ (.A1(net1383),
    .A2(net871),
    .Y(_2032_),
    .B1(net896));
 sg13g2_o21ai_1 _5231_ (.B1(_2032_),
    .Y(_0416_),
    .A1(_0881_),
    .A2(net871));
 sg13g2_a21oi_1 _5232_ (.A1(\uart_inst.uart_rx_inst.SIGNAL_Q[2] ),
    .A2(net871),
    .Y(_2033_),
    .B1(net897));
 sg13g2_o21ai_1 _5233_ (.B1(_2033_),
    .Y(_0417_),
    .A1(_0880_),
    .A2(net871));
 sg13g2_a21oi_1 _5234_ (.A1(\uart_inst.uart_rx_inst.SIGNAL_Q[3] ),
    .A2(net871),
    .Y(_2034_),
    .B1(net897));
 sg13g2_o21ai_1 _5235_ (.B1(_2034_),
    .Y(_0418_),
    .A1(_0879_),
    .A2(net871));
 sg13g2_a21oi_1 _5236_ (.A1(net1552),
    .A2(_2031_),
    .Y(_2035_),
    .B1(net897));
 sg13g2_o21ai_1 _5237_ (.B1(_2035_),
    .Y(_0419_),
    .A1(_0878_),
    .A2(_2031_));
 sg13g2_a21oi_1 _5238_ (.A1(net1),
    .A2(net871),
    .Y(_2036_),
    .B1(net897));
 sg13g2_o21ai_1 _5239_ (.B1(_2036_),
    .Y(_0420_),
    .A1(_0877_),
    .A2(net871));
 sg13g2_nor3_1 _5240_ (.A(_1218_),
    .B(_1219_),
    .C(_0705_),
    .Y(_0421_));
 sg13g2_nor2_1 _5241_ (.A(\uart_inst.uart_tx_inst.state[0] ),
    .B(\uart_inst.uart_tx_inst.state[1] ),
    .Y(_2037_));
 sg13g2_a21oi_1 _5242_ (.A1(\uart_inst.uart_tx_inst.state[1] ),
    .A2(_0998_),
    .Y(_2038_),
    .B1(_2037_));
 sg13g2_and3_1 _5243_ (.X(_2039_),
    .A(net808),
    .B(_1006_),
    .C(_2038_));
 sg13g2_nand3_1 _5244_ (.B(_1006_),
    .C(_2038_),
    .A(net808),
    .Y(_2040_));
 sg13g2_and2_1 _5245_ (.A(net1575),
    .B(_2039_),
    .X(_2041_));
 sg13g2_o21ai_1 _5246_ (.B1(net953),
    .Y(_2042_),
    .A1(net1703),
    .A2(_2041_));
 sg13g2_a21oi_1 _5247_ (.A1(net1703),
    .A2(_2039_),
    .Y(_0423_),
    .B1(_2042_));
 sg13g2_xor2_1 _5248_ (.B(net1780),
    .A(net1661),
    .X(_2043_));
 sg13g2_a22oi_1 _5249_ (.Y(_2044_),
    .B1(_2041_),
    .B2(_2043_),
    .A2(_2040_),
    .A1(net1661));
 sg13g2_nor2_1 _5250_ (.A(net908),
    .B(_2044_),
    .Y(_0424_));
 sg13g2_xor2_1 _5251_ (.B(_0997_),
    .A(_0108_),
    .X(_2045_));
 sg13g2_a22oi_1 _5252_ (.Y(_2046_),
    .B1(_2041_),
    .B2(_2045_),
    .A2(_2040_),
    .A1(net1346));
 sg13g2_nor2_1 _5253_ (.A(net908),
    .B(net1347),
    .Y(_0425_));
 sg13g2_a21oi_1 _5254_ (.A1(_0109_),
    .A2(_2037_),
    .Y(_2047_),
    .B1(net914));
 sg13g2_nor2b_2 _5255_ (.A(_0995_),
    .B_N(_2047_),
    .Y(_2048_));
 sg13g2_nor2b_1 _5256_ (.A(_1004_),
    .B_N(_2047_),
    .Y(_2049_));
 sg13g2_o21ai_1 _5257_ (.B1(_1005_),
    .Y(_2050_),
    .A1(_2048_),
    .A2(_2049_));
 sg13g2_a21oi_2 _5258_ (.B1(_2048_),
    .Y(_2051_),
    .A2(_2049_),
    .A1(_1005_));
 sg13g2_inv_2 _5259_ (.Y(_2052_),
    .A(_2051_));
 sg13g2_nand2_1 _5260_ (.Y(_2053_),
    .A(net1546),
    .B(_0995_));
 sg13g2_o21ai_1 _5261_ (.B1(net1530),
    .Y(_2054_),
    .A1(_0992_),
    .A2(_0994_));
 sg13g2_and2_1 _5262_ (.A(_2053_),
    .B(_2054_),
    .X(_2055_));
 sg13g2_o21ai_1 _5263_ (.B1(net954),
    .Y(_2056_),
    .A1(\uart_inst.uart_tx_inst.CLK_CNT[0] ),
    .A2(_2052_));
 sg13g2_a21oi_1 _5264_ (.A1(_2052_),
    .A2(net1531),
    .Y(_0426_),
    .B1(_2056_));
 sg13g2_nor2_1 _5265_ (.A(\uart_inst.uart_tx_inst.CLK_CNT[0] ),
    .B(_2051_),
    .Y(_2057_));
 sg13g2_o21ai_1 _5266_ (.B1(net954),
    .Y(_2058_),
    .A1(net1361),
    .A2(_2057_));
 sg13g2_a21oi_1 _5267_ (.A1(net1361),
    .A2(_2057_),
    .Y(_0427_),
    .B1(_2058_));
 sg13g2_xor2_1 _5268_ (.B(_0990_),
    .A(net1553),
    .X(_2059_));
 sg13g2_a22oi_1 _5269_ (.Y(_2060_),
    .B1(_2059_),
    .B2(_2048_),
    .A2(_2051_),
    .A1(net1553));
 sg13g2_nor2_1 _5270_ (.A(net896),
    .B(net1554),
    .Y(_0428_));
 sg13g2_nor4_1 _5271_ (.A(\uart_inst.uart_tx_inst.CLK_CNT[2] ),
    .B(\uart_inst.uart_tx_inst.CLK_CNT[1] ),
    .C(\uart_inst.uart_tx_inst.CLK_CNT[0] ),
    .D(_2051_),
    .Y(_2061_));
 sg13g2_nand2b_1 _5272_ (.Y(_2062_),
    .B(net1651),
    .A_N(_2061_));
 sg13g2_nor4_1 _5273_ (.A(\uart_inst.uart_tx_inst.CLK_CNT[5] ),
    .B(\uart_inst.uart_tx_inst.CLK_CNT[4] ),
    .C(\uart_inst.uart_tx_inst.state[2] ),
    .D(_0992_),
    .Y(_2063_));
 sg13g2_nand2_2 _5274_ (.Y(_2064_),
    .A(_0991_),
    .B(_2052_));
 sg13g2_o21ai_1 _5275_ (.B1(_2062_),
    .Y(_2065_),
    .A1(_2063_),
    .A2(_2064_));
 sg13g2_and2_1 _5276_ (.A(net954),
    .B(net1652),
    .X(_0429_));
 sg13g2_nor3_1 _5277_ (.A(net1564),
    .B(net1444),
    .C(_0992_),
    .Y(_2066_));
 sg13g2_nor3_1 _5278_ (.A(net1573),
    .B(_2064_),
    .C(_2066_),
    .Y(_2067_));
 sg13g2_a21oi_1 _5279_ (.A1(net1573),
    .A2(_2064_),
    .Y(_2068_),
    .B1(_2067_));
 sg13g2_nor2_1 _5280_ (.A(net896),
    .B(net1574),
    .Y(_0430_));
 sg13g2_o21ai_1 _5281_ (.B1(net1564),
    .Y(_2069_),
    .A1(\uart_inst.uart_tx_inst.CLK_CNT[4] ),
    .A2(_2064_));
 sg13g2_nor3_1 _5282_ (.A(net1564),
    .B(\uart_inst.uart_tx_inst.CLK_CNT[4] ),
    .C(_2064_),
    .Y(_2070_));
 sg13g2_o21ai_1 _5283_ (.B1(_2070_),
    .Y(_2071_),
    .A1(net1444),
    .A2(_0992_));
 sg13g2_a21oi_1 _5284_ (.A1(net1565),
    .A2(_2071_),
    .Y(_0431_),
    .B1(net896));
 sg13g2_o21ai_1 _5285_ (.B1(net1521),
    .Y(_2072_),
    .A1(_0994_),
    .A2(_2051_));
 sg13g2_or3_1 _5286_ (.A(net1521),
    .B(_0994_),
    .C(_2051_),
    .X(_2073_));
 sg13g2_a221oi_1 _5287_ (.B2(_2073_),
    .C1(net897),
    .B1(_2072_),
    .A1(_0995_),
    .Y(_0432_),
    .A2(_2052_));
 sg13g2_nand2_1 _5288_ (.Y(_2074_),
    .A(net1104),
    .B(_2073_));
 sg13g2_or4_1 _5289_ (.A(net1104),
    .B(\uart_inst.uart_tx_inst.CLK_CNT[6] ),
    .C(_0994_),
    .D(_2051_),
    .X(_2075_));
 sg13g2_a21oi_1 _5290_ (.A1(net1105),
    .A2(_2075_),
    .Y(_0433_),
    .B1(net896));
 sg13g2_xor2_1 _5291_ (.B(_2075_),
    .A(\uart_inst.uart_tx_inst.CLK_CNT[8] ),
    .X(_2076_));
 sg13g2_nor3_1 _5292_ (.A(\uart_inst.uart_tx_inst.CLK_CNT[9] ),
    .B(\uart_inst.uart_tx_inst.CLK_CNT[8] ),
    .C(net1444),
    .Y(_2077_));
 sg13g2_nor3_1 _5293_ (.A(net908),
    .B(_2076_),
    .C(net1445),
    .Y(_0434_));
 sg13g2_o21ai_1 _5294_ (.B1(net1673),
    .Y(_2078_),
    .A1(\uart_inst.uart_tx_inst.CLK_CNT[8] ),
    .A2(_2075_));
 sg13g2_o21ai_1 _5295_ (.B1(net1674),
    .Y(_2079_),
    .A1(_2050_),
    .A2(_2053_));
 sg13g2_and2_1 _5296_ (.A(net954),
    .B(_2079_),
    .X(_0435_));
 sg13g2_nor3_1 _5297_ (.A(\uart_inst.uart_tx_inst.state[0] ),
    .B(\uart_inst.uart_tx_inst.state[1] ),
    .C(\uart_inst.uart_tx_inst.state[2] ),
    .Y(_2080_));
 sg13g2_o21ai_1 _5298_ (.B1(_2052_),
    .Y(_2081_),
    .A1(_0995_),
    .A2(_2080_));
 sg13g2_mux4_1 _5299_ (.S0(\uart_inst.uart_tx_inst.DATA_CNT[0] ),
    .A0(\uart_inst.uart_tx_inst.DATA_REG[0] ),
    .A1(\uart_inst.uart_tx_inst.DATA_REG[1] ),
    .A2(\uart_inst.uart_tx_inst.DATA_REG[2] ),
    .A3(\uart_inst.uart_tx_inst.DATA_REG[3] ),
    .S1(\uart_inst.uart_tx_inst.DATA_CNT[1] ),
    .X(_2082_));
 sg13g2_nor2_1 _5300_ (.A(net1346),
    .B(_2082_),
    .Y(_2083_));
 sg13g2_nor2b_1 _5301_ (.A(\uart_inst.uart_tx_inst.DATA_REG[5] ),
    .B_N(\uart_inst.uart_tx_inst.DATA_CNT[0] ),
    .Y(_2084_));
 sg13g2_nor2_1 _5302_ (.A(\uart_inst.uart_tx_inst.DATA_REG[4] ),
    .B(\uart_inst.uart_tx_inst.DATA_CNT[0] ),
    .Y(_2085_));
 sg13g2_nor3_1 _5303_ (.A(\uart_inst.uart_tx_inst.DATA_CNT[1] ),
    .B(_2084_),
    .C(_2085_),
    .Y(_2086_));
 sg13g2_nand2_1 _5304_ (.Y(_2087_),
    .A(\uart_inst.uart_tx_inst.DATA_REG[6] ),
    .B(\uart_inst.uart_tx_inst.DATA_CNT[1] ));
 sg13g2_o21ai_1 _5305_ (.B1(\uart_inst.uart_tx_inst.DATA_CNT[2] ),
    .Y(_2088_),
    .A1(\uart_inst.uart_tx_inst.DATA_CNT[0] ),
    .A2(_2087_));
 sg13g2_o21ai_1 _5306_ (.B1(\uart_inst.uart_tx_inst.state[1] ),
    .Y(_2089_),
    .A1(_2086_),
    .A2(_2088_));
 sg13g2_nor2_1 _5307_ (.A(_2083_),
    .B(_2089_),
    .Y(_2090_));
 sg13g2_nor2_1 _5308_ (.A(\uart_inst.uart_tx_inst.state[2] ),
    .B(_2090_),
    .Y(_2091_));
 sg13g2_a21oi_1 _5309_ (.A1(net1377),
    .A2(_2081_),
    .Y(_2092_),
    .B1(net897));
 sg13g2_o21ai_1 _5310_ (.B1(_2092_),
    .Y(_0436_),
    .A1(_2081_),
    .A2(_2091_));
 sg13g2_nor2_1 _5311_ (.A(_0876_),
    .B(_1008_),
    .Y(_2093_));
 sg13g2_a21oi_1 _5312_ (.A1(\uart_inst.uart_tx_inst.state[0] ),
    .A2(_0996_),
    .Y(_2094_),
    .B1(net1222));
 sg13g2_o21ai_1 _5313_ (.B1(net952),
    .Y(_0437_),
    .A1(net764),
    .A2(net1223));
 sg13g2_and2_2 _5314_ (.A(net964),
    .B(rx_valid),
    .X(_2095_));
 sg13g2_nand2_1 _5315_ (.Y(_2096_),
    .A(net964),
    .B(net1301));
 sg13g2_o21ai_1 _5316_ (.B1(net938),
    .Y(_2097_),
    .A1(\input_value_check_inst.character_buff[9][0] ),
    .A2(net863));
 sg13g2_a21oi_1 _5317_ (.A1(_0873_),
    .A2(net863),
    .Y(_0438_),
    .B1(_2097_));
 sg13g2_o21ai_1 _5318_ (.B1(net938),
    .Y(_2098_),
    .A1(\input_value_check_inst.character_buff[8][1] ),
    .A2(net848));
 sg13g2_a21oi_1 _5319_ (.A1(_0875_),
    .A2(net848),
    .Y(_0439_),
    .B1(_2098_));
 sg13g2_o21ai_1 _5320_ (.B1(net917),
    .Y(_2099_),
    .A1(net1304),
    .A2(net861));
 sg13g2_a21oi_1 _5321_ (.A1(_0872_),
    .A2(net861),
    .Y(_0440_),
    .B1(_2099_));
 sg13g2_o21ai_1 _5322_ (.B1(net918),
    .Y(_2100_),
    .A1(\input_value_check_inst.character_buff[9][3] ),
    .A2(net861));
 sg13g2_a21oi_1 _5323_ (.A1(_0871_),
    .A2(net861),
    .Y(_0441_),
    .B1(_2100_));
 sg13g2_o21ai_1 _5324_ (.B1(net938),
    .Y(_2101_),
    .A1(\input_value_check_inst.character_buff[9][4] ),
    .A2(net864));
 sg13g2_a21oi_1 _5325_ (.A1(_0870_),
    .A2(net863),
    .Y(_0442_),
    .B1(_2101_));
 sg13g2_o21ai_1 _5326_ (.B1(net929),
    .Y(_2102_),
    .A1(\input_value_check_inst.character_buff[9][5] ),
    .A2(net863));
 sg13g2_a21oi_1 _5327_ (.A1(_0869_),
    .A2(net862),
    .Y(_0443_),
    .B1(_2102_));
 sg13g2_o21ai_1 _5328_ (.B1(net917),
    .Y(_2103_),
    .A1(\input_value_check_inst.character_buff[8][6] ),
    .A2(net847));
 sg13g2_a21oi_1 _5329_ (.A1(_0874_),
    .A2(net847),
    .Y(_0444_),
    .B1(_2103_));
 sg13g2_o21ai_1 _5330_ (.B1(net917),
    .Y(_2104_),
    .A1(\input_value_check_inst.character_buff[9][7] ),
    .A2(net861));
 sg13g2_a21oi_1 _5331_ (.A1(_0868_),
    .A2(net861),
    .Y(_0445_),
    .B1(_2104_));
 sg13g2_o21ai_1 _5332_ (.B1(net929),
    .Y(_2105_),
    .A1(\input_value_check_inst.character_buff[8][0] ),
    .A2(net863));
 sg13g2_a21oi_1 _5333_ (.A1(_0867_),
    .A2(net863),
    .Y(_0446_),
    .B1(_2105_));
 sg13g2_o21ai_1 _5334_ (.B1(net929),
    .Y(_2106_),
    .A1(\input_value_check_inst.character_buff[8][1] ),
    .A2(net864));
 sg13g2_a21oi_1 _5335_ (.A1(_0866_),
    .A2(net864),
    .Y(_0447_),
    .B1(_2106_));
 sg13g2_o21ai_1 _5336_ (.B1(net917),
    .Y(_2107_),
    .A1(net1176),
    .A2(net847));
 sg13g2_a21oi_1 _5337_ (.A1(_0872_),
    .A2(net847),
    .Y(_0448_),
    .B1(_2107_));
 sg13g2_o21ai_1 _5338_ (.B1(net917),
    .Y(_2108_),
    .A1(net1153),
    .A2(net861));
 sg13g2_a21oi_1 _5339_ (.A1(_0865_),
    .A2(net861),
    .Y(_0449_),
    .B1(_2108_));
 sg13g2_o21ai_1 _5340_ (.B1(net917),
    .Y(_2109_),
    .A1(net1382),
    .A2(net846));
 sg13g2_a21oi_1 _5341_ (.A1(_0870_),
    .A2(net847),
    .Y(_0450_),
    .B1(_2109_));
 sg13g2_o21ai_1 _5342_ (.B1(net915),
    .Y(_2110_),
    .A1(net1319),
    .A2(net844));
 sg13g2_a21oi_1 _5343_ (.A1(_0869_),
    .A2(net847),
    .Y(_0451_),
    .B1(_2110_));
 sg13g2_o21ai_1 _5344_ (.B1(net915),
    .Y(_2111_),
    .A1(\input_value_check_inst.character_buff[8][6] ),
    .A2(net855));
 sg13g2_a21oi_1 _5345_ (.A1(_0864_),
    .A2(net855),
    .Y(_0452_),
    .B1(_2111_));
 sg13g2_o21ai_1 _5346_ (.B1(net915),
    .Y(_2112_),
    .A1(net1252),
    .A2(net855));
 sg13g2_a21oi_1 _5347_ (.A1(_0863_),
    .A2(net860),
    .Y(_0453_),
    .B1(_2112_));
 sg13g2_o21ai_1 _5348_ (.B1(net929),
    .Y(_2113_),
    .A1(net1260),
    .A2(net847));
 sg13g2_a21oi_1 _5349_ (.A1(_0867_),
    .A2(net847),
    .Y(_0454_),
    .B1(_2113_));
 sg13g2_o21ai_1 _5350_ (.B1(net930),
    .Y(_2114_),
    .A1(net1215),
    .A2(net864));
 sg13g2_a21oi_1 _5351_ (.A1(_0862_),
    .A2(net864),
    .Y(_0455_),
    .B1(_2114_));
 sg13g2_o21ai_1 _5352_ (.B1(net917),
    .Y(_2115_),
    .A1(net1176),
    .A2(net862));
 sg13g2_a21oi_1 _5353_ (.A1(_0861_),
    .A2(net862),
    .Y(_0456_),
    .B1(_2115_));
 sg13g2_o21ai_1 _5354_ (.B1(net916),
    .Y(_2116_),
    .A1(net1295),
    .A2(net855));
 sg13g2_a21oi_1 _5355_ (.A1(_0860_),
    .A2(net855),
    .Y(_0457_),
    .B1(_2116_));
 sg13g2_o21ai_1 _5356_ (.B1(net915),
    .Y(_2117_),
    .A1(\input_value_check_inst.character_buff[7][4] ),
    .A2(net860));
 sg13g2_a21oi_1 _5357_ (.A1(_0859_),
    .A2(net860),
    .Y(_0458_),
    .B1(_2117_));
 sg13g2_o21ai_1 _5358_ (.B1(net915),
    .Y(_2118_),
    .A1(net1319),
    .A2(net854));
 sg13g2_a21oi_1 _5359_ (.A1(_0858_),
    .A2(net854),
    .Y(_0459_),
    .B1(_2118_));
 sg13g2_o21ai_1 _5360_ (.B1(net915),
    .Y(_2119_),
    .A1(\input_value_check_inst.character_buff[7][6] ),
    .A2(net854));
 sg13g2_a21oi_1 _5361_ (.A1(_0857_),
    .A2(net854),
    .Y(_0460_),
    .B1(_2119_));
 sg13g2_o21ai_1 _5362_ (.B1(net915),
    .Y(_2120_),
    .A1(net1271),
    .A2(net844));
 sg13g2_a21oi_1 _5363_ (.A1(_0863_),
    .A2(net844),
    .Y(_0461_),
    .B1(_2120_));
 sg13g2_o21ai_1 _5364_ (.B1(net929),
    .Y(_2121_),
    .A1(net1260),
    .A2(net862));
 sg13g2_a21oi_1 _5365_ (.A1(_0856_),
    .A2(net864),
    .Y(_0462_),
    .B1(_2121_));
 sg13g2_o21ai_1 _5366_ (.B1(net929),
    .Y(_2122_),
    .A1(net1335),
    .A2(net848));
 sg13g2_a21oi_1 _5367_ (.A1(_0862_),
    .A2(net848),
    .Y(_0463_),
    .B1(_2122_));
 sg13g2_o21ai_1 _5368_ (.B1(net926),
    .Y(_2123_),
    .A1(\input_value_check_inst.character_buff[5][2] ),
    .A2(net846));
 sg13g2_a21oi_1 _5369_ (.A1(_0861_),
    .A2(net844),
    .Y(_0464_),
    .B1(_2123_));
 sg13g2_o21ai_1 _5370_ (.B1(net926),
    .Y(_2124_),
    .A1(\input_value_check_inst.character_buff[5][3] ),
    .A2(net844));
 sg13g2_a21oi_1 _5371_ (.A1(_0860_),
    .A2(net844),
    .Y(_0465_),
    .B1(_2124_));
 sg13g2_o21ai_1 _5372_ (.B1(net925),
    .Y(_2125_),
    .A1(net1168),
    .A2(net855));
 sg13g2_a21oi_1 _5373_ (.A1(_0855_),
    .A2(net855),
    .Y(_0466_),
    .B1(_2125_));
 sg13g2_o21ai_1 _5374_ (.B1(net925),
    .Y(_2126_),
    .A1(net1330),
    .A2(net854));
 sg13g2_a21oi_1 _5375_ (.A1(_0854_),
    .A2(net854),
    .Y(_0467_),
    .B1(_2126_));
 sg13g2_o21ai_1 _5376_ (.B1(net925),
    .Y(_2127_),
    .A1(net1375),
    .A2(net844));
 sg13g2_a21oi_1 _5377_ (.A1(_0857_),
    .A2(net844),
    .Y(_0468_),
    .B1(_2127_));
 sg13g2_o21ai_1 _5378_ (.B1(net915),
    .Y(_2128_),
    .A1(net1271),
    .A2(net854));
 sg13g2_a21oi_1 _5379_ (.A1(_0853_),
    .A2(net854),
    .Y(_0469_),
    .B1(_2128_));
 sg13g2_o21ai_1 _5380_ (.B1(net929),
    .Y(_2129_),
    .A1(\input_value_check_inst.character_buff[4][0] ),
    .A2(net848));
 sg13g2_a21oi_1 _5381_ (.A1(_0856_),
    .A2(net848),
    .Y(_0470_),
    .B1(_2129_));
 sg13g2_o21ai_1 _5382_ (.B1(net926),
    .Y(_2130_),
    .A1(\input_value_check_inst.character_buff[5][1] ),
    .A2(net858));
 sg13g2_a21oi_1 _5383_ (.A1(_0852_),
    .A2(net858),
    .Y(_0471_),
    .B1(_2130_));
 sg13g2_o21ai_1 _5384_ (.B1(net926),
    .Y(_2131_),
    .A1(\input_value_check_inst.character_buff[5][2] ),
    .A2(net858));
 sg13g2_a21oi_1 _5385_ (.A1(_0851_),
    .A2(net858),
    .Y(_0472_),
    .B1(_2131_));
 sg13g2_o21ai_1 _5386_ (.B1(net926),
    .Y(_2132_),
    .A1(net1334),
    .A2(net858));
 sg13g2_a21oi_1 _5387_ (.A1(_0850_),
    .A2(net858),
    .Y(_0473_),
    .B1(_2132_));
 sg13g2_o21ai_1 _5388_ (.B1(net925),
    .Y(_2133_),
    .A1(net1233),
    .A2(net856));
 sg13g2_a21oi_1 _5389_ (.A1(_0849_),
    .A2(net856),
    .Y(_0474_),
    .B1(_2133_));
 sg13g2_o21ai_1 _5390_ (.B1(net925),
    .Y(_2134_),
    .A1(\input_value_check_inst.character_buff[5][5] ),
    .A2(net856));
 sg13g2_a21oi_1 _5391_ (.A1(_0848_),
    .A2(net856),
    .Y(_0475_),
    .B1(_2134_));
 sg13g2_o21ai_1 _5392_ (.B1(net925),
    .Y(_2135_),
    .A1(\input_value_check_inst.character_buff[5][6] ),
    .A2(net856));
 sg13g2_a21oi_1 _5393_ (.A1(_0847_),
    .A2(net856),
    .Y(_0476_),
    .B1(_2135_));
 sg13g2_o21ai_1 _5394_ (.B1(net925),
    .Y(_2136_),
    .A1(\input_value_check_inst.character_buff[4][7] ),
    .A2(net845));
 sg13g2_a21oi_1 _5395_ (.A1(_0853_),
    .A2(net845),
    .Y(_0477_),
    .B1(_2136_));
 sg13g2_o21ai_1 _5396_ (.B1(net929),
    .Y(_2137_),
    .A1(net1538),
    .A2(net858));
 sg13g2_a21oi_1 _5397_ (.A1(_0846_),
    .A2(net859),
    .Y(_0478_),
    .B1(_2137_));
 sg13g2_o21ai_1 _5398_ (.B1(net926),
    .Y(_2138_),
    .A1(net1160),
    .A2(net845));
 sg13g2_a21oi_1 _5399_ (.A1(_0852_),
    .A2(net845),
    .Y(_0479_),
    .B1(_2138_));
 sg13g2_o21ai_1 _5400_ (.B1(net925),
    .Y(_2139_),
    .A1(net1261),
    .A2(net845));
 sg13g2_a21oi_1 _5401_ (.A1(_0851_),
    .A2(net845),
    .Y(_0480_),
    .B1(_2139_));
 sg13g2_o21ai_1 _5402_ (.B1(net928),
    .Y(_2140_),
    .A1(\input_value_check_inst.character_buff[3][3] ),
    .A2(net845));
 sg13g2_a21oi_1 _5403_ (.A1(_0850_),
    .A2(net845),
    .Y(_0481_),
    .B1(_2140_));
 sg13g2_o21ai_1 _5404_ (.B1(net927),
    .Y(_2141_),
    .A1(net1241),
    .A2(net857));
 sg13g2_a21oi_1 _5405_ (.A1(_0845_),
    .A2(net857),
    .Y(_0482_),
    .B1(_2141_));
 sg13g2_o21ai_1 _5406_ (.B1(net927),
    .Y(_2142_),
    .A1(net1206),
    .A2(net857));
 sg13g2_a21oi_1 _5407_ (.A1(_0844_),
    .A2(net856),
    .Y(_0483_),
    .B1(_2142_));
 sg13g2_o21ai_1 _5408_ (.B1(net927),
    .Y(_2143_),
    .A1(\input_value_check_inst.character_buff[4][6] ),
    .A2(net865));
 sg13g2_a21oi_1 _5409_ (.A1(_0843_),
    .A2(net865),
    .Y(_0484_),
    .B1(_2143_));
 sg13g2_o21ai_1 _5410_ (.B1(net927),
    .Y(_2144_),
    .A1(\input_value_check_inst.character_buff[4][7] ),
    .A2(net857));
 sg13g2_a21oi_1 _5411_ (.A1(_0842_),
    .A2(net856),
    .Y(_0485_),
    .B1(_2144_));
 sg13g2_o21ai_1 _5412_ (.B1(net930),
    .Y(_2145_),
    .A1(net1655),
    .A2(net858));
 sg13g2_a21oi_1 _5413_ (.A1(_0841_),
    .A2(net869),
    .Y(_0486_),
    .B1(_2145_));
 sg13g2_o21ai_1 _5414_ (.B1(net930),
    .Y(_2146_),
    .A1(net1160),
    .A2(net869));
 sg13g2_a21oi_1 _5415_ (.A1(_0840_),
    .A2(net869),
    .Y(_0487_),
    .B1(_2146_));
 sg13g2_o21ai_1 _5416_ (.B1(net928),
    .Y(_2147_),
    .A1(net1261),
    .A2(net866));
 sg13g2_a21oi_1 _5417_ (.A1(_0839_),
    .A2(net866),
    .Y(_0488_),
    .B1(_2147_));
 sg13g2_o21ai_1 _5418_ (.B1(net928),
    .Y(_2148_),
    .A1(net1588),
    .A2(net859));
 sg13g2_a21oi_1 _5419_ (.A1(_0838_),
    .A2(net866),
    .Y(_0489_),
    .B1(_2148_));
 sg13g2_o21ai_1 _5420_ (.B1(net927),
    .Y(_2149_),
    .A1(net1545),
    .A2(net849));
 sg13g2_a21oi_1 _5421_ (.A1(_0845_),
    .A2(net849),
    .Y(_0490_),
    .B1(_2149_));
 sg13g2_o21ai_1 _5422_ (.B1(net927),
    .Y(_2150_),
    .A1(net1189),
    .A2(net849));
 sg13g2_a21oi_1 _5423_ (.A1(_0844_),
    .A2(net849),
    .Y(_0491_),
    .B1(_2150_));
 sg13g2_o21ai_1 _5424_ (.B1(net927),
    .Y(_2151_),
    .A1(net1336),
    .A2(net849));
 sg13g2_a21oi_1 _5425_ (.A1(_0843_),
    .A2(net849),
    .Y(_0492_),
    .B1(_2151_));
 sg13g2_o21ai_1 _5426_ (.B1(net927),
    .Y(_2152_),
    .A1(net1327),
    .A2(net849));
 sg13g2_a21oi_1 _5427_ (.A1(_0842_),
    .A2(net849),
    .Y(_0493_),
    .B1(_2152_));
 sg13g2_o21ai_1 _5428_ (.B1(net936),
    .Y(_2153_),
    .A1(net1612),
    .A2(net853));
 sg13g2_a21oi_1 _5429_ (.A1(_0841_),
    .A2(net853),
    .Y(_0494_),
    .B1(_2153_));
 sg13g2_o21ai_1 _5430_ (.B1(net936),
    .Y(_2154_),
    .A1(net1597),
    .A2(net851));
 sg13g2_a21oi_1 _5431_ (.A1(_0840_),
    .A2(net852),
    .Y(_0495_),
    .B1(_2154_));
 sg13g2_o21ai_1 _5432_ (.B1(net931),
    .Y(_2155_),
    .A1(net1381),
    .A2(net850));
 sg13g2_a21oi_1 _5433_ (.A1(_0839_),
    .A2(net852),
    .Y(_0496_),
    .B1(_2155_));
 sg13g2_o21ai_1 _5434_ (.B1(net932),
    .Y(_2156_),
    .A1(net1493),
    .A2(net866));
 sg13g2_a21oi_1 _5435_ (.A1(_0837_),
    .A2(net866),
    .Y(_0497_),
    .B1(_2156_));
 sg13g2_o21ai_1 _5436_ (.B1(net932),
    .Y(_2157_),
    .A1(\input_value_check_inst.character_buff[2][4] ),
    .A2(net865));
 sg13g2_a21oi_1 _5437_ (.A1(_0836_),
    .A2(net866),
    .Y(_0498_),
    .B1(_2157_));
 sg13g2_o21ai_1 _5438_ (.B1(net931),
    .Y(_2158_),
    .A1(net1189),
    .A2(net865));
 sg13g2_a21oi_1 _5439_ (.A1(_0835_),
    .A2(net866),
    .Y(_0499_),
    .B1(_2158_));
 sg13g2_o21ai_1 _5440_ (.B1(net931),
    .Y(_2159_),
    .A1(net1336),
    .A2(net865));
 sg13g2_a21oi_1 _5441_ (.A1(_0834_),
    .A2(net865),
    .Y(_0500_),
    .B1(_2159_));
 sg13g2_o21ai_1 _5442_ (.B1(net931),
    .Y(_2160_),
    .A1(net1327),
    .A2(net865));
 sg13g2_a21oi_1 _5443_ (.A1(_0833_),
    .A2(net865),
    .Y(_0501_),
    .B1(_2160_));
 sg13g2_o21ai_1 _5444_ (.B1(net936),
    .Y(_2161_),
    .A1(net1612),
    .A2(net870));
 sg13g2_a21oi_1 _5445_ (.A1(_0831_),
    .A2(net870),
    .Y(_0502_),
    .B1(_2161_));
 sg13g2_o21ai_1 _5446_ (.B1(net936),
    .Y(_2162_),
    .A1(net1597),
    .A2(net867));
 sg13g2_a21oi_1 _5447_ (.A1(_0829_),
    .A2(net867),
    .Y(_0503_),
    .B1(_2162_));
 sg13g2_o21ai_1 _5448_ (.B1(net932),
    .Y(_2163_),
    .A1(net1381),
    .A2(net867));
 sg13g2_a21oi_1 _5449_ (.A1(_0827_),
    .A2(net867),
    .Y(_0504_),
    .B1(_2163_));
 sg13g2_o21ai_1 _5450_ (.B1(net932),
    .Y(_2164_),
    .A1(\input_value_check_inst.character_buff[0][3] ),
    .A2(net851));
 sg13g2_a21oi_1 _5451_ (.A1(_0837_),
    .A2(net851),
    .Y(_0505_),
    .B1(_2164_));
 sg13g2_o21ai_1 _5452_ (.B1(net932),
    .Y(_2165_),
    .A1(net1523),
    .A2(net850));
 sg13g2_a21oi_1 _5453_ (.A1(_0836_),
    .A2(net851),
    .Y(_0506_),
    .B1(_2165_));
 sg13g2_o21ai_1 _5454_ (.B1(net931),
    .Y(_2166_),
    .A1(\input_value_check_inst.character_buff[0][5] ),
    .A2(net850));
 sg13g2_a21oi_1 _5455_ (.A1(_0835_),
    .A2(net850),
    .Y(_0507_),
    .B1(_2166_));
 sg13g2_o21ai_1 _5456_ (.B1(net931),
    .Y(_2167_),
    .A1(net1267),
    .A2(net850));
 sg13g2_a21oi_1 _5457_ (.A1(_0834_),
    .A2(net850),
    .Y(_0508_),
    .B1(_2167_));
 sg13g2_o21ai_1 _5458_ (.B1(net931),
    .Y(_2168_),
    .A1(\input_value_check_inst.character_buff[0][7] ),
    .A2(net850));
 sg13g2_a21oi_1 _5459_ (.A1(_0833_),
    .A2(net850),
    .Y(_0509_),
    .B1(_2168_));
 sg13g2_o21ai_1 _5460_ (.B1(net937),
    .Y(_2169_),
    .A1(net997),
    .A2(net870));
 sg13g2_a21oi_1 _5461_ (.A1(_0832_),
    .A2(net870),
    .Y(_0510_),
    .B1(_2169_));
 sg13g2_o21ai_1 _5462_ (.B1(net934),
    .Y(_2170_),
    .A1(net989),
    .A2(net867));
 sg13g2_a21oi_1 _5463_ (.A1(_0830_),
    .A2(net869),
    .Y(_0511_),
    .B1(_2170_));
 sg13g2_o21ai_1 _5464_ (.B1(net934),
    .Y(_2171_),
    .A1(net1041),
    .A2(net867));
 sg13g2_a21oi_1 _5465_ (.A1(_0828_),
    .A2(net867),
    .Y(_0512_),
    .B1(_2171_));
 sg13g2_o21ai_1 _5466_ (.B1(net935),
    .Y(_2172_),
    .A1(\input_value_check_inst.character_buff[0][3] ),
    .A2(net867));
 sg13g2_a21oi_1 _5467_ (.A1(_0826_),
    .A2(net869),
    .Y(_0513_),
    .B1(_2172_));
 sg13g2_o21ai_1 _5468_ (.B1(net933),
    .Y(_2173_),
    .A1(\input_value_check_inst.character_buff[0][4] ),
    .A2(net868));
 sg13g2_a21oi_1 _5469_ (.A1(_0825_),
    .A2(net868),
    .Y(_0514_),
    .B1(_2173_));
 sg13g2_o21ai_1 _5470_ (.B1(net933),
    .Y(_2174_),
    .A1(\input_value_check_inst.character_buff[0][5] ),
    .A2(net868));
 sg13g2_a21oi_1 _5471_ (.A1(_0824_),
    .A2(net868),
    .Y(_0515_),
    .B1(_2174_));
 sg13g2_o21ai_1 _5472_ (.B1(net931),
    .Y(_2175_),
    .A1(net1267),
    .A2(net868));
 sg13g2_a21oi_1 _5473_ (.A1(_0823_),
    .A2(net868),
    .Y(_0516_),
    .B1(_2175_));
 sg13g2_o21ai_1 _5474_ (.B1(net933),
    .Y(_2176_),
    .A1(\input_value_check_inst.character_buff[0][7] ),
    .A2(net868));
 sg13g2_a21oi_1 _5475_ (.A1(_0822_),
    .A2(net868),
    .Y(_0517_),
    .B1(_2176_));
 sg13g2_and3_1 _5476_ (.X(_0518_),
    .A(_1376_),
    .B(_1379_),
    .C(_1382_));
 sg13g2_nand2_2 _5477_ (.Y(_2177_),
    .A(_1419_),
    .B(_1421_));
 sg13g2_nor3_2 _5478_ (.A(_0876_),
    .B(_1397_),
    .C(_2177_),
    .Y(_2178_));
 sg13g2_nand2_1 _5479_ (.Y(_2179_),
    .A(net880),
    .B(net962));
 sg13g2_nor2_2 _5480_ (.A(_0771_),
    .B(_0985_),
    .Y(_2180_));
 sg13g2_a221oi_1 _5481_ (.B2(_0821_),
    .C1(net908),
    .B1(_2179_),
    .A1(net743),
    .Y(_0520_),
    .A2(_2178_));
 sg13g2_a21oi_1 _5482_ (.A1(_1416_),
    .A2(_2179_),
    .Y(_2181_),
    .B1(net1507));
 sg13g2_a21oi_1 _5483_ (.A1(\uart_tx_fifo_inst.fifo_valid[1] ),
    .A2(net953),
    .Y(_2182_),
    .B1(net825));
 sg13g2_nor2_1 _5484_ (.A(_2181_),
    .B(_2182_),
    .Y(_0521_));
 sg13g2_a21oi_1 _5485_ (.A1(_0821_),
    .A2(net889),
    .Y(_2183_),
    .B1(net880));
 sg13g2_nor3_1 _5486_ (.A(net914),
    .B(\uart_tx_fifo_inst.fifo_valid[1] ),
    .C(_2183_),
    .Y(_2184_));
 sg13g2_a21oi_1 _5487_ (.A1(net1473),
    .A2(net953),
    .Y(_2185_),
    .B1(net825));
 sg13g2_nor2_1 _5488_ (.A(_2184_),
    .B(_2185_),
    .Y(_0522_));
 sg13g2_and2_1 _5489_ (.A(_1405_),
    .B(_1411_),
    .X(_2186_));
 sg13g2_inv_1 _5490_ (.Y(_2187_),
    .A(net759));
 sg13g2_o21ai_1 _5491_ (.B1(_0984_),
    .Y(_2188_),
    .A1(net879),
    .A2(net1496));
 sg13g2_a221oi_1 _5492_ (.B2(net761),
    .C1(_2188_),
    .B1(net889),
    .A1(net879),
    .Y(_2189_),
    .A2(_0820_));
 sg13g2_a21o_1 _5493_ (.A2(net872),
    .A1(net1496),
    .B1(_2189_),
    .X(_0523_));
 sg13g2_and2_2 _5494_ (.A(_1419_),
    .B(_1420_),
    .X(_2190_));
 sg13g2_nand2_1 _5495_ (.Y(_2191_),
    .A(net889),
    .B(_2190_));
 sg13g2_inv_1 _5496_ (.Y(_2192_),
    .A(_2191_));
 sg13g2_o21ai_1 _5497_ (.B1(_0984_),
    .Y(_2193_),
    .A1(net880),
    .A2(net1339));
 sg13g2_a221oi_1 _5498_ (.B2(_2192_),
    .C1(_2193_),
    .B1(net743),
    .A1(net879),
    .Y(_2194_),
    .A2(_0819_));
 sg13g2_a21o_1 _5499_ (.A2(net872),
    .A1(net1339),
    .B1(_2194_),
    .X(_0524_));
 sg13g2_nor2_1 _5500_ (.A(net770),
    .B(_1411_),
    .Y(_2195_));
 sg13g2_inv_2 _5501_ (.Y(_2196_),
    .A(net738));
 sg13g2_o21ai_1 _5502_ (.B1(_0984_),
    .Y(_2197_),
    .A1(net880),
    .A2(net1582));
 sg13g2_a221oi_1 _5503_ (.B2(net738),
    .C1(_2197_),
    .B1(_2192_),
    .A1(net879),
    .Y(_2198_),
    .A2(_0818_));
 sg13g2_a21o_1 _5504_ (.A2(_2027_),
    .A1(net1582),
    .B1(_2198_),
    .X(_0525_));
 sg13g2_nor2_1 _5505_ (.A(_1405_),
    .B(_1412_),
    .Y(_2199_));
 sg13g2_inv_1 _5506_ (.Y(_2200_),
    .A(net756));
 sg13g2_o21ai_1 _5507_ (.B1(_0984_),
    .Y(_2201_),
    .A1(net879),
    .A2(net1595));
 sg13g2_a221oi_1 _5508_ (.B2(net758),
    .C1(_2201_),
    .B1(_2192_),
    .A1(net879),
    .Y(_2202_),
    .A2(_0817_));
 sg13g2_a21o_1 _5509_ (.A2(net872),
    .A1(net1595),
    .B1(_2202_),
    .X(_0526_));
 sg13g2_o21ai_1 _5510_ (.B1(_0984_),
    .Y(_2203_),
    .A1(_0771_),
    .A2(\uart_tx_fifo_inst.fifo_valid[6] ));
 sg13g2_a221oi_1 _5511_ (.B2(_2192_),
    .C1(_2203_),
    .B1(net761),
    .A1(_0771_),
    .Y(_2204_),
    .A2(_0816_));
 sg13g2_a21o_1 _5512_ (.A2(net872),
    .A1(net1578),
    .B1(_2204_),
    .X(_0527_));
 sg13g2_and2_2 _5513_ (.A(net953),
    .B(_2179_),
    .X(_2205_));
 sg13g2_a22oi_1 _5514_ (.Y(_2206_),
    .B1(_2205_),
    .B2(net1420),
    .A2(net825),
    .A1(\uart_tx_fifo_inst.fifo_valid[7] ));
 sg13g2_a21oi_1 _5515_ (.A1(_1415_),
    .A2(_1422_),
    .Y(_0528_),
    .B1(net1421));
 sg13g2_o21ai_1 _5516_ (.B1(_0984_),
    .Y(_2207_),
    .A1(net879),
    .A2(net1427));
 sg13g2_a21oi_1 _5517_ (.A1(net880),
    .A2(_0815_),
    .Y(_2208_),
    .B1(_2207_));
 sg13g2_nand3_1 _5518_ (.B(_1422_),
    .C(net738),
    .A(net889),
    .Y(_2209_));
 sg13g2_a22oi_1 _5519_ (.Y(_2210_),
    .B1(_2208_),
    .B2(_2209_),
    .A2(net872),
    .A1(net1427));
 sg13g2_inv_1 _5520_ (.Y(_0529_),
    .A(_2210_));
 sg13g2_nand2_1 _5521_ (.Y(_2211_),
    .A(net1213),
    .B(net872));
 sg13g2_nand2_1 _5522_ (.Y(_0530_),
    .A(_1418_),
    .B(_2211_));
 sg13g2_nor3_1 _5523_ (.A(_0380_),
    .B(_0381_),
    .C(_0382_),
    .Y(_0531_));
 sg13g2_nor3_1 _5524_ (.A(net1647),
    .B(_1162_),
    .C(_0709_),
    .Y(_0532_));
 sg13g2_nor3_1 _5525_ (.A(_1306_),
    .B(_0692_),
    .C(_0693_),
    .Y(_0534_));
 sg13g2_nand2_1 _5526_ (.Y(_2212_),
    .A(net883),
    .B(net963));
 sg13g2_nor3_1 _5527_ (.A(net887),
    .B(\output_value_inst.send_element_data ),
    .C(_0099_),
    .Y(_2213_));
 sg13g2_a21oi_1 _5528_ (.A1(_1416_),
    .A2(_2212_),
    .Y(_2214_),
    .B1(_2213_));
 sg13g2_a21o_1 _5529_ (.A2(_2212_),
    .A1(_1416_),
    .B1(_2213_),
    .X(_2215_));
 sg13g2_nor2_1 _5530_ (.A(net882),
    .B(net812),
    .Y(_2216_));
 sg13g2_nor2_1 _5531_ (.A(net885),
    .B(_0091_),
    .Y(_2217_));
 sg13g2_o21ai_1 _5532_ (.B1(net881),
    .Y(_2218_),
    .A1(net873),
    .A2(_0067_));
 sg13g2_nor3_1 _5533_ (.A(net810),
    .B(_2217_),
    .C(_2218_),
    .Y(_2219_));
 sg13g2_a221oi_1 _5534_ (.B2(net1629),
    .C1(_2219_),
    .B1(net800),
    .A1(net1616),
    .Y(_2220_),
    .A2(net810));
 sg13g2_nor2_1 _5535_ (.A(net905),
    .B(net1630),
    .Y(_0536_));
 sg13g2_nor2_1 _5536_ (.A(net873),
    .B(_0068_),
    .Y(_2221_));
 sg13g2_o21ai_1 _5537_ (.B1(net881),
    .Y(_2222_),
    .A1(net885),
    .A2(_0092_));
 sg13g2_nor3_1 _5538_ (.A(net810),
    .B(_2221_),
    .C(_2222_),
    .Y(_2223_));
 sg13g2_a221oi_1 _5539_ (.B2(net1670),
    .C1(_2223_),
    .B1(net800),
    .A1(net1625),
    .Y(_2224_),
    .A2(net810));
 sg13g2_nor2_1 _5540_ (.A(net895),
    .B(net1671),
    .Y(_0537_));
 sg13g2_nor2_1 _5541_ (.A(net873),
    .B(_0069_),
    .Y(_2225_));
 sg13g2_o21ai_1 _5542_ (.B1(net881),
    .Y(_2226_),
    .A1(net885),
    .A2(_0093_));
 sg13g2_nor3_1 _5543_ (.A(net809),
    .B(_2225_),
    .C(_2226_),
    .Y(_2227_));
 sg13g2_a221oi_1 _5544_ (.B2(net1602),
    .C1(_2227_),
    .B1(net800),
    .A1(\output_value_inst.character_buff[8][2] ),
    .Y(_2228_),
    .A2(net809));
 sg13g2_nor2_1 _5545_ (.A(net900),
    .B(net1603),
    .Y(_0538_));
 sg13g2_nor2_1 _5546_ (.A(net873),
    .B(_0070_),
    .Y(_2229_));
 sg13g2_o21ai_1 _5547_ (.B1(net881),
    .Y(_2230_),
    .A1(net885),
    .A2(_0094_));
 sg13g2_nor3_1 _5548_ (.A(net809),
    .B(_2229_),
    .C(_2230_),
    .Y(_2231_));
 sg13g2_a221oi_1 _5549_ (.B2(\output_value_inst.character_buff[9][3] ),
    .C1(_2231_),
    .B1(net800),
    .A1(net1653),
    .Y(_2232_),
    .A2(net809));
 sg13g2_nor2_1 _5550_ (.A(net900),
    .B(net1654),
    .Y(_0539_));
 sg13g2_nor2_1 _5551_ (.A(net873),
    .B(_0071_),
    .Y(_2233_));
 sg13g2_o21ai_1 _5552_ (.B1(net881),
    .Y(_2234_),
    .A1(net885),
    .A2(_0095_));
 sg13g2_nor3_1 _5553_ (.A(net809),
    .B(_2233_),
    .C(_2234_),
    .Y(_2235_));
 sg13g2_a221oi_1 _5554_ (.B2(net1643),
    .C1(_2235_),
    .B1(net800),
    .A1(net1608),
    .Y(_2236_),
    .A2(net811));
 sg13g2_nor2_1 _5555_ (.A(net905),
    .B(net1644),
    .Y(_0540_));
 sg13g2_nor2_1 _5556_ (.A(net873),
    .B(_0072_),
    .Y(_2237_));
 sg13g2_o21ai_1 _5557_ (.B1(net881),
    .Y(_2238_),
    .A1(net885),
    .A2(_0096_));
 sg13g2_nor3_1 _5558_ (.A(net809),
    .B(_2237_),
    .C(_2238_),
    .Y(_2239_));
 sg13g2_a221oi_1 _5559_ (.B2(net1610),
    .C1(_2239_),
    .B1(net800),
    .A1(net1586),
    .Y(_2240_),
    .A2(net811));
 sg13g2_nor2_1 _5560_ (.A(net905),
    .B(net1611),
    .Y(_0541_));
 sg13g2_nand3_1 _5561_ (.B(net1562),
    .C(net1494),
    .A(net1552),
    .Y(_2241_));
 sg13g2_nand3_1 _5562_ (.B(_0878_),
    .C(_0152_),
    .A(_0877_),
    .Y(_2242_));
 sg13g2_o21ai_1 _5563_ (.B1(_2242_),
    .Y(_2243_),
    .A1(\uart_inst.uart_rx_inst.SIGNAL_Q[1] ),
    .A2(\uart_inst.uart_rx_inst.SIGNAL_Q[0] ));
 sg13g2_o21ai_1 _5564_ (.B1(net1552),
    .Y(_2244_),
    .A1(\uart_inst.uart_rx_inst.SIGNAL_Q[3] ),
    .A2(\uart_inst.uart_rx_inst.SIGNAL_Q[2] ));
 sg13g2_a22oi_1 _5565_ (.Y(_2245_),
    .B1(net1383),
    .B2(net1385),
    .A2(\uart_inst.uart_rx_inst.SIGNAL_Q[2] ),
    .A1(net1624));
 sg13g2_a221oi_1 _5566_ (.B2(_2245_),
    .C1(net913),
    .B1(_2244_),
    .A1(_2241_),
    .Y(_2246_),
    .A2(_2243_));
 sg13g2_a21oi_1 _5567_ (.A1(net913),
    .A2(net1356),
    .Y(_2247_),
    .B1(net893));
 sg13g2_nand2b_1 _5568_ (.Y(_0542_),
    .B(_2247_),
    .A_N(_2246_));
 sg13g2_nor3_1 _5569_ (.A(_1292_),
    .B(_1295_),
    .C(_1298_),
    .Y(_0543_));
 sg13g2_a22oi_1 _5570_ (.Y(_2248_),
    .B1(net775),
    .B2(net1200),
    .A2(net748),
    .A1(net1190));
 sg13g2_nand2_2 _5571_ (.Y(_2249_),
    .A(net959),
    .B(_2178_));
 sg13g2_nor2_2 _5572_ (.A(_2196_),
    .B(_2249_),
    .Y(_2250_));
 sg13g2_nor2_1 _5573_ (.A(_2248_),
    .B(_2250_),
    .Y(_0545_));
 sg13g2_a22oi_1 _5574_ (.Y(_2251_),
    .B1(net775),
    .B2(net992),
    .A2(net748),
    .A1(net1097));
 sg13g2_nor2_1 _5575_ (.A(_2250_),
    .B(_2251_),
    .Y(_0546_));
 sg13g2_a22oi_1 _5576_ (.Y(_2252_),
    .B1(net772),
    .B2(net1087),
    .A2(net745),
    .A1(net1062));
 sg13g2_nor2_1 _5577_ (.A(_2250_),
    .B(_2252_),
    .Y(_0547_));
 sg13g2_a22oi_1 _5578_ (.Y(_2253_),
    .B1(net771),
    .B2(net1118),
    .A2(net744),
    .A1(net702));
 sg13g2_nor2_1 _5579_ (.A(_2250_),
    .B(_2253_),
    .Y(_0548_));
 sg13g2_a22oi_1 _5580_ (.Y(_2254_),
    .B1(net771),
    .B2(net1059),
    .A2(net744),
    .A1(net697));
 sg13g2_nor2_1 _5581_ (.A(_2250_),
    .B(_2254_),
    .Y(_0549_));
 sg13g2_a22oi_1 _5582_ (.Y(_2255_),
    .B1(net777),
    .B2(net1132),
    .A2(net750),
    .A1(net1178));
 sg13g2_nor2_1 _5583_ (.A(_2250_),
    .B(_2255_),
    .Y(_0550_));
 sg13g2_a22oi_1 _5584_ (.Y(_2256_),
    .B1(net777),
    .B2(net1133),
    .A2(net750),
    .A1(net974));
 sg13g2_nor2_1 _5585_ (.A(_2250_),
    .B(_2256_),
    .Y(_0551_));
 sg13g2_a22oi_1 _5586_ (.Y(_2257_),
    .B1(net775),
    .B2(net1190),
    .A2(net748),
    .A1(\uart_tx_fifo_inst.fifo[2][0] ));
 sg13g2_nor2_2 _5587_ (.A(_2200_),
    .B(_2249_),
    .Y(_2258_));
 sg13g2_nor2_1 _5588_ (.A(net1191),
    .B(_2258_),
    .Y(_0552_));
 sg13g2_a22oi_1 _5589_ (.Y(_2259_),
    .B1(net775),
    .B2(net1097),
    .A2(net748),
    .A1(net1050));
 sg13g2_nor2_1 _5590_ (.A(_2258_),
    .B(_2259_),
    .Y(_0553_));
 sg13g2_a22oi_1 _5591_ (.Y(_2260_),
    .B1(net772),
    .B2(net1062),
    .A2(net745),
    .A1(\uart_tx_fifo_inst.fifo[2][2] ));
 sg13g2_nor2_1 _5592_ (.A(_2258_),
    .B(net1063),
    .Y(_0554_));
 sg13g2_a22oi_1 _5593_ (.Y(_2261_),
    .B1(net771),
    .B2(net702),
    .A2(net744),
    .A1(\uart_tx_fifo_inst.fifo[2][3] ));
 sg13g2_nor2_1 _5594_ (.A(_2258_),
    .B(net703),
    .Y(_0555_));
 sg13g2_a22oi_1 _5595_ (.Y(_2262_),
    .B1(net771),
    .B2(net697),
    .A2(net744),
    .A1(\uart_tx_fifo_inst.fifo[2][4] ));
 sg13g2_nor2_1 _5596_ (.A(_2258_),
    .B(net698),
    .Y(_0556_));
 sg13g2_a22oi_1 _5597_ (.Y(_2263_),
    .B1(net777),
    .B2(net1178),
    .A2(net750),
    .A1(net690));
 sg13g2_nor2_1 _5598_ (.A(_2258_),
    .B(_2263_),
    .Y(_0557_));
 sg13g2_a22oi_1 _5599_ (.Y(_2264_),
    .B1(net775),
    .B2(net974),
    .A2(net748),
    .A1(\uart_tx_fifo_inst.fifo[2][6] ));
 sg13g2_nor2_1 _5600_ (.A(_2258_),
    .B(net975),
    .Y(_0558_));
 sg13g2_a22oi_1 _5601_ (.Y(_2265_),
    .B1(net775),
    .B2(net1418),
    .A2(net748),
    .A1(net607));
 sg13g2_nor2_2 _5602_ (.A(_2187_),
    .B(_2249_),
    .Y(_2266_));
 sg13g2_nor2_1 _5603_ (.A(_2265_),
    .B(_2266_),
    .Y(_0559_));
 sg13g2_a22oi_1 _5604_ (.Y(_2267_),
    .B1(net775),
    .B2(net1050),
    .A2(net748),
    .A1(\uart_tx_fifo_inst.fifo[3][1] ));
 sg13g2_nor2_1 _5605_ (.A(_2266_),
    .B(net1051),
    .Y(_0560_));
 sg13g2_a22oi_1 _5606_ (.Y(_2268_),
    .B1(net772),
    .B2(net1159),
    .A2(net745),
    .A1(net1057));
 sg13g2_nor2_1 _5607_ (.A(_2266_),
    .B(_2268_),
    .Y(_0561_));
 sg13g2_a22oi_1 _5608_ (.Y(_2269_),
    .B1(net771),
    .B2(net1016),
    .A2(net744),
    .A1(\uart_tx_fifo_inst.fifo[3][3] ));
 sg13g2_nor2_1 _5609_ (.A(_2266_),
    .B(net1017),
    .Y(_0562_));
 sg13g2_a22oi_1 _5610_ (.Y(_2270_),
    .B1(net771),
    .B2(net1058),
    .A2(net744),
    .A1(net993));
 sg13g2_nor2_1 _5611_ (.A(_2266_),
    .B(_2270_),
    .Y(_0563_));
 sg13g2_a22oi_1 _5612_ (.Y(_2271_),
    .B1(net777),
    .B2(net690),
    .A2(net750),
    .A1(\uart_tx_fifo_inst.fifo[3][5] ));
 sg13g2_nor2_1 _5613_ (.A(_2266_),
    .B(net691),
    .Y(_0564_));
 sg13g2_a22oi_1 _5614_ (.Y(_2272_),
    .B1(net776),
    .B2(net1010),
    .A2(net749),
    .A1(\uart_tx_fifo_inst.fifo[3][6] ));
 sg13g2_nor2_1 _5615_ (.A(_2266_),
    .B(net1011),
    .Y(_0565_));
 sg13g2_a22oi_1 _5616_ (.Y(_2273_),
    .B1(net776),
    .B2(net607),
    .A2(net749),
    .A1(\uart_tx_fifo_inst.fifo[4][0] ));
 sg13g2_nor2b_2 _5617_ (.A(net740),
    .B_N(_2190_),
    .Y(_2274_));
 sg13g2_nand3_1 _5618_ (.B(_1417_),
    .C(_2190_),
    .A(net959),
    .Y(_2275_));
 sg13g2_nor2_2 _5619_ (.A(_1414_),
    .B(_2275_),
    .Y(_2276_));
 sg13g2_nor2_1 _5620_ (.A(net608),
    .B(_2276_),
    .Y(_0566_));
 sg13g2_a22oi_1 _5621_ (.Y(_2277_),
    .B1(net776),
    .B2(net1286),
    .A2(net749),
    .A1(net1008));
 sg13g2_nor2_1 _5622_ (.A(_2276_),
    .B(_2277_),
    .Y(_0567_));
 sg13g2_a22oi_1 _5623_ (.Y(_2278_),
    .B1(net772),
    .B2(net1057),
    .A2(net745),
    .A1(net998));
 sg13g2_nor2_1 _5624_ (.A(_2276_),
    .B(_2278_),
    .Y(_0568_));
 sg13g2_a22oi_1 _5625_ (.Y(_2279_),
    .B1(net771),
    .B2(net1093),
    .A2(net744),
    .A1(\uart_tx_fifo_inst.fifo[4][3] ));
 sg13g2_nor2_1 _5626_ (.A(_2276_),
    .B(net1094),
    .Y(_0569_));
 sg13g2_a22oi_1 _5627_ (.Y(_2280_),
    .B1(net772),
    .B2(net993),
    .A2(net745),
    .A1(\uart_tx_fifo_inst.fifo[4][4] ));
 sg13g2_nor2_1 _5628_ (.A(_2276_),
    .B(net994),
    .Y(_0570_));
 sg13g2_a22oi_1 _5629_ (.Y(_2281_),
    .B1(net777),
    .B2(net1055),
    .A2(net750),
    .A1(\uart_tx_fifo_inst.fifo[4][5] ));
 sg13g2_nor2_1 _5630_ (.A(_2276_),
    .B(net1056),
    .Y(_0571_));
 sg13g2_a22oi_1 _5631_ (.Y(_2282_),
    .B1(net776),
    .B2(net1195),
    .A2(net749),
    .A1(net1177));
 sg13g2_nor2_1 _5632_ (.A(_2276_),
    .B(_2282_),
    .Y(_0572_));
 sg13g2_a22oi_1 _5633_ (.Y(_2283_),
    .B1(net778),
    .B2(net1090),
    .A2(net751),
    .A1(\uart_tx_fifo_inst.fifo[5][0] ));
 sg13g2_nor2_2 _5634_ (.A(_2196_),
    .B(_2275_),
    .Y(_2284_));
 sg13g2_nor2_1 _5635_ (.A(net1091),
    .B(_2284_),
    .Y(_0573_));
 sg13g2_a22oi_1 _5636_ (.Y(_2285_),
    .B1(net778),
    .B2(net1008),
    .A2(net751),
    .A1(\uart_tx_fifo_inst.fifo[5][1] ));
 sg13g2_nor2_1 _5637_ (.A(_2284_),
    .B(net1009),
    .Y(_0574_));
 sg13g2_a22oi_1 _5638_ (.Y(_2286_),
    .B1(net773),
    .B2(net998),
    .A2(net746),
    .A1(\uart_tx_fifo_inst.fifo[5][2] ));
 sg13g2_nor2_1 _5639_ (.A(_2284_),
    .B(net999),
    .Y(_0575_));
 sg13g2_a22oi_1 _5640_ (.Y(_2287_),
    .B1(net771),
    .B2(net1126),
    .A2(net744),
    .A1(net1116));
 sg13g2_nor2_1 _5641_ (.A(_2284_),
    .B(_2287_),
    .Y(_0576_));
 sg13g2_a22oi_1 _5642_ (.Y(_2288_),
    .B1(net777),
    .B2(net1147),
    .A2(net750),
    .A1(\uart_tx_fifo_inst.fifo[5][4] ));
 sg13g2_nor2_1 _5643_ (.A(_2284_),
    .B(net1148),
    .Y(_0577_));
 sg13g2_a22oi_1 _5644_ (.Y(_2289_),
    .B1(net777),
    .B2(net1157),
    .A2(net750),
    .A1(\uart_tx_fifo_inst.fifo[5][5] ));
 sg13g2_nor2_1 _5645_ (.A(_2284_),
    .B(net1158),
    .Y(_0578_));
 sg13g2_a22oi_1 _5646_ (.Y(_2290_),
    .B1(net775),
    .B2(net1177),
    .A2(net748),
    .A1(net1102));
 sg13g2_nor2_1 _5647_ (.A(_2284_),
    .B(_2290_),
    .Y(_0579_));
 sg13g2_a22oi_1 _5648_ (.Y(_2291_),
    .B1(net779),
    .B2(net1265),
    .A2(net752),
    .A1(net718));
 sg13g2_nor2_2 _5649_ (.A(_2200_),
    .B(_2275_),
    .Y(_2292_));
 sg13g2_nor2_1 _5650_ (.A(_2291_),
    .B(_2292_),
    .Y(_0580_));
 sg13g2_a22oi_1 _5651_ (.Y(_2293_),
    .B1(net779),
    .B2(net1281),
    .A2(net752),
    .A1(net1006));
 sg13g2_nor2_1 _5652_ (.A(_2292_),
    .B(_2293_),
    .Y(_0581_));
 sg13g2_a22oi_1 _5653_ (.Y(_2294_),
    .B1(net773),
    .B2(net1052),
    .A2(net746),
    .A1(net1039));
 sg13g2_nor2_1 _5654_ (.A(_2292_),
    .B(_2294_),
    .Y(_0582_));
 sg13g2_a22oi_1 _5655_ (.Y(_2295_),
    .B1(net773),
    .B2(net1116),
    .A2(net746),
    .A1(\uart_tx_fifo_inst.fifo[6][3] ));
 sg13g2_nor2_1 _5656_ (.A(_2292_),
    .B(net1117),
    .Y(_0583_));
 sg13g2_a22oi_1 _5657_ (.Y(_2296_),
    .B1(net780),
    .B2(net1318),
    .A2(net753),
    .A1(net968));
 sg13g2_nor2_1 _5658_ (.A(_2292_),
    .B(_2296_),
    .Y(_0584_));
 sg13g2_a22oi_1 _5659_ (.Y(_2297_),
    .B1(net778),
    .B2(net1170),
    .A2(net751),
    .A1(net966));
 sg13g2_nor2_1 _5660_ (.A(_2292_),
    .B(_2297_),
    .Y(_0585_));
 sg13g2_a22oi_1 _5661_ (.Y(_2298_),
    .B1(net778),
    .B2(net1102),
    .A2(net751),
    .A1(net724));
 sg13g2_nor2_1 _5662_ (.A(_2292_),
    .B(_2298_),
    .Y(_0586_));
 sg13g2_a22oi_1 _5663_ (.Y(_2299_),
    .B1(net778),
    .B2(net718),
    .A2(net751),
    .A1(\uart_tx_fifo_inst.fifo[7][0] ));
 sg13g2_nor2_2 _5664_ (.A(_2187_),
    .B(_2275_),
    .Y(_2300_));
 sg13g2_nor2_1 _5665_ (.A(net719),
    .B(_2300_),
    .Y(_0587_));
 sg13g2_a22oi_1 _5666_ (.Y(_2301_),
    .B1(net778),
    .B2(net1006),
    .A2(net751),
    .A1(\uart_tx_fifo_inst.fifo[7][1] ));
 sg13g2_nor2_1 _5667_ (.A(_2300_),
    .B(net1007),
    .Y(_0588_));
 sg13g2_a22oi_1 _5668_ (.Y(_2302_),
    .B1(net773),
    .B2(net1039),
    .A2(net746),
    .A1(\uart_tx_fifo_inst.fifo[7][2] ));
 sg13g2_nor2_1 _5669_ (.A(_2300_),
    .B(net1040),
    .Y(_0589_));
 sg13g2_a22oi_1 _5670_ (.Y(_2303_),
    .B1(net773),
    .B2(net1257),
    .A2(net746),
    .A1(net695));
 sg13g2_nor2_1 _5671_ (.A(_2300_),
    .B(_2303_),
    .Y(_0590_));
 sg13g2_a22oi_1 _5672_ (.Y(_2304_),
    .B1(net780),
    .B2(net968),
    .A2(net753),
    .A1(\uart_tx_fifo_inst.fifo[7][4] ));
 sg13g2_nor2_1 _5673_ (.A(_2300_),
    .B(net969),
    .Y(_0591_));
 sg13g2_a22oi_1 _5674_ (.Y(_2305_),
    .B1(net780),
    .B2(net966),
    .A2(net753),
    .A1(\uart_tx_fifo_inst.fifo[7][5] ));
 sg13g2_nor2_1 _5675_ (.A(_2300_),
    .B(net967),
    .Y(_0592_));
 sg13g2_a22oi_1 _5676_ (.Y(_2306_),
    .B1(net778),
    .B2(net724),
    .A2(net751),
    .A1(\uart_tx_fifo_inst.fifo[7][6] ));
 sg13g2_nor2_1 _5677_ (.A(_2300_),
    .B(net965),
    .Y(_0593_));
 sg13g2_nor2_2 _5678_ (.A(net878),
    .B(net875),
    .Y(_2307_));
 sg13g2_a21oi_1 _5679_ (.A1(net1312),
    .A2(_2307_),
    .Y(_2308_),
    .B1(net811));
 sg13g2_o21ai_1 _5680_ (.B1(net945),
    .Y(_2309_),
    .A1(\output_value_inst.character_buff[9][0] ),
    .A2(net824));
 sg13g2_nor2_1 _5681_ (.A(_2308_),
    .B(_2309_),
    .Y(_0594_));
 sg13g2_a21oi_1 _5682_ (.A1(net1451),
    .A2(_2307_),
    .Y(_2310_),
    .B1(net812));
 sg13g2_o21ai_1 _5683_ (.B1(net960),
    .Y(_2311_),
    .A1(\output_value_inst.character_buff[9][1] ),
    .A2(net824));
 sg13g2_nor2_1 _5684_ (.A(_2310_),
    .B(_2311_),
    .Y(_0595_));
 sg13g2_a21oi_1 _5685_ (.A1(net1193),
    .A2(_2307_),
    .Y(_2312_),
    .B1(net811));
 sg13g2_o21ai_1 _5686_ (.B1(net946),
    .Y(_2313_),
    .A1(\output_value_inst.character_buff[9][2] ),
    .A2(net824));
 sg13g2_nor2_1 _5687_ (.A(_2312_),
    .B(_2313_),
    .Y(_0596_));
 sg13g2_a21oi_1 _5688_ (.A1(net1263),
    .A2(_2307_),
    .Y(_2314_),
    .B1(net811));
 sg13g2_o21ai_1 _5689_ (.B1(net946),
    .Y(_2315_),
    .A1(\output_value_inst.character_buff[9][3] ),
    .A2(net824));
 sg13g2_nor2_1 _5690_ (.A(_2314_),
    .B(_2315_),
    .Y(_0597_));
 sg13g2_o21ai_1 _5691_ (.B1(net883),
    .Y(_2316_),
    .A1(net875),
    .A2(net1455));
 sg13g2_o21ai_1 _5692_ (.B1(net951),
    .Y(_2317_),
    .A1(\output_value_inst.character_buff[9][4] ),
    .A2(net824));
 sg13g2_a21oi_1 _5693_ (.A1(net824),
    .A2(_2316_),
    .Y(_0598_),
    .B1(_2317_));
 sg13g2_a21oi_1 _5694_ (.A1(net1291),
    .A2(_2307_),
    .Y(_2318_),
    .B1(net811));
 sg13g2_o21ai_1 _5695_ (.B1(net945),
    .Y(_2319_),
    .A1(\output_value_inst.character_buff[9][6] ),
    .A2(net824));
 sg13g2_nor2_1 _5696_ (.A(_2318_),
    .B(_2319_),
    .Y(_0599_));
 sg13g2_nand2_1 _5697_ (.Y(_2320_),
    .A(net1437),
    .B(net783));
 sg13g2_a21oi_1 _5698_ (.A1(_1342_),
    .A2(_2320_),
    .Y(_0600_),
    .B1(net893));
 sg13g2_nand2_1 _5699_ (.Y(_2321_),
    .A(net1475),
    .B(net783));
 sg13g2_a21oi_1 _5700_ (.A1(_1336_),
    .A2(_2321_),
    .Y(_0601_),
    .B1(net893));
 sg13g2_nand2_1 _5701_ (.Y(_2322_),
    .A(uo_out[7]),
    .B(net783));
 sg13g2_a21oi_1 _5702_ (.A1(_1043_),
    .A2(_2322_),
    .Y(_0607_),
    .B1(net893));
 sg13g2_a21oi_1 _5703_ (.A1(net711),
    .A2(net782),
    .Y(_2323_),
    .B1(_1142_));
 sg13g2_nor2_1 _5704_ (.A(net894),
    .B(net712),
    .Y(_0608_));
 sg13g2_a21oi_1 _5705_ (.A1(net720),
    .A2(net782),
    .Y(_2324_),
    .B1(_1126_));
 sg13g2_nor2_1 _5706_ (.A(net894),
    .B(net721),
    .Y(_0609_));
 sg13g2_nand2_1 _5707_ (.Y(_2325_),
    .A(net976),
    .B(net782));
 sg13g2_a21oi_1 _5708_ (.A1(_1197_),
    .A2(_2325_),
    .Y(_0612_),
    .B1(net894));
 sg13g2_nand2_1 _5709_ (.Y(_2326_),
    .A(net982),
    .B(net782));
 sg13g2_a21oi_1 _5710_ (.A1(_1191_),
    .A2(_2326_),
    .Y(_0613_),
    .B1(net894));
 sg13g2_nor3_1 _5711_ (.A(\input_value_check_inst.character_buff[9][4] ),
    .B(_0875_),
    .C(\input_value_check_inst.character_buff[9][0] ),
    .Y(_2327_));
 sg13g2_nor2_1 _5712_ (.A(\input_value_check_inst.character_buff[8][1] ),
    .B(\input_value_check_inst.character_buff[8][0] ),
    .Y(_2328_));
 sg13g2_nand3_1 _5713_ (.B(_2327_),
    .C(_2328_),
    .A(_1013_),
    .Y(_2329_));
 sg13g2_nor4_2 _5714_ (.A(_1024_),
    .B(_1026_),
    .C(_1027_),
    .Y(_2330_),
    .D(_2329_));
 sg13g2_nor2_1 _5715_ (.A(net1443),
    .B(net784),
    .Y(_2331_));
 sg13g2_nor2b_1 _5716_ (.A(_1341_),
    .B_N(_2330_),
    .Y(_2332_));
 sg13g2_nor3_1 _5717_ (.A(net892),
    .B(_2331_),
    .C(_2332_),
    .Y(_0616_));
 sg13g2_nor2_1 _5718_ (.A(net1467),
    .B(net784),
    .Y(_2333_));
 sg13g2_nor2b_1 _5719_ (.A(_1335_),
    .B_N(_2330_),
    .Y(_2334_));
 sg13g2_nor3_1 _5720_ (.A(net891),
    .B(_2333_),
    .C(_2334_),
    .Y(_0617_));
 sg13g2_nand2_1 _5721_ (.Y(_2335_),
    .A(_1331_),
    .B(net784));
 sg13g2_o21ai_1 _5722_ (.B1(_2335_),
    .Y(_2336_),
    .A1(net1672),
    .A2(net784));
 sg13g2_nor2_1 _5723_ (.A(net891),
    .B(_2336_),
    .Y(_0618_));
 sg13g2_nor2_1 _5724_ (.A(net1662),
    .B(net784),
    .Y(_2337_));
 sg13g2_and2_1 _5725_ (.A(_1330_),
    .B(net784),
    .X(_2338_));
 sg13g2_nor3_1 _5726_ (.A(net891),
    .B(_2337_),
    .C(_2338_),
    .Y(_0619_));
 sg13g2_nor2_1 _5727_ (.A(net1302),
    .B(net784),
    .Y(_2339_));
 sg13g2_and2_1 _5728_ (.A(_1056_),
    .B(net784),
    .X(_2340_));
 sg13g2_nor3_1 _5729_ (.A(net891),
    .B(_2339_),
    .C(_2340_),
    .Y(_0620_));
 sg13g2_nor2_1 _5730_ (.A(net874),
    .B(_0061_),
    .Y(_2341_));
 sg13g2_o21ai_1 _5731_ (.B1(net882),
    .Y(_2342_),
    .A1(net886),
    .A2(_0085_));
 sg13g2_nor3_1 _5732_ (.A(net810),
    .B(_2341_),
    .C(_2342_),
    .Y(_2343_));
 sg13g2_a221oi_1 _5733_ (.B2(net1616),
    .C1(_2343_),
    .B1(net801),
    .A1(net1548),
    .Y(_2344_),
    .A2(net813));
 sg13g2_nor2_1 _5734_ (.A(net905),
    .B(net1617),
    .Y(_0621_));
 sg13g2_nor2_1 _5735_ (.A(net873),
    .B(_0062_),
    .Y(_2345_));
 sg13g2_o21ai_1 _5736_ (.B1(net882),
    .Y(_2346_),
    .A1(net886),
    .A2(_0086_));
 sg13g2_nor3_1 _5737_ (.A(net810),
    .B(_2345_),
    .C(_2346_),
    .Y(_2347_));
 sg13g2_a221oi_1 _5738_ (.B2(net1625),
    .C1(_2347_),
    .B1(net801),
    .A1(\output_value_inst.character_buff[7][1] ),
    .Y(_2348_),
    .A2(net812));
 sg13g2_nor2_1 _5739_ (.A(net905),
    .B(net1626),
    .Y(_0622_));
 sg13g2_nor2_1 _5740_ (.A(net874),
    .B(_0063_),
    .Y(_2349_));
 sg13g2_o21ai_1 _5741_ (.B1(net881),
    .Y(_2350_),
    .A1(net886),
    .A2(_0087_));
 sg13g2_nor3_1 _5742_ (.A(net809),
    .B(_2349_),
    .C(_2350_),
    .Y(_2351_));
 sg13g2_a221oi_1 _5743_ (.B2(net1638),
    .C1(_2351_),
    .B1(net800),
    .A1(net1604),
    .Y(_2352_),
    .A2(net811));
 sg13g2_nor2_1 _5744_ (.A(net905),
    .B(net1639),
    .Y(_0623_));
 sg13g2_nor2_1 _5745_ (.A(net873),
    .B(net1664),
    .Y(_2353_));
 sg13g2_o21ai_1 _5746_ (.B1(net881),
    .Y(_2354_),
    .A1(net885),
    .A2(_0088_));
 sg13g2_nor3_1 _5747_ (.A(net809),
    .B(_2353_),
    .C(_2354_),
    .Y(_2355_));
 sg13g2_a221oi_1 _5748_ (.B2(net1653),
    .C1(_2355_),
    .B1(net800),
    .A1(net1622),
    .Y(_2356_),
    .A2(net811));
 sg13g2_nor2_1 _5749_ (.A(net905),
    .B(_2356_),
    .Y(_0624_));
 sg13g2_nor2_1 _5750_ (.A(net874),
    .B(_0065_),
    .Y(_2357_));
 sg13g2_o21ai_1 _5751_ (.B1(net882),
    .Y(_2358_),
    .A1(net886),
    .A2(_0089_));
 sg13g2_nor3_1 _5752_ (.A(net810),
    .B(_2357_),
    .C(_2358_),
    .Y(_2359_));
 sg13g2_a221oi_1 _5753_ (.B2(net1608),
    .C1(_2359_),
    .B1(net801),
    .A1(\output_value_inst.character_buff[7][4] ),
    .Y(_2360_),
    .A2(net812));
 sg13g2_nor2_1 _5754_ (.A(net906),
    .B(net1609),
    .Y(_0625_));
 sg13g2_nor2_1 _5755_ (.A(net874),
    .B(_0066_),
    .Y(_2361_));
 sg13g2_o21ai_1 _5756_ (.B1(net882),
    .Y(_2362_),
    .A1(net886),
    .A2(_0090_));
 sg13g2_nor3_1 _5757_ (.A(net810),
    .B(_2361_),
    .C(_2362_),
    .Y(_2363_));
 sg13g2_a221oi_1 _5758_ (.B2(net1586),
    .C1(_2363_),
    .B1(net801),
    .A1(\output_value_inst.character_buff[7][6] ),
    .Y(_2364_),
    .A2(net812));
 sg13g2_nor2_1 _5759_ (.A(net905),
    .B(net1587),
    .Y(_0626_));
 sg13g2_nor2_1 _5760_ (.A(net876),
    .B(_0055_),
    .Y(_2365_));
 sg13g2_o21ai_1 _5761_ (.B1(net883),
    .Y(_2366_),
    .A1(net888),
    .A2(_0079_));
 sg13g2_nor3_1 _5762_ (.A(net814),
    .B(_2365_),
    .C(_2366_),
    .Y(_2367_));
 sg13g2_a221oi_1 _5763_ (.B2(net1548),
    .C1(_2367_),
    .B1(net802),
    .A1(net1192),
    .Y(_2368_),
    .A2(net814));
 sg13g2_nor2_1 _5764_ (.A(net907),
    .B(net1549),
    .Y(_0627_));
 sg13g2_nor2_1 _5765_ (.A(net875),
    .B(_0056_),
    .Y(_2369_));
 sg13g2_o21ai_1 _5766_ (.B1(net884),
    .Y(_2370_),
    .A1(net888),
    .A2(_0080_));
 sg13g2_nor3_1 _5767_ (.A(net812),
    .B(_2369_),
    .C(_2370_),
    .Y(_2371_));
 sg13g2_a221oi_1 _5768_ (.B2(net1627),
    .C1(_2371_),
    .B1(net802),
    .A1(net1240),
    .Y(_2372_),
    .A2(net814));
 sg13g2_nor2_1 _5769_ (.A(net907),
    .B(net1628),
    .Y(_0628_));
 sg13g2_nor2_1 _5770_ (.A(net875),
    .B(_0057_),
    .Y(_2373_));
 sg13g2_o21ai_1 _5771_ (.B1(net883),
    .Y(_2374_),
    .A1(net887),
    .A2(_0081_));
 sg13g2_nor3_1 _5772_ (.A(net815),
    .B(_2373_),
    .C(_2374_),
    .Y(_2375_));
 sg13g2_a221oi_1 _5773_ (.B2(net1604),
    .C1(_2375_),
    .B1(net802),
    .A1(net1251),
    .Y(_2376_),
    .A2(net815));
 sg13g2_nor2_1 _5774_ (.A(net907),
    .B(net1605),
    .Y(_0629_));
 sg13g2_nor2_1 _5775_ (.A(net875),
    .B(_0058_),
    .Y(_2377_));
 sg13g2_o21ai_1 _5776_ (.B1(net883),
    .Y(_2378_),
    .A1(net887),
    .A2(_0082_));
 sg13g2_nor3_1 _5777_ (.A(net812),
    .B(_2377_),
    .C(_2378_),
    .Y(_2379_));
 sg13g2_a221oi_1 _5778_ (.B2(net1622),
    .C1(_2379_),
    .B1(net802),
    .A1(net1296),
    .Y(_2380_),
    .A2(net815));
 sg13g2_nor2_1 _5779_ (.A(net907),
    .B(net1623),
    .Y(_0630_));
 sg13g2_nor2_1 _5780_ (.A(net875),
    .B(_0059_),
    .Y(_2381_));
 sg13g2_o21ai_1 _5781_ (.B1(net884),
    .Y(_2382_),
    .A1(net887),
    .A2(_0083_));
 sg13g2_nor3_1 _5782_ (.A(net814),
    .B(_2381_),
    .C(_2382_),
    .Y(_2383_));
 sg13g2_a221oi_1 _5783_ (.B2(net1659),
    .C1(_2383_),
    .B1(net804),
    .A1(net1282),
    .Y(_2384_),
    .A2(net814));
 sg13g2_nor2_1 _5784_ (.A(net909),
    .B(net1660),
    .Y(_0631_));
 sg13g2_nor2_1 _5785_ (.A(net875),
    .B(_0060_),
    .Y(_2385_));
 sg13g2_o21ai_1 _5786_ (.B1(net883),
    .Y(_2386_),
    .A1(net887),
    .A2(_0084_));
 sg13g2_nor3_1 _5787_ (.A(net814),
    .B(_2385_),
    .C(_2386_),
    .Y(_2387_));
 sg13g2_a221oi_1 _5788_ (.B2(net1636),
    .C1(_2387_),
    .B1(net804),
    .A1(net1187),
    .Y(_2388_),
    .A2(net814));
 sg13g2_nor2_1 _5789_ (.A(net909),
    .B(net1637),
    .Y(_0632_));
 sg13g2_a22oi_1 _5790_ (.Y(_2389_),
    .B1(net803),
    .B2(net1192),
    .A2(net819),
    .A1(net1053));
 sg13g2_nor2_1 _5791_ (.A(net909),
    .B(_2389_),
    .Y(_0633_));
 sg13g2_a22oi_1 _5792_ (.Y(_2390_),
    .B1(net803),
    .B2(net1240),
    .A2(net815),
    .A1(net985));
 sg13g2_nor2_1 _5793_ (.A(net902),
    .B(_2390_),
    .Y(_0634_));
 sg13g2_a22oi_1 _5794_ (.Y(_2391_),
    .B1(net803),
    .B2(net1251),
    .A2(net815),
    .A1(net1203));
 sg13g2_nor2_1 _5795_ (.A(net902),
    .B(_2391_),
    .Y(_0635_));
 sg13g2_o21ai_1 _5796_ (.B1(net949),
    .Y(_2392_),
    .A1(net1114),
    .A2(net823));
 sg13g2_a21oi_1 _5797_ (.A1(_0813_),
    .A2(net803),
    .Y(_0636_),
    .B1(_2392_));
 sg13g2_a221oi_1 _5798_ (.B2(_0812_),
    .C1(net909),
    .B1(net803),
    .A1(_0810_),
    .Y(_0637_),
    .A2(net819));
 sg13g2_o21ai_1 _5799_ (.B1(net957),
    .Y(_2393_),
    .A1(\output_value_inst.character_buff[5][6] ),
    .A2(net823));
 sg13g2_a21oi_1 _5800_ (.A1(_0811_),
    .A2(net803),
    .Y(_0638_),
    .B1(_2393_));
 sg13g2_a22oi_1 _5801_ (.Y(_2394_),
    .B1(net803),
    .B2(net1053),
    .A2(net815),
    .A1(\output_value_inst.character_buff[4][0] ));
 sg13g2_nor2_1 _5802_ (.A(net902),
    .B(net1054),
    .Y(_0639_));
 sg13g2_a22oi_1 _5803_ (.Y(_2395_),
    .B1(net803),
    .B2(net985),
    .A2(net815),
    .A1(\output_value_inst.character_buff[4][1] ));
 sg13g2_nor2_1 _5804_ (.A(net902),
    .B(net986),
    .Y(_0640_));
 sg13g2_a22oi_1 _5805_ (.Y(_2396_),
    .B1(net804),
    .B2(net1203),
    .A2(net816),
    .A1(net1046));
 sg13g2_nor2_1 _5806_ (.A(net903),
    .B(_2396_),
    .Y(_0641_));
 sg13g2_a22oi_1 _5807_ (.Y(_2397_),
    .B1(net804),
    .B2(net1114),
    .A2(net816),
    .A1(\output_value_inst.character_buff[4][3] ));
 sg13g2_nor2_1 _5808_ (.A(net902),
    .B(net1115),
    .Y(_0642_));
 sg13g2_a221oi_1 _5809_ (.B2(_0810_),
    .C1(net910),
    .B1(net806),
    .A1(_0809_),
    .Y(_0643_),
    .A2(net816));
 sg13g2_a22oi_1 _5810_ (.Y(_2398_),
    .B1(net805),
    .B2(net1229),
    .A2(net817),
    .A1(net970));
 sg13g2_nor2_1 _5811_ (.A(net903),
    .B(_2398_),
    .Y(_0644_));
 sg13g2_a22oi_1 _5812_ (.Y(_2399_),
    .B1(net805),
    .B2(net1214),
    .A2(net816),
    .A1(net1031));
 sg13g2_nor2_1 _5813_ (.A(net903),
    .B(_2399_),
    .Y(_0645_));
 sg13g2_a22oi_1 _5814_ (.Y(_2400_),
    .B1(net804),
    .B2(net1181),
    .A2(net816),
    .A1(net987));
 sg13g2_nor2_1 _5815_ (.A(net903),
    .B(_2400_),
    .Y(_0646_));
 sg13g2_a22oi_1 _5816_ (.Y(_2401_),
    .B1(net805),
    .B2(net1046),
    .A2(net817),
    .A1(net1012));
 sg13g2_nor2_1 _5817_ (.A(net903),
    .B(_2401_),
    .Y(_0647_));
 sg13g2_a22oi_1 _5818_ (.Y(_2402_),
    .B1(net805),
    .B2(net1258),
    .A2(net816),
    .A1(\output_value_inst.character_buff[3][3] ));
 sg13g2_nor2_1 _5819_ (.A(net902),
    .B(net1259),
    .Y(_0648_));
 sg13g2_a22oi_1 _5820_ (.Y(_2403_),
    .B1(net805),
    .B2(net1266),
    .A2(net817),
    .A1(net1081));
 sg13g2_nor2_1 _5821_ (.A(net910),
    .B(_2403_),
    .Y(_0649_));
 sg13g2_a221oi_1 _5822_ (.B2(_0809_),
    .C1(net909),
    .B1(net806),
    .A1(_0805_),
    .Y(_0650_),
    .A2(net816));
 sg13g2_a22oi_1 _5823_ (.Y(_2404_),
    .B1(net805),
    .B2(net970),
    .A2(net817),
    .A1(\output_value_inst.character_buff[3][6] ));
 sg13g2_nor2_1 _5824_ (.A(net902),
    .B(net971),
    .Y(_0651_));
 sg13g2_a22oi_1 _5825_ (.Y(_2405_),
    .B1(net805),
    .B2(net1031),
    .A2(net816),
    .A1(\output_value_inst.character_buff[2][0] ));
 sg13g2_nor2_1 _5826_ (.A(net910),
    .B(net1032),
    .Y(_0652_));
 sg13g2_o21ai_1 _5827_ (.B1(net957),
    .Y(_2406_),
    .A1(\output_value_inst.character_buff[2][1] ),
    .A2(net822));
 sg13g2_a21oi_1 _5828_ (.A1(_0808_),
    .A2(net807),
    .Y(_0653_),
    .B1(_2406_));
 sg13g2_a22oi_1 _5829_ (.Y(_2407_),
    .B1(net805),
    .B2(net1012),
    .A2(net817),
    .A1(\output_value_inst.character_buff[2][2] ));
 sg13g2_nor2_1 _5830_ (.A(net910),
    .B(net1013),
    .Y(_0654_));
 sg13g2_o21ai_1 _5831_ (.B1(net957),
    .Y(_2408_),
    .A1(net1136),
    .A2(net822));
 sg13g2_a21oi_1 _5832_ (.A1(_0807_),
    .A2(net807),
    .Y(_0655_),
    .B1(_2408_));
 sg13g2_o21ai_1 _5833_ (.B1(net957),
    .Y(_2409_),
    .A1(\output_value_inst.character_buff[2][4] ),
    .A2(net820));
 sg13g2_a21oi_1 _5834_ (.A1(_0806_),
    .A2(net806),
    .Y(_0656_),
    .B1(_2409_));
 sg13g2_o21ai_1 _5835_ (.B1(net957),
    .Y(_2410_),
    .A1(\output_value_inst.character_buff[2][5] ),
    .A2(net821));
 sg13g2_a21oi_1 _5836_ (.A1(_0805_),
    .A2(net806),
    .Y(_0657_),
    .B1(_2410_));
 sg13g2_a22oi_1 _5837_ (.Y(_2411_),
    .B1(net806),
    .B2(net1000),
    .A2(net818),
    .A1(\output_value_inst.character_buff[2][6] ));
 sg13g2_nor2_1 _5838_ (.A(net909),
    .B(net1001),
    .Y(_0658_));
 sg13g2_a21o_2 _5839_ (.A2(_0165_),
    .A1(net884),
    .B1(net814),
    .X(_2412_));
 sg13g2_a21oi_1 _5840_ (.A1(net877),
    .A2(net1497),
    .Y(_2413_),
    .B1(_2412_));
 sg13g2_o21ai_1 _5841_ (.B1(net957),
    .Y(_2414_),
    .A1(\output_value_inst.character_buff[1][0] ),
    .A2(net821));
 sg13g2_nor2_1 _5842_ (.A(net1498),
    .B(_2414_),
    .Y(_0659_));
 sg13g2_a21oi_1 _5843_ (.A1(net877),
    .A2(net1509),
    .Y(_2415_),
    .B1(_2412_));
 sg13g2_o21ai_1 _5844_ (.B1(net957),
    .Y(_2416_),
    .A1(net1440),
    .A2(net821));
 sg13g2_nor2_1 _5845_ (.A(net1510),
    .B(_2416_),
    .Y(_0660_));
 sg13g2_a21oi_1 _5846_ (.A1(net877),
    .A2(net1540),
    .Y(_2417_),
    .B1(_2307_));
 sg13g2_o21ai_1 _5847_ (.B1(net957),
    .Y(_2418_),
    .A1(net1145),
    .A2(net820));
 sg13g2_a21oi_1 _5848_ (.A1(net820),
    .A2(_2417_),
    .Y(_0661_),
    .B1(_2418_));
 sg13g2_a22oi_1 _5849_ (.Y(_2419_),
    .B1(net804),
    .B2(net1136),
    .A2(net818),
    .A1(\output_value_inst.character_buff[1][3] ));
 sg13g2_nor2_1 _5850_ (.A(net909),
    .B(net1137),
    .Y(_0662_));
 sg13g2_a21oi_1 _5851_ (.A1(net877),
    .A2(net1541),
    .Y(_2420_),
    .B1(_2412_));
 sg13g2_o21ai_1 _5852_ (.B1(net955),
    .Y(_2421_),
    .A1(net1457),
    .A2(net823));
 sg13g2_nor2_1 _5853_ (.A(net1542),
    .B(_2421_),
    .Y(_0663_));
 sg13g2_a22oi_1 _5854_ (.Y(_2422_),
    .B1(net807),
    .B2(net1316),
    .A2(net818),
    .A1(\output_value_inst.character_buff[1][5] ));
 sg13g2_nor2_1 _5855_ (.A(net909),
    .B(net1317),
    .Y(_0664_));
 sg13g2_o21ai_1 _5856_ (.B1(net956),
    .Y(_2423_),
    .A1(\output_value_inst.character_buff[1][6] ),
    .A2(net821));
 sg13g2_a21oi_1 _5857_ (.A1(_0804_),
    .A2(net806),
    .Y(_0665_),
    .B1(_2423_));
 sg13g2_a21oi_1 _5858_ (.A1(net878),
    .A2(net1513),
    .Y(_2424_),
    .B1(_2412_));
 sg13g2_o21ai_1 _5859_ (.B1(net956),
    .Y(_2425_),
    .A1(\output_value_inst.character_buff[0][0] ),
    .A2(net821));
 sg13g2_nor2_1 _5860_ (.A(net1514),
    .B(_2425_),
    .Y(_0666_));
 sg13g2_a21oi_1 _5861_ (.A1(net877),
    .A2(net1440),
    .Y(_2426_),
    .B1(_2412_));
 sg13g2_o21ai_1 _5862_ (.B1(net956),
    .Y(_2427_),
    .A1(\output_value_inst.character_buff[0][1] ),
    .A2(net820));
 sg13g2_nor2_1 _5863_ (.A(net1441),
    .B(_2427_),
    .Y(_0667_));
 sg13g2_o21ai_1 _5864_ (.B1(net955),
    .Y(_2428_),
    .A1(\output_value_inst.character_buff[0][2] ),
    .A2(net820));
 sg13g2_a21oi_1 _5865_ (.A1(_0803_),
    .A2(net806),
    .Y(_0668_),
    .B1(_2428_));
 sg13g2_a21oi_1 _5866_ (.A1(net877),
    .A2(\output_value_inst.character_buff[1][3] ),
    .Y(_2429_),
    .B1(_2307_));
 sg13g2_o21ai_1 _5867_ (.B1(net958),
    .Y(_2430_),
    .A1(net1580),
    .A2(net823));
 sg13g2_a21oi_1 _5868_ (.A1(net823),
    .A2(_2429_),
    .Y(_0669_),
    .B1(_2430_));
 sg13g2_a21oi_1 _5869_ (.A1(net877),
    .A2(net1457),
    .Y(_2431_),
    .B1(_2412_));
 sg13g2_o21ai_1 _5870_ (.B1(net955),
    .Y(_2432_),
    .A1(\output_value_inst.character_buff[0][4] ),
    .A2(net823));
 sg13g2_nor2_1 _5871_ (.A(net1458),
    .B(_2432_),
    .Y(_0670_));
 sg13g2_a21oi_1 _5872_ (.A1(net878),
    .A2(net1488),
    .Y(_2433_),
    .B1(_2412_));
 sg13g2_o21ai_1 _5873_ (.B1(net955),
    .Y(_2434_),
    .A1(\output_value_inst.character_buff[0][5] ),
    .A2(net820));
 sg13g2_nor2_1 _5874_ (.A(net1489),
    .B(_2434_),
    .Y(_0671_));
 sg13g2_a21oi_1 _5875_ (.A1(net877),
    .A2(\output_value_inst.character_buff[1][6] ),
    .Y(_2435_),
    .B1(_2307_));
 sg13g2_o21ai_1 _5876_ (.B1(net955),
    .Y(_2436_),
    .A1(net1567),
    .A2(net820));
 sg13g2_a21oi_1 _5877_ (.A1(net820),
    .A2(_2435_),
    .Y(_0672_),
    .B1(_2436_));
 sg13g2_nand3_1 _5878_ (.B(net889),
    .C(net1535),
    .A(net962),
    .Y(_2437_));
 sg13g2_o21ai_1 _5879_ (.B1(net956),
    .Y(_2438_),
    .A1(\output_value_inst.character_buff[0][0] ),
    .A2(net842));
 sg13g2_a21oi_1 _5880_ (.A1(_0802_),
    .A2(net842),
    .Y(_0673_),
    .B1(_2438_));
 sg13g2_o21ai_1 _5881_ (.B1(net956),
    .Y(_2439_),
    .A1(\output_value_inst.character_buff[0][1] ),
    .A2(net842));
 sg13g2_a21oi_1 _5882_ (.A1(_0801_),
    .A2(net842),
    .Y(_0674_),
    .B1(_2439_));
 sg13g2_o21ai_1 _5883_ (.B1(net955),
    .Y(_2440_),
    .A1(\output_value_inst.character_buff[0][2] ),
    .A2(net842));
 sg13g2_a21oi_1 _5884_ (.A1(_0800_),
    .A2(net842),
    .Y(_0675_),
    .B1(_2440_));
 sg13g2_o21ai_1 _5885_ (.B1(net958),
    .Y(_2441_),
    .A1(\output_value_inst.character_buff[0][3] ),
    .A2(net843));
 sg13g2_a21oi_1 _5886_ (.A1(_0799_),
    .A2(net843),
    .Y(_0676_),
    .B1(_2441_));
 sg13g2_o21ai_1 _5887_ (.B1(net958),
    .Y(_2442_),
    .A1(\output_value_inst.character_buff[0][4] ),
    .A2(net843));
 sg13g2_a21oi_1 _5888_ (.A1(_0798_),
    .A2(net843),
    .Y(_0677_),
    .B1(_2442_));
 sg13g2_o21ai_1 _5889_ (.B1(net955),
    .Y(_2443_),
    .A1(\output_value_inst.character_buff[0][5] ),
    .A2(net842));
 sg13g2_a21oi_1 _5890_ (.A1(_0797_),
    .A2(_2437_),
    .Y(_0678_),
    .B1(_2443_));
 sg13g2_o21ai_1 _5891_ (.B1(net955),
    .Y(_2444_),
    .A1(\output_value_inst.character_buff[0][6] ),
    .A2(net843));
 sg13g2_a21oi_1 _5892_ (.A1(_0796_),
    .A2(net842),
    .Y(_0679_),
    .B1(_2444_));
 sg13g2_nor2_1 _5893_ (.A(net887),
    .B(_2212_),
    .Y(_2445_));
 sg13g2_o21ai_1 _5894_ (.B1(net951),
    .Y(_2446_),
    .A1(net1047),
    .A2(net735));
 sg13g2_a21oi_1 _5895_ (.A1(net1047),
    .A2(_2445_),
    .Y(_0680_),
    .B1(_2446_));
 sg13g2_nand2_1 _5896_ (.Y(_2447_),
    .A(net963),
    .B(net887));
 sg13g2_o21ai_1 _5897_ (.B1(net951),
    .Y(_2448_),
    .A1(net1535),
    .A2(_2447_));
 sg13g2_a21oi_1 _5898_ (.A1(net875),
    .A2(_1094_),
    .Y(_0681_),
    .B1(_2448_));
 sg13g2_nor4_1 _5899_ (.A(\output_value_inst.character_buff[2][0] ),
    .B(\output_value_inst.character_buff[3][6] ),
    .C(\output_value_inst.character_buff[3][5] ),
    .D(\output_value_inst.character_buff[3][4] ),
    .Y(_2449_));
 sg13g2_nor4_1 _5900_ (.A(\output_value_inst.character_buff[2][4] ),
    .B(\output_value_inst.character_buff[2][3] ),
    .C(\output_value_inst.character_buff[2][2] ),
    .D(\output_value_inst.character_buff[2][1] ),
    .Y(_2450_));
 sg13g2_or4_1 _5901_ (.A(\output_value_inst.character_buff[3][3] ),
    .B(\output_value_inst.character_buff[3][2] ),
    .C(\output_value_inst.character_buff[3][1] ),
    .D(\output_value_inst.character_buff[3][0] ),
    .X(_2451_));
 sg13g2_nor4_1 _5902_ (.A(\output_value_inst.character_buff[4][6] ),
    .B(\output_value_inst.character_buff[4][4] ),
    .C(\output_value_inst.character_buff[4][3] ),
    .D(\output_value_inst.character_buff[4][2] ),
    .Y(_2452_));
 sg13g2_nand3_1 _5903_ (.B(_2450_),
    .C(_2452_),
    .A(_2449_),
    .Y(_2453_));
 sg13g2_nor4_1 _5904_ (.A(\output_value_inst.character_buff[0][2] ),
    .B(\output_value_inst.character_buff[0][1] ),
    .C(\output_value_inst.character_buff[0][0] ),
    .D(\output_value_inst.character_buff[1][6] ),
    .Y(_2454_));
 sg13g2_nor4_1 _5905_ (.A(\output_value_inst.character_buff[0][6] ),
    .B(\output_value_inst.character_buff[0][5] ),
    .C(\output_value_inst.character_buff[0][4] ),
    .D(\output_value_inst.character_buff[0][3] ),
    .Y(_2455_));
 sg13g2_nor4_1 _5906_ (.A(\output_value_inst.character_buff[1][5] ),
    .B(\output_value_inst.character_buff[1][4] ),
    .C(\output_value_inst.character_buff[1][3] ),
    .D(\output_value_inst.character_buff[1][2] ),
    .Y(_2456_));
 sg13g2_nor4_1 _5907_ (.A(\output_value_inst.character_buff[1][1] ),
    .B(\output_value_inst.character_buff[1][0] ),
    .C(\output_value_inst.character_buff[2][6] ),
    .D(\output_value_inst.character_buff[2][5] ),
    .Y(_2457_));
 sg13g2_nand4_1 _5908_ (.B(_2455_),
    .C(_2456_),
    .A(_2454_),
    .Y(_2458_),
    .D(_2457_));
 sg13g2_nor4_1 _5909_ (.A(\output_value_inst.character_buff[5][3] ),
    .B(\output_value_inst.character_buff[5][2] ),
    .C(\output_value_inst.character_buff[5][1] ),
    .D(\output_value_inst.character_buff[5][0] ),
    .Y(_2459_));
 sg13g2_nor4_1 _5910_ (.A(\output_value_inst.character_buff[4][1] ),
    .B(\output_value_inst.character_buff[4][0] ),
    .C(\output_value_inst.character_buff[5][6] ),
    .D(\output_value_inst.character_buff[5][4] ),
    .Y(_2460_));
 sg13g2_and2_1 _5911_ (.A(_2459_),
    .B(_2460_),
    .X(_2461_));
 sg13g2_nor4_1 _5912_ (.A(\output_value_inst.character_buff[6][6] ),
    .B(\output_value_inst.character_buff[6][4] ),
    .C(\output_value_inst.character_buff[6][3] ),
    .D(net1771),
    .Y(_2462_));
 sg13g2_nor4_1 _5913_ (.A(\output_value_inst.character_buff[6][1] ),
    .B(\output_value_inst.character_buff[6][0] ),
    .C(\output_value_inst.character_buff[7][6] ),
    .D(\output_value_inst.character_buff[7][4] ),
    .Y(_2463_));
 sg13g2_nor4_1 _5914_ (.A(\output_value_inst.character_buff[9][6] ),
    .B(\output_value_inst.character_buff[9][4] ),
    .C(\output_value_inst.character_buff[9][3] ),
    .D(\output_value_inst.character_buff[9][2] ),
    .Y(_2464_));
 sg13g2_nor4_1 _5915_ (.A(\output_value_inst.character_buff[7][3] ),
    .B(\output_value_inst.character_buff[7][2] ),
    .C(\output_value_inst.character_buff[7][1] ),
    .D(\output_value_inst.character_buff[7][0] ),
    .Y(_2465_));
 sg13g2_and2_1 _5916_ (.A(_2464_),
    .B(_2465_),
    .X(_2466_));
 sg13g2_nor4_1 _5917_ (.A(\output_value_inst.character_buff[9][1] ),
    .B(\output_value_inst.character_buff[9][0] ),
    .C(\output_value_inst.character_buff[8][6] ),
    .D(\output_value_inst.character_buff[8][4] ),
    .Y(_2467_));
 sg13g2_nor4_1 _5918_ (.A(\output_value_inst.character_buff[8][3] ),
    .B(\output_value_inst.character_buff[8][2] ),
    .C(\output_value_inst.character_buff[8][1] ),
    .D(\output_value_inst.character_buff[8][0] ),
    .Y(_2468_));
 sg13g2_nand3_1 _5919_ (.B(_2467_),
    .C(_2468_),
    .A(_2466_),
    .Y(_2469_));
 sg13g2_nor4_1 _5920_ (.A(_2451_),
    .B(_2453_),
    .C(_2458_),
    .D(_2469_),
    .Y(_2470_));
 sg13g2_nand4_1 _5921_ (.B(net1772),
    .C(_2463_),
    .A(_2461_),
    .Y(_2471_),
    .D(_2470_));
 sg13g2_nor3_1 _5922_ (.A(net883),
    .B(net1704),
    .C(_2471_),
    .Y(_2472_));
 sg13g2_nor3_1 _5923_ (.A(net878),
    .B(net887),
    .C(net1047),
    .Y(_2473_));
 sg13g2_nor3_1 _5924_ (.A(_0985_),
    .B(_2472_),
    .C(_2473_),
    .Y(_2474_));
 sg13g2_a21oi_1 _5925_ (.A1(net878),
    .A2(net872),
    .Y(_0682_),
    .B1(_2474_));
 sg13g2_mux2_1 _5926_ (.A0(_0792_),
    .A1(_1260_),
    .S(net734),
    .X(_2475_));
 sg13g2_nor2_1 _5927_ (.A(net895),
    .B(_2475_),
    .Y(_0683_));
 sg13g2_nand2b_1 _5928_ (.Y(_2476_),
    .B(net1028),
    .A_N(net734));
 sg13g2_a21oi_1 _5929_ (.A1(_1374_),
    .A2(_2476_),
    .Y(_0684_),
    .B1(net896));
 sg13g2_nand2b_1 _5930_ (.Y(_2477_),
    .B(net978),
    .A_N(net735));
 sg13g2_a21oi_1 _5931_ (.A1(_1377_),
    .A2(_2477_),
    .Y(_0685_),
    .B1(net906));
 sg13g2_nand2b_1 _5932_ (.Y(_2478_),
    .B(net984),
    .A_N(net734));
 sg13g2_a21oi_1 _5933_ (.A1(_1371_),
    .A2(_2478_),
    .Y(_0686_),
    .B1(net906));
 sg13g2_nand2b_1 _5934_ (.Y(_2479_),
    .B(net1033),
    .A_N(net732));
 sg13g2_a21oi_1 _5935_ (.A1(_1299_),
    .A2(_2479_),
    .Y(_0687_),
    .B1(net896));
 sg13g2_nand2b_1 _5936_ (.Y(_2480_),
    .B(net1014),
    .A_N(net733));
 sg13g2_a21oi_1 _5937_ (.A1(_1293_),
    .A2(_2480_),
    .Y(_0688_),
    .B1(net898));
 sg13g2_nand2b_1 _5938_ (.Y(_2481_),
    .B(net715),
    .A_N(net732));
 sg13g2_a21oi_1 _5939_ (.A1(_1296_),
    .A2(_2481_),
    .Y(_0689_),
    .B1(net895));
 sg13g2_o21ai_1 _5940_ (.B1(net939),
    .Y(_2482_),
    .A1(net1522),
    .A2(net730));
 sg13g2_a21oi_1 _5941_ (.A1(_0791_),
    .A2(net730),
    .Y(_0690_),
    .B1(_2482_));
 sg13g2_o21ai_1 _5942_ (.B1(net938),
    .Y(_2483_),
    .A1(net1583),
    .A2(net731));
 sg13g2_a21oi_1 _5943_ (.A1(_0790_),
    .A2(net731),
    .Y(_0691_),
    .B1(_2483_));
 sg13g2_o21ai_1 _5944_ (.B1(net941),
    .Y(_2484_),
    .A1(net1465),
    .A2(net731));
 sg13g2_a21oi_1 _5945_ (.A1(_0788_),
    .A2(net730),
    .Y(_0694_),
    .B1(_2484_));
 sg13g2_o21ai_1 _5946_ (.B1(net949),
    .Y(_2485_),
    .A1(\Led_Cycle_inst.genblk1[0].pwm_unit.pwm_out ),
    .A2(net793));
 sg13g2_a21oi_1 _5947_ (.A1(_0787_),
    .A2(net793),
    .Y(_0695_),
    .B1(_2485_));
 sg13g2_o21ai_1 _5948_ (.B1(net945),
    .Y(_2486_),
    .A1(\Led_Cycle_inst.genblk1[3].pwm_unit.pwm_out ),
    .A2(net794));
 sg13g2_a21oi_1 _5949_ (.A1(_0782_),
    .A2(net794),
    .Y(_0698_),
    .B1(_2486_));
 sg13g2_o21ai_1 _5950_ (.B1(net946),
    .Y(_2487_),
    .A1(\Led_Cycle_inst.genblk1[4].pwm_unit.pwm_out ),
    .A2(net790));
 sg13g2_a21oi_1 _5951_ (.A1(_0781_),
    .A2(net790),
    .Y(_0699_),
    .B1(_2487_));
 sg13g2_o21ai_1 _5952_ (.B1(net923),
    .Y(_2488_),
    .A1(\Led_Cycle_inst.genblk1[7].pwm_unit.pwm_out ),
    .A2(net789));
 sg13g2_a21oi_1 _5953_ (.A1(_0779_),
    .A2(net789),
    .Y(_0702_),
    .B1(_2488_));
 sg13g2_o21ai_1 _5954_ (.B1(net922),
    .Y(_2489_),
    .A1(\Led_Cycle_inst.genblk1[8].pwm_unit.pwm_out ),
    .A2(net788));
 sg13g2_a21oi_1 _5955_ (.A1(_0778_),
    .A2(net788),
    .Y(_0703_),
    .B1(_2489_));
 sg13g2_o21ai_1 _5956_ (.B1(net922),
    .Y(_2490_),
    .A1(\Led_Cycle_inst.genblk1[11].pwm_unit.pwm_out ),
    .A2(net788));
 sg13g2_a21oi_1 _5957_ (.A1(_0776_),
    .A2(net788),
    .Y(_0706_),
    .B1(_2490_));
 sg13g2_o21ai_1 _5958_ (.B1(net946),
    .Y(_2491_),
    .A1(\Led_Cycle_inst.genblk1[12].pwm_unit.pwm_out ),
    .A2(net789));
 sg13g2_a21oi_1 _5959_ (.A1(_0775_),
    .A2(net789),
    .Y(_0707_),
    .B1(_2491_));
 sg13g2_o21ai_1 _5960_ (.B1(net945),
    .Y(_2492_),
    .A1(\Led_Cycle_inst.genblk1[15].pwm_unit.pwm_out ),
    .A2(net792));
 sg13g2_a21oi_1 _5961_ (.A1(_0772_),
    .A2(net792),
    .Y(_0710_),
    .B1(_2492_));
 sg13g2_o21ai_1 _5962_ (.B1(net951),
    .Y(_2493_),
    .A1(net843),
    .A2(net1773));
 sg13g2_a21oi_1 _5963_ (.A1(_0771_),
    .A2(net843),
    .Y(_0711_),
    .B1(_2493_));
 sg13g2_a22oi_1 _5964_ (.Y(_2494_),
    .B1(_2205_),
    .B2(net1200),
    .A2(_2180_),
    .A1(net1026));
 sg13g2_nor2_2 _5965_ (.A(_1414_),
    .B(_2249_),
    .Y(_2495_));
 sg13g2_nor2_1 _5966_ (.A(_2494_),
    .B(_2495_),
    .Y(_0712_));
 sg13g2_a22oi_1 _5967_ (.Y(_2496_),
    .B1(_2205_),
    .B2(net992),
    .A2(_2180_),
    .A1(net713));
 sg13g2_nor2_1 _5968_ (.A(_2495_),
    .B(_2496_),
    .Y(_0713_));
 sg13g2_a22oi_1 _5969_ (.Y(_2497_),
    .B1(_2205_),
    .B2(net1087),
    .A2(net825),
    .A1(net972));
 sg13g2_nor2_1 _5970_ (.A(_2495_),
    .B(_2497_),
    .Y(_0714_));
 sg13g2_a22oi_1 _5971_ (.Y(_2498_),
    .B1(_2205_),
    .B2(net1118),
    .A2(net825),
    .A1(net716));
 sg13g2_nor2_1 _5972_ (.A(_2495_),
    .B(_2498_),
    .Y(_0715_));
 sg13g2_a22oi_1 _5973_ (.Y(_2499_),
    .B1(_2205_),
    .B2(net1059),
    .A2(net825),
    .A1(net688));
 sg13g2_nor2_1 _5974_ (.A(_2495_),
    .B(_2499_),
    .Y(_0716_));
 sg13g2_a22oi_1 _5975_ (.Y(_2500_),
    .B1(_2205_),
    .B2(net1132),
    .A2(net825),
    .A1(net722));
 sg13g2_nor2_1 _5976_ (.A(_2495_),
    .B(_2500_),
    .Y(_0717_));
 sg13g2_a22oi_1 _5977_ (.Y(_2501_),
    .B1(_2205_),
    .B2(net1133),
    .A2(net825),
    .A1(net707));
 sg13g2_nor2_1 _5978_ (.A(_2495_),
    .B(_2501_),
    .Y(_0718_));
 sg13g2_nor3_1 _5979_ (.A(net1657),
    .B(_1097_),
    .C(_0697_),
    .Y(_0719_));
 sg13g2_o21ai_1 _5980_ (.B1(net959),
    .Y(_2502_),
    .A1(\uart_inst.uart_tx_inst.DATA_REG[0] ),
    .A2(net763));
 sg13g2_a21oi_1 _5981_ (.A1(_0770_),
    .A2(net762),
    .Y(_0721_),
    .B1(_2502_));
 sg13g2_o21ai_1 _5982_ (.B1(net960),
    .Y(_2503_),
    .A1(\uart_inst.uart_tx_inst.DATA_REG[1] ),
    .A2(net763));
 sg13g2_a21oi_1 _5983_ (.A1(_0769_),
    .A2(net762),
    .Y(_0722_),
    .B1(_2503_));
 sg13g2_o21ai_1 _5984_ (.B1(net959),
    .Y(_2504_),
    .A1(\uart_inst.uart_tx_inst.DATA_REG[2] ),
    .A2(net763));
 sg13g2_a21oi_1 _5985_ (.A1(_0768_),
    .A2(net762),
    .Y(_0723_),
    .B1(_2504_));
 sg13g2_o21ai_1 _5986_ (.B1(net959),
    .Y(_2505_),
    .A1(net1386),
    .A2(net763));
 sg13g2_a21oi_1 _5987_ (.A1(_0767_),
    .A2(net762),
    .Y(_0724_),
    .B1(_2505_));
 sg13g2_o21ai_1 _5988_ (.B1(net952),
    .Y(_2506_),
    .A1(\uart_inst.uart_tx_inst.DATA_REG[4] ),
    .A2(net762));
 sg13g2_a21oi_1 _5989_ (.A1(_0766_),
    .A2(net762),
    .Y(_0725_),
    .B1(_2506_));
 sg13g2_o21ai_1 _5990_ (.B1(net952),
    .Y(_2507_),
    .A1(\uart_inst.uart_tx_inst.DATA_REG[5] ),
    .A2(net762));
 sg13g2_a21oi_1 _5991_ (.A1(_0765_),
    .A2(net762),
    .Y(_0726_),
    .B1(_2507_));
 sg13g2_o21ai_1 _5992_ (.B1(net952),
    .Y(_2508_),
    .A1(\uart_inst.uart_tx_inst.DATA_REG[6] ),
    .A2(net764));
 sg13g2_a21oi_1 _5993_ (.A1(_0764_),
    .A2(net764),
    .Y(_0727_),
    .B1(_2508_));
 sg13g2_nor2_1 _5994_ (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[0] ),
    .B(net1559),
    .Y(_2509_));
 sg13g2_nor4_1 _5995_ (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[12] ),
    .B(\SegmentDisplay.seg_driver.clk_reducer.counter[3] ),
    .C(\SegmentDisplay.seg_driver.clk_reducer.counter[2] ),
    .D(\SegmentDisplay.seg_driver.clk_reducer.counter[5] ),
    .Y(_2510_));
 sg13g2_nor3_1 _5996_ (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[8] ),
    .B(\SegmentDisplay.seg_driver.clk_reducer.counter[11] ),
    .C(\SegmentDisplay.seg_driver.clk_reducer.counter[10] ),
    .Y(_2511_));
 sg13g2_nor4_1 _5997_ (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[4] ),
    .B(\SegmentDisplay.seg_driver.clk_reducer.counter[7] ),
    .C(\SegmentDisplay.seg_driver.clk_reducer.counter[6] ),
    .D(\SegmentDisplay.seg_driver.clk_reducer.counter[9] ),
    .Y(_2512_));
 sg13g2_nand4_1 _5998_ (.B(_2510_),
    .C(_2511_),
    .A(_2509_),
    .Y(_2513_),
    .D(_2512_));
 sg13g2_nand2_2 _5999_ (.Y(_2514_),
    .A(net918),
    .B(_2513_));
 sg13g2_and3_1 _6000_ (.X(_0728_),
    .A(net918),
    .B(net633),
    .C(_2513_));
 sg13g2_and2_1 _6001_ (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[0] ),
    .B(net1559),
    .X(_2515_));
 sg13g2_nor3_1 _6002_ (.A(net891),
    .B(net1560),
    .C(_2515_),
    .Y(_0729_));
 sg13g2_xnor2_1 _6003_ (.Y(_2516_),
    .A(net1516),
    .B(_2515_));
 sg13g2_nor2_1 _6004_ (.A(_2514_),
    .B(net1517),
    .Y(_0730_));
 sg13g2_and4_1 _6005_ (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[0] ),
    .B(\SegmentDisplay.seg_driver.clk_reducer.counter[1] ),
    .C(net1074),
    .D(\SegmentDisplay.seg_driver.clk_reducer.counter[2] ),
    .X(_2517_));
 sg13g2_a21oi_1 _6006_ (.A1(\SegmentDisplay.seg_driver.clk_reducer.counter[2] ),
    .A2(_2515_),
    .Y(_2518_),
    .B1(net1074));
 sg13g2_nor3_1 _6007_ (.A(_2514_),
    .B(_2517_),
    .C(net1075),
    .Y(_0731_));
 sg13g2_and2_1 _6008_ (.A(net1354),
    .B(_2517_),
    .X(_2519_));
 sg13g2_nor2_1 _6009_ (.A(net1354),
    .B(_2517_),
    .Y(_2520_));
 sg13g2_nor3_1 _6010_ (.A(net799),
    .B(_2519_),
    .C(net1355),
    .Y(_0732_));
 sg13g2_and2_1 _6011_ (.A(net1293),
    .B(_2519_),
    .X(_2521_));
 sg13g2_nor2_1 _6012_ (.A(net1293),
    .B(_2519_),
    .Y(_2522_));
 sg13g2_nor3_1 _6013_ (.A(net799),
    .B(_2521_),
    .C(net1294),
    .Y(_0733_));
 sg13g2_xnor2_1 _6014_ (.Y(_2523_),
    .A(net1524),
    .B(_2521_));
 sg13g2_nor2_1 _6015_ (.A(net799),
    .B(_2523_),
    .Y(_0734_));
 sg13g2_a21oi_1 _6016_ (.A1(\SegmentDisplay.seg_driver.clk_reducer.counter[6] ),
    .A2(_2521_),
    .Y(_2524_),
    .B1(net1139));
 sg13g2_and3_1 _6017_ (.X(_2525_),
    .A(net1139),
    .B(\SegmentDisplay.seg_driver.clk_reducer.counter[6] ),
    .C(_2521_));
 sg13g2_nor3_1 _6018_ (.A(net799),
    .B(net1140),
    .C(_2525_),
    .Y(_0735_));
 sg13g2_nor2_1 _6019_ (.A(net1359),
    .B(_2525_),
    .Y(_2526_));
 sg13g2_and2_1 _6020_ (.A(net1359),
    .B(_2525_),
    .X(_2527_));
 sg13g2_nor3_1 _6021_ (.A(net799),
    .B(net1360),
    .C(_2527_),
    .Y(_0736_));
 sg13g2_nor2_1 _6022_ (.A(net1376),
    .B(_2527_),
    .Y(_2528_));
 sg13g2_and2_1 _6023_ (.A(net1376),
    .B(_2527_),
    .X(_2529_));
 sg13g2_nor3_1 _6024_ (.A(net799),
    .B(_2528_),
    .C(_2529_),
    .Y(_0737_));
 sg13g2_nor2_1 _6025_ (.A(net1422),
    .B(_2529_),
    .Y(_2530_));
 sg13g2_and2_1 _6026_ (.A(net1422),
    .B(_2529_),
    .X(_2531_));
 sg13g2_nor3_1 _6027_ (.A(net799),
    .B(_2530_),
    .C(_2531_),
    .Y(_0738_));
 sg13g2_nor2_1 _6028_ (.A(net1392),
    .B(_2531_),
    .Y(_2532_));
 sg13g2_and2_1 _6029_ (.A(net1392),
    .B(_2531_),
    .X(_2533_));
 sg13g2_nor3_1 _6030_ (.A(_2514_),
    .B(net1393),
    .C(_2533_),
    .Y(_0739_));
 sg13g2_nor2_1 _6031_ (.A(net1409),
    .B(_2533_),
    .Y(_2534_));
 sg13g2_a21oi_1 _6032_ (.A1(net1409),
    .A2(_2533_),
    .Y(_2535_),
    .B1(net799));
 sg13g2_nor2b_1 _6033_ (.A(_2534_),
    .B_N(_2535_),
    .Y(_0740_));
 sg13g2_and2_2 _6034_ (.A(net918),
    .B(net981),
    .X(_0741_));
 sg13g2_and3_1 _6035_ (.X(_2536_),
    .A(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[0] ),
    .B(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[1] ),
    .C(net1127));
 sg13g2_and2_1 _6036_ (.A(net1414),
    .B(_2536_),
    .X(_2537_));
 sg13g2_nand2_1 _6037_ (.Y(_2538_),
    .A(net1685),
    .B(_2537_));
 sg13g2_o21ai_1 _6038_ (.B1(net921),
    .Y(_2539_),
    .A1(_0911_),
    .A2(_2538_));
 sg13g2_nor2_1 _6039_ (.A(_0947_),
    .B(_2539_),
    .Y(_0742_));
 sg13g2_or2_1 _6040_ (.X(_2540_),
    .B(net1716),
    .A(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[0] ));
 sg13g2_and3_1 _6041_ (.X(_0743_),
    .A(net920),
    .B(net1717),
    .C(_2540_));
 sg13g2_a21oi_1 _6042_ (.A1(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[0] ),
    .A2(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[1] ),
    .Y(_2541_),
    .B1(net1127));
 sg13g2_nor3_1 _6043_ (.A(net892),
    .B(_2536_),
    .C(net1128),
    .Y(_0744_));
 sg13g2_o21ai_1 _6044_ (.B1(net920),
    .Y(_2542_),
    .A1(net1414),
    .A2(_2536_));
 sg13g2_nor2_1 _6045_ (.A(_2537_),
    .B(net1415),
    .Y(_0745_));
 sg13g2_or2_1 _6046_ (.X(_2543_),
    .B(_2537_),
    .A(net1685));
 sg13g2_and3_1 _6047_ (.X(_0746_),
    .A(net921),
    .B(_2538_),
    .C(_2543_));
 sg13g2_a21oi_1 _6048_ (.A1(_0911_),
    .A2(_2538_),
    .Y(_0747_),
    .B1(_2539_));
 sg13g2_a22oi_1 _6049_ (.Y(_2544_),
    .B1(net757),
    .B2(net718),
    .A2(net760),
    .A1(\uart_tx_fifo_inst.fifo[7][0] ));
 sg13g2_a21oi_1 _6050_ (.A1(_0895_),
    .A2(net770),
    .Y(_2545_),
    .B1(_1423_));
 sg13g2_o21ai_1 _6051_ (.B1(_2545_),
    .Y(_2546_),
    .A1(net1174),
    .A2(net770));
 sg13g2_a22oi_1 _6052_ (.Y(_2547_),
    .B1(net757),
    .B2(\uart_tx_fifo_inst.fifo[2][0] ),
    .A2(net760),
    .A1(net1520));
 sg13g2_inv_1 _6053_ (.Y(_2548_),
    .A(_2547_));
 sg13g2_a221oi_1 _6054_ (.B2(\uart_tx_fifo_inst.fifo[1][0] ),
    .C1(_2548_),
    .B1(net737),
    .A1(\uart_tx_fifo_inst.fifo[0][0] ),
    .Y(_2549_),
    .A2(net741));
 sg13g2_o21ai_1 _6055_ (.B1(_2546_),
    .Y(_2550_),
    .A1(_2249_),
    .A2(_2549_));
 sg13g2_a22oi_1 _6056_ (.Y(_2551_),
    .B1(net737),
    .B2(net1265),
    .A2(net742),
    .A1(\uart_tx_fifo_inst.fifo[4][0] ));
 sg13g2_nand2_1 _6057_ (.Y(_2552_),
    .A(_2544_),
    .B(_2551_));
 sg13g2_a22oi_1 _6058_ (.Y(_2553_),
    .B1(_2274_),
    .B2(_2552_),
    .A2(net739),
    .A1(net1350));
 sg13g2_nand2b_1 _6059_ (.Y(_0748_),
    .B(_2553_),
    .A_N(_2550_));
 sg13g2_a22oi_1 _6060_ (.Y(_2554_),
    .B1(net757),
    .B2(net1006),
    .A2(net759),
    .A1(net1112));
 sg13g2_a21oi_1 _6061_ (.A1(_0894_),
    .A2(net769),
    .Y(_2555_),
    .B1(_1423_));
 sg13g2_o21ai_1 _6062_ (.B1(_2555_),
    .Y(_2556_),
    .A1(net1201),
    .A2(net769));
 sg13g2_a22oi_1 _6063_ (.Y(_2557_),
    .B1(net757),
    .B2(\uart_tx_fifo_inst.fifo[2][1] ),
    .A2(net760),
    .A1(\uart_tx_fifo_inst.fifo[3][1] ));
 sg13g2_inv_1 _6064_ (.Y(_2558_),
    .A(_2557_));
 sg13g2_a221oi_1 _6065_ (.B2(\uart_tx_fifo_inst.fifo[1][1] ),
    .C1(_2558_),
    .B1(net737),
    .A1(\uart_tx_fifo_inst.fifo[0][1] ),
    .Y(_2559_),
    .A2(net741));
 sg13g2_o21ai_1 _6066_ (.B1(_2556_),
    .Y(_2560_),
    .A1(_2249_),
    .A2(_2559_));
 sg13g2_a22oi_1 _6067_ (.Y(_2561_),
    .B1(net736),
    .B2(net1281),
    .A2(net742),
    .A1(net1425));
 sg13g2_nand2_1 _6068_ (.Y(_2562_),
    .A(_2554_),
    .B(_2561_));
 sg13g2_a22oi_1 _6069_ (.Y(_2563_),
    .B1(_2274_),
    .B2(_2562_),
    .A2(net739),
    .A1(net1320));
 sg13g2_nand2b_1 _6070_ (.Y(_0749_),
    .B(_2563_),
    .A_N(_2560_));
 sg13g2_a22oi_1 _6071_ (.Y(_2564_),
    .B1(net756),
    .B2(\uart_tx_fifo_inst.fifo[6][2] ),
    .A2(net759),
    .A1(\uart_tx_fifo_inst.fifo[7][2] ));
 sg13g2_inv_1 _6072_ (.Y(_2565_),
    .A(_2564_));
 sg13g2_a221oi_1 _6073_ (.B2(\uart_tx_fifo_inst.fifo[5][2] ),
    .C1(_2565_),
    .B1(net736),
    .A1(\uart_tx_fifo_inst.fifo[4][2] ),
    .Y(_2566_),
    .A2(net741));
 sg13g2_nand2b_1 _6074_ (.Y(_2567_),
    .B(_2190_),
    .A_N(_2566_));
 sg13g2_o21ai_1 _6075_ (.B1(_1422_),
    .Y(_2568_),
    .A1(net1107),
    .A2(net769));
 sg13g2_a21oi_1 _6076_ (.A1(_0893_),
    .A2(net769),
    .Y(_2569_),
    .B1(_2568_));
 sg13g2_nand2_1 _6077_ (.Y(_2570_),
    .A(\uart_tx_fifo_inst.fifo[1][2] ),
    .B(net736));
 sg13g2_and2_1 _6078_ (.A(\uart_tx_fifo_inst.fifo[3][2] ),
    .B(net759),
    .X(_2571_));
 sg13g2_a221oi_1 _6079_ (.B2(\uart_tx_fifo_inst.fifo[2][2] ),
    .C1(_2571_),
    .B1(net756),
    .A1(\uart_tx_fifo_inst.fifo[0][2] ),
    .Y(_2572_),
    .A2(net741));
 sg13g2_a21oi_1 _6080_ (.A1(_2570_),
    .A2(_2572_),
    .Y(_2573_),
    .B1(_2177_));
 sg13g2_nor3_1 _6081_ (.A(net740),
    .B(_2569_),
    .C(_2573_),
    .Y(_2574_));
 sg13g2_a22oi_1 _6082_ (.Y(_0750_),
    .B1(_2567_),
    .B2(_2574_),
    .A2(net739),
    .A1(_0768_));
 sg13g2_a22oi_1 _6083_ (.Y(_2575_),
    .B1(net756),
    .B2(\uart_tx_fifo_inst.fifo[6][3] ),
    .A2(net759),
    .A1(\uart_tx_fifo_inst.fifo[7][3] ));
 sg13g2_inv_1 _6084_ (.Y(_2576_),
    .A(_2575_));
 sg13g2_a221oi_1 _6085_ (.B2(\uart_tx_fifo_inst.fifo[5][3] ),
    .C1(_2576_),
    .B1(net736),
    .A1(\uart_tx_fifo_inst.fifo[4][3] ),
    .Y(_2577_),
    .A2(net741));
 sg13g2_nand2b_1 _6086_ (.Y(_2578_),
    .B(_2190_),
    .A_N(_2577_));
 sg13g2_o21ai_1 _6087_ (.B1(_1422_),
    .Y(_2579_),
    .A1(\uart_tx_fifo_inst.fifo[8][3] ),
    .A2(_1407_));
 sg13g2_a21oi_1 _6088_ (.A1(_0763_),
    .A2(_1407_),
    .Y(_2580_),
    .B1(_2579_));
 sg13g2_nand2_1 _6089_ (.Y(_2581_),
    .A(\uart_tx_fifo_inst.fifo[1][3] ),
    .B(net738));
 sg13g2_and2_1 _6090_ (.A(\uart_tx_fifo_inst.fifo[3][3] ),
    .B(net761),
    .X(_2582_));
 sg13g2_a221oi_1 _6091_ (.B2(\uart_tx_fifo_inst.fifo[2][3] ),
    .C1(_2582_),
    .B1(net758),
    .A1(\uart_tx_fifo_inst.fifo[0][3] ),
    .Y(_2583_),
    .A2(net743));
 sg13g2_a21oi_1 _6092_ (.A1(_2581_),
    .A2(_2583_),
    .Y(_2584_),
    .B1(_2177_));
 sg13g2_nor3_1 _6093_ (.A(net739),
    .B(_2580_),
    .C(_2584_),
    .Y(_2585_));
 sg13g2_a22oi_1 _6094_ (.Y(_0751_),
    .B1(_2578_),
    .B2(_2585_),
    .A2(net739),
    .A1(_0767_));
 sg13g2_a22oi_1 _6095_ (.Y(_2586_),
    .B1(net756),
    .B2(\uart_tx_fifo_inst.fifo[6][4] ),
    .A2(net759),
    .A1(\uart_tx_fifo_inst.fifo[7][4] ));
 sg13g2_inv_1 _6096_ (.Y(_2587_),
    .A(_2586_));
 sg13g2_a221oi_1 _6097_ (.B2(\uart_tx_fifo_inst.fifo[5][4] ),
    .C1(_2587_),
    .B1(net736),
    .A1(\uart_tx_fifo_inst.fifo[4][4] ),
    .Y(_2588_),
    .A2(net741));
 sg13g2_nand2b_1 _6098_ (.Y(_2589_),
    .B(_2190_),
    .A_N(_2588_));
 sg13g2_nand2_1 _6099_ (.Y(_2590_),
    .A(\uart_tx_fifo_inst.fifo[0][4] ),
    .B(net743));
 sg13g2_and2_1 _6100_ (.A(\uart_tx_fifo_inst.fifo[3][4] ),
    .B(net761),
    .X(_2591_));
 sg13g2_a221oi_1 _6101_ (.B2(\uart_tx_fifo_inst.fifo[2][4] ),
    .C1(_2591_),
    .B1(net758),
    .A1(\uart_tx_fifo_inst.fifo[1][4] ),
    .Y(_2592_),
    .A2(net738));
 sg13g2_a21oi_1 _6102_ (.A1(_2590_),
    .A2(_2592_),
    .Y(_2593_),
    .B1(_2177_));
 sg13g2_o21ai_1 _6103_ (.B1(_1422_),
    .Y(_2594_),
    .A1(net1196),
    .A2(net769));
 sg13g2_a21oi_1 _6104_ (.A1(_0892_),
    .A2(net769),
    .Y(_2595_),
    .B1(_2594_));
 sg13g2_nor3_1 _6105_ (.A(net740),
    .B(_2593_),
    .C(_2595_),
    .Y(_2596_));
 sg13g2_a22oi_1 _6106_ (.Y(_0752_),
    .B1(_2589_),
    .B2(_2596_),
    .A2(net739),
    .A1(_0766_));
 sg13g2_nand2_1 _6107_ (.Y(_2597_),
    .A(net1372),
    .B(net741));
 sg13g2_and2_1 _6108_ (.A(\uart_tx_fifo_inst.fifo[3][5] ),
    .B(net760),
    .X(_2598_));
 sg13g2_a221oi_1 _6109_ (.B2(\uart_tx_fifo_inst.fifo[2][5] ),
    .C1(_2598_),
    .B1(net756),
    .A1(\uart_tx_fifo_inst.fifo[1][5] ),
    .Y(_2599_),
    .A2(net737));
 sg13g2_a21oi_1 _6110_ (.A1(_2597_),
    .A2(_2599_),
    .Y(_2600_),
    .B1(_2177_));
 sg13g2_o21ai_1 _6111_ (.B1(_1422_),
    .Y(_2601_),
    .A1(\uart_tx_fifo_inst.fifo[8][5] ),
    .A2(_1407_));
 sg13g2_a21oi_1 _6112_ (.A1(_0762_),
    .A2(_1407_),
    .Y(_2602_),
    .B1(_2601_));
 sg13g2_nor2_1 _6113_ (.A(_2600_),
    .B(_2602_),
    .Y(_2603_));
 sg13g2_nand2_1 _6114_ (.Y(_2604_),
    .A(net1170),
    .B(net736));
 sg13g2_nand2_1 _6115_ (.Y(_2605_),
    .A(\uart_tx_fifo_inst.fifo[4][5] ),
    .B(net741));
 sg13g2_a22oi_1 _6116_ (.Y(_2606_),
    .B1(net756),
    .B2(\uart_tx_fifo_inst.fifo[6][5] ),
    .A2(net759),
    .A1(\uart_tx_fifo_inst.fifo[7][5] ));
 sg13g2_nand3_1 _6117_ (.B(_2605_),
    .C(_2606_),
    .A(_2604_),
    .Y(_2607_));
 sg13g2_a22oi_1 _6118_ (.Y(_2608_),
    .B1(_2274_),
    .B2(_2607_),
    .A2(net739),
    .A1(net1227));
 sg13g2_o21ai_1 _6119_ (.B1(_2608_),
    .Y(_0753_),
    .A1(net740),
    .A2(net1373));
 sg13g2_a22oi_1 _6120_ (.Y(_2609_),
    .B1(net757),
    .B2(\uart_tx_fifo_inst.fifo[2][6] ),
    .A2(net760),
    .A1(\uart_tx_fifo_inst.fifo[3][6] ));
 sg13g2_inv_1 _6121_ (.Y(_2610_),
    .A(_2609_));
 sg13g2_a21oi_1 _6122_ (.A1(_0891_),
    .A2(net769),
    .Y(_2611_),
    .B1(_1423_));
 sg13g2_o21ai_1 _6123_ (.B1(_2611_),
    .Y(_2612_),
    .A1(net1166),
    .A2(net769));
 sg13g2_a221oi_1 _6124_ (.B2(\uart_tx_fifo_inst.fifo[1][6] ),
    .C1(_2610_),
    .B1(net736),
    .A1(\uart_tx_fifo_inst.fifo[0][6] ),
    .Y(_2613_),
    .A2(net742));
 sg13g2_o21ai_1 _6125_ (.B1(_2612_),
    .Y(_2614_),
    .A1(_2249_),
    .A2(_2613_));
 sg13g2_a22oi_1 _6126_ (.Y(_2615_),
    .B1(net756),
    .B2(net724),
    .A2(net759),
    .A1(net1018));
 sg13g2_a22oi_1 _6127_ (.Y(_2616_),
    .B1(net736),
    .B2(net1102),
    .A2(net742),
    .A1(net1439));
 sg13g2_nand2_1 _6128_ (.Y(_2617_),
    .A(_2615_),
    .B(_2616_));
 sg13g2_a22oi_1 _6129_ (.Y(_2618_),
    .B1(_2274_),
    .B2(_2617_),
    .A2(net739),
    .A1(net1323));
 sg13g2_nand2b_1 _6130_ (.Y(_0754_),
    .B(_2618_),
    .A_N(_2614_));
 sg13g2_a22oi_1 _6131_ (.Y(_2619_),
    .B1(net774),
    .B2(\uart_tx_fifo_inst.fifo[8][0] ),
    .A2(net747),
    .A1(net1174));
 sg13g2_nor2_2 _6132_ (.A(_1423_),
    .B(_2196_),
    .Y(_2620_));
 sg13g2_nor2_1 _6133_ (.A(net1175),
    .B(_2620_),
    .Y(_0755_));
 sg13g2_a22oi_1 _6134_ (.Y(_2621_),
    .B1(net774),
    .B2(\uart_tx_fifo_inst.fifo[8][1] ),
    .A2(net747),
    .A1(net1201));
 sg13g2_nor2_1 _6135_ (.A(_2620_),
    .B(net1202),
    .Y(_0756_));
 sg13g2_a22oi_1 _6136_ (.Y(_2622_),
    .B1(net774),
    .B2(\uart_tx_fifo_inst.fifo[8][2] ),
    .A2(net747),
    .A1(net1107));
 sg13g2_nor2_1 _6137_ (.A(_2620_),
    .B(net1108),
    .Y(_0757_));
 sg13g2_a22oi_1 _6138_ (.Y(_2623_),
    .B1(net774),
    .B2(\uart_tx_fifo_inst.fifo[8][3] ),
    .A2(net747),
    .A1(net1119));
 sg13g2_nor2_1 _6139_ (.A(_2620_),
    .B(net1120),
    .Y(_0758_));
 sg13g2_a22oi_1 _6140_ (.Y(_2624_),
    .B1(net774),
    .B2(\uart_tx_fifo_inst.fifo[8][4] ),
    .A2(net747),
    .A1(net1196));
 sg13g2_nor2_1 _6141_ (.A(_2620_),
    .B(net1197),
    .Y(_0759_));
 sg13g2_a22oi_1 _6142_ (.Y(_2625_),
    .B1(net774),
    .B2(\uart_tx_fifo_inst.fifo[8][5] ),
    .A2(net747),
    .A1(net1198));
 sg13g2_nor2_1 _6143_ (.A(_2620_),
    .B(net1199),
    .Y(_0760_));
 sg13g2_a22oi_1 _6144_ (.Y(_2626_),
    .B1(net773),
    .B2(\uart_tx_fifo_inst.fifo[8][6] ),
    .A2(net746),
    .A1(net1166));
 sg13g2_nor2_1 _6145_ (.A(_2620_),
    .B(net1167),
    .Y(_0761_));
 sg13g2_dfrbp_1 _6146_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net158),
    .D(_0225_),
    .Q_N(_3037_),
    .Q(\uart_tx_fifo_inst.fifo[8][0] ));
 sg13g2_dfrbp_1 _6147_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net258),
    .D(_0226_),
    .Q_N(_3036_),
    .Q(\uart_tx_fifo_inst.fifo[8][1] ));
 sg13g2_dfrbp_1 _6148_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net256),
    .D(_0227_),
    .Q_N(_3035_),
    .Q(\uart_tx_fifo_inst.fifo[8][2] ));
 sg13g2_dfrbp_1 _6149_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net254),
    .D(_0228_),
    .Q_N(_3034_),
    .Q(\uart_tx_fifo_inst.fifo[8][3] ));
 sg13g2_dfrbp_1 _6150_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net252),
    .D(_0229_),
    .Q_N(_3033_),
    .Q(\uart_tx_fifo_inst.fifo[8][4] ));
 sg13g2_dfrbp_1 _6151_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net250),
    .D(_0230_),
    .Q_N(_3032_),
    .Q(\uart_tx_fifo_inst.fifo[8][5] ));
 sg13g2_dfrbp_1 _6152_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net248),
    .D(_0231_),
    .Q_N(_3031_),
    .Q(\uart_tx_fifo_inst.fifo[8][6] ));
 sg13g2_dfrbp_1 _6153_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net246),
    .D(net652),
    .Q_N(_0224_),
    .Q(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[0] ));
 sg13g2_dfrbp_1 _6154_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net245),
    .D(_0233_),
    .Q_N(_3030_),
    .Q(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[1] ));
 sg13g2_dfrbp_1 _6155_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net244),
    .D(net1163),
    .Q_N(_3029_),
    .Q(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[2] ));
 sg13g2_dfrbp_1 _6156_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net243),
    .D(_0235_),
    .Q_N(_0198_),
    .Q(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[3] ));
 sg13g2_dfrbp_1 _6157_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net242),
    .D(_0236_),
    .Q_N(_3028_),
    .Q(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[4] ));
 sg13g2_dfrbp_1 _6158_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net241),
    .D(net1096),
    .Q_N(_0197_),
    .Q(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[5] ));
 sg13g2_dfrbp_1 _6159_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net240),
    .D(net636),
    .Q_N(_0140_),
    .Q(\Led_Cycle_inst.genblk1[15].pwm_unit.pwm_out ));
 sg13g2_dfrbp_1 _6160_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net239),
    .D(net625),
    .Q_N(_0223_),
    .Q(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[0] ));
 sg13g2_dfrbp_1 _6161_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net238),
    .D(_0240_),
    .Q_N(_3027_),
    .Q(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[1] ));
 sg13g2_dfrbp_1 _6162_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net237),
    .D(net1279),
    .Q_N(_3026_),
    .Q(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[2] ));
 sg13g2_dfrbp_1 _6163_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net236),
    .D(_0242_),
    .Q_N(_0196_),
    .Q(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[3] ));
 sg13g2_dfrbp_1 _6164_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net235),
    .D(_0243_),
    .Q_N(_3025_),
    .Q(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[4] ));
 sg13g2_dfrbp_1 _6165_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net234),
    .D(net1078),
    .Q_N(_0195_),
    .Q(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[5] ));
 sg13g2_dfrbp_1 _6166_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net233),
    .D(net648),
    .Q_N(_3024_),
    .Q(\Led_Cycle_inst.genblk1[14].pwm_unit.pwm_out ));
 sg13g2_dfrbp_1 _6167_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net232),
    .D(net662),
    .Q_N(_0222_),
    .Q(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[0] ));
 sg13g2_dfrbp_1 _6168_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net231),
    .D(_0247_),
    .Q_N(_0194_),
    .Q(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[1] ));
 sg13g2_dfrbp_1 _6169_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net230),
    .D(net1276),
    .Q_N(_3023_),
    .Q(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[2] ));
 sg13g2_dfrbp_1 _6170_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net229),
    .D(_0249_),
    .Q_N(_0193_),
    .Q(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[3] ));
 sg13g2_dfrbp_1 _6171_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net228),
    .D(_0250_),
    .Q_N(_3022_),
    .Q(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[4] ));
 sg13g2_dfrbp_1 _6172_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net227),
    .D(net1005),
    .Q_N(_0192_),
    .Q(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[5] ));
 sg13g2_dfrbp_1 _6173_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net226),
    .D(net666),
    .Q_N(_3021_),
    .Q(\Led_Cycle_inst.genblk1[13].pwm_unit.pwm_out ));
 sg13g2_dfrbp_1 _6174_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net225),
    .D(net619),
    .Q_N(_0221_),
    .Q(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[0] ));
 sg13g2_dfrbp_1 _6175_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net224),
    .D(_0254_),
    .Q_N(_3020_),
    .Q(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[1] ));
 sg13g2_dfrbp_1 _6176_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net223),
    .D(net694),
    .Q_N(_3019_),
    .Q(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[2] ));
 sg13g2_dfrbp_1 _6177_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net222),
    .D(_0256_),
    .Q_N(_3018_),
    .Q(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[3] ));
 sg13g2_dfrbp_1 _6178_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net221),
    .D(_0257_),
    .Q_N(_3017_),
    .Q(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[4] ));
 sg13g2_dfrbp_1 _6179_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net220),
    .D(net1043),
    .Q_N(_0191_),
    .Q(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[5] ));
 sg13g2_dfrbp_1 _6180_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net216),
    .D(net684),
    .Q_N(_0142_),
    .Q(\Led_Cycle_inst.genblk1[12].pwm_unit.pwm_out ));
 sg13g2_dfrbp_1 _6181_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net215),
    .D(net686),
    .Q_N(_0220_),
    .Q(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[0] ));
 sg13g2_dfrbp_1 _6182_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net214),
    .D(_0261_),
    .Q_N(_0190_),
    .Q(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[1] ));
 sg13g2_dfrbp_1 _6183_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net213),
    .D(net1397),
    .Q_N(_3016_),
    .Q(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[2] ));
 sg13g2_dfrbp_1 _6184_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net212),
    .D(_0263_),
    .Q_N(_3015_),
    .Q(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[3] ));
 sg13g2_dfrbp_1 _6185_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net211),
    .D(_0264_),
    .Q_N(_3014_),
    .Q(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[4] ));
 sg13g2_dfrbp_1 _6186_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net210),
    .D(net1086),
    .Q_N(_0189_),
    .Q(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[5] ));
 sg13g2_dfrbp_1 _6187_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net209),
    .D(net676),
    .Q_N(_0146_),
    .Q(\Led_Cycle_inst.genblk1[11].pwm_unit.pwm_out ));
 sg13g2_dfrbp_1 _6188_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net208),
    .D(net668),
    .Q_N(_0219_),
    .Q(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[0] ));
 sg13g2_dfrbp_1 _6189_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net207),
    .D(_0268_),
    .Q_N(_0185_),
    .Q(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[1] ));
 sg13g2_dfrbp_1 _6190_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net206),
    .D(net1232),
    .Q_N(_3013_),
    .Q(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[2] ));
 sg13g2_dfrbp_1 _6191_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net205),
    .D(_0270_),
    .Q_N(_0184_),
    .Q(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[3] ));
 sg13g2_dfrbp_1 _6192_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net204),
    .D(_0271_),
    .Q_N(_3012_),
    .Q(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[4] ));
 sg13g2_dfrbp_1 _6193_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net203),
    .D(net1037),
    .Q_N(_0183_),
    .Q(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[5] ));
 sg13g2_dfrbp_1 _6194_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net202),
    .D(net664),
    .Q_N(_3011_),
    .Q(\Led_Cycle_inst.genblk1[10].pwm_unit.pwm_out ));
 sg13g2_dfrbp_1 _6195_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net201),
    .D(net632),
    .Q_N(_0218_),
    .Q(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[0] ));
 sg13g2_dfrbp_1 _6196_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net200),
    .D(_0275_),
    .Q_N(_3010_),
    .Q(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[1] ));
 sg13g2_dfrbp_1 _6197_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net199),
    .D(net1219),
    .Q_N(_3009_),
    .Q(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[2] ));
 sg13g2_dfrbp_1 _6198_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net198),
    .D(_0277_),
    .Q_N(_0179_),
    .Q(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[3] ));
 sg13g2_dfrbp_1 _6199_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net197),
    .D(_0278_),
    .Q_N(_3008_),
    .Q(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[4] ));
 sg13g2_dfrbp_1 _6200_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net196),
    .D(net1101),
    .Q_N(_0178_),
    .Q(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[5] ));
 sg13g2_dfrbp_1 _6201_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net195),
    .D(net656),
    .Q_N(_3007_),
    .Q(\Led_Cycle_inst.genblk1[9].pwm_unit.pwm_out ));
 sg13g2_dfrbp_1 _6202_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net194),
    .D(net615),
    .Q_N(_0217_),
    .Q(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[0] ));
 sg13g2_dfrbp_1 _6203_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net193),
    .D(_0282_),
    .Q_N(_0188_),
    .Q(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[1] ));
 sg13g2_dfrbp_1 _6204_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net192),
    .D(net1345),
    .Q_N(_3006_),
    .Q(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[2] ));
 sg13g2_dfrbp_1 _6205_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net191),
    .D(_0284_),
    .Q_N(_0187_),
    .Q(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[3] ));
 sg13g2_dfrbp_1 _6206_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net190),
    .D(_0285_),
    .Q_N(_3005_),
    .Q(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[4] ));
 sg13g2_dfrbp_1 _6207_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net189),
    .D(net1035),
    .Q_N(_0186_),
    .Q(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[5] ));
 sg13g2_dfrbp_1 _6208_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net188),
    .D(net650),
    .Q_N(_0148_),
    .Q(\Led_Cycle_inst.genblk1[8].pwm_unit.pwm_out ));
 sg13g2_dfrbp_1 _6209_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net187),
    .D(net617),
    .Q_N(_0216_),
    .Q(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[0] ));
 sg13g2_dfrbp_1 _6210_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net186),
    .D(_0289_),
    .Q_N(_3004_),
    .Q(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[1] ));
 sg13g2_dfrbp_1 _6211_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net185),
    .D(net701),
    .Q_N(_3003_),
    .Q(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[2] ));
 sg13g2_dfrbp_1 _6212_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net184),
    .D(_0291_),
    .Q_N(_0175_),
    .Q(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[3] ));
 sg13g2_dfrbp_1 _6213_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net183),
    .D(_0292_),
    .Q_N(_3002_),
    .Q(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[4] ));
 sg13g2_dfrbp_1 _6214_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net182),
    .D(net1021),
    .Q_N(_0174_),
    .Q(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[5] ));
 sg13g2_dfrbp_1 _6215_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net181),
    .D(net630),
    .Q_N(_0161_),
    .Q(\Led_Cycle_inst.genblk1[7].pwm_unit.pwm_out ));
 sg13g2_dfrbp_1 _6216_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net180),
    .D(net670),
    .Q_N(_0215_),
    .Q(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[0] ));
 sg13g2_dfrbp_1 _6217_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net179),
    .D(_0296_),
    .Q_N(_0173_),
    .Q(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[1] ));
 sg13g2_dfrbp_1 _6218_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net169),
    .D(net1236),
    .Q_N(_3001_),
    .Q(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[2] ));
 sg13g2_dfrbp_1 _6219_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net168),
    .D(_0298_),
    .Q_N(_3000_),
    .Q(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[3] ));
 sg13g2_dfrbp_1 _6220_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net167),
    .D(_0299_),
    .Q_N(_2999_),
    .Q(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[4] ));
 sg13g2_dfrbp_1 _6221_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net166),
    .D(net1080),
    .Q_N(_0172_),
    .Q(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[5] ));
 sg13g2_dfrbp_1 _6222_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net165),
    .D(net641),
    .Q_N(_2998_),
    .Q(\Led_Cycle_inst.genblk1[6].pwm_unit.pwm_out ));
 sg13g2_dfrbp_1 _6223_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net164),
    .D(net623),
    .Q_N(_0214_),
    .Q(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[0] ));
 sg13g2_dfrbp_1 _6224_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net163),
    .D(_0303_),
    .Q_N(_2997_),
    .Q(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[1] ));
 sg13g2_dfrbp_1 _6225_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net162),
    .D(net1125),
    .Q_N(_2996_),
    .Q(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[2] ));
 sg13g2_dfrbp_1 _6226_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net161),
    .D(_0305_),
    .Q_N(_2995_),
    .Q(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[3] ));
 sg13g2_dfrbp_1 _6227_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net160),
    .D(_0306_),
    .Q_N(_2994_),
    .Q(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[4] ));
 sg13g2_dfrbp_1 _6228_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net157),
    .D(net1069),
    .Q_N(_0171_),
    .Q(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[5] ));
 sg13g2_dfrbp_1 _6229_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net156),
    .D(net660),
    .Q_N(_2993_),
    .Q(\Led_Cycle_inst.genblk1[5].pwm_unit.pwm_out ));
 sg13g2_dfrbp_1 _6230_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net155),
    .D(net643),
    .Q_N(_0213_),
    .Q(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[0] ));
 sg13g2_dfrbp_1 _6231_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net154),
    .D(net1696),
    .Q_N(_2992_),
    .Q(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[1] ));
 sg13g2_dfrbp_1 _6232_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net153),
    .D(net1186),
    .Q_N(_2991_),
    .Q(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[2] ));
 sg13g2_dfrbp_1 _6233_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net152),
    .D(_0312_),
    .Q_N(_0170_),
    .Q(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[3] ));
 sg13g2_dfrbp_1 _6234_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net151),
    .D(_0313_),
    .Q_N(_2990_),
    .Q(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[4] ));
 sg13g2_dfrbp_1 _6235_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net150),
    .D(net1049),
    .Q_N(_0169_),
    .Q(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[5] ));
 sg13g2_dfrbp_1 _6236_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net149),
    .D(net1487),
    .Q_N(_0163_),
    .Q(\Led_Cycle_inst.genblk1[4].pwm_unit.pwm_out ));
 sg13g2_dfrbp_1 _6237_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net148),
    .D(net639),
    .Q_N(_0212_),
    .Q(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[0] ));
 sg13g2_dfrbp_1 _6238_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net147),
    .D(_0317_),
    .Q_N(_2989_),
    .Q(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[1] ));
 sg13g2_dfrbp_1 _6239_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net146),
    .D(net1299),
    .Q_N(_2988_),
    .Q(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[2] ));
 sg13g2_dfrbp_1 _6240_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net145),
    .D(_0319_),
    .Q_N(_0168_),
    .Q(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[3] ));
 sg13g2_dfrbp_1 _6241_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net144),
    .D(_0320_),
    .Q_N(_2987_),
    .Q(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[4] ));
 sg13g2_dfrbp_1 _6242_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net143),
    .D(net991),
    .Q_N(_0166_),
    .Q(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[5] ));
 sg13g2_dfrbp_1 _6243_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net142),
    .D(net673),
    .Q_N(_0123_),
    .Q(\Led_Cycle_inst.genblk1[3].pwm_unit.pwm_out ));
 sg13g2_dfrbp_1 _6244_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net141),
    .D(net621),
    .Q_N(_0211_),
    .Q(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[0] ));
 sg13g2_dfrbp_1 _6245_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net140),
    .D(_0324_),
    .Q_N(_2986_),
    .Q(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[1] ));
 sg13g2_dfrbp_1 _6246_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net139),
    .D(net1239),
    .Q_N(_2985_),
    .Q(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[2] ));
 sg13g2_dfrbp_1 _6247_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net138),
    .D(_0326_),
    .Q_N(_0202_),
    .Q(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[3] ));
 sg13g2_dfrbp_1 _6248_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net137),
    .D(_0327_),
    .Q_N(_2984_),
    .Q(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[4] ));
 sg13g2_dfrbp_1 _6249_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net136),
    .D(net1071),
    .Q_N(_0201_),
    .Q(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[5] ));
 sg13g2_dfrbp_1 _6250_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net135),
    .D(net628),
    .Q_N(_2983_),
    .Q(\Led_Cycle_inst.genblk1[2].pwm_unit.pwm_out ));
 sg13g2_dfrbp_1 _6251_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net134),
    .D(_0330_),
    .Q_N(_0210_),
    .Q(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[0] ));
 sg13g2_dfrbp_1 _6252_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net133),
    .D(net613),
    .Q_N(_2982_),
    .Q(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[1] ));
 sg13g2_dfrbp_1 _6253_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net132),
    .D(net611),
    .Q_N(_2981_),
    .Q(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[2] ));
 sg13g2_dfrbp_1 _6254_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net131),
    .D(_0333_),
    .Q_N(_0200_),
    .Q(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[3] ));
 sg13g2_dfrbp_1 _6255_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net130),
    .D(_0334_),
    .Q_N(_2980_),
    .Q(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[4] ));
 sg13g2_dfrbp_1 _6256_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net129),
    .D(net1025),
    .Q_N(_0199_),
    .Q(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[5] ));
 sg13g2_dfrbp_1 _6257_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net128),
    .D(net654),
    .Q_N(_2979_),
    .Q(\Led_Cycle_inst.genblk1[1].pwm_unit.pwm_out ));
 sg13g2_dfrbp_1 _6258_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net127),
    .D(_0337_),
    .Q_N(_0209_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[0] ));
 sg13g2_dfrbp_1 _6259_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net126),
    .D(_0338_),
    .Q_N(_2978_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[1] ));
 sg13g2_dfrbp_1 _6260_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net125),
    .D(net1311),
    .Q_N(_2977_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[2] ));
 sg13g2_dfrbp_1 _6261_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net124),
    .D(_0340_),
    .Q_N(_2976_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[3] ));
 sg13g2_dfrbp_1 _6262_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net123),
    .D(_0341_),
    .Q_N(_2975_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[4] ));
 sg13g2_dfrbp_1 _6263_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net122),
    .D(_0342_),
    .Q_N(_0182_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[5] ));
 sg13g2_dfrbp_1 _6264_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net121),
    .D(_0343_),
    .Q_N(_0110_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[6] ));
 sg13g2_dfrbp_1 _6265_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net120),
    .D(_0344_),
    .Q_N(_2974_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[7] ));
 sg13g2_dfrbp_1 _6266_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net119),
    .D(_0345_),
    .Q_N(_0112_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[8] ));
 sg13g2_dfrbp_1 _6267_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net118),
    .D(_0346_),
    .Q_N(_0113_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[9] ));
 sg13g2_dfrbp_1 _6268_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net117),
    .D(_0347_),
    .Q_N(_2973_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[10] ));
 sg13g2_dfrbp_1 _6269_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net116),
    .D(_0348_),
    .Q_N(_0114_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[11] ));
 sg13g2_dfrbp_1 _6270_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net115),
    .D(net1402),
    .Q_N(_2972_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[12] ));
 sg13g2_dfrbp_1 _6271_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net114),
    .D(_0350_),
    .Q_N(_2971_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[13] ));
 sg13g2_dfrbp_1 _6272_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net113),
    .D(_0351_),
    .Q_N(_0115_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[14] ));
 sg13g2_dfrbp_1 _6273_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net112),
    .D(_0352_),
    .Q_N(_0181_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[15] ));
 sg13g2_dfrbp_1 _6274_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net111),
    .D(_0353_),
    .Q_N(_2970_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[16] ));
 sg13g2_dfrbp_1 _6275_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net110),
    .D(_0354_),
    .Q_N(_2969_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[17] ));
 sg13g2_dfrbp_1 _6276_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net109),
    .D(_0355_),
    .Q_N(_0180_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[18] ));
 sg13g2_dfrbp_1 _6277_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net108),
    .D(_0356_),
    .Q_N(_2968_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[19] ));
 sg13g2_dfrbp_1 _6278_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net107),
    .D(_0357_),
    .Q_N(_2967_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[20] ));
 sg13g2_dfrbp_1 _6279_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net106),
    .D(_0358_),
    .Q_N(_2966_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[21] ));
 sg13g2_dfrbp_1 _6280_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net105),
    .D(_0359_),
    .Q_N(_2965_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[22] ));
 sg13g2_dfrbp_1 _6281_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net104),
    .D(_0360_),
    .Q_N(_2964_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[23] ));
 sg13g2_dfrbp_1 _6282_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net103),
    .D(_0361_),
    .Q_N(_2963_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[24] ));
 sg13g2_dfrbp_1 _6283_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net102),
    .D(_0362_),
    .Q_N(_2962_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[25] ));
 sg13g2_dfrbp_1 _6284_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net101),
    .D(net1435),
    .Q_N(_2961_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[26] ));
 sg13g2_dfrbp_1 _6285_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net100),
    .D(_0364_),
    .Q_N(_2960_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[27] ));
 sg13g2_dfrbp_1 _6286_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net99),
    .D(_0365_),
    .Q_N(_2959_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[28] ));
 sg13g2_dfrbp_1 _6287_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net98),
    .D(_0366_),
    .Q_N(_2958_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[29] ));
 sg13g2_dfrbp_1 _6288_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net97),
    .D(net1210),
    .Q_N(_2957_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[30] ));
 sg13g2_dfrbp_1 _6289_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net96),
    .D(_0368_),
    .Q_N(_2956_),
    .Q(\Led_Cycle_inst.clk_reducer.counter[31] ));
 sg13g2_dfrbp_1 _6290_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net95),
    .D(net679),
    .Q_N(_0125_),
    .Q(\Led_Cycle_inst.genblk1[0].pwm_unit.pwm_out ));
 sg13g2_dfrbp_1 _6291_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net94),
    .D(_0370_),
    .Q_N(_2955_),
    .Q(\Led_Cycle_inst.clk_reduced ));
 sg13g2_dfrbp_1 _6292_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net93),
    .D(net1677),
    .Q_N(_2954_),
    .Q(_0064_));
 sg13g2_dfrbp_1 _6293_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net159),
    .D(net1709),
    .Q_N(_3038_),
    .Q(_0066_));
 sg13g2_dfrbp_1 _6294_ (.CLK(\Led_Cycle_inst.clk_reduced ),
    .RESET_B(net920),
    .D(_2628_),
    .Q_N(_2628_),
    .Q(\Led_Cycle_inst.csr.read_ptr[0] ));
 sg13g2_dfrbp_1 _6295_ (.CLK(\Led_Cycle_inst.clk_reduced ),
    .RESET_B(net920),
    .D(_0203_),
    .Q_N(_3039_),
    .Q(\Led_Cycle_inst.csr.read_ptr[1] ));
 sg13g2_dfrbp_1 _6296_ (.CLK(\Led_Cycle_inst.clk_reduced ),
    .RESET_B(net944),
    .D(_0204_),
    .Q_N(_0097_),
    .Q(\Led_Cycle_inst.csr.read_ptr[2] ));
 sg13g2_dfrbp_1 _6297_ (.CLK(\Led_Cycle_inst.clk_reduced ),
    .RESET_B(net944),
    .D(_0205_),
    .Q_N(_0167_),
    .Q(\Led_Cycle_inst.csr.read_ptr[3] ));
 sg13g2_dfrbp_1 _6298_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net92),
    .D(_0373_),
    .Q_N(_2953_),
    .Q(_0095_));
 sg13g2_dfrbp_1 _6299_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net91),
    .D(_0374_),
    .Q_N(_2952_),
    .Q(_0083_));
 sg13g2_dfrbp_1 _6300_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net90),
    .D(_0375_),
    .Q_N(_2951_),
    .Q(_0089_));
 sg13g2_dfrbp_1 _6301_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net89),
    .D(_0376_),
    .Q_N(_2950_),
    .Q(_0071_));
 sg13g2_dfrbp_1 _6302_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net88),
    .D(_0377_),
    .Q_N(_2949_),
    .Q(_0065_));
 sg13g2_dfrbp_1 _6303_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net87),
    .D(_0378_),
    .Q_N(_2948_),
    .Q(_0059_));
 sg13g2_dfrbp_1 _6304_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net86),
    .D(_0379_),
    .Q_N(_2947_),
    .Q(_0077_));
 sg13g2_dfrbp_1 _6305_ (.CLK(\SegmentDisplay.seg_driver.clk_reduced ),
    .RESET_B(net85),
    .D(_0380_),
    .Q_N(\SegmentDisplay.an[3] ),
    .Q(\SegmentDisplay.out_sel[3] ));
 sg13g2_dfrbp_1 _6306_ (.CLK(\SegmentDisplay.seg_driver.clk_reduced ),
    .RESET_B(net84),
    .D(_0381_),
    .Q_N(\SegmentDisplay.an[2] ),
    .Q(\SegmentDisplay.out_sel[2] ));
 sg13g2_dfrbp_1 _6307_ (.CLK(\SegmentDisplay.seg_driver.clk_reduced ),
    .RESET_B(net170),
    .D(_0382_),
    .Q_N(\SegmentDisplay.an[1] ),
    .Q(\SegmentDisplay.out_sel[1] ));
 sg13g2_dfrbp_1 _6308_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net171),
    .D(_0014_),
    .Q_N(_3040_),
    .Q(\SegmentDisplay.digit2[0] ));
 sg13g2_dfrbp_1 _6309_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net172),
    .D(_0015_),
    .Q_N(_3041_),
    .Q(\SegmentDisplay.digit2[1] ));
 sg13g2_dfrbp_1 _6310_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net173),
    .D(_0016_),
    .Q_N(_3042_),
    .Q(\SegmentDisplay.digit2[2] ));
 sg13g2_dfrbp_1 _6311_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net174),
    .D(_0017_),
    .Q_N(_3043_),
    .Q(\SegmentDisplay.digit2[3] ));
 sg13g2_dfrbp_1 _6312_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net175),
    .D(net1669),
    .Q_N(_3044_),
    .Q(\SegmentDisplay.digit2[4] ));
 sg13g2_dfrbp_1 _6313_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net176),
    .D(_0019_),
    .Q_N(_3045_),
    .Q(\SegmentDisplay.digit2[5] ));
 sg13g2_dfrbp_1 _6314_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net177),
    .D(_0020_),
    .Q_N(_3046_),
    .Q(\SegmentDisplay.digit2[6] ));
 sg13g2_dfrbp_1 _6315_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net178),
    .D(_0049_),
    .Q_N(_3047_),
    .Q(\uart_inst.uart_rx_inst.state[0] ));
 sg13g2_dfrbp_1 _6316_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net217),
    .D(_0050_),
    .Q_N(_3048_),
    .Q(\uart_inst.uart_rx_inst.state[1] ));
 sg13g2_dfrbp_1 _6317_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net83),
    .D(_0051_),
    .Q_N(_0106_),
    .Q(\uart_inst.uart_rx_inst.state[2] ));
 sg13g2_dfrbp_1 _6318_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net82),
    .D(net996),
    .Q_N(_2946_),
    .Q(\rx_data[0] ));
 sg13g2_dfrbp_1 _6319_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net80),
    .D(net980),
    .Q_N(_2945_),
    .Q(\rx_data[1] ));
 sg13g2_dfrbp_1 _6320_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net78),
    .D(net1023),
    .Q_N(_2944_),
    .Q(\rx_data[2] ));
 sg13g2_dfrbp_1 _6321_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net76),
    .D(_0386_),
    .Q_N(_2943_),
    .Q(\rx_data[3] ));
 sg13g2_dfrbp_1 _6322_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net74),
    .D(_0387_),
    .Q_N(_2942_),
    .Q(\rx_data[4] ));
 sg13g2_dfrbp_1 _6323_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net72),
    .D(_0388_),
    .Q_N(_2941_),
    .Q(\rx_data[5] ));
 sg13g2_dfrbp_1 _6324_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net70),
    .D(_0389_),
    .Q_N(_2940_),
    .Q(\rx_data[6] ));
 sg13g2_dfrbp_1 _6325_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net68),
    .D(_0390_),
    .Q_N(_2939_),
    .Q(\rx_data[7] ));
 sg13g2_dfrbp_1 _6326_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net66),
    .D(_0391_),
    .Q_N(_2938_),
    .Q(rx_valid));
 sg13g2_dfrbp_1 _6327_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net64),
    .D(net710),
    .Q_N(_2937_),
    .Q(\uart_inst.uart_rx_inst.DATA_TEMP_REG[0] ));
 sg13g2_dfrbp_1 _6328_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net62),
    .D(net1180),
    .Q_N(_2936_),
    .Q(\uart_inst.uart_rx_inst.DATA_TEMP_REG[1] ));
 sg13g2_dfrbp_1 _6329_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net60),
    .D(_0394_),
    .Q_N(_2935_),
    .Q(\uart_inst.uart_rx_inst.DATA_TEMP_REG[2] ));
 sg13g2_dfrbp_1 _6330_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net58),
    .D(_0395_),
    .Q_N(_2934_),
    .Q(\uart_inst.uart_rx_inst.DATA_TEMP_REG[3] ));
 sg13g2_dfrbp_1 _6331_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net56),
    .D(_0396_),
    .Q_N(_2933_),
    .Q(\uart_inst.uart_rx_inst.DATA_TEMP_REG[4] ));
 sg13g2_dfrbp_1 _6332_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net54),
    .D(_0397_),
    .Q_N(_2932_),
    .Q(\uart_inst.uart_rx_inst.DATA_TEMP_REG[5] ));
 sg13g2_dfrbp_1 _6333_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net52),
    .D(net1073),
    .Q_N(_2931_),
    .Q(\uart_inst.uart_rx_inst.DATA_TEMP_REG[6] ));
 sg13g2_dfrbp_1 _6334_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net50),
    .D(_0399_),
    .Q_N(_2930_),
    .Q(\uart_inst.uart_rx_inst.DATA_TEMP_REG[7] ));
 sg13g2_dfrbp_1 _6335_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net48),
    .D(_0400_),
    .Q_N(_2929_),
    .Q(\uart_inst.uart_rx_inst.DATA_CNT[0] ));
 sg13g2_dfrbp_1 _6336_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net46),
    .D(_0401_),
    .Q_N(_2928_),
    .Q(\uart_inst.uart_rx_inst.DATA_CNT[1] ));
 sg13g2_dfrbp_1 _6337_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net44),
    .D(_0402_),
    .Q_N(_2927_),
    .Q(\uart_inst.uart_rx_inst.DATA_CNT[2] ));
 sg13g2_dfrbp_1 _6338_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net42),
    .D(net681),
    .Q_N(_2926_),
    .Q(\uart_inst.uart_rx_inst.DATA_CNT[3] ));
 sg13g2_dfrbp_1 _6339_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net40),
    .D(net1572),
    .Q_N(_2925_),
    .Q(\uart_inst.uart_rx_inst.CLK_CNT[0] ));
 sg13g2_dfrbp_1 _6340_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net38),
    .D(net1333),
    .Q_N(_2924_),
    .Q(\uart_inst.uart_rx_inst.CLK_CNT[1] ));
 sg13g2_dfrbp_1 _6341_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net36),
    .D(net1502),
    .Q_N(_0126_),
    .Q(\uart_inst.uart_rx_inst.CLK_CNT[2] ));
 sg13g2_dfrbp_1 _6342_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net34),
    .D(net1621),
    .Q_N(_2923_),
    .Q(\uart_inst.uart_rx_inst.CLK_CNT[3] ));
 sg13g2_dfrbp_1 _6343_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net32),
    .D(_0408_),
    .Q_N(_2922_),
    .Q(\uart_inst.uart_rx_inst.CLK_CNT[4] ));
 sg13g2_dfrbp_1 _6344_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net30),
    .D(_0409_),
    .Q_N(_2921_),
    .Q(\uart_inst.uart_rx_inst.CLK_CNT[5] ));
 sg13g2_dfrbp_1 _6345_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net28),
    .D(_0410_),
    .Q_N(_2920_),
    .Q(\uart_inst.uart_rx_inst.CLK_CNT[6] ));
 sg13g2_dfrbp_1 _6346_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net26),
    .D(_0411_),
    .Q_N(_2919_),
    .Q(\uart_inst.uart_rx_inst.CLK_CNT[7] ));
 sg13g2_dfrbp_1 _6347_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net24),
    .D(_0412_),
    .Q_N(_2918_),
    .Q(\uart_inst.uart_rx_inst.CLK_CNT[8] ));
 sg13g2_dfrbp_1 _6348_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net22),
    .D(net1432),
    .Q_N(_2917_),
    .Q(\uart_inst.uart_rx_inst.CLK_CNT[9] ));
 sg13g2_dfrbp_1 _6349_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net20),
    .D(_0414_),
    .Q_N(_0208_),
    .Q(\uart_inst.uart_rx_inst.SAMPLING_COUNT[0] ));
 sg13g2_dfrbp_1 _6350_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net18),
    .D(net1256),
    .Q_N(_2916_),
    .Q(\uart_inst.uart_rx_inst.SAMPLING_COUNT[1] ));
 sg13g2_dfrbp_1 _6351_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net16),
    .D(_0416_),
    .Q_N(_2915_),
    .Q(\uart_inst.uart_rx_inst.SIGNAL_Q[0] ));
 sg13g2_dfrbp_1 _6352_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net14),
    .D(net1384),
    .Q_N(_2914_),
    .Q(\uart_inst.uart_rx_inst.SIGNAL_Q[1] ));
 sg13g2_dfrbp_1 _6353_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net12),
    .D(net1495),
    .Q_N(_0152_),
    .Q(\uart_inst.uart_rx_inst.SIGNAL_Q[2] ));
 sg13g2_dfrbp_1 _6354_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net595),
    .D(net1563),
    .Q_N(_2913_),
    .Q(\uart_inst.uart_rx_inst.SIGNAL_Q[3] ));
 sg13g2_dfrbp_1 _6355_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net218),
    .D(_0420_),
    .Q_N(_3049_),
    .Q(\uart_inst.uart_rx_inst.SIGNAL_Q[4] ));
 sg13g2_dfrbp_1 _6356_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net219),
    .D(_0046_),
    .Q_N(_3050_),
    .Q(_0091_));
 sg13g2_dfrbp_1 _6357_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net319),
    .D(_0047_),
    .Q_N(_3051_),
    .Q(_0092_));
 sg13g2_dfrbp_1 _6358_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net593),
    .D(net1768),
    .Q_N(_2912_),
    .Q(_0093_));
 sg13g2_dfrbp_1 _6359_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net591),
    .D(net1691),
    .Q_N(_2911_),
    .Q(_0070_));
 sg13g2_dfrbp_1 _6360_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net590),
    .D(_0422_),
    .Q_N(_2910_),
    .Q(_0072_));
 sg13g2_dfrbp_1 _6361_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net589),
    .D(_0423_),
    .Q_N(_2909_),
    .Q(\uart_inst.uart_tx_inst.DATA_CNT[0] ));
 sg13g2_dfrbp_1 _6362_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net587),
    .D(_0424_),
    .Q_N(_2908_),
    .Q(\uart_inst.uart_tx_inst.DATA_CNT[1] ));
 sg13g2_dfrbp_1 _6363_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net585),
    .D(_0425_),
    .Q_N(_0108_),
    .Q(\uart_inst.uart_tx_inst.DATA_CNT[2] ));
 sg13g2_dfrbp_1 _6364_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net583),
    .D(net1532),
    .Q_N(_0134_),
    .Q(\uart_inst.uart_tx_inst.CLK_CNT[0] ));
 sg13g2_dfrbp_1 _6365_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net581),
    .D(net1362),
    .Q_N(_2907_),
    .Q(\uart_inst.uart_tx_inst.CLK_CNT[1] ));
 sg13g2_dfrbp_1 _6366_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net579),
    .D(_0428_),
    .Q_N(_2906_),
    .Q(\uart_inst.uart_tx_inst.CLK_CNT[2] ));
 sg13g2_dfrbp_1 _6367_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net577),
    .D(_0429_),
    .Q_N(_2905_),
    .Q(\uart_inst.uart_tx_inst.CLK_CNT[3] ));
 sg13g2_dfrbp_1 _6368_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net575),
    .D(_0430_),
    .Q_N(_2904_),
    .Q(\uart_inst.uart_tx_inst.CLK_CNT[4] ));
 sg13g2_dfrbp_1 _6369_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net573),
    .D(net1566),
    .Q_N(_2903_),
    .Q(\uart_inst.uart_tx_inst.CLK_CNT[5] ));
 sg13g2_dfrbp_1 _6370_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net571),
    .D(_0432_),
    .Q_N(_2902_),
    .Q(\uart_inst.uart_tx_inst.CLK_CNT[6] ));
 sg13g2_dfrbp_1 _6371_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net569),
    .D(net1106),
    .Q_N(_2901_),
    .Q(\uart_inst.uart_tx_inst.CLK_CNT[7] ));
 sg13g2_dfrbp_1 _6372_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net567),
    .D(net1446),
    .Q_N(_2900_),
    .Q(\uart_inst.uart_tx_inst.CLK_CNT[8] ));
 sg13g2_dfrbp_1 _6373_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net565),
    .D(_0435_),
    .Q_N(_2899_),
    .Q(\uart_inst.uart_tx_inst.CLK_CNT[9] ));
 sg13g2_dfrbp_1 _6374_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net563),
    .D(net1378),
    .Q_N(_2898_),
    .Q(tx_signal));
 sg13g2_dfrbp_1 _6375_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net561),
    .D(_0437_),
    .Q_N(_0107_),
    .Q(\output_value_inst.tx_ready ));
 sg13g2_dfrbp_1 _6376_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net559),
    .D(net1391),
    .Q_N(_2897_),
    .Q(\input_value_check_inst.character_buff[9][0] ));
 sg13g2_dfrbp_1 _6377_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net557),
    .D(net1152),
    .Q_N(_2896_),
    .Q(\input_value_check_inst.character_buff[9][1] ));
 sg13g2_dfrbp_1 _6378_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net555),
    .D(_0440_),
    .Q_N(_2895_),
    .Q(\input_value_check_inst.character_buff[9][2] ));
 sg13g2_dfrbp_1 _6379_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net553),
    .D(net1154),
    .Q_N(_2894_),
    .Q(\input_value_check_inst.character_buff[9][3] ));
 sg13g2_dfrbp_1 _6380_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net551),
    .D(net1342),
    .Q_N(_2893_),
    .Q(\input_value_check_inst.character_buff[9][4] ));
 sg13g2_dfrbp_1 _6381_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net549),
    .D(net1247),
    .Q_N(_2892_),
    .Q(\input_value_check_inst.character_buff[9][5] ));
 sg13g2_dfrbp_1 _6382_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net547),
    .D(net1045),
    .Q_N(_2891_),
    .Q(\input_value_check_inst.character_buff[9][6] ));
 sg13g2_dfrbp_1 _6383_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net545),
    .D(net1253),
    .Q_N(_2890_),
    .Q(\input_value_check_inst.character_buff[9][7] ));
 sg13g2_dfrbp_1 _6384_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net543),
    .D(net1135),
    .Q_N(_2889_),
    .Q(\input_value_check_inst.character_buff[8][0] ));
 sg13g2_dfrbp_1 _6385_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net541),
    .D(net1216),
    .Q_N(_2888_),
    .Q(\input_value_check_inst.character_buff[8][1] ));
 sg13g2_dfrbp_1 _6386_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net539),
    .D(_0448_),
    .Q_N(_2887_),
    .Q(\input_value_check_inst.character_buff[8][2] ));
 sg13g2_dfrbp_1 _6387_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net537),
    .D(_0449_),
    .Q_N(_2886_),
    .Q(\input_value_check_inst.character_buff[8][3] ));
 sg13g2_dfrbp_1 _6388_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net535),
    .D(_0450_),
    .Q_N(_2885_),
    .Q(\input_value_check_inst.character_buff[8][4] ));
 sg13g2_dfrbp_1 _6389_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net533),
    .D(_0451_),
    .Q_N(_2884_),
    .Q(\input_value_check_inst.character_buff[8][5] ));
 sg13g2_dfrbp_1 _6390_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net531),
    .D(net1367),
    .Q_N(_2883_),
    .Q(\input_value_check_inst.character_buff[8][6] ));
 sg13g2_dfrbp_1 _6391_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net529),
    .D(_0453_),
    .Q_N(_2882_),
    .Q(\input_value_check_inst.character_buff[8][7] ));
 sg13g2_dfrbp_1 _6392_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net527),
    .D(_0454_),
    .Q_N(_2881_),
    .Q(\input_value_check_inst.character_buff[7][0] ));
 sg13g2_dfrbp_1 _6393_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net525),
    .D(_0455_),
    .Q_N(_2880_),
    .Q(\input_value_check_inst.character_buff[7][1] ));
 sg13g2_dfrbp_1 _6394_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net523),
    .D(_0456_),
    .Q_N(_2879_),
    .Q(\input_value_check_inst.character_buff[7][2] ));
 sg13g2_dfrbp_1 _6395_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net521),
    .D(_0457_),
    .Q_N(_2878_),
    .Q(\input_value_check_inst.character_buff[7][3] ));
 sg13g2_dfrbp_1 _6396_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net519),
    .D(net1169),
    .Q_N(_2877_),
    .Q(\input_value_check_inst.character_buff[7][4] ));
 sg13g2_dfrbp_1 _6397_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net517),
    .D(_0459_),
    .Q_N(_2876_),
    .Q(\input_value_check_inst.character_buff[7][5] ));
 sg13g2_dfrbp_1 _6398_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net515),
    .D(net1212),
    .Q_N(_2875_),
    .Q(\input_value_check_inst.character_buff[7][6] ));
 sg13g2_dfrbp_1 _6399_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net513),
    .D(_0461_),
    .Q_N(_2874_),
    .Q(\input_value_check_inst.character_buff[7][7] ));
 sg13g2_dfrbp_1 _6400_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net511),
    .D(_0462_),
    .Q_N(_2873_),
    .Q(\input_value_check_inst.character_buff[6][0] ));
 sg13g2_dfrbp_1 _6401_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net509),
    .D(_0463_),
    .Q_N(_2872_),
    .Q(\input_value_check_inst.character_buff[6][1] ));
 sg13g2_dfrbp_1 _6402_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net507),
    .D(net1131),
    .Q_N(_2871_),
    .Q(\input_value_check_inst.character_buff[6][2] ));
 sg13g2_dfrbp_1 _6403_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net505),
    .D(net1306),
    .Q_N(_2870_),
    .Q(\input_value_check_inst.character_buff[6][3] ));
 sg13g2_dfrbp_1 _6404_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net503),
    .D(_0466_),
    .Q_N(_2869_),
    .Q(\input_value_check_inst.character_buff[6][4] ));
 sg13g2_dfrbp_1 _6405_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net501),
    .D(_0467_),
    .Q_N(_2868_),
    .Q(\input_value_check_inst.character_buff[6][5] ));
 sg13g2_dfrbp_1 _6406_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net499),
    .D(_0468_),
    .Q_N(_2867_),
    .Q(\input_value_check_inst.character_buff[6][6] ));
 sg13g2_dfrbp_1 _6407_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net497),
    .D(_0469_),
    .Q_N(_2866_),
    .Q(\input_value_check_inst.character_buff[6][7] ));
 sg13g2_dfrbp_1 _6408_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net495),
    .D(net1269),
    .Q_N(_2865_),
    .Q(\input_value_check_inst.character_buff[5][0] ));
 sg13g2_dfrbp_1 _6409_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net493),
    .D(net1143),
    .Q_N(_2864_),
    .Q(\input_value_check_inst.character_buff[5][1] ));
 sg13g2_dfrbp_1 _6410_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net491),
    .D(net1250),
    .Q_N(_2863_),
    .Q(\input_value_check_inst.character_buff[5][2] ));
 sg13g2_dfrbp_1 _6411_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net489),
    .D(_0473_),
    .Q_N(_2862_),
    .Q(\input_value_check_inst.character_buff[5][3] ));
 sg13g2_dfrbp_1 _6412_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net487),
    .D(_0474_),
    .Q_N(_2861_),
    .Q(\input_value_check_inst.character_buff[5][4] ));
 sg13g2_dfrbp_1 _6413_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net485),
    .D(net1207),
    .Q_N(_2860_),
    .Q(\input_value_check_inst.character_buff[5][5] ));
 sg13g2_dfrbp_1 _6414_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net483),
    .D(net1349),
    .Q_N(_2859_),
    .Q(\input_value_check_inst.character_buff[5][6] ));
 sg13g2_dfrbp_1 _6415_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net481),
    .D(net1172),
    .Q_N(_2858_),
    .Q(\input_value_check_inst.character_buff[5][7] ));
 sg13g2_dfrbp_1 _6416_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net479),
    .D(net1539),
    .Q_N(_2857_),
    .Q(\input_value_check_inst.character_buff[4][0] ));
 sg13g2_dfrbp_1 _6417_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net477),
    .D(_0479_),
    .Q_N(_2856_),
    .Q(\input_value_check_inst.character_buff[4][1] ));
 sg13g2_dfrbp_1 _6418_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net475),
    .D(_0480_),
    .Q_N(_2855_),
    .Q(\input_value_check_inst.character_buff[4][2] ));
 sg13g2_dfrbp_1 _6419_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net473),
    .D(net1285),
    .Q_N(_2854_),
    .Q(\input_value_check_inst.character_buff[4][3] ));
 sg13g2_dfrbp_1 _6420_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net471),
    .D(_0482_),
    .Q_N(_2853_),
    .Q(\input_value_check_inst.character_buff[4][4] ));
 sg13g2_dfrbp_1 _6421_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net469),
    .D(_0483_),
    .Q_N(_2852_),
    .Q(\input_value_check_inst.character_buff[4][5] ));
 sg13g2_dfrbp_1 _6422_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net467),
    .D(net1326),
    .Q_N(_2851_),
    .Q(\input_value_check_inst.character_buff[4][6] ));
 sg13g2_dfrbp_1 _6423_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net465),
    .D(net1290),
    .Q_N(_2850_),
    .Q(\input_value_check_inst.character_buff[4][7] ));
 sg13g2_dfrbp_1 _6424_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net463),
    .D(_0486_),
    .Q_N(_0135_),
    .Q(\input_value_check_inst.character_buff[3][0] ));
 sg13g2_dfrbp_1 _6425_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net461),
    .D(_0487_),
    .Q_N(_0136_),
    .Q(\input_value_check_inst.character_buff[3][1] ));
 sg13g2_dfrbp_1 _6426_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net459),
    .D(_0488_),
    .Q_N(_0137_),
    .Q(\input_value_check_inst.character_buff[3][2] ));
 sg13g2_dfrbp_1 _6427_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net457),
    .D(_0489_),
    .Q_N(_0138_),
    .Q(\input_value_check_inst.character_buff[3][3] ));
 sg13g2_dfrbp_1 _6428_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net455),
    .D(_0490_),
    .Q_N(_2849_),
    .Q(\input_value_check_inst.character_buff[3][4] ));
 sg13g2_dfrbp_1 _6429_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net453),
    .D(_0491_),
    .Q_N(_2848_),
    .Q(\input_value_check_inst.character_buff[3][5] ));
 sg13g2_dfrbp_1 _6430_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net451),
    .D(_0492_),
    .Q_N(_2847_),
    .Q(\input_value_check_inst.character_buff[3][6] ));
 sg13g2_dfrbp_1 _6431_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net449),
    .D(_0493_),
    .Q_N(_2846_),
    .Q(\input_value_check_inst.character_buff[3][7] ));
 sg13g2_dfrbp_1 _6432_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net447),
    .D(_0494_),
    .Q_N(_0131_),
    .Q(\input_value_check_inst.character_buff[2][0] ));
 sg13g2_dfrbp_1 _6433_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net445),
    .D(_0495_),
    .Q_N(_0128_),
    .Q(\input_value_check_inst.character_buff[2][1] ));
 sg13g2_dfrbp_1 _6434_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net443),
    .D(_0496_),
    .Q_N(_0132_),
    .Q(\input_value_check_inst.character_buff[2][2] ));
 sg13g2_dfrbp_1 _6435_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net441),
    .D(_0497_),
    .Q_N(_0133_),
    .Q(\input_value_check_inst.character_buff[2][3] ));
 sg13g2_dfrbp_1 _6436_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net439),
    .D(net1506),
    .Q_N(_2845_),
    .Q(\input_value_check_inst.character_buff[2][4] ));
 sg13g2_dfrbp_1 _6437_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net437),
    .D(_0499_),
    .Q_N(_2844_),
    .Q(\input_value_check_inst.character_buff[2][5] ));
 sg13g2_dfrbp_1 _6438_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net435),
    .D(_0500_),
    .Q_N(_2843_),
    .Q(\input_value_check_inst.character_buff[2][6] ));
 sg13g2_dfrbp_1 _6439_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net433),
    .D(_0501_),
    .Q_N(_0129_),
    .Q(\input_value_check_inst.character_buff[2][7] ));
 sg13g2_dfrbp_1 _6440_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net431),
    .D(_0502_),
    .Q_N(_0117_),
    .Q(\input_value_check_inst.character_buff[1][0] ));
 sg13g2_dfrbp_1 _6441_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net429),
    .D(_0503_),
    .Q_N(_0118_),
    .Q(\input_value_check_inst.character_buff[1][1] ));
 sg13g2_dfrbp_1 _6442_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net427),
    .D(_0504_),
    .Q_N(_0116_),
    .Q(\input_value_check_inst.character_buff[1][2] ));
 sg13g2_dfrbp_1 _6443_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net425),
    .D(net1448),
    .Q_N(_0120_),
    .Q(\input_value_check_inst.character_buff[1][3] ));
 sg13g2_dfrbp_1 _6444_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net423),
    .D(_0506_),
    .Q_N(_2842_),
    .Q(\input_value_check_inst.character_buff[1][4] ));
 sg13g2_dfrbp_1 _6445_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net421),
    .D(net1150),
    .Q_N(_2841_),
    .Q(\input_value_check_inst.character_buff[1][5] ));
 sg13g2_dfrbp_1 _6446_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net419),
    .D(_0508_),
    .Q_N(_2840_),
    .Q(\input_value_check_inst.character_buff[1][6] ));
 sg13g2_dfrbp_1 _6447_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net417),
    .D(net1369),
    .Q_N(_2839_),
    .Q(\input_value_check_inst.character_buff[1][7] ));
 sg13g2_dfrbp_1 _6448_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net415),
    .D(_0510_),
    .Q_N(_0156_),
    .Q(\input_value_check_inst.character_buff[0][0] ));
 sg13g2_dfrbp_1 _6449_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net413),
    .D(_0511_),
    .Q_N(_0154_),
    .Q(\input_value_check_inst.character_buff[0][1] ));
 sg13g2_dfrbp_1 _6450_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net411),
    .D(_0512_),
    .Q_N(_0157_),
    .Q(\input_value_check_inst.character_buff[0][2] ));
 sg13g2_dfrbp_1 _6451_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net409),
    .D(net1003),
    .Q_N(_0158_),
    .Q(\input_value_check_inst.character_buff[0][3] ));
 sg13g2_dfrbp_1 _6452_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net407),
    .D(net1084),
    .Q_N(_2838_),
    .Q(\input_value_check_inst.character_buff[0][4] ));
 sg13g2_dfrbp_1 _6453_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net405),
    .D(net1067),
    .Q_N(_2837_),
    .Q(\input_value_check_inst.character_buff[0][5] ));
 sg13g2_dfrbp_1 _6454_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net403),
    .D(_0516_),
    .Q_N(_2836_),
    .Q(\input_value_check_inst.character_buff[0][6] ));
 sg13g2_dfrbp_1 _6455_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net401),
    .D(net1030),
    .Q_N(_2835_),
    .Q(\input_value_check_inst.character_buff[0][7] ));
 sg13g2_dfrbp_1 _6456_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net399),
    .D(_0518_),
    .Q_N(_2834_),
    .Q(_0082_));
 sg13g2_dfrbp_1 _6457_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net320),
    .D(_0519_),
    .Q_N(_3052_),
    .Q(_0084_));
 sg13g2_dfrbp_1 _6458_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net321),
    .D(_0040_),
    .Q_N(_3053_),
    .Q(_0079_));
 sg13g2_dfrbp_1 _6459_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net322),
    .D(_0041_),
    .Q_N(_3054_),
    .Q(_0080_));
 sg13g2_dfrbp_1 _6460_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net323),
    .D(net1739),
    .Q_N(_3055_),
    .Q(_0081_));
 sg13g2_dfrbp_1 _6461_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net324),
    .D(_0021_),
    .Q_N(_3056_),
    .Q(\SegmentDisplay.digit3[0] ));
 sg13g2_dfrbp_1 _6462_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net325),
    .D(_0022_),
    .Q_N(_3057_),
    .Q(\SegmentDisplay.digit3[1] ));
 sg13g2_dfrbp_1 _6463_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net326),
    .D(_0023_),
    .Q_N(_3058_),
    .Q(\SegmentDisplay.digit3[2] ));
 sg13g2_dfrbp_1 _6464_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net327),
    .D(_0024_),
    .Q_N(_3059_),
    .Q(\SegmentDisplay.digit3[3] ));
 sg13g2_dfrbp_1 _6465_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net328),
    .D(_0025_),
    .Q_N(_3060_),
    .Q(\SegmentDisplay.digit3[4] ));
 sg13g2_dfrbp_1 _6466_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net329),
    .D(_0026_),
    .Q_N(_3061_),
    .Q(\SegmentDisplay.digit3[5] ));
 sg13g2_dfrbp_1 _6467_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net330),
    .D(_0027_),
    .Q_N(_3062_),
    .Q(\SegmentDisplay.digit3[6] ));
 sg13g2_dfrbp_1 _6468_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net331),
    .D(net1679),
    .Q_N(_3063_),
    .Q(\uart_inst.uart_tx_inst.state[0] ));
 sg13g2_dfrbp_1 _6469_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net346),
    .D(net1577),
    .Q_N(_3064_),
    .Q(\uart_inst.uart_tx_inst.state[1] ));
 sg13g2_dfrbp_1 _6470_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net398),
    .D(net1547),
    .Q_N(_0109_),
    .Q(\uart_inst.uart_tx_inst.state[2] ));
 sg13g2_dfrbp_1 _6471_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net397),
    .D(_0520_),
    .Q_N(_2833_),
    .Q(\uart_tx_fifo_inst.fifo_valid[0] ));
 sg13g2_dfrbp_1 _6472_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net395),
    .D(net1508),
    .Q_N(_2832_),
    .Q(\uart_tx_fifo_inst.fifo_valid[1] ));
 sg13g2_dfrbp_1 _6473_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net393),
    .D(net1474),
    .Q_N(_2831_),
    .Q(\uart_tx_fifo_inst.fifo_valid[2] ));
 sg13g2_dfrbp_1 _6474_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net391),
    .D(_0523_),
    .Q_N(_2830_),
    .Q(\uart_tx_fifo_inst.fifo_valid[3] ));
 sg13g2_dfrbp_1 _6475_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net389),
    .D(net1340),
    .Q_N(_0121_),
    .Q(\uart_tx_fifo_inst.fifo_valid[4] ));
 sg13g2_dfrbp_1 _6476_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net387),
    .D(_0525_),
    .Q_N(_2829_),
    .Q(\uart_tx_fifo_inst.fifo_valid[5] ));
 sg13g2_dfrbp_1 _6477_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net385),
    .D(_0526_),
    .Q_N(_2828_),
    .Q(\uart_tx_fifo_inst.fifo_valid[6] ));
 sg13g2_dfrbp_1 _6478_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net383),
    .D(net1579),
    .Q_N(_2827_),
    .Q(\uart_tx_fifo_inst.fifo_valid[7] ));
 sg13g2_dfrbp_1 _6479_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net381),
    .D(_0528_),
    .Q_N(_2826_),
    .Q(\uart_tx_fifo_inst.fifo_valid[8] ));
 sg13g2_dfrbp_1 _6480_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net379),
    .D(_0529_),
    .Q_N(_2825_),
    .Q(\uart_tx_fifo_inst.fifo_valid[9] ));
 sg13g2_dfrbp_1 _6481_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net374),
    .D(_0530_),
    .Q_N(_2824_),
    .Q(tx_valid));
 sg13g2_dfrbp_1 _6482_ (.CLK(\SegmentDisplay.seg_driver.clk_reduced ),
    .RESET_B(net369),
    .D(_0531_),
    .Q_N(\SegmentDisplay.an[0] ),
    .Q(\SegmentDisplay.out_sel[0] ));
 sg13g2_dfrbp_1 _6483_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net368),
    .D(net1648),
    .Q_N(_2823_),
    .Q(_0076_));
 sg13g2_dfrbp_1 _6484_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net347),
    .D(net1689),
    .Q_N(_3065_),
    .Q(_0078_));
 sg13g2_dfrbp_1 _6485_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net348),
    .D(_0043_),
    .Q_N(_3066_),
    .Q(_0085_));
 sg13g2_dfrbp_1 _6486_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net349),
    .D(_0044_),
    .Q_N(_3067_),
    .Q(_0086_));
 sg13g2_dfrbp_1 _6487_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net350),
    .D(_0045_),
    .Q_N(_3068_),
    .Q(_0087_));
 sg13g2_dfrbp_1 _6488_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net351),
    .D(_0034_),
    .Q_N(_3069_),
    .Q(_0067_));
 sg13g2_dfrbp_1 _6489_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net354),
    .D(_0035_),
    .Q_N(_3070_),
    .Q(_0068_));
 sg13g2_dfrbp_1 _6490_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net367),
    .D(_0036_),
    .Q_N(_2822_),
    .Q(_0069_));
 sg13g2_dfrbp_1 _6491_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net366),
    .D(net1766),
    .Q_N(_2821_),
    .Q(_0094_));
 sg13g2_dfrbp_1 _6492_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net355),
    .D(_0535_),
    .Q_N(_3071_),
    .Q(_0096_));
 sg13g2_dfrbp_1 _6493_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net356),
    .D(_0000_),
    .Q_N(_3072_),
    .Q(\SegmentDisplay.digit0[0] ));
 sg13g2_dfrbp_1 _6494_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net357),
    .D(_0001_),
    .Q_N(_3073_),
    .Q(\SegmentDisplay.digit0[1] ));
 sg13g2_dfrbp_1 _6495_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net358),
    .D(_0002_),
    .Q_N(_3074_),
    .Q(\SegmentDisplay.digit0[2] ));
 sg13g2_dfrbp_1 _6496_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net359),
    .D(_0003_),
    .Q_N(_3075_),
    .Q(\SegmentDisplay.digit0[3] ));
 sg13g2_dfrbp_1 _6497_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net360),
    .D(_0004_),
    .Q_N(_3076_),
    .Q(\SegmentDisplay.digit0[4] ));
 sg13g2_dfrbp_1 _6498_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net361),
    .D(_0005_),
    .Q_N(_3077_),
    .Q(\SegmentDisplay.digit0[5] ));
 sg13g2_dfrbp_1 _6499_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net362),
    .D(_0006_),
    .Q_N(_3078_),
    .Q(\SegmentDisplay.digit0[6] ));
 sg13g2_dfrbp_1 _6500_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net363),
    .D(_0031_),
    .Q_N(_3079_),
    .Q(_0061_));
 sg13g2_dfrbp_1 _6501_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net370),
    .D(net1731),
    .Q_N(_3080_),
    .Q(_0062_));
 sg13g2_dfrbp_1 _6502_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net365),
    .D(net1750),
    .Q_N(_2820_),
    .Q(_0063_));
 sg13g2_dfrbp_1 _6503_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net364),
    .D(_0536_),
    .Q_N(_2819_),
    .Q(\output_value_inst.character_buff[8][0] ));
 sg13g2_dfrbp_1 _6504_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net352),
    .D(_0537_),
    .Q_N(_2818_),
    .Q(\output_value_inst.character_buff[8][1] ));
 sg13g2_dfrbp_1 _6505_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net344),
    .D(_0538_),
    .Q_N(_2817_),
    .Q(\output_value_inst.character_buff[8][2] ));
 sg13g2_dfrbp_1 _6506_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net342),
    .D(_0539_),
    .Q_N(_2816_),
    .Q(\output_value_inst.character_buff[8][3] ));
 sg13g2_dfrbp_1 _6507_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net340),
    .D(_0540_),
    .Q_N(_2815_),
    .Q(\output_value_inst.character_buff[8][4] ));
 sg13g2_dfrbp_1 _6508_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net371),
    .D(_0541_),
    .Q_N(_3081_),
    .Q(\output_value_inst.character_buff[8][6] ));
 sg13g2_dfrbp_1 _6509_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net372),
    .D(_0028_),
    .Q_N(_3082_),
    .Q(_0055_));
 sg13g2_dfrbp_1 _6510_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net376),
    .D(net1700),
    .Q_N(_3083_),
    .Q(_0056_));
 sg13g2_dfrbp_1 _6511_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net338),
    .D(_0030_),
    .Q_N(_2814_),
    .Q(_0057_));
 sg13g2_dfrbp_1 _6512_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net336),
    .D(_0542_),
    .Q_N(_0098_),
    .Q(\uart_inst.uart_rx_inst.SIGNAL_R ));
 sg13g2_dfrbp_1 _6513_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net334),
    .D(net1243),
    .Q_N(_2813_),
    .Q(_0088_));
 sg13g2_dfrbp_1 _6514_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net377),
    .D(_0544_),
    .Q_N(_3084_),
    .Q(_0090_));
 sg13g2_dfrbp_1 _6515_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net378),
    .D(_0037_),
    .Q_N(_3085_),
    .Q(_0073_));
 sg13g2_dfrbp_1 _6516_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net596),
    .D(net1722),
    .Q_N(_3086_),
    .Q(_0074_));
 sg13g2_dfrbp_1 _6517_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net333),
    .D(_0039_),
    .Q_N(_2812_),
    .Q(_0075_));
 sg13g2_dfrbp_1 _6518_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net332),
    .D(_0545_),
    .Q_N(_2811_),
    .Q(\uart_tx_fifo_inst.fifo[1][0] ));
 sg13g2_dfrbp_1 _6519_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net317),
    .D(_0546_),
    .Q_N(_2810_),
    .Q(\uart_tx_fifo_inst.fifo[1][1] ));
 sg13g2_dfrbp_1 _6520_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net315),
    .D(_0547_),
    .Q_N(_2809_),
    .Q(\uart_tx_fifo_inst.fifo[1][2] ));
 sg13g2_dfrbp_1 _6521_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net313),
    .D(_0548_),
    .Q_N(_2808_),
    .Q(\uart_tx_fifo_inst.fifo[1][3] ));
 sg13g2_dfrbp_1 _6522_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net311),
    .D(_0549_),
    .Q_N(_2807_),
    .Q(\uart_tx_fifo_inst.fifo[1][4] ));
 sg13g2_dfrbp_1 _6523_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net309),
    .D(_0550_),
    .Q_N(_2806_),
    .Q(\uart_tx_fifo_inst.fifo[1][5] ));
 sg13g2_dfrbp_1 _6524_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net307),
    .D(_0551_),
    .Q_N(_2805_),
    .Q(\uart_tx_fifo_inst.fifo[1][6] ));
 sg13g2_dfrbp_1 _6525_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net305),
    .D(_0552_),
    .Q_N(_2804_),
    .Q(\uart_tx_fifo_inst.fifo[2][0] ));
 sg13g2_dfrbp_1 _6526_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net303),
    .D(_0553_),
    .Q_N(_2803_),
    .Q(\uart_tx_fifo_inst.fifo[2][1] ));
 sg13g2_dfrbp_1 _6527_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net301),
    .D(_0554_),
    .Q_N(_2802_),
    .Q(\uart_tx_fifo_inst.fifo[2][2] ));
 sg13g2_dfrbp_1 _6528_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net299),
    .D(_0555_),
    .Q_N(_2801_),
    .Q(\uart_tx_fifo_inst.fifo[2][3] ));
 sg13g2_dfrbp_1 _6529_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net297),
    .D(_0556_),
    .Q_N(_2800_),
    .Q(\uart_tx_fifo_inst.fifo[2][4] ));
 sg13g2_dfrbp_1 _6530_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net295),
    .D(_0557_),
    .Q_N(_2799_),
    .Q(\uart_tx_fifo_inst.fifo[2][5] ));
 sg13g2_dfrbp_1 _6531_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net293),
    .D(_0558_),
    .Q_N(_2798_),
    .Q(\uart_tx_fifo_inst.fifo[2][6] ));
 sg13g2_dfrbp_1 _6532_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net291),
    .D(_0559_),
    .Q_N(_2797_),
    .Q(\uart_tx_fifo_inst.fifo[3][0] ));
 sg13g2_dfrbp_1 _6533_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net289),
    .D(_0560_),
    .Q_N(_2796_),
    .Q(\uart_tx_fifo_inst.fifo[3][1] ));
 sg13g2_dfrbp_1 _6534_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net287),
    .D(_0561_),
    .Q_N(_2795_),
    .Q(\uart_tx_fifo_inst.fifo[3][2] ));
 sg13g2_dfrbp_1 _6535_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net285),
    .D(_0562_),
    .Q_N(_2794_),
    .Q(\uart_tx_fifo_inst.fifo[3][3] ));
 sg13g2_dfrbp_1 _6536_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net283),
    .D(_0563_),
    .Q_N(_2793_),
    .Q(\uart_tx_fifo_inst.fifo[3][4] ));
 sg13g2_dfrbp_1 _6537_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net281),
    .D(_0564_),
    .Q_N(_2792_),
    .Q(\uart_tx_fifo_inst.fifo[3][5] ));
 sg13g2_dfrbp_1 _6538_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net279),
    .D(_0565_),
    .Q_N(_2791_),
    .Q(\uart_tx_fifo_inst.fifo[3][6] ));
 sg13g2_dfrbp_1 _6539_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net277),
    .D(_0566_),
    .Q_N(_2790_),
    .Q(\uart_tx_fifo_inst.fifo[4][0] ));
 sg13g2_dfrbp_1 _6540_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net275),
    .D(_0567_),
    .Q_N(_2789_),
    .Q(\uart_tx_fifo_inst.fifo[4][1] ));
 sg13g2_dfrbp_1 _6541_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net273),
    .D(_0568_),
    .Q_N(_2788_),
    .Q(\uart_tx_fifo_inst.fifo[4][2] ));
 sg13g2_dfrbp_1 _6542_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net271),
    .D(_0569_),
    .Q_N(_2787_),
    .Q(\uart_tx_fifo_inst.fifo[4][3] ));
 sg13g2_dfrbp_1 _6543_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net269),
    .D(_0570_),
    .Q_N(_2786_),
    .Q(\uart_tx_fifo_inst.fifo[4][4] ));
 sg13g2_dfrbp_1 _6544_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net267),
    .D(_0571_),
    .Q_N(_2785_),
    .Q(\uart_tx_fifo_inst.fifo[4][5] ));
 sg13g2_dfrbp_1 _6545_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net265),
    .D(_0572_),
    .Q_N(_2784_),
    .Q(\uart_tx_fifo_inst.fifo[4][6] ));
 sg13g2_dfrbp_1 _6546_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net263),
    .D(_0573_),
    .Q_N(_2783_),
    .Q(\uart_tx_fifo_inst.fifo[5][0] ));
 sg13g2_dfrbp_1 _6547_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net261),
    .D(_0574_),
    .Q_N(_2782_),
    .Q(\uart_tx_fifo_inst.fifo[5][1] ));
 sg13g2_dfrbp_1 _6548_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net259),
    .D(_0575_),
    .Q_N(_2781_),
    .Q(\uart_tx_fifo_inst.fifo[5][2] ));
 sg13g2_dfrbp_1 _6549_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net255),
    .D(_0576_),
    .Q_N(_2780_),
    .Q(\uart_tx_fifo_inst.fifo[5][3] ));
 sg13g2_dfrbp_1 _6550_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net251),
    .D(_0577_),
    .Q_N(_2779_),
    .Q(\uart_tx_fifo_inst.fifo[5][4] ));
 sg13g2_dfrbp_1 _6551_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net247),
    .D(_0578_),
    .Q_N(_2778_),
    .Q(\uart_tx_fifo_inst.fifo[5][5] ));
 sg13g2_dfrbp_1 _6552_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net79),
    .D(_0579_),
    .Q_N(_2777_),
    .Q(\uart_tx_fifo_inst.fifo[5][6] ));
 sg13g2_dfrbp_1 _6553_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net75),
    .D(_0580_),
    .Q_N(_2776_),
    .Q(\uart_tx_fifo_inst.fifo[6][0] ));
 sg13g2_dfrbp_1 _6554_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net71),
    .D(_0581_),
    .Q_N(_2775_),
    .Q(\uart_tx_fifo_inst.fifo[6][1] ));
 sg13g2_dfrbp_1 _6555_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net67),
    .D(_0582_),
    .Q_N(_2774_),
    .Q(\uart_tx_fifo_inst.fifo[6][2] ));
 sg13g2_dfrbp_1 _6556_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net63),
    .D(_0583_),
    .Q_N(_2773_),
    .Q(\uart_tx_fifo_inst.fifo[6][3] ));
 sg13g2_dfrbp_1 _6557_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net59),
    .D(_0584_),
    .Q_N(_2772_),
    .Q(\uart_tx_fifo_inst.fifo[6][4] ));
 sg13g2_dfrbp_1 _6558_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net55),
    .D(_0585_),
    .Q_N(_2771_),
    .Q(\uart_tx_fifo_inst.fifo[6][5] ));
 sg13g2_dfrbp_1 _6559_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net51),
    .D(_0586_),
    .Q_N(_2770_),
    .Q(\uart_tx_fifo_inst.fifo[6][6] ));
 sg13g2_dfrbp_1 _6560_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net47),
    .D(_0587_),
    .Q_N(_2769_),
    .Q(\uart_tx_fifo_inst.fifo[7][0] ));
 sg13g2_dfrbp_1 _6561_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net43),
    .D(_0588_),
    .Q_N(_2768_),
    .Q(\uart_tx_fifo_inst.fifo[7][1] ));
 sg13g2_dfrbp_1 _6562_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net39),
    .D(_0589_),
    .Q_N(_2767_),
    .Q(\uart_tx_fifo_inst.fifo[7][2] ));
 sg13g2_dfrbp_1 _6563_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net35),
    .D(_0590_),
    .Q_N(_2766_),
    .Q(\uart_tx_fifo_inst.fifo[7][3] ));
 sg13g2_dfrbp_1 _6564_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net31),
    .D(_0591_),
    .Q_N(_2765_),
    .Q(\uart_tx_fifo_inst.fifo[7][4] ));
 sg13g2_dfrbp_1 _6565_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net27),
    .D(_0592_),
    .Q_N(_2764_),
    .Q(\uart_tx_fifo_inst.fifo[7][5] ));
 sg13g2_dfrbp_1 _6566_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net23),
    .D(_0593_),
    .Q_N(_2763_),
    .Q(\uart_tx_fifo_inst.fifo[7][6] ));
 sg13g2_dfrbp_1 _6567_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net19),
    .D(net1313),
    .Q_N(_2762_),
    .Q(\output_value_inst.character_buff[9][0] ));
 sg13g2_dfrbp_1 _6568_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net15),
    .D(net1452),
    .Q_N(_2761_),
    .Q(\output_value_inst.character_buff[9][1] ));
 sg13g2_dfrbp_1 _6569_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net11),
    .D(net1194),
    .Q_N(_2760_),
    .Q(\output_value_inst.character_buff[9][2] ));
 sg13g2_dfrbp_1 _6570_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net592),
    .D(net1264),
    .Q_N(_2759_),
    .Q(\output_value_inst.character_buff[9][3] ));
 sg13g2_dfrbp_1 _6571_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net586),
    .D(net1456),
    .Q_N(_2758_),
    .Q(\output_value_inst.character_buff[9][4] ));
 sg13g2_dfrbp_1 _6572_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net582),
    .D(net1292),
    .Q_N(_2757_),
    .Q(\output_value_inst.character_buff[9][6] ));
 sg13g2_dfrbp_1 _6573_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net578),
    .D(net1438),
    .Q_N(_0155_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _6574_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net574),
    .D(net1476),
    .Q_N(_0153_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _6575_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net570),
    .D(_0602_),
    .Q_N(_2756_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _6576_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net566),
    .D(net755),
    .Q_N(_2755_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _6577_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net562),
    .D(_0604_),
    .Q_N(_2754_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _6578_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net558),
    .D(_0605_),
    .Q_N(_2753_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _6579_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net554),
    .D(_0606_),
    .Q_N(_2752_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _6580_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net550),
    .D(net1570),
    .Q_N(_0119_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _6581_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net546),
    .D(_0608_),
    .Q_N(_0130_),
    .Q(\SegmentDisplay.bcd2[0] ));
 sg13g2_dfrbp_1 _6582_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net542),
    .D(_0609_),
    .Q_N(_0127_),
    .Q(\SegmentDisplay.bcd2[1] ));
 sg13g2_dfrbp_1 _6583_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net538),
    .D(_0610_),
    .Q_N(_2751_),
    .Q(\SegmentDisplay.bcd2[2] ));
 sg13g2_dfrbp_1 _6584_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net534),
    .D(_0611_),
    .Q_N(_2750_),
    .Q(\SegmentDisplay.bcd2[3] ));
 sg13g2_dfrbp_1 _6585_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net530),
    .D(net977),
    .Q_N(_0144_),
    .Q(\SegmentDisplay.bcd3[0] ));
 sg13g2_dfrbp_1 _6586_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net526),
    .D(net983),
    .Q_N(_0143_),
    .Q(\SegmentDisplay.bcd3[1] ));
 sg13g2_dfrbp_1 _6587_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net522),
    .D(_0614_),
    .Q_N(_2749_),
    .Q(\SegmentDisplay.bcd3[2] ));
 sg13g2_dfrbp_1 _6588_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net518),
    .D(_0615_),
    .Q_N(_2748_),
    .Q(\SegmentDisplay.bcd3[3] ));
 sg13g2_dfrbp_1 _6589_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net514),
    .D(_0616_),
    .Q_N(_2747_),
    .Q(\Led_Cycle_inst.buttons[0] ));
 sg13g2_dfrbp_1 _6590_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net510),
    .D(_0617_),
    .Q_N(_2746_),
    .Q(\Led_Cycle_inst.buttons[1] ));
 sg13g2_dfrbp_1 _6591_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net506),
    .D(_0618_),
    .Q_N(_2745_),
    .Q(\Led_Cycle_inst.buttons[2] ));
 sg13g2_dfrbp_1 _6592_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net502),
    .D(_0619_),
    .Q_N(_2744_),
    .Q(\Led_Cycle_inst.buttons[3] ));
 sg13g2_dfrbp_1 _6593_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net498),
    .D(net1303),
    .Q_N(_0111_),
    .Q(\Led_Cycle_inst.buttons[4] ));
 sg13g2_dfrbp_1 _6594_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net494),
    .D(_0621_),
    .Q_N(_2743_),
    .Q(\output_value_inst.character_buff[7][0] ));
 sg13g2_dfrbp_1 _6595_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net490),
    .D(_0622_),
    .Q_N(_2742_),
    .Q(\output_value_inst.character_buff[7][1] ));
 sg13g2_dfrbp_1 _6596_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net486),
    .D(_0623_),
    .Q_N(_2741_),
    .Q(\output_value_inst.character_buff[7][2] ));
 sg13g2_dfrbp_1 _6597_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net482),
    .D(_0624_),
    .Q_N(_2740_),
    .Q(\output_value_inst.character_buff[7][3] ));
 sg13g2_dfrbp_1 _6598_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net478),
    .D(_0625_),
    .Q_N(_2739_),
    .Q(\output_value_inst.character_buff[7][4] ));
 sg13g2_dfrbp_1 _6599_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net474),
    .D(_0626_),
    .Q_N(_2738_),
    .Q(\output_value_inst.character_buff[7][6] ));
 sg13g2_dfrbp_1 _6600_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net470),
    .D(_0627_),
    .Q_N(_2737_),
    .Q(\output_value_inst.character_buff[6][0] ));
 sg13g2_dfrbp_1 _6601_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net466),
    .D(_0628_),
    .Q_N(_2736_),
    .Q(\output_value_inst.character_buff[6][1] ));
 sg13g2_dfrbp_1 _6602_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net462),
    .D(_0629_),
    .Q_N(_2735_),
    .Q(\output_value_inst.character_buff[6][2] ));
 sg13g2_dfrbp_1 _6603_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net458),
    .D(_0630_),
    .Q_N(_2734_),
    .Q(\output_value_inst.character_buff[6][3] ));
 sg13g2_dfrbp_1 _6604_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net454),
    .D(_0631_),
    .Q_N(_2733_),
    .Q(\output_value_inst.character_buff[6][4] ));
 sg13g2_dfrbp_1 _6605_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net450),
    .D(_0632_),
    .Q_N(_2732_),
    .Q(\output_value_inst.character_buff[6][6] ));
 sg13g2_dfrbp_1 _6606_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net446),
    .D(_0633_),
    .Q_N(_2731_),
    .Q(\output_value_inst.character_buff[5][0] ));
 sg13g2_dfrbp_1 _6607_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net442),
    .D(_0634_),
    .Q_N(_2730_),
    .Q(\output_value_inst.character_buff[5][1] ));
 sg13g2_dfrbp_1 _6608_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net438),
    .D(_0635_),
    .Q_N(_2729_),
    .Q(\output_value_inst.character_buff[5][2] ));
 sg13g2_dfrbp_1 _6609_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net434),
    .D(_0636_),
    .Q_N(_2728_),
    .Q(\output_value_inst.character_buff[5][3] ));
 sg13g2_dfrbp_1 _6610_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net430),
    .D(net1283),
    .Q_N(_2727_),
    .Q(\output_value_inst.character_buff[5][4] ));
 sg13g2_dfrbp_1 _6611_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net426),
    .D(net1188),
    .Q_N(_2726_),
    .Q(\output_value_inst.character_buff[5][6] ));
 sg13g2_dfrbp_1 _6612_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net422),
    .D(_0639_),
    .Q_N(_2725_),
    .Q(\output_value_inst.character_buff[4][0] ));
 sg13g2_dfrbp_1 _6613_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net418),
    .D(_0640_),
    .Q_N(_2724_),
    .Q(\output_value_inst.character_buff[4][1] ));
 sg13g2_dfrbp_1 _6614_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net414),
    .D(_0641_),
    .Q_N(_2723_),
    .Q(\output_value_inst.character_buff[4][2] ));
 sg13g2_dfrbp_1 _6615_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net410),
    .D(_0642_),
    .Q_N(_2722_),
    .Q(\output_value_inst.character_buff[4][3] ));
 sg13g2_dfrbp_1 _6616_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net406),
    .D(_0643_),
    .Q_N(_2721_),
    .Q(\output_value_inst.character_buff[4][4] ));
 sg13g2_dfrbp_1 _6617_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net402),
    .D(_0644_),
    .Q_N(_2720_),
    .Q(\output_value_inst.character_buff[4][6] ));
 sg13g2_dfrbp_1 _6618_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net396),
    .D(_0645_),
    .Q_N(_2719_),
    .Q(\output_value_inst.character_buff[3][0] ));
 sg13g2_dfrbp_1 _6619_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net392),
    .D(_0646_),
    .Q_N(_2718_),
    .Q(\output_value_inst.character_buff[3][1] ));
 sg13g2_dfrbp_1 _6620_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net388),
    .D(_0647_),
    .Q_N(_2717_),
    .Q(\output_value_inst.character_buff[3][2] ));
 sg13g2_dfrbp_1 _6621_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net384),
    .D(_0648_),
    .Q_N(_2716_),
    .Q(\output_value_inst.character_buff[3][3] ));
 sg13g2_dfrbp_1 _6622_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net380),
    .D(_0649_),
    .Q_N(_2715_),
    .Q(\output_value_inst.character_buff[3][4] ));
 sg13g2_dfrbp_1 _6623_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net373),
    .D(_0650_),
    .Q_N(_2714_),
    .Q(\output_value_inst.character_buff[3][5] ));
 sg13g2_dfrbp_1 _6624_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net345),
    .D(_0651_),
    .Q_N(_2713_),
    .Q(\output_value_inst.character_buff[3][6] ));
 sg13g2_dfrbp_1 _6625_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net341),
    .D(_0652_),
    .Q_N(_2712_),
    .Q(\output_value_inst.character_buff[2][0] ));
 sg13g2_dfrbp_1 _6626_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net337),
    .D(net988),
    .Q_N(_2711_),
    .Q(\output_value_inst.character_buff[2][1] ));
 sg13g2_dfrbp_1 _6627_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net318),
    .D(_0654_),
    .Q_N(_2710_),
    .Q(\output_value_inst.character_buff[2][2] ));
 sg13g2_dfrbp_1 _6628_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net314),
    .D(_0655_),
    .Q_N(_2709_),
    .Q(\output_value_inst.character_buff[2][3] ));
 sg13g2_dfrbp_1 _6629_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net310),
    .D(net1082),
    .Q_N(_2708_),
    .Q(\output_value_inst.character_buff[2][4] ));
 sg13g2_dfrbp_1 _6630_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net306),
    .D(net1226),
    .Q_N(_2707_),
    .Q(\output_value_inst.character_buff[2][5] ));
 sg13g2_dfrbp_1 _6631_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net302),
    .D(_0658_),
    .Q_N(_2706_),
    .Q(\output_value_inst.character_buff[2][6] ));
 sg13g2_dfrbp_1 _6632_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net298),
    .D(net1499),
    .Q_N(_2705_),
    .Q(\output_value_inst.character_buff[1][0] ));
 sg13g2_dfrbp_1 _6633_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net294),
    .D(_0660_),
    .Q_N(_2704_),
    .Q(\output_value_inst.character_buff[1][1] ));
 sg13g2_dfrbp_1 _6634_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net290),
    .D(_0661_),
    .Q_N(_2703_),
    .Q(\output_value_inst.character_buff[1][2] ));
 sg13g2_dfrbp_1 _6635_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net286),
    .D(_0662_),
    .Q_N(_2702_),
    .Q(\output_value_inst.character_buff[1][3] ));
 sg13g2_dfrbp_1 _6636_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net282),
    .D(_0663_),
    .Q_N(_2701_),
    .Q(\output_value_inst.character_buff[1][4] ));
 sg13g2_dfrbp_1 _6637_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net278),
    .D(_0664_),
    .Q_N(_2700_),
    .Q(\output_value_inst.character_buff[1][5] ));
 sg13g2_dfrbp_1 _6638_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net274),
    .D(net1221),
    .Q_N(_2699_),
    .Q(\output_value_inst.character_buff[1][6] ));
 sg13g2_dfrbp_1 _6639_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net270),
    .D(net1515),
    .Q_N(_2698_),
    .Q(\output_value_inst.character_buff[0][0] ));
 sg13g2_dfrbp_1 _6640_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net266),
    .D(net1442),
    .Q_N(_2697_),
    .Q(\output_value_inst.character_buff[0][1] ));
 sg13g2_dfrbp_1 _6641_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net262),
    .D(net1146),
    .Q_N(_2696_),
    .Q(\output_value_inst.character_buff[0][2] ));
 sg13g2_dfrbp_1 _6642_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net257),
    .D(net1581),
    .Q_N(_2695_),
    .Q(\output_value_inst.character_buff[0][3] ));
 sg13g2_dfrbp_1 _6643_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net249),
    .D(net1459),
    .Q_N(_2694_),
    .Q(\output_value_inst.character_buff[0][4] ));
 sg13g2_dfrbp_1 _6644_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net77),
    .D(net1490),
    .Q_N(_2693_),
    .Q(\output_value_inst.character_buff[0][5] ));
 sg13g2_dfrbp_1 _6645_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net69),
    .D(net1568),
    .Q_N(_2692_),
    .Q(\output_value_inst.character_buff[0][6] ));
 sg13g2_dfrbp_1 _6646_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net61),
    .D(net1027),
    .Q_N(_2691_),
    .Q(\output_value_inst.output_data[0] ));
 sg13g2_dfrbp_1 _6647_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net53),
    .D(net714),
    .Q_N(_2690_),
    .Q(\output_value_inst.output_data[1] ));
 sg13g2_dfrbp_1 _6648_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net45),
    .D(net973),
    .Q_N(_2689_),
    .Q(\output_value_inst.output_data[2] ));
 sg13g2_dfrbp_1 _6649_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net37),
    .D(net717),
    .Q_N(_2688_),
    .Q(\output_value_inst.output_data[3] ));
 sg13g2_dfrbp_1 _6650_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net29),
    .D(net689),
    .Q_N(_2687_),
    .Q(\output_value_inst.output_data[4] ));
 sg13g2_dfrbp_1 _6651_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net21),
    .D(net723),
    .Q_N(_2686_),
    .Q(\output_value_inst.output_data[5] ));
 sg13g2_dfrbp_1 _6652_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net13),
    .D(net708),
    .Q_N(_2685_),
    .Q(\output_value_inst.output_data[6] ));
 sg13g2_dfrbp_1 _6653_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net588),
    .D(_0680_),
    .Q_N(_2684_),
    .Q(\output_value_inst.send_element_data ));
 sg13g2_dfrbp_1 _6654_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net580),
    .D(_0681_),
    .Q_N(_0165_),
    .Q(\output_value_inst.send_led_data ));
 sg13g2_dfrbp_1 _6655_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net572),
    .D(_0682_),
    .Q_N(_0099_),
    .Q(\output_value_inst.ready_to_send ));
 sg13g2_dfrbp_1 _6656_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net564),
    .D(_0683_),
    .Q_N(_0164_),
    .Q(\output_value_inst.element_data_reg[0] ));
 sg13g2_dfrbp_1 _6657_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net556),
    .D(_0684_),
    .Q_N(_0100_),
    .Q(\output_value_inst.element_data_reg[1] ));
 sg13g2_dfrbp_1 _6658_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net548),
    .D(_0685_),
    .Q_N(_0101_),
    .Q(\output_value_inst.element_data_reg[2] ));
 sg13g2_dfrbp_1 _6659_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net540),
    .D(_0686_),
    .Q_N(_0102_),
    .Q(\output_value_inst.element_data_reg[3] ));
 sg13g2_dfrbp_1 _6660_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net532),
    .D(_0687_),
    .Q_N(_0103_),
    .Q(\output_value_inst.element_data_reg[4] ));
 sg13g2_dfrbp_1 _6661_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net524),
    .D(net1015),
    .Q_N(_0104_),
    .Q(\output_value_inst.element_data_reg[5] ));
 sg13g2_dfrbp_1 _6662_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net516),
    .D(_0689_),
    .Q_N(_0105_),
    .Q(\output_value_inst.element_data_reg[6] ));
 sg13g2_dfrbp_1 _6663_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net508),
    .D(_0690_),
    .Q_N(_0149_),
    .Q(\output_value_inst.element_data_reg[7] ));
 sg13g2_dfrbp_1 _6664_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net500),
    .D(_0691_),
    .Q_N(_0151_),
    .Q(\output_value_inst.element_data_reg[8] ));
 sg13g2_dfrbp_1 _6665_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net492),
    .D(_0692_),
    .Q_N(_2683_),
    .Q(\output_value_inst.element_data_reg[9] ));
 sg13g2_dfrbp_1 _6666_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net484),
    .D(_0693_),
    .Q_N(_2682_),
    .Q(\output_value_inst.element_data_reg[10] ));
 sg13g2_dfrbp_1 _6667_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net476),
    .D(net1466),
    .Q_N(_0150_),
    .Q(\output_value_inst.element_data_reg[11] ));
 sg13g2_dfrbp_1 _6668_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net468),
    .D(net1156),
    .Q_N(_0124_),
    .Q(\output_value_inst.led_data_reg[0] ));
 sg13g2_dfrbp_1 _6669_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net460),
    .D(_0696_),
    .Q_N(_2681_),
    .Q(\output_value_inst.led_data_reg[1] ));
 sg13g2_dfrbp_1 _6670_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net452),
    .D(_0697_),
    .Q_N(_2680_),
    .Q(\output_value_inst.led_data_reg[2] ));
 sg13g2_dfrbp_1 _6671_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net444),
    .D(net1089),
    .Q_N(_0122_),
    .Q(\output_value_inst.led_data_reg[3] ));
 sg13g2_dfrbp_1 _6672_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net436),
    .D(net1165),
    .Q_N(_0162_),
    .Q(\output_value_inst.led_data_reg[4] ));
 sg13g2_dfrbp_1 _6673_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net428),
    .D(_0700_),
    .Q_N(_2679_),
    .Q(\output_value_inst.led_data_reg[5] ));
 sg13g2_dfrbp_1 _6674_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net420),
    .D(_0701_),
    .Q_N(_2678_),
    .Q(\output_value_inst.led_data_reg[6] ));
 sg13g2_dfrbp_1 _6675_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net412),
    .D(net1065),
    .Q_N(_0160_),
    .Q(\output_value_inst.led_data_reg[7] ));
 sg13g2_dfrbp_1 _6676_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net404),
    .D(net1122),
    .Q_N(_0147_),
    .Q(\output_value_inst.led_data_reg[8] ));
 sg13g2_dfrbp_1 _6677_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net394),
    .D(_0704_),
    .Q_N(_2677_),
    .Q(\output_value_inst.led_data_reg[9] ));
 sg13g2_dfrbp_1 _6678_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net386),
    .D(_0705_),
    .Q_N(_2676_),
    .Q(\output_value_inst.led_data_reg[10] ));
 sg13g2_dfrbp_1 _6679_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net375),
    .D(net1110),
    .Q_N(_0145_),
    .Q(\output_value_inst.led_data_reg[11] ));
 sg13g2_dfrbp_1 _6680_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net343),
    .D(net1183),
    .Q_N(_0141_),
    .Q(\output_value_inst.led_data_reg[12] ));
 sg13g2_dfrbp_1 _6681_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net335),
    .D(_0708_),
    .Q_N(_2675_),
    .Q(\output_value_inst.led_data_reg[13] ));
 sg13g2_dfrbp_1 _6682_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net312),
    .D(_0709_),
    .Q_N(_2674_),
    .Q(\output_value_inst.led_data_reg[14] ));
 sg13g2_dfrbp_1 _6683_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net304),
    .D(net1273),
    .Q_N(_0139_),
    .Q(\output_value_inst.led_data_reg[15] ));
 sg13g2_dfrbp_1 _6684_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net296),
    .D(_0711_),
    .Q_N(_0159_),
    .Q(\output_value_inst.output_valid ));
 sg13g2_dfrbp_1 _6685_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net288),
    .D(_0712_),
    .Q_N(_2673_),
    .Q(\uart_tx_fifo_inst.fifo[0][0] ));
 sg13g2_dfrbp_1 _6686_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net280),
    .D(_0713_),
    .Q_N(_2672_),
    .Q(\uart_tx_fifo_inst.fifo[0][1] ));
 sg13g2_dfrbp_1 _6687_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net272),
    .D(_0714_),
    .Q_N(_2671_),
    .Q(\uart_tx_fifo_inst.fifo[0][2] ));
 sg13g2_dfrbp_1 _6688_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net264),
    .D(_0715_),
    .Q_N(_2670_),
    .Q(\uart_tx_fifo_inst.fifo[0][3] ));
 sg13g2_dfrbp_1 _6689_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net253),
    .D(_0716_),
    .Q_N(_2669_),
    .Q(\uart_tx_fifo_inst.fifo[0][4] ));
 sg13g2_dfrbp_1 _6690_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net73),
    .D(_0717_),
    .Q_N(_2668_),
    .Q(\uart_tx_fifo_inst.fifo[0][5] ));
 sg13g2_dfrbp_1 _6691_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net57),
    .D(_0718_),
    .Q_N(_2667_),
    .Q(\uart_tx_fifo_inst.fifo[0][6] ));
 sg13g2_dfrbp_1 _6692_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net41),
    .D(net1658),
    .Q_N(_2666_),
    .Q(_0058_));
 sg13g2_dfrbp_1 _6693_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net33),
    .D(net1683),
    .Q_N(_2665_),
    .Q(_0060_));
 sg13g2_dfrbp_1 _6694_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net25),
    .D(net1351),
    .Q_N(_2664_),
    .Q(\uart_inst.uart_tx_inst.DATA_REG[0] ));
 sg13g2_dfrbp_1 _6695_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net594),
    .D(net1321),
    .Q_N(_2663_),
    .Q(\uart_inst.uart_tx_inst.DATA_REG[1] ));
 sg13g2_dfrbp_1 _6696_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net576),
    .D(net1308),
    .Q_N(_2662_),
    .Q(\uart_inst.uart_tx_inst.DATA_REG[2] ));
 sg13g2_dfrbp_1 _6697_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net560),
    .D(_0724_),
    .Q_N(_2661_),
    .Q(\uart_inst.uart_tx_inst.DATA_REG[3] ));
 sg13g2_dfrbp_1 _6698_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net544),
    .D(net1408),
    .Q_N(_2660_),
    .Q(\uart_inst.uart_tx_inst.DATA_REG[4] ));
 sg13g2_dfrbp_1 _6699_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net528),
    .D(net1228),
    .Q_N(_2659_),
    .Q(\uart_inst.uart_tx_inst.DATA_REG[5] ));
 sg13g2_dfrbp_1 _6700_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net512),
    .D(net1324),
    .Q_N(_2658_),
    .Q(\uart_inst.uart_tx_inst.DATA_REG[6] ));
 sg13g2_dfrbp_1 _6701_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net496),
    .D(net634),
    .Q_N(_0207_),
    .Q(\SegmentDisplay.seg_driver.clk_reducer.counter[0] ));
 sg13g2_dfrbp_1 _6702_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net488),
    .D(net1561),
    .Q_N(_2657_),
    .Q(\SegmentDisplay.seg_driver.clk_reducer.counter[1] ));
 sg13g2_dfrbp_1 _6703_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net480),
    .D(_0730_),
    .Q_N(_2656_),
    .Q(\SegmentDisplay.seg_driver.clk_reducer.counter[2] ));
 sg13g2_dfrbp_1 _6704_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net472),
    .D(net1076),
    .Q_N(_2655_),
    .Q(\SegmentDisplay.seg_driver.clk_reducer.counter[3] ));
 sg13g2_dfrbp_1 _6705_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net464),
    .D(_0732_),
    .Q_N(_2654_),
    .Q(\SegmentDisplay.seg_driver.clk_reducer.counter[4] ));
 sg13g2_dfrbp_1 _6706_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net456),
    .D(_0733_),
    .Q_N(_2653_),
    .Q(\SegmentDisplay.seg_driver.clk_reducer.counter[5] ));
 sg13g2_dfrbp_1 _6707_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net448),
    .D(_0734_),
    .Q_N(_2652_),
    .Q(\SegmentDisplay.seg_driver.clk_reducer.counter[6] ));
 sg13g2_dfrbp_1 _6708_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net440),
    .D(net1141),
    .Q_N(_2651_),
    .Q(\SegmentDisplay.seg_driver.clk_reducer.counter[7] ));
 sg13g2_dfrbp_1 _6709_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net432),
    .D(_0736_),
    .Q_N(_2650_),
    .Q(\SegmentDisplay.seg_driver.clk_reducer.counter[8] ));
 sg13g2_dfrbp_1 _6710_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net424),
    .D(_0737_),
    .Q_N(_2649_),
    .Q(\SegmentDisplay.seg_driver.clk_reducer.counter[9] ));
 sg13g2_dfrbp_1 _6711_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net416),
    .D(_0738_),
    .Q_N(_2648_),
    .Q(\SegmentDisplay.seg_driver.clk_reducer.counter[10] ));
 sg13g2_dfrbp_1 _6712_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net408),
    .D(net1394),
    .Q_N(_2647_),
    .Q(\SegmentDisplay.seg_driver.clk_reducer.counter[11] ));
 sg13g2_dfrbp_1 _6713_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net400),
    .D(_0740_),
    .Q_N(_2627_),
    .Q(\SegmentDisplay.seg_driver.clk_reducer.counter[12] ));
 sg13g2_dfrbp_1 _6714_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net390),
    .D(_0741_),
    .Q_N(_2646_),
    .Q(\SegmentDisplay.seg_driver.clk_reduced ));
 sg13g2_dfrbp_1 _6715_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net382),
    .D(net645),
    .Q_N(_0206_),
    .Q(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[0] ));
 sg13g2_dfrbp_1 _6716_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net353),
    .D(net1718),
    .Q_N(_2645_),
    .Q(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[1] ));
 sg13g2_dfrbp_1 _6717_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net339),
    .D(net1129),
    .Q_N(_2644_),
    .Q(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[2] ));
 sg13g2_dfrbp_1 _6718_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net316),
    .D(_0745_),
    .Q_N(_0177_),
    .Q(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[3] ));
 sg13g2_dfrbp_1 _6719_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net308),
    .D(_0746_),
    .Q_N(_2643_),
    .Q(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[4] ));
 sg13g2_dfrbp_1 _6720_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net300),
    .D(net1061),
    .Q_N(_0176_),
    .Q(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[5] ));
 sg13g2_dfrbp_1 _6721_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net292),
    .D(_0748_),
    .Q_N(_2642_),
    .Q(\tx_data[0] ));
 sg13g2_dfrbp_1 _6722_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net284),
    .D(_0749_),
    .Q_N(_2641_),
    .Q(\tx_data[1] ));
 sg13g2_dfrbp_1 _6723_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net276),
    .D(_0750_),
    .Q_N(_2640_),
    .Q(\tx_data[2] ));
 sg13g2_dfrbp_1 _6724_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net268),
    .D(net1315),
    .Q_N(_2639_),
    .Q(\tx_data[3] ));
 sg13g2_dfrbp_1 _6725_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net260),
    .D(_0752_),
    .Q_N(_2638_),
    .Q(\uart_inst.tx_data[4] ));
 sg13g2_dfrbp_1 _6726_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net81),
    .D(net1374),
    .Q_N(_2637_),
    .Q(\uart_inst.tx_data[5] ));
 sg13g2_dfrbp_1 _6727_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net65),
    .D(_0754_),
    .Q_N(_2636_),
    .Q(\uart_inst.tx_data[6] ));
 sg13g2_dfrbp_1 _6728_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net49),
    .D(_0755_),
    .Q_N(_2635_),
    .Q(\uart_tx_fifo_inst.fifo[9][0] ));
 sg13g2_dfrbp_1 _6729_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net584),
    .D(_0756_),
    .Q_N(_2634_),
    .Q(\uart_tx_fifo_inst.fifo[9][1] ));
 sg13g2_dfrbp_1 _6730_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net552),
    .D(_0757_),
    .Q_N(_2633_),
    .Q(\uart_tx_fifo_inst.fifo[9][2] ));
 sg13g2_dfrbp_1 _6731_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net520),
    .D(_0758_),
    .Q_N(_2632_),
    .Q(\uart_tx_fifo_inst.fifo[9][3] ));
 sg13g2_dfrbp_1 _6732_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net17),
    .D(_0759_),
    .Q_N(_2631_),
    .Q(\uart_tx_fifo_inst.fifo[9][4] ));
 sg13g2_dfrbp_1 _6733_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net536),
    .D(_0760_),
    .Q_N(_2630_),
    .Q(\uart_tx_fifo_inst.fifo[9][5] ));
 sg13g2_dfrbp_1 _6734_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net597),
    .D(_0761_),
    .Q_N(_3087_),
    .Q(\uart_tx_fifo_inst.fifo[9][6] ));
 sg13g2_dfrbp_1 _6735_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net598),
    .D(_0007_),
    .Q_N(_3088_),
    .Q(\SegmentDisplay.digit1[0] ));
 sg13g2_dfrbp_1 _6736_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net599),
    .D(_0008_),
    .Q_N(_3089_),
    .Q(\SegmentDisplay.digit1[1] ));
 sg13g2_dfrbp_1 _6737_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net600),
    .D(_0009_),
    .Q_N(_3090_),
    .Q(\SegmentDisplay.digit1[2] ));
 sg13g2_dfrbp_1 _6738_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net601),
    .D(_0010_),
    .Q_N(_3091_),
    .Q(\SegmentDisplay.digit1[3] ));
 sg13g2_dfrbp_1 _6739_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net602),
    .D(_0011_),
    .Q_N(_3092_),
    .Q(\SegmentDisplay.digit1[4] ));
 sg13g2_dfrbp_1 _6740_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net504),
    .D(_0012_),
    .Q_N(_3093_),
    .Q(\SegmentDisplay.digit1[5] ));
 sg13g2_dfrbp_1 _6741_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net568),
    .D(_0013_),
    .Q_N(_2629_),
    .Q(\SegmentDisplay.digit1[6] ));
 sg13g2_tiehi _6353__12 (.L_HI(net12));
 sg13g2_tiehi _6652__13 (.L_HI(net13));
 sg13g2_tiehi _6352__14 (.L_HI(net14));
 sg13g2_tiehi _6568__15 (.L_HI(net15));
 sg13g2_tiehi _6351__16 (.L_HI(net16));
 sg13g2_tiehi _6732__17 (.L_HI(net17));
 sg13g2_tiehi _6350__18 (.L_HI(net18));
 sg13g2_tiehi _6567__19 (.L_HI(net19));
 sg13g2_tiehi _6349__20 (.L_HI(net20));
 sg13g2_tiehi _6651__21 (.L_HI(net21));
 sg13g2_tiehi _6348__22 (.L_HI(net22));
 sg13g2_tiehi _6566__23 (.L_HI(net23));
 sg13g2_tiehi _6347__24 (.L_HI(net24));
 sg13g2_tiehi _6694__25 (.L_HI(net25));
 sg13g2_tiehi _6346__26 (.L_HI(net26));
 sg13g2_tiehi _6565__27 (.L_HI(net27));
 sg13g2_tiehi _6345__28 (.L_HI(net28));
 sg13g2_tiehi _6650__29 (.L_HI(net29));
 sg13g2_tiehi _6344__30 (.L_HI(net30));
 sg13g2_tiehi _6564__31 (.L_HI(net31));
 sg13g2_tiehi _6343__32 (.L_HI(net32));
 sg13g2_tiehi _6693__33 (.L_HI(net33));
 sg13g2_tiehi _6342__34 (.L_HI(net34));
 sg13g2_tiehi _6563__35 (.L_HI(net35));
 sg13g2_tiehi _6341__36 (.L_HI(net36));
 sg13g2_tiehi _6649__37 (.L_HI(net37));
 sg13g2_tiehi _6340__38 (.L_HI(net38));
 sg13g2_tiehi _6562__39 (.L_HI(net39));
 sg13g2_tiehi _6339__40 (.L_HI(net40));
 sg13g2_tiehi _6692__41 (.L_HI(net41));
 sg13g2_tiehi _6338__42 (.L_HI(net42));
 sg13g2_tiehi _6561__43 (.L_HI(net43));
 sg13g2_tiehi _6337__44 (.L_HI(net44));
 sg13g2_tiehi _6648__45 (.L_HI(net45));
 sg13g2_tiehi _6336__46 (.L_HI(net46));
 sg13g2_tiehi _6560__47 (.L_HI(net47));
 sg13g2_tiehi _6335__48 (.L_HI(net48));
 sg13g2_tiehi _6728__49 (.L_HI(net49));
 sg13g2_tiehi _6334__50 (.L_HI(net50));
 sg13g2_tiehi _6559__51 (.L_HI(net51));
 sg13g2_tiehi _6333__52 (.L_HI(net52));
 sg13g2_tiehi _6647__53 (.L_HI(net53));
 sg13g2_tiehi _6332__54 (.L_HI(net54));
 sg13g2_tiehi _6558__55 (.L_HI(net55));
 sg13g2_tiehi _6331__56 (.L_HI(net56));
 sg13g2_tiehi _6691__57 (.L_HI(net57));
 sg13g2_tiehi _6330__58 (.L_HI(net58));
 sg13g2_tiehi _6557__59 (.L_HI(net59));
 sg13g2_tiehi _6329__60 (.L_HI(net60));
 sg13g2_tiehi _6646__61 (.L_HI(net61));
 sg13g2_tiehi _6328__62 (.L_HI(net62));
 sg13g2_tiehi _6556__63 (.L_HI(net63));
 sg13g2_tiehi _6327__64 (.L_HI(net64));
 sg13g2_tiehi _6727__65 (.L_HI(net65));
 sg13g2_tiehi _6326__66 (.L_HI(net66));
 sg13g2_tiehi _6555__67 (.L_HI(net67));
 sg13g2_tiehi _6325__68 (.L_HI(net68));
 sg13g2_tiehi _6645__69 (.L_HI(net69));
 sg13g2_tiehi _6324__70 (.L_HI(net70));
 sg13g2_tiehi _6554__71 (.L_HI(net71));
 sg13g2_tiehi _6323__72 (.L_HI(net72));
 sg13g2_tiehi _6690__73 (.L_HI(net73));
 sg13g2_tiehi _6322__74 (.L_HI(net74));
 sg13g2_tiehi _6553__75 (.L_HI(net75));
 sg13g2_tiehi _6321__76 (.L_HI(net76));
 sg13g2_tiehi _6644__77 (.L_HI(net77));
 sg13g2_tiehi _6320__78 (.L_HI(net78));
 sg13g2_tiehi _6552__79 (.L_HI(net79));
 sg13g2_tiehi _6319__80 (.L_HI(net80));
 sg13g2_tiehi _6726__81 (.L_HI(net81));
 sg13g2_tiehi _6318__82 (.L_HI(net82));
 sg13g2_tiehi _6317__83 (.L_HI(net83));
 sg13g2_tiehi _6306__84 (.L_HI(net84));
 sg13g2_tiehi _6305__85 (.L_HI(net85));
 sg13g2_tiehi _6304__86 (.L_HI(net86));
 sg13g2_tiehi _6303__87 (.L_HI(net87));
 sg13g2_tiehi _6302__88 (.L_HI(net88));
 sg13g2_tiehi _6301__89 (.L_HI(net89));
 sg13g2_tiehi _6300__90 (.L_HI(net90));
 sg13g2_tiehi _6299__91 (.L_HI(net91));
 sg13g2_tiehi _6298__92 (.L_HI(net92));
 sg13g2_tiehi _6292__93 (.L_HI(net93));
 sg13g2_tiehi _6291__94 (.L_HI(net94));
 sg13g2_tiehi _6290__95 (.L_HI(net95));
 sg13g2_tiehi _6289__96 (.L_HI(net96));
 sg13g2_tiehi _6288__97 (.L_HI(net97));
 sg13g2_tiehi _6287__98 (.L_HI(net98));
 sg13g2_tiehi _6286__99 (.L_HI(net99));
 sg13g2_tiehi _6285__100 (.L_HI(net100));
 sg13g2_tiehi _6284__101 (.L_HI(net101));
 sg13g2_tiehi _6283__102 (.L_HI(net102));
 sg13g2_tiehi _6282__103 (.L_HI(net103));
 sg13g2_tiehi _6281__104 (.L_HI(net104));
 sg13g2_tiehi _6280__105 (.L_HI(net105));
 sg13g2_tiehi _6279__106 (.L_HI(net106));
 sg13g2_tiehi _6278__107 (.L_HI(net107));
 sg13g2_tiehi _6277__108 (.L_HI(net108));
 sg13g2_tiehi _6276__109 (.L_HI(net109));
 sg13g2_tiehi _6275__110 (.L_HI(net110));
 sg13g2_tiehi _6274__111 (.L_HI(net111));
 sg13g2_tiehi _6273__112 (.L_HI(net112));
 sg13g2_tiehi _6272__113 (.L_HI(net113));
 sg13g2_tiehi _6271__114 (.L_HI(net114));
 sg13g2_tiehi _6270__115 (.L_HI(net115));
 sg13g2_tiehi _6269__116 (.L_HI(net116));
 sg13g2_tiehi _6268__117 (.L_HI(net117));
 sg13g2_tiehi _6267__118 (.L_HI(net118));
 sg13g2_tiehi _6266__119 (.L_HI(net119));
 sg13g2_tiehi _6265__120 (.L_HI(net120));
 sg13g2_tiehi _6264__121 (.L_HI(net121));
 sg13g2_tiehi _6263__122 (.L_HI(net122));
 sg13g2_tiehi _6262__123 (.L_HI(net123));
 sg13g2_tiehi _6261__124 (.L_HI(net124));
 sg13g2_tiehi _6260__125 (.L_HI(net125));
 sg13g2_tiehi _6259__126 (.L_HI(net126));
 sg13g2_tiehi _6258__127 (.L_HI(net127));
 sg13g2_tiehi _6257__128 (.L_HI(net128));
 sg13g2_tiehi _6256__129 (.L_HI(net129));
 sg13g2_tiehi _6255__130 (.L_HI(net130));
 sg13g2_tiehi _6254__131 (.L_HI(net131));
 sg13g2_tiehi _6253__132 (.L_HI(net132));
 sg13g2_tiehi _6252__133 (.L_HI(net133));
 sg13g2_tiehi _6251__134 (.L_HI(net134));
 sg13g2_tiehi _6250__135 (.L_HI(net135));
 sg13g2_tiehi _6249__136 (.L_HI(net136));
 sg13g2_tiehi _6248__137 (.L_HI(net137));
 sg13g2_tiehi _6247__138 (.L_HI(net138));
 sg13g2_tiehi _6246__139 (.L_HI(net139));
 sg13g2_tiehi _6245__140 (.L_HI(net140));
 sg13g2_tiehi _6244__141 (.L_HI(net141));
 sg13g2_tiehi _6243__142 (.L_HI(net142));
 sg13g2_tiehi _6242__143 (.L_HI(net143));
 sg13g2_tiehi _6241__144 (.L_HI(net144));
 sg13g2_tiehi _6240__145 (.L_HI(net145));
 sg13g2_tiehi _6239__146 (.L_HI(net146));
 sg13g2_tiehi _6238__147 (.L_HI(net147));
 sg13g2_tiehi _6237__148 (.L_HI(net148));
 sg13g2_tiehi _6236__149 (.L_HI(net149));
 sg13g2_tiehi _6235__150 (.L_HI(net150));
 sg13g2_tiehi _6234__151 (.L_HI(net151));
 sg13g2_tiehi _6233__152 (.L_HI(net152));
 sg13g2_tiehi _6232__153 (.L_HI(net153));
 sg13g2_tiehi _6231__154 (.L_HI(net154));
 sg13g2_tiehi _6230__155 (.L_HI(net155));
 sg13g2_tiehi _6229__156 (.L_HI(net156));
 sg13g2_tiehi _6228__157 (.L_HI(net157));
 sg13g2_tiehi _6146__158 (.L_HI(net158));
 sg13g2_tiehi _6293__159 (.L_HI(net159));
 sg13g2_tiehi _6227__160 (.L_HI(net160));
 sg13g2_tiehi _6226__161 (.L_HI(net161));
 sg13g2_tiehi _6225__162 (.L_HI(net162));
 sg13g2_tiehi _6224__163 (.L_HI(net163));
 sg13g2_tiehi _6223__164 (.L_HI(net164));
 sg13g2_tiehi _6222__165 (.L_HI(net165));
 sg13g2_tiehi _6221__166 (.L_HI(net166));
 sg13g2_tiehi _6220__167 (.L_HI(net167));
 sg13g2_tiehi _6219__168 (.L_HI(net168));
 sg13g2_tiehi _6218__169 (.L_HI(net169));
 sg13g2_tiehi _6307__170 (.L_HI(net170));
 sg13g2_tiehi _6308__171 (.L_HI(net171));
 sg13g2_tiehi _6309__172 (.L_HI(net172));
 sg13g2_tiehi _6310__173 (.L_HI(net173));
 sg13g2_tiehi _6311__174 (.L_HI(net174));
 sg13g2_tiehi _6312__175 (.L_HI(net175));
 sg13g2_tiehi _6313__176 (.L_HI(net176));
 sg13g2_tiehi _6314__177 (.L_HI(net177));
 sg13g2_tiehi _6315__178 (.L_HI(net178));
 sg13g2_tiehi _6217__179 (.L_HI(net179));
 sg13g2_tiehi _6216__180 (.L_HI(net180));
 sg13g2_tiehi _6215__181 (.L_HI(net181));
 sg13g2_tiehi _6214__182 (.L_HI(net182));
 sg13g2_tiehi _6213__183 (.L_HI(net183));
 sg13g2_tiehi _6212__184 (.L_HI(net184));
 sg13g2_tiehi _6211__185 (.L_HI(net185));
 sg13g2_tiehi _6210__186 (.L_HI(net186));
 sg13g2_tiehi _6209__187 (.L_HI(net187));
 sg13g2_tiehi _6208__188 (.L_HI(net188));
 sg13g2_tiehi _6207__189 (.L_HI(net189));
 sg13g2_tiehi _6206__190 (.L_HI(net190));
 sg13g2_tiehi _6205__191 (.L_HI(net191));
 sg13g2_tiehi _6204__192 (.L_HI(net192));
 sg13g2_tiehi _6203__193 (.L_HI(net193));
 sg13g2_tiehi _6202__194 (.L_HI(net194));
 sg13g2_tiehi _6201__195 (.L_HI(net195));
 sg13g2_tiehi _6200__196 (.L_HI(net196));
 sg13g2_tiehi _6199__197 (.L_HI(net197));
 sg13g2_tiehi _6198__198 (.L_HI(net198));
 sg13g2_tiehi _6197__199 (.L_HI(net199));
 sg13g2_tiehi _6196__200 (.L_HI(net200));
 sg13g2_tiehi _6195__201 (.L_HI(net201));
 sg13g2_tiehi _6194__202 (.L_HI(net202));
 sg13g2_tiehi _6193__203 (.L_HI(net203));
 sg13g2_tiehi _6192__204 (.L_HI(net204));
 sg13g2_tiehi _6191__205 (.L_HI(net205));
 sg13g2_tiehi _6190__206 (.L_HI(net206));
 sg13g2_tiehi _6189__207 (.L_HI(net207));
 sg13g2_tiehi _6188__208 (.L_HI(net208));
 sg13g2_tiehi _6187__209 (.L_HI(net209));
 sg13g2_tiehi _6186__210 (.L_HI(net210));
 sg13g2_tiehi _6185__211 (.L_HI(net211));
 sg13g2_tiehi _6184__212 (.L_HI(net212));
 sg13g2_tiehi _6183__213 (.L_HI(net213));
 sg13g2_tiehi _6182__214 (.L_HI(net214));
 sg13g2_tiehi _6181__215 (.L_HI(net215));
 sg13g2_tiehi _6180__216 (.L_HI(net216));
 sg13g2_tiehi _6316__217 (.L_HI(net217));
 sg13g2_tiehi _6355__218 (.L_HI(net218));
 sg13g2_tiehi _6356__219 (.L_HI(net219));
 sg13g2_tiehi _6179__220 (.L_HI(net220));
 sg13g2_tiehi _6178__221 (.L_HI(net221));
 sg13g2_tiehi _6177__222 (.L_HI(net222));
 sg13g2_tiehi _6176__223 (.L_HI(net223));
 sg13g2_tiehi _6175__224 (.L_HI(net224));
 sg13g2_tiehi _6174__225 (.L_HI(net225));
 sg13g2_tiehi _6173__226 (.L_HI(net226));
 sg13g2_tiehi _6172__227 (.L_HI(net227));
 sg13g2_tiehi _6171__228 (.L_HI(net228));
 sg13g2_tiehi _6170__229 (.L_HI(net229));
 sg13g2_tiehi _6169__230 (.L_HI(net230));
 sg13g2_tiehi _6168__231 (.L_HI(net231));
 sg13g2_tiehi _6167__232 (.L_HI(net232));
 sg13g2_tiehi _6166__233 (.L_HI(net233));
 sg13g2_tiehi _6165__234 (.L_HI(net234));
 sg13g2_tiehi _6164__235 (.L_HI(net235));
 sg13g2_tiehi _6163__236 (.L_HI(net236));
 sg13g2_tiehi _6162__237 (.L_HI(net237));
 sg13g2_tiehi _6161__238 (.L_HI(net238));
 sg13g2_tiehi _6160__239 (.L_HI(net239));
 sg13g2_tiehi _6159__240 (.L_HI(net240));
 sg13g2_tiehi _6158__241 (.L_HI(net241));
 sg13g2_tiehi _6157__242 (.L_HI(net242));
 sg13g2_tiehi _6156__243 (.L_HI(net243));
 sg13g2_tiehi _6155__244 (.L_HI(net244));
 sg13g2_tiehi _6154__245 (.L_HI(net245));
 sg13g2_tiehi _6153__246 (.L_HI(net246));
 sg13g2_tiehi _6551__247 (.L_HI(net247));
 sg13g2_tiehi _6152__248 (.L_HI(net248));
 sg13g2_tiehi _6643__249 (.L_HI(net249));
 sg13g2_tiehi _6151__250 (.L_HI(net250));
 sg13g2_tiehi _6550__251 (.L_HI(net251));
 sg13g2_tiehi _6150__252 (.L_HI(net252));
 sg13g2_tiehi _6689__253 (.L_HI(net253));
 sg13g2_tiehi _6149__254 (.L_HI(net254));
 sg13g2_tiehi _6549__255 (.L_HI(net255));
 sg13g2_tiehi _6148__256 (.L_HI(net256));
 sg13g2_tiehi _6642__257 (.L_HI(net257));
 sg13g2_tiehi _6147__258 (.L_HI(net258));
 sg13g2_tiehi _6548__259 (.L_HI(net259));
 sg13g2_tiehi _6725__260 (.L_HI(net260));
 sg13g2_tiehi _6547__261 (.L_HI(net261));
 sg13g2_tiehi _6641__262 (.L_HI(net262));
 sg13g2_tiehi _6546__263 (.L_HI(net263));
 sg13g2_tiehi _6688__264 (.L_HI(net264));
 sg13g2_tiehi _6545__265 (.L_HI(net265));
 sg13g2_tiehi _6640__266 (.L_HI(net266));
 sg13g2_tiehi _6544__267 (.L_HI(net267));
 sg13g2_tiehi _6724__268 (.L_HI(net268));
 sg13g2_tiehi _6543__269 (.L_HI(net269));
 sg13g2_tiehi _6639__270 (.L_HI(net270));
 sg13g2_tiehi _6542__271 (.L_HI(net271));
 sg13g2_tiehi _6687__272 (.L_HI(net272));
 sg13g2_tiehi _6541__273 (.L_HI(net273));
 sg13g2_tiehi _6638__274 (.L_HI(net274));
 sg13g2_tiehi _6540__275 (.L_HI(net275));
 sg13g2_tiehi _6723__276 (.L_HI(net276));
 sg13g2_tiehi _6539__277 (.L_HI(net277));
 sg13g2_tiehi _6637__278 (.L_HI(net278));
 sg13g2_tiehi _6538__279 (.L_HI(net279));
 sg13g2_tiehi _6686__280 (.L_HI(net280));
 sg13g2_tiehi _6537__281 (.L_HI(net281));
 sg13g2_tiehi _6636__282 (.L_HI(net282));
 sg13g2_tiehi _6536__283 (.L_HI(net283));
 sg13g2_tiehi _6722__284 (.L_HI(net284));
 sg13g2_tiehi _6535__285 (.L_HI(net285));
 sg13g2_tiehi _6635__286 (.L_HI(net286));
 sg13g2_tiehi _6534__287 (.L_HI(net287));
 sg13g2_tiehi _6685__288 (.L_HI(net288));
 sg13g2_tiehi _6533__289 (.L_HI(net289));
 sg13g2_tiehi _6634__290 (.L_HI(net290));
 sg13g2_tiehi _6532__291 (.L_HI(net291));
 sg13g2_tiehi _6721__292 (.L_HI(net292));
 sg13g2_tiehi _6531__293 (.L_HI(net293));
 sg13g2_tiehi _6633__294 (.L_HI(net294));
 sg13g2_tiehi _6530__295 (.L_HI(net295));
 sg13g2_tiehi _6684__296 (.L_HI(net296));
 sg13g2_tiehi _6529__297 (.L_HI(net297));
 sg13g2_tiehi _6632__298 (.L_HI(net298));
 sg13g2_tiehi _6528__299 (.L_HI(net299));
 sg13g2_tiehi _6720__300 (.L_HI(net300));
 sg13g2_tiehi _6527__301 (.L_HI(net301));
 sg13g2_tiehi _6631__302 (.L_HI(net302));
 sg13g2_tiehi _6526__303 (.L_HI(net303));
 sg13g2_tiehi _6683__304 (.L_HI(net304));
 sg13g2_tiehi _6525__305 (.L_HI(net305));
 sg13g2_tiehi _6630__306 (.L_HI(net306));
 sg13g2_tiehi _6524__307 (.L_HI(net307));
 sg13g2_tiehi _6719__308 (.L_HI(net308));
 sg13g2_tiehi _6523__309 (.L_HI(net309));
 sg13g2_tiehi _6629__310 (.L_HI(net310));
 sg13g2_tiehi _6522__311 (.L_HI(net311));
 sg13g2_tiehi _6682__312 (.L_HI(net312));
 sg13g2_tiehi _6521__313 (.L_HI(net313));
 sg13g2_tiehi _6628__314 (.L_HI(net314));
 sg13g2_tiehi _6520__315 (.L_HI(net315));
 sg13g2_tiehi _6718__316 (.L_HI(net316));
 sg13g2_tiehi _6519__317 (.L_HI(net317));
 sg13g2_tiehi _6627__318 (.L_HI(net318));
 sg13g2_tiehi _6357__319 (.L_HI(net319));
 sg13g2_tiehi _6457__320 (.L_HI(net320));
 sg13g2_tiehi _6458__321 (.L_HI(net321));
 sg13g2_tiehi _6459__322 (.L_HI(net322));
 sg13g2_tiehi _6460__323 (.L_HI(net323));
 sg13g2_tiehi _6461__324 (.L_HI(net324));
 sg13g2_tiehi _6462__325 (.L_HI(net325));
 sg13g2_tiehi _6463__326 (.L_HI(net326));
 sg13g2_tiehi _6464__327 (.L_HI(net327));
 sg13g2_tiehi _6465__328 (.L_HI(net328));
 sg13g2_tiehi _6466__329 (.L_HI(net329));
 sg13g2_tiehi _6467__330 (.L_HI(net330));
 sg13g2_tiehi _6468__331 (.L_HI(net331));
 sg13g2_tiehi _6518__332 (.L_HI(net332));
 sg13g2_tiehi _6517__333 (.L_HI(net333));
 sg13g2_tiehi _6513__334 (.L_HI(net334));
 sg13g2_tiehi _6681__335 (.L_HI(net335));
 sg13g2_tiehi _6512__336 (.L_HI(net336));
 sg13g2_tiehi _6626__337 (.L_HI(net337));
 sg13g2_tiehi _6511__338 (.L_HI(net338));
 sg13g2_tiehi _6717__339 (.L_HI(net339));
 sg13g2_tiehi _6507__340 (.L_HI(net340));
 sg13g2_tiehi _6625__341 (.L_HI(net341));
 sg13g2_tiehi _6506__342 (.L_HI(net342));
 sg13g2_tiehi _6680__343 (.L_HI(net343));
 sg13g2_tiehi _6505__344 (.L_HI(net344));
 sg13g2_tiehi _6624__345 (.L_HI(net345));
 sg13g2_tiehi _6469__346 (.L_HI(net346));
 sg13g2_tiehi _6484__347 (.L_HI(net347));
 sg13g2_tiehi _6485__348 (.L_HI(net348));
 sg13g2_tiehi _6486__349 (.L_HI(net349));
 sg13g2_tiehi _6487__350 (.L_HI(net350));
 sg13g2_tiehi _6488__351 (.L_HI(net351));
 sg13g2_tiehi _6504__352 (.L_HI(net352));
 sg13g2_tiehi _6716__353 (.L_HI(net353));
 sg13g2_tiehi _6489__354 (.L_HI(net354));
 sg13g2_tiehi _6492__355 (.L_HI(net355));
 sg13g2_tiehi _6493__356 (.L_HI(net356));
 sg13g2_tiehi _6494__357 (.L_HI(net357));
 sg13g2_tiehi _6495__358 (.L_HI(net358));
 sg13g2_tiehi _6496__359 (.L_HI(net359));
 sg13g2_tiehi _6497__360 (.L_HI(net360));
 sg13g2_tiehi _6498__361 (.L_HI(net361));
 sg13g2_tiehi _6499__362 (.L_HI(net362));
 sg13g2_tiehi _6500__363 (.L_HI(net363));
 sg13g2_tiehi _6503__364 (.L_HI(net364));
 sg13g2_tiehi _6502__365 (.L_HI(net365));
 sg13g2_tiehi _6491__366 (.L_HI(net366));
 sg13g2_tiehi _6490__367 (.L_HI(net367));
 sg13g2_tiehi _6483__368 (.L_HI(net368));
 sg13g2_tiehi _6482__369 (.L_HI(net369));
 sg13g2_tiehi _6501__370 (.L_HI(net370));
 sg13g2_tiehi _6508__371 (.L_HI(net371));
 sg13g2_tiehi _6509__372 (.L_HI(net372));
 sg13g2_tiehi _6623__373 (.L_HI(net373));
 sg13g2_tiehi _6481__374 (.L_HI(net374));
 sg13g2_tiehi _6679__375 (.L_HI(net375));
 sg13g2_tiehi _6510__376 (.L_HI(net376));
 sg13g2_tiehi _6514__377 (.L_HI(net377));
 sg13g2_tiehi _6515__378 (.L_HI(net378));
 sg13g2_tiehi _6480__379 (.L_HI(net379));
 sg13g2_tiehi _6622__380 (.L_HI(net380));
 sg13g2_tiehi _6479__381 (.L_HI(net381));
 sg13g2_tiehi _6715__382 (.L_HI(net382));
 sg13g2_tiehi _6478__383 (.L_HI(net383));
 sg13g2_tiehi _6621__384 (.L_HI(net384));
 sg13g2_tiehi _6477__385 (.L_HI(net385));
 sg13g2_tiehi _6678__386 (.L_HI(net386));
 sg13g2_tiehi _6476__387 (.L_HI(net387));
 sg13g2_tiehi _6620__388 (.L_HI(net388));
 sg13g2_tiehi _6475__389 (.L_HI(net389));
 sg13g2_tiehi _6714__390 (.L_HI(net390));
 sg13g2_tiehi _6474__391 (.L_HI(net391));
 sg13g2_tiehi _6619__392 (.L_HI(net392));
 sg13g2_tiehi _6473__393 (.L_HI(net393));
 sg13g2_tiehi _6677__394 (.L_HI(net394));
 sg13g2_tiehi _6472__395 (.L_HI(net395));
 sg13g2_tiehi _6618__396 (.L_HI(net396));
 sg13g2_tiehi _6471__397 (.L_HI(net397));
 sg13g2_tiehi _6470__398 (.L_HI(net398));
 sg13g2_tiehi _6456__399 (.L_HI(net399));
 sg13g2_tiehi _6713__400 (.L_HI(net400));
 sg13g2_tiehi _6455__401 (.L_HI(net401));
 sg13g2_tiehi _6617__402 (.L_HI(net402));
 sg13g2_tiehi _6454__403 (.L_HI(net403));
 sg13g2_tiehi _6676__404 (.L_HI(net404));
 sg13g2_tiehi _6453__405 (.L_HI(net405));
 sg13g2_tiehi _6616__406 (.L_HI(net406));
 sg13g2_tiehi _6452__407 (.L_HI(net407));
 sg13g2_tiehi _6712__408 (.L_HI(net408));
 sg13g2_tiehi _6451__409 (.L_HI(net409));
 sg13g2_tiehi _6615__410 (.L_HI(net410));
 sg13g2_tiehi _6450__411 (.L_HI(net411));
 sg13g2_tiehi _6675__412 (.L_HI(net412));
 sg13g2_tiehi _6449__413 (.L_HI(net413));
 sg13g2_tiehi _6614__414 (.L_HI(net414));
 sg13g2_tiehi _6448__415 (.L_HI(net415));
 sg13g2_tiehi _6711__416 (.L_HI(net416));
 sg13g2_tiehi _6447__417 (.L_HI(net417));
 sg13g2_tiehi _6613__418 (.L_HI(net418));
 sg13g2_tiehi _6446__419 (.L_HI(net419));
 sg13g2_tiehi _6674__420 (.L_HI(net420));
 sg13g2_tiehi _6445__421 (.L_HI(net421));
 sg13g2_tiehi _6612__422 (.L_HI(net422));
 sg13g2_tiehi _6444__423 (.L_HI(net423));
 sg13g2_tiehi _6710__424 (.L_HI(net424));
 sg13g2_tiehi _6443__425 (.L_HI(net425));
 sg13g2_tiehi _6611__426 (.L_HI(net426));
 sg13g2_tiehi _6442__427 (.L_HI(net427));
 sg13g2_tiehi _6673__428 (.L_HI(net428));
 sg13g2_tiehi _6441__429 (.L_HI(net429));
 sg13g2_tiehi _6610__430 (.L_HI(net430));
 sg13g2_tiehi _6440__431 (.L_HI(net431));
 sg13g2_tiehi _6709__432 (.L_HI(net432));
 sg13g2_tiehi _6439__433 (.L_HI(net433));
 sg13g2_tiehi _6609__434 (.L_HI(net434));
 sg13g2_tiehi _6438__435 (.L_HI(net435));
 sg13g2_tiehi _6672__436 (.L_HI(net436));
 sg13g2_tiehi _6437__437 (.L_HI(net437));
 sg13g2_tiehi _6608__438 (.L_HI(net438));
 sg13g2_tiehi _6436__439 (.L_HI(net439));
 sg13g2_tiehi _6708__440 (.L_HI(net440));
 sg13g2_tiehi _6435__441 (.L_HI(net441));
 sg13g2_tiehi _6607__442 (.L_HI(net442));
 sg13g2_tiehi _6434__443 (.L_HI(net443));
 sg13g2_tiehi _6671__444 (.L_HI(net444));
 sg13g2_tiehi _6433__445 (.L_HI(net445));
 sg13g2_tiehi _6606__446 (.L_HI(net446));
 sg13g2_tiehi _6432__447 (.L_HI(net447));
 sg13g2_tiehi _6707__448 (.L_HI(net448));
 sg13g2_tiehi _6431__449 (.L_HI(net449));
 sg13g2_tiehi _6605__450 (.L_HI(net450));
 sg13g2_tiehi _6430__451 (.L_HI(net451));
 sg13g2_tiehi _6670__452 (.L_HI(net452));
 sg13g2_tiehi _6429__453 (.L_HI(net453));
 sg13g2_tiehi _6604__454 (.L_HI(net454));
 sg13g2_tiehi _6428__455 (.L_HI(net455));
 sg13g2_tiehi _6706__456 (.L_HI(net456));
 sg13g2_tiehi _6427__457 (.L_HI(net457));
 sg13g2_tiehi _6603__458 (.L_HI(net458));
 sg13g2_tiehi _6426__459 (.L_HI(net459));
 sg13g2_tiehi _6669__460 (.L_HI(net460));
 sg13g2_tiehi _6425__461 (.L_HI(net461));
 sg13g2_tiehi _6602__462 (.L_HI(net462));
 sg13g2_tiehi _6424__463 (.L_HI(net463));
 sg13g2_tiehi _6705__464 (.L_HI(net464));
 sg13g2_tiehi _6423__465 (.L_HI(net465));
 sg13g2_tiehi _6601__466 (.L_HI(net466));
 sg13g2_tiehi _6422__467 (.L_HI(net467));
 sg13g2_tiehi _6668__468 (.L_HI(net468));
 sg13g2_tiehi _6421__469 (.L_HI(net469));
 sg13g2_tiehi _6600__470 (.L_HI(net470));
 sg13g2_tiehi _6420__471 (.L_HI(net471));
 sg13g2_tiehi _6704__472 (.L_HI(net472));
 sg13g2_tiehi _6419__473 (.L_HI(net473));
 sg13g2_tiehi _6599__474 (.L_HI(net474));
 sg13g2_tiehi _6418__475 (.L_HI(net475));
 sg13g2_tiehi _6667__476 (.L_HI(net476));
 sg13g2_tiehi _6417__477 (.L_HI(net477));
 sg13g2_tiehi _6598__478 (.L_HI(net478));
 sg13g2_tiehi _6416__479 (.L_HI(net479));
 sg13g2_tiehi _6703__480 (.L_HI(net480));
 sg13g2_tiehi _6415__481 (.L_HI(net481));
 sg13g2_tiehi _6597__482 (.L_HI(net482));
 sg13g2_tiehi _6414__483 (.L_HI(net483));
 sg13g2_tiehi _6666__484 (.L_HI(net484));
 sg13g2_tiehi _6413__485 (.L_HI(net485));
 sg13g2_tiehi _6596__486 (.L_HI(net486));
 sg13g2_tiehi _6412__487 (.L_HI(net487));
 sg13g2_tiehi _6702__488 (.L_HI(net488));
 sg13g2_tiehi _6411__489 (.L_HI(net489));
 sg13g2_tiehi _6595__490 (.L_HI(net490));
 sg13g2_tiehi _6410__491 (.L_HI(net491));
 sg13g2_tiehi _6665__492 (.L_HI(net492));
 sg13g2_tiehi _6409__493 (.L_HI(net493));
 sg13g2_tiehi _6594__494 (.L_HI(net494));
 sg13g2_tiehi _6408__495 (.L_HI(net495));
 sg13g2_tiehi _6701__496 (.L_HI(net496));
 sg13g2_tiehi _6407__497 (.L_HI(net497));
 sg13g2_tiehi _6593__498 (.L_HI(net498));
 sg13g2_tiehi _6406__499 (.L_HI(net499));
 sg13g2_tiehi _6664__500 (.L_HI(net500));
 sg13g2_tiehi _6405__501 (.L_HI(net501));
 sg13g2_tiehi _6592__502 (.L_HI(net502));
 sg13g2_tiehi _6404__503 (.L_HI(net503));
 sg13g2_tiehi _6740__504 (.L_HI(net504));
 sg13g2_tiehi _6403__505 (.L_HI(net505));
 sg13g2_tiehi _6591__506 (.L_HI(net506));
 sg13g2_tiehi _6402__507 (.L_HI(net507));
 sg13g2_tiehi _6663__508 (.L_HI(net508));
 sg13g2_tiehi _6401__509 (.L_HI(net509));
 sg13g2_tiehi _6590__510 (.L_HI(net510));
 sg13g2_tiehi _6400__511 (.L_HI(net511));
 sg13g2_tiehi _6700__512 (.L_HI(net512));
 sg13g2_tiehi _6399__513 (.L_HI(net513));
 sg13g2_tiehi _6589__514 (.L_HI(net514));
 sg13g2_tiehi _6398__515 (.L_HI(net515));
 sg13g2_tiehi _6662__516 (.L_HI(net516));
 sg13g2_tiehi _6397__517 (.L_HI(net517));
 sg13g2_tiehi _6588__518 (.L_HI(net518));
 sg13g2_tiehi _6396__519 (.L_HI(net519));
 sg13g2_tiehi _6731__520 (.L_HI(net520));
 sg13g2_tiehi _6395__521 (.L_HI(net521));
 sg13g2_tiehi _6587__522 (.L_HI(net522));
 sg13g2_tiehi _6394__523 (.L_HI(net523));
 sg13g2_tiehi _6661__524 (.L_HI(net524));
 sg13g2_tiehi _6393__525 (.L_HI(net525));
 sg13g2_tiehi _6586__526 (.L_HI(net526));
 sg13g2_tiehi _6392__527 (.L_HI(net527));
 sg13g2_tiehi _6699__528 (.L_HI(net528));
 sg13g2_tiehi _6391__529 (.L_HI(net529));
 sg13g2_tiehi _6585__530 (.L_HI(net530));
 sg13g2_tiehi _6390__531 (.L_HI(net531));
 sg13g2_tiehi _6660__532 (.L_HI(net532));
 sg13g2_tiehi _6389__533 (.L_HI(net533));
 sg13g2_tiehi _6584__534 (.L_HI(net534));
 sg13g2_tiehi _6388__535 (.L_HI(net535));
 sg13g2_tiehi _6733__536 (.L_HI(net536));
 sg13g2_tiehi _6387__537 (.L_HI(net537));
 sg13g2_tiehi _6583__538 (.L_HI(net538));
 sg13g2_tiehi _6386__539 (.L_HI(net539));
 sg13g2_tiehi _6659__540 (.L_HI(net540));
 sg13g2_tiehi _6385__541 (.L_HI(net541));
 sg13g2_tiehi _6582__542 (.L_HI(net542));
 sg13g2_tiehi _6384__543 (.L_HI(net543));
 sg13g2_tiehi _6698__544 (.L_HI(net544));
 sg13g2_tiehi _6383__545 (.L_HI(net545));
 sg13g2_tiehi _6581__546 (.L_HI(net546));
 sg13g2_tiehi _6382__547 (.L_HI(net547));
 sg13g2_tiehi _6658__548 (.L_HI(net548));
 sg13g2_tiehi _6381__549 (.L_HI(net549));
 sg13g2_tiehi _6580__550 (.L_HI(net550));
 sg13g2_tiehi _6380__551 (.L_HI(net551));
 sg13g2_tiehi _6730__552 (.L_HI(net552));
 sg13g2_tiehi _6379__553 (.L_HI(net553));
 sg13g2_tiehi _6579__554 (.L_HI(net554));
 sg13g2_tiehi _6378__555 (.L_HI(net555));
 sg13g2_tiehi _6657__556 (.L_HI(net556));
 sg13g2_tiehi _6377__557 (.L_HI(net557));
 sg13g2_tiehi _6578__558 (.L_HI(net558));
 sg13g2_tiehi _6376__559 (.L_HI(net559));
 sg13g2_tiehi _6697__560 (.L_HI(net560));
 sg13g2_tiehi _6375__561 (.L_HI(net561));
 sg13g2_tiehi _6577__562 (.L_HI(net562));
 sg13g2_tiehi _6374__563 (.L_HI(net563));
 sg13g2_tiehi _6656__564 (.L_HI(net564));
 sg13g2_tiehi _6373__565 (.L_HI(net565));
 sg13g2_tiehi _6576__566 (.L_HI(net566));
 sg13g2_tiehi _6372__567 (.L_HI(net567));
 sg13g2_tiehi _6741__568 (.L_HI(net568));
 sg13g2_tiehi _6371__569 (.L_HI(net569));
 sg13g2_tiehi _6575__570 (.L_HI(net570));
 sg13g2_tiehi _6370__571 (.L_HI(net571));
 sg13g2_tiehi _6655__572 (.L_HI(net572));
 sg13g2_tiehi _6369__573 (.L_HI(net573));
 sg13g2_tiehi _6574__574 (.L_HI(net574));
 sg13g2_tiehi _6368__575 (.L_HI(net575));
 sg13g2_tiehi _6696__576 (.L_HI(net576));
 sg13g2_tiehi _6367__577 (.L_HI(net577));
 sg13g2_tiehi _6573__578 (.L_HI(net578));
 sg13g2_tiehi _6366__579 (.L_HI(net579));
 sg13g2_tiehi _6654__580 (.L_HI(net580));
 sg13g2_tiehi _6365__581 (.L_HI(net581));
 sg13g2_tiehi _6572__582 (.L_HI(net582));
 sg13g2_tiehi _6364__583 (.L_HI(net583));
 sg13g2_tiehi _6729__584 (.L_HI(net584));
 sg13g2_tiehi _6363__585 (.L_HI(net585));
 sg13g2_tiehi _6571__586 (.L_HI(net586));
 sg13g2_tiehi _6362__587 (.L_HI(net587));
 sg13g2_tiehi _6653__588 (.L_HI(net588));
 sg13g2_tiehi _6361__589 (.L_HI(net589));
 sg13g2_tiehi _6360__590 (.L_HI(net590));
 sg13g2_tiehi _6359__591 (.L_HI(net591));
 sg13g2_tiehi _6570__592 (.L_HI(net592));
 sg13g2_tiehi _6358__593 (.L_HI(net593));
 sg13g2_tiehi _6695__594 (.L_HI(net594));
 sg13g2_tiehi _6354__595 (.L_HI(net595));
 sg13g2_tiehi _6516__596 (.L_HI(net596));
 sg13g2_tiehi _6734__597 (.L_HI(net597));
 sg13g2_tiehi _6735__598 (.L_HI(net598));
 sg13g2_tiehi _6736__599 (.L_HI(net599));
 sg13g2_tiehi _6737__600 (.L_HI(net600));
 sg13g2_tiehi _6738__601 (.L_HI(net601));
 sg13g2_tiehi _6739__602 (.L_HI(net602));
 sg13g2_tiehi tt_um_devinatkin_basys3_uart_603 (.L_HI(net603));
 sg13g2_tiehi tt_um_devinatkin_basys3_uart_604 (.L_HI(net604));
 sg13g2_tiehi tt_um_devinatkin_basys3_uart_605 (.L_HI(net605));
 sg13g2_tiehi tt_um_devinatkin_basys3_uart_606 (.L_HI(net606));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_devinatkin_basys3_uart_4 (.L_LO(net4));
 sg13g2_tielo tt_um_devinatkin_basys3_uart_5 (.L_LO(net5));
 sg13g2_tielo tt_um_devinatkin_basys3_uart_6 (.L_LO(net6));
 sg13g2_tielo tt_um_devinatkin_basys3_uart_7 (.L_LO(net7));
 sg13g2_tielo tt_um_devinatkin_basys3_uart_8 (.L_LO(net8));
 sg13g2_tielo tt_um_devinatkin_basys3_uart_9 (.L_LO(net9));
 sg13g2_tielo tt_um_devinatkin_basys3_uart_10 (.L_LO(net10));
 sg13g2_tiehi _6569__11 (.L_HI(net11));
 sg13g2_buf_1 _7346_ (.A(tx_signal),
    .X(uio_out[0]));
 sg13g2_buf_2 _7347_ (.A(net889),
    .X(uio_out[2]));
 sg13g2_buf_2 _7348_ (.A(tx_valid),
    .X(uio_out[3]));
 sg13g2_buf_1 _7349_ (.A(rx_valid),
    .X(uio_out[5]));
 sg13g2_buf_2 fanout725 (.A(net726),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(net729),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(net729),
    .X(net727));
 sg13g2_buf_1 fanout728 (.A(net729),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(_1837_),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(net733),
    .X(net730));
 sg13g2_buf_1 fanout731 (.A(net733),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(net733),
    .X(net732));
 sg13g2_buf_1 fanout733 (.A(_1288_),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(net735),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(_1288_),
    .X(net735));
 sg13g2_buf_4 fanout736 (.X(net736),
    .A(net738));
 sg13g2_buf_2 fanout737 (.A(net738),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_2195_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(_1418_),
    .X(net739));
 sg13g2_buf_1 fanout740 (.A(_1418_),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(net743),
    .X(net741));
 sg13g2_buf_1 fanout742 (.A(net743),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(_1413_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(net754),
    .X(net744));
 sg13g2_buf_1 fanout745 (.A(net754),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(net747),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(net754),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(net754),
    .X(net748));
 sg13g2_buf_1 fanout749 (.A(net750),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(net754),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(net753),
    .X(net751));
 sg13g2_buf_1 fanout752 (.A(net753),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(net754),
    .X(net753));
 sg13g2_buf_4 fanout754 (.X(net754),
    .A(_1399_));
 sg13g2_buf_2 fanout755 (.A(_0603_),
    .X(net755));
 sg13g2_buf_4 fanout756 (.X(net756),
    .A(net758));
 sg13g2_buf_2 fanout757 (.A(net758),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(_2199_),
    .X(net758));
 sg13g2_buf_4 fanout759 (.X(net759),
    .A(net761));
 sg13g2_buf_2 fanout760 (.A(net761),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_2186_),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(net764),
    .X(net762));
 sg13g2_buf_1 fanout763 (.A(net764),
    .X(net763));
 sg13g2_buf_1 fanout764 (.A(_2093_),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(_1999_),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(net768),
    .X(net766));
 sg13g2_buf_1 fanout767 (.A(net768),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(_1973_),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(net770),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(_1408_),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(net781),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(net781),
    .X(net772));
 sg13g2_buf_4 fanout773 (.X(net773),
    .A(net774));
 sg13g2_buf_4 fanout774 (.X(net774),
    .A(net781));
 sg13g2_buf_4 fanout775 (.X(net775),
    .A(net781));
 sg13g2_buf_1 fanout776 (.A(net777),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(net781),
    .X(net777));
 sg13g2_buf_4 fanout778 (.X(net778),
    .A(net780));
 sg13g2_buf_2 fanout779 (.A(net780),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(net781),
    .X(net780));
 sg13g2_buf_4 fanout781 (.X(net781),
    .A(_1400_));
 sg13g2_buf_2 fanout782 (.A(net783),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_1029_),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(_2330_),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(net787),
    .X(net785));
 sg13g2_buf_1 fanout786 (.A(net787),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(_1963_),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(net789),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(net791),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(net791),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(_1094_),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(net794),
    .X(net792));
 sg13g2_buf_2 fanout793 (.A(net794),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(_1094_),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(_1028_),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(net797),
    .X(net796));
 sg13g2_buf_1 fanout797 (.A(net798),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(_1028_),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(_2514_),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(net802),
    .X(net800));
 sg13g2_buf_1 fanout801 (.A(net802),
    .X(net801));
 sg13g2_buf_2 fanout802 (.A(_2216_),
    .X(net802));
 sg13g2_buf_2 fanout803 (.A(net804),
    .X(net803));
 sg13g2_buf_2 fanout804 (.A(net807),
    .X(net804));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(net806));
 sg13g2_buf_2 fanout806 (.A(net807),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(_2216_),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(_0996_),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(net813),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(net813),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(net812),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(net813),
    .X(net812));
 sg13g2_buf_1 fanout813 (.A(_2215_),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(net815),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(net819),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(net818),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(net818),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(net819),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(_2215_),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(net822),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(net822),
    .X(net821));
 sg13g2_buf_1 fanout822 (.A(net823),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(net824),
    .X(net823));
 sg13g2_buf_4 fanout824 (.X(net824),
    .A(_2214_));
 sg13g2_buf_2 fanout825 (.A(_2180_),
    .X(net825));
 sg13g2_buf_4 fanout826 (.X(net826),
    .A(_0899_));
 sg13g2_buf_2 fanout827 (.A(net828),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(\SegmentDisplay.out_sel[1] ),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(net830),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(\SegmentDisplay.out_sel[2] ),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(_0167_),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(net833),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(\Led_Cycle_inst.csr.read_ptr[3] ),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(_0097_),
    .X(net834));
 sg13g2_buf_1 fanout835 (.A(_0097_),
    .X(net835));
 sg13g2_buf_4 fanout836 (.X(net836),
    .A(net837));
 sg13g2_buf_2 fanout837 (.A(\Led_Cycle_inst.csr.read_ptr[2] ),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(net839),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(\Led_Cycle_inst.csr.read_ptr[1] ),
    .X(net839));
 sg13g2_buf_4 fanout840 (.X(net840),
    .A(net841));
 sg13g2_buf_2 fanout841 (.A(\Led_Cycle_inst.csr.read_ptr[0] ),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(net843),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(_2437_),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(net846),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(net846),
    .X(net845));
 sg13g2_buf_1 fanout846 (.A(net853),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(net853),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(net853),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(net852),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(net852),
    .X(net850));
 sg13g2_buf_1 fanout851 (.A(net852),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(net853),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_2096_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(net855),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(net860),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(net859),
    .X(net856));
 sg13g2_buf_1 fanout857 (.A(net859),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(net859),
    .X(net858));
 sg13g2_buf_1 fanout859 (.A(net860),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_2095_),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(net863),
    .X(net861));
 sg13g2_buf_1 fanout862 (.A(net863),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(net864),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(_2095_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(net866),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(net869),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(net869),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(net869),
    .X(net868));
 sg13g2_buf_4 fanout869 (.X(net869),
    .A(net870));
 sg13g2_buf_1 fanout870 (.A(_2095_),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(_2031_),
    .X(net871));
 sg13g2_buf_4 fanout872 (.X(net872),
    .A(_2027_));
 sg13g2_buf_2 fanout873 (.A(net876),
    .X(net873));
 sg13g2_buf_1 fanout874 (.A(net876),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(net876),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(_0795_),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(net878),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(_0793_),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(net880),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(net1204),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(net882),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(net884),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(net884),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(\output_value_inst.ready_to_send ),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(net888),
    .X(net885));
 sg13g2_buf_1 fanout886 (.A(net888),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(net888),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(\output_value_inst.send_led_data ),
    .X(net888));
 sg13g2_buf_4 fanout889 (.X(net889),
    .A(net1222));
 sg13g2_buf_2 fanout890 (.A(net1173),
    .X(net890));
 sg13g2_buf_4 fanout891 (.X(net891),
    .A(net892));
 sg13g2_buf_4 fanout892 (.X(net892),
    .A(net899));
 sg13g2_buf_2 fanout893 (.A(net898),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(net898),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(net898),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(net897),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(net898),
    .X(net897));
 sg13g2_buf_4 fanout898 (.X(net898),
    .A(net899));
 sg13g2_buf_4 fanout899 (.X(net899),
    .A(_0900_));
 sg13g2_buf_4 fanout900 (.X(net900),
    .A(net912));
 sg13g2_buf_1 fanout901 (.A(net912),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(net904),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(net904),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(net912),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(net906),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(net907),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(net908),
    .X(net907));
 sg13g2_buf_4 fanout908 (.X(net908),
    .A(net912));
 sg13g2_buf_2 fanout909 (.A(net911),
    .X(net909));
 sg13g2_buf_1 fanout910 (.A(net911),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(net912),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(_0900_),
    .X(net912));
 sg13g2_buf_4 fanout913 (.X(net913),
    .A(_0794_));
 sg13g2_buf_4 fanout914 (.X(net914),
    .A(_0794_));
 sg13g2_buf_2 fanout915 (.A(net916),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(net917),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(net918),
    .X(net917));
 sg13g2_buf_4 fanout918 (.X(net918),
    .A(net924));
 sg13g2_buf_2 fanout919 (.A(net920),
    .X(net919));
 sg13g2_buf_4 fanout920 (.X(net920),
    .A(net924));
 sg13g2_buf_2 fanout921 (.A(net924),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(net923),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(net924),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(net961),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(net928),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(net928),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(net928),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(net937),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(net930),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(net937),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(net935),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(net935),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(net934),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(net935),
    .X(net934));
 sg13g2_buf_2 fanout935 (.A(net937),
    .X(net935));
 sg13g2_buf_4 fanout936 (.X(net936),
    .A(net937));
 sg13g2_buf_2 fanout937 (.A(net961),
    .X(net937));
 sg13g2_buf_4 fanout938 (.X(net938),
    .A(net942));
 sg13g2_buf_2 fanout939 (.A(net942),
    .X(net939));
 sg13g2_buf_4 fanout940 (.X(net940),
    .A(net941));
 sg13g2_buf_4 fanout941 (.X(net941),
    .A(net942));
 sg13g2_buf_2 fanout942 (.A(net961),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(net944),
    .X(net943));
 sg13g2_buf_4 fanout944 (.X(net944),
    .A(net947));
 sg13g2_buf_2 fanout945 (.A(net946),
    .X(net945));
 sg13g2_buf_4 fanout946 (.X(net946),
    .A(net947));
 sg13g2_buf_2 fanout947 (.A(net961),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(net950),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(net950),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(net961),
    .X(net950));
 sg13g2_buf_4 fanout951 (.X(net951),
    .A(net960));
 sg13g2_buf_2 fanout952 (.A(net953),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(net954),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(net960),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(net958),
    .X(net955));
 sg13g2_buf_1 fanout956 (.A(net958),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(net958),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(net959),
    .X(net958));
 sg13g2_buf_4 fanout959 (.X(net959),
    .A(net960));
 sg13g2_buf_2 fanout960 (.A(net961),
    .X(net960));
 sg13g2_buf_4 fanout961 (.X(net961),
    .A(rst_n));
 sg13g2_buf_4 fanout962 (.X(net962),
    .A(net963));
 sg13g2_buf_2 fanout963 (.A(net964),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(ena),
    .X(net964));
 sg13g2_buf_1 input1 (.A(uio_in[1]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(uio_in[4]),
    .X(net2));
 sg13g2_tielo tt_um_devinatkin_basys3_uart_3 (.L_LO(net3));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_72_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_75_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_2 clkbuf_leaf_76_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_2 clkbuf_leaf_77_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_2 clkbuf_leaf_78_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_2 clkbuf_leaf_79_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_2 clkbuf_leaf_80_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_2 clkbuf_leaf_81_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_4_4_0_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_4_5_0_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_4_6_0_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_buf_2 clkload7 (.A(clknet_4_9_0_clk));
 sg13g2_buf_2 clkload8 (.A(clknet_4_10_0_clk));
 sg13g2_buf_2 clkload9 (.A(clknet_4_11_0_clk));
 sg13g2_buf_2 clkload10 (.A(clknet_4_12_0_clk));
 sg13g2_buf_2 clkload11 (.A(clknet_4_13_0_clk));
 sg13g2_buf_1 clkload12 (.A(clknet_4_14_0_clk));
 sg13g2_buf_2 clkload13 (.A(clknet_4_15_0_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_1_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_81_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_2_clk));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_73_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_78_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_72_clk));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_20_clk));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_14_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_25_clk));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_27_clk));
 sg13g2_inv_4 clkload24 (.A(clknet_leaf_33_clk));
 sg13g2_inv_1 clkload25 (.A(clknet_leaf_66_clk));
 sg13g2_inv_1 clkload26 (.A(clknet_leaf_53_clk));
 sg13g2_inv_2 clkload27 (.A(clknet_leaf_54_clk));
 sg13g2_inv_2 clkload28 (.A(clknet_leaf_30_clk));
 sg13g2_inv_1 clkload29 (.A(clknet_leaf_31_clk));
 sg13g2_inv_4 clkload30 (.A(clknet_leaf_38_clk));
 sg13g2_inv_2 clkload31 (.A(clknet_leaf_43_clk));
 sg13g2_inv_4 clkload32 (.A(clknet_leaf_29_clk));
 sg13g2_inv_4 clkload33 (.A(clknet_leaf_40_clk));
 sg13g2_inv_1 clkload34 (.A(clknet_leaf_41_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\uart_tx_fifo_inst.fifo[3][0] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold2 (.A(_2273_),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold3 (.A(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[0] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold4 (.A(_1783_),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0332_),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold6 (.A(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[1] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0331_),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0217_),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0281_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0216_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0288_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0221_),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0253_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0211_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0323_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0214_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0302_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0223_),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0239_),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0166_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold21 (.A(_1777_),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0329_),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0186_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0294_),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0218_),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0274_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0207_),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0728_),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0199_),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0238_),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0209_),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0212_),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0316_),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0174_),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0301_),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0213_),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0309_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0206_),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0742_),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0197_),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold41 (.A(_1510_),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0245_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0178_),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0287_),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0224_),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0232_),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0201_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0336_),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0176_),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0280_),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0208_),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold52 (.A(_2028_),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0172_),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0308_),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0222_),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0246_),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0189_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0273_),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0195_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0252_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0219_),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0267_),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0215_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0295_),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0169_),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold66 (.A(_1748_),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0322_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0191_),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold69 (.A(_1572_),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0266_),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0183_),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold72 (.A(_1907_),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0369_),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold74 (.A(\uart_inst.uart_rx_inst.DATA_CNT[3] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0403_),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0192_),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold77 (.A(_1547_),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0259_),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0220_),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0260_),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0210_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold82 (.A(\output_value_inst.output_data[4] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0677_),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold84 (.A(\uart_tx_fifo_inst.fifo[2][5] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold85 (.A(_2271_),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold86 (.A(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[2] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold87 (.A(_1537_),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0255_),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold89 (.A(\uart_tx_fifo_inst.fifo[7][3] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold90 (.A(_1427_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold91 (.A(\uart_tx_fifo_inst.fifo[1][4] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold92 (.A(_2262_),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold93 (.A(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[2] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold94 (.A(_1655_),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0290_),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold96 (.A(\uart_tx_fifo_inst.fifo[1][3] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold97 (.A(_2261_),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0098_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0988_),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0989_),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold101 (.A(\output_value_inst.output_data[6] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0679_),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold103 (.A(\uart_inst.uart_rx_inst.DATA_TEMP_REG[0] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0392_),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold105 (.A(\SegmentDisplay.bcd2[0] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold106 (.A(_2323_),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold107 (.A(\output_value_inst.output_data[1] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0674_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold109 (.A(\output_value_inst.element_data_reg[6] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold110 (.A(\output_value_inst.output_data[3] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0676_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold112 (.A(\uart_tx_fifo_inst.fifo[6][0] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold113 (.A(_2299_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold114 (.A(\SegmentDisplay.bcd2[1] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold115 (.A(_2324_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold116 (.A(\output_value_inst.output_data[5] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0678_),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold118 (.A(\uart_tx_fifo_inst.fifo[6][6] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold119 (.A(_2306_),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold120 (.A(\uart_tx_fifo_inst.fifo[6][5] ),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold121 (.A(_2305_),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold122 (.A(\uart_tx_fifo_inst.fifo[6][4] ),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold123 (.A(_2304_),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold124 (.A(\output_value_inst.character_buff[4][6] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold125 (.A(_2404_),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold126 (.A(\output_value_inst.output_data[2] ),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0675_),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold128 (.A(\uart_tx_fifo_inst.fifo[1][6] ),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold129 (.A(_2264_),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold130 (.A(\SegmentDisplay.bcd3[0] ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0612_),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold132 (.A(\output_value_inst.element_data_reg[2] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold133 (.A(\rx_data[1] ),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0384_),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold135 (.A(_2627_),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold136 (.A(\SegmentDisplay.bcd3[1] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0613_),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold138 (.A(\output_value_inst.element_data_reg[3] ),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold139 (.A(\output_value_inst.character_buff[5][1] ),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold140 (.A(_2395_),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold141 (.A(\output_value_inst.character_buff[3][1] ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0653_),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold143 (.A(\input_value_check_inst.character_buff[0][1] ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold144 (.A(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[5] ),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0321_),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold146 (.A(\uart_tx_fifo_inst.fifo[0][1] ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold147 (.A(\uart_tx_fifo_inst.fifo[3][4] ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold148 (.A(_2280_),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold149 (.A(\rx_data[0] ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0383_),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold151 (.A(\input_value_check_inst.character_buff[0][0] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold152 (.A(\uart_tx_fifo_inst.fifo[4][2] ),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold153 (.A(_2286_),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold154 (.A(\output_value_inst.character_buff[3][6] ),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold155 (.A(_2411_),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold156 (.A(\rx_data[3] ),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0513_),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold158 (.A(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[5] ),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0251_),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold160 (.A(\uart_tx_fifo_inst.fifo[6][1] ),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold161 (.A(_2301_),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold162 (.A(\uart_tx_fifo_inst.fifo[4][1] ),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold163 (.A(_2285_),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold164 (.A(\uart_tx_fifo_inst.fifo[2][6] ),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold165 (.A(_2272_),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold166 (.A(\output_value_inst.character_buff[3][2] ),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold167 (.A(_2407_),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold168 (.A(\output_value_inst.element_data_reg[5] ),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0688_),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold170 (.A(\uart_tx_fifo_inst.fifo[2][3] ),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold171 (.A(_2269_),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold172 (.A(\uart_tx_fifo_inst.fifo[7][6] ),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold173 (.A(_1430_),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold174 (.A(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[5] ),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0293_),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold176 (.A(\rx_data[2] ),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0385_),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold178 (.A(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[5] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0335_),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold180 (.A(\output_value_inst.output_data[0] ),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0673_),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold182 (.A(\output_value_inst.element_data_reg[1] ),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold183 (.A(\rx_data[7] ),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0517_),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold185 (.A(\output_value_inst.character_buff[3][0] ),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold186 (.A(_2405_),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold187 (.A(\output_value_inst.element_data_reg[4] ),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold188 (.A(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[5] ),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0286_),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold190 (.A(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[5] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0272_),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold192 (.A(\uart_inst.uart_rx_inst.DATA_TEMP_REG[3] ),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold193 (.A(\uart_tx_fifo_inst.fifo[6][2] ),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold194 (.A(_2302_),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold195 (.A(\input_value_check_inst.character_buff[0][2] ),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold196 (.A(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[5] ),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0258_),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold198 (.A(\input_value_check_inst.character_buff[9][6] ),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0444_),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold200 (.A(\output_value_inst.character_buff[4][2] ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold201 (.A(\output_value_inst.send_element_data ),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold202 (.A(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[5] ),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0314_),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold204 (.A(\uart_tx_fifo_inst.fifo[2][1] ),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold205 (.A(_2267_),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold206 (.A(\uart_tx_fifo_inst.fifo[5][2] ),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold207 (.A(\output_value_inst.character_buff[5][0] ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold208 (.A(_2394_),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold209 (.A(\uart_tx_fifo_inst.fifo[3][5] ),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold210 (.A(_2281_),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold211 (.A(\uart_tx_fifo_inst.fifo[3][2] ),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold212 (.A(\uart_tx_fifo_inst.fifo[2][4] ),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold213 (.A(\uart_tx_fifo_inst.fifo[0][4] ),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold214 (.A(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[5] ),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0747_),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold216 (.A(\uart_tx_fifo_inst.fifo[1][2] ),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold217 (.A(_2260_),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold218 (.A(\output_value_inst.led_data_reg[7] ),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0702_),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold220 (.A(\rx_data[5] ),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0515_),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold222 (.A(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[5] ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0307_),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold224 (.A(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[5] ),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0328_),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold226 (.A(\uart_inst.uart_rx_inst.DATA_TEMP_REG[6] ),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0398_),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold228 (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[3] ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold229 (.A(_2518_),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0731_),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold231 (.A(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[5] ),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0244_),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold233 (.A(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[5] ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0300_),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold235 (.A(\output_value_inst.character_buff[3][4] ),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0656_),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold237 (.A(\rx_data[4] ),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0514_),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold239 (.A(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[5] ),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0265_),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold241 (.A(\uart_tx_fifo_inst.fifo[0][2] ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold242 (.A(\output_value_inst.led_data_reg[3] ),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0698_),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold244 (.A(\uart_tx_fifo_inst.fifo[4][0] ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold245 (.A(_2283_),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold246 (.A(\uart_inst.uart_rx_inst.DATA_TEMP_REG[5] ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold247 (.A(\uart_tx_fifo_inst.fifo[3][3] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold248 (.A(_2279_),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold249 (.A(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[5] ),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0237_),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold251 (.A(\uart_tx_fifo_inst.fifo[1][1] ),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold252 (.A(\uart_tx_fifo_inst.fifo[7][4] ),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold253 (.A(_1428_),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold254 (.A(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[5] ),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0279_),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold256 (.A(\uart_tx_fifo_inst.fifo[5][6] ),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold257 (.A(\uart_inst.uart_rx_inst.CLK_CNT[6] ),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold258 (.A(\uart_inst.uart_tx_inst.CLK_CNT[7] ),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold259 (.A(_2074_),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0433_),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold261 (.A(\uart_tx_fifo_inst.fifo[9][2] ),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold262 (.A(_2622_),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold263 (.A(\output_value_inst.led_data_reg[11] ),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0706_),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold265 (.A(\uart_inst.uart_rx_inst.DATA_TEMP_REG[7] ),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold266 (.A(\uart_tx_fifo_inst.fifo[7][1] ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold267 (.A(_1425_),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold268 (.A(\output_value_inst.character_buff[5][3] ),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold269 (.A(_2397_),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold270 (.A(\uart_tx_fifo_inst.fifo[5][3] ),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold271 (.A(_2295_),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold272 (.A(\uart_tx_fifo_inst.fifo[0][3] ),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold273 (.A(\uart_tx_fifo_inst.fifo[9][3] ),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold274 (.A(_2623_),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold275 (.A(\output_value_inst.led_data_reg[8] ),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0703_),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold277 (.A(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[2] ),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold278 (.A(_1688_),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0304_),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold280 (.A(\uart_tx_fifo_inst.fifo[4][3] ),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold281 (.A(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[2] ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold282 (.A(_2541_),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0744_),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold284 (.A(\input_value_check_inst.character_buff[6][2] ),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0464_),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold286 (.A(\uart_tx_fifo_inst.fifo[0][5] ),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold287 (.A(\uart_tx_fifo_inst.fifo[0][6] ),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold288 (.A(\input_value_check_inst.character_buff[7][0] ),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0446_),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold290 (.A(\output_value_inst.character_buff[2][3] ),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold291 (.A(_2419_),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold292 (.A(\uart_inst.uart_rx_inst.DATA_TEMP_REG[4] ),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold293 (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[7] ),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold294 (.A(_2524_),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0735_),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold296 (.A(\input_value_check_inst.character_buff[4][1] ),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0471_),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0106_),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold299 (.A(\output_value_inst.character_buff[1][2] ),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0668_),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold301 (.A(\uart_tx_fifo_inst.fifo[4][4] ),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold302 (.A(_2288_),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold303 (.A(\input_value_check_inst.character_buff[1][5] ),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0507_),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold305 (.A(\input_value_check_inst.character_buff[9][1] ),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0439_),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold307 (.A(\input_value_check_inst.character_buff[8][3] ),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0441_),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold309 (.A(\output_value_inst.led_data_reg[0] ),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0695_),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold311 (.A(\uart_tx_fifo_inst.fifo[4][5] ),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold312 (.A(_2289_),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold313 (.A(\uart_tx_fifo_inst.fifo[2][2] ),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold314 (.A(\input_value_check_inst.character_buff[3][1] ),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold315 (.A(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[2] ),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold316 (.A(_1436_),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0234_),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold318 (.A(\output_value_inst.led_data_reg[4] ),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0699_),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold320 (.A(\uart_tx_fifo_inst.fifo[9][6] ),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold321 (.A(_2626_),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold322 (.A(\input_value_check_inst.character_buff[6][4] ),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0458_),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold324 (.A(\uart_tx_fifo_inst.fifo[5][5] ),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold325 (.A(\input_value_check_inst.character_buff[5][7] ),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0477_),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold327 (.A(\uart_inst.uart_rx_inst.state[1] ),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold328 (.A(\uart_tx_fifo_inst.fifo[9][0] ),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold329 (.A(_2619_),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold330 (.A(\input_value_check_inst.character_buff[7][2] ),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold331 (.A(\uart_tx_fifo_inst.fifo[4][6] ),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold332 (.A(\uart_tx_fifo_inst.fifo[1][5] ),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold333 (.A(\uart_inst.uart_rx_inst.DATA_TEMP_REG[1] ),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0393_),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold335 (.A(\output_value_inst.character_buff[4][1] ),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold336 (.A(\output_value_inst.led_data_reg[12] ),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0707_),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold338 (.A(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[2] ),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold339 (.A(_1708_),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0311_),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold341 (.A(\output_value_inst.character_buff[6][6] ),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0638_),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold343 (.A(\input_value_check_inst.character_buff[2][5] ),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold344 (.A(\uart_tx_fifo_inst.fifo[1][0] ),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold345 (.A(_2257_),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold346 (.A(\output_value_inst.character_buff[6][0] ),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold347 (.A(_0075_),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0596_),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold349 (.A(\uart_tx_fifo_inst.fifo[3][6] ),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold350 (.A(\uart_tx_fifo_inst.fifo[9][4] ),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold351 (.A(_2624_),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold352 (.A(\uart_tx_fifo_inst.fifo[9][5] ),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold353 (.A(_2625_),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold354 (.A(\uart_tx_fifo_inst.fifo[0][0] ),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold355 (.A(\uart_tx_fifo_inst.fifo[9][1] ),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold356 (.A(_2621_),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold357 (.A(\output_value_inst.character_buff[5][2] ),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold358 (.A(\output_value_inst.output_valid ),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold359 (.A(\rx_data[6] ),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold360 (.A(\input_value_check_inst.character_buff[4][5] ),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold361 (.A(_0475_),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold362 (.A(\Led_Cycle_inst.clk_reducer.counter[30] ),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold363 (.A(_1896_),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0367_),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold365 (.A(\input_value_check_inst.character_buff[6][6] ),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0460_),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold367 (.A(tx_valid),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold368 (.A(\output_value_inst.character_buff[4][0] ),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold369 (.A(\input_value_check_inst.character_buff[7][1] ),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0447_),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold371 (.A(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[2] ),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold372 (.A(_1599_),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0276_),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold374 (.A(\output_value_inst.character_buff[2][6] ),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0665_),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold376 (.A(\output_value_inst.tx_ready ),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold377 (.A(_2094_),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold378 (.A(\uart_inst.uart_rx_inst.DATA_TEMP_REG[2] ),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold379 (.A(\output_value_inst.character_buff[3][5] ),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0657_),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold381 (.A(\uart_inst.tx_data[5] ),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0726_),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold383 (.A(\output_value_inst.character_buff[5][6] ),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold384 (.A(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[2] ),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold385 (.A(_1578_),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0269_),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold387 (.A(\input_value_check_inst.character_buff[5][4] ),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold388 (.A(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[2] ),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold389 (.A(_1677_),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0297_),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold391 (.A(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[2] ),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold392 (.A(_1754_),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0325_),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold394 (.A(\output_value_inst.character_buff[6][1] ),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold395 (.A(\input_value_check_inst.character_buff[4][4] ),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0149_),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0543_),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold398 (.A(_0180_),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold399 (.A(_1875_),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold400 (.A(\input_value_check_inst.character_buff[8][5] ),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0443_),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold402 (.A(\input_value_check_inst.character_buff[8][2] ),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold403 (.A(\input_value_check_inst.character_buff[4][2] ),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0472_),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold405 (.A(\output_value_inst.character_buff[6][2] ),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold406 (.A(\input_value_check_inst.character_buff[8][7] ),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0445_),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold408 (.A(\uart_inst.uart_rx_inst.SAMPLING_COUNT[1] ),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold409 (.A(_2029_),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0415_),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold411 (.A(\uart_tx_fifo_inst.fifo[6][3] ),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold412 (.A(\output_value_inst.character_buff[4][3] ),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold413 (.A(_2402_),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold414 (.A(\input_value_check_inst.character_buff[6][0] ),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold415 (.A(\input_value_check_inst.character_buff[3][2] ),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold416 (.A(\output_value_inst.character_buff[3][3] ),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0076_),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold418 (.A(_0597_),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold419 (.A(\uart_tx_fifo_inst.fifo[5][0] ),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold420 (.A(\output_value_inst.character_buff[4][4] ),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold421 (.A(\input_value_check_inst.character_buff[0][6] ),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold422 (.A(\input_value_check_inst.character_buff[5][0] ),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0470_),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold424 (.A(\input_value_check_inst.character_buff[7][7] ),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold425 (.A(\input_value_check_inst.character_buff[6][7] ),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold426 (.A(\output_value_inst.led_data_reg[15] ),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0710_),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold428 (.A(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[2] ),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold429 (.A(_1516_),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0248_),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold431 (.A(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[2] ),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold432 (.A(_1474_),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold433 (.A(_0241_),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold434 (.A(\uart_inst.uart_rx_inst.DATA_CNT[0] ),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold435 (.A(\uart_tx_fifo_inst.fifo[5][1] ),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold436 (.A(\output_value_inst.character_buff[6][4] ),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold437 (.A(_0637_),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold438 (.A(\input_value_check_inst.character_buff[4][3] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold439 (.A(_0481_),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold440 (.A(\uart_tx_fifo_inst.fifo[3][1] ),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold441 (.A(\uart_tx_fifo_inst.fifo[7][0] ),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold442 (.A(_1401_),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold443 (.A(\input_value_check_inst.character_buff[3][7] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold444 (.A(_0485_),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold445 (.A(_0078_),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0599_),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold447 (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[5] ),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold448 (.A(_2522_),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold449 (.A(\input_value_check_inst.character_buff[7][3] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold450 (.A(\output_value_inst.character_buff[6][3] ),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold451 (.A(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[2] ),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold452 (.A(_1728_),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold453 (.A(_0318_),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold454 (.A(\input_value_check_inst.character_buff[1][6] ),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold455 (.A(rx_valid),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold456 (.A(\Led_Cycle_inst.buttons[4] ),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold457 (.A(_0620_),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold458 (.A(\input_value_check_inst.character_buff[9][2] ),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold459 (.A(\input_value_check_inst.character_buff[6][3] ),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold460 (.A(_0465_),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold461 (.A(\tx_data[2] ),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold462 (.A(_0723_),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold463 (.A(\Led_Cycle_inst.clk_reducer.counter[2] ),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold464 (.A(_1840_),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold465 (.A(_0339_),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold466 (.A(_0073_),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold467 (.A(_0594_),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold468 (.A(\tx_data[3] ),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold469 (.A(_0751_),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold470 (.A(\output_value_inst.character_buff[2][5] ),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold471 (.A(_2422_),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold472 (.A(\uart_tx_fifo_inst.fifo[5][4] ),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold473 (.A(\input_value_check_inst.character_buff[7][5] ),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold474 (.A(\tx_data[1] ),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold475 (.A(_0722_),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold476 (.A(\input_value_check_inst.character_buff[6][1] ),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold477 (.A(\uart_inst.tx_data[6] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold478 (.A(_0727_),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold479 (.A(\input_value_check_inst.character_buff[3][6] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold480 (.A(_0484_),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold481 (.A(\input_value_check_inst.character_buff[2][7] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold482 (.A(\uart_tx_fifo_inst.fifo[7][5] ),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold483 (.A(_1429_),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold484 (.A(\input_value_check_inst.character_buff[6][5] ),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold485 (.A(\uart_inst.uart_rx_inst.CLK_CNT[1] ),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold486 (.A(_2001_),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold487 (.A(_0405_),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold488 (.A(\input_value_check_inst.character_buff[5][3] ),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold489 (.A(\input_value_check_inst.character_buff[5][1] ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold490 (.A(\input_value_check_inst.character_buff[2][6] ),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold491 (.A(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[1] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold492 (.A(_1687_),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold493 (.A(\uart_tx_fifo_inst.fifo_valid[4] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold494 (.A(_0524_),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold495 (.A(\input_value_check_inst.character_buff[8][4] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold496 (.A(_0442_),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold497 (.A(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[2] ),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold498 (.A(_1630_),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold499 (.A(_0283_),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold500 (.A(\uart_inst.uart_tx_inst.DATA_CNT[2] ),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold501 (.A(_2046_),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold502 (.A(\input_value_check_inst.character_buff[4][6] ),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold503 (.A(_0476_),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold504 (.A(\tx_data[0] ),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold505 (.A(_0721_),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold506 (.A(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[1] ),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold507 (.A(_1552_),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold508 (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[4] ),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold509 (.A(_2520_),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold510 (.A(\uart_inst.uart_rx_inst.SIGNAL_R ),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold511 (.A(\uart_tx_fifo_inst.fifo[8][2] ),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold512 (.A(_1426_),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold513 (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[8] ),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold514 (.A(_2526_),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold515 (.A(\uart_inst.uart_tx_inst.CLK_CNT[1] ),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold516 (.A(_0427_),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold517 (.A(\input_value_check_inst.character_buff[5][5] ),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold518 (.A(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[1] ),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold519 (.A(_1577_),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold520 (.A(\input_value_check_inst.character_buff[7][6] ),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold521 (.A(_0452_),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold522 (.A(\input_value_check_inst.character_buff[1][7] ),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold523 (.A(_0509_),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold524 (.A(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[1] ),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold525 (.A(_1536_),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold526 (.A(\uart_tx_fifo_inst.fifo[0][5] ),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold527 (.A(_2603_),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold528 (.A(_0753_),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold529 (.A(\input_value_check_inst.character_buff[5][6] ),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold530 (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[9] ),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold531 (.A(tx_signal),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold532 (.A(_0436_),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold533 (.A(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[1] ),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold534 (.A(_1654_),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold535 (.A(\input_value_check_inst.character_buff[1][2] ),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold536 (.A(\input_value_check_inst.character_buff[7][4] ),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold537 (.A(\uart_inst.uart_rx_inst.SIGNAL_Q[1] ),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold538 (.A(_0417_),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold539 (.A(\uart_inst.uart_rx_inst.SIGNAL_Q[0] ),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold540 (.A(\uart_inst.uart_tx_inst.DATA_REG[3] ),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold541 (.A(\uart_inst.uart_rx_inst.DATA_CNT[1] ),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold542 (.A(\Led_Cycle_inst.clk_reducer.counter[3] ),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold543 (.A(_1842_),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold544 (.A(\input_value_check_inst.character_buff[8][0] ),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold545 (.A(_0438_),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold546 (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[11] ),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold547 (.A(_2532_),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold548 (.A(_0739_),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold549 (.A(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[2] ),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold550 (.A(_1553_),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold551 (.A(_0262_),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold552 (.A(\Led_Cycle_inst.clk_reducer.counter[9] ),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold553 (.A(_1854_),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold554 (.A(\Led_Cycle_inst.clk_reducer.counter[12] ),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold555 (.A(_1862_),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold556 (.A(_0349_),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold557 (.A(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[3] ),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold558 (.A(_1517_),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold559 (.A(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[3] ),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold560 (.A(_1755_),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold561 (.A(\uart_inst.tx_data[4] ),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold562 (.A(_0725_),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold563 (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[12] ),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold564 (.A(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[3] ),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold565 (.A(_1631_),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold566 (.A(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[1] ),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold567 (.A(_1629_),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold568 (.A(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[3] ),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold569 (.A(_2542_),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold570 (.A(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[1] ),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold571 (.A(_1676_),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold572 (.A(\uart_tx_fifo_inst.fifo[2][0] ),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold573 (.A(\uart_tx_fifo_inst.fifo[8][4] ),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold574 (.A(\uart_tx_fifo_inst.fifo_valid[8] ),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold575 (.A(_2206_),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold576 (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[10] ),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold577 (.A(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[1] ),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold578 (.A(_1515_),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold579 (.A(\uart_tx_fifo_inst.fifo[4][1] ),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold580 (.A(\input_value_check_inst.character_buff[3][5] ),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold581 (.A(\uart_tx_fifo_inst.fifo_valid[9] ),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold582 (.A(\Led_Cycle_inst.clk_reducer.counter[31] ),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold583 (.A(_1898_),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold584 (.A(\uart_inst.uart_rx_inst.CLK_CNT[9] ),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold585 (.A(_2024_),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold586 (.A(_0413_),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold587 (.A(\Led_Cycle_inst.clk_reducer.counter[26] ),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold588 (.A(_1888_),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold589 (.A(_0363_),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold590 (.A(\input_value_check_inst.character_buff[3][4] ),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold591 (.A(uo_out[0]),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold592 (.A(_0600_),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold593 (.A(\uart_tx_fifo_inst.fifo[4][6] ),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold594 (.A(\output_value_inst.character_buff[1][1] ),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold595 (.A(_2426_),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold596 (.A(_0667_),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold597 (.A(\Led_Cycle_inst.buttons[0] ),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold598 (.A(_0109_),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold599 (.A(_2077_),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold600 (.A(_0434_),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold601 (.A(\input_value_check_inst.character_buff[1][3] ),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold602 (.A(_0505_),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold603 (.A(\uart_inst.uart_rx_inst.CLK_CNT[5] ),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold604 (.A(_2017_),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold605 (.A(_0074_),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold606 (.A(_0595_),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold607 (.A(\Led_Cycle_inst.clk_reducer.counter[27] ),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold608 (.A(_1890_),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold609 (.A(_0077_),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold610 (.A(_0598_),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold611 (.A(\output_value_inst.character_buff[1][4] ),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold612 (.A(_2431_),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold613 (.A(_0670_),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold614 (.A(\input_value_check_inst.character_buff[2][2] ),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold615 (.A(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[3] ),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold616 (.A(_1579_),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold617 (.A(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[3] ),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold618 (.A(_1784_),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold619 (.A(\output_value_inst.element_data_reg[11] ),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold620 (.A(_0694_),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold621 (.A(\Led_Cycle_inst.buttons[1] ),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold622 (.A(\Led_Cycle_inst.clk_reducer.counter[24] ),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold623 (.A(_1885_),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold624 (.A(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[3] ),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold625 (.A(_1729_),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold626 (.A(\output_value_inst.character_buff[5][4] ),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold627 (.A(\uart_tx_fifo_inst.fifo_valid[2] ),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold628 (.A(_0522_),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold629 (.A(uo_out[1]),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold630 (.A(_0601_),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold631 (.A(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[3] ),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold632 (.A(_1600_),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold633 (.A(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[3] ),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold634 (.A(_1709_),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold635 (.A(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[3] ),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold636 (.A(_1656_),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold637 (.A(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[3] ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold638 (.A(_1475_),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold639 (.A(_0171_),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold640 (.A(_1722_),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold641 (.A(_0315_),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold642 (.A(\output_value_inst.character_buff[1][5] ),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold643 (.A(_2433_),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold644 (.A(_0671_),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold645 (.A(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[3] ),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold646 (.A(_1437_),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold647 (.A(\input_value_check_inst.character_buff[2][3] ),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold648 (.A(\uart_inst.uart_rx_inst.SIGNAL_Q[2] ),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold649 (.A(_0418_),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold650 (.A(\uart_tx_fifo_inst.fifo_valid[3] ),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold651 (.A(\output_value_inst.character_buff[2][0] ),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold652 (.A(_2413_),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold653 (.A(_0659_),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold654 (.A(\uart_inst.uart_rx_inst.DATA_CNT[2] ),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold655 (.A(\uart_inst.uart_rx_inst.CLK_CNT[2] ),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold656 (.A(_0406_),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold657 (.A(\Led_Cycle_inst.clk_reducer.counter[15] ),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold658 (.A(_1867_),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold659 (.A(\input_value_check_inst.character_buff[1][4] ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold660 (.A(_0498_),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold661 (.A(\uart_tx_fifo_inst.fifo_valid[0] ),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold662 (.A(_0521_),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold663 (.A(\output_value_inst.character_buff[2][1] ),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold664 (.A(_2415_),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold665 (.A(\Led_Cycle_inst.clk_reducer.counter[28] ),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold666 (.A(_1892_),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold667 (.A(\output_value_inst.character_buff[1][0] ),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold668 (.A(_2424_),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold669 (.A(_0666_),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold670 (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[2] ),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold671 (.A(_2516_),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold672 (.A(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[0] ),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold673 (.A(_1753_),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold674 (.A(\uart_tx_fifo_inst.fifo[3][0] ),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold675 (.A(\uart_inst.uart_tx_inst.CLK_CNT[6] ),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold676 (.A(\output_value_inst.element_data_reg[7] ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold677 (.A(\input_value_check_inst.character_buff[0][4] ),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold678 (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[6] ),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold679 (.A(\Led_Cycle_inst.clk_reducer.counter[20] ),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold680 (.A(_1877_),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold681 (.A(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[3] ),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold682 (.A(_1689_),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold683 (.A(\uart_inst.uart_rx_inst.state[0] ),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold684 (.A(_0134_),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold685 (.A(_2055_),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold686 (.A(_0426_),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold687 (.A(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[1] ),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold688 (.A(_1598_),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold689 (.A(_0099_),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold690 (.A(\Led_Cycle_inst.clk_reducer.counter[4] ),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold691 (.A(_1844_),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold692 (.A(\input_value_check_inst.character_buff[4][0] ),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold693 (.A(_0478_),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold694 (.A(\output_value_inst.character_buff[2][2] ),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold695 (.A(\output_value_inst.character_buff[2][4] ),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold696 (.A(_2420_),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold697 (.A(\Led_Cycle_inst.clk_reducer.counter[14] ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold698 (.A(_1865_),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold699 (.A(\input_value_check_inst.character_buff[2][4] ),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold700 (.A(\uart_inst.uart_tx_inst.state[2] ),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold701 (.A(_0054_),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold702 (.A(\output_value_inst.character_buff[7][0] ),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold703 (.A(_2368_),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold704 (.A(\Led_Cycle_inst.clk_reducer.counter[11] ),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold705 (.A(_1859_),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold706 (.A(\uart_inst.uart_rx_inst.SIGNAL_Q[4] ),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold707 (.A(\uart_inst.uart_tx_inst.CLK_CNT[2] ),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold708 (.A(_2060_),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold709 (.A(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[0] ),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold710 (.A(_1473_),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold711 (.A(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[1] ),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold712 (.A(_1435_),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold713 (.A(\SegmentDisplay.seg_driver.clk_reducer.counter[1] ),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold714 (.A(_2509_),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold715 (.A(_0729_),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold716 (.A(\uart_inst.uart_rx_inst.SIGNAL_Q[3] ),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold717 (.A(_0419_),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold718 (.A(\uart_inst.uart_tx_inst.CLK_CNT[5] ),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold719 (.A(_2069_),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold720 (.A(_0431_),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold721 (.A(\output_value_inst.character_buff[0][6] ),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold722 (.A(_0672_),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold723 (.A(_0120_),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold724 (.A(_0607_),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold725 (.A(\uart_inst.uart_rx_inst.CLK_CNT[0] ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold726 (.A(_0404_),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold727 (.A(\uart_inst.uart_tx_inst.CLK_CNT[4] ),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold728 (.A(_2068_),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold729 (.A(\uart_inst.uart_tx_inst.state[1] ),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold730 (.A(_1007_),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold731 (.A(_0053_),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold732 (.A(\uart_tx_fifo_inst.fifo_valid[7] ),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold733 (.A(_0527_),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold734 (.A(\output_value_inst.character_buff[0][3] ),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold735 (.A(_0669_),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold736 (.A(\uart_tx_fifo_inst.fifo_valid[5] ),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold737 (.A(\output_value_inst.element_data_reg[8] ),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold738 (.A(\uart_inst.uart_rx_inst.CLK_CNT[7] ),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold739 (.A(\Led_Cycle_inst.clk_reducer.counter[29] ),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold740 (.A(\output_value_inst.character_buff[8][6] ),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold741 (.A(_2364_),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold742 (.A(\input_value_check_inst.character_buff[3][3] ),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold743 (.A(\Led_Cycle_inst.clk_reducer.counter[6] ),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold744 (.A(_1847_),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold745 (.A(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[1] ),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold746 (.A(_1727_),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold747 (.A(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[3] ),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold748 (.A(_1538_),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold749 (.A(\uart_tx_fifo_inst.fifo_valid[6] ),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold750 (.A(\Led_Cycle_inst.clk_reducer.counter[5] ),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold751 (.A(\input_value_check_inst.character_buff[1][1] ),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold752 (.A(\uart_inst.uart_rx_inst.state[2] ),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold753 (.A(\Led_Cycle_inst.clk_reducer.counter[25] ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold754 (.A(\Led_Cycle_inst.clk_reducer.counter[1] ),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold755 (.A(_1838_),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold756 (.A(\output_value_inst.character_buff[9][2] ),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold757 (.A(_2228_),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold758 (.A(\output_value_inst.character_buff[7][2] ),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold759 (.A(_2376_),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold760 (.A(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[3] ),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold761 (.A(_1554_),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold762 (.A(\output_value_inst.character_buff[8][4] ),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold763 (.A(_2360_),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold764 (.A(\output_value_inst.character_buff[9][6] ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold765 (.A(_2240_),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold766 (.A(\input_value_check_inst.character_buff[1][0] ),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold767 (.A(\Led_Cycle_inst.clk_reducer.counter[10] ),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold768 (.A(_1858_),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold769 (.A(\uart_inst.uart_rx_inst.CLK_CNT[8] ),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold770 (.A(\output_value_inst.character_buff[8][0] ),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold771 (.A(_2344_),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold772 (.A(\SegmentDisplay.bcd3[3] ),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold773 (.A(_1185_),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold774 (.A(\uart_inst.uart_rx_inst.CLK_CNT[3] ),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold775 (.A(_0407_),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold776 (.A(\output_value_inst.character_buff[7][3] ),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold777 (.A(_2380_),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold778 (.A(\uart_inst.uart_rx_inst.SIGNAL_Q[3] ),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold779 (.A(\output_value_inst.character_buff[8][1] ),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold780 (.A(_2348_),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold781 (.A(\output_value_inst.character_buff[7][1] ),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold782 (.A(_2372_),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold783 (.A(\output_value_inst.character_buff[9][0] ),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold784 (.A(_2220_),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold785 (.A(\Led_Cycle_inst.clk_reducer.counter[21] ),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold786 (.A(_0110_),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold787 (.A(_1849_),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold788 (.A(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[3] ),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold789 (.A(_1678_),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold790 (.A(\output_value_inst.character_buff[7][6] ),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold791 (.A(_2388_),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold792 (.A(\output_value_inst.character_buff[8][2] ),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold793 (.A(_2352_),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold794 (.A(\Led_Cycle_inst.clk_reducer.counter[13] ),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold795 (.A(_1864_),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold796 (.A(\Led_Cycle_inst.clk_reducer.counter[16] ),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold797 (.A(\output_value_inst.character_buff[9][4] ),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold798 (.A(_2236_),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold799 (.A(\input_value_check_inst.character_buff[2][1] ),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold800 (.A(_0139_),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold801 (.A(_1161_),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold802 (.A(_0532_),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold803 (.A(\output_value_inst.element_data_reg[0] ),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold804 (.A(\input_value_check_inst.character_buff[2][0] ),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold805 (.A(\uart_inst.uart_tx_inst.CLK_CNT[3] ),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold806 (.A(_2065_),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold807 (.A(\output_value_inst.character_buff[8][3] ),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold808 (.A(_2232_),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold809 (.A(\input_value_check_inst.character_buff[3][0] ),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold810 (.A(_0122_),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold811 (.A(_1096_),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold812 (.A(_0719_),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold813 (.A(\output_value_inst.character_buff[7][4] ),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold814 (.A(_2384_),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold815 (.A(\uart_inst.uart_tx_inst.DATA_CNT[1] ),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold816 (.A(\Led_Cycle_inst.buttons[3] ),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold817 (.A(_0144_),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold818 (.A(_0064_),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold819 (.A(\Led_Cycle_inst.clk_reducer.counter[18] ),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold820 (.A(_1873_),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold821 (.A(_0130_),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold822 (.A(_1157_),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold823 (.A(_0018_),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold824 (.A(\output_value_inst.character_buff[9][1] ),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold825 (.A(_2224_),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold826 (.A(\Led_Cycle_inst.buttons[2] ),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold827 (.A(\uart_inst.uart_tx_inst.CLK_CNT[9] ),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold828 (.A(_2078_),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold829 (.A(\output_value_inst.led_data_reg[5] ),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold830 (.A(_1361_),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold831 (.A(_0371_),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold832 (.A(\uart_inst.uart_tx_inst.state[0] ),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold833 (.A(_0052_),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold834 (.A(\Led_Cycle_inst.clk_reducer.counter[23] ),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold835 (.A(\output_value_inst.led_data_reg[2] ),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold836 (.A(_1100_),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold837 (.A(_0720_),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold838 (.A(\uart_inst.uart_rx_inst.CLK_CNT[4] ),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold839 (.A(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[4] ),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold840 (.A(_0164_),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold841 (.A(\output_value_inst.led_data_reg[14] ),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold842 (.A(_1165_),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold843 (.A(_0533_),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold844 (.A(_0145_),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold845 (.A(_0421_),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold846 (.A(\Led_Cycle_inst.clk_reducer.counter[22] ),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold847 (.A(\Led_Cycle_inst.genblk1[4].pwm_unit.counter[4] ),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold848 (.A(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[0] ),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold849 (.A(_1702_),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold850 (.A(_0310_),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold851 (.A(_0125_),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold852 (.A(_1102_),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold853 (.A(_1105_),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold854 (.A(_0029_),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold855 (.A(\Led_Cycle_inst.clk_reducer.counter[8] ),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold856 (.A(\Led_Cycle_inst.genblk1[8].pwm_unit.counter[4] ),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold857 (.A(\uart_inst.uart_tx_inst.DATA_CNT[0] ),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold858 (.A(_0107_),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold859 (.A(\Led_Cycle_inst.genblk1[10].pwm_unit.counter[4] ),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold860 (.A(\Led_Cycle_inst.genblk1[3].pwm_unit.counter[4] ),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold861 (.A(_0160_),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold862 (.A(_1360_),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold863 (.A(_0372_),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold864 (.A(\Led_Cycle_inst.genblk1[13].pwm_unit.counter[4] ),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold865 (.A(\Led_Cycle_inst.genblk1[2].pwm_unit.counter[4] ),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold866 (.A(_0105_),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold867 (.A(\Led_Cycle_inst.genblk1[15].pwm_unit.counter[4] ),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold868 (.A(\Led_Cycle_inst.genblk1[1].pwm_unit.counter[4] ),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold869 (.A(\Led_Cycle_inst.genblk1[14].pwm_unit.counter[4] ),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold870 (.A(\Led_Cycle_inst.genblk1[9].pwm_unit.counter[1] ),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold871 (.A(_1612_),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold872 (.A(_0743_),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold873 (.A(_0142_),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold874 (.A(_1167_),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold875 (.A(_1170_),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold876 (.A(_0038_),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold877 (.A(\Led_Cycle_inst.genblk1[11].pwm_unit.counter[4] ),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold878 (.A(\Led_Cycle_inst.genblk1[6].pwm_unit.counter[4] ),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold879 (.A(\Led_Cycle_inst.genblk1[7].pwm_unit.counter[4] ),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold880 (.A(\Led_Cycle_inst.genblk1[5].pwm_unit.counter[4] ),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold881 (.A(\Led_Cycle_inst.genblk1[12].pwm_unit.counter[4] ),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold882 (.A(_0163_),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold883 (.A(_1366_),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold884 (.A(_1369_),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold885 (.A(_0032_),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold886 (.A(\Led_Cycle_inst.genblk1[0].pwm_unit.counter[4] ),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold887 (.A(_0102_),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold888 (.A(_0124_),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold889 (.A(_1104_),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold890 (.A(\SegmentDisplay.bcd3[2] ),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold891 (.A(uo_out[2]),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold892 (.A(_0101_),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold893 (.A(_0042_),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold894 (.A(_0161_),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold895 (.A(_0147_),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold896 (.A(_1224_),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold897 (.A(_0103_),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold898 (.A(_0127_),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold899 (.A(\Led_Cycle_inst.clk_reducer.counter[17] ),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold900 (.A(\SegmentDisplay.bcd2[3] ),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold901 (.A(_1139_),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold902 (.A(\output_value_inst.led_data_reg[6] ),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold903 (.A(_1364_),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold904 (.A(_0033_),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold905 (.A(_0155_),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold906 (.A(_0148_),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold907 (.A(\output_value_inst.led_data_reg[10] ),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold908 (.A(_1222_),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold909 (.A(_1219_),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold910 (.A(_0140_),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold911 (.A(_1171_),
    .X(net1757));
 sg13g2_dlygate4sd3_1 hold912 (.A(\output_value_inst.element_data_reg[9] ),
    .X(net1758));
 sg13g2_dlygate4sd3_1 hold913 (.A(\Led_Cycle_inst.genblk1[1].pwm_unit.pwm_out ),
    .X(net1759));
 sg13g2_dlygate4sd3_1 hold914 (.A(_1097_),
    .X(net1760));
 sg13g2_dlygate4sd3_1 hold915 (.A(_0118_),
    .X(net1761));
 sg13g2_dlygate4sd3_1 hold916 (.A(\Led_Cycle_inst.genblk1[13].pwm_unit.pwm_out ),
    .X(net1762));
 sg13g2_dlygate4sd3_1 hold917 (.A(_1162_),
    .X(net1763));
 sg13g2_dlygate4sd3_1 hold918 (.A(\SegmentDisplay.bcd2[2] ),
    .X(net1764));
 sg13g2_dlygate4sd3_1 hold919 (.A(_0119_),
    .X(net1765));
 sg13g2_dlygate4sd3_1 hold920 (.A(_0534_),
    .X(net1766));
 sg13g2_dlygate4sd3_1 hold921 (.A(\output_value_inst.element_data_reg[10] ),
    .X(net1767));
 sg13g2_dlygate4sd3_1 hold922 (.A(_0048_),
    .X(net1768));
 sg13g2_dlygate4sd3_1 hold923 (.A(uo_out[4]),
    .X(net1769));
 sg13g2_dlygate4sd3_1 hold924 (.A(_0151_),
    .X(net1770));
 sg13g2_dlygate4sd3_1 hold925 (.A(\output_value_inst.character_buff[6][2] ),
    .X(net1771));
 sg13g2_dlygate4sd3_1 hold926 (.A(_2462_),
    .X(net1772));
 sg13g2_dlygate4sd3_1 hold927 (.A(_2471_),
    .X(net1773));
 sg13g2_dlygate4sd3_1 hold928 (.A(\Led_Cycle_inst.clk_reducer.counter[23] ),
    .X(net1774));
 sg13g2_dlygate4sd3_1 hold929 (.A(_1886_),
    .X(net1775));
 sg13g2_dlygate4sd3_1 hold930 (.A(\uart_inst.uart_rx_inst.state[2] ),
    .X(net1776));
 sg13g2_dlygate4sd3_1 hold931 (.A(\Led_Cycle_inst.clk_reducer.counter[22] ),
    .X(net1777));
 sg13g2_dlygate4sd3_1 hold932 (.A(\Led_Cycle_inst.clk_reducer.counter[25] ),
    .X(net1778));
 sg13g2_dlygate4sd3_1 hold933 (.A(_0119_),
    .X(net1779));
 sg13g2_dlygate4sd3_1 hold934 (.A(\uart_inst.uart_tx_inst.DATA_CNT[0] ),
    .X(net1780));
 sg13g2_dlygate4sd3_1 hold935 (.A(\Led_Cycle_inst.clk_reducer.counter[8] ),
    .X(net1781));
 sg13g2_dlygate4sd3_1 hold936 (.A(\Led_Cycle_inst.genblk1[10].pwm_unit.pwm_out ),
    .X(net1782));
 sg13g2_dlygate4sd3_1 hold937 (.A(\uart_inst.uart_rx_inst.CLK_CNT[4] ),
    .X(net1783));
 sg13g2_dlygate4sd3_1 hold938 (.A(_0975_),
    .X(net1784));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_fill_1 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_138 ();
 sg13g2_decap_8 FILLER_14_145 ();
 sg13g2_decap_8 FILLER_14_152 ();
 sg13g2_decap_8 FILLER_14_159 ();
 sg13g2_decap_8 FILLER_14_166 ();
 sg13g2_decap_8 FILLER_14_173 ();
 sg13g2_decap_8 FILLER_14_180 ();
 sg13g2_decap_8 FILLER_14_187 ();
 sg13g2_decap_8 FILLER_14_194 ();
 sg13g2_decap_8 FILLER_14_201 ();
 sg13g2_decap_8 FILLER_14_208 ();
 sg13g2_decap_8 FILLER_14_215 ();
 sg13g2_decap_8 FILLER_14_222 ();
 sg13g2_decap_8 FILLER_14_229 ();
 sg13g2_decap_8 FILLER_14_236 ();
 sg13g2_decap_8 FILLER_14_243 ();
 sg13g2_decap_8 FILLER_14_250 ();
 sg13g2_decap_8 FILLER_14_257 ();
 sg13g2_decap_8 FILLER_14_264 ();
 sg13g2_decap_8 FILLER_14_271 ();
 sg13g2_decap_8 FILLER_14_278 ();
 sg13g2_decap_8 FILLER_14_285 ();
 sg13g2_decap_8 FILLER_14_292 ();
 sg13g2_decap_8 FILLER_14_299 ();
 sg13g2_decap_8 FILLER_14_306 ();
 sg13g2_decap_8 FILLER_14_313 ();
 sg13g2_decap_8 FILLER_14_320 ();
 sg13g2_decap_8 FILLER_14_327 ();
 sg13g2_decap_8 FILLER_14_334 ();
 sg13g2_decap_8 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_348 ();
 sg13g2_decap_8 FILLER_14_355 ();
 sg13g2_decap_8 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_8 FILLER_14_404 ();
 sg13g2_decap_8 FILLER_14_411 ();
 sg13g2_decap_8 FILLER_14_418 ();
 sg13g2_decap_8 FILLER_14_425 ();
 sg13g2_decap_8 FILLER_14_432 ();
 sg13g2_decap_8 FILLER_14_439 ();
 sg13g2_decap_8 FILLER_14_446 ();
 sg13g2_decap_8 FILLER_14_453 ();
 sg13g2_decap_8 FILLER_14_460 ();
 sg13g2_decap_8 FILLER_14_467 ();
 sg13g2_decap_8 FILLER_14_474 ();
 sg13g2_decap_8 FILLER_14_481 ();
 sg13g2_decap_8 FILLER_14_488 ();
 sg13g2_decap_8 FILLER_14_495 ();
 sg13g2_decap_8 FILLER_14_502 ();
 sg13g2_decap_8 FILLER_14_509 ();
 sg13g2_decap_8 FILLER_14_516 ();
 sg13g2_decap_8 FILLER_14_523 ();
 sg13g2_decap_8 FILLER_14_530 ();
 sg13g2_decap_8 FILLER_14_537 ();
 sg13g2_decap_8 FILLER_14_544 ();
 sg13g2_decap_8 FILLER_14_551 ();
 sg13g2_decap_8 FILLER_14_558 ();
 sg13g2_decap_8 FILLER_14_565 ();
 sg13g2_decap_8 FILLER_14_572 ();
 sg13g2_decap_8 FILLER_14_579 ();
 sg13g2_decap_8 FILLER_14_586 ();
 sg13g2_decap_8 FILLER_14_593 ();
 sg13g2_decap_8 FILLER_14_600 ();
 sg13g2_decap_8 FILLER_14_607 ();
 sg13g2_decap_8 FILLER_14_614 ();
 sg13g2_decap_8 FILLER_14_621 ();
 sg13g2_decap_8 FILLER_14_628 ();
 sg13g2_decap_8 FILLER_14_635 ();
 sg13g2_decap_8 FILLER_14_642 ();
 sg13g2_decap_8 FILLER_14_649 ();
 sg13g2_decap_8 FILLER_14_656 ();
 sg13g2_decap_8 FILLER_14_663 ();
 sg13g2_decap_8 FILLER_14_670 ();
 sg13g2_decap_8 FILLER_14_677 ();
 sg13g2_decap_8 FILLER_14_684 ();
 sg13g2_decap_8 FILLER_14_691 ();
 sg13g2_decap_8 FILLER_14_698 ();
 sg13g2_decap_8 FILLER_14_705 ();
 sg13g2_decap_8 FILLER_14_712 ();
 sg13g2_decap_8 FILLER_14_719 ();
 sg13g2_decap_8 FILLER_14_726 ();
 sg13g2_decap_8 FILLER_14_733 ();
 sg13g2_decap_8 FILLER_14_740 ();
 sg13g2_decap_8 FILLER_14_747 ();
 sg13g2_decap_8 FILLER_14_754 ();
 sg13g2_decap_8 FILLER_14_761 ();
 sg13g2_decap_8 FILLER_14_768 ();
 sg13g2_decap_8 FILLER_14_775 ();
 sg13g2_decap_8 FILLER_14_782 ();
 sg13g2_decap_8 FILLER_14_789 ();
 sg13g2_decap_8 FILLER_14_796 ();
 sg13g2_decap_8 FILLER_14_803 ();
 sg13g2_decap_8 FILLER_14_810 ();
 sg13g2_decap_8 FILLER_14_817 ();
 sg13g2_decap_8 FILLER_14_824 ();
 sg13g2_decap_8 FILLER_14_831 ();
 sg13g2_decap_8 FILLER_14_838 ();
 sg13g2_decap_8 FILLER_14_845 ();
 sg13g2_decap_8 FILLER_14_852 ();
 sg13g2_fill_2 FILLER_14_859 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_4 FILLER_15_77 ();
 sg13g2_fill_1 FILLER_15_81 ();
 sg13g2_fill_1 FILLER_15_87 ();
 sg13g2_fill_1 FILLER_15_97 ();
 sg13g2_fill_2 FILLER_15_103 ();
 sg13g2_fill_1 FILLER_15_105 ();
 sg13g2_fill_1 FILLER_15_114 ();
 sg13g2_fill_2 FILLER_15_151 ();
 sg13g2_decap_8 FILLER_15_157 ();
 sg13g2_decap_8 FILLER_15_164 ();
 sg13g2_decap_8 FILLER_15_171 ();
 sg13g2_decap_8 FILLER_15_178 ();
 sg13g2_decap_8 FILLER_15_185 ();
 sg13g2_decap_8 FILLER_15_192 ();
 sg13g2_decap_8 FILLER_15_199 ();
 sg13g2_decap_8 FILLER_15_206 ();
 sg13g2_decap_8 FILLER_15_213 ();
 sg13g2_decap_8 FILLER_15_220 ();
 sg13g2_decap_8 FILLER_15_227 ();
 sg13g2_decap_8 FILLER_15_234 ();
 sg13g2_decap_8 FILLER_15_241 ();
 sg13g2_decap_8 FILLER_15_248 ();
 sg13g2_decap_8 FILLER_15_255 ();
 sg13g2_decap_8 FILLER_15_262 ();
 sg13g2_fill_2 FILLER_15_269 ();
 sg13g2_fill_1 FILLER_15_271 ();
 sg13g2_fill_2 FILLER_15_276 ();
 sg13g2_decap_8 FILLER_15_282 ();
 sg13g2_decap_8 FILLER_15_289 ();
 sg13g2_decap_8 FILLER_15_296 ();
 sg13g2_decap_8 FILLER_15_303 ();
 sg13g2_decap_8 FILLER_15_310 ();
 sg13g2_decap_4 FILLER_15_317 ();
 sg13g2_fill_1 FILLER_15_321 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_4 FILLER_16_70 ();
 sg13g2_fill_1 FILLER_16_126 ();
 sg13g2_fill_2 FILLER_16_166 ();
 sg13g2_fill_1 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_173 ();
 sg13g2_decap_8 FILLER_16_180 ();
 sg13g2_decap_8 FILLER_16_187 ();
 sg13g2_decap_8 FILLER_16_194 ();
 sg13g2_decap_8 FILLER_16_201 ();
 sg13g2_decap_8 FILLER_16_208 ();
 sg13g2_decap_8 FILLER_16_215 ();
 sg13g2_decap_8 FILLER_16_222 ();
 sg13g2_decap_8 FILLER_16_229 ();
 sg13g2_decap_8 FILLER_16_236 ();
 sg13g2_fill_2 FILLER_16_243 ();
 sg13g2_fill_2 FILLER_16_258 ();
 sg13g2_fill_1 FILLER_16_260 ();
 sg13g2_fill_1 FILLER_16_276 ();
 sg13g2_fill_1 FILLER_16_282 ();
 sg13g2_decap_8 FILLER_16_291 ();
 sg13g2_decap_8 FILLER_16_298 ();
 sg13g2_decap_8 FILLER_16_305 ();
 sg13g2_decap_8 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_decap_8 FILLER_16_361 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_4 FILLER_16_382 ();
 sg13g2_fill_1 FILLER_16_386 ();
 sg13g2_decap_4 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_16_415 ();
 sg13g2_decap_8 FILLER_16_422 ();
 sg13g2_decap_8 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_16_436 ();
 sg13g2_decap_8 FILLER_16_443 ();
 sg13g2_decap_8 FILLER_16_450 ();
 sg13g2_decap_8 FILLER_16_457 ();
 sg13g2_decap_8 FILLER_16_464 ();
 sg13g2_decap_8 FILLER_16_471 ();
 sg13g2_decap_8 FILLER_16_478 ();
 sg13g2_decap_8 FILLER_16_485 ();
 sg13g2_decap_8 FILLER_16_492 ();
 sg13g2_decap_8 FILLER_16_499 ();
 sg13g2_decap_8 FILLER_16_506 ();
 sg13g2_decap_8 FILLER_16_513 ();
 sg13g2_decap_8 FILLER_16_520 ();
 sg13g2_decap_8 FILLER_16_527 ();
 sg13g2_decap_8 FILLER_16_534 ();
 sg13g2_decap_8 FILLER_16_541 ();
 sg13g2_decap_8 FILLER_16_548 ();
 sg13g2_decap_8 FILLER_16_555 ();
 sg13g2_decap_8 FILLER_16_562 ();
 sg13g2_decap_8 FILLER_16_569 ();
 sg13g2_decap_8 FILLER_16_576 ();
 sg13g2_decap_8 FILLER_16_583 ();
 sg13g2_decap_8 FILLER_16_590 ();
 sg13g2_decap_8 FILLER_16_597 ();
 sg13g2_decap_8 FILLER_16_604 ();
 sg13g2_decap_8 FILLER_16_611 ();
 sg13g2_decap_8 FILLER_16_618 ();
 sg13g2_decap_8 FILLER_16_625 ();
 sg13g2_decap_8 FILLER_16_632 ();
 sg13g2_decap_8 FILLER_16_639 ();
 sg13g2_decap_8 FILLER_16_646 ();
 sg13g2_decap_8 FILLER_16_653 ();
 sg13g2_decap_8 FILLER_16_660 ();
 sg13g2_decap_8 FILLER_16_667 ();
 sg13g2_decap_8 FILLER_16_674 ();
 sg13g2_decap_8 FILLER_16_681 ();
 sg13g2_decap_8 FILLER_16_688 ();
 sg13g2_decap_8 FILLER_16_695 ();
 sg13g2_decap_8 FILLER_16_702 ();
 sg13g2_decap_8 FILLER_16_709 ();
 sg13g2_decap_8 FILLER_16_716 ();
 sg13g2_decap_8 FILLER_16_723 ();
 sg13g2_decap_8 FILLER_16_730 ();
 sg13g2_decap_8 FILLER_16_737 ();
 sg13g2_decap_8 FILLER_16_744 ();
 sg13g2_decap_8 FILLER_16_751 ();
 sg13g2_decap_8 FILLER_16_758 ();
 sg13g2_decap_8 FILLER_16_765 ();
 sg13g2_decap_8 FILLER_16_772 ();
 sg13g2_decap_8 FILLER_16_779 ();
 sg13g2_decap_8 FILLER_16_786 ();
 sg13g2_decap_8 FILLER_16_793 ();
 sg13g2_decap_8 FILLER_16_800 ();
 sg13g2_decap_8 FILLER_16_807 ();
 sg13g2_decap_8 FILLER_16_814 ();
 sg13g2_decap_8 FILLER_16_821 ();
 sg13g2_decap_8 FILLER_16_828 ();
 sg13g2_decap_8 FILLER_16_835 ();
 sg13g2_decap_8 FILLER_16_842 ();
 sg13g2_decap_8 FILLER_16_849 ();
 sg13g2_decap_4 FILLER_16_856 ();
 sg13g2_fill_2 FILLER_16_860 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_fill_2 FILLER_17_89 ();
 sg13g2_fill_2 FILLER_17_96 ();
 sg13g2_fill_1 FILLER_17_98 ();
 sg13g2_fill_2 FILLER_17_177 ();
 sg13g2_decap_8 FILLER_17_183 ();
 sg13g2_decap_8 FILLER_17_190 ();
 sg13g2_decap_8 FILLER_17_197 ();
 sg13g2_decap_8 FILLER_17_204 ();
 sg13g2_decap_4 FILLER_17_211 ();
 sg13g2_fill_2 FILLER_17_215 ();
 sg13g2_fill_2 FILLER_17_243 ();
 sg13g2_fill_2 FILLER_17_254 ();
 sg13g2_fill_1 FILLER_17_256 ();
 sg13g2_fill_1 FILLER_17_266 ();
 sg13g2_fill_1 FILLER_17_272 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_fill_2 FILLER_17_371 ();
 sg13g2_fill_1 FILLER_17_373 ();
 sg13g2_fill_2 FILLER_17_400 ();
 sg13g2_fill_2 FILLER_17_411 ();
 sg13g2_decap_8 FILLER_17_417 ();
 sg13g2_decap_8 FILLER_17_424 ();
 sg13g2_decap_8 FILLER_17_431 ();
 sg13g2_decap_8 FILLER_17_438 ();
 sg13g2_decap_8 FILLER_17_445 ();
 sg13g2_decap_8 FILLER_17_452 ();
 sg13g2_decap_8 FILLER_17_459 ();
 sg13g2_decap_8 FILLER_17_466 ();
 sg13g2_decap_8 FILLER_17_473 ();
 sg13g2_decap_8 FILLER_17_480 ();
 sg13g2_decap_8 FILLER_17_487 ();
 sg13g2_decap_8 FILLER_17_494 ();
 sg13g2_decap_8 FILLER_17_501 ();
 sg13g2_decap_8 FILLER_17_508 ();
 sg13g2_decap_8 FILLER_17_515 ();
 sg13g2_decap_8 FILLER_17_522 ();
 sg13g2_decap_8 FILLER_17_529 ();
 sg13g2_decap_8 FILLER_17_536 ();
 sg13g2_decap_8 FILLER_17_543 ();
 sg13g2_decap_8 FILLER_17_550 ();
 sg13g2_decap_8 FILLER_17_557 ();
 sg13g2_decap_8 FILLER_17_564 ();
 sg13g2_decap_8 FILLER_17_571 ();
 sg13g2_decap_8 FILLER_17_578 ();
 sg13g2_decap_8 FILLER_17_585 ();
 sg13g2_decap_8 FILLER_17_592 ();
 sg13g2_decap_8 FILLER_17_599 ();
 sg13g2_decap_8 FILLER_17_606 ();
 sg13g2_decap_8 FILLER_17_613 ();
 sg13g2_decap_8 FILLER_17_620 ();
 sg13g2_decap_8 FILLER_17_627 ();
 sg13g2_decap_8 FILLER_17_634 ();
 sg13g2_decap_8 FILLER_17_641 ();
 sg13g2_decap_8 FILLER_17_648 ();
 sg13g2_decap_8 FILLER_17_655 ();
 sg13g2_decap_8 FILLER_17_662 ();
 sg13g2_decap_8 FILLER_17_669 ();
 sg13g2_decap_8 FILLER_17_676 ();
 sg13g2_decap_8 FILLER_17_683 ();
 sg13g2_decap_8 FILLER_17_690 ();
 sg13g2_decap_8 FILLER_17_697 ();
 sg13g2_decap_8 FILLER_17_704 ();
 sg13g2_decap_8 FILLER_17_711 ();
 sg13g2_decap_8 FILLER_17_718 ();
 sg13g2_decap_8 FILLER_17_725 ();
 sg13g2_decap_8 FILLER_17_732 ();
 sg13g2_decap_8 FILLER_17_739 ();
 sg13g2_decap_8 FILLER_17_746 ();
 sg13g2_decap_8 FILLER_17_753 ();
 sg13g2_decap_8 FILLER_17_760 ();
 sg13g2_decap_8 FILLER_17_767 ();
 sg13g2_decap_8 FILLER_17_774 ();
 sg13g2_decap_8 FILLER_17_781 ();
 sg13g2_decap_8 FILLER_17_788 ();
 sg13g2_decap_8 FILLER_17_795 ();
 sg13g2_decap_8 FILLER_17_802 ();
 sg13g2_decap_8 FILLER_17_809 ();
 sg13g2_decap_8 FILLER_17_816 ();
 sg13g2_decap_8 FILLER_17_823 ();
 sg13g2_decap_8 FILLER_17_830 ();
 sg13g2_decap_8 FILLER_17_837 ();
 sg13g2_decap_8 FILLER_17_844 ();
 sg13g2_decap_8 FILLER_17_851 ();
 sg13g2_decap_4 FILLER_17_858 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_4 FILLER_18_49 ();
 sg13g2_fill_2 FILLER_18_79 ();
 sg13g2_fill_1 FILLER_18_148 ();
 sg13g2_fill_1 FILLER_18_184 ();
 sg13g2_decap_8 FILLER_18_193 ();
 sg13g2_decap_4 FILLER_18_200 ();
 sg13g2_fill_2 FILLER_18_204 ();
 sg13g2_fill_2 FILLER_18_235 ();
 sg13g2_fill_2 FILLER_18_272 ();
 sg13g2_fill_1 FILLER_18_274 ();
 sg13g2_fill_2 FILLER_18_280 ();
 sg13g2_fill_2 FILLER_18_361 ();
 sg13g2_fill_2 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_18_436 ();
 sg13g2_decap_8 FILLER_18_443 ();
 sg13g2_decap_4 FILLER_18_450 ();
 sg13g2_fill_1 FILLER_18_454 ();
 sg13g2_decap_4 FILLER_18_458 ();
 sg13g2_fill_1 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_471 ();
 sg13g2_decap_8 FILLER_18_478 ();
 sg13g2_decap_8 FILLER_18_485 ();
 sg13g2_decap_8 FILLER_18_492 ();
 sg13g2_decap_8 FILLER_18_499 ();
 sg13g2_decap_8 FILLER_18_506 ();
 sg13g2_decap_8 FILLER_18_513 ();
 sg13g2_decap_8 FILLER_18_520 ();
 sg13g2_decap_8 FILLER_18_527 ();
 sg13g2_decap_8 FILLER_18_534 ();
 sg13g2_decap_8 FILLER_18_541 ();
 sg13g2_decap_8 FILLER_18_548 ();
 sg13g2_decap_8 FILLER_18_555 ();
 sg13g2_decap_8 FILLER_18_562 ();
 sg13g2_decap_8 FILLER_18_569 ();
 sg13g2_decap_8 FILLER_18_576 ();
 sg13g2_decap_8 FILLER_18_583 ();
 sg13g2_decap_8 FILLER_18_590 ();
 sg13g2_decap_8 FILLER_18_597 ();
 sg13g2_decap_8 FILLER_18_604 ();
 sg13g2_decap_8 FILLER_18_611 ();
 sg13g2_decap_8 FILLER_18_618 ();
 sg13g2_decap_8 FILLER_18_625 ();
 sg13g2_decap_8 FILLER_18_632 ();
 sg13g2_decap_8 FILLER_18_639 ();
 sg13g2_decap_8 FILLER_18_646 ();
 sg13g2_decap_8 FILLER_18_653 ();
 sg13g2_decap_8 FILLER_18_660 ();
 sg13g2_decap_8 FILLER_18_667 ();
 sg13g2_decap_8 FILLER_18_674 ();
 sg13g2_decap_8 FILLER_18_681 ();
 sg13g2_decap_8 FILLER_18_688 ();
 sg13g2_decap_8 FILLER_18_695 ();
 sg13g2_decap_8 FILLER_18_702 ();
 sg13g2_decap_8 FILLER_18_709 ();
 sg13g2_decap_8 FILLER_18_716 ();
 sg13g2_decap_8 FILLER_18_723 ();
 sg13g2_decap_8 FILLER_18_730 ();
 sg13g2_decap_8 FILLER_18_737 ();
 sg13g2_decap_8 FILLER_18_744 ();
 sg13g2_decap_8 FILLER_18_751 ();
 sg13g2_decap_8 FILLER_18_758 ();
 sg13g2_decap_8 FILLER_18_765 ();
 sg13g2_decap_8 FILLER_18_772 ();
 sg13g2_decap_8 FILLER_18_779 ();
 sg13g2_decap_8 FILLER_18_786 ();
 sg13g2_decap_8 FILLER_18_793 ();
 sg13g2_decap_8 FILLER_18_800 ();
 sg13g2_decap_8 FILLER_18_807 ();
 sg13g2_decap_8 FILLER_18_814 ();
 sg13g2_decap_8 FILLER_18_821 ();
 sg13g2_decap_8 FILLER_18_828 ();
 sg13g2_decap_8 FILLER_18_835 ();
 sg13g2_decap_8 FILLER_18_842 ();
 sg13g2_decap_8 FILLER_18_849 ();
 sg13g2_decap_4 FILLER_18_856 ();
 sg13g2_fill_2 FILLER_18_860 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_fill_1 FILLER_19_86 ();
 sg13g2_fill_2 FILLER_19_130 ();
 sg13g2_fill_1 FILLER_19_132 ();
 sg13g2_fill_2 FILLER_19_150 ();
 sg13g2_fill_2 FILLER_19_161 ();
 sg13g2_fill_1 FILLER_19_206 ();
 sg13g2_fill_1 FILLER_19_211 ();
 sg13g2_fill_1 FILLER_19_261 ();
 sg13g2_fill_1 FILLER_19_267 ();
 sg13g2_fill_1 FILLER_19_321 ();
 sg13g2_fill_1 FILLER_19_366 ();
 sg13g2_fill_1 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_435 ();
 sg13g2_decap_4 FILLER_19_442 ();
 sg13g2_decap_8 FILLER_19_491 ();
 sg13g2_fill_2 FILLER_19_498 ();
 sg13g2_fill_1 FILLER_19_500 ();
 sg13g2_decap_8 FILLER_19_509 ();
 sg13g2_decap_8 FILLER_19_516 ();
 sg13g2_decap_8 FILLER_19_523 ();
 sg13g2_decap_8 FILLER_19_530 ();
 sg13g2_decap_8 FILLER_19_537 ();
 sg13g2_decap_8 FILLER_19_544 ();
 sg13g2_decap_8 FILLER_19_551 ();
 sg13g2_decap_8 FILLER_19_558 ();
 sg13g2_decap_8 FILLER_19_565 ();
 sg13g2_decap_8 FILLER_19_572 ();
 sg13g2_decap_8 FILLER_19_579 ();
 sg13g2_decap_8 FILLER_19_586 ();
 sg13g2_decap_8 FILLER_19_593 ();
 sg13g2_decap_8 FILLER_19_600 ();
 sg13g2_decap_8 FILLER_19_607 ();
 sg13g2_decap_8 FILLER_19_614 ();
 sg13g2_decap_8 FILLER_19_621 ();
 sg13g2_decap_8 FILLER_19_628 ();
 sg13g2_decap_8 FILLER_19_635 ();
 sg13g2_decap_8 FILLER_19_642 ();
 sg13g2_decap_8 FILLER_19_649 ();
 sg13g2_decap_8 FILLER_19_656 ();
 sg13g2_decap_8 FILLER_19_663 ();
 sg13g2_decap_8 FILLER_19_670 ();
 sg13g2_decap_8 FILLER_19_677 ();
 sg13g2_decap_8 FILLER_19_684 ();
 sg13g2_decap_8 FILLER_19_691 ();
 sg13g2_decap_8 FILLER_19_698 ();
 sg13g2_decap_8 FILLER_19_705 ();
 sg13g2_decap_8 FILLER_19_712 ();
 sg13g2_decap_8 FILLER_19_719 ();
 sg13g2_decap_8 FILLER_19_726 ();
 sg13g2_decap_8 FILLER_19_733 ();
 sg13g2_decap_8 FILLER_19_740 ();
 sg13g2_decap_8 FILLER_19_747 ();
 sg13g2_decap_8 FILLER_19_754 ();
 sg13g2_decap_8 FILLER_19_761 ();
 sg13g2_decap_8 FILLER_19_768 ();
 sg13g2_decap_8 FILLER_19_775 ();
 sg13g2_decap_8 FILLER_19_782 ();
 sg13g2_decap_8 FILLER_19_789 ();
 sg13g2_decap_8 FILLER_19_796 ();
 sg13g2_decap_8 FILLER_19_803 ();
 sg13g2_decap_8 FILLER_19_810 ();
 sg13g2_decap_8 FILLER_19_817 ();
 sg13g2_decap_8 FILLER_19_824 ();
 sg13g2_decap_8 FILLER_19_831 ();
 sg13g2_decap_8 FILLER_19_838 ();
 sg13g2_decap_8 FILLER_19_845 ();
 sg13g2_decap_8 FILLER_19_852 ();
 sg13g2_fill_2 FILLER_19_859 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_fill_1 FILLER_20_49 ();
 sg13g2_fill_2 FILLER_20_76 ();
 sg13g2_fill_1 FILLER_20_78 ();
 sg13g2_fill_2 FILLER_20_93 ();
 sg13g2_fill_2 FILLER_20_110 ();
 sg13g2_fill_1 FILLER_20_112 ();
 sg13g2_fill_2 FILLER_20_128 ();
 sg13g2_fill_2 FILLER_20_139 ();
 sg13g2_fill_1 FILLER_20_141 ();
 sg13g2_fill_1 FILLER_20_214 ();
 sg13g2_fill_2 FILLER_20_344 ();
 sg13g2_fill_1 FILLER_20_369 ();
 sg13g2_fill_2 FILLER_20_393 ();
 sg13g2_decap_4 FILLER_20_437 ();
 sg13g2_fill_2 FILLER_20_472 ();
 sg13g2_decap_8 FILLER_20_517 ();
 sg13g2_decap_8 FILLER_20_524 ();
 sg13g2_decap_4 FILLER_20_531 ();
 sg13g2_fill_1 FILLER_20_535 ();
 sg13g2_decap_4 FILLER_20_551 ();
 sg13g2_fill_1 FILLER_20_555 ();
 sg13g2_fill_2 FILLER_20_570 ();
 sg13g2_fill_1 FILLER_20_572 ();
 sg13g2_decap_8 FILLER_20_590 ();
 sg13g2_decap_8 FILLER_20_597 ();
 sg13g2_decap_8 FILLER_20_604 ();
 sg13g2_decap_8 FILLER_20_611 ();
 sg13g2_decap_8 FILLER_20_618 ();
 sg13g2_decap_8 FILLER_20_625 ();
 sg13g2_decap_8 FILLER_20_632 ();
 sg13g2_decap_8 FILLER_20_639 ();
 sg13g2_decap_8 FILLER_20_646 ();
 sg13g2_decap_8 FILLER_20_653 ();
 sg13g2_decap_8 FILLER_20_660 ();
 sg13g2_decap_8 FILLER_20_667 ();
 sg13g2_decap_8 FILLER_20_674 ();
 sg13g2_decap_8 FILLER_20_681 ();
 sg13g2_decap_8 FILLER_20_688 ();
 sg13g2_decap_8 FILLER_20_695 ();
 sg13g2_decap_8 FILLER_20_702 ();
 sg13g2_decap_8 FILLER_20_709 ();
 sg13g2_decap_8 FILLER_20_716 ();
 sg13g2_decap_8 FILLER_20_723 ();
 sg13g2_decap_8 FILLER_20_730 ();
 sg13g2_decap_8 FILLER_20_737 ();
 sg13g2_decap_8 FILLER_20_744 ();
 sg13g2_decap_8 FILLER_20_751 ();
 sg13g2_decap_8 FILLER_20_758 ();
 sg13g2_decap_8 FILLER_20_765 ();
 sg13g2_decap_8 FILLER_20_772 ();
 sg13g2_decap_8 FILLER_20_779 ();
 sg13g2_decap_8 FILLER_20_786 ();
 sg13g2_decap_8 FILLER_20_793 ();
 sg13g2_decap_8 FILLER_20_800 ();
 sg13g2_decap_8 FILLER_20_807 ();
 sg13g2_decap_8 FILLER_20_814 ();
 sg13g2_decap_8 FILLER_20_821 ();
 sg13g2_decap_8 FILLER_20_828 ();
 sg13g2_decap_8 FILLER_20_835 ();
 sg13g2_decap_8 FILLER_20_842 ();
 sg13g2_decap_8 FILLER_20_849 ();
 sg13g2_decap_4 FILLER_20_856 ();
 sg13g2_fill_2 FILLER_20_860 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_37 ();
 sg13g2_fill_2 FILLER_21_66 ();
 sg13g2_fill_1 FILLER_21_107 ();
 sg13g2_fill_1 FILLER_21_139 ();
 sg13g2_fill_1 FILLER_21_172 ();
 sg13g2_fill_1 FILLER_21_225 ();
 sg13g2_fill_1 FILLER_21_270 ();
 sg13g2_fill_2 FILLER_21_304 ();
 sg13g2_fill_2 FILLER_21_329 ();
 sg13g2_fill_1 FILLER_21_331 ();
 sg13g2_fill_1 FILLER_21_423 ();
 sg13g2_fill_1 FILLER_21_459 ();
 sg13g2_fill_2 FILLER_21_529 ();
 sg13g2_fill_2 FILLER_21_580 ();
 sg13g2_decap_8 FILLER_21_604 ();
 sg13g2_decap_8 FILLER_21_611 ();
 sg13g2_decap_8 FILLER_21_618 ();
 sg13g2_decap_8 FILLER_21_625 ();
 sg13g2_decap_8 FILLER_21_632 ();
 sg13g2_decap_8 FILLER_21_639 ();
 sg13g2_decap_8 FILLER_21_646 ();
 sg13g2_decap_8 FILLER_21_653 ();
 sg13g2_decap_8 FILLER_21_660 ();
 sg13g2_decap_8 FILLER_21_667 ();
 sg13g2_decap_8 FILLER_21_674 ();
 sg13g2_decap_8 FILLER_21_681 ();
 sg13g2_decap_8 FILLER_21_688 ();
 sg13g2_decap_8 FILLER_21_695 ();
 sg13g2_decap_8 FILLER_21_702 ();
 sg13g2_decap_8 FILLER_21_709 ();
 sg13g2_decap_8 FILLER_21_716 ();
 sg13g2_decap_8 FILLER_21_723 ();
 sg13g2_decap_8 FILLER_21_730 ();
 sg13g2_decap_8 FILLER_21_737 ();
 sg13g2_decap_8 FILLER_21_744 ();
 sg13g2_decap_8 FILLER_21_751 ();
 sg13g2_decap_8 FILLER_21_758 ();
 sg13g2_decap_8 FILLER_21_765 ();
 sg13g2_decap_8 FILLER_21_772 ();
 sg13g2_decap_8 FILLER_21_779 ();
 sg13g2_decap_8 FILLER_21_786 ();
 sg13g2_decap_8 FILLER_21_793 ();
 sg13g2_decap_8 FILLER_21_800 ();
 sg13g2_decap_8 FILLER_21_807 ();
 sg13g2_decap_8 FILLER_21_814 ();
 sg13g2_decap_8 FILLER_21_821 ();
 sg13g2_decap_8 FILLER_21_828 ();
 sg13g2_decap_8 FILLER_21_835 ();
 sg13g2_decap_8 FILLER_21_842 ();
 sg13g2_decap_8 FILLER_21_849 ();
 sg13g2_decap_4 FILLER_21_856 ();
 sg13g2_fill_2 FILLER_21_860 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_4 FILLER_22_21 ();
 sg13g2_fill_2 FILLER_22_89 ();
 sg13g2_fill_2 FILLER_22_138 ();
 sg13g2_fill_2 FILLER_22_166 ();
 sg13g2_fill_1 FILLER_22_168 ();
 sg13g2_fill_1 FILLER_22_237 ();
 sg13g2_fill_1 FILLER_22_252 ();
 sg13g2_fill_1 FILLER_22_293 ();
 sg13g2_fill_2 FILLER_22_343 ();
 sg13g2_decap_4 FILLER_22_359 ();
 sg13g2_fill_1 FILLER_22_363 ();
 sg13g2_fill_2 FILLER_22_430 ();
 sg13g2_fill_2 FILLER_22_478 ();
 sg13g2_fill_1 FILLER_22_523 ();
 sg13g2_decap_8 FILLER_22_612 ();
 sg13g2_decap_8 FILLER_22_619 ();
 sg13g2_decap_8 FILLER_22_626 ();
 sg13g2_decap_8 FILLER_22_633 ();
 sg13g2_decap_8 FILLER_22_640 ();
 sg13g2_decap_8 FILLER_22_647 ();
 sg13g2_decap_8 FILLER_22_654 ();
 sg13g2_decap_8 FILLER_22_661 ();
 sg13g2_decap_8 FILLER_22_668 ();
 sg13g2_decap_8 FILLER_22_675 ();
 sg13g2_decap_8 FILLER_22_682 ();
 sg13g2_decap_8 FILLER_22_689 ();
 sg13g2_decap_8 FILLER_22_696 ();
 sg13g2_decap_8 FILLER_22_703 ();
 sg13g2_decap_8 FILLER_22_710 ();
 sg13g2_decap_8 FILLER_22_717 ();
 sg13g2_decap_8 FILLER_22_724 ();
 sg13g2_decap_8 FILLER_22_731 ();
 sg13g2_decap_8 FILLER_22_738 ();
 sg13g2_decap_8 FILLER_22_745 ();
 sg13g2_decap_8 FILLER_22_752 ();
 sg13g2_decap_8 FILLER_22_759 ();
 sg13g2_decap_8 FILLER_22_766 ();
 sg13g2_decap_8 FILLER_22_773 ();
 sg13g2_decap_8 FILLER_22_780 ();
 sg13g2_decap_8 FILLER_22_787 ();
 sg13g2_decap_8 FILLER_22_794 ();
 sg13g2_decap_8 FILLER_22_801 ();
 sg13g2_decap_8 FILLER_22_808 ();
 sg13g2_decap_8 FILLER_22_815 ();
 sg13g2_decap_8 FILLER_22_822 ();
 sg13g2_decap_8 FILLER_22_829 ();
 sg13g2_decap_8 FILLER_22_836 ();
 sg13g2_decap_8 FILLER_22_843 ();
 sg13g2_decap_8 FILLER_22_850 ();
 sg13g2_decap_4 FILLER_22_857 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_4 FILLER_23_14 ();
 sg13g2_fill_1 FILLER_23_18 ();
 sg13g2_fill_1 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_95 ();
 sg13g2_fill_2 FILLER_23_101 ();
 sg13g2_fill_1 FILLER_23_103 ();
 sg13g2_fill_2 FILLER_23_109 ();
 sg13g2_fill_1 FILLER_23_281 ();
 sg13g2_decap_8 FILLER_23_352 ();
 sg13g2_fill_1 FILLER_23_359 ();
 sg13g2_decap_4 FILLER_23_365 ();
 sg13g2_fill_1 FILLER_23_373 ();
 sg13g2_fill_2 FILLER_23_383 ();
 sg13g2_decap_8 FILLER_23_408 ();
 sg13g2_fill_1 FILLER_23_428 ();
 sg13g2_fill_2 FILLER_23_525 ();
 sg13g2_fill_2 FILLER_23_540 ();
 sg13g2_fill_1 FILLER_23_597 ();
 sg13g2_decap_8 FILLER_23_615 ();
 sg13g2_decap_8 FILLER_23_622 ();
 sg13g2_decap_8 FILLER_23_629 ();
 sg13g2_decap_8 FILLER_23_636 ();
 sg13g2_decap_8 FILLER_23_643 ();
 sg13g2_decap_8 FILLER_23_650 ();
 sg13g2_decap_8 FILLER_23_657 ();
 sg13g2_decap_8 FILLER_23_664 ();
 sg13g2_decap_8 FILLER_23_671 ();
 sg13g2_decap_8 FILLER_23_678 ();
 sg13g2_decap_8 FILLER_23_685 ();
 sg13g2_decap_8 FILLER_23_692 ();
 sg13g2_decap_8 FILLER_23_699 ();
 sg13g2_decap_8 FILLER_23_706 ();
 sg13g2_decap_8 FILLER_23_713 ();
 sg13g2_decap_8 FILLER_23_720 ();
 sg13g2_decap_8 FILLER_23_727 ();
 sg13g2_decap_8 FILLER_23_734 ();
 sg13g2_decap_8 FILLER_23_741 ();
 sg13g2_decap_8 FILLER_23_748 ();
 sg13g2_decap_8 FILLER_23_755 ();
 sg13g2_decap_8 FILLER_23_762 ();
 sg13g2_decap_8 FILLER_23_769 ();
 sg13g2_decap_8 FILLER_23_776 ();
 sg13g2_decap_8 FILLER_23_783 ();
 sg13g2_decap_8 FILLER_23_790 ();
 sg13g2_decap_8 FILLER_23_797 ();
 sg13g2_decap_8 FILLER_23_804 ();
 sg13g2_decap_8 FILLER_23_811 ();
 sg13g2_decap_8 FILLER_23_818 ();
 sg13g2_decap_8 FILLER_23_825 ();
 sg13g2_decap_8 FILLER_23_832 ();
 sg13g2_decap_8 FILLER_23_839 ();
 sg13g2_decap_8 FILLER_23_846 ();
 sg13g2_decap_8 FILLER_23_853 ();
 sg13g2_fill_2 FILLER_23_860 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_99 ();
 sg13g2_fill_1 FILLER_24_101 ();
 sg13g2_fill_2 FILLER_24_141 ();
 sg13g2_fill_1 FILLER_24_143 ();
 sg13g2_fill_1 FILLER_24_159 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_fill_1 FILLER_24_207 ();
 sg13g2_fill_1 FILLER_24_267 ();
 sg13g2_fill_2 FILLER_24_301 ();
 sg13g2_fill_1 FILLER_24_308 ();
 sg13g2_fill_2 FILLER_24_318 ();
 sg13g2_fill_1 FILLER_24_324 ();
 sg13g2_fill_2 FILLER_24_333 ();
 sg13g2_fill_1 FILLER_24_335 ();
 sg13g2_decap_4 FILLER_24_340 ();
 sg13g2_fill_1 FILLER_24_344 ();
 sg13g2_decap_4 FILLER_24_351 ();
 sg13g2_fill_1 FILLER_24_355 ();
 sg13g2_decap_4 FILLER_24_373 ();
 sg13g2_fill_1 FILLER_24_377 ();
 sg13g2_fill_1 FILLER_24_390 ();
 sg13g2_fill_2 FILLER_24_396 ();
 sg13g2_fill_1 FILLER_24_403 ();
 sg13g2_decap_4 FILLER_24_408 ();
 sg13g2_fill_1 FILLER_24_412 ();
 sg13g2_decap_4 FILLER_24_427 ();
 sg13g2_fill_1 FILLER_24_431 ();
 sg13g2_fill_1 FILLER_24_437 ();
 sg13g2_fill_1 FILLER_24_520 ();
 sg13g2_decap_8 FILLER_24_622 ();
 sg13g2_decap_8 FILLER_24_629 ();
 sg13g2_decap_8 FILLER_24_636 ();
 sg13g2_decap_8 FILLER_24_643 ();
 sg13g2_decap_8 FILLER_24_650 ();
 sg13g2_decap_8 FILLER_24_657 ();
 sg13g2_decap_8 FILLER_24_664 ();
 sg13g2_decap_8 FILLER_24_671 ();
 sg13g2_decap_8 FILLER_24_678 ();
 sg13g2_decap_8 FILLER_24_685 ();
 sg13g2_decap_8 FILLER_24_692 ();
 sg13g2_decap_8 FILLER_24_699 ();
 sg13g2_decap_8 FILLER_24_706 ();
 sg13g2_decap_8 FILLER_24_713 ();
 sg13g2_decap_8 FILLER_24_720 ();
 sg13g2_decap_8 FILLER_24_727 ();
 sg13g2_decap_8 FILLER_24_734 ();
 sg13g2_decap_8 FILLER_24_741 ();
 sg13g2_decap_8 FILLER_24_748 ();
 sg13g2_decap_8 FILLER_24_755 ();
 sg13g2_decap_8 FILLER_24_762 ();
 sg13g2_decap_8 FILLER_24_769 ();
 sg13g2_decap_8 FILLER_24_776 ();
 sg13g2_decap_8 FILLER_24_783 ();
 sg13g2_decap_8 FILLER_24_790 ();
 sg13g2_decap_8 FILLER_24_797 ();
 sg13g2_decap_8 FILLER_24_804 ();
 sg13g2_decap_8 FILLER_24_811 ();
 sg13g2_decap_8 FILLER_24_818 ();
 sg13g2_decap_8 FILLER_24_825 ();
 sg13g2_decap_8 FILLER_24_832 ();
 sg13g2_decap_8 FILLER_24_839 ();
 sg13g2_decap_8 FILLER_24_846 ();
 sg13g2_decap_8 FILLER_24_853 ();
 sg13g2_fill_2 FILLER_24_860 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_2 ();
 sg13g2_fill_1 FILLER_25_52 ();
 sg13g2_fill_2 FILLER_25_70 ();
 sg13g2_fill_1 FILLER_25_129 ();
 sg13g2_fill_2 FILLER_25_197 ();
 sg13g2_fill_1 FILLER_25_244 ();
 sg13g2_fill_1 FILLER_25_284 ();
 sg13g2_fill_1 FILLER_25_297 ();
 sg13g2_fill_2 FILLER_25_313 ();
 sg13g2_fill_1 FILLER_25_315 ();
 sg13g2_decap_4 FILLER_25_331 ();
 sg13g2_fill_2 FILLER_25_335 ();
 sg13g2_fill_2 FILLER_25_350 ();
 sg13g2_fill_2 FILLER_25_394 ();
 sg13g2_fill_2 FILLER_25_427 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_25_437 ();
 sg13g2_fill_1 FILLER_25_444 ();
 sg13g2_fill_1 FILLER_25_491 ();
 sg13g2_fill_1 FILLER_25_528 ();
 sg13g2_fill_2 FILLER_25_547 ();
 sg13g2_fill_1 FILLER_25_589 ();
 sg13g2_decap_8 FILLER_25_616 ();
 sg13g2_decap_8 FILLER_25_623 ();
 sg13g2_decap_8 FILLER_25_630 ();
 sg13g2_decap_8 FILLER_25_637 ();
 sg13g2_decap_8 FILLER_25_644 ();
 sg13g2_decap_8 FILLER_25_651 ();
 sg13g2_decap_8 FILLER_25_658 ();
 sg13g2_decap_8 FILLER_25_665 ();
 sg13g2_decap_8 FILLER_25_672 ();
 sg13g2_decap_8 FILLER_25_679 ();
 sg13g2_decap_8 FILLER_25_686 ();
 sg13g2_decap_8 FILLER_25_693 ();
 sg13g2_decap_8 FILLER_25_700 ();
 sg13g2_decap_8 FILLER_25_707 ();
 sg13g2_decap_8 FILLER_25_714 ();
 sg13g2_decap_8 FILLER_25_721 ();
 sg13g2_decap_8 FILLER_25_728 ();
 sg13g2_decap_8 FILLER_25_735 ();
 sg13g2_decap_8 FILLER_25_742 ();
 sg13g2_decap_8 FILLER_25_749 ();
 sg13g2_decap_8 FILLER_25_756 ();
 sg13g2_decap_8 FILLER_25_763 ();
 sg13g2_decap_8 FILLER_25_770 ();
 sg13g2_decap_8 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_784 ();
 sg13g2_decap_8 FILLER_25_791 ();
 sg13g2_decap_8 FILLER_25_798 ();
 sg13g2_decap_8 FILLER_25_805 ();
 sg13g2_decap_8 FILLER_25_812 ();
 sg13g2_decap_8 FILLER_25_819 ();
 sg13g2_decap_8 FILLER_25_826 ();
 sg13g2_decap_8 FILLER_25_833 ();
 sg13g2_decap_8 FILLER_25_840 ();
 sg13g2_decap_8 FILLER_25_847 ();
 sg13g2_decap_8 FILLER_25_854 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_65 ();
 sg13g2_fill_1 FILLER_26_67 ();
 sg13g2_fill_2 FILLER_26_86 ();
 sg13g2_fill_1 FILLER_26_88 ();
 sg13g2_fill_2 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_208 ();
 sg13g2_fill_2 FILLER_26_223 ();
 sg13g2_fill_1 FILLER_26_291 ();
 sg13g2_fill_2 FILLER_26_307 ();
 sg13g2_fill_1 FILLER_26_309 ();
 sg13g2_fill_2 FILLER_26_328 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_fill_2 FILLER_26_411 ();
 sg13g2_fill_1 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_427 ();
 sg13g2_fill_2 FILLER_26_454 ();
 sg13g2_fill_1 FILLER_26_456 ();
 sg13g2_fill_2 FILLER_26_484 ();
 sg13g2_fill_2 FILLER_26_551 ();
 sg13g2_decap_8 FILLER_26_609 ();
 sg13g2_decap_8 FILLER_26_616 ();
 sg13g2_decap_8 FILLER_26_623 ();
 sg13g2_decap_8 FILLER_26_630 ();
 sg13g2_decap_8 FILLER_26_637 ();
 sg13g2_decap_8 FILLER_26_644 ();
 sg13g2_decap_8 FILLER_26_651 ();
 sg13g2_decap_8 FILLER_26_658 ();
 sg13g2_decap_8 FILLER_26_665 ();
 sg13g2_decap_8 FILLER_26_672 ();
 sg13g2_decap_8 FILLER_26_679 ();
 sg13g2_decap_8 FILLER_26_686 ();
 sg13g2_decap_8 FILLER_26_693 ();
 sg13g2_decap_8 FILLER_26_700 ();
 sg13g2_decap_8 FILLER_26_707 ();
 sg13g2_decap_8 FILLER_26_714 ();
 sg13g2_decap_8 FILLER_26_721 ();
 sg13g2_decap_8 FILLER_26_728 ();
 sg13g2_decap_8 FILLER_26_735 ();
 sg13g2_decap_8 FILLER_26_742 ();
 sg13g2_decap_8 FILLER_26_749 ();
 sg13g2_decap_8 FILLER_26_756 ();
 sg13g2_decap_8 FILLER_26_763 ();
 sg13g2_decap_8 FILLER_26_770 ();
 sg13g2_decap_8 FILLER_26_777 ();
 sg13g2_decap_8 FILLER_26_784 ();
 sg13g2_decap_8 FILLER_26_791 ();
 sg13g2_decap_8 FILLER_26_798 ();
 sg13g2_decap_8 FILLER_26_805 ();
 sg13g2_decap_8 FILLER_26_812 ();
 sg13g2_decap_8 FILLER_26_819 ();
 sg13g2_decap_8 FILLER_26_826 ();
 sg13g2_decap_8 FILLER_26_833 ();
 sg13g2_decap_8 FILLER_26_840 ();
 sg13g2_decap_8 FILLER_26_847 ();
 sg13g2_decap_8 FILLER_26_854 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_41 ();
 sg13g2_fill_2 FILLER_27_139 ();
 sg13g2_fill_1 FILLER_27_141 ();
 sg13g2_fill_1 FILLER_27_165 ();
 sg13g2_fill_1 FILLER_27_174 ();
 sg13g2_fill_2 FILLER_27_242 ();
 sg13g2_fill_2 FILLER_27_306 ();
 sg13g2_decap_4 FILLER_27_331 ();
 sg13g2_decap_8 FILLER_27_340 ();
 sg13g2_decap_4 FILLER_27_347 ();
 sg13g2_fill_1 FILLER_27_351 ();
 sg13g2_decap_8 FILLER_27_365 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_decap_4 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_4 FILLER_27_409 ();
 sg13g2_fill_1 FILLER_27_418 ();
 sg13g2_fill_1 FILLER_27_435 ();
 sg13g2_fill_2 FILLER_27_462 ();
 sg13g2_fill_2 FILLER_27_484 ();
 sg13g2_fill_2 FILLER_27_493 ();
 sg13g2_fill_1 FILLER_27_504 ();
 sg13g2_fill_1 FILLER_27_549 ();
 sg13g2_decap_8 FILLER_27_616 ();
 sg13g2_decap_8 FILLER_27_623 ();
 sg13g2_decap_8 FILLER_27_630 ();
 sg13g2_decap_8 FILLER_27_637 ();
 sg13g2_decap_8 FILLER_27_644 ();
 sg13g2_decap_8 FILLER_27_651 ();
 sg13g2_decap_8 FILLER_27_658 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_decap_8 FILLER_27_672 ();
 sg13g2_decap_8 FILLER_27_679 ();
 sg13g2_decap_8 FILLER_27_686 ();
 sg13g2_decap_8 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_700 ();
 sg13g2_decap_8 FILLER_27_707 ();
 sg13g2_decap_8 FILLER_27_714 ();
 sg13g2_decap_8 FILLER_27_721 ();
 sg13g2_decap_8 FILLER_27_728 ();
 sg13g2_decap_8 FILLER_27_735 ();
 sg13g2_decap_8 FILLER_27_742 ();
 sg13g2_decap_8 FILLER_27_749 ();
 sg13g2_decap_8 FILLER_27_756 ();
 sg13g2_decap_8 FILLER_27_763 ();
 sg13g2_decap_8 FILLER_27_770 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_decap_8 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_798 ();
 sg13g2_decap_8 FILLER_27_805 ();
 sg13g2_decap_8 FILLER_27_812 ();
 sg13g2_decap_8 FILLER_27_819 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_8 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_fill_1 FILLER_27_861 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_28 ();
 sg13g2_fill_1 FILLER_28_61 ();
 sg13g2_fill_2 FILLER_28_79 ();
 sg13g2_fill_1 FILLER_28_81 ();
 sg13g2_fill_1 FILLER_28_130 ();
 sg13g2_fill_1 FILLER_28_218 ();
 sg13g2_decap_4 FILLER_28_299 ();
 sg13g2_fill_1 FILLER_28_303 ();
 sg13g2_decap_8 FILLER_28_318 ();
 sg13g2_decap_8 FILLER_28_325 ();
 sg13g2_decap_4 FILLER_28_332 ();
 sg13g2_fill_1 FILLER_28_356 ();
 sg13g2_fill_2 FILLER_28_368 ();
 sg13g2_fill_1 FILLER_28_370 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_fill_1 FILLER_28_409 ();
 sg13g2_fill_2 FILLER_28_438 ();
 sg13g2_fill_1 FILLER_28_465 ();
 sg13g2_fill_1 FILLER_28_590 ();
 sg13g2_decap_8 FILLER_28_622 ();
 sg13g2_decap_8 FILLER_28_629 ();
 sg13g2_decap_8 FILLER_28_636 ();
 sg13g2_decap_8 FILLER_28_643 ();
 sg13g2_decap_8 FILLER_28_650 ();
 sg13g2_decap_8 FILLER_28_657 ();
 sg13g2_decap_8 FILLER_28_664 ();
 sg13g2_decap_8 FILLER_28_671 ();
 sg13g2_decap_8 FILLER_28_678 ();
 sg13g2_decap_8 FILLER_28_685 ();
 sg13g2_decap_8 FILLER_28_692 ();
 sg13g2_decap_8 FILLER_28_699 ();
 sg13g2_decap_8 FILLER_28_706 ();
 sg13g2_decap_8 FILLER_28_713 ();
 sg13g2_decap_8 FILLER_28_720 ();
 sg13g2_decap_8 FILLER_28_727 ();
 sg13g2_decap_8 FILLER_28_734 ();
 sg13g2_decap_8 FILLER_28_741 ();
 sg13g2_decap_8 FILLER_28_748 ();
 sg13g2_decap_8 FILLER_28_755 ();
 sg13g2_decap_8 FILLER_28_762 ();
 sg13g2_decap_8 FILLER_28_769 ();
 sg13g2_decap_8 FILLER_28_776 ();
 sg13g2_decap_8 FILLER_28_783 ();
 sg13g2_decap_8 FILLER_28_790 ();
 sg13g2_decap_8 FILLER_28_797 ();
 sg13g2_decap_8 FILLER_28_804 ();
 sg13g2_decap_8 FILLER_28_811 ();
 sg13g2_decap_8 FILLER_28_818 ();
 sg13g2_decap_8 FILLER_28_825 ();
 sg13g2_decap_8 FILLER_28_832 ();
 sg13g2_decap_8 FILLER_28_839 ();
 sg13g2_decap_8 FILLER_28_846 ();
 sg13g2_decap_8 FILLER_28_853 ();
 sg13g2_fill_2 FILLER_28_860 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_9 ();
 sg13g2_fill_1 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_97 ();
 sg13g2_fill_1 FILLER_29_103 ();
 sg13g2_fill_1 FILLER_29_132 ();
 sg13g2_fill_1 FILLER_29_138 ();
 sg13g2_fill_1 FILLER_29_144 ();
 sg13g2_fill_1 FILLER_29_150 ();
 sg13g2_fill_2 FILLER_29_177 ();
 sg13g2_fill_2 FILLER_29_233 ();
 sg13g2_fill_1 FILLER_29_253 ();
 sg13g2_fill_2 FILLER_29_280 ();
 sg13g2_fill_1 FILLER_29_298 ();
 sg13g2_fill_2 FILLER_29_353 ();
 sg13g2_fill_1 FILLER_29_355 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_decap_8 FILLER_29_408 ();
 sg13g2_fill_2 FILLER_29_424 ();
 sg13g2_fill_2 FILLER_29_436 ();
 sg13g2_fill_2 FILLER_29_441 ();
 sg13g2_fill_1 FILLER_29_448 ();
 sg13g2_fill_2 FILLER_29_454 ();
 sg13g2_fill_1 FILLER_29_456 ();
 sg13g2_decap_8 FILLER_29_616 ();
 sg13g2_decap_8 FILLER_29_623 ();
 sg13g2_decap_8 FILLER_29_630 ();
 sg13g2_decap_8 FILLER_29_637 ();
 sg13g2_decap_8 FILLER_29_644 ();
 sg13g2_decap_8 FILLER_29_651 ();
 sg13g2_decap_8 FILLER_29_658 ();
 sg13g2_decap_8 FILLER_29_665 ();
 sg13g2_decap_8 FILLER_29_672 ();
 sg13g2_decap_8 FILLER_29_679 ();
 sg13g2_decap_8 FILLER_29_686 ();
 sg13g2_decap_8 FILLER_29_693 ();
 sg13g2_decap_8 FILLER_29_700 ();
 sg13g2_decap_8 FILLER_29_707 ();
 sg13g2_decap_8 FILLER_29_714 ();
 sg13g2_decap_8 FILLER_29_721 ();
 sg13g2_decap_8 FILLER_29_728 ();
 sg13g2_decap_8 FILLER_29_735 ();
 sg13g2_decap_8 FILLER_29_742 ();
 sg13g2_decap_8 FILLER_29_749 ();
 sg13g2_decap_8 FILLER_29_756 ();
 sg13g2_decap_8 FILLER_29_763 ();
 sg13g2_decap_8 FILLER_29_770 ();
 sg13g2_decap_8 FILLER_29_777 ();
 sg13g2_decap_8 FILLER_29_784 ();
 sg13g2_decap_8 FILLER_29_791 ();
 sg13g2_decap_8 FILLER_29_798 ();
 sg13g2_decap_8 FILLER_29_805 ();
 sg13g2_decap_8 FILLER_29_812 ();
 sg13g2_decap_8 FILLER_29_819 ();
 sg13g2_decap_8 FILLER_29_826 ();
 sg13g2_decap_8 FILLER_29_833 ();
 sg13g2_decap_8 FILLER_29_840 ();
 sg13g2_decap_8 FILLER_29_847 ();
 sg13g2_decap_8 FILLER_29_854 ();
 sg13g2_fill_1 FILLER_29_861 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_4 FILLER_30_14 ();
 sg13g2_fill_1 FILLER_30_18 ();
 sg13g2_fill_2 FILLER_30_76 ();
 sg13g2_fill_2 FILLER_30_100 ();
 sg13g2_fill_2 FILLER_30_107 ();
 sg13g2_fill_1 FILLER_30_109 ();
 sg13g2_fill_1 FILLER_30_149 ();
 sg13g2_fill_1 FILLER_30_219 ();
 sg13g2_fill_2 FILLER_30_303 ();
 sg13g2_fill_1 FILLER_30_331 ();
 sg13g2_fill_2 FILLER_30_338 ();
 sg13g2_fill_1 FILLER_30_340 ();
 sg13g2_fill_2 FILLER_30_356 ();
 sg13g2_fill_1 FILLER_30_364 ();
 sg13g2_decap_4 FILLER_30_402 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_2 FILLER_30_422 ();
 sg13g2_fill_1 FILLER_30_424 ();
 sg13g2_decap_4 FILLER_30_432 ();
 sg13g2_fill_2 FILLER_30_465 ();
 sg13g2_fill_1 FILLER_30_474 ();
 sg13g2_fill_1 FILLER_30_503 ();
 sg13g2_fill_2 FILLER_30_527 ();
 sg13g2_fill_1 FILLER_30_538 ();
 sg13g2_fill_1 FILLER_30_561 ();
 sg13g2_fill_1 FILLER_30_571 ();
 sg13g2_fill_1 FILLER_30_603 ();
 sg13g2_decap_8 FILLER_30_617 ();
 sg13g2_decap_8 FILLER_30_624 ();
 sg13g2_decap_8 FILLER_30_631 ();
 sg13g2_decap_8 FILLER_30_638 ();
 sg13g2_decap_8 FILLER_30_645 ();
 sg13g2_decap_8 FILLER_30_652 ();
 sg13g2_decap_8 FILLER_30_659 ();
 sg13g2_decap_8 FILLER_30_666 ();
 sg13g2_decap_8 FILLER_30_673 ();
 sg13g2_decap_8 FILLER_30_680 ();
 sg13g2_decap_8 FILLER_30_687 ();
 sg13g2_decap_8 FILLER_30_694 ();
 sg13g2_decap_8 FILLER_30_701 ();
 sg13g2_decap_8 FILLER_30_708 ();
 sg13g2_decap_8 FILLER_30_715 ();
 sg13g2_decap_8 FILLER_30_722 ();
 sg13g2_decap_8 FILLER_30_729 ();
 sg13g2_decap_8 FILLER_30_736 ();
 sg13g2_decap_8 FILLER_30_743 ();
 sg13g2_decap_8 FILLER_30_750 ();
 sg13g2_decap_8 FILLER_30_757 ();
 sg13g2_decap_8 FILLER_30_764 ();
 sg13g2_decap_8 FILLER_30_771 ();
 sg13g2_decap_8 FILLER_30_778 ();
 sg13g2_decap_8 FILLER_30_785 ();
 sg13g2_decap_8 FILLER_30_792 ();
 sg13g2_decap_8 FILLER_30_799 ();
 sg13g2_decap_8 FILLER_30_806 ();
 sg13g2_decap_8 FILLER_30_813 ();
 sg13g2_decap_8 FILLER_30_820 ();
 sg13g2_decap_8 FILLER_30_827 ();
 sg13g2_decap_8 FILLER_30_834 ();
 sg13g2_decap_8 FILLER_30_841 ();
 sg13g2_decap_8 FILLER_30_848 ();
 sg13g2_decap_8 FILLER_30_855 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_11 ();
 sg13g2_fill_1 FILLER_31_46 ();
 sg13g2_fill_2 FILLER_31_79 ();
 sg13g2_fill_1 FILLER_31_81 ();
 sg13g2_decap_4 FILLER_31_113 ();
 sg13g2_fill_2 FILLER_31_117 ();
 sg13g2_fill_1 FILLER_31_152 ();
 sg13g2_fill_1 FILLER_31_166 ();
 sg13g2_fill_2 FILLER_31_195 ();
 sg13g2_fill_1 FILLER_31_215 ();
 sg13g2_fill_2 FILLER_31_229 ();
 sg13g2_fill_1 FILLER_31_316 ();
 sg13g2_fill_1 FILLER_31_327 ();
 sg13g2_fill_1 FILLER_31_364 ();
 sg13g2_fill_1 FILLER_31_384 ();
 sg13g2_decap_4 FILLER_31_411 ();
 sg13g2_fill_1 FILLER_31_441 ();
 sg13g2_fill_2 FILLER_31_451 ();
 sg13g2_fill_2 FILLER_31_509 ();
 sg13g2_decap_8 FILLER_31_608 ();
 sg13g2_decap_8 FILLER_31_615 ();
 sg13g2_decap_8 FILLER_31_622 ();
 sg13g2_decap_8 FILLER_31_629 ();
 sg13g2_decap_8 FILLER_31_636 ();
 sg13g2_decap_8 FILLER_31_643 ();
 sg13g2_decap_8 FILLER_31_650 ();
 sg13g2_decap_8 FILLER_31_657 ();
 sg13g2_decap_8 FILLER_31_664 ();
 sg13g2_decap_8 FILLER_31_671 ();
 sg13g2_decap_8 FILLER_31_678 ();
 sg13g2_decap_8 FILLER_31_685 ();
 sg13g2_decap_8 FILLER_31_692 ();
 sg13g2_decap_8 FILLER_31_699 ();
 sg13g2_decap_8 FILLER_31_706 ();
 sg13g2_decap_8 FILLER_31_713 ();
 sg13g2_decap_8 FILLER_31_720 ();
 sg13g2_decap_8 FILLER_31_727 ();
 sg13g2_decap_8 FILLER_31_734 ();
 sg13g2_decap_8 FILLER_31_741 ();
 sg13g2_decap_8 FILLER_31_748 ();
 sg13g2_decap_8 FILLER_31_755 ();
 sg13g2_decap_8 FILLER_31_762 ();
 sg13g2_decap_8 FILLER_31_769 ();
 sg13g2_decap_8 FILLER_31_776 ();
 sg13g2_decap_8 FILLER_31_783 ();
 sg13g2_decap_8 FILLER_31_790 ();
 sg13g2_decap_8 FILLER_31_797 ();
 sg13g2_decap_8 FILLER_31_804 ();
 sg13g2_decap_8 FILLER_31_811 ();
 sg13g2_decap_8 FILLER_31_818 ();
 sg13g2_decap_8 FILLER_31_825 ();
 sg13g2_decap_8 FILLER_31_832 ();
 sg13g2_decap_8 FILLER_31_839 ();
 sg13g2_decap_8 FILLER_31_846 ();
 sg13g2_decap_8 FILLER_31_853 ();
 sg13g2_fill_2 FILLER_31_860 ();
 sg13g2_fill_2 FILLER_32_31 ();
 sg13g2_fill_2 FILLER_32_59 ();
 sg13g2_fill_2 FILLER_32_76 ();
 sg13g2_fill_1 FILLER_32_78 ();
 sg13g2_fill_1 FILLER_32_89 ();
 sg13g2_fill_2 FILLER_32_94 ();
 sg13g2_decap_4 FILLER_32_106 ();
 sg13g2_fill_1 FILLER_32_115 ();
 sg13g2_fill_1 FILLER_32_129 ();
 sg13g2_fill_2 FILLER_32_148 ();
 sg13g2_fill_1 FILLER_32_150 ();
 sg13g2_fill_1 FILLER_32_324 ();
 sg13g2_decap_8 FILLER_32_334 ();
 sg13g2_decap_4 FILLER_32_341 ();
 sg13g2_fill_1 FILLER_32_345 ();
 sg13g2_fill_2 FILLER_32_365 ();
 sg13g2_fill_1 FILLER_32_403 ();
 sg13g2_decap_8 FILLER_32_418 ();
 sg13g2_fill_1 FILLER_32_425 ();
 sg13g2_fill_1 FILLER_32_430 ();
 sg13g2_fill_1 FILLER_32_546 ();
 sg13g2_fill_2 FILLER_32_580 ();
 sg13g2_fill_2 FILLER_32_591 ();
 sg13g2_decap_8 FILLER_32_615 ();
 sg13g2_decap_8 FILLER_32_622 ();
 sg13g2_decap_8 FILLER_32_629 ();
 sg13g2_decap_8 FILLER_32_636 ();
 sg13g2_decap_8 FILLER_32_643 ();
 sg13g2_decap_8 FILLER_32_650 ();
 sg13g2_decap_8 FILLER_32_657 ();
 sg13g2_decap_8 FILLER_32_664 ();
 sg13g2_decap_8 FILLER_32_671 ();
 sg13g2_decap_8 FILLER_32_678 ();
 sg13g2_decap_8 FILLER_32_685 ();
 sg13g2_decap_8 FILLER_32_692 ();
 sg13g2_decap_8 FILLER_32_699 ();
 sg13g2_decap_8 FILLER_32_706 ();
 sg13g2_decap_8 FILLER_32_713 ();
 sg13g2_decap_8 FILLER_32_720 ();
 sg13g2_decap_8 FILLER_32_727 ();
 sg13g2_decap_8 FILLER_32_734 ();
 sg13g2_decap_8 FILLER_32_741 ();
 sg13g2_decap_8 FILLER_32_748 ();
 sg13g2_decap_8 FILLER_32_755 ();
 sg13g2_decap_8 FILLER_32_762 ();
 sg13g2_decap_8 FILLER_32_769 ();
 sg13g2_decap_8 FILLER_32_776 ();
 sg13g2_decap_8 FILLER_32_783 ();
 sg13g2_decap_8 FILLER_32_790 ();
 sg13g2_decap_8 FILLER_32_797 ();
 sg13g2_decap_8 FILLER_32_804 ();
 sg13g2_decap_8 FILLER_32_811 ();
 sg13g2_decap_8 FILLER_32_818 ();
 sg13g2_decap_8 FILLER_32_825 ();
 sg13g2_decap_8 FILLER_32_832 ();
 sg13g2_decap_8 FILLER_32_839 ();
 sg13g2_decap_8 FILLER_32_846 ();
 sg13g2_decap_8 FILLER_32_853 ();
 sg13g2_fill_2 FILLER_32_860 ();
 sg13g2_fill_1 FILLER_33_40 ();
 sg13g2_fill_2 FILLER_33_50 ();
 sg13g2_fill_2 FILLER_33_61 ();
 sg13g2_fill_2 FILLER_33_76 ();
 sg13g2_decap_8 FILLER_33_101 ();
 sg13g2_decap_8 FILLER_33_108 ();
 sg13g2_fill_1 FILLER_33_115 ();
 sg13g2_fill_2 FILLER_33_127 ();
 sg13g2_fill_1 FILLER_33_129 ();
 sg13g2_fill_2 FILLER_33_134 ();
 sg13g2_fill_1 FILLER_33_144 ();
 sg13g2_fill_1 FILLER_33_184 ();
 sg13g2_fill_1 FILLER_33_216 ();
 sg13g2_fill_1 FILLER_33_237 ();
 sg13g2_fill_2 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_fill_2 FILLER_33_341 ();
 sg13g2_fill_1 FILLER_33_343 ();
 sg13g2_fill_2 FILLER_33_357 ();
 sg13g2_fill_2 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_33_434 ();
 sg13g2_fill_1 FILLER_33_479 ();
 sg13g2_fill_2 FILLER_33_506 ();
 sg13g2_fill_2 FILLER_33_552 ();
 sg13g2_fill_2 FILLER_33_580 ();
 sg13g2_fill_1 FILLER_33_582 ();
 sg13g2_fill_1 FILLER_33_592 ();
 sg13g2_fill_2 FILLER_33_603 ();
 sg13g2_decap_8 FILLER_33_618 ();
 sg13g2_decap_8 FILLER_33_625 ();
 sg13g2_decap_8 FILLER_33_632 ();
 sg13g2_decap_8 FILLER_33_639 ();
 sg13g2_decap_8 FILLER_33_646 ();
 sg13g2_decap_8 FILLER_33_653 ();
 sg13g2_decap_8 FILLER_33_660 ();
 sg13g2_decap_8 FILLER_33_667 ();
 sg13g2_decap_8 FILLER_33_674 ();
 sg13g2_decap_8 FILLER_33_681 ();
 sg13g2_decap_8 FILLER_33_688 ();
 sg13g2_decap_8 FILLER_33_695 ();
 sg13g2_decap_8 FILLER_33_702 ();
 sg13g2_decap_8 FILLER_33_709 ();
 sg13g2_decap_8 FILLER_33_716 ();
 sg13g2_decap_8 FILLER_33_723 ();
 sg13g2_decap_8 FILLER_33_730 ();
 sg13g2_decap_8 FILLER_33_737 ();
 sg13g2_decap_8 FILLER_33_744 ();
 sg13g2_decap_8 FILLER_33_751 ();
 sg13g2_decap_8 FILLER_33_758 ();
 sg13g2_decap_8 FILLER_33_765 ();
 sg13g2_decap_8 FILLER_33_772 ();
 sg13g2_decap_8 FILLER_33_779 ();
 sg13g2_decap_8 FILLER_33_786 ();
 sg13g2_decap_8 FILLER_33_793 ();
 sg13g2_decap_8 FILLER_33_800 ();
 sg13g2_decap_8 FILLER_33_807 ();
 sg13g2_decap_8 FILLER_33_814 ();
 sg13g2_decap_8 FILLER_33_821 ();
 sg13g2_decap_8 FILLER_33_828 ();
 sg13g2_decap_8 FILLER_33_835 ();
 sg13g2_decap_8 FILLER_33_842 ();
 sg13g2_decap_8 FILLER_33_849 ();
 sg13g2_decap_4 FILLER_33_856 ();
 sg13g2_fill_2 FILLER_33_860 ();
 sg13g2_fill_1 FILLER_34_72 ();
 sg13g2_decap_8 FILLER_34_104 ();
 sg13g2_fill_2 FILLER_34_122 ();
 sg13g2_fill_2 FILLER_34_144 ();
 sg13g2_fill_2 FILLER_34_186 ();
 sg13g2_fill_1 FILLER_34_215 ();
 sg13g2_fill_2 FILLER_34_226 ();
 sg13g2_fill_2 FILLER_34_243 ();
 sg13g2_fill_1 FILLER_34_267 ();
 sg13g2_fill_2 FILLER_34_277 ();
 sg13g2_fill_1 FILLER_34_329 ();
 sg13g2_fill_2 FILLER_34_376 ();
 sg13g2_fill_1 FILLER_34_435 ();
 sg13g2_fill_1 FILLER_34_444 ();
 sg13g2_fill_2 FILLER_34_464 ();
 sg13g2_fill_2 FILLER_34_503 ();
 sg13g2_fill_2 FILLER_34_532 ();
 sg13g2_fill_1 FILLER_34_559 ();
 sg13g2_fill_2 FILLER_34_579 ();
 sg13g2_decap_8 FILLER_34_621 ();
 sg13g2_decap_8 FILLER_34_628 ();
 sg13g2_decap_8 FILLER_34_635 ();
 sg13g2_decap_8 FILLER_34_642 ();
 sg13g2_decap_8 FILLER_34_649 ();
 sg13g2_decap_8 FILLER_34_656 ();
 sg13g2_decap_8 FILLER_34_663 ();
 sg13g2_decap_8 FILLER_34_670 ();
 sg13g2_decap_8 FILLER_34_677 ();
 sg13g2_decap_8 FILLER_34_684 ();
 sg13g2_decap_8 FILLER_34_691 ();
 sg13g2_decap_8 FILLER_34_698 ();
 sg13g2_decap_8 FILLER_34_705 ();
 sg13g2_decap_8 FILLER_34_712 ();
 sg13g2_decap_8 FILLER_34_719 ();
 sg13g2_decap_8 FILLER_34_726 ();
 sg13g2_decap_8 FILLER_34_733 ();
 sg13g2_decap_8 FILLER_34_740 ();
 sg13g2_decap_8 FILLER_34_747 ();
 sg13g2_decap_8 FILLER_34_754 ();
 sg13g2_decap_8 FILLER_34_761 ();
 sg13g2_decap_8 FILLER_34_768 ();
 sg13g2_decap_8 FILLER_34_775 ();
 sg13g2_decap_8 FILLER_34_782 ();
 sg13g2_decap_8 FILLER_34_789 ();
 sg13g2_decap_8 FILLER_34_796 ();
 sg13g2_decap_8 FILLER_34_803 ();
 sg13g2_decap_8 FILLER_34_810 ();
 sg13g2_decap_8 FILLER_34_817 ();
 sg13g2_decap_8 FILLER_34_824 ();
 sg13g2_decap_8 FILLER_34_831 ();
 sg13g2_decap_8 FILLER_34_838 ();
 sg13g2_decap_8 FILLER_34_845 ();
 sg13g2_decap_8 FILLER_34_852 ();
 sg13g2_fill_2 FILLER_34_859 ();
 sg13g2_fill_1 FILLER_34_861 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_37 ();
 sg13g2_fill_1 FILLER_35_63 ();
 sg13g2_fill_2 FILLER_35_68 ();
 sg13g2_fill_1 FILLER_35_70 ();
 sg13g2_fill_1 FILLER_35_80 ();
 sg13g2_fill_2 FILLER_35_108 ();
 sg13g2_fill_1 FILLER_35_134 ();
 sg13g2_fill_1 FILLER_35_154 ();
 sg13g2_fill_2 FILLER_35_168 ();
 sg13g2_fill_1 FILLER_35_178 ();
 sg13g2_fill_2 FILLER_35_273 ();
 sg13g2_fill_1 FILLER_35_301 ();
 sg13g2_fill_2 FILLER_35_307 ();
 sg13g2_fill_1 FILLER_35_347 ();
 sg13g2_fill_2 FILLER_35_376 ();
 sg13g2_fill_2 FILLER_35_392 ();
 sg13g2_fill_2 FILLER_35_433 ();
 sg13g2_fill_1 FILLER_35_435 ();
 sg13g2_fill_1 FILLER_35_471 ();
 sg13g2_fill_2 FILLER_35_533 ();
 sg13g2_fill_2 FILLER_35_570 ();
 sg13g2_fill_2 FILLER_35_606 ();
 sg13g2_fill_1 FILLER_35_608 ();
 sg13g2_decap_8 FILLER_35_631 ();
 sg13g2_decap_8 FILLER_35_638 ();
 sg13g2_decap_8 FILLER_35_645 ();
 sg13g2_decap_8 FILLER_35_652 ();
 sg13g2_decap_8 FILLER_35_659 ();
 sg13g2_decap_8 FILLER_35_666 ();
 sg13g2_decap_8 FILLER_35_673 ();
 sg13g2_decap_8 FILLER_35_680 ();
 sg13g2_decap_8 FILLER_35_687 ();
 sg13g2_decap_8 FILLER_35_694 ();
 sg13g2_decap_8 FILLER_35_701 ();
 sg13g2_decap_8 FILLER_35_708 ();
 sg13g2_decap_8 FILLER_35_715 ();
 sg13g2_decap_8 FILLER_35_722 ();
 sg13g2_decap_8 FILLER_35_729 ();
 sg13g2_decap_8 FILLER_35_736 ();
 sg13g2_decap_8 FILLER_35_743 ();
 sg13g2_decap_8 FILLER_35_750 ();
 sg13g2_decap_8 FILLER_35_757 ();
 sg13g2_decap_8 FILLER_35_764 ();
 sg13g2_decap_8 FILLER_35_771 ();
 sg13g2_decap_8 FILLER_35_778 ();
 sg13g2_decap_8 FILLER_35_785 ();
 sg13g2_decap_8 FILLER_35_792 ();
 sg13g2_decap_8 FILLER_35_799 ();
 sg13g2_decap_8 FILLER_35_806 ();
 sg13g2_decap_8 FILLER_35_813 ();
 sg13g2_decap_8 FILLER_35_820 ();
 sg13g2_decap_8 FILLER_35_827 ();
 sg13g2_decap_8 FILLER_35_834 ();
 sg13g2_decap_8 FILLER_35_841 ();
 sg13g2_decap_8 FILLER_35_848 ();
 sg13g2_decap_8 FILLER_35_855 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_41 ();
 sg13g2_fill_2 FILLER_36_57 ();
 sg13g2_fill_1 FILLER_36_59 ();
 sg13g2_fill_1 FILLER_36_86 ();
 sg13g2_fill_2 FILLER_36_104 ();
 sg13g2_fill_1 FILLER_36_106 ();
 sg13g2_fill_2 FILLER_36_130 ();
 sg13g2_fill_1 FILLER_36_149 ();
 sg13g2_fill_2 FILLER_36_187 ();
 sg13g2_fill_1 FILLER_36_189 ();
 sg13g2_fill_1 FILLER_36_216 ();
 sg13g2_fill_2 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_262 ();
 sg13g2_fill_2 FILLER_36_375 ();
 sg13g2_fill_2 FILLER_36_417 ();
 sg13g2_fill_1 FILLER_36_424 ();
 sg13g2_fill_1 FILLER_36_443 ();
 sg13g2_fill_2 FILLER_36_530 ();
 sg13g2_fill_2 FILLER_36_562 ();
 sg13g2_decap_8 FILLER_36_634 ();
 sg13g2_decap_8 FILLER_36_641 ();
 sg13g2_decap_8 FILLER_36_648 ();
 sg13g2_decap_8 FILLER_36_655 ();
 sg13g2_decap_8 FILLER_36_662 ();
 sg13g2_decap_8 FILLER_36_669 ();
 sg13g2_decap_8 FILLER_36_676 ();
 sg13g2_decap_8 FILLER_36_683 ();
 sg13g2_decap_8 FILLER_36_690 ();
 sg13g2_decap_8 FILLER_36_697 ();
 sg13g2_decap_8 FILLER_36_704 ();
 sg13g2_decap_8 FILLER_36_711 ();
 sg13g2_decap_8 FILLER_36_718 ();
 sg13g2_decap_8 FILLER_36_725 ();
 sg13g2_decap_8 FILLER_36_732 ();
 sg13g2_decap_8 FILLER_36_739 ();
 sg13g2_decap_8 FILLER_36_746 ();
 sg13g2_decap_8 FILLER_36_753 ();
 sg13g2_decap_8 FILLER_36_760 ();
 sg13g2_decap_8 FILLER_36_767 ();
 sg13g2_decap_8 FILLER_36_774 ();
 sg13g2_decap_8 FILLER_36_781 ();
 sg13g2_decap_8 FILLER_36_788 ();
 sg13g2_decap_8 FILLER_36_795 ();
 sg13g2_decap_8 FILLER_36_802 ();
 sg13g2_decap_8 FILLER_36_809 ();
 sg13g2_decap_8 FILLER_36_816 ();
 sg13g2_decap_8 FILLER_36_823 ();
 sg13g2_decap_8 FILLER_36_830 ();
 sg13g2_decap_8 FILLER_36_837 ();
 sg13g2_decap_8 FILLER_36_844 ();
 sg13g2_decap_8 FILLER_36_851 ();
 sg13g2_decap_4 FILLER_36_858 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_4 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_15 ();
 sg13g2_fill_1 FILLER_37_45 ();
 sg13g2_fill_1 FILLER_37_60 ();
 sg13g2_fill_1 FILLER_37_65 ();
 sg13g2_fill_1 FILLER_37_97 ();
 sg13g2_decap_4 FILLER_37_102 ();
 sg13g2_fill_1 FILLER_37_110 ();
 sg13g2_fill_2 FILLER_37_119 ();
 sg13g2_fill_2 FILLER_37_125 ();
 sg13g2_fill_1 FILLER_37_127 ();
 sg13g2_fill_1 FILLER_37_163 ();
 sg13g2_fill_2 FILLER_37_190 ();
 sg13g2_fill_1 FILLER_37_192 ();
 sg13g2_fill_2 FILLER_37_339 ();
 sg13g2_fill_2 FILLER_37_367 ();
 sg13g2_fill_1 FILLER_37_455 ();
 sg13g2_fill_1 FILLER_37_521 ();
 sg13g2_fill_2 FILLER_37_584 ();
 sg13g2_fill_1 FILLER_37_600 ();
 sg13g2_fill_1 FILLER_37_622 ();
 sg13g2_decap_8 FILLER_37_636 ();
 sg13g2_decap_8 FILLER_37_643 ();
 sg13g2_decap_8 FILLER_37_650 ();
 sg13g2_decap_8 FILLER_37_657 ();
 sg13g2_decap_8 FILLER_37_664 ();
 sg13g2_decap_8 FILLER_37_671 ();
 sg13g2_decap_8 FILLER_37_678 ();
 sg13g2_decap_8 FILLER_37_685 ();
 sg13g2_decap_8 FILLER_37_692 ();
 sg13g2_decap_8 FILLER_37_699 ();
 sg13g2_decap_8 FILLER_37_706 ();
 sg13g2_decap_8 FILLER_37_713 ();
 sg13g2_decap_8 FILLER_37_720 ();
 sg13g2_decap_8 FILLER_37_727 ();
 sg13g2_decap_8 FILLER_37_734 ();
 sg13g2_decap_8 FILLER_37_741 ();
 sg13g2_decap_8 FILLER_37_748 ();
 sg13g2_decap_8 FILLER_37_755 ();
 sg13g2_decap_8 FILLER_37_762 ();
 sg13g2_decap_8 FILLER_37_769 ();
 sg13g2_decap_8 FILLER_37_776 ();
 sg13g2_decap_8 FILLER_37_783 ();
 sg13g2_decap_8 FILLER_37_790 ();
 sg13g2_decap_8 FILLER_37_797 ();
 sg13g2_decap_8 FILLER_37_804 ();
 sg13g2_decap_8 FILLER_37_811 ();
 sg13g2_decap_8 FILLER_37_818 ();
 sg13g2_decap_8 FILLER_37_825 ();
 sg13g2_decap_8 FILLER_37_832 ();
 sg13g2_decap_8 FILLER_37_839 ();
 sg13g2_decap_8 FILLER_37_846 ();
 sg13g2_decap_8 FILLER_37_853 ();
 sg13g2_fill_2 FILLER_37_860 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_fill_2 FILLER_38_28 ();
 sg13g2_fill_1 FILLER_38_30 ();
 sg13g2_fill_1 FILLER_38_57 ();
 sg13g2_fill_1 FILLER_38_84 ();
 sg13g2_fill_1 FILLER_38_94 ();
 sg13g2_decap_4 FILLER_38_121 ();
 sg13g2_fill_1 FILLER_38_125 ();
 sg13g2_fill_2 FILLER_38_158 ();
 sg13g2_fill_1 FILLER_38_160 ();
 sg13g2_fill_1 FILLER_38_225 ();
 sg13g2_fill_2 FILLER_38_265 ();
 sg13g2_fill_1 FILLER_38_402 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_fill_2 FILLER_38_426 ();
 sg13g2_decap_8 FILLER_38_442 ();
 sg13g2_fill_2 FILLER_38_449 ();
 sg13g2_fill_2 FILLER_38_495 ();
 sg13g2_fill_1 FILLER_38_497 ();
 sg13g2_fill_1 FILLER_38_575 ();
 sg13g2_decap_8 FILLER_38_637 ();
 sg13g2_decap_8 FILLER_38_644 ();
 sg13g2_decap_8 FILLER_38_651 ();
 sg13g2_decap_8 FILLER_38_658 ();
 sg13g2_decap_8 FILLER_38_665 ();
 sg13g2_decap_8 FILLER_38_672 ();
 sg13g2_decap_8 FILLER_38_679 ();
 sg13g2_decap_8 FILLER_38_686 ();
 sg13g2_decap_8 FILLER_38_693 ();
 sg13g2_decap_8 FILLER_38_700 ();
 sg13g2_decap_8 FILLER_38_707 ();
 sg13g2_decap_8 FILLER_38_714 ();
 sg13g2_decap_8 FILLER_38_721 ();
 sg13g2_decap_8 FILLER_38_728 ();
 sg13g2_decap_8 FILLER_38_735 ();
 sg13g2_decap_8 FILLER_38_742 ();
 sg13g2_decap_8 FILLER_38_749 ();
 sg13g2_decap_8 FILLER_38_756 ();
 sg13g2_decap_8 FILLER_38_763 ();
 sg13g2_decap_8 FILLER_38_770 ();
 sg13g2_decap_8 FILLER_38_777 ();
 sg13g2_decap_8 FILLER_38_784 ();
 sg13g2_decap_8 FILLER_38_791 ();
 sg13g2_decap_8 FILLER_38_798 ();
 sg13g2_decap_8 FILLER_38_805 ();
 sg13g2_decap_8 FILLER_38_812 ();
 sg13g2_decap_8 FILLER_38_819 ();
 sg13g2_decap_8 FILLER_38_826 ();
 sg13g2_decap_8 FILLER_38_833 ();
 sg13g2_decap_8 FILLER_38_840 ();
 sg13g2_decap_8 FILLER_38_847 ();
 sg13g2_decap_8 FILLER_38_854 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_46 ();
 sg13g2_decap_8 FILLER_39_53 ();
 sg13g2_decap_8 FILLER_39_60 ();
 sg13g2_fill_2 FILLER_39_67 ();
 sg13g2_decap_8 FILLER_39_73 ();
 sg13g2_decap_8 FILLER_39_80 ();
 sg13g2_fill_1 FILLER_39_87 ();
 sg13g2_fill_1 FILLER_39_93 ();
 sg13g2_fill_1 FILLER_39_103 ();
 sg13g2_decap_8 FILLER_39_117 ();
 sg13g2_fill_2 FILLER_39_124 ();
 sg13g2_fill_1 FILLER_39_126 ();
 sg13g2_fill_1 FILLER_39_131 ();
 sg13g2_fill_1 FILLER_39_160 ();
 sg13g2_decap_4 FILLER_39_188 ();
 sg13g2_fill_2 FILLER_39_192 ();
 sg13g2_fill_1 FILLER_39_258 ();
 sg13g2_fill_2 FILLER_39_310 ();
 sg13g2_fill_2 FILLER_39_347 ();
 sg13g2_fill_2 FILLER_39_426 ();
 sg13g2_fill_1 FILLER_39_454 ();
 sg13g2_fill_2 FILLER_39_496 ();
 sg13g2_fill_1 FILLER_39_498 ();
 sg13g2_fill_2 FILLER_39_512 ();
 sg13g2_fill_2 FILLER_39_530 ();
 sg13g2_fill_2 FILLER_39_585 ();
 sg13g2_fill_1 FILLER_39_601 ();
 sg13g2_decap_8 FILLER_39_636 ();
 sg13g2_decap_8 FILLER_39_643 ();
 sg13g2_decap_8 FILLER_39_650 ();
 sg13g2_decap_8 FILLER_39_657 ();
 sg13g2_decap_8 FILLER_39_664 ();
 sg13g2_decap_8 FILLER_39_671 ();
 sg13g2_decap_8 FILLER_39_678 ();
 sg13g2_decap_8 FILLER_39_685 ();
 sg13g2_decap_8 FILLER_39_692 ();
 sg13g2_decap_8 FILLER_39_699 ();
 sg13g2_decap_8 FILLER_39_706 ();
 sg13g2_decap_8 FILLER_39_713 ();
 sg13g2_decap_8 FILLER_39_720 ();
 sg13g2_decap_8 FILLER_39_727 ();
 sg13g2_decap_8 FILLER_39_734 ();
 sg13g2_decap_8 FILLER_39_741 ();
 sg13g2_decap_8 FILLER_39_748 ();
 sg13g2_decap_8 FILLER_39_755 ();
 sg13g2_decap_8 FILLER_39_762 ();
 sg13g2_decap_8 FILLER_39_769 ();
 sg13g2_decap_8 FILLER_39_776 ();
 sg13g2_decap_8 FILLER_39_783 ();
 sg13g2_decap_8 FILLER_39_790 ();
 sg13g2_decap_8 FILLER_39_797 ();
 sg13g2_decap_8 FILLER_39_804 ();
 sg13g2_decap_8 FILLER_39_811 ();
 sg13g2_decap_8 FILLER_39_818 ();
 sg13g2_decap_8 FILLER_39_825 ();
 sg13g2_decap_8 FILLER_39_832 ();
 sg13g2_decap_8 FILLER_39_839 ();
 sg13g2_decap_8 FILLER_39_846 ();
 sg13g2_decap_8 FILLER_39_853 ();
 sg13g2_fill_2 FILLER_39_860 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_fill_2 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_97 ();
 sg13g2_decap_8 FILLER_40_104 ();
 sg13g2_decap_4 FILLER_40_111 ();
 sg13g2_fill_1 FILLER_40_115 ();
 sg13g2_fill_2 FILLER_40_155 ();
 sg13g2_decap_4 FILLER_40_197 ();
 sg13g2_fill_2 FILLER_40_201 ();
 sg13g2_fill_1 FILLER_40_306 ();
 sg13g2_fill_2 FILLER_40_328 ();
 sg13g2_fill_2 FILLER_40_388 ();
 sg13g2_fill_1 FILLER_40_390 ();
 sg13g2_fill_1 FILLER_40_403 ();
 sg13g2_fill_2 FILLER_40_413 ();
 sg13g2_fill_2 FILLER_40_474 ();
 sg13g2_decap_8 FILLER_40_488 ();
 sg13g2_fill_2 FILLER_40_495 ();
 sg13g2_fill_1 FILLER_40_497 ();
 sg13g2_fill_2 FILLER_40_554 ();
 sg13g2_fill_2 FILLER_40_582 ();
 sg13g2_fill_1 FILLER_40_584 ();
 sg13g2_decap_8 FILLER_40_637 ();
 sg13g2_decap_8 FILLER_40_644 ();
 sg13g2_decap_8 FILLER_40_651 ();
 sg13g2_decap_8 FILLER_40_658 ();
 sg13g2_decap_8 FILLER_40_665 ();
 sg13g2_decap_8 FILLER_40_672 ();
 sg13g2_decap_8 FILLER_40_679 ();
 sg13g2_decap_8 FILLER_40_686 ();
 sg13g2_decap_8 FILLER_40_693 ();
 sg13g2_decap_8 FILLER_40_700 ();
 sg13g2_decap_8 FILLER_40_707 ();
 sg13g2_decap_8 FILLER_40_714 ();
 sg13g2_decap_8 FILLER_40_721 ();
 sg13g2_decap_8 FILLER_40_728 ();
 sg13g2_decap_8 FILLER_40_735 ();
 sg13g2_decap_8 FILLER_40_742 ();
 sg13g2_decap_8 FILLER_40_749 ();
 sg13g2_decap_8 FILLER_40_756 ();
 sg13g2_decap_8 FILLER_40_763 ();
 sg13g2_decap_8 FILLER_40_770 ();
 sg13g2_decap_8 FILLER_40_777 ();
 sg13g2_decap_8 FILLER_40_784 ();
 sg13g2_decap_8 FILLER_40_791 ();
 sg13g2_decap_8 FILLER_40_798 ();
 sg13g2_decap_8 FILLER_40_805 ();
 sg13g2_decap_8 FILLER_40_812 ();
 sg13g2_decap_8 FILLER_40_819 ();
 sg13g2_decap_8 FILLER_40_826 ();
 sg13g2_decap_8 FILLER_40_833 ();
 sg13g2_decap_8 FILLER_40_840 ();
 sg13g2_decap_8 FILLER_40_847 ();
 sg13g2_decap_8 FILLER_40_854 ();
 sg13g2_fill_1 FILLER_40_861 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_fill_1 FILLER_41_133 ();
 sg13g2_fill_2 FILLER_41_155 ();
 sg13g2_fill_1 FILLER_41_157 ();
 sg13g2_fill_2 FILLER_41_167 ();
 sg13g2_decap_8 FILLER_41_195 ();
 sg13g2_decap_8 FILLER_41_202 ();
 sg13g2_fill_2 FILLER_41_209 ();
 sg13g2_fill_1 FILLER_41_211 ();
 sg13g2_fill_1 FILLER_41_221 ();
 sg13g2_decap_4 FILLER_41_235 ();
 sg13g2_fill_1 FILLER_41_278 ();
 sg13g2_fill_2 FILLER_41_309 ();
 sg13g2_fill_1 FILLER_41_321 ();
 sg13g2_decap_4 FILLER_41_345 ();
 sg13g2_fill_1 FILLER_41_349 ();
 sg13g2_fill_1 FILLER_41_422 ();
 sg13g2_fill_1 FILLER_41_438 ();
 sg13g2_fill_1 FILLER_41_448 ();
 sg13g2_decap_4 FILLER_41_462 ();
 sg13g2_fill_2 FILLER_41_466 ();
 sg13g2_fill_1 FILLER_41_511 ();
 sg13g2_fill_1 FILLER_41_549 ();
 sg13g2_fill_2 FILLER_41_562 ();
 sg13g2_fill_1 FILLER_41_564 ();
 sg13g2_decap_8 FILLER_41_626 ();
 sg13g2_decap_8 FILLER_41_633 ();
 sg13g2_decap_8 FILLER_41_640 ();
 sg13g2_decap_8 FILLER_41_647 ();
 sg13g2_decap_8 FILLER_41_654 ();
 sg13g2_decap_8 FILLER_41_661 ();
 sg13g2_decap_8 FILLER_41_668 ();
 sg13g2_decap_8 FILLER_41_675 ();
 sg13g2_decap_8 FILLER_41_682 ();
 sg13g2_decap_8 FILLER_41_689 ();
 sg13g2_decap_8 FILLER_41_696 ();
 sg13g2_decap_8 FILLER_41_703 ();
 sg13g2_decap_8 FILLER_41_710 ();
 sg13g2_decap_8 FILLER_41_717 ();
 sg13g2_decap_8 FILLER_41_724 ();
 sg13g2_decap_8 FILLER_41_731 ();
 sg13g2_decap_8 FILLER_41_738 ();
 sg13g2_decap_8 FILLER_41_745 ();
 sg13g2_decap_8 FILLER_41_752 ();
 sg13g2_decap_8 FILLER_41_759 ();
 sg13g2_decap_8 FILLER_41_766 ();
 sg13g2_decap_8 FILLER_41_773 ();
 sg13g2_decap_8 FILLER_41_780 ();
 sg13g2_decap_8 FILLER_41_787 ();
 sg13g2_decap_8 FILLER_41_794 ();
 sg13g2_decap_8 FILLER_41_801 ();
 sg13g2_decap_8 FILLER_41_808 ();
 sg13g2_decap_8 FILLER_41_815 ();
 sg13g2_decap_8 FILLER_41_822 ();
 sg13g2_decap_8 FILLER_41_829 ();
 sg13g2_decap_8 FILLER_41_836 ();
 sg13g2_decap_8 FILLER_41_843 ();
 sg13g2_decap_8 FILLER_41_850 ();
 sg13g2_decap_4 FILLER_41_857 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_4 FILLER_42_126 ();
 sg13g2_fill_2 FILLER_42_174 ();
 sg13g2_fill_1 FILLER_42_176 ();
 sg13g2_decap_4 FILLER_42_204 ();
 sg13g2_fill_2 FILLER_42_208 ();
 sg13g2_fill_1 FILLER_42_215 ();
 sg13g2_decap_4 FILLER_42_242 ();
 sg13g2_fill_2 FILLER_42_279 ();
 sg13g2_fill_2 FILLER_42_290 ();
 sg13g2_fill_1 FILLER_42_318 ();
 sg13g2_fill_2 FILLER_42_332 ();
 sg13g2_fill_2 FILLER_42_347 ();
 sg13g2_fill_1 FILLER_42_349 ();
 sg13g2_fill_1 FILLER_42_401 ();
 sg13g2_fill_1 FILLER_42_410 ();
 sg13g2_fill_2 FILLER_42_477 ();
 sg13g2_fill_1 FILLER_42_488 ();
 sg13g2_fill_1 FILLER_42_498 ();
 sg13g2_fill_2 FILLER_42_513 ();
 sg13g2_fill_1 FILLER_42_599 ();
 sg13g2_decap_8 FILLER_42_604 ();
 sg13g2_fill_2 FILLER_42_611 ();
 sg13g2_fill_1 FILLER_42_613 ();
 sg13g2_decap_4 FILLER_42_619 ();
 sg13g2_decap_8 FILLER_42_642 ();
 sg13g2_fill_2 FILLER_42_653 ();
 sg13g2_fill_1 FILLER_42_655 ();
 sg13g2_decap_8 FILLER_42_664 ();
 sg13g2_decap_8 FILLER_42_671 ();
 sg13g2_decap_8 FILLER_42_678 ();
 sg13g2_decap_8 FILLER_42_685 ();
 sg13g2_decap_8 FILLER_42_692 ();
 sg13g2_decap_8 FILLER_42_699 ();
 sg13g2_decap_8 FILLER_42_706 ();
 sg13g2_decap_8 FILLER_42_713 ();
 sg13g2_decap_8 FILLER_42_720 ();
 sg13g2_decap_8 FILLER_42_727 ();
 sg13g2_decap_8 FILLER_42_734 ();
 sg13g2_decap_8 FILLER_42_741 ();
 sg13g2_decap_8 FILLER_42_748 ();
 sg13g2_decap_8 FILLER_42_755 ();
 sg13g2_decap_8 FILLER_42_762 ();
 sg13g2_decap_8 FILLER_42_769 ();
 sg13g2_decap_8 FILLER_42_776 ();
 sg13g2_decap_8 FILLER_42_783 ();
 sg13g2_decap_8 FILLER_42_790 ();
 sg13g2_decap_8 FILLER_42_797 ();
 sg13g2_decap_8 FILLER_42_804 ();
 sg13g2_decap_8 FILLER_42_811 ();
 sg13g2_decap_8 FILLER_42_818 ();
 sg13g2_decap_8 FILLER_42_825 ();
 sg13g2_decap_8 FILLER_42_832 ();
 sg13g2_decap_8 FILLER_42_839 ();
 sg13g2_decap_8 FILLER_42_846 ();
 sg13g2_decap_8 FILLER_42_853 ();
 sg13g2_fill_2 FILLER_42_860 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_fill_2 FILLER_43_63 ();
 sg13g2_fill_1 FILLER_43_65 ();
 sg13g2_decap_8 FILLER_43_71 ();
 sg13g2_decap_8 FILLER_43_78 ();
 sg13g2_decap_8 FILLER_43_85 ();
 sg13g2_decap_8 FILLER_43_108 ();
 sg13g2_fill_1 FILLER_43_115 ();
 sg13g2_decap_8 FILLER_43_121 ();
 sg13g2_decap_4 FILLER_43_128 ();
 sg13g2_fill_2 FILLER_43_132 ();
 sg13g2_decap_8 FILLER_43_153 ();
 sg13g2_decap_4 FILLER_43_160 ();
 sg13g2_fill_2 FILLER_43_183 ();
 sg13g2_fill_1 FILLER_43_185 ();
 sg13g2_fill_1 FILLER_43_218 ();
 sg13g2_fill_1 FILLER_43_254 ();
 sg13g2_fill_2 FILLER_43_273 ();
 sg13g2_fill_2 FILLER_43_284 ();
 sg13g2_fill_1 FILLER_43_301 ();
 sg13g2_fill_1 FILLER_43_405 ();
 sg13g2_fill_1 FILLER_43_486 ();
 sg13g2_decap_8 FILLER_43_575 ();
 sg13g2_decap_8 FILLER_43_582 ();
 sg13g2_fill_1 FILLER_43_589 ();
 sg13g2_fill_1 FILLER_43_594 ();
 sg13g2_fill_2 FILLER_43_621 ();
 sg13g2_decap_8 FILLER_43_679 ();
 sg13g2_decap_8 FILLER_43_686 ();
 sg13g2_decap_8 FILLER_43_693 ();
 sg13g2_decap_8 FILLER_43_700 ();
 sg13g2_decap_8 FILLER_43_707 ();
 sg13g2_decap_8 FILLER_43_714 ();
 sg13g2_decap_8 FILLER_43_721 ();
 sg13g2_decap_8 FILLER_43_728 ();
 sg13g2_decap_8 FILLER_43_735 ();
 sg13g2_decap_8 FILLER_43_742 ();
 sg13g2_decap_8 FILLER_43_749 ();
 sg13g2_decap_8 FILLER_43_756 ();
 sg13g2_decap_8 FILLER_43_763 ();
 sg13g2_decap_8 FILLER_43_770 ();
 sg13g2_decap_8 FILLER_43_777 ();
 sg13g2_decap_8 FILLER_43_784 ();
 sg13g2_decap_8 FILLER_43_791 ();
 sg13g2_decap_8 FILLER_43_798 ();
 sg13g2_decap_8 FILLER_43_805 ();
 sg13g2_decap_8 FILLER_43_812 ();
 sg13g2_decap_8 FILLER_43_819 ();
 sg13g2_decap_8 FILLER_43_826 ();
 sg13g2_decap_8 FILLER_43_833 ();
 sg13g2_decap_8 FILLER_43_840 ();
 sg13g2_decap_8 FILLER_43_847 ();
 sg13g2_decap_8 FILLER_43_854 ();
 sg13g2_fill_1 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_4 FILLER_44_35 ();
 sg13g2_fill_1 FILLER_44_65 ();
 sg13g2_fill_1 FILLER_44_149 ();
 sg13g2_fill_1 FILLER_44_193 ();
 sg13g2_fill_2 FILLER_44_257 ();
 sg13g2_fill_1 FILLER_44_259 ();
 sg13g2_fill_2 FILLER_44_325 ();
 sg13g2_fill_2 FILLER_44_356 ();
 sg13g2_fill_1 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_416 ();
 sg13g2_fill_2 FILLER_44_447 ();
 sg13g2_fill_2 FILLER_44_458 ();
 sg13g2_decap_4 FILLER_44_503 ();
 sg13g2_fill_2 FILLER_44_507 ();
 sg13g2_decap_4 FILLER_44_513 ();
 sg13g2_fill_2 FILLER_44_517 ();
 sg13g2_decap_4 FILLER_44_545 ();
 sg13g2_fill_1 FILLER_44_549 ();
 sg13g2_fill_1 FILLER_44_576 ();
 sg13g2_fill_1 FILLER_44_644 ();
 sg13g2_decap_8 FILLER_44_698 ();
 sg13g2_decap_8 FILLER_44_705 ();
 sg13g2_decap_8 FILLER_44_712 ();
 sg13g2_decap_8 FILLER_44_719 ();
 sg13g2_decap_8 FILLER_44_726 ();
 sg13g2_decap_8 FILLER_44_733 ();
 sg13g2_decap_8 FILLER_44_740 ();
 sg13g2_decap_8 FILLER_44_747 ();
 sg13g2_decap_8 FILLER_44_754 ();
 sg13g2_decap_8 FILLER_44_761 ();
 sg13g2_decap_8 FILLER_44_768 ();
 sg13g2_decap_8 FILLER_44_775 ();
 sg13g2_decap_8 FILLER_44_782 ();
 sg13g2_decap_8 FILLER_44_789 ();
 sg13g2_decap_8 FILLER_44_796 ();
 sg13g2_decap_8 FILLER_44_803 ();
 sg13g2_decap_8 FILLER_44_810 ();
 sg13g2_decap_8 FILLER_44_817 ();
 sg13g2_decap_8 FILLER_44_824 ();
 sg13g2_decap_8 FILLER_44_831 ();
 sg13g2_decap_8 FILLER_44_838 ();
 sg13g2_decap_8 FILLER_44_845 ();
 sg13g2_decap_8 FILLER_44_852 ();
 sg13g2_fill_2 FILLER_44_859 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_4 FILLER_45_35 ();
 sg13g2_fill_1 FILLER_45_39 ();
 sg13g2_fill_1 FILLER_45_59 ();
 sg13g2_fill_1 FILLER_45_69 ();
 sg13g2_fill_2 FILLER_45_75 ();
 sg13g2_fill_1 FILLER_45_77 ();
 sg13g2_fill_1 FILLER_45_94 ();
 sg13g2_decap_4 FILLER_45_117 ();
 sg13g2_fill_2 FILLER_45_126 ();
 sg13g2_fill_1 FILLER_45_189 ();
 sg13g2_decap_4 FILLER_45_199 ();
 sg13g2_fill_2 FILLER_45_267 ();
 sg13g2_fill_1 FILLER_45_269 ();
 sg13g2_fill_1 FILLER_45_273 ();
 sg13g2_fill_1 FILLER_45_308 ();
 sg13g2_fill_2 FILLER_45_349 ();
 sg13g2_fill_1 FILLER_45_366 ();
 sg13g2_fill_1 FILLER_45_376 ();
 sg13g2_fill_1 FILLER_45_386 ();
 sg13g2_fill_1 FILLER_45_392 ();
 sg13g2_fill_2 FILLER_45_445 ();
 sg13g2_fill_1 FILLER_45_447 ();
 sg13g2_fill_1 FILLER_45_524 ();
 sg13g2_fill_1 FILLER_45_529 ();
 sg13g2_fill_2 FILLER_45_534 ();
 sg13g2_fill_1 FILLER_45_536 ();
 sg13g2_fill_1 FILLER_45_576 ();
 sg13g2_fill_2 FILLER_45_594 ();
 sg13g2_fill_1 FILLER_45_601 ();
 sg13g2_fill_1 FILLER_45_661 ();
 sg13g2_fill_2 FILLER_45_671 ();
 sg13g2_decap_8 FILLER_45_725 ();
 sg13g2_decap_8 FILLER_45_732 ();
 sg13g2_decap_8 FILLER_45_739 ();
 sg13g2_decap_8 FILLER_45_746 ();
 sg13g2_decap_8 FILLER_45_753 ();
 sg13g2_decap_8 FILLER_45_760 ();
 sg13g2_decap_8 FILLER_45_767 ();
 sg13g2_decap_8 FILLER_45_774 ();
 sg13g2_decap_8 FILLER_45_781 ();
 sg13g2_decap_8 FILLER_45_788 ();
 sg13g2_decap_8 FILLER_45_795 ();
 sg13g2_decap_8 FILLER_45_802 ();
 sg13g2_decap_8 FILLER_45_809 ();
 sg13g2_decap_8 FILLER_45_816 ();
 sg13g2_decap_8 FILLER_45_823 ();
 sg13g2_decap_8 FILLER_45_830 ();
 sg13g2_decap_8 FILLER_45_837 ();
 sg13g2_decap_8 FILLER_45_844 ();
 sg13g2_decap_8 FILLER_45_851 ();
 sg13g2_decap_4 FILLER_45_858 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_54 ();
 sg13g2_fill_1 FILLER_46_107 ();
 sg13g2_decap_8 FILLER_46_131 ();
 sg13g2_fill_2 FILLER_46_138 ();
 sg13g2_fill_1 FILLER_46_140 ();
 sg13g2_fill_1 FILLER_46_213 ();
 sg13g2_fill_1 FILLER_46_228 ();
 sg13g2_fill_2 FILLER_46_246 ();
 sg13g2_decap_8 FILLER_46_255 ();
 sg13g2_fill_2 FILLER_46_262 ();
 sg13g2_fill_1 FILLER_46_264 ();
 sg13g2_decap_4 FILLER_46_278 ();
 sg13g2_decap_4 FILLER_46_285 ();
 sg13g2_fill_2 FILLER_46_289 ();
 sg13g2_fill_2 FILLER_46_312 ();
 sg13g2_fill_1 FILLER_46_314 ();
 sg13g2_fill_1 FILLER_46_333 ();
 sg13g2_decap_8 FILLER_46_338 ();
 sg13g2_fill_2 FILLER_46_345 ();
 sg13g2_fill_1 FILLER_46_403 ();
 sg13g2_fill_2 FILLER_46_408 ();
 sg13g2_decap_4 FILLER_46_515 ();
 sg13g2_fill_2 FILLER_46_523 ();
 sg13g2_fill_1 FILLER_46_525 ();
 sg13g2_fill_1 FILLER_46_552 ();
 sg13g2_fill_1 FILLER_46_557 ();
 sg13g2_fill_1 FILLER_46_604 ();
 sg13g2_decap_8 FILLER_46_723 ();
 sg13g2_decap_8 FILLER_46_730 ();
 sg13g2_decap_8 FILLER_46_737 ();
 sg13g2_decap_8 FILLER_46_744 ();
 sg13g2_decap_8 FILLER_46_751 ();
 sg13g2_decap_8 FILLER_46_758 ();
 sg13g2_decap_8 FILLER_46_765 ();
 sg13g2_decap_8 FILLER_46_772 ();
 sg13g2_decap_8 FILLER_46_779 ();
 sg13g2_decap_8 FILLER_46_786 ();
 sg13g2_decap_8 FILLER_46_793 ();
 sg13g2_decap_8 FILLER_46_800 ();
 sg13g2_decap_8 FILLER_46_807 ();
 sg13g2_decap_8 FILLER_46_814 ();
 sg13g2_decap_8 FILLER_46_821 ();
 sg13g2_decap_8 FILLER_46_828 ();
 sg13g2_decap_8 FILLER_46_835 ();
 sg13g2_decap_8 FILLER_46_842 ();
 sg13g2_decap_8 FILLER_46_849 ();
 sg13g2_decap_4 FILLER_46_856 ();
 sg13g2_fill_2 FILLER_46_860 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_14 ();
 sg13g2_fill_1 FILLER_47_16 ();
 sg13g2_fill_2 FILLER_47_21 ();
 sg13g2_fill_2 FILLER_47_41 ();
 sg13g2_fill_2 FILLER_47_62 ();
 sg13g2_decap_4 FILLER_47_82 ();
 sg13g2_fill_1 FILLER_47_86 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_fill_1 FILLER_47_98 ();
 sg13g2_fill_2 FILLER_47_138 ();
 sg13g2_fill_1 FILLER_47_140 ();
 sg13g2_fill_2 FILLER_47_164 ();
 sg13g2_fill_2 FILLER_47_196 ();
 sg13g2_fill_2 FILLER_47_202 ();
 sg13g2_fill_1 FILLER_47_204 ();
 sg13g2_fill_1 FILLER_47_225 ();
 sg13g2_decap_4 FILLER_47_286 ();
 sg13g2_fill_1 FILLER_47_388 ();
 sg13g2_fill_2 FILLER_47_416 ();
 sg13g2_fill_2 FILLER_47_452 ();
 sg13g2_fill_1 FILLER_47_563 ();
 sg13g2_fill_1 FILLER_47_573 ();
 sg13g2_fill_1 FILLER_47_637 ();
 sg13g2_fill_1 FILLER_47_668 ();
 sg13g2_fill_2 FILLER_47_695 ();
 sg13g2_decap_8 FILLER_47_732 ();
 sg13g2_decap_8 FILLER_47_739 ();
 sg13g2_decap_8 FILLER_47_746 ();
 sg13g2_decap_8 FILLER_47_753 ();
 sg13g2_decap_8 FILLER_47_760 ();
 sg13g2_decap_8 FILLER_47_767 ();
 sg13g2_decap_8 FILLER_47_774 ();
 sg13g2_decap_8 FILLER_47_781 ();
 sg13g2_decap_8 FILLER_47_788 ();
 sg13g2_decap_8 FILLER_47_795 ();
 sg13g2_decap_8 FILLER_47_802 ();
 sg13g2_decap_8 FILLER_47_809 ();
 sg13g2_decap_8 FILLER_47_816 ();
 sg13g2_decap_8 FILLER_47_823 ();
 sg13g2_decap_8 FILLER_47_830 ();
 sg13g2_decap_8 FILLER_47_837 ();
 sg13g2_decap_8 FILLER_47_844 ();
 sg13g2_decap_8 FILLER_47_851 ();
 sg13g2_decap_4 FILLER_47_858 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_fill_2 FILLER_48_49 ();
 sg13g2_fill_1 FILLER_48_65 ();
 sg13g2_fill_1 FILLER_48_76 ();
 sg13g2_fill_1 FILLER_48_112 ();
 sg13g2_fill_1 FILLER_48_122 ();
 sg13g2_fill_2 FILLER_48_226 ();
 sg13g2_fill_2 FILLER_48_251 ();
 sg13g2_decap_8 FILLER_48_257 ();
 sg13g2_fill_1 FILLER_48_264 ();
 sg13g2_fill_1 FILLER_48_279 ();
 sg13g2_fill_1 FILLER_48_293 ();
 sg13g2_fill_1 FILLER_48_328 ();
 sg13g2_fill_2 FILLER_48_333 ();
 sg13g2_fill_2 FILLER_48_361 ();
 sg13g2_fill_2 FILLER_48_426 ();
 sg13g2_fill_2 FILLER_48_524 ();
 sg13g2_fill_2 FILLER_48_535 ();
 sg13g2_fill_1 FILLER_48_537 ();
 sg13g2_fill_2 FILLER_48_598 ();
 sg13g2_fill_2 FILLER_48_631 ();
 sg13g2_fill_2 FILLER_48_643 ();
 sg13g2_fill_2 FILLER_48_662 ();
 sg13g2_fill_1 FILLER_48_690 ();
 sg13g2_decap_8 FILLER_48_742 ();
 sg13g2_decap_8 FILLER_48_749 ();
 sg13g2_decap_8 FILLER_48_756 ();
 sg13g2_decap_8 FILLER_48_763 ();
 sg13g2_decap_8 FILLER_48_770 ();
 sg13g2_decap_8 FILLER_48_777 ();
 sg13g2_decap_8 FILLER_48_784 ();
 sg13g2_decap_8 FILLER_48_791 ();
 sg13g2_decap_8 FILLER_48_798 ();
 sg13g2_decap_8 FILLER_48_805 ();
 sg13g2_decap_8 FILLER_48_812 ();
 sg13g2_decap_8 FILLER_48_819 ();
 sg13g2_decap_8 FILLER_48_826 ();
 sg13g2_decap_8 FILLER_48_833 ();
 sg13g2_decap_8 FILLER_48_840 ();
 sg13g2_decap_8 FILLER_48_847 ();
 sg13g2_decap_8 FILLER_48_854 ();
 sg13g2_fill_1 FILLER_48_861 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_36 ();
 sg13g2_fill_2 FILLER_49_89 ();
 sg13g2_fill_1 FILLER_49_91 ();
 sg13g2_fill_1 FILLER_49_100 ();
 sg13g2_fill_2 FILLER_49_150 ();
 sg13g2_fill_1 FILLER_49_161 ();
 sg13g2_fill_2 FILLER_49_166 ();
 sg13g2_fill_2 FILLER_49_239 ();
 sg13g2_fill_1 FILLER_49_241 ();
 sg13g2_fill_2 FILLER_49_268 ();
 sg13g2_decap_8 FILLER_49_296 ();
 sg13g2_fill_1 FILLER_49_303 ();
 sg13g2_decap_8 FILLER_49_308 ();
 sg13g2_fill_2 FILLER_49_315 ();
 sg13g2_fill_1 FILLER_49_317 ();
 sg13g2_decap_4 FILLER_49_344 ();
 sg13g2_fill_2 FILLER_49_352 ();
 sg13g2_fill_2 FILLER_49_363 ();
 sg13g2_fill_1 FILLER_49_482 ();
 sg13g2_fill_2 FILLER_49_512 ();
 sg13g2_fill_2 FILLER_49_608 ();
 sg13g2_fill_2 FILLER_49_636 ();
 sg13g2_fill_1 FILLER_49_672 ();
 sg13g2_fill_2 FILLER_49_708 ();
 sg13g2_fill_2 FILLER_49_733 ();
 sg13g2_decap_8 FILLER_49_752 ();
 sg13g2_decap_8 FILLER_49_759 ();
 sg13g2_decap_8 FILLER_49_766 ();
 sg13g2_decap_8 FILLER_49_773 ();
 sg13g2_decap_8 FILLER_49_780 ();
 sg13g2_decap_8 FILLER_49_787 ();
 sg13g2_decap_8 FILLER_49_794 ();
 sg13g2_decap_8 FILLER_49_801 ();
 sg13g2_decap_8 FILLER_49_808 ();
 sg13g2_decap_8 FILLER_49_815 ();
 sg13g2_decap_8 FILLER_49_822 ();
 sg13g2_decap_8 FILLER_49_829 ();
 sg13g2_decap_8 FILLER_49_836 ();
 sg13g2_decap_8 FILLER_49_843 ();
 sg13g2_decap_8 FILLER_49_850 ();
 sg13g2_decap_4 FILLER_49_857 ();
 sg13g2_fill_1 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_7 ();
 sg13g2_fill_2 FILLER_50_51 ();
 sg13g2_fill_2 FILLER_50_79 ();
 sg13g2_fill_2 FILLER_50_107 ();
 sg13g2_fill_1 FILLER_50_120 ();
 sg13g2_fill_2 FILLER_50_126 ();
 sg13g2_fill_2 FILLER_50_134 ();
 sg13g2_fill_1 FILLER_50_140 ();
 sg13g2_fill_1 FILLER_50_145 ();
 sg13g2_fill_2 FILLER_50_172 ();
 sg13g2_fill_2 FILLER_50_186 ();
 sg13g2_fill_1 FILLER_50_223 ();
 sg13g2_fill_1 FILLER_50_239 ();
 sg13g2_fill_2 FILLER_50_249 ();
 sg13g2_fill_1 FILLER_50_251 ();
 sg13g2_fill_1 FILLER_50_324 ();
 sg13g2_decap_4 FILLER_50_329 ();
 sg13g2_fill_1 FILLER_50_333 ();
 sg13g2_fill_1 FILLER_50_360 ();
 sg13g2_decap_8 FILLER_50_374 ();
 sg13g2_fill_1 FILLER_50_425 ();
 sg13g2_fill_2 FILLER_50_436 ();
 sg13g2_fill_1 FILLER_50_438 ();
 sg13g2_fill_2 FILLER_50_448 ();
 sg13g2_fill_1 FILLER_50_450 ();
 sg13g2_fill_2 FILLER_50_475 ();
 sg13g2_fill_2 FILLER_50_486 ();
 sg13g2_fill_2 FILLER_50_519 ();
 sg13g2_fill_1 FILLER_50_521 ();
 sg13g2_fill_1 FILLER_50_536 ();
 sg13g2_fill_1 FILLER_50_597 ();
 sg13g2_fill_2 FILLER_50_628 ();
 sg13g2_fill_1 FILLER_50_635 ();
 sg13g2_fill_1 FILLER_50_645 ();
 sg13g2_decap_8 FILLER_50_747 ();
 sg13g2_decap_8 FILLER_50_754 ();
 sg13g2_decap_8 FILLER_50_761 ();
 sg13g2_decap_8 FILLER_50_768 ();
 sg13g2_decap_8 FILLER_50_775 ();
 sg13g2_decap_8 FILLER_50_782 ();
 sg13g2_decap_8 FILLER_50_789 ();
 sg13g2_decap_8 FILLER_50_796 ();
 sg13g2_decap_8 FILLER_50_803 ();
 sg13g2_decap_8 FILLER_50_810 ();
 sg13g2_decap_8 FILLER_50_817 ();
 sg13g2_decap_8 FILLER_50_824 ();
 sg13g2_decap_8 FILLER_50_831 ();
 sg13g2_decap_8 FILLER_50_838 ();
 sg13g2_decap_8 FILLER_50_845 ();
 sg13g2_decap_8 FILLER_50_852 ();
 sg13g2_fill_2 FILLER_50_859 ();
 sg13g2_fill_1 FILLER_50_861 ();
 sg13g2_fill_1 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_36 ();
 sg13g2_fill_2 FILLER_51_64 ();
 sg13g2_fill_2 FILLER_51_69 ();
 sg13g2_fill_2 FILLER_51_97 ();
 sg13g2_fill_1 FILLER_51_151 ();
 sg13g2_fill_1 FILLER_51_180 ();
 sg13g2_fill_2 FILLER_51_226 ();
 sg13g2_fill_1 FILLER_51_228 ();
 sg13g2_fill_2 FILLER_51_265 ();
 sg13g2_fill_1 FILLER_51_282 ();
 sg13g2_decap_8 FILLER_51_296 ();
 sg13g2_decap_4 FILLER_51_303 ();
 sg13g2_fill_2 FILLER_51_307 ();
 sg13g2_fill_2 FILLER_51_313 ();
 sg13g2_decap_4 FILLER_51_341 ();
 sg13g2_decap_4 FILLER_51_349 ();
 sg13g2_fill_1 FILLER_51_353 ();
 sg13g2_decap_8 FILLER_51_359 ();
 sg13g2_decap_8 FILLER_51_366 ();
 sg13g2_decap_4 FILLER_51_373 ();
 sg13g2_fill_2 FILLER_51_377 ();
 sg13g2_decap_4 FILLER_51_388 ();
 sg13g2_decap_4 FILLER_51_396 ();
 sg13g2_fill_1 FILLER_51_412 ();
 sg13g2_fill_2 FILLER_51_426 ();
 sg13g2_fill_1 FILLER_51_438 ();
 sg13g2_fill_2 FILLER_51_447 ();
 sg13g2_fill_1 FILLER_51_449 ();
 sg13g2_fill_2 FILLER_51_470 ();
 sg13g2_fill_1 FILLER_51_486 ();
 sg13g2_fill_1 FILLER_51_496 ();
 sg13g2_fill_2 FILLER_51_523 ();
 sg13g2_fill_1 FILLER_51_525 ();
 sg13g2_fill_2 FILLER_51_567 ();
 sg13g2_fill_2 FILLER_51_595 ();
 sg13g2_fill_2 FILLER_51_692 ();
 sg13g2_fill_2 FILLER_51_740 ();
 sg13g2_decap_8 FILLER_51_755 ();
 sg13g2_decap_8 FILLER_51_762 ();
 sg13g2_decap_8 FILLER_51_769 ();
 sg13g2_decap_8 FILLER_51_776 ();
 sg13g2_decap_8 FILLER_51_783 ();
 sg13g2_decap_8 FILLER_51_790 ();
 sg13g2_decap_8 FILLER_51_797 ();
 sg13g2_decap_8 FILLER_51_804 ();
 sg13g2_decap_8 FILLER_51_811 ();
 sg13g2_decap_8 FILLER_51_818 ();
 sg13g2_decap_8 FILLER_51_825 ();
 sg13g2_decap_8 FILLER_51_832 ();
 sg13g2_decap_8 FILLER_51_839 ();
 sg13g2_decap_8 FILLER_51_846 ();
 sg13g2_decap_8 FILLER_51_853 ();
 sg13g2_fill_2 FILLER_51_860 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_2 ();
 sg13g2_fill_2 FILLER_52_19 ();
 sg13g2_fill_1 FILLER_52_35 ();
 sg13g2_fill_1 FILLER_52_41 ();
 sg13g2_decap_4 FILLER_52_45 ();
 sg13g2_decap_4 FILLER_52_53 ();
 sg13g2_decap_8 FILLER_52_62 ();
 sg13g2_fill_2 FILLER_52_69 ();
 sg13g2_fill_1 FILLER_52_76 ();
 sg13g2_fill_2 FILLER_52_87 ();
 sg13g2_fill_1 FILLER_52_118 ();
 sg13g2_fill_1 FILLER_52_138 ();
 sg13g2_fill_1 FILLER_52_187 ();
 sg13g2_fill_2 FILLER_52_240 ();
 sg13g2_fill_1 FILLER_52_268 ();
 sg13g2_fill_2 FILLER_52_282 ();
 sg13g2_fill_1 FILLER_52_310 ();
 sg13g2_decap_8 FILLER_52_337 ();
 sg13g2_decap_8 FILLER_52_348 ();
 sg13g2_fill_2 FILLER_52_355 ();
 sg13g2_decap_8 FILLER_52_367 ();
 sg13g2_fill_2 FILLER_52_374 ();
 sg13g2_fill_1 FILLER_52_376 ();
 sg13g2_decap_8 FILLER_52_395 ();
 sg13g2_fill_2 FILLER_52_402 ();
 sg13g2_decap_4 FILLER_52_409 ();
 sg13g2_fill_1 FILLER_52_413 ();
 sg13g2_fill_2 FILLER_52_428 ();
 sg13g2_fill_1 FILLER_52_430 ();
 sg13g2_fill_2 FILLER_52_478 ();
 sg13g2_fill_1 FILLER_52_480 ();
 sg13g2_fill_2 FILLER_52_520 ();
 sg13g2_fill_1 FILLER_52_545 ();
 sg13g2_fill_2 FILLER_52_572 ();
 sg13g2_fill_1 FILLER_52_640 ();
 sg13g2_fill_1 FILLER_52_716 ();
 sg13g2_decap_8 FILLER_52_760 ();
 sg13g2_decap_8 FILLER_52_767 ();
 sg13g2_decap_8 FILLER_52_774 ();
 sg13g2_decap_8 FILLER_52_781 ();
 sg13g2_decap_8 FILLER_52_788 ();
 sg13g2_decap_8 FILLER_52_795 ();
 sg13g2_decap_8 FILLER_52_802 ();
 sg13g2_decap_8 FILLER_52_809 ();
 sg13g2_decap_8 FILLER_52_816 ();
 sg13g2_decap_8 FILLER_52_823 ();
 sg13g2_decap_8 FILLER_52_830 ();
 sg13g2_decap_8 FILLER_52_837 ();
 sg13g2_decap_8 FILLER_52_844 ();
 sg13g2_decap_8 FILLER_52_851 ();
 sg13g2_decap_4 FILLER_52_858 ();
 sg13g2_fill_2 FILLER_53_60 ();
 sg13g2_fill_1 FILLER_53_62 ();
 sg13g2_decap_8 FILLER_53_162 ();
 sg13g2_decap_4 FILLER_53_173 ();
 sg13g2_fill_1 FILLER_53_177 ();
 sg13g2_fill_2 FILLER_53_183 ();
 sg13g2_fill_1 FILLER_53_185 ();
 sg13g2_fill_2 FILLER_53_196 ();
 sg13g2_fill_2 FILLER_53_202 ();
 sg13g2_fill_1 FILLER_53_204 ();
 sg13g2_fill_2 FILLER_53_209 ();
 sg13g2_fill_1 FILLER_53_211 ();
 sg13g2_decap_4 FILLER_53_221 ();
 sg13g2_decap_4 FILLER_53_233 ();
 sg13g2_fill_1 FILLER_53_237 ();
 sg13g2_fill_1 FILLER_53_261 ();
 sg13g2_decap_8 FILLER_53_288 ();
 sg13g2_decap_8 FILLER_53_299 ();
 sg13g2_decap_4 FILLER_53_306 ();
 sg13g2_fill_1 FILLER_53_310 ();
 sg13g2_fill_2 FILLER_53_319 ();
 sg13g2_fill_1 FILLER_53_321 ();
 sg13g2_fill_2 FILLER_53_326 ();
 sg13g2_decap_4 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_425 ();
 sg13g2_fill_2 FILLER_53_436 ();
 sg13g2_fill_2 FILLER_53_456 ();
 sg13g2_fill_1 FILLER_53_458 ();
 sg13g2_fill_1 FILLER_53_545 ();
 sg13g2_fill_1 FILLER_53_560 ();
 sg13g2_fill_1 FILLER_53_571 ();
 sg13g2_fill_1 FILLER_53_611 ();
 sg13g2_fill_1 FILLER_53_644 ();
 sg13g2_fill_2 FILLER_53_663 ();
 sg13g2_fill_2 FILLER_53_679 ();
 sg13g2_decap_8 FILLER_53_757 ();
 sg13g2_decap_8 FILLER_53_764 ();
 sg13g2_decap_8 FILLER_53_771 ();
 sg13g2_decap_8 FILLER_53_778 ();
 sg13g2_decap_8 FILLER_53_785 ();
 sg13g2_decap_8 FILLER_53_792 ();
 sg13g2_decap_8 FILLER_53_799 ();
 sg13g2_decap_8 FILLER_53_806 ();
 sg13g2_decap_8 FILLER_53_813 ();
 sg13g2_decap_8 FILLER_53_820 ();
 sg13g2_decap_8 FILLER_53_827 ();
 sg13g2_decap_8 FILLER_53_834 ();
 sg13g2_decap_8 FILLER_53_841 ();
 sg13g2_decap_8 FILLER_53_848 ();
 sg13g2_decap_8 FILLER_53_855 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_7 ();
 sg13g2_fill_2 FILLER_54_48 ();
 sg13g2_fill_1 FILLER_54_50 ();
 sg13g2_fill_1 FILLER_54_83 ();
 sg13g2_fill_1 FILLER_54_140 ();
 sg13g2_fill_1 FILLER_54_150 ();
 sg13g2_fill_1 FILLER_54_165 ();
 sg13g2_decap_4 FILLER_54_179 ();
 sg13g2_fill_2 FILLER_54_183 ();
 sg13g2_fill_1 FILLER_54_223 ();
 sg13g2_decap_8 FILLER_54_262 ();
 sg13g2_decap_8 FILLER_54_269 ();
 sg13g2_decap_4 FILLER_54_276 ();
 sg13g2_fill_1 FILLER_54_280 ();
 sg13g2_fill_2 FILLER_54_285 ();
 sg13g2_decap_4 FILLER_54_313 ();
 sg13g2_fill_2 FILLER_54_317 ();
 sg13g2_decap_4 FILLER_54_323 ();
 sg13g2_fill_1 FILLER_54_327 ();
 sg13g2_fill_1 FILLER_54_345 ();
 sg13g2_fill_2 FILLER_54_364 ();
 sg13g2_decap_8 FILLER_54_377 ();
 sg13g2_decap_8 FILLER_54_384 ();
 sg13g2_fill_1 FILLER_54_417 ();
 sg13g2_fill_2 FILLER_54_423 ();
 sg13g2_fill_1 FILLER_54_461 ();
 sg13g2_fill_2 FILLER_54_524 ();
 sg13g2_fill_1 FILLER_54_526 ();
 sg13g2_fill_1 FILLER_54_604 ();
 sg13g2_fill_2 FILLER_54_640 ();
 sg13g2_fill_1 FILLER_54_647 ();
 sg13g2_fill_1 FILLER_54_723 ();
 sg13g2_decap_8 FILLER_54_757 ();
 sg13g2_decap_8 FILLER_54_764 ();
 sg13g2_decap_8 FILLER_54_771 ();
 sg13g2_decap_8 FILLER_54_778 ();
 sg13g2_decap_8 FILLER_54_785 ();
 sg13g2_decap_8 FILLER_54_792 ();
 sg13g2_decap_8 FILLER_54_799 ();
 sg13g2_decap_8 FILLER_54_806 ();
 sg13g2_decap_8 FILLER_54_813 ();
 sg13g2_decap_8 FILLER_54_820 ();
 sg13g2_decap_8 FILLER_54_827 ();
 sg13g2_decap_8 FILLER_54_834 ();
 sg13g2_decap_8 FILLER_54_841 ();
 sg13g2_decap_8 FILLER_54_848 ();
 sg13g2_decap_8 FILLER_54_855 ();
 sg13g2_fill_2 FILLER_55_53 ();
 sg13g2_fill_2 FILLER_55_64 ();
 sg13g2_fill_1 FILLER_55_66 ();
 sg13g2_fill_2 FILLER_55_98 ();
 sg13g2_fill_2 FILLER_55_119 ();
 sg13g2_fill_2 FILLER_55_217 ();
 sg13g2_fill_2 FILLER_55_242 ();
 sg13g2_fill_1 FILLER_55_269 ();
 sg13g2_fill_2 FILLER_55_296 ();
 sg13g2_decap_4 FILLER_55_302 ();
 sg13g2_fill_2 FILLER_55_306 ();
 sg13g2_fill_1 FILLER_55_334 ();
 sg13g2_fill_2 FILLER_55_357 ();
 sg13g2_decap_4 FILLER_55_398 ();
 sg13g2_decap_8 FILLER_55_406 ();
 sg13g2_decap_8 FILLER_55_413 ();
 sg13g2_fill_2 FILLER_55_420 ();
 sg13g2_fill_1 FILLER_55_430 ();
 sg13g2_fill_2 FILLER_55_462 ();
 sg13g2_fill_1 FILLER_55_464 ();
 sg13g2_fill_1 FILLER_55_474 ();
 sg13g2_decap_4 FILLER_55_501 ();
 sg13g2_fill_1 FILLER_55_505 ();
 sg13g2_decap_8 FILLER_55_510 ();
 sg13g2_fill_2 FILLER_55_530 ();
 sg13g2_fill_2 FILLER_55_555 ();
 sg13g2_fill_1 FILLER_55_561 ();
 sg13g2_fill_2 FILLER_55_575 ();
 sg13g2_fill_2 FILLER_55_586 ();
 sg13g2_fill_1 FILLER_55_593 ();
 sg13g2_fill_1 FILLER_55_607 ();
 sg13g2_fill_2 FILLER_55_620 ();
 sg13g2_fill_2 FILLER_55_666 ();
 sg13g2_fill_1 FILLER_55_691 ();
 sg13g2_fill_1 FILLER_55_706 ();
 sg13g2_decap_8 FILLER_55_763 ();
 sg13g2_decap_8 FILLER_55_770 ();
 sg13g2_decap_8 FILLER_55_777 ();
 sg13g2_decap_8 FILLER_55_784 ();
 sg13g2_decap_8 FILLER_55_791 ();
 sg13g2_decap_8 FILLER_55_798 ();
 sg13g2_decap_8 FILLER_55_805 ();
 sg13g2_decap_8 FILLER_55_812 ();
 sg13g2_decap_8 FILLER_55_819 ();
 sg13g2_decap_8 FILLER_55_826 ();
 sg13g2_decap_8 FILLER_55_833 ();
 sg13g2_decap_8 FILLER_55_840 ();
 sg13g2_decap_8 FILLER_55_847 ();
 sg13g2_decap_8 FILLER_55_854 ();
 sg13g2_fill_1 FILLER_55_861 ();
 sg13g2_decap_4 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_4 ();
 sg13g2_fill_1 FILLER_56_111 ();
 sg13g2_fill_2 FILLER_56_153 ();
 sg13g2_fill_1 FILLER_56_155 ();
 sg13g2_fill_2 FILLER_56_210 ();
 sg13g2_fill_1 FILLER_56_225 ();
 sg13g2_decap_4 FILLER_56_241 ();
 sg13g2_fill_2 FILLER_56_259 ();
 sg13g2_fill_1 FILLER_56_264 ();
 sg13g2_decap_8 FILLER_56_275 ();
 sg13g2_decap_4 FILLER_56_282 ();
 sg13g2_fill_2 FILLER_56_286 ();
 sg13g2_decap_8 FILLER_56_314 ();
 sg13g2_decap_4 FILLER_56_321 ();
 sg13g2_fill_2 FILLER_56_378 ();
 sg13g2_fill_1 FILLER_56_385 ();
 sg13g2_fill_2 FILLER_56_438 ();
 sg13g2_fill_2 FILLER_56_444 ();
 sg13g2_fill_1 FILLER_56_446 ();
 sg13g2_decap_4 FILLER_56_491 ();
 sg13g2_fill_1 FILLER_56_521 ();
 sg13g2_fill_1 FILLER_56_527 ();
 sg13g2_fill_1 FILLER_56_533 ();
 sg13g2_fill_1 FILLER_56_538 ();
 sg13g2_fill_1 FILLER_56_570 ();
 sg13g2_fill_2 FILLER_56_585 ();
 sg13g2_fill_2 FILLER_56_650 ();
 sg13g2_fill_1 FILLER_56_689 ();
 sg13g2_decap_8 FILLER_56_760 ();
 sg13g2_decap_8 FILLER_56_767 ();
 sg13g2_decap_8 FILLER_56_774 ();
 sg13g2_decap_8 FILLER_56_781 ();
 sg13g2_decap_8 FILLER_56_788 ();
 sg13g2_decap_8 FILLER_56_795 ();
 sg13g2_decap_8 FILLER_56_802 ();
 sg13g2_decap_8 FILLER_56_809 ();
 sg13g2_decap_8 FILLER_56_816 ();
 sg13g2_decap_8 FILLER_56_823 ();
 sg13g2_decap_8 FILLER_56_830 ();
 sg13g2_decap_8 FILLER_56_837 ();
 sg13g2_decap_8 FILLER_56_844 ();
 sg13g2_decap_8 FILLER_56_851 ();
 sg13g2_decap_4 FILLER_56_858 ();
 sg13g2_fill_1 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_47 ();
 sg13g2_fill_1 FILLER_57_49 ();
 sg13g2_fill_1 FILLER_57_54 ();
 sg13g2_fill_2 FILLER_57_64 ();
 sg13g2_fill_1 FILLER_57_66 ();
 sg13g2_decap_8 FILLER_57_72 ();
 sg13g2_fill_2 FILLER_57_84 ();
 sg13g2_fill_1 FILLER_57_86 ();
 sg13g2_fill_2 FILLER_57_91 ();
 sg13g2_fill_1 FILLER_57_93 ();
 sg13g2_fill_1 FILLER_57_99 ();
 sg13g2_decap_4 FILLER_57_105 ();
 sg13g2_fill_2 FILLER_57_114 ();
 sg13g2_fill_1 FILLER_57_116 ();
 sg13g2_decap_4 FILLER_57_143 ();
 sg13g2_fill_1 FILLER_57_147 ();
 sg13g2_fill_2 FILLER_57_170 ();
 sg13g2_fill_1 FILLER_57_172 ();
 sg13g2_fill_1 FILLER_57_191 ();
 sg13g2_fill_2 FILLER_57_196 ();
 sg13g2_fill_1 FILLER_57_198 ();
 sg13g2_fill_2 FILLER_57_233 ();
 sg13g2_fill_2 FILLER_57_261 ();
 sg13g2_fill_2 FILLER_57_270 ();
 sg13g2_fill_1 FILLER_57_272 ();
 sg13g2_decap_8 FILLER_57_303 ();
 sg13g2_fill_1 FILLER_57_310 ();
 sg13g2_fill_2 FILLER_57_361 ();
 sg13g2_fill_2 FILLER_57_376 ();
 sg13g2_fill_1 FILLER_57_378 ();
 sg13g2_decap_8 FILLER_57_429 ();
 sg13g2_decap_4 FILLER_57_436 ();
 sg13g2_fill_1 FILLER_57_488 ();
 sg13g2_decap_4 FILLER_57_515 ();
 sg13g2_fill_1 FILLER_57_519 ();
 sg13g2_decap_4 FILLER_57_537 ();
 sg13g2_fill_2 FILLER_57_541 ();
 sg13g2_decap_8 FILLER_57_576 ();
 sg13g2_fill_2 FILLER_57_609 ();
 sg13g2_fill_1 FILLER_57_611 ();
 sg13g2_fill_2 FILLER_57_642 ();
 sg13g2_fill_1 FILLER_57_676 ();
 sg13g2_fill_1 FILLER_57_712 ();
 sg13g2_decap_8 FILLER_57_765 ();
 sg13g2_decap_8 FILLER_57_772 ();
 sg13g2_decap_8 FILLER_57_779 ();
 sg13g2_decap_8 FILLER_57_786 ();
 sg13g2_decap_8 FILLER_57_793 ();
 sg13g2_decap_8 FILLER_57_800 ();
 sg13g2_decap_8 FILLER_57_807 ();
 sg13g2_decap_8 FILLER_57_814 ();
 sg13g2_decap_8 FILLER_57_821 ();
 sg13g2_decap_8 FILLER_57_828 ();
 sg13g2_decap_8 FILLER_57_835 ();
 sg13g2_decap_8 FILLER_57_842 ();
 sg13g2_decap_8 FILLER_57_849 ();
 sg13g2_decap_4 FILLER_57_856 ();
 sg13g2_fill_2 FILLER_57_860 ();
 sg13g2_fill_1 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_27 ();
 sg13g2_fill_1 FILLER_58_33 ();
 sg13g2_fill_1 FILLER_58_70 ();
 sg13g2_fill_2 FILLER_58_102 ();
 sg13g2_fill_1 FILLER_58_109 ();
 sg13g2_decap_4 FILLER_58_136 ();
 sg13g2_fill_1 FILLER_58_140 ();
 sg13g2_fill_1 FILLER_58_207 ();
 sg13g2_decap_4 FILLER_58_217 ();
 sg13g2_decap_8 FILLER_58_231 ();
 sg13g2_decap_4 FILLER_58_238 ();
 sg13g2_fill_1 FILLER_58_242 ();
 sg13g2_decap_4 FILLER_58_278 ();
 sg13g2_fill_2 FILLER_58_282 ();
 sg13g2_decap_8 FILLER_58_288 ();
 sg13g2_decap_4 FILLER_58_295 ();
 sg13g2_decap_4 FILLER_58_304 ();
 sg13g2_fill_1 FILLER_58_308 ();
 sg13g2_fill_2 FILLER_58_319 ();
 sg13g2_fill_1 FILLER_58_321 ();
 sg13g2_decap_4 FILLER_58_326 ();
 sg13g2_fill_2 FILLER_58_330 ();
 sg13g2_decap_4 FILLER_58_345 ();
 sg13g2_fill_2 FILLER_58_349 ();
 sg13g2_fill_1 FILLER_58_359 ();
 sg13g2_fill_1 FILLER_58_373 ();
 sg13g2_fill_2 FILLER_58_406 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_58_435 ();
 sg13g2_decap_8 FILLER_58_442 ();
 sg13g2_fill_2 FILLER_58_449 ();
 sg13g2_fill_2 FILLER_58_486 ();
 sg13g2_fill_1 FILLER_58_488 ();
 sg13g2_fill_2 FILLER_58_497 ();
 sg13g2_fill_1 FILLER_58_499 ();
 sg13g2_decap_8 FILLER_58_504 ();
 sg13g2_decap_4 FILLER_58_511 ();
 sg13g2_fill_2 FILLER_58_546 ();
 sg13g2_fill_1 FILLER_58_548 ();
 sg13g2_fill_2 FILLER_58_558 ();
 sg13g2_decap_8 FILLER_58_572 ();
 sg13g2_fill_2 FILLER_58_579 ();
 sg13g2_fill_1 FILLER_58_581 ();
 sg13g2_fill_1 FILLER_58_592 ();
 sg13g2_fill_1 FILLER_58_664 ();
 sg13g2_decap_8 FILLER_58_771 ();
 sg13g2_decap_8 FILLER_58_778 ();
 sg13g2_decap_8 FILLER_58_785 ();
 sg13g2_decap_8 FILLER_58_792 ();
 sg13g2_decap_8 FILLER_58_799 ();
 sg13g2_decap_8 FILLER_58_806 ();
 sg13g2_decap_8 FILLER_58_813 ();
 sg13g2_decap_8 FILLER_58_820 ();
 sg13g2_decap_8 FILLER_58_827 ();
 sg13g2_decap_8 FILLER_58_834 ();
 sg13g2_decap_8 FILLER_58_841 ();
 sg13g2_decap_8 FILLER_58_848 ();
 sg13g2_decap_8 FILLER_58_855 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_2 ();
 sg13g2_fill_2 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_46 ();
 sg13g2_decap_4 FILLER_59_53 ();
 sg13g2_fill_2 FILLER_59_57 ();
 sg13g2_fill_2 FILLER_59_71 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_fill_2 FILLER_59_98 ();
 sg13g2_fill_2 FILLER_59_110 ();
 sg13g2_fill_1 FILLER_59_112 ();
 sg13g2_decap_4 FILLER_59_118 ();
 sg13g2_decap_8 FILLER_59_131 ();
 sg13g2_fill_2 FILLER_59_138 ();
 sg13g2_fill_2 FILLER_59_204 ();
 sg13g2_decap_8 FILLER_59_263 ();
 sg13g2_fill_2 FILLER_59_270 ();
 sg13g2_fill_2 FILLER_59_292 ();
 sg13g2_decap_4 FILLER_59_323 ();
 sg13g2_fill_2 FILLER_59_327 ();
 sg13g2_fill_1 FILLER_59_359 ();
 sg13g2_decap_8 FILLER_59_364 ();
 sg13g2_decap_4 FILLER_59_371 ();
 sg13g2_fill_1 FILLER_59_375 ();
 sg13g2_decap_8 FILLER_59_396 ();
 sg13g2_decap_8 FILLER_59_403 ();
 sg13g2_fill_2 FILLER_59_418 ();
 sg13g2_fill_2 FILLER_59_424 ();
 sg13g2_fill_1 FILLER_59_426 ();
 sg13g2_fill_2 FILLER_59_440 ();
 sg13g2_fill_1 FILLER_59_451 ();
 sg13g2_fill_2 FILLER_59_468 ();
 sg13g2_fill_2 FILLER_59_519 ();
 sg13g2_fill_1 FILLER_59_521 ();
 sg13g2_fill_1 FILLER_59_540 ();
 sg13g2_fill_1 FILLER_59_577 ();
 sg13g2_fill_1 FILLER_59_604 ();
 sg13g2_fill_1 FILLER_59_662 ();
 sg13g2_fill_2 FILLER_59_700 ();
 sg13g2_decap_8 FILLER_59_760 ();
 sg13g2_decap_8 FILLER_59_767 ();
 sg13g2_decap_8 FILLER_59_774 ();
 sg13g2_decap_8 FILLER_59_781 ();
 sg13g2_decap_8 FILLER_59_788 ();
 sg13g2_decap_8 FILLER_59_795 ();
 sg13g2_decap_8 FILLER_59_802 ();
 sg13g2_decap_8 FILLER_59_809 ();
 sg13g2_decap_8 FILLER_59_816 ();
 sg13g2_decap_8 FILLER_59_823 ();
 sg13g2_decap_8 FILLER_59_830 ();
 sg13g2_decap_8 FILLER_59_837 ();
 sg13g2_decap_8 FILLER_59_844 ();
 sg13g2_decap_8 FILLER_59_851 ();
 sg13g2_decap_4 FILLER_59_858 ();
 sg13g2_fill_2 FILLER_60_26 ();
 sg13g2_fill_1 FILLER_60_28 ();
 sg13g2_fill_1 FILLER_60_38 ();
 sg13g2_fill_2 FILLER_60_53 ();
 sg13g2_fill_2 FILLER_60_125 ();
 sg13g2_fill_1 FILLER_60_133 ();
 sg13g2_fill_1 FILLER_60_200 ();
 sg13g2_fill_1 FILLER_60_206 ();
 sg13g2_decap_8 FILLER_60_236 ();
 sg13g2_fill_2 FILLER_60_243 ();
 sg13g2_fill_1 FILLER_60_275 ();
 sg13g2_decap_8 FILLER_60_292 ();
 sg13g2_fill_1 FILLER_60_299 ();
 sg13g2_decap_8 FILLER_60_327 ();
 sg13g2_decap_4 FILLER_60_334 ();
 sg13g2_fill_1 FILLER_60_338 ();
 sg13g2_decap_4 FILLER_60_343 ();
 sg13g2_decap_8 FILLER_60_365 ();
 sg13g2_fill_2 FILLER_60_372 ();
 sg13g2_decap_8 FILLER_60_388 ();
 sg13g2_fill_2 FILLER_60_417 ();
 sg13g2_fill_2 FILLER_60_455 ();
 sg13g2_fill_2 FILLER_60_461 ();
 sg13g2_fill_2 FILLER_60_484 ();
 sg13g2_fill_2 FILLER_60_499 ();
 sg13g2_fill_1 FILLER_60_501 ();
 sg13g2_decap_4 FILLER_60_546 ();
 sg13g2_fill_1 FILLER_60_550 ();
 sg13g2_decap_8 FILLER_60_555 ();
 sg13g2_decap_4 FILLER_60_572 ();
 sg13g2_fill_2 FILLER_60_576 ();
 sg13g2_fill_2 FILLER_60_583 ();
 sg13g2_fill_2 FILLER_60_599 ();
 sg13g2_fill_1 FILLER_60_601 ();
 sg13g2_fill_1 FILLER_60_660 ();
 sg13g2_fill_1 FILLER_60_713 ();
 sg13g2_decap_8 FILLER_60_770 ();
 sg13g2_decap_8 FILLER_60_777 ();
 sg13g2_decap_8 FILLER_60_784 ();
 sg13g2_decap_8 FILLER_60_791 ();
 sg13g2_decap_8 FILLER_60_798 ();
 sg13g2_decap_8 FILLER_60_805 ();
 sg13g2_decap_8 FILLER_60_812 ();
 sg13g2_decap_8 FILLER_60_819 ();
 sg13g2_decap_8 FILLER_60_826 ();
 sg13g2_decap_8 FILLER_60_833 ();
 sg13g2_decap_8 FILLER_60_840 ();
 sg13g2_decap_8 FILLER_60_847 ();
 sg13g2_decap_8 FILLER_60_854 ();
 sg13g2_fill_1 FILLER_60_861 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_2 ();
 sg13g2_fill_2 FILLER_61_26 ();
 sg13g2_fill_1 FILLER_61_28 ();
 sg13g2_fill_1 FILLER_61_55 ();
 sg13g2_decap_4 FILLER_61_87 ();
 sg13g2_fill_1 FILLER_61_91 ();
 sg13g2_fill_1 FILLER_61_122 ();
 sg13g2_fill_1 FILLER_61_137 ();
 sg13g2_fill_1 FILLER_61_172 ();
 sg13g2_fill_1 FILLER_61_182 ();
 sg13g2_fill_1 FILLER_61_188 ();
 sg13g2_fill_1 FILLER_61_214 ();
 sg13g2_decap_8 FILLER_61_241 ();
 sg13g2_decap_8 FILLER_61_248 ();
 sg13g2_decap_4 FILLER_61_255 ();
 sg13g2_fill_1 FILLER_61_259 ();
 sg13g2_decap_8 FILLER_61_264 ();
 sg13g2_decap_8 FILLER_61_271 ();
 sg13g2_decap_8 FILLER_61_288 ();
 sg13g2_fill_2 FILLER_61_295 ();
 sg13g2_fill_1 FILLER_61_297 ();
 sg13g2_fill_2 FILLER_61_324 ();
 sg13g2_fill_1 FILLER_61_326 ();
 sg13g2_fill_1 FILLER_61_384 ();
 sg13g2_fill_1 FILLER_61_425 ();
 sg13g2_fill_2 FILLER_61_438 ();
 sg13g2_fill_1 FILLER_61_440 ();
 sg13g2_fill_2 FILLER_61_465 ();
 sg13g2_fill_1 FILLER_61_467 ();
 sg13g2_decap_8 FILLER_61_506 ();
 sg13g2_decap_8 FILLER_61_513 ();
 sg13g2_fill_1 FILLER_61_520 ();
 sg13g2_fill_1 FILLER_61_529 ();
 sg13g2_fill_2 FILLER_61_534 ();
 sg13g2_decap_8 FILLER_61_554 ();
 sg13g2_fill_1 FILLER_61_561 ();
 sg13g2_decap_8 FILLER_61_578 ();
 sg13g2_decap_8 FILLER_61_585 ();
 sg13g2_fill_1 FILLER_61_592 ();
 sg13g2_decap_4 FILLER_61_597 ();
 sg13g2_fill_2 FILLER_61_620 ();
 sg13g2_fill_2 FILLER_61_677 ();
 sg13g2_fill_2 FILLER_61_697 ();
 sg13g2_fill_2 FILLER_61_717 ();
 sg13g2_fill_1 FILLER_61_719 ();
 sg13g2_fill_2 FILLER_61_740 ();
 sg13g2_decap_8 FILLER_61_768 ();
 sg13g2_decap_8 FILLER_61_775 ();
 sg13g2_decap_8 FILLER_61_782 ();
 sg13g2_decap_8 FILLER_61_789 ();
 sg13g2_decap_8 FILLER_61_796 ();
 sg13g2_decap_8 FILLER_61_803 ();
 sg13g2_decap_8 FILLER_61_810 ();
 sg13g2_decap_8 FILLER_61_817 ();
 sg13g2_decap_8 FILLER_61_824 ();
 sg13g2_decap_8 FILLER_61_831 ();
 sg13g2_decap_8 FILLER_61_838 ();
 sg13g2_decap_8 FILLER_61_845 ();
 sg13g2_decap_8 FILLER_61_852 ();
 sg13g2_fill_2 FILLER_61_859 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_decap_4 FILLER_62_45 ();
 sg13g2_fill_2 FILLER_62_77 ();
 sg13g2_fill_1 FILLER_62_79 ();
 sg13g2_fill_1 FILLER_62_106 ();
 sg13g2_fill_2 FILLER_62_123 ();
 sg13g2_fill_2 FILLER_62_176 ();
 sg13g2_fill_1 FILLER_62_205 ();
 sg13g2_decap_4 FILLER_62_215 ();
 sg13g2_fill_2 FILLER_62_219 ();
 sg13g2_fill_2 FILLER_62_273 ();
 sg13g2_fill_2 FILLER_62_306 ();
 sg13g2_fill_1 FILLER_62_308 ();
 sg13g2_decap_8 FILLER_62_329 ();
 sg13g2_fill_1 FILLER_62_351 ();
 sg13g2_decap_4 FILLER_62_365 ();
 sg13g2_fill_1 FILLER_62_373 ();
 sg13g2_decap_8 FILLER_62_421 ();
 sg13g2_decap_4 FILLER_62_428 ();
 sg13g2_fill_1 FILLER_62_432 ();
 sg13g2_decap_4 FILLER_62_459 ();
 sg13g2_fill_2 FILLER_62_530 ();
 sg13g2_fill_1 FILLER_62_532 ();
 sg13g2_fill_2 FILLER_62_564 ();
 sg13g2_fill_2 FILLER_62_729 ();
 sg13g2_fill_1 FILLER_62_766 ();
 sg13g2_decap_8 FILLER_62_771 ();
 sg13g2_decap_8 FILLER_62_808 ();
 sg13g2_decap_8 FILLER_62_815 ();
 sg13g2_decap_8 FILLER_62_822 ();
 sg13g2_decap_8 FILLER_62_829 ();
 sg13g2_decap_8 FILLER_62_836 ();
 sg13g2_decap_8 FILLER_62_843 ();
 sg13g2_decap_8 FILLER_62_850 ();
 sg13g2_decap_4 FILLER_62_857 ();
 sg13g2_fill_1 FILLER_62_861 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_7 ();
 sg13g2_fill_2 FILLER_63_35 ();
 sg13g2_fill_1 FILLER_63_37 ();
 sg13g2_fill_2 FILLER_63_74 ();
 sg13g2_fill_1 FILLER_63_76 ();
 sg13g2_fill_1 FILLER_63_95 ();
 sg13g2_decap_4 FILLER_63_205 ();
 sg13g2_fill_2 FILLER_63_209 ();
 sg13g2_decap_8 FILLER_63_215 ();
 sg13g2_decap_4 FILLER_63_222 ();
 sg13g2_decap_4 FILLER_63_230 ();
 sg13g2_fill_2 FILLER_63_234 ();
 sg13g2_decap_8 FILLER_63_240 ();
 sg13g2_fill_2 FILLER_63_273 ();
 sg13g2_decap_4 FILLER_63_297 ();
 sg13g2_fill_2 FILLER_63_306 ();
 sg13g2_decap_4 FILLER_63_319 ();
 sg13g2_decap_8 FILLER_63_369 ();
 sg13g2_decap_4 FILLER_63_420 ();
 sg13g2_fill_2 FILLER_63_442 ();
 sg13g2_decap_4 FILLER_63_472 ();
 sg13g2_fill_2 FILLER_63_502 ();
 sg13g2_fill_1 FILLER_63_509 ();
 sg13g2_fill_1 FILLER_63_527 ();
 sg13g2_fill_2 FILLER_63_564 ();
 sg13g2_fill_1 FILLER_63_566 ();
 sg13g2_fill_2 FILLER_63_580 ();
 sg13g2_fill_2 FILLER_63_587 ();
 sg13g2_decap_4 FILLER_63_623 ();
 sg13g2_fill_1 FILLER_63_631 ();
 sg13g2_fill_2 FILLER_63_669 ();
 sg13g2_fill_1 FILLER_63_671 ();
 sg13g2_fill_2 FILLER_63_676 ();
 sg13g2_fill_1 FILLER_63_678 ();
 sg13g2_fill_1 FILLER_63_684 ();
 sg13g2_fill_1 FILLER_63_724 ();
 sg13g2_fill_2 FILLER_63_747 ();
 sg13g2_decap_8 FILLER_63_805 ();
 sg13g2_decap_8 FILLER_63_812 ();
 sg13g2_decap_8 FILLER_63_819 ();
 sg13g2_decap_8 FILLER_63_826 ();
 sg13g2_decap_8 FILLER_63_833 ();
 sg13g2_decap_8 FILLER_63_840 ();
 sg13g2_decap_8 FILLER_63_847 ();
 sg13g2_decap_8 FILLER_63_854 ();
 sg13g2_fill_1 FILLER_63_861 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_7 ();
 sg13g2_fill_1 FILLER_64_44 ();
 sg13g2_fill_1 FILLER_64_50 ();
 sg13g2_decap_8 FILLER_64_69 ();
 sg13g2_decap_4 FILLER_64_76 ();
 sg13g2_fill_1 FILLER_64_80 ();
 sg13g2_fill_1 FILLER_64_113 ();
 sg13g2_fill_1 FILLER_64_128 ();
 sg13g2_fill_2 FILLER_64_133 ();
 sg13g2_fill_2 FILLER_64_143 ();
 sg13g2_fill_1 FILLER_64_145 ();
 sg13g2_fill_1 FILLER_64_172 ();
 sg13g2_fill_2 FILLER_64_188 ();
 sg13g2_fill_2 FILLER_64_194 ();
 sg13g2_fill_1 FILLER_64_196 ();
 sg13g2_fill_2 FILLER_64_226 ();
 sg13g2_fill_1 FILLER_64_228 ();
 sg13g2_fill_2 FILLER_64_255 ();
 sg13g2_fill_2 FILLER_64_302 ();
 sg13g2_decap_8 FILLER_64_324 ();
 sg13g2_decap_4 FILLER_64_331 ();
 sg13g2_fill_1 FILLER_64_349 ();
 sg13g2_fill_1 FILLER_64_354 ();
 sg13g2_fill_2 FILLER_64_363 ();
 sg13g2_fill_2 FILLER_64_370 ();
 sg13g2_fill_1 FILLER_64_405 ();
 sg13g2_fill_1 FILLER_64_415 ();
 sg13g2_fill_2 FILLER_64_425 ();
 sg13g2_fill_1 FILLER_64_448 ();
 sg13g2_decap_4 FILLER_64_491 ();
 sg13g2_fill_1 FILLER_64_548 ();
 sg13g2_fill_1 FILLER_64_587 ();
 sg13g2_fill_1 FILLER_64_662 ();
 sg13g2_fill_2 FILLER_64_710 ();
 sg13g2_fill_1 FILLER_64_712 ();
 sg13g2_decap_4 FILLER_64_739 ();
 sg13g2_fill_2 FILLER_64_743 ();
 sg13g2_fill_1 FILLER_64_785 ();
 sg13g2_decap_8 FILLER_64_830 ();
 sg13g2_decap_8 FILLER_64_837 ();
 sg13g2_decap_8 FILLER_64_844 ();
 sg13g2_decap_8 FILLER_64_851 ();
 sg13g2_decap_4 FILLER_64_858 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_36 ();
 sg13g2_fill_2 FILLER_65_122 ();
 sg13g2_fill_1 FILLER_65_135 ();
 sg13g2_fill_1 FILLER_65_141 ();
 sg13g2_decap_8 FILLER_65_150 ();
 sg13g2_decap_4 FILLER_65_161 ();
 sg13g2_fill_2 FILLER_65_165 ();
 sg13g2_decap_4 FILLER_65_172 ();
 sg13g2_fill_1 FILLER_65_176 ();
 sg13g2_fill_1 FILLER_65_183 ();
 sg13g2_fill_2 FILLER_65_190 ();
 sg13g2_fill_2 FILLER_65_207 ();
 sg13g2_fill_2 FILLER_65_224 ();
 sg13g2_fill_1 FILLER_65_226 ();
 sg13g2_decap_8 FILLER_65_248 ();
 sg13g2_fill_2 FILLER_65_255 ();
 sg13g2_fill_1 FILLER_65_257 ();
 sg13g2_decap_8 FILLER_65_262 ();
 sg13g2_decap_4 FILLER_65_269 ();
 sg13g2_fill_1 FILLER_65_273 ();
 sg13g2_fill_2 FILLER_65_309 ();
 sg13g2_decap_8 FILLER_65_319 ();
 sg13g2_fill_2 FILLER_65_326 ();
 sg13g2_fill_2 FILLER_65_456 ();
 sg13g2_decap_8 FILLER_65_488 ();
 sg13g2_fill_1 FILLER_65_528 ();
 sg13g2_fill_2 FILLER_65_547 ();
 sg13g2_decap_8 FILLER_65_574 ();
 sg13g2_fill_2 FILLER_65_581 ();
 sg13g2_fill_1 FILLER_65_583 ();
 sg13g2_fill_2 FILLER_65_615 ();
 sg13g2_fill_1 FILLER_65_617 ();
 sg13g2_fill_2 FILLER_65_665 ();
 sg13g2_fill_1 FILLER_65_667 ();
 sg13g2_fill_1 FILLER_65_723 ();
 sg13g2_fill_1 FILLER_65_729 ();
 sg13g2_fill_1 FILLER_65_761 ();
 sg13g2_decap_8 FILLER_65_826 ();
 sg13g2_decap_8 FILLER_65_833 ();
 sg13g2_decap_8 FILLER_65_840 ();
 sg13g2_decap_8 FILLER_65_847 ();
 sg13g2_decap_8 FILLER_65_854 ();
 sg13g2_fill_1 FILLER_65_861 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_4 FILLER_66_7 ();
 sg13g2_fill_2 FILLER_66_11 ();
 sg13g2_fill_2 FILLER_66_17 ();
 sg13g2_fill_1 FILLER_66_28 ();
 sg13g2_decap_4 FILLER_66_41 ();
 sg13g2_fill_1 FILLER_66_55 ();
 sg13g2_fill_2 FILLER_66_78 ();
 sg13g2_fill_2 FILLER_66_94 ();
 sg13g2_fill_1 FILLER_66_96 ();
 sg13g2_fill_2 FILLER_66_154 ();
 sg13g2_decap_8 FILLER_66_170 ();
 sg13g2_fill_1 FILLER_66_177 ();
 sg13g2_fill_2 FILLER_66_191 ();
 sg13g2_fill_2 FILLER_66_201 ();
 sg13g2_fill_2 FILLER_66_235 ();
 sg13g2_decap_8 FILLER_66_250 ();
 sg13g2_decap_4 FILLER_66_257 ();
 sg13g2_fill_2 FILLER_66_265 ();
 sg13g2_fill_1 FILLER_66_267 ();
 sg13g2_decap_8 FILLER_66_277 ();
 sg13g2_decap_8 FILLER_66_284 ();
 sg13g2_fill_2 FILLER_66_291 ();
 sg13g2_decap_8 FILLER_66_319 ();
 sg13g2_fill_2 FILLER_66_326 ();
 sg13g2_fill_1 FILLER_66_328 ();
 sg13g2_fill_2 FILLER_66_337 ();
 sg13g2_decap_8 FILLER_66_382 ();
 sg13g2_fill_2 FILLER_66_389 ();
 sg13g2_decap_8 FILLER_66_400 ();
 sg13g2_decap_4 FILLER_66_407 ();
 sg13g2_fill_2 FILLER_66_411 ();
 sg13g2_fill_2 FILLER_66_423 ();
 sg13g2_fill_1 FILLER_66_425 ();
 sg13g2_fill_2 FILLER_66_442 ();
 sg13g2_fill_2 FILLER_66_470 ();
 sg13g2_fill_1 FILLER_66_472 ();
 sg13g2_fill_2 FILLER_66_499 ();
 sg13g2_fill_2 FILLER_66_531 ();
 sg13g2_fill_2 FILLER_66_558 ();
 sg13g2_fill_2 FILLER_66_575 ();
 sg13g2_decap_8 FILLER_66_587 ();
 sg13g2_fill_1 FILLER_66_594 ();
 sg13g2_fill_1 FILLER_66_607 ();
 sg13g2_fill_1 FILLER_66_614 ();
 sg13g2_decap_4 FILLER_66_619 ();
 sg13g2_fill_2 FILLER_66_623 ();
 sg13g2_fill_1 FILLER_66_712 ();
 sg13g2_decap_4 FILLER_66_732 ();
 sg13g2_decap_4 FILLER_66_741 ();
 sg13g2_fill_1 FILLER_66_745 ();
 sg13g2_decap_4 FILLER_66_750 ();
 sg13g2_fill_2 FILLER_66_765 ();
 sg13g2_fill_2 FILLER_66_799 ();
 sg13g2_fill_2 FILLER_66_810 ();
 sg13g2_fill_1 FILLER_66_812 ();
 sg13g2_decap_8 FILLER_66_826 ();
 sg13g2_decap_8 FILLER_66_833 ();
 sg13g2_decap_8 FILLER_66_840 ();
 sg13g2_decap_8 FILLER_66_847 ();
 sg13g2_decap_8 FILLER_66_854 ();
 sg13g2_fill_1 FILLER_66_861 ();
 sg13g2_fill_1 FILLER_67_31 ();
 sg13g2_fill_2 FILLER_67_181 ();
 sg13g2_fill_1 FILLER_67_193 ();
 sg13g2_fill_1 FILLER_67_218 ();
 sg13g2_fill_2 FILLER_67_234 ();
 sg13g2_decap_8 FILLER_67_276 ();
 sg13g2_decap_8 FILLER_67_283 ();
 sg13g2_decap_8 FILLER_67_294 ();
 sg13g2_decap_4 FILLER_67_301 ();
 sg13g2_fill_1 FILLER_67_305 ();
 sg13g2_fill_2 FILLER_67_350 ();
 sg13g2_fill_2 FILLER_67_371 ();
 sg13g2_fill_1 FILLER_67_385 ();
 sg13g2_decap_4 FILLER_67_391 ();
 sg13g2_fill_1 FILLER_67_395 ();
 sg13g2_fill_2 FILLER_67_459 ();
 sg13g2_fill_2 FILLER_67_481 ();
 sg13g2_fill_1 FILLER_67_538 ();
 sg13g2_fill_2 FILLER_67_550 ();
 sg13g2_fill_2 FILLER_67_556 ();
 sg13g2_fill_2 FILLER_67_573 ();
 sg13g2_fill_2 FILLER_67_592 ();
 sg13g2_fill_1 FILLER_67_594 ();
 sg13g2_fill_2 FILLER_67_623 ();
 sg13g2_decap_8 FILLER_67_634 ();
 sg13g2_fill_1 FILLER_67_667 ();
 sg13g2_fill_2 FILLER_67_695 ();
 sg13g2_fill_2 FILLER_67_710 ();
 sg13g2_fill_2 FILLER_67_746 ();
 sg13g2_fill_1 FILLER_67_748 ();
 sg13g2_fill_2 FILLER_67_775 ();
 sg13g2_fill_1 FILLER_67_777 ();
 sg13g2_fill_1 FILLER_67_810 ();
 sg13g2_decap_8 FILLER_67_837 ();
 sg13g2_decap_8 FILLER_67_844 ();
 sg13g2_decap_8 FILLER_67_851 ();
 sg13g2_decap_4 FILLER_67_858 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_4 ();
 sg13g2_fill_2 FILLER_68_23 ();
 sg13g2_fill_1 FILLER_68_25 ();
 sg13g2_fill_2 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_55 ();
 sg13g2_fill_1 FILLER_68_62 ();
 sg13g2_decap_4 FILLER_68_68 ();
 sg13g2_fill_2 FILLER_68_94 ();
 sg13g2_fill_2 FILLER_68_150 ();
 sg13g2_decap_8 FILLER_68_160 ();
 sg13g2_decap_4 FILLER_68_167 ();
 sg13g2_fill_1 FILLER_68_175 ();
 sg13g2_fill_1 FILLER_68_181 ();
 sg13g2_fill_2 FILLER_68_218 ();
 sg13g2_fill_1 FILLER_68_220 ();
 sg13g2_fill_2 FILLER_68_330 ();
 sg13g2_fill_2 FILLER_68_341 ();
 sg13g2_fill_2 FILLER_68_426 ();
 sg13g2_fill_2 FILLER_68_446 ();
 sg13g2_fill_1 FILLER_68_448 ();
 sg13g2_fill_1 FILLER_68_462 ();
 sg13g2_fill_1 FILLER_68_515 ();
 sg13g2_fill_2 FILLER_68_521 ();
 sg13g2_fill_1 FILLER_68_532 ();
 sg13g2_fill_2 FILLER_68_547 ();
 sg13g2_fill_2 FILLER_68_561 ();
 sg13g2_decap_8 FILLER_68_567 ();
 sg13g2_decap_4 FILLER_68_574 ();
 sg13g2_fill_1 FILLER_68_609 ();
 sg13g2_fill_2 FILLER_68_616 ();
 sg13g2_fill_1 FILLER_68_644 ();
 sg13g2_fill_2 FILLER_68_649 ();
 sg13g2_fill_1 FILLER_68_651 ();
 sg13g2_fill_2 FILLER_68_656 ();
 sg13g2_fill_1 FILLER_68_722 ();
 sg13g2_fill_1 FILLER_68_728 ();
 sg13g2_fill_2 FILLER_68_742 ();
 sg13g2_fill_2 FILLER_68_767 ();
 sg13g2_fill_2 FILLER_68_799 ();
 sg13g2_decap_8 FILLER_68_844 ();
 sg13g2_decap_8 FILLER_68_851 ();
 sg13g2_decap_4 FILLER_68_858 ();
 sg13g2_fill_2 FILLER_69_26 ();
 sg13g2_decap_8 FILLER_69_59 ();
 sg13g2_fill_1 FILLER_69_66 ();
 sg13g2_fill_1 FILLER_69_82 ();
 sg13g2_fill_2 FILLER_69_87 ();
 sg13g2_fill_2 FILLER_69_96 ();
 sg13g2_fill_1 FILLER_69_108 ();
 sg13g2_fill_2 FILLER_69_127 ();
 sg13g2_fill_2 FILLER_69_134 ();
 sg13g2_decap_8 FILLER_69_188 ();
 sg13g2_decap_4 FILLER_69_198 ();
 sg13g2_fill_1 FILLER_69_202 ();
 sg13g2_fill_1 FILLER_69_211 ();
 sg13g2_decap_4 FILLER_69_226 ();
 sg13g2_fill_1 FILLER_69_230 ();
 sg13g2_decap_4 FILLER_69_242 ();
 sg13g2_fill_2 FILLER_69_246 ();
 sg13g2_fill_1 FILLER_69_257 ();
 sg13g2_decap_4 FILLER_69_263 ();
 sg13g2_fill_1 FILLER_69_267 ();
 sg13g2_decap_8 FILLER_69_272 ();
 sg13g2_decap_8 FILLER_69_279 ();
 sg13g2_fill_2 FILLER_69_286 ();
 sg13g2_fill_1 FILLER_69_288 ();
 sg13g2_decap_4 FILLER_69_293 ();
 sg13g2_fill_2 FILLER_69_297 ();
 sg13g2_decap_4 FILLER_69_303 ();
 sg13g2_fill_1 FILLER_69_307 ();
 sg13g2_fill_2 FILLER_69_320 ();
 sg13g2_fill_1 FILLER_69_357 ();
 sg13g2_fill_1 FILLER_69_375 ();
 sg13g2_fill_1 FILLER_69_385 ();
 sg13g2_decap_8 FILLER_69_394 ();
 sg13g2_decap_8 FILLER_69_401 ();
 sg13g2_fill_2 FILLER_69_408 ();
 sg13g2_fill_1 FILLER_69_410 ();
 sg13g2_fill_1 FILLER_69_419 ();
 sg13g2_fill_2 FILLER_69_472 ();
 sg13g2_decap_8 FILLER_69_478 ();
 sg13g2_fill_2 FILLER_69_485 ();
 sg13g2_fill_1 FILLER_69_558 ();
 sg13g2_fill_1 FILLER_69_568 ();
 sg13g2_decap_4 FILLER_69_575 ();
 sg13g2_fill_1 FILLER_69_703 ();
 sg13g2_fill_1 FILLER_69_762 ();
 sg13g2_fill_1 FILLER_69_810 ();
 sg13g2_decap_8 FILLER_69_855 ();
 sg13g2_decap_4 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_37 ();
 sg13g2_fill_2 FILLER_70_75 ();
 sg13g2_fill_1 FILLER_70_77 ();
 sg13g2_fill_2 FILLER_70_91 ();
 sg13g2_fill_2 FILLER_70_105 ();
 sg13g2_fill_2 FILLER_70_122 ();
 sg13g2_fill_1 FILLER_70_127 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_fill_1 FILLER_70_161 ();
 sg13g2_fill_1 FILLER_70_175 ();
 sg13g2_fill_2 FILLER_70_189 ();
 sg13g2_fill_1 FILLER_70_191 ();
 sg13g2_fill_1 FILLER_70_259 ();
 sg13g2_fill_2 FILLER_70_407 ();
 sg13g2_fill_2 FILLER_70_418 ();
 sg13g2_fill_2 FILLER_70_459 ();
 sg13g2_decap_8 FILLER_70_542 ();
 sg13g2_decap_8 FILLER_70_549 ();
 sg13g2_fill_2 FILLER_70_556 ();
 sg13g2_fill_2 FILLER_70_566 ();
 sg13g2_fill_1 FILLER_70_568 ();
 sg13g2_decap_8 FILLER_70_574 ();
 sg13g2_decap_8 FILLER_70_581 ();
 sg13g2_fill_2 FILLER_70_588 ();
 sg13g2_fill_2 FILLER_70_594 ();
 sg13g2_fill_1 FILLER_70_596 ();
 sg13g2_fill_1 FILLER_70_648 ();
 sg13g2_fill_2 FILLER_70_668 ();
 sg13g2_fill_2 FILLER_70_696 ();
 sg13g2_fill_1 FILLER_70_698 ();
 sg13g2_fill_2 FILLER_70_743 ();
 sg13g2_fill_1 FILLER_70_745 ();
 sg13g2_fill_1 FILLER_70_798 ();
 sg13g2_fill_1 FILLER_70_814 ();
 sg13g2_decap_8 FILLER_70_850 ();
 sg13g2_decap_4 FILLER_70_857 ();
 sg13g2_fill_1 FILLER_70_861 ();
 sg13g2_fill_2 FILLER_71_89 ();
 sg13g2_fill_1 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_120 ();
 sg13g2_decap_4 FILLER_71_127 ();
 sg13g2_fill_2 FILLER_71_136 ();
 sg13g2_fill_1 FILLER_71_138 ();
 sg13g2_fill_2 FILLER_71_148 ();
 sg13g2_fill_1 FILLER_71_150 ();
 sg13g2_fill_1 FILLER_71_184 ();
 sg13g2_fill_2 FILLER_71_202 ();
 sg13g2_fill_1 FILLER_71_218 ();
 sg13g2_fill_2 FILLER_71_229 ();
 sg13g2_fill_2 FILLER_71_249 ();
 sg13g2_fill_1 FILLER_71_251 ();
 sg13g2_decap_4 FILLER_71_271 ();
 sg13g2_fill_1 FILLER_71_275 ();
 sg13g2_decap_8 FILLER_71_288 ();
 sg13g2_decap_8 FILLER_71_295 ();
 sg13g2_fill_2 FILLER_71_306 ();
 sg13g2_fill_1 FILLER_71_308 ();
 sg13g2_fill_1 FILLER_71_367 ();
 sg13g2_fill_2 FILLER_71_439 ();
 sg13g2_fill_1 FILLER_71_441 ();
 sg13g2_fill_1 FILLER_71_469 ();
 sg13g2_fill_1 FILLER_71_496 ();
 sg13g2_decap_4 FILLER_71_551 ();
 sg13g2_fill_2 FILLER_71_555 ();
 sg13g2_decap_4 FILLER_71_605 ();
 sg13g2_fill_2 FILLER_71_650 ();
 sg13g2_fill_2 FILLER_71_658 ();
 sg13g2_fill_1 FILLER_71_677 ();
 sg13g2_fill_2 FILLER_71_690 ();
 sg13g2_fill_1 FILLER_71_692 ();
 sg13g2_fill_1 FILLER_71_768 ();
 sg13g2_fill_2 FILLER_71_779 ();
 sg13g2_fill_1 FILLER_71_781 ();
 sg13g2_decap_8 FILLER_71_843 ();
 sg13g2_decap_8 FILLER_71_850 ();
 sg13g2_decap_4 FILLER_71_857 ();
 sg13g2_fill_1 FILLER_71_861 ();
 sg13g2_fill_2 FILLER_72_38 ();
 sg13g2_fill_2 FILLER_72_66 ();
 sg13g2_fill_1 FILLER_72_111 ();
 sg13g2_fill_2 FILLER_72_143 ();
 sg13g2_fill_1 FILLER_72_181 ();
 sg13g2_fill_2 FILLER_72_217 ();
 sg13g2_fill_2 FILLER_72_263 ();
 sg13g2_fill_1 FILLER_72_265 ();
 sg13g2_fill_2 FILLER_72_395 ();
 sg13g2_fill_1 FILLER_72_397 ();
 sg13g2_fill_2 FILLER_72_442 ();
 sg13g2_fill_1 FILLER_72_444 ();
 sg13g2_fill_1 FILLER_72_455 ();
 sg13g2_fill_2 FILLER_72_492 ();
 sg13g2_decap_4 FILLER_72_520 ();
 sg13g2_fill_1 FILLER_72_553 ();
 sg13g2_fill_1 FILLER_72_581 ();
 sg13g2_fill_2 FILLER_72_586 ();
 sg13g2_fill_2 FILLER_72_609 ();
 sg13g2_decap_4 FILLER_72_615 ();
 sg13g2_fill_1 FILLER_72_619 ();
 sg13g2_fill_1 FILLER_72_665 ();
 sg13g2_fill_2 FILLER_72_728 ();
 sg13g2_fill_1 FILLER_72_730 ();
 sg13g2_fill_2 FILLER_72_735 ();
 sg13g2_fill_1 FILLER_72_737 ();
 sg13g2_fill_1 FILLER_72_753 ();
 sg13g2_fill_2 FILLER_72_763 ();
 sg13g2_fill_2 FILLER_72_810 ();
 sg13g2_decap_8 FILLER_72_842 ();
 sg13g2_decap_8 FILLER_72_849 ();
 sg13g2_decap_4 FILLER_72_856 ();
 sg13g2_fill_2 FILLER_72_860 ();
 sg13g2_decap_4 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_4 ();
 sg13g2_fill_2 FILLER_73_18 ();
 sg13g2_decap_4 FILLER_73_54 ();
 sg13g2_fill_2 FILLER_73_58 ();
 sg13g2_fill_1 FILLER_73_92 ();
 sg13g2_fill_2 FILLER_73_102 ();
 sg13g2_fill_1 FILLER_73_127 ();
 sg13g2_fill_1 FILLER_73_153 ();
 sg13g2_fill_1 FILLER_73_197 ();
 sg13g2_fill_2 FILLER_73_203 ();
 sg13g2_fill_2 FILLER_73_218 ();
 sg13g2_fill_1 FILLER_73_246 ();
 sg13g2_fill_1 FILLER_73_277 ();
 sg13g2_fill_2 FILLER_73_287 ();
 sg13g2_fill_2 FILLER_73_299 ();
 sg13g2_fill_2 FILLER_73_309 ();
 sg13g2_fill_2 FILLER_73_315 ();
 sg13g2_fill_1 FILLER_73_317 ();
 sg13g2_fill_2 FILLER_73_348 ();
 sg13g2_fill_2 FILLER_73_376 ();
 sg13g2_fill_2 FILLER_73_408 ();
 sg13g2_fill_2 FILLER_73_416 ();
 sg13g2_fill_1 FILLER_73_488 ();
 sg13g2_fill_2 FILLER_73_508 ();
 sg13g2_decap_4 FILLER_73_513 ();
 sg13g2_fill_2 FILLER_73_517 ();
 sg13g2_fill_1 FILLER_73_552 ();
 sg13g2_fill_1 FILLER_73_593 ();
 sg13g2_fill_1 FILLER_73_705 ();
 sg13g2_fill_2 FILLER_73_723 ();
 sg13g2_fill_2 FILLER_73_784 ();
 sg13g2_decap_8 FILLER_73_841 ();
 sg13g2_decap_8 FILLER_73_848 ();
 sg13g2_decap_8 FILLER_73_855 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_4 FILLER_74_7 ();
 sg13g2_fill_1 FILLER_74_15 ();
 sg13g2_fill_2 FILLER_74_40 ();
 sg13g2_fill_1 FILLER_74_158 ();
 sg13g2_fill_2 FILLER_74_190 ();
 sg13g2_fill_1 FILLER_74_223 ();
 sg13g2_fill_1 FILLER_74_255 ();
 sg13g2_fill_1 FILLER_74_278 ();
 sg13g2_fill_1 FILLER_74_288 ();
 sg13g2_fill_2 FILLER_74_375 ();
 sg13g2_fill_1 FILLER_74_377 ();
 sg13g2_fill_1 FILLER_74_386 ();
 sg13g2_fill_2 FILLER_74_413 ();
 sg13g2_fill_2 FILLER_74_429 ();
 sg13g2_fill_1 FILLER_74_431 ();
 sg13g2_fill_1 FILLER_74_558 ();
 sg13g2_fill_2 FILLER_74_568 ();
 sg13g2_fill_1 FILLER_74_611 ();
 sg13g2_fill_1 FILLER_74_625 ();
 sg13g2_fill_2 FILLER_74_631 ();
 sg13g2_fill_2 FILLER_74_750 ();
 sg13g2_fill_1 FILLER_74_752 ();
 sg13g2_decap_8 FILLER_74_841 ();
 sg13g2_decap_8 FILLER_74_848 ();
 sg13g2_decap_8 FILLER_74_855 ();
 sg13g2_fill_2 FILLER_75_39 ();
 sg13g2_decap_4 FILLER_75_59 ();
 sg13g2_fill_2 FILLER_75_145 ();
 sg13g2_fill_1 FILLER_75_147 ();
 sg13g2_fill_1 FILLER_75_156 ();
 sg13g2_fill_1 FILLER_75_169 ();
 sg13g2_fill_2 FILLER_75_200 ();
 sg13g2_fill_1 FILLER_75_202 ();
 sg13g2_fill_2 FILLER_75_212 ();
 sg13g2_fill_1 FILLER_75_214 ();
 sg13g2_fill_1 FILLER_75_289 ();
 sg13g2_fill_1 FILLER_75_299 ();
 sg13g2_fill_1 FILLER_75_361 ();
 sg13g2_fill_2 FILLER_75_371 ();
 sg13g2_fill_1 FILLER_75_373 ();
 sg13g2_fill_1 FILLER_75_382 ();
 sg13g2_fill_1 FILLER_75_397 ();
 sg13g2_fill_1 FILLER_75_403 ();
 sg13g2_fill_2 FILLER_75_430 ();
 sg13g2_fill_1 FILLER_75_432 ();
 sg13g2_fill_2 FILLER_75_442 ();
 sg13g2_fill_1 FILLER_75_444 ();
 sg13g2_fill_2 FILLER_75_452 ();
 sg13g2_fill_2 FILLER_75_495 ();
 sg13g2_fill_2 FILLER_75_502 ();
 sg13g2_fill_2 FILLER_75_541 ();
 sg13g2_fill_1 FILLER_75_567 ();
 sg13g2_fill_1 FILLER_75_587 ();
 sg13g2_fill_1 FILLER_75_646 ();
 sg13g2_decap_8 FILLER_75_831 ();
 sg13g2_decap_8 FILLER_75_838 ();
 sg13g2_decap_8 FILLER_75_845 ();
 sg13g2_decap_8 FILLER_75_852 ();
 sg13g2_fill_2 FILLER_75_859 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_decap_4 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_4 ();
 sg13g2_fill_1 FILLER_76_21 ();
 sg13g2_fill_1 FILLER_76_37 ();
 sg13g2_decap_4 FILLER_76_64 ();
 sg13g2_fill_2 FILLER_76_68 ();
 sg13g2_fill_1 FILLER_76_178 ();
 sg13g2_fill_2 FILLER_76_231 ();
 sg13g2_fill_1 FILLER_76_250 ();
 sg13g2_fill_1 FILLER_76_266 ();
 sg13g2_fill_2 FILLER_76_299 ();
 sg13g2_fill_1 FILLER_76_331 ();
 sg13g2_fill_2 FILLER_76_416 ();
 sg13g2_fill_2 FILLER_76_427 ();
 sg13g2_fill_1 FILLER_76_429 ();
 sg13g2_fill_2 FILLER_76_449 ();
 sg13g2_fill_1 FILLER_76_457 ();
 sg13g2_fill_2 FILLER_76_517 ();
 sg13g2_fill_2 FILLER_76_564 ();
 sg13g2_fill_1 FILLER_76_654 ();
 sg13g2_fill_1 FILLER_76_688 ();
 sg13g2_fill_1 FILLER_76_725 ();
 sg13g2_decap_8 FILLER_76_835 ();
 sg13g2_decap_8 FILLER_76_842 ();
 sg13g2_decap_8 FILLER_76_849 ();
 sg13g2_decap_4 FILLER_76_856 ();
 sg13g2_fill_2 FILLER_76_860 ();
 sg13g2_fill_1 FILLER_77_36 ();
 sg13g2_fill_1 FILLER_77_42 ();
 sg13g2_fill_2 FILLER_77_52 ();
 sg13g2_fill_1 FILLER_77_68 ();
 sg13g2_fill_1 FILLER_77_134 ();
 sg13g2_fill_2 FILLER_77_153 ();
 sg13g2_fill_2 FILLER_77_168 ();
 sg13g2_fill_2 FILLER_77_179 ();
 sg13g2_fill_1 FILLER_77_215 ();
 sg13g2_fill_1 FILLER_77_226 ();
 sg13g2_fill_1 FILLER_77_261 ();
 sg13g2_fill_1 FILLER_77_267 ();
 sg13g2_fill_1 FILLER_77_400 ();
 sg13g2_fill_2 FILLER_77_413 ();
 sg13g2_fill_1 FILLER_77_415 ();
 sg13g2_fill_1 FILLER_77_426 ();
 sg13g2_fill_1 FILLER_77_482 ();
 sg13g2_fill_2 FILLER_77_492 ();
 sg13g2_fill_2 FILLER_77_518 ();
 sg13g2_fill_2 FILLER_77_559 ();
 sg13g2_fill_1 FILLER_77_620 ();
 sg13g2_fill_2 FILLER_77_798 ();
 sg13g2_fill_1 FILLER_77_800 ();
 sg13g2_decap_8 FILLER_77_827 ();
 sg13g2_decap_8 FILLER_77_834 ();
 sg13g2_decap_8 FILLER_77_841 ();
 sg13g2_decap_8 FILLER_77_848 ();
 sg13g2_decap_8 FILLER_77_855 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_7 ();
 sg13g2_fill_1 FILLER_78_26 ();
 sg13g2_fill_2 FILLER_78_36 ();
 sg13g2_fill_1 FILLER_78_47 ();
 sg13g2_fill_2 FILLER_78_53 ();
 sg13g2_fill_2 FILLER_78_60 ();
 sg13g2_fill_1 FILLER_78_65 ();
 sg13g2_fill_2 FILLER_78_70 ();
 sg13g2_fill_1 FILLER_78_72 ();
 sg13g2_fill_1 FILLER_78_105 ();
 sg13g2_decap_4 FILLER_78_113 ();
 sg13g2_fill_2 FILLER_78_117 ();
 sg13g2_fill_1 FILLER_78_190 ();
 sg13g2_fill_1 FILLER_78_262 ();
 sg13g2_fill_2 FILLER_78_271 ();
 sg13g2_fill_2 FILLER_78_287 ();
 sg13g2_fill_1 FILLER_78_341 ();
 sg13g2_fill_2 FILLER_78_384 ();
 sg13g2_fill_2 FILLER_78_403 ();
 sg13g2_fill_1 FILLER_78_405 ();
 sg13g2_fill_1 FILLER_78_439 ();
 sg13g2_fill_1 FILLER_78_528 ();
 sg13g2_fill_2 FILLER_78_547 ();
 sg13g2_fill_1 FILLER_78_553 ();
 sg13g2_fill_1 FILLER_78_585 ();
 sg13g2_fill_1 FILLER_78_613 ();
 sg13g2_fill_2 FILLER_78_623 ();
 sg13g2_fill_2 FILLER_78_634 ();
 sg13g2_fill_2 FILLER_78_756 ();
 sg13g2_fill_1 FILLER_78_783 ();
 sg13g2_fill_1 FILLER_78_788 ();
 sg13g2_fill_1 FILLER_78_793 ();
 sg13g2_decap_8 FILLER_78_823 ();
 sg13g2_decap_8 FILLER_78_830 ();
 sg13g2_decap_8 FILLER_78_837 ();
 sg13g2_decap_8 FILLER_78_844 ();
 sg13g2_decap_8 FILLER_78_851 ();
 sg13g2_decap_4 FILLER_78_858 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_4 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_11 ();
 sg13g2_fill_1 FILLER_79_38 ();
 sg13g2_fill_2 FILLER_79_44 ();
 sg13g2_fill_2 FILLER_79_53 ();
 sg13g2_fill_1 FILLER_79_81 ();
 sg13g2_decap_4 FILLER_79_89 ();
 sg13g2_fill_2 FILLER_79_93 ();
 sg13g2_decap_8 FILLER_79_100 ();
 sg13g2_decap_4 FILLER_79_107 ();
 sg13g2_fill_2 FILLER_79_111 ();
 sg13g2_fill_1 FILLER_79_171 ();
 sg13g2_fill_2 FILLER_79_224 ();
 sg13g2_fill_2 FILLER_79_262 ();
 sg13g2_fill_1 FILLER_79_387 ();
 sg13g2_fill_2 FILLER_79_450 ();
 sg13g2_fill_1 FILLER_79_499 ();
 sg13g2_fill_2 FILLER_79_559 ();
 sg13g2_fill_1 FILLER_79_570 ();
 sg13g2_fill_2 FILLER_79_655 ();
 sg13g2_fill_1 FILLER_79_657 ();
 sg13g2_fill_2 FILLER_79_710 ();
 sg13g2_fill_1 FILLER_79_749 ();
 sg13g2_decap_8 FILLER_79_784 ();
 sg13g2_decap_8 FILLER_79_791 ();
 sg13g2_decap_8 FILLER_79_798 ();
 sg13g2_decap_8 FILLER_79_805 ();
 sg13g2_decap_8 FILLER_79_816 ();
 sg13g2_decap_8 FILLER_79_823 ();
 sg13g2_decap_8 FILLER_79_830 ();
 sg13g2_decap_8 FILLER_79_837 ();
 sg13g2_decap_8 FILLER_79_844 ();
 sg13g2_decap_8 FILLER_79_851 ();
 sg13g2_decap_4 FILLER_79_858 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_fill_2 FILLER_80_21 ();
 sg13g2_decap_4 FILLER_80_27 ();
 sg13g2_fill_1 FILLER_80_31 ();
 sg13g2_fill_2 FILLER_80_70 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_fill_2 FILLER_80_159 ();
 sg13g2_fill_1 FILLER_80_161 ();
 sg13g2_fill_1 FILLER_80_235 ();
 sg13g2_fill_1 FILLER_80_272 ();
 sg13g2_fill_1 FILLER_80_302 ();
 sg13g2_fill_2 FILLER_80_334 ();
 sg13g2_fill_2 FILLER_80_428 ();
 sg13g2_fill_1 FILLER_80_430 ();
 sg13g2_fill_1 FILLER_80_448 ();
 sg13g2_fill_1 FILLER_80_483 ();
 sg13g2_fill_1 FILLER_80_522 ();
 sg13g2_fill_2 FILLER_80_536 ();
 sg13g2_fill_1 FILLER_80_594 ();
 sg13g2_fill_2 FILLER_80_656 ();
 sg13g2_fill_1 FILLER_80_671 ();
 sg13g2_fill_2 FILLER_80_701 ();
 sg13g2_decap_8 FILLER_80_765 ();
 sg13g2_decap_8 FILLER_80_772 ();
 sg13g2_decap_8 FILLER_80_779 ();
 sg13g2_decap_8 FILLER_80_786 ();
 sg13g2_decap_8 FILLER_80_793 ();
 sg13g2_decap_8 FILLER_80_800 ();
 sg13g2_decap_8 FILLER_80_807 ();
 sg13g2_decap_8 FILLER_80_814 ();
 sg13g2_decap_8 FILLER_80_821 ();
 sg13g2_decap_8 FILLER_80_828 ();
 sg13g2_decap_8 FILLER_80_835 ();
 sg13g2_decap_8 FILLER_80_842 ();
 sg13g2_decap_8 FILLER_80_849 ();
 sg13g2_decap_4 FILLER_80_856 ();
 sg13g2_fill_2 FILLER_80_860 ();
 assign uio_oe[0] = net603;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net604;
 assign uio_oe[3] = net605;
 assign uio_oe[4] = net606;
 assign uio_oe[5] = net4;
 assign uio_oe[6] = net5;
 assign uio_oe[7] = net6;
 assign uio_out[1] = net7;
 assign uio_out[4] = net8;
 assign uio_out[6] = net9;
 assign uio_out[7] = net10;
endmodule

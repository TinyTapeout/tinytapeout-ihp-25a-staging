module tt_um_save_buffer_hash_table (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire \tb.cursor[0] ;
 wire \tb.cursor[1] ;
 wire \tb.cursor[2] ;
 wire \tb.cursor[3] ;
 wire \tb.go_ok ;
 wire \tb.hash_saved[0] ;
 wire \tb.hash_saved[1] ;
 wire \tb.hash_saved[2] ;
 wire \tb.key_saved[0] ;
 wire \tb.key_saved[1] ;
 wire \tb.key_saved[2] ;
 wire \tb.key_saved[3] ;
 wire \tb.mem[0][0] ;
 wire \tb.mem[0][1] ;
 wire \tb.mem[0][2] ;
 wire \tb.mem[0][3] ;
 wire \tb.mem[0][4] ;
 wire \tb.mem[0][5] ;
 wire \tb.mem[0][6] ;
 wire \tb.mem[0][7] ;
 wire \tb.mem[0][8] ;
 wire \tb.mem[1][0] ;
 wire \tb.mem[1][1] ;
 wire \tb.mem[1][2] ;
 wire \tb.mem[1][3] ;
 wire \tb.mem[1][4] ;
 wire \tb.mem[1][5] ;
 wire \tb.mem[1][6] ;
 wire \tb.mem[1][7] ;
 wire \tb.mem[1][8] ;
 wire \tb.mem[2][0] ;
 wire \tb.mem[2][1] ;
 wire \tb.mem[2][2] ;
 wire \tb.mem[2][3] ;
 wire \tb.mem[2][4] ;
 wire \tb.mem[2][5] ;
 wire \tb.mem[2][6] ;
 wire \tb.mem[2][7] ;
 wire \tb.mem[2][8] ;
 wire \tb.mem[3][0] ;
 wire \tb.mem[3][1] ;
 wire \tb.mem[3][2] ;
 wire \tb.mem[3][3] ;
 wire \tb.mem[3][4] ;
 wire \tb.mem[3][5] ;
 wire \tb.mem[3][6] ;
 wire \tb.mem[3][7] ;
 wire \tb.mem[3][8] ;
 wire \tb.mem[4][0] ;
 wire \tb.mem[4][1] ;
 wire \tb.mem[4][2] ;
 wire \tb.mem[4][3] ;
 wire \tb.mem[4][4] ;
 wire \tb.mem[4][5] ;
 wire \tb.mem[4][6] ;
 wire \tb.mem[4][7] ;
 wire \tb.mem[4][8] ;
 wire \tb.mem[5][0] ;
 wire \tb.mem[5][1] ;
 wire \tb.mem[5][2] ;
 wire \tb.mem[5][3] ;
 wire \tb.mem[5][4] ;
 wire \tb.mem[5][5] ;
 wire \tb.mem[5][6] ;
 wire \tb.mem[5][7] ;
 wire \tb.mem[5][8] ;
 wire \tb.mem[6][0] ;
 wire \tb.mem[6][1] ;
 wire \tb.mem[6][2] ;
 wire \tb.mem[6][3] ;
 wire \tb.mem[6][4] ;
 wire \tb.mem[6][5] ;
 wire \tb.mem[6][6] ;
 wire \tb.mem[6][7] ;
 wire \tb.mem[6][8] ;
 wire \tb.mem[7][0] ;
 wire \tb.mem[7][1] ;
 wire \tb.mem[7][2] ;
 wire \tb.mem[7][3] ;
 wire \tb.mem[7][4] ;
 wire \tb.mem[7][5] ;
 wire \tb.mem[7][6] ;
 wire \tb.mem[7][7] ;
 wire \tb.mem[7][8] ;
 wire \tb.state ;
 wire \tb.val_saved[0] ;
 wire \tb.val_saved[1] ;
 wire \tb.val_saved[2] ;
 wire \tb.val_saved[3] ;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net167;
 wire clknet_0_clk;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;

 sg13g2_inv_1 _0597_ (.Y(_0103_),
    .A(net4));
 sg13g2_inv_1 _0598_ (.Y(_0104_),
    .A(net3));
 sg13g2_inv_1 _0599_ (.Y(_0105_),
    .A(net2));
 sg13g2_inv_1 _0600_ (.Y(_0106_),
    .A(net1));
 sg13g2_inv_1 _0601_ (.Y(_0107_),
    .A(net8));
 sg13g2_inv_1 _0602_ (.Y(_0108_),
    .A(net7));
 sg13g2_inv_1 _0603_ (.Y(_0109_),
    .A(net6));
 sg13g2_inv_1 _0604_ (.Y(_0110_),
    .A(net5));
 sg13g2_inv_1 _0605_ (.Y(_0111_),
    .A(net282));
 sg13g2_inv_1 _0606_ (.Y(_0112_),
    .A(net140));
 sg13g2_inv_1 _0607_ (.Y(_0113_),
    .A(net141));
 sg13g2_inv_1 _0608_ (.Y(_0114_),
    .A(net285));
 sg13g2_inv_1 _0609_ (.Y(_0115_),
    .A(net284));
 sg13g2_inv_1 _0610_ (.Y(_0116_),
    .A(net286));
 sg13g2_inv_1 _0611_ (.Y(_0117_),
    .A(net287));
 sg13g2_inv_1 _0612_ (.Y(_0118_),
    .A(net142));
 sg13g2_inv_1 _0613_ (.Y(_0119_),
    .A(net146));
 sg13g2_inv_1 _0614_ (.Y(_0120_),
    .A(net234));
 sg13g2_inv_1 _0615_ (.Y(_0121_),
    .A(net221));
 sg13g2_inv_1 _0616_ (.Y(_0122_),
    .A(net178));
 sg13g2_inv_1 _0617_ (.Y(_0123_),
    .A(net182));
 sg13g2_inv_1 _0618_ (.Y(_0124_),
    .A(net242));
 sg13g2_inv_1 _0619_ (.Y(_0125_),
    .A(net277));
 sg13g2_inv_1 _0620_ (.Y(_0126_),
    .A(net271));
 sg13g2_inv_1 _0621_ (.Y(_0127_),
    .A(net255));
 sg13g2_inv_1 _0622_ (.Y(_0128_),
    .A(net248));
 sg13g2_inv_1 _0623_ (.Y(_0129_),
    .A(net175));
 sg13g2_inv_1 _0624_ (.Y(_0130_),
    .A(net190));
 sg13g2_inv_1 _0625_ (.Y(_0131_),
    .A(net218));
 sg13g2_inv_1 _0626_ (.Y(_0132_),
    .A(net258));
 sg13g2_inv_1 _0627_ (.Y(_0133_),
    .A(net253));
 sg13g2_inv_1 _0628_ (.Y(_0134_),
    .A(net172));
 sg13g2_inv_1 _0629_ (.Y(_0135_),
    .A(net180));
 sg13g2_inv_1 _0630_ (.Y(_0136_),
    .A(net236));
 sg13g2_inv_1 _0631_ (.Y(_0137_),
    .A(net214));
 sg13g2_inv_1 _0632_ (.Y(_0138_),
    .A(net251));
 sg13g2_inv_1 _0633_ (.Y(_0139_),
    .A(net223));
 sg13g2_inv_1 _0634_ (.Y(_0140_),
    .A(net228));
 sg13g2_inv_1 _0635_ (.Y(_0141_),
    .A(net232));
 sg13g2_inv_1 _0636_ (.Y(_0142_),
    .A(net273));
 sg13g2_inv_1 _0637_ (.Y(_0143_),
    .A(net226));
 sg13g2_inv_1 _0638_ (.Y(_0144_),
    .A(net275));
 sg13g2_inv_1 _0639_ (.Y(_0145_),
    .A(net244));
 sg13g2_inv_1 _0640_ (.Y(_0146_),
    .A(net212));
 sg13g2_inv_1 _0641_ (.Y(_0147_),
    .A(net210));
 sg13g2_inv_1 _0642_ (.Y(_0148_),
    .A(net240));
 sg13g2_inv_1 _0643_ (.Y(_0149_),
    .A(net230));
 sg13g2_inv_1 _0644_ (.Y(_0150_),
    .A(net187));
 sg13g2_inv_1 _0645_ (.Y(_0151_),
    .A(net184));
 sg13g2_inv_2 _0646_ (.Y(_0152_),
    .A(net152));
 sg13g2_inv_1 _0647_ (.Y(_0153_),
    .A(net199));
 sg13g2_inv_1 _0648_ (.Y(_0154_),
    .A(net225));
 sg13g2_inv_1 _0649_ (.Y(_0155_),
    .A(net194));
 sg13g2_inv_1 _0650_ (.Y(_0156_),
    .A(\tb.mem[3][0] ));
 sg13g2_inv_1 _0651_ (.Y(_0157_),
    .A(net204));
 sg13g2_inv_1 _0652_ (.Y(_0158_),
    .A(net192));
 sg13g2_inv_1 _0653_ (.Y(_0159_),
    .A(net250));
 sg13g2_inv_1 _0654_ (.Y(_0160_),
    .A(net262));
 sg13g2_inv_1 _0655_ (.Y(_0161_),
    .A(net246));
 sg13g2_inv_1 _0656_ (.Y(_0162_),
    .A(net207));
 sg13g2_inv_1 _0657_ (.Y(_0163_),
    .A(net238));
 sg13g2_inv_1 _0658_ (.Y(_0164_),
    .A(net201));
 sg13g2_inv_1 _0659_ (.Y(_0165_),
    .A(net269));
 sg13g2_inv_1 _0660_ (.Y(_0166_),
    .A(net196));
 sg13g2_inv_1 _0661_ (.Y(_0167_),
    .A(net267));
 sg13g2_inv_1 _0662_ (.Y(_0168_),
    .A(net263));
 sg13g2_inv_1 _0663_ (.Y(_0169_),
    .A(net257));
 sg13g2_inv_1 _0664_ (.Y(_0170_),
    .A(net206));
 sg13g2_inv_1 _0665_ (.Y(_0171_),
    .A(net220));
 sg13g2_inv_1 _0666_ (.Y(_0172_),
    .A(\tb.mem[3][2] ));
 sg13g2_inv_1 _0667_ (.Y(_0173_),
    .A(net198));
 sg13g2_inv_1 _0668_ (.Y(_0174_),
    .A(net209));
 sg13g2_inv_1 _0669_ (.Y(_0175_),
    .A(net203));
 sg13g2_inv_1 _0670_ (.Y(_0176_),
    .A(net189));
 sg13g2_inv_1 _0671_ (.Y(_0177_),
    .A(\tb.mem[0][3] ));
 sg13g2_inv_1 _0672_ (.Y(_0178_),
    .A(net260));
 sg13g2_inv_1 _0673_ (.Y(_0179_),
    .A(net261));
 sg13g2_inv_1 _0674_ (.Y(_0180_),
    .A(net265));
 sg13g2_inv_1 _0675_ (.Y(_0181_),
    .A(net174));
 sg13g2_inv_1 _0676_ (.Y(_0182_),
    .A(net186));
 sg13g2_inv_1 _0677_ (.Y(_0183_),
    .A(net177));
 sg13g2_inv_1 _0678_ (.Y(_0184_),
    .A(net266));
 sg13g2_nand2b_2 _0679_ (.Y(_0185_),
    .B(net9),
    .A_N(net10));
 sg13g2_mux4_1 _0680_ (.S0(net150),
    .A0(\tb.mem[0][5] ),
    .A1(\tb.mem[1][5] ),
    .A2(\tb.mem[2][5] ),
    .A3(\tb.mem[3][5] ),
    .S1(net146),
    .X(_0186_));
 sg13g2_mux4_1 _0681_ (.S0(net150),
    .A0(\tb.mem[4][5] ),
    .A1(\tb.mem[5][5] ),
    .A2(\tb.mem[6][5] ),
    .A3(\tb.mem[7][5] ),
    .S1(net147),
    .X(_0187_));
 sg13g2_mux2_1 _0682_ (.A0(_0186_),
    .A1(_0187_),
    .S(net143),
    .X(_0188_));
 sg13g2_xnor2_1 _0683_ (.Y(_0189_),
    .A(net138),
    .B(_0188_));
 sg13g2_mux4_1 _0684_ (.S0(net150),
    .A0(\tb.mem[0][4] ),
    .A1(\tb.mem[1][4] ),
    .A2(\tb.mem[2][4] ),
    .A3(\tb.mem[3][4] ),
    .S1(net147),
    .X(_0190_));
 sg13g2_mux4_1 _0685_ (.S0(net150),
    .A0(\tb.mem[4][4] ),
    .A1(\tb.mem[5][4] ),
    .A2(\tb.mem[6][4] ),
    .A3(\tb.mem[7][4] ),
    .S1(net145),
    .X(_0191_));
 sg13g2_mux2_1 _0686_ (.A0(_0190_),
    .A1(_0191_),
    .S(net143),
    .X(_0192_));
 sg13g2_xnor2_1 _0687_ (.Y(_0193_),
    .A(net139),
    .B(_0192_));
 sg13g2_mux4_1 _0688_ (.S0(net150),
    .A0(\tb.mem[0][6] ),
    .A1(\tb.mem[1][6] ),
    .A2(\tb.mem[2][6] ),
    .A3(\tb.mem[3][6] ),
    .S1(net146),
    .X(_0194_));
 sg13g2_mux4_1 _0689_ (.S0(net148),
    .A0(\tb.mem[4][6] ),
    .A1(\tb.mem[5][6] ),
    .A2(\tb.mem[6][6] ),
    .A3(\tb.mem[7][6] ),
    .S1(net145),
    .X(_0195_));
 sg13g2_mux2_1 _0690_ (.A0(_0194_),
    .A1(_0195_),
    .S(net143),
    .X(_0196_));
 sg13g2_xnor2_1 _0691_ (.Y(_0197_),
    .A(\tb.key_saved[2] ),
    .B(_0196_));
 sg13g2_mux4_1 _0692_ (.S0(net148),
    .A0(\tb.mem[4][7] ),
    .A1(\tb.mem[5][7] ),
    .A2(\tb.mem[6][7] ),
    .A3(\tb.mem[7][7] ),
    .S1(net145),
    .X(_0198_));
 sg13g2_mux4_1 _0693_ (.S0(net149),
    .A0(\tb.mem[0][7] ),
    .A1(\tb.mem[1][7] ),
    .A2(\tb.mem[2][7] ),
    .A3(\tb.mem[3][7] ),
    .S1(net146),
    .X(_0199_));
 sg13g2_mux2_1 _0694_ (.A0(_0199_),
    .A1(_0198_),
    .S(net143),
    .X(_0200_));
 sg13g2_xnor2_1 _0695_ (.Y(_0201_),
    .A(\tb.key_saved[3] ),
    .B(_0200_));
 sg13g2_nand4_1 _0696_ (.B(_0193_),
    .C(_0197_),
    .A(_0189_),
    .Y(_0202_),
    .D(_0201_));
 sg13g2_mux2_1 _0697_ (.A0(\tb.mem[4][8] ),
    .A1(\tb.mem[5][8] ),
    .S(net148),
    .X(_0203_));
 sg13g2_nor2b_1 _0698_ (.A(\tb.mem[7][8] ),
    .B_N(net150),
    .Y(_0204_));
 sg13g2_o21ai_1 _0699_ (.B1(net145),
    .Y(_0205_),
    .A1(net148),
    .A2(\tb.mem[6][8] ));
 sg13g2_o21ai_1 _0700_ (.B1(net144),
    .Y(_0206_),
    .A1(_0204_),
    .A2(_0205_));
 sg13g2_a21oi_1 _0701_ (.A1(_0119_),
    .A2(_0203_),
    .Y(_0207_),
    .B1(_0206_));
 sg13g2_mux2_1 _0702_ (.A0(\tb.mem[0][8] ),
    .A1(\tb.mem[1][8] ),
    .S(net149),
    .X(_0208_));
 sg13g2_nand2b_1 _0703_ (.Y(_0209_),
    .B(net149),
    .A_N(\tb.mem[3][8] ));
 sg13g2_nor2_1 _0704_ (.A(net149),
    .B(\tb.mem[2][8] ),
    .Y(_0210_));
 sg13g2_nor2_1 _0705_ (.A(_0119_),
    .B(_0210_),
    .Y(_0211_));
 sg13g2_a221oi_1 _0706_ (.B2(_0211_),
    .C1(net144),
    .B1(_0209_),
    .A1(_0119_),
    .Y(_0212_),
    .A2(_0208_));
 sg13g2_nor2_1 _0707_ (.A(_0207_),
    .B(_0212_),
    .Y(_0213_));
 sg13g2_a21oi_1 _0708_ (.A1(_0202_),
    .A2(_0213_),
    .Y(_0214_),
    .B1(_0185_));
 sg13g2_a21o_1 _0709_ (.A2(_0213_),
    .A1(_0202_),
    .B1(_0185_),
    .X(_0215_));
 sg13g2_nand2b_1 _0710_ (.Y(_0216_),
    .B(\tb.cursor[2] ),
    .A_N(\tb.hash_saved[2] ));
 sg13g2_a21o_1 _0711_ (.A2(_0112_),
    .A1(\tb.hash_saved[2] ),
    .B1(_0111_),
    .X(_0217_));
 sg13g2_xor2_1 _0712_ (.B(\tb.cursor[0] ),
    .A(\tb.hash_saved[0] ),
    .X(_0218_));
 sg13g2_nor2b_1 _0713_ (.A(net141),
    .B_N(\tb.hash_saved[1] ),
    .Y(_0219_));
 sg13g2_o21ai_1 _0714_ (.B1(_0216_),
    .Y(_0220_),
    .A1(\tb.hash_saved[1] ),
    .A2(_0113_));
 sg13g2_nor4_2 _0715_ (.A(_0217_),
    .B(_0218_),
    .C(_0219_),
    .Y(_0221_),
    .D(_0220_));
 sg13g2_inv_1 _0716_ (.Y(_0222_),
    .A(_0221_));
 sg13g2_nor2_2 _0717_ (.A(_0004_),
    .B(_0221_),
    .Y(_0223_));
 sg13g2_or2_2 _0718_ (.X(_0224_),
    .B(_0221_),
    .A(_0004_));
 sg13g2_nand3_1 _0719_ (.B(net141),
    .C(_0003_),
    .A(net140),
    .Y(_0225_));
 sg13g2_nor4_2 _0720_ (.A(_0152_),
    .B(_0215_),
    .C(_0224_),
    .Y(_0226_),
    .D(_0225_));
 sg13g2_nor4_2 _0721_ (.A(net9),
    .B(_0202_),
    .C(_0207_),
    .Y(_0227_),
    .D(_0212_));
 sg13g2_and3_2 _0722_ (.X(_0228_),
    .A(net10),
    .B(_0223_),
    .C(_0227_));
 sg13g2_nand2b_1 _0723_ (.Y(_0229_),
    .B(_0228_),
    .A_N(_0225_));
 sg13g2_and2_1 _0724_ (.A(net304),
    .B(net151),
    .X(_0230_));
 sg13g2_a21o_1 _0725_ (.A2(_0230_),
    .A1(_0229_),
    .B1(net126),
    .X(_0005_));
 sg13g2_nor2_1 _0726_ (.A(\tb.cursor[1] ),
    .B(\tb.cursor[0] ),
    .Y(_0231_));
 sg13g2_nand2_1 _0727_ (.Y(_0232_),
    .A(net140),
    .B(_0231_));
 sg13g2_nor4_2 _0728_ (.A(_0152_),
    .B(_0215_),
    .C(_0224_),
    .Y(_0233_),
    .D(_0232_));
 sg13g2_nand2_1 _0729_ (.Y(_0234_),
    .A(net135),
    .B(net125));
 sg13g2_nand2b_2 _0730_ (.Y(_0235_),
    .B(net151),
    .A_N(net125));
 sg13g2_o21ai_1 _0731_ (.B1(_0234_),
    .Y(_0006_),
    .A1(_0157_),
    .A2(_0235_));
 sg13g2_nand2_1 _0732_ (.Y(_0236_),
    .A(net134),
    .B(net125));
 sg13g2_o21ai_1 _0733_ (.B1(_0236_),
    .Y(_0007_),
    .A1(_0165_),
    .A2(_0235_));
 sg13g2_nand2_1 _0734_ (.Y(_0237_),
    .A(net133),
    .B(net125));
 sg13g2_o21ai_1 _0735_ (.B1(_0237_),
    .Y(_0008_),
    .A1(_0173_),
    .A2(_0235_));
 sg13g2_nand2_1 _0736_ (.Y(_0238_),
    .A(net132),
    .B(net125));
 sg13g2_o21ai_1 _0737_ (.B1(_0238_),
    .Y(_0009_),
    .A1(_0181_),
    .A2(_0235_));
 sg13g2_nand2_1 _0738_ (.Y(_0239_),
    .A(net139),
    .B(_0233_));
 sg13g2_o21ai_1 _0739_ (.B1(_0239_),
    .Y(_0010_),
    .A1(_0124_),
    .A2(_0235_));
 sg13g2_nand2_1 _0740_ (.Y(_0240_),
    .A(net138),
    .B(_0233_));
 sg13g2_o21ai_1 _0741_ (.B1(_0240_),
    .Y(_0011_),
    .A1(_0132_),
    .A2(_0235_));
 sg13g2_nand2_1 _0742_ (.Y(_0241_),
    .A(net137),
    .B(net125));
 sg13g2_o21ai_1 _0743_ (.B1(_0241_),
    .Y(_0012_),
    .A1(_0140_),
    .A2(_0235_));
 sg13g2_nand2_1 _0744_ (.Y(_0242_),
    .A(net136),
    .B(net125));
 sg13g2_o21ai_1 _0745_ (.B1(_0242_),
    .Y(_0013_),
    .A1(_0148_),
    .A2(_0235_));
 sg13g2_nand2_1 _0746_ (.Y(_0243_),
    .A(_0112_),
    .B(net141));
 sg13g2_nor2_1 _0747_ (.A(net310),
    .B(_0243_),
    .Y(_0244_));
 sg13g2_and4_1 _0748_ (.A(net156),
    .B(_0214_),
    .C(_0223_),
    .D(_0244_),
    .X(_0245_));
 sg13g2_nand2_1 _0749_ (.Y(_0246_),
    .A(net216),
    .B(net124));
 sg13g2_nand2b_2 _0750_ (.Y(_0247_),
    .B(net155),
    .A_N(_0245_));
 sg13g2_o21ai_1 _0751_ (.B1(_0246_),
    .Y(_0014_),
    .A1(_0156_),
    .A2(_0247_));
 sg13g2_nand2_1 _0752_ (.Y(_0248_),
    .A(\tb.val_saved[1] ),
    .B(net124));
 sg13g2_o21ai_1 _0753_ (.B1(_0248_),
    .Y(_0015_),
    .A1(_0164_),
    .A2(_0247_));
 sg13g2_nand2_1 _0754_ (.Y(_0249_),
    .A(net168),
    .B(net124));
 sg13g2_o21ai_1 _0755_ (.B1(_0249_),
    .Y(_0016_),
    .A1(_0172_),
    .A2(_0247_));
 sg13g2_nand2_1 _0756_ (.Y(_0250_),
    .A(net132),
    .B(net124));
 sg13g2_o21ai_1 _0757_ (.B1(_0250_),
    .Y(_0017_),
    .A1(_0180_),
    .A2(_0247_));
 sg13g2_nand2_1 _0758_ (.Y(_0251_),
    .A(\tb.key_saved[0] ),
    .B(net124));
 sg13g2_o21ai_1 _0759_ (.B1(_0251_),
    .Y(_0018_),
    .A1(_0123_),
    .A2(_0247_));
 sg13g2_nand2_1 _0760_ (.Y(_0252_),
    .A(\tb.key_saved[1] ),
    .B(net124));
 sg13g2_o21ai_1 _0761_ (.B1(_0252_),
    .Y(_0019_),
    .A1(_0131_),
    .A2(_0247_));
 sg13g2_nand2_1 _0762_ (.Y(_0253_),
    .A(\tb.key_saved[2] ),
    .B(net124));
 sg13g2_o21ai_1 _0763_ (.B1(_0253_),
    .Y(_0020_),
    .A1(_0139_),
    .A2(_0247_));
 sg13g2_nand2_1 _0764_ (.Y(_0254_),
    .A(\tb.key_saved[3] ),
    .B(net124));
 sg13g2_o21ai_1 _0765_ (.B1(_0254_),
    .Y(_0021_),
    .A1(_0147_),
    .A2(_0247_));
 sg13g2_nor2_1 _0766_ (.A(\tb.cursor[0] ),
    .B(_0243_),
    .Y(_0255_));
 sg13g2_and4_2 _0767_ (.A(net156),
    .B(_0214_),
    .C(_0223_),
    .D(_0255_),
    .X(_0256_));
 sg13g2_nand2_1 _0768_ (.Y(_0257_),
    .A(net135),
    .B(net123));
 sg13g2_nand2b_2 _0769_ (.Y(_0258_),
    .B(net155),
    .A_N(net123));
 sg13g2_o21ai_1 _0770_ (.B1(_0257_),
    .Y(_0022_),
    .A1(_0155_),
    .A2(_0258_));
 sg13g2_nand2_1 _0771_ (.Y(_0259_),
    .A(net134),
    .B(_0256_));
 sg13g2_o21ai_1 _0772_ (.B1(_0259_),
    .Y(_0023_),
    .A1(_0163_),
    .A2(_0258_));
 sg13g2_nand2_1 _0773_ (.Y(_0260_),
    .A(net133),
    .B(net123));
 sg13g2_o21ai_1 _0774_ (.B1(_0260_),
    .Y(_0024_),
    .A1(_0171_),
    .A2(_0258_));
 sg13g2_nand2_1 _0775_ (.Y(_0261_),
    .A(net132),
    .B(net123));
 sg13g2_o21ai_1 _0776_ (.B1(_0261_),
    .Y(_0025_),
    .A1(_0179_),
    .A2(_0258_));
 sg13g2_nand2_1 _0777_ (.Y(_0262_),
    .A(\tb.key_saved[0] ),
    .B(_0256_));
 sg13g2_o21ai_1 _0778_ (.B1(_0262_),
    .Y(_0026_),
    .A1(_0122_),
    .A2(_0258_));
 sg13g2_nand2_1 _0779_ (.Y(_0263_),
    .A(\tb.key_saved[1] ),
    .B(net123));
 sg13g2_o21ai_1 _0780_ (.B1(_0263_),
    .Y(_0027_),
    .A1(_0130_),
    .A2(_0258_));
 sg13g2_nand2_1 _0781_ (.Y(_0264_),
    .A(net137),
    .B(net123));
 sg13g2_o21ai_1 _0782_ (.B1(_0264_),
    .Y(_0028_),
    .A1(_0138_),
    .A2(_0258_));
 sg13g2_nand2_1 _0783_ (.Y(_0265_),
    .A(net136),
    .B(net123));
 sg13g2_o21ai_1 _0784_ (.B1(_0265_),
    .Y(_0029_),
    .A1(_0146_),
    .A2(_0258_));
 sg13g2_nor3_1 _0785_ (.A(_0112_),
    .B(_0113_),
    .C(net310),
    .Y(_0266_));
 sg13g2_and4_1 _0786_ (.A(net153),
    .B(net127),
    .C(_0223_),
    .D(_0266_),
    .X(_0267_));
 sg13g2_nand2_1 _0787_ (.Y(_0268_),
    .A(net135),
    .B(_0267_));
 sg13g2_nand2b_2 _0788_ (.Y(_0269_),
    .B(net151),
    .A_N(_0267_));
 sg13g2_o21ai_1 _0789_ (.B1(_0268_),
    .Y(_0030_),
    .A1(_0160_),
    .A2(_0269_));
 sg13g2_nand2_1 _0790_ (.Y(_0270_),
    .A(net134),
    .B(net122));
 sg13g2_o21ai_1 _0791_ (.B1(_0270_),
    .Y(_0031_),
    .A1(_0168_),
    .A2(_0269_));
 sg13g2_nand2_1 _0792_ (.Y(_0271_),
    .A(net133),
    .B(net122));
 sg13g2_o21ai_1 _0793_ (.B1(_0271_),
    .Y(_0032_),
    .A1(_0176_),
    .A2(_0269_));
 sg13g2_nand2_1 _0794_ (.Y(_0272_),
    .A(net132),
    .B(net122));
 sg13g2_o21ai_1 _0795_ (.B1(_0272_),
    .Y(_0033_),
    .A1(_0184_),
    .A2(_0269_));
 sg13g2_nand2_1 _0796_ (.Y(_0273_),
    .A(net139),
    .B(net122));
 sg13g2_o21ai_1 _0797_ (.B1(_0273_),
    .Y(_0034_),
    .A1(_0127_),
    .A2(_0269_));
 sg13g2_nand2_1 _0798_ (.Y(_0274_),
    .A(net138),
    .B(net122));
 sg13g2_o21ai_1 _0799_ (.B1(_0274_),
    .Y(_0035_),
    .A1(_0135_),
    .A2(_0269_));
 sg13g2_nand2_1 _0800_ (.Y(_0275_),
    .A(net137),
    .B(net122));
 sg13g2_o21ai_1 _0801_ (.B1(_0275_),
    .Y(_0036_),
    .A1(_0143_),
    .A2(_0269_));
 sg13g2_nand2_1 _0802_ (.Y(_0276_),
    .A(net136),
    .B(net122));
 sg13g2_o21ai_1 _0803_ (.B1(_0276_),
    .Y(_0037_),
    .A1(_0151_),
    .A2(_0269_));
 sg13g2_nand2_1 _0804_ (.Y(_0277_),
    .A(net135),
    .B(net126));
 sg13g2_nand2b_2 _0805_ (.Y(_0278_),
    .B(net151),
    .A_N(_0226_));
 sg13g2_o21ai_1 _0806_ (.B1(_0277_),
    .Y(_0038_),
    .A1(_0159_),
    .A2(_0278_));
 sg13g2_nand2_1 _0807_ (.Y(_0279_),
    .A(net134),
    .B(net126));
 sg13g2_o21ai_1 _0808_ (.B1(_0279_),
    .Y(_0039_),
    .A1(_0167_),
    .A2(_0278_));
 sg13g2_nand2_1 _0809_ (.Y(_0280_),
    .A(net133),
    .B(net126));
 sg13g2_o21ai_1 _0810_ (.B1(_0280_),
    .Y(_0040_),
    .A1(_0175_),
    .A2(_0278_));
 sg13g2_nand2_1 _0811_ (.Y(_0281_),
    .A(net132),
    .B(net126));
 sg13g2_o21ai_1 _0812_ (.B1(_0281_),
    .Y(_0041_),
    .A1(_0183_),
    .A2(_0278_));
 sg13g2_nand2_1 _0813_ (.Y(_0282_),
    .A(net139),
    .B(_0226_));
 sg13g2_o21ai_1 _0814_ (.B1(_0282_),
    .Y(_0042_),
    .A1(_0126_),
    .A2(_0278_));
 sg13g2_nand2_1 _0815_ (.Y(_0283_),
    .A(net138),
    .B(net126));
 sg13g2_o21ai_1 _0816_ (.B1(_0283_),
    .Y(_0043_),
    .A1(_0134_),
    .A2(_0278_));
 sg13g2_nand2_1 _0817_ (.Y(_0284_),
    .A(net137),
    .B(net126));
 sg13g2_o21ai_1 _0818_ (.B1(_0284_),
    .Y(_0044_),
    .A1(_0142_),
    .A2(_0278_));
 sg13g2_nand2_1 _0819_ (.Y(_0285_),
    .A(net136),
    .B(net126));
 sg13g2_o21ai_1 _0820_ (.B1(_0285_),
    .Y(_0045_),
    .A1(_0150_),
    .A2(_0278_));
 sg13g2_nor3_1 _0821_ (.A(\tb.cursor[2] ),
    .B(net141),
    .C(net310),
    .Y(_0286_));
 sg13g2_and4_1 _0822_ (.A(net153),
    .B(net127),
    .C(_0223_),
    .D(_0286_),
    .X(_0287_));
 sg13g2_nand2_1 _0823_ (.Y(_0288_),
    .A(net299),
    .B(net153));
 sg13g2_a21oi_1 _0824_ (.A1(_0228_),
    .A2(_0286_),
    .Y(_0289_),
    .B1(_0288_));
 sg13g2_or2_1 _0825_ (.X(_0046_),
    .B(_0289_),
    .A(net121));
 sg13g2_nor2_1 _0826_ (.A(_0118_),
    .B(_0221_),
    .Y(_0290_));
 sg13g2_a21oi_1 _0827_ (.A1(net290),
    .A2(net11),
    .Y(_0291_),
    .B1(net142));
 sg13g2_a21o_1 _0828_ (.A2(net11),
    .A1(\tb.go_ok ),
    .B1(net142),
    .X(_0292_));
 sg13g2_o21ai_1 _0829_ (.B1(_0292_),
    .Y(_0293_),
    .A1(_0004_),
    .A2(_0222_));
 sg13g2_a221oi_1 _0830_ (.B2(_0290_),
    .C1(_0293_),
    .B1(_0227_),
    .A1(net127),
    .Y(_0294_),
    .A2(_0223_));
 sg13g2_nand2_1 _0831_ (.Y(_0295_),
    .A(net8),
    .B(net6));
 sg13g2_o21ai_1 _0832_ (.B1(_0109_),
    .Y(_0296_),
    .A1(_0107_),
    .A2(_0110_));
 sg13g2_o21ai_1 _0833_ (.B1(_0296_),
    .Y(_0297_),
    .A1(_0110_),
    .A2(_0295_));
 sg13g2_nor2_1 _0834_ (.A(net303),
    .B(_0297_),
    .Y(_0298_));
 sg13g2_a21oi_1 _0835_ (.A1(net305),
    .A2(net142),
    .Y(_0299_),
    .B1(_0298_));
 sg13g2_o21ai_1 _0836_ (.B1(net156),
    .Y(_0300_),
    .A1(net307),
    .A2(net120));
 sg13g2_a21oi_1 _0837_ (.A1(net120),
    .A2(_0299_),
    .Y(_0047_),
    .B1(_0300_));
 sg13g2_and2_1 _0838_ (.A(net141),
    .B(\tb.cursor[0] ),
    .X(_0301_));
 sg13g2_xnor2_1 _0839_ (.Y(_0302_),
    .A(_0108_),
    .B(_0295_));
 sg13g2_or3_1 _0840_ (.A(_0118_),
    .B(_0231_),
    .C(_0301_),
    .X(_0303_));
 sg13g2_o21ai_1 _0841_ (.B1(_0303_),
    .Y(_0304_),
    .A1(net142),
    .A2(_0302_));
 sg13g2_nor2b_1 _0842_ (.A(_0304_),
    .B_N(net120),
    .Y(_0305_));
 sg13g2_o21ai_1 _0843_ (.B1(net152),
    .Y(_0306_),
    .A1(net141),
    .A2(net120));
 sg13g2_nor2_1 _0844_ (.A(_0305_),
    .B(_0306_),
    .Y(_0048_));
 sg13g2_nor2_1 _0845_ (.A(_0107_),
    .B(net7),
    .Y(_0307_));
 sg13g2_nand2_1 _0846_ (.Y(_0308_),
    .A(net140),
    .B(_0301_));
 sg13g2_xnor2_1 _0847_ (.Y(_0309_),
    .A(net140),
    .B(_0301_));
 sg13g2_nand2_1 _0848_ (.Y(_0310_),
    .A(net142),
    .B(_0309_));
 sg13g2_o21ai_1 _0849_ (.B1(_0310_),
    .Y(_0311_),
    .A1(net142),
    .A2(_0307_));
 sg13g2_o21ai_1 _0850_ (.B1(net153),
    .Y(_0312_),
    .A1(net140),
    .A2(_0294_));
 sg13g2_a21oi_1 _0851_ (.A1(net120),
    .A2(_0311_),
    .Y(_0049_),
    .B1(_0312_));
 sg13g2_nor3_1 _0852_ (.A(_0112_),
    .B(\tb.cursor[1] ),
    .C(_0003_),
    .Y(_0313_));
 sg13g2_and4_1 _0853_ (.A(net151),
    .B(net127),
    .C(_0223_),
    .D(_0313_),
    .X(_0314_));
 sg13g2_nand2_1 _0854_ (.Y(_0315_),
    .A(net135),
    .B(_0314_));
 sg13g2_nand2b_2 _0855_ (.Y(_0316_),
    .B(net151),
    .A_N(_0314_));
 sg13g2_o21ai_1 _0856_ (.B1(_0315_),
    .Y(_0050_),
    .A1(_0158_),
    .A2(_0316_));
 sg13g2_nand2_1 _0857_ (.Y(_0317_),
    .A(net134),
    .B(net119));
 sg13g2_o21ai_1 _0858_ (.B1(_0317_),
    .Y(_0051_),
    .A1(_0166_),
    .A2(_0316_));
 sg13g2_nand2_1 _0859_ (.Y(_0318_),
    .A(net133),
    .B(net119));
 sg13g2_o21ai_1 _0860_ (.B1(_0318_),
    .Y(_0052_),
    .A1(_0174_),
    .A2(_0316_));
 sg13g2_nand2_1 _0861_ (.Y(_0319_),
    .A(net132),
    .B(net119));
 sg13g2_o21ai_1 _0862_ (.B1(_0319_),
    .Y(_0053_),
    .A1(_0182_),
    .A2(_0316_));
 sg13g2_nand2_1 _0863_ (.Y(_0320_),
    .A(net139),
    .B(net119));
 sg13g2_o21ai_1 _0864_ (.B1(_0320_),
    .Y(_0054_),
    .A1(_0125_),
    .A2(_0316_));
 sg13g2_nand2_1 _0865_ (.Y(_0321_),
    .A(net138),
    .B(net119));
 sg13g2_o21ai_1 _0866_ (.B1(_0321_),
    .Y(_0055_),
    .A1(_0133_),
    .A2(_0316_));
 sg13g2_nand2_1 _0867_ (.Y(_0322_),
    .A(net137),
    .B(net119));
 sg13g2_o21ai_1 _0868_ (.B1(_0322_),
    .Y(_0056_),
    .A1(_0141_),
    .A2(_0316_));
 sg13g2_nand2_1 _0869_ (.Y(_0323_),
    .A(net136),
    .B(net119));
 sg13g2_o21ai_1 _0870_ (.B1(_0323_),
    .Y(_0057_),
    .A1(_0149_),
    .A2(_0316_));
 sg13g2_nand2_1 _0871_ (.Y(_0324_),
    .A(net135),
    .B(net121));
 sg13g2_nand2b_2 _0872_ (.Y(_0325_),
    .B(net155),
    .A_N(_0287_));
 sg13g2_o21ai_1 _0873_ (.B1(_0324_),
    .Y(_0058_),
    .A1(_0154_),
    .A2(_0325_));
 sg13g2_nand2_1 _0874_ (.Y(_0326_),
    .A(net134),
    .B(_0287_));
 sg13g2_o21ai_1 _0875_ (.B1(_0326_),
    .Y(_0059_),
    .A1(_0162_),
    .A2(_0325_));
 sg13g2_nand2_1 _0876_ (.Y(_0327_),
    .A(net133),
    .B(net121));
 sg13g2_o21ai_1 _0877_ (.B1(_0327_),
    .Y(_0060_),
    .A1(_0170_),
    .A2(_0325_));
 sg13g2_nand2_1 _0878_ (.Y(_0328_),
    .A(net132),
    .B(net121));
 sg13g2_o21ai_1 _0879_ (.B1(_0328_),
    .Y(_0061_),
    .A1(_0178_),
    .A2(_0325_));
 sg13g2_nand2_1 _0880_ (.Y(_0329_),
    .A(net139),
    .B(net121));
 sg13g2_o21ai_1 _0881_ (.B1(_0329_),
    .Y(_0062_),
    .A1(_0121_),
    .A2(_0325_));
 sg13g2_nand2_1 _0882_ (.Y(_0330_),
    .A(net138),
    .B(net121));
 sg13g2_o21ai_1 _0883_ (.B1(_0330_),
    .Y(_0063_),
    .A1(_0129_),
    .A2(_0325_));
 sg13g2_nand2_1 _0884_ (.Y(_0331_),
    .A(net137),
    .B(net121));
 sg13g2_o21ai_1 _0885_ (.B1(_0331_),
    .Y(_0064_),
    .A1(_0137_),
    .A2(_0325_));
 sg13g2_nand2_1 _0886_ (.Y(_0332_),
    .A(net136),
    .B(net121));
 sg13g2_o21ai_1 _0887_ (.B1(_0332_),
    .Y(_0065_),
    .A1(_0145_),
    .A2(_0325_));
 sg13g2_nand3_1 _0888_ (.B(_0228_),
    .C(_0231_),
    .A(net140),
    .Y(_0333_));
 sg13g2_and2_1 _0889_ (.A(net301),
    .B(net151),
    .X(_0334_));
 sg13g2_a21o_1 _0890_ (.A2(_0334_),
    .A1(_0333_),
    .B1(net125),
    .X(_0066_));
 sg13g2_nor3_1 _0891_ (.A(\tb.cursor[2] ),
    .B(net141),
    .C(\tb.cursor[0] ),
    .Y(_0335_));
 sg13g2_and4_1 _0892_ (.A(net153),
    .B(net127),
    .C(_0223_),
    .D(_0335_),
    .X(_0336_));
 sg13g2_nand2_1 _0893_ (.Y(_0337_),
    .A(net293),
    .B(net153));
 sg13g2_a21oi_1 _0894_ (.A1(_0228_),
    .A2(_0335_),
    .Y(_0338_),
    .B1(_0337_));
 sg13g2_or2_1 _0895_ (.X(_0067_),
    .B(_0338_),
    .A(net118));
 sg13g2_nor3_1 _0896_ (.A(net127),
    .B(_0221_),
    .C(_0227_),
    .Y(_0339_));
 sg13g2_o21ai_1 _0897_ (.B1(net152),
    .Y(_0340_),
    .A1(_0118_),
    .A2(_0339_));
 sg13g2_nor2_1 _0898_ (.A(_0291_),
    .B(_0340_),
    .Y(_0068_));
 sg13g2_nand2_1 _0899_ (.Y(_0341_),
    .A(net296),
    .B(net156));
 sg13g2_a21oi_1 _0900_ (.A1(_0228_),
    .A2(_0255_),
    .Y(_0342_),
    .B1(_0341_));
 sg13g2_or2_1 _0901_ (.X(_0069_),
    .B(_0342_),
    .A(net123));
 sg13g2_nand2_1 _0902_ (.Y(_0343_),
    .A(net297),
    .B(net151));
 sg13g2_a21oi_1 _0903_ (.A1(_0228_),
    .A2(_0313_),
    .Y(_0344_),
    .B1(_0343_));
 sg13g2_or2_1 _0904_ (.X(_0070_),
    .B(net298),
    .A(net119));
 sg13g2_nand2_1 _0905_ (.Y(_0345_),
    .A(net295),
    .B(net156));
 sg13g2_a21oi_1 _0906_ (.A1(_0228_),
    .A2(_0244_),
    .Y(_0346_),
    .B1(_0345_));
 sg13g2_or2_1 _0907_ (.X(_0071_),
    .B(_0346_),
    .A(_0245_));
 sg13g2_nor3_1 _0908_ (.A(net127),
    .B(_0224_),
    .C(_0227_),
    .Y(_0347_));
 sg13g2_o21ai_1 _0909_ (.B1(net279),
    .Y(_0348_),
    .A1(_0291_),
    .A2(_0347_));
 sg13g2_nand2b_1 _0910_ (.Y(_0349_),
    .B(_0185_),
    .A_N(_0004_));
 sg13g2_nand3_1 _0911_ (.B(_0292_),
    .C(_0349_),
    .A(_0224_),
    .Y(_0350_));
 sg13g2_a21oi_1 _0912_ (.A1(_0348_),
    .A2(_0350_),
    .Y(_0072_),
    .B1(_0152_));
 sg13g2_o21ai_1 _0913_ (.B1(_0292_),
    .Y(_0351_),
    .A1(_0004_),
    .A2(_0185_));
 sg13g2_nand2b_1 _0914_ (.Y(_0352_),
    .B(_0224_),
    .A_N(_0351_));
 sg13g2_o21ai_1 _0915_ (.B1(net281),
    .Y(_0353_),
    .A1(_0291_),
    .A2(_0347_));
 sg13g2_a21oi_1 _0916_ (.A1(_0352_),
    .A2(_0353_),
    .Y(_0073_),
    .B1(_0152_));
 sg13g2_o21ai_1 _0917_ (.B1(_0290_),
    .Y(_0354_),
    .A1(net127),
    .A2(_0227_));
 sg13g2_mux4_1 _0918_ (.S0(net149),
    .A0(_0153_),
    .A1(_0154_),
    .A2(_0155_),
    .A3(_0156_),
    .S1(net146),
    .X(_0355_));
 sg13g2_mux4_1 _0919_ (.S0(net148),
    .A0(\tb.mem[4][0] ),
    .A1(\tb.mem[5][0] ),
    .A2(\tb.mem[6][0] ),
    .A3(\tb.mem[7][0] ),
    .S1(net145),
    .X(_0356_));
 sg13g2_nand2_1 _0920_ (.Y(_0357_),
    .A(net143),
    .B(_0356_));
 sg13g2_o21ai_1 _0921_ (.B1(_0357_),
    .Y(_0358_),
    .A1(net143),
    .A2(_0355_));
 sg13g2_o21ai_1 _0922_ (.B1(net152),
    .Y(_0359_),
    .A1(_0354_),
    .A2(_0358_));
 sg13g2_a21oi_1 _0923_ (.A1(_0117_),
    .A2(_0354_),
    .Y(_0074_),
    .B1(_0359_));
 sg13g2_mux4_1 _0924_ (.S0(net149),
    .A0(_0161_),
    .A1(_0162_),
    .A2(_0163_),
    .A3(_0164_),
    .S1(net146),
    .X(_0360_));
 sg13g2_mux4_1 _0925_ (.S0(net148),
    .A0(\tb.mem[4][1] ),
    .A1(\tb.mem[5][1] ),
    .A2(\tb.mem[6][1] ),
    .A3(\tb.mem[7][1] ),
    .S1(net145),
    .X(_0361_));
 sg13g2_nand2_1 _0926_ (.Y(_0362_),
    .A(net143),
    .B(_0361_));
 sg13g2_o21ai_1 _0927_ (.B1(_0362_),
    .Y(_0363_),
    .A1(net143),
    .A2(_0360_));
 sg13g2_o21ai_1 _0928_ (.B1(net152),
    .Y(_0364_),
    .A1(_0354_),
    .A2(_0363_));
 sg13g2_a21oi_1 _0929_ (.A1(_0116_),
    .A2(_0354_),
    .Y(_0075_),
    .B1(_0364_));
 sg13g2_mux4_1 _0930_ (.S0(net149),
    .A0(_0169_),
    .A1(_0170_),
    .A2(_0171_),
    .A3(_0172_),
    .S1(net146),
    .X(_0365_));
 sg13g2_mux4_1 _0931_ (.S0(net148),
    .A0(\tb.mem[4][2] ),
    .A1(\tb.mem[5][2] ),
    .A2(\tb.mem[6][2] ),
    .A3(\tb.mem[7][2] ),
    .S1(net145),
    .X(_0366_));
 sg13g2_nand2_1 _0932_ (.Y(_0367_),
    .A(net144),
    .B(_0366_));
 sg13g2_o21ai_1 _0933_ (.B1(_0367_),
    .Y(_0368_),
    .A1(net144),
    .A2(_0365_));
 sg13g2_o21ai_1 _0934_ (.B1(net152),
    .Y(_0369_),
    .A1(_0354_),
    .A2(_0368_));
 sg13g2_a21oi_1 _0935_ (.A1(_0115_),
    .A2(_0354_),
    .Y(_0076_),
    .B1(_0369_));
 sg13g2_mux4_1 _0936_ (.S0(net149),
    .A0(_0177_),
    .A1(_0178_),
    .A2(_0179_),
    .A3(_0180_),
    .S1(net146),
    .X(_0370_));
 sg13g2_mux4_1 _0937_ (.S0(net148),
    .A0(\tb.mem[4][3] ),
    .A1(\tb.mem[5][3] ),
    .A2(\tb.mem[6][3] ),
    .A3(\tb.mem[7][3] ),
    .S1(net145),
    .X(_0371_));
 sg13g2_nand2_1 _0938_ (.Y(_0372_),
    .A(net144),
    .B(_0371_));
 sg13g2_o21ai_1 _0939_ (.B1(_0372_),
    .Y(_0373_),
    .A1(net144),
    .A2(_0370_));
 sg13g2_o21ai_1 _0940_ (.B1(net152),
    .Y(_0374_),
    .A1(_0354_),
    .A2(_0373_));
 sg13g2_a21oi_1 _0941_ (.A1(_0114_),
    .A2(_0354_),
    .Y(_0077_),
    .B1(_0374_));
 sg13g2_nand3_1 _0942_ (.B(net120),
    .C(_0301_),
    .A(net140),
    .Y(_0375_));
 sg13g2_o21ai_1 _0943_ (.B1(net142),
    .Y(_0376_),
    .A1(_0111_),
    .A2(_0308_));
 sg13g2_a221oi_1 _0944_ (.B2(net120),
    .C1(_0152_),
    .B1(_0376_),
    .A1(_0111_),
    .Y(_0081_),
    .A2(_0375_));
 sg13g2_nand2b_1 _0945_ (.Y(_0377_),
    .B(_0004_),
    .A_N(net11));
 sg13g2_nand2b_1 _0946_ (.Y(_0378_),
    .B(net290),
    .A_N(_0004_));
 sg13g2_nand3_1 _0947_ (.B(_0377_),
    .C(net291),
    .A(net154),
    .Y(_0082_));
 sg13g2_and3_1 _0948_ (.X(_0379_),
    .A(\tb.go_ok ),
    .B(net11),
    .C(_0004_));
 sg13g2_o21ai_1 _0949_ (.B1(net157),
    .Y(_0380_),
    .A1(net139),
    .A2(net129));
 sg13g2_a21oi_1 _0950_ (.A1(_0110_),
    .A2(net129),
    .Y(_0083_),
    .B1(_0380_));
 sg13g2_o21ai_1 _0951_ (.B1(net155),
    .Y(_0381_),
    .A1(net138),
    .A2(net129));
 sg13g2_a21oi_1 _0952_ (.A1(_0109_),
    .A2(net129),
    .Y(_0084_),
    .B1(_0381_));
 sg13g2_o21ai_1 _0953_ (.B1(net156),
    .Y(_0382_),
    .A1(net137),
    .A2(net131));
 sg13g2_a21oi_1 _0954_ (.A1(_0108_),
    .A2(net131),
    .Y(_0085_),
    .B1(_0382_));
 sg13g2_o21ai_1 _0955_ (.B1(net156),
    .Y(_0383_),
    .A1(net136),
    .A2(net128));
 sg13g2_a21oi_1 _0956_ (.A1(_0107_),
    .A2(net128),
    .Y(_0086_),
    .B1(_0383_));
 sg13g2_o21ai_1 _0957_ (.B1(net157),
    .Y(_0384_),
    .A1(net135),
    .A2(net130));
 sg13g2_a21oi_1 _0958_ (.A1(_0106_),
    .A2(net130),
    .Y(_0087_),
    .B1(_0384_));
 sg13g2_o21ai_1 _0959_ (.B1(net155),
    .Y(_0385_),
    .A1(net134),
    .A2(net130));
 sg13g2_a21oi_1 _0960_ (.A1(_0105_),
    .A2(net130),
    .Y(_0088_),
    .B1(_0385_));
 sg13g2_o21ai_1 _0961_ (.B1(net155),
    .Y(_0386_),
    .A1(net133),
    .A2(net129));
 sg13g2_a21oi_1 _0962_ (.A1(_0104_),
    .A2(net129),
    .Y(_0089_),
    .B1(_0386_));
 sg13g2_o21ai_1 _0963_ (.B1(net155),
    .Y(_0387_),
    .A1(net132),
    .A2(net129));
 sg13g2_a21oi_1 _0964_ (.A1(_0103_),
    .A2(net129),
    .Y(_0090_),
    .B1(_0387_));
 sg13g2_o21ai_1 _0965_ (.B1(net156),
    .Y(_0388_),
    .A1(net288),
    .A2(net128));
 sg13g2_a21oi_1 _0966_ (.A1(_0297_),
    .A2(net128),
    .Y(_0091_),
    .B1(_0388_));
 sg13g2_o21ai_1 _0967_ (.B1(net153),
    .Y(_0389_),
    .A1(net289),
    .A2(net128));
 sg13g2_a21oi_1 _0968_ (.A1(_0302_),
    .A2(net128),
    .Y(_0092_),
    .B1(_0389_));
 sg13g2_o21ai_1 _0969_ (.B1(net128),
    .Y(_0390_),
    .A1(_0107_),
    .A2(net7));
 sg13g2_o21ai_1 _0970_ (.B1(_0390_),
    .Y(_0391_),
    .A1(net300),
    .A2(net128));
 sg13g2_nor2_1 _0971_ (.A(_0152_),
    .B(_0391_),
    .Y(_0093_));
 sg13g2_nand2_1 _0972_ (.Y(_0392_),
    .A(net135),
    .B(net118));
 sg13g2_nand2b_2 _0973_ (.Y(_0393_),
    .B(net155),
    .A_N(_0336_));
 sg13g2_o21ai_1 _0974_ (.B1(_0392_),
    .Y(_0094_),
    .A1(_0153_),
    .A2(_0393_));
 sg13g2_nand2_1 _0975_ (.Y(_0394_),
    .A(net134),
    .B(net118));
 sg13g2_o21ai_1 _0976_ (.B1(_0394_),
    .Y(_0095_),
    .A1(_0161_),
    .A2(_0393_));
 sg13g2_nand2_1 _0977_ (.Y(_0395_),
    .A(net133),
    .B(net118));
 sg13g2_o21ai_1 _0978_ (.B1(_0395_),
    .Y(_0096_),
    .A1(_0169_),
    .A2(_0393_));
 sg13g2_nand2_1 _0979_ (.Y(_0396_),
    .A(net170),
    .B(_0336_));
 sg13g2_o21ai_1 _0980_ (.B1(_0396_),
    .Y(_0097_),
    .A1(_0177_),
    .A2(_0393_));
 sg13g2_nand2_1 _0981_ (.Y(_0397_),
    .A(net139),
    .B(net118));
 sg13g2_o21ai_1 _0982_ (.B1(_0397_),
    .Y(_0098_),
    .A1(_0120_),
    .A2(_0393_));
 sg13g2_nand2_1 _0983_ (.Y(_0398_),
    .A(net138),
    .B(net118));
 sg13g2_o21ai_1 _0984_ (.B1(_0398_),
    .Y(_0099_),
    .A1(_0128_),
    .A2(_0393_));
 sg13g2_nand2_1 _0985_ (.Y(_0399_),
    .A(net137),
    .B(net118));
 sg13g2_o21ai_1 _0986_ (.B1(_0399_),
    .Y(_0100_),
    .A1(_0136_),
    .A2(_0393_));
 sg13g2_nand2_1 _0987_ (.Y(_0400_),
    .A(net136),
    .B(net118));
 sg13g2_o21ai_1 _0988_ (.B1(_0400_),
    .Y(_0101_),
    .A1(_0144_),
    .A2(_0393_));
 sg13g2_nand2_1 _0989_ (.Y(_0401_),
    .A(net294),
    .B(net153));
 sg13g2_a21oi_1 _0990_ (.A1(_0228_),
    .A2(_0266_),
    .Y(_0402_),
    .B1(_0401_));
 sg13g2_or2_1 _0991_ (.X(_0102_),
    .B(_0402_),
    .A(net122));
 sg13g2_a21oi_1 _0992_ (.A1(net120),
    .A2(_0299_),
    .Y(_0078_),
    .B1(_0300_));
 sg13g2_nor2_1 _0993_ (.A(_0305_),
    .B(_0306_),
    .Y(_0079_));
 sg13g2_a21oi_1 _0994_ (.A1(_0294_),
    .A2(_0311_),
    .Y(_0080_),
    .B1(_0312_));
 sg13g2_dfrbp_1 _0995_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net73),
    .D(_0005_),
    .Q_N(_0498_),
    .Q(\tb.mem[6][8] ));
 sg13g2_dfrbp_1 _0996_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net34),
    .D(net205),
    .Q_N(_0497_),
    .Q(\tb.mem[4][0] ));
 sg13g2_dfrbp_1 _0997_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net32),
    .D(net270),
    .Q_N(_0496_),
    .Q(\tb.mem[4][1] ));
 sg13g2_dfrbp_1 _0998_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net30),
    .D(_0008_),
    .Q_N(_0495_),
    .Q(\tb.mem[4][2] ));
 sg13g2_dfrbp_1 _0999_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net28),
    .D(_0009_),
    .Q_N(_0494_),
    .Q(\tb.mem[4][3] ));
 sg13g2_dfrbp_1 _1000_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net164),
    .D(net243),
    .Q_N(_0493_),
    .Q(\tb.mem[4][4] ));
 sg13g2_dfrbp_1 _1001_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net162),
    .D(net259),
    .Q_N(_0492_),
    .Q(\tb.mem[4][5] ));
 sg13g2_dfrbp_1 _1002_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net160),
    .D(net229),
    .Q_N(_0491_),
    .Q(\tb.mem[4][6] ));
 sg13g2_dfrbp_1 _1003_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net158),
    .D(net241),
    .Q_N(_0490_),
    .Q(\tb.mem[4][7] ));
 sg13g2_dfrbp_1 _1004_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net116),
    .D(net217),
    .Q_N(_0489_),
    .Q(\tb.mem[3][0] ));
 sg13g2_dfrbp_1 _1005_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net114),
    .D(net202),
    .Q_N(_0488_),
    .Q(\tb.mem[3][1] ));
 sg13g2_dfrbp_1 _1006_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net112),
    .D(net169),
    .Q_N(_0487_),
    .Q(\tb.mem[3][2] ));
 sg13g2_dfrbp_1 _1007_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net110),
    .D(_0017_),
    .Q_N(_0486_),
    .Q(\tb.mem[3][3] ));
 sg13g2_dfrbp_1 _1008_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net108),
    .D(net183),
    .Q_N(_0485_),
    .Q(\tb.mem[3][4] ));
 sg13g2_dfrbp_1 _1009_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net106),
    .D(net219),
    .Q_N(_0484_),
    .Q(\tb.mem[3][5] ));
 sg13g2_dfrbp_1 _1010_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net104),
    .D(net224),
    .Q_N(_0483_),
    .Q(\tb.mem[3][6] ));
 sg13g2_dfrbp_1 _1011_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net102),
    .D(net211),
    .Q_N(_0482_),
    .Q(\tb.mem[3][7] ));
 sg13g2_dfrbp_1 _1012_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net100),
    .D(net195),
    .Q_N(_0481_),
    .Q(\tb.mem[2][0] ));
 sg13g2_dfrbp_1 _1013_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net98),
    .D(net239),
    .Q_N(_0480_),
    .Q(\tb.mem[2][1] ));
 sg13g2_dfrbp_1 _1014_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net96),
    .D(_0024_),
    .Q_N(_0479_),
    .Q(\tb.mem[2][2] ));
 sg13g2_dfrbp_1 _1015_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net94),
    .D(_0025_),
    .Q_N(_0478_),
    .Q(\tb.mem[2][3] ));
 sg13g2_dfrbp_1 _1016_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net92),
    .D(net179),
    .Q_N(_0477_),
    .Q(\tb.mem[2][4] ));
 sg13g2_dfrbp_1 _1017_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net90),
    .D(net191),
    .Q_N(_0476_),
    .Q(\tb.mem[2][5] ));
 sg13g2_dfrbp_1 _1018_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net88),
    .D(net252),
    .Q_N(_0475_),
    .Q(\tb.mem[2][6] ));
 sg13g2_dfrbp_1 _1019_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net86),
    .D(net213),
    .Q_N(_0474_),
    .Q(\tb.mem[2][7] ));
 sg13g2_dfrbp_1 _1020_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net84),
    .D(_0030_),
    .Q_N(_0473_),
    .Q(\tb.mem[7][0] ));
 sg13g2_dfrbp_1 _1021_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net82),
    .D(net264),
    .Q_N(_0472_),
    .Q(\tb.mem[7][1] ));
 sg13g2_dfrbp_1 _1022_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net80),
    .D(_0032_),
    .Q_N(_0471_),
    .Q(\tb.mem[7][2] ));
 sg13g2_dfrbp_1 _1023_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net78),
    .D(_0033_),
    .Q_N(_0470_),
    .Q(\tb.mem[7][3] ));
 sg13g2_dfrbp_1 _1024_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net76),
    .D(net256),
    .Q_N(_0469_),
    .Q(\tb.mem[7][4] ));
 sg13g2_dfrbp_1 _1025_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net74),
    .D(net181),
    .Q_N(_0468_),
    .Q(\tb.mem[7][5] ));
 sg13g2_dfrbp_1 _1026_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net72),
    .D(net227),
    .Q_N(_0467_),
    .Q(\tb.mem[7][6] ));
 sg13g2_dfrbp_1 _1027_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net70),
    .D(net185),
    .Q_N(_0466_),
    .Q(\tb.mem[7][7] ));
 sg13g2_dfrbp_1 _1028_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net68),
    .D(_0038_),
    .Q_N(_0465_),
    .Q(\tb.mem[6][0] ));
 sg13g2_dfrbp_1 _1029_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net66),
    .D(net268),
    .Q_N(_0464_),
    .Q(\tb.mem[6][1] ));
 sg13g2_dfrbp_1 _1030_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net64),
    .D(_0040_),
    .Q_N(_0463_),
    .Q(\tb.mem[6][2] ));
 sg13g2_dfrbp_1 _1031_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net62),
    .D(_0041_),
    .Q_N(_0462_),
    .Q(\tb.mem[6][3] ));
 sg13g2_dfrbp_1 _1032_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net60),
    .D(net272),
    .Q_N(_0461_),
    .Q(\tb.mem[6][4] ));
 sg13g2_dfrbp_1 _1033_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net58),
    .D(net173),
    .Q_N(_0460_),
    .Q(\tb.mem[6][5] ));
 sg13g2_dfrbp_1 _1034_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net56),
    .D(net274),
    .Q_N(_0459_),
    .Q(\tb.mem[6][6] ));
 sg13g2_dfrbp_1 _1035_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net54),
    .D(net188),
    .Q_N(_0458_),
    .Q(\tb.mem[6][7] ));
 sg13g2_dfrbp_1 _1036_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net52),
    .D(_0046_),
    .Q_N(_0457_),
    .Q(\tb.mem[1][8] ));
 sg13g2_dfrbp_1 _1037_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net50),
    .D(_0047_),
    .Q_N(_0456_),
    .Q(_0000_));
 sg13g2_dfrbp_1 _1038_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net49),
    .D(_0048_),
    .Q_N(_0455_),
    .Q(_0001_));
 sg13g2_dfrbp_1 _1039_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net48),
    .D(_0049_),
    .Q_N(_0454_),
    .Q(_0002_));
 sg13g2_dfrbp_1 _1040_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net47),
    .D(net193),
    .Q_N(_0453_),
    .Q(\tb.mem[5][0] ));
 sg13g2_dfrbp_1 _1041_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net45),
    .D(net197),
    .Q_N(_0452_),
    .Q(\tb.mem[5][1] ));
 sg13g2_dfrbp_1 _1042_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net43),
    .D(_0052_),
    .Q_N(_0451_),
    .Q(\tb.mem[5][2] ));
 sg13g2_dfrbp_1 _1043_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net41),
    .D(_0053_),
    .Q_N(_0450_),
    .Q(\tb.mem[5][3] ));
 sg13g2_dfrbp_1 _1044_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net39),
    .D(net278),
    .Q_N(_0449_),
    .Q(\tb.mem[5][4] ));
 sg13g2_dfrbp_1 _1045_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net37),
    .D(net254),
    .Q_N(_0448_),
    .Q(\tb.mem[5][5] ));
 sg13g2_dfrbp_1 _1046_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net35),
    .D(net233),
    .Q_N(_0447_),
    .Q(\tb.mem[5][6] ));
 sg13g2_dfrbp_1 _1047_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net31),
    .D(net231),
    .Q_N(_0446_),
    .Q(\tb.mem[5][7] ));
 sg13g2_dfrbp_1 _1048_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net165),
    .D(_0058_),
    .Q_N(_0445_),
    .Q(\tb.mem[1][0] ));
 sg13g2_dfrbp_1 _1049_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net161),
    .D(net208),
    .Q_N(_0444_),
    .Q(\tb.mem[1][1] ));
 sg13g2_dfrbp_1 _1050_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net117),
    .D(_0060_),
    .Q_N(_0443_),
    .Q(\tb.mem[1][2] ));
 sg13g2_dfrbp_1 _1051_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net113),
    .D(_0061_),
    .Q_N(_0442_),
    .Q(\tb.mem[1][3] ));
 sg13g2_dfrbp_1 _1052_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net109),
    .D(net222),
    .Q_N(_0441_),
    .Q(\tb.mem[1][4] ));
 sg13g2_dfrbp_1 _1053_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net105),
    .D(net176),
    .Q_N(_0440_),
    .Q(\tb.mem[1][5] ));
 sg13g2_dfrbp_1 _1054_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net101),
    .D(net215),
    .Q_N(_0439_),
    .Q(\tb.mem[1][6] ));
 sg13g2_dfrbp_1 _1055_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net97),
    .D(net245),
    .Q_N(_0438_),
    .Q(\tb.mem[1][7] ));
 sg13g2_dfrbp_1 _1056_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net93),
    .D(net302),
    .Q_N(_0437_),
    .Q(\tb.mem[4][8] ));
 sg13g2_dfrbp_1 _1057_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net89),
    .D(_0067_),
    .Q_N(_0436_),
    .Q(\tb.mem[0][8] ));
 sg13g2_dfrbp_1 _1058_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net85),
    .D(_0068_),
    .Q_N(_0004_),
    .Q(\tb.state ));
 sg13g2_dfrbp_1 _1059_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net83),
    .D(_0069_),
    .Q_N(_0435_),
    .Q(\tb.mem[2][8] ));
 sg13g2_dfrbp_1 _1060_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net79),
    .D(_0070_),
    .Q_N(_0434_),
    .Q(\tb.mem[5][8] ));
 sg13g2_dfrbp_1 _1061_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net75),
    .D(_0071_),
    .Q_N(_0433_),
    .Q(\tb.mem[3][8] ));
 sg13g2_dfrbp_1 _1062_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net71),
    .D(net280),
    .Q_N(_0432_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _1063_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net67),
    .D(_0073_),
    .Q_N(_0431_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _1064_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net63),
    .D(_0074_),
    .Q_N(_0430_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _1065_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net59),
    .D(_0075_),
    .Q_N(_0429_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1066_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net55),
    .D(_0076_),
    .Q_N(_0428_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1067_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net51),
    .D(_0077_),
    .Q_N(_0427_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _1068_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net44),
    .D(net306),
    .Q_N(_0003_),
    .Q(\tb.cursor[0] ));
 sg13g2_dfrbp_1 _1069_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net40),
    .D(_0079_),
    .Q_N(_0426_),
    .Q(\tb.cursor[1] ));
 sg13g2_dfrbp_1 _1070_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net36),
    .D(_0080_),
    .Q_N(_0425_),
    .Q(\tb.cursor[2] ));
 sg13g2_dfrbp_1 _1071_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net29),
    .D(net283),
    .Q_N(_0424_),
    .Q(\tb.cursor[3] ));
 sg13g2_dfrbp_1 _1072_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net159),
    .D(net292),
    .Q_N(_0423_),
    .Q(\tb.go_ok ));
 sg13g2_dfrbp_1 _1073_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net111),
    .D(_0083_),
    .Q_N(_0422_),
    .Q(\tb.key_saved[0] ));
 sg13g2_dfrbp_1 _1074_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net103),
    .D(_0084_),
    .Q_N(_0421_),
    .Q(\tb.key_saved[1] ));
 sg13g2_dfrbp_1 _1075_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net95),
    .D(_0085_),
    .Q_N(_0420_),
    .Q(\tb.key_saved[2] ));
 sg13g2_dfrbp_1 _1076_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net87),
    .D(_0086_),
    .Q_N(_0419_),
    .Q(\tb.key_saved[3] ));
 sg13g2_dfrbp_1 _1077_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net77),
    .D(_0087_),
    .Q_N(_0418_),
    .Q(\tb.val_saved[0] ));
 sg13g2_dfrbp_1 _1078_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net69),
    .D(_0088_),
    .Q_N(_0417_),
    .Q(\tb.val_saved[1] ));
 sg13g2_dfrbp_1 _1079_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net61),
    .D(_0089_),
    .Q_N(_0416_),
    .Q(\tb.val_saved[2] ));
 sg13g2_dfrbp_1 _1080_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net53),
    .D(_0090_),
    .Q_N(_0415_),
    .Q(\tb.val_saved[3] ));
 sg13g2_dfrbp_1 _1081_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net42),
    .D(_0091_),
    .Q_N(_0414_),
    .Q(\tb.hash_saved[0] ));
 sg13g2_dfrbp_1 _1082_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net33),
    .D(_0092_),
    .Q_N(_0413_),
    .Q(\tb.hash_saved[1] ));
 sg13g2_dfrbp_1 _1083_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net115),
    .D(_0093_),
    .Q_N(_0412_),
    .Q(\tb.hash_saved[2] ));
 sg13g2_dfrbp_1 _1084_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net99),
    .D(net200),
    .Q_N(_0411_),
    .Q(\tb.mem[0][0] ));
 sg13g2_dfrbp_1 _1085_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net81),
    .D(net247),
    .Q_N(_0410_),
    .Q(\tb.mem[0][1] ));
 sg13g2_dfrbp_1 _1086_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net65),
    .D(_0096_),
    .Q_N(_0409_),
    .Q(\tb.mem[0][2] ));
 sg13g2_dfrbp_1 _1087_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net46),
    .D(net171),
    .Q_N(_0408_),
    .Q(\tb.mem[0][3] ));
 sg13g2_dfrbp_1 _1088_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net163),
    .D(net235),
    .Q_N(_0407_),
    .Q(\tb.mem[0][4] ));
 sg13g2_dfrbp_1 _1089_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net91),
    .D(net249),
    .Q_N(_0406_),
    .Q(\tb.mem[0][5] ));
 sg13g2_dfrbp_1 _1090_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net57),
    .D(net237),
    .Q_N(_0405_),
    .Q(\tb.mem[0][6] ));
 sg13g2_dfrbp_1 _1091_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net107),
    .D(net276),
    .Q_N(_0404_),
    .Q(\tb.mem[0][7] ));
 sg13g2_dfrbp_1 _1092_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net38),
    .D(_0102_),
    .Q_N(_0403_),
    .Q(\tb.mem[7][8] ));
 sg13g2_tiehi _1071__29 (.L_HI(net29));
 sg13g2_tiehi _0998__30 (.L_HI(net30));
 sg13g2_tiehi _1047__31 (.L_HI(net31));
 sg13g2_tiehi _0997__32 (.L_HI(net32));
 sg13g2_tiehi _1082__33 (.L_HI(net33));
 sg13g2_tiehi _0996__34 (.L_HI(net34));
 sg13g2_tiehi _1046__35 (.L_HI(net35));
 sg13g2_tiehi _1070__36 (.L_HI(net36));
 sg13g2_tiehi _1045__37 (.L_HI(net37));
 sg13g2_tiehi _1092__38 (.L_HI(net38));
 sg13g2_tiehi _1044__39 (.L_HI(net39));
 sg13g2_tiehi _1069__40 (.L_HI(net40));
 sg13g2_tiehi _1043__41 (.L_HI(net41));
 sg13g2_tiehi _1081__42 (.L_HI(net42));
 sg13g2_tiehi _1042__43 (.L_HI(net43));
 sg13g2_tiehi _1068__44 (.L_HI(net44));
 sg13g2_tiehi _1041__45 (.L_HI(net45));
 sg13g2_tiehi _1087__46 (.L_HI(net46));
 sg13g2_tiehi _1040__47 (.L_HI(net47));
 sg13g2_tiehi _1039__48 (.L_HI(net48));
 sg13g2_tiehi _1038__49 (.L_HI(net49));
 sg13g2_tiehi _1037__50 (.L_HI(net50));
 sg13g2_tiehi _1067__51 (.L_HI(net51));
 sg13g2_tiehi _1036__52 (.L_HI(net52));
 sg13g2_tiehi _1080__53 (.L_HI(net53));
 sg13g2_tiehi _1035__54 (.L_HI(net54));
 sg13g2_tiehi _1066__55 (.L_HI(net55));
 sg13g2_tiehi _1034__56 (.L_HI(net56));
 sg13g2_tiehi _1090__57 (.L_HI(net57));
 sg13g2_tiehi _1033__58 (.L_HI(net58));
 sg13g2_tiehi _1065__59 (.L_HI(net59));
 sg13g2_tiehi _1032__60 (.L_HI(net60));
 sg13g2_tiehi _1079__61 (.L_HI(net61));
 sg13g2_tiehi _1031__62 (.L_HI(net62));
 sg13g2_tiehi _1064__63 (.L_HI(net63));
 sg13g2_tiehi _1030__64 (.L_HI(net64));
 sg13g2_tiehi _1086__65 (.L_HI(net65));
 sg13g2_tiehi _1029__66 (.L_HI(net66));
 sg13g2_tiehi _1063__67 (.L_HI(net67));
 sg13g2_tiehi _1028__68 (.L_HI(net68));
 sg13g2_tiehi _1078__69 (.L_HI(net69));
 sg13g2_tiehi _1027__70 (.L_HI(net70));
 sg13g2_tiehi _1062__71 (.L_HI(net71));
 sg13g2_tiehi _1026__72 (.L_HI(net72));
 sg13g2_tiehi _0995__73 (.L_HI(net73));
 sg13g2_tiehi _1025__74 (.L_HI(net74));
 sg13g2_tiehi _1061__75 (.L_HI(net75));
 sg13g2_tiehi _1024__76 (.L_HI(net76));
 sg13g2_tiehi _1077__77 (.L_HI(net77));
 sg13g2_tiehi _1023__78 (.L_HI(net78));
 sg13g2_tiehi _1060__79 (.L_HI(net79));
 sg13g2_tiehi _1022__80 (.L_HI(net80));
 sg13g2_tiehi _1085__81 (.L_HI(net81));
 sg13g2_tiehi _1021__82 (.L_HI(net82));
 sg13g2_tiehi _1059__83 (.L_HI(net83));
 sg13g2_tiehi _1020__84 (.L_HI(net84));
 sg13g2_tiehi _1058__85 (.L_HI(net85));
 sg13g2_tiehi _1019__86 (.L_HI(net86));
 sg13g2_tiehi _1076__87 (.L_HI(net87));
 sg13g2_tiehi _1018__88 (.L_HI(net88));
 sg13g2_tiehi _1057__89 (.L_HI(net89));
 sg13g2_tiehi _1017__90 (.L_HI(net90));
 sg13g2_tiehi _1089__91 (.L_HI(net91));
 sg13g2_tiehi _1016__92 (.L_HI(net92));
 sg13g2_tiehi _1056__93 (.L_HI(net93));
 sg13g2_tiehi _1015__94 (.L_HI(net94));
 sg13g2_tiehi _1075__95 (.L_HI(net95));
 sg13g2_tiehi _1014__96 (.L_HI(net96));
 sg13g2_tiehi _1055__97 (.L_HI(net97));
 sg13g2_tiehi _1013__98 (.L_HI(net98));
 sg13g2_tiehi _1084__99 (.L_HI(net99));
 sg13g2_tiehi _1012__100 (.L_HI(net100));
 sg13g2_tiehi _1054__101 (.L_HI(net101));
 sg13g2_tiehi _1011__102 (.L_HI(net102));
 sg13g2_tiehi _1074__103 (.L_HI(net103));
 sg13g2_tiehi _1010__104 (.L_HI(net104));
 sg13g2_tiehi _1053__105 (.L_HI(net105));
 sg13g2_tiehi _1009__106 (.L_HI(net106));
 sg13g2_tiehi _1091__107 (.L_HI(net107));
 sg13g2_tiehi _1008__108 (.L_HI(net108));
 sg13g2_tiehi _1052__109 (.L_HI(net109));
 sg13g2_tiehi _1007__110 (.L_HI(net110));
 sg13g2_tiehi _1073__111 (.L_HI(net111));
 sg13g2_tiehi _1006__112 (.L_HI(net112));
 sg13g2_tiehi _1051__113 (.L_HI(net113));
 sg13g2_tiehi _1005__114 (.L_HI(net114));
 sg13g2_tiehi _1083__115 (.L_HI(net115));
 sg13g2_tiehi _1004__116 (.L_HI(net116));
 sg13g2_tiehi _1050__117 (.L_HI(net117));
 sg13g2_tiehi _1003__118 (.L_HI(net158));
 sg13g2_tiehi _1072__119 (.L_HI(net159));
 sg13g2_tiehi _1002__120 (.L_HI(net160));
 sg13g2_tiehi _1049__121 (.L_HI(net161));
 sg13g2_tiehi _1001__122 (.L_HI(net162));
 sg13g2_tiehi _1088__123 (.L_HI(net163));
 sg13g2_tiehi _1000__124 (.L_HI(net164));
 sg13g2_tiehi _1048__125 (.L_HI(net165));
 sg13g2_tiehi tt_um_save_buffer_hash_table_126 (.L_HI(net166));
 sg13g2_tiehi tt_um_save_buffer_hash_table_127 (.L_HI(net167));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_save_buffer_hash_table_13 (.L_LO(net13));
 sg13g2_tielo tt_um_save_buffer_hash_table_14 (.L_LO(net14));
 sg13g2_tielo tt_um_save_buffer_hash_table_15 (.L_LO(net15));
 sg13g2_tielo tt_um_save_buffer_hash_table_16 (.L_LO(net16));
 sg13g2_tielo tt_um_save_buffer_hash_table_17 (.L_LO(net17));
 sg13g2_tielo tt_um_save_buffer_hash_table_18 (.L_LO(net18));
 sg13g2_tielo tt_um_save_buffer_hash_table_19 (.L_LO(net19));
 sg13g2_tielo tt_um_save_buffer_hash_table_20 (.L_LO(net20));
 sg13g2_tielo tt_um_save_buffer_hash_table_21 (.L_LO(net21));
 sg13g2_tielo tt_um_save_buffer_hash_table_22 (.L_LO(net22));
 sg13g2_tielo tt_um_save_buffer_hash_table_23 (.L_LO(net23));
 sg13g2_tielo tt_um_save_buffer_hash_table_24 (.L_LO(net24));
 sg13g2_tielo tt_um_save_buffer_hash_table_25 (.L_LO(net25));
 sg13g2_tielo tt_um_save_buffer_hash_table_26 (.L_LO(net26));
 sg13g2_tielo tt_um_save_buffer_hash_table_27 (.L_LO(net27));
 sg13g2_tiehi _0999__28 (.L_HI(net28));
 sg13g2_buf_4 fanout118 (.X(net118),
    .A(_0336_));
 sg13g2_buf_4 fanout119 (.X(net119),
    .A(_0314_));
 sg13g2_buf_2 fanout120 (.A(_0294_),
    .X(net120));
 sg13g2_buf_4 fanout121 (.X(net121),
    .A(_0287_));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(_0267_));
 sg13g2_buf_2 fanout123 (.A(_0256_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_0245_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_0233_),
    .X(net125));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(_0226_));
 sg13g2_buf_2 fanout127 (.A(_0214_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(net131),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(net131),
    .X(net129));
 sg13g2_buf_1 fanout130 (.A(net131),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_0379_),
    .X(net131));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(net170));
 sg13g2_buf_4 fanout133 (.X(net133),
    .A(net168));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(net308));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(net216));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(\tb.key_saved[3] ));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(\tb.key_saved[2] ));
 sg13g2_buf_4 fanout138 (.X(net138),
    .A(\tb.key_saved[1] ));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(net309));
 sg13g2_buf_2 fanout140 (.A(\tb.cursor[2] ),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(\tb.cursor[1] ),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(net303),
    .X(net142));
 sg13g2_buf_4 fanout143 (.X(net143),
    .A(_0002_));
 sg13g2_buf_2 fanout144 (.A(_0002_),
    .X(net144));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(net147));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(net147));
 sg13g2_buf_2 fanout147 (.A(_0001_),
    .X(net147));
 sg13g2_buf_8 fanout148 (.A(net150),
    .X(net148));
 sg13g2_buf_4 fanout149 (.X(net149),
    .A(net150));
 sg13g2_buf_8 fanout150 (.A(_0000_),
    .X(net150));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(net154));
 sg13g2_buf_2 fanout152 (.A(net154),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(net154),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(net157),
    .X(net154));
 sg13g2_buf_4 fanout155 (.X(net155),
    .A(net157));
 sg13g2_buf_2 fanout156 (.A(net157),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(rst_n),
    .X(net157));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_tielo tt_um_save_buffer_hash_table_12 (.L_LO(net12));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_4_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_12_0_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\tb.val_saved[2] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0016_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold3 (.A(\tb.val_saved[3] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0097_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold5 (.A(\tb.mem[6][5] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0043_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold7 (.A(\tb.mem[4][3] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold8 (.A(\tb.mem[1][5] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0063_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold10 (.A(\tb.mem[6][3] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold11 (.A(\tb.mem[2][4] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0026_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold13 (.A(\tb.mem[7][5] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0035_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold15 (.A(\tb.mem[3][4] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0018_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold17 (.A(\tb.mem[7][7] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0037_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold19 (.A(\tb.mem[5][3] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold20 (.A(\tb.mem[6][7] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0045_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold22 (.A(\tb.mem[7][2] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold23 (.A(\tb.mem[2][5] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0027_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold25 (.A(\tb.mem[5][0] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0050_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold27 (.A(\tb.mem[2][0] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0022_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold29 (.A(\tb.mem[5][1] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0051_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold31 (.A(\tb.mem[4][2] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold32 (.A(\tb.mem[0][0] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0094_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold34 (.A(\tb.mem[3][1] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0015_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold36 (.A(\tb.mem[6][2] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold37 (.A(\tb.mem[4][0] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0006_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold39 (.A(\tb.mem[1][2] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold40 (.A(\tb.mem[1][1] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0059_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold42 (.A(\tb.mem[5][2] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold43 (.A(\tb.mem[3][7] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0021_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold45 (.A(\tb.mem[2][7] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0029_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold47 (.A(\tb.mem[1][6] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0064_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold49 (.A(\tb.val_saved[0] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0014_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold51 (.A(\tb.mem[3][5] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0019_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold53 (.A(\tb.mem[2][2] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold54 (.A(\tb.mem[1][4] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0062_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold56 (.A(\tb.mem[3][6] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0020_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold58 (.A(\tb.mem[1][0] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold59 (.A(\tb.mem[7][6] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0036_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold61 (.A(\tb.mem[4][6] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0012_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold63 (.A(\tb.mem[5][7] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0057_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold65 (.A(\tb.mem[5][6] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0056_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold67 (.A(\tb.mem[0][4] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0098_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold69 (.A(\tb.mem[0][6] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0100_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold71 (.A(\tb.mem[2][1] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0023_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold73 (.A(\tb.mem[4][7] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0013_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold75 (.A(\tb.mem[4][4] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0010_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold77 (.A(\tb.mem[1][7] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0065_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold79 (.A(\tb.mem[0][1] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0095_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold81 (.A(\tb.mem[0][5] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0099_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold83 (.A(\tb.mem[6][0] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold84 (.A(\tb.mem[2][6] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0028_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold86 (.A(\tb.mem[5][5] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0055_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold88 (.A(\tb.mem[7][4] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0034_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold90 (.A(\tb.mem[0][2] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold91 (.A(\tb.mem[4][5] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0011_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold93 (.A(\tb.mem[1][3] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold94 (.A(\tb.mem[2][3] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold95 (.A(\tb.mem[7][0] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold96 (.A(\tb.mem[7][1] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0031_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold98 (.A(\tb.mem[3][3] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold99 (.A(\tb.mem[7][3] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold100 (.A(\tb.mem[6][1] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0039_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold102 (.A(\tb.mem[4][1] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0007_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold104 (.A(\tb.mem[6][4] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0042_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold106 (.A(\tb.mem[6][6] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0044_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold108 (.A(\tb.mem[0][7] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0101_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold110 (.A(\tb.mem[5][4] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0054_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold112 (.A(uio_out[6]),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0072_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold114 (.A(uio_out[7]),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold115 (.A(\tb.cursor[3] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0081_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold117 (.A(uo_out[2]),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold118 (.A(uo_out[3]),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold119 (.A(uo_out[1]),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold120 (.A(uo_out[0]),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold121 (.A(\tb.hash_saved[0] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold122 (.A(\tb.hash_saved[1] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold123 (.A(\tb.go_ok ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0378_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0082_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold126 (.A(\tb.mem[0][8] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold127 (.A(\tb.mem[7][8] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold128 (.A(\tb.mem[3][8] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold129 (.A(\tb.mem[2][8] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold130 (.A(\tb.mem[5][8] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0344_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold132 (.A(\tb.mem[1][8] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold133 (.A(\tb.hash_saved[2] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold134 (.A(\tb.mem[4][8] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0066_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold136 (.A(\tb.state ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold137 (.A(\tb.mem[6][8] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0003_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0078_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold140 (.A(\tb.cursor[0] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold141 (.A(\tb.val_saved[1] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold142 (.A(\tb.key_saved[0] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0003_),
    .X(net310));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_4 FILLER_16_161 ();
 sg13g2_fill_1 FILLER_16_165 ();
 sg13g2_decap_8 FILLER_16_170 ();
 sg13g2_decap_8 FILLER_16_177 ();
 sg13g2_decap_8 FILLER_16_184 ();
 sg13g2_decap_8 FILLER_16_191 ();
 sg13g2_decap_8 FILLER_16_198 ();
 sg13g2_decap_8 FILLER_16_205 ();
 sg13g2_decap_8 FILLER_16_212 ();
 sg13g2_decap_8 FILLER_16_219 ();
 sg13g2_decap_8 FILLER_16_226 ();
 sg13g2_decap_8 FILLER_16_233 ();
 sg13g2_decap_8 FILLER_16_240 ();
 sg13g2_decap_8 FILLER_16_247 ();
 sg13g2_decap_8 FILLER_16_254 ();
 sg13g2_decap_8 FILLER_16_261 ();
 sg13g2_decap_8 FILLER_16_268 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_fill_2 FILLER_16_308 ();
 sg13g2_fill_1 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_decap_8 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_349 ();
 sg13g2_decap_8 FILLER_16_356 ();
 sg13g2_decap_8 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_decap_8 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_75 ();
 sg13g2_decap_8 FILLER_17_82 ();
 sg13g2_fill_2 FILLER_17_89 ();
 sg13g2_fill_1 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_95 ();
 sg13g2_decap_8 FILLER_17_102 ();
 sg13g2_decap_8 FILLER_17_109 ();
 sg13g2_decap_8 FILLER_17_116 ();
 sg13g2_decap_8 FILLER_17_123 ();
 sg13g2_decap_8 FILLER_17_130 ();
 sg13g2_decap_4 FILLER_17_137 ();
 sg13g2_fill_2 FILLER_17_141 ();
 sg13g2_decap_8 FILLER_17_150 ();
 sg13g2_decap_4 FILLER_17_157 ();
 sg13g2_decap_8 FILLER_17_187 ();
 sg13g2_fill_2 FILLER_17_194 ();
 sg13g2_decap_8 FILLER_17_199 ();
 sg13g2_fill_1 FILLER_17_206 ();
 sg13g2_fill_2 FILLER_17_212 ();
 sg13g2_fill_1 FILLER_17_214 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_4 FILLER_17_259 ();
 sg13g2_fill_1 FILLER_17_263 ();
 sg13g2_fill_1 FILLER_17_267 ();
 sg13g2_decap_8 FILLER_17_298 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_fill_2 FILLER_17_353 ();
 sg13g2_fill_2 FILLER_17_358 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_fill_1 FILLER_18_63 ();
 sg13g2_fill_1 FILLER_18_73 ();
 sg13g2_fill_1 FILLER_18_100 ();
 sg13g2_fill_2 FILLER_18_110 ();
 sg13g2_fill_1 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_131 ();
 sg13g2_fill_1 FILLER_18_164 ();
 sg13g2_fill_2 FILLER_18_205 ();
 sg13g2_decap_8 FILLER_18_242 ();
 sg13g2_decap_4 FILLER_18_249 ();
 sg13g2_fill_2 FILLER_18_337 ();
 sg13g2_fill_1 FILLER_18_379 ();
 sg13g2_decap_8 FILLER_18_393 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_4 FILLER_19_49 ();
 sg13g2_fill_2 FILLER_19_53 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_fill_2 FILLER_19_161 ();
 sg13g2_fill_1 FILLER_19_186 ();
 sg13g2_fill_2 FILLER_19_282 ();
 sg13g2_fill_1 FILLER_19_310 ();
 sg13g2_fill_1 FILLER_19_342 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_fill_2 FILLER_20_70 ();
 sg13g2_fill_2 FILLER_20_76 ();
 sg13g2_fill_1 FILLER_20_94 ();
 sg13g2_decap_4 FILLER_20_99 ();
 sg13g2_fill_1 FILLER_20_103 ();
 sg13g2_fill_2 FILLER_20_120 ();
 sg13g2_fill_1 FILLER_20_194 ();
 sg13g2_fill_2 FILLER_20_233 ();
 sg13g2_fill_1 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_250 ();
 sg13g2_decap_8 FILLER_20_257 ();
 sg13g2_decap_4 FILLER_20_264 ();
 sg13g2_fill_1 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_316 ();
 sg13g2_fill_2 FILLER_20_326 ();
 sg13g2_fill_2 FILLER_20_381 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_fill_1 FILLER_21_56 ();
 sg13g2_fill_1 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_100 ();
 sg13g2_decap_8 FILLER_21_138 ();
 sg13g2_fill_2 FILLER_21_145 ();
 sg13g2_fill_1 FILLER_21_147 ();
 sg13g2_fill_2 FILLER_21_174 ();
 sg13g2_fill_1 FILLER_21_223 ();
 sg13g2_fill_1 FILLER_21_234 ();
 sg13g2_fill_2 FILLER_21_356 ();
 sg13g2_fill_1 FILLER_21_396 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_fill_1 FILLER_22_49 ();
 sg13g2_fill_2 FILLER_22_126 ();
 sg13g2_fill_2 FILLER_22_137 ();
 sg13g2_fill_1 FILLER_22_139 ();
 sg13g2_decap_4 FILLER_22_145 ();
 sg13g2_fill_2 FILLER_22_149 ();
 sg13g2_decap_8 FILLER_22_209 ();
 sg13g2_decap_8 FILLER_22_216 ();
 sg13g2_decap_8 FILLER_22_223 ();
 sg13g2_fill_2 FILLER_22_230 ();
 sg13g2_fill_2 FILLER_22_240 ();
 sg13g2_fill_1 FILLER_22_242 ();
 sg13g2_fill_1 FILLER_22_310 ();
 sg13g2_fill_1 FILLER_22_375 ();
 sg13g2_fill_2 FILLER_22_381 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_104 ();
 sg13g2_decap_4 FILLER_23_136 ();
 sg13g2_fill_1 FILLER_23_171 ();
 sg13g2_fill_1 FILLER_23_198 ();
 sg13g2_fill_1 FILLER_23_208 ();
 sg13g2_fill_2 FILLER_23_230 ();
 sg13g2_fill_1 FILLER_23_250 ();
 sg13g2_fill_1 FILLER_23_335 ();
 sg13g2_fill_1 FILLER_23_349 ();
 sg13g2_fill_1 FILLER_23_359 ();
 sg13g2_fill_1 FILLER_23_374 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_35 ();
 sg13g2_fill_1 FILLER_24_111 ();
 sg13g2_fill_1 FILLER_24_116 ();
 sg13g2_fill_1 FILLER_24_120 ();
 sg13g2_fill_2 FILLER_24_125 ();
 sg13g2_fill_2 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_fill_2 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_255 ();
 sg13g2_fill_1 FILLER_24_343 ();
 sg13g2_fill_1 FILLER_24_375 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_fill_2 FILLER_25_28 ();
 sg13g2_fill_1 FILLER_25_30 ();
 sg13g2_fill_2 FILLER_25_78 ();
 sg13g2_fill_2 FILLER_25_94 ();
 sg13g2_fill_1 FILLER_25_109 ();
 sg13g2_fill_1 FILLER_25_151 ();
 sg13g2_fill_2 FILLER_25_190 ();
 sg13g2_fill_2 FILLER_25_196 ();
 sg13g2_fill_2 FILLER_25_201 ();
 sg13g2_decap_4 FILLER_25_238 ();
 sg13g2_fill_1 FILLER_25_242 ();
 sg13g2_decap_4 FILLER_25_248 ();
 sg13g2_fill_1 FILLER_25_252 ();
 sg13g2_fill_1 FILLER_25_279 ();
 sg13g2_fill_2 FILLER_25_289 ();
 sg13g2_fill_2 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_4 FILLER_26_35 ();
 sg13g2_fill_1 FILLER_26_86 ();
 sg13g2_fill_1 FILLER_26_158 ();
 sg13g2_fill_1 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_178 ();
 sg13g2_fill_1 FILLER_26_180 ();
 sg13g2_fill_1 FILLER_26_207 ();
 sg13g2_decap_4 FILLER_26_219 ();
 sg13g2_fill_2 FILLER_26_257 ();
 sg13g2_fill_1 FILLER_26_259 ();
 sg13g2_fill_1 FILLER_26_273 ();
 sg13g2_fill_2 FILLER_26_284 ();
 sg13g2_fill_1 FILLER_26_286 ();
 sg13g2_fill_2 FILLER_26_338 ();
 sg13g2_fill_2 FILLER_26_366 ();
 sg13g2_fill_2 FILLER_26_381 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_4 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_32 ();
 sg13g2_fill_2 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_111 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_fill_1 FILLER_27_181 ();
 sg13g2_fill_2 FILLER_27_189 ();
 sg13g2_fill_1 FILLER_27_191 ();
 sg13g2_fill_2 FILLER_27_196 ();
 sg13g2_fill_1 FILLER_27_203 ();
 sg13g2_decap_4 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_240 ();
 sg13g2_fill_2 FILLER_27_247 ();
 sg13g2_fill_1 FILLER_27_249 ();
 sg13g2_fill_2 FILLER_27_279 ();
 sg13g2_fill_1 FILLER_27_281 ();
 sg13g2_fill_1 FILLER_27_306 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_fill_2 FILLER_27_376 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_fill_1 FILLER_28_87 ();
 sg13g2_fill_2 FILLER_28_148 ();
 sg13g2_fill_1 FILLER_28_209 ();
 sg13g2_fill_1 FILLER_28_304 ();
 sg13g2_fill_1 FILLER_28_313 ();
 sg13g2_fill_1 FILLER_28_344 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_fill_2 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_97 ();
 sg13g2_fill_1 FILLER_29_131 ();
 sg13g2_decap_8 FILLER_29_136 ();
 sg13g2_fill_2 FILLER_29_143 ();
 sg13g2_fill_2 FILLER_29_157 ();
 sg13g2_fill_1 FILLER_29_225 ();
 sg13g2_fill_2 FILLER_29_234 ();
 sg13g2_decap_4 FILLER_29_250 ();
 sg13g2_fill_1 FILLER_29_272 ();
 sg13g2_decap_8 FILLER_29_303 ();
 sg13g2_fill_2 FILLER_29_310 ();
 sg13g2_fill_1 FILLER_29_328 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_fill_2 FILLER_30_42 ();
 sg13g2_fill_1 FILLER_30_44 ();
 sg13g2_fill_1 FILLER_30_74 ();
 sg13g2_fill_1 FILLER_30_79 ();
 sg13g2_fill_2 FILLER_30_88 ();
 sg13g2_fill_1 FILLER_30_103 ();
 sg13g2_fill_2 FILLER_30_132 ();
 sg13g2_decap_8 FILLER_30_150 ();
 sg13g2_fill_2 FILLER_30_203 ();
 sg13g2_fill_1 FILLER_30_205 ();
 sg13g2_decap_4 FILLER_30_210 ();
 sg13g2_fill_2 FILLER_30_214 ();
 sg13g2_decap_8 FILLER_30_229 ();
 sg13g2_decap_4 FILLER_30_252 ();
 sg13g2_fill_1 FILLER_30_268 ();
 sg13g2_decap_4 FILLER_30_320 ();
 sg13g2_fill_1 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_fill_1 FILLER_31_49 ();
 sg13g2_fill_2 FILLER_31_81 ();
 sg13g2_fill_1 FILLER_31_109 ();
 sg13g2_fill_2 FILLER_31_122 ();
 sg13g2_fill_1 FILLER_31_168 ();
 sg13g2_decap_4 FILLER_31_221 ();
 sg13g2_fill_1 FILLER_31_225 ();
 sg13g2_fill_2 FILLER_31_263 ();
 sg13g2_decap_8 FILLER_31_300 ();
 sg13g2_fill_2 FILLER_31_307 ();
 sg13g2_fill_1 FILLER_31_309 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_4 FILLER_32_56 ();
 sg13g2_fill_1 FILLER_32_60 ();
 sg13g2_fill_2 FILLER_32_65 ();
 sg13g2_fill_1 FILLER_32_67 ();
 sg13g2_fill_2 FILLER_32_97 ();
 sg13g2_decap_4 FILLER_32_104 ();
 sg13g2_fill_2 FILLER_32_108 ();
 sg13g2_fill_1 FILLER_32_113 ();
 sg13g2_fill_2 FILLER_32_132 ();
 sg13g2_fill_1 FILLER_32_134 ();
 sg13g2_decap_4 FILLER_32_139 ();
 sg13g2_fill_2 FILLER_32_143 ();
 sg13g2_decap_8 FILLER_32_149 ();
 sg13g2_fill_2 FILLER_32_156 ();
 sg13g2_decap_8 FILLER_32_163 ();
 sg13g2_decap_4 FILLER_32_170 ();
 sg13g2_fill_2 FILLER_32_188 ();
 sg13g2_decap_8 FILLER_32_204 ();
 sg13g2_decap_4 FILLER_32_211 ();
 sg13g2_fill_2 FILLER_32_215 ();
 sg13g2_decap_8 FILLER_32_227 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_fill_2 FILLER_32_245 ();
 sg13g2_fill_1 FILLER_32_247 ();
 sg13g2_fill_2 FILLER_32_263 ();
 sg13g2_fill_1 FILLER_32_313 ();
 sg13g2_fill_1 FILLER_32_349 ();
 sg13g2_fill_2 FILLER_32_375 ();
 sg13g2_fill_2 FILLER_32_398 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_fill_2 FILLER_33_77 ();
 sg13g2_fill_2 FILLER_33_92 ();
 sg13g2_fill_1 FILLER_33_133 ();
 sg13g2_fill_2 FILLER_33_165 ();
 sg13g2_fill_2 FILLER_33_179 ();
 sg13g2_decap_4 FILLER_33_211 ();
 sg13g2_fill_1 FILLER_33_249 ();
 sg13g2_fill_1 FILLER_33_268 ();
 sg13g2_fill_1 FILLER_33_308 ();
 sg13g2_decap_4 FILLER_33_317 ();
 sg13g2_fill_1 FILLER_33_321 ();
 sg13g2_decap_4 FILLER_33_335 ();
 sg13g2_fill_2 FILLER_33_339 ();
 sg13g2_fill_2 FILLER_33_370 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_4 FILLER_34_70 ();
 sg13g2_fill_1 FILLER_34_122 ();
 sg13g2_fill_1 FILLER_34_186 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_fill_1 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_233 ();
 sg13g2_decap_4 FILLER_34_240 ();
 sg13g2_fill_2 FILLER_34_301 ();
 sg13g2_fill_1 FILLER_34_303 ();
 sg13g2_fill_2 FILLER_34_317 ();
 sg13g2_fill_2 FILLER_34_329 ();
 sg13g2_fill_1 FILLER_34_335 ();
 sg13g2_fill_2 FILLER_34_358 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_fill_1 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_89 ();
 sg13g2_decap_4 FILLER_35_96 ();
 sg13g2_fill_2 FILLER_35_100 ();
 sg13g2_fill_2 FILLER_35_157 ();
 sg13g2_fill_1 FILLER_35_159 ();
 sg13g2_fill_2 FILLER_35_197 ();
 sg13g2_fill_1 FILLER_35_204 ();
 sg13g2_fill_2 FILLER_35_223 ();
 sg13g2_fill_2 FILLER_35_255 ();
 sg13g2_decap_8 FILLER_35_274 ();
 sg13g2_fill_1 FILLER_35_284 ();
 sg13g2_fill_1 FILLER_35_346 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_fill_2 FILLER_36_105 ();
 sg13g2_fill_1 FILLER_36_107 ();
 sg13g2_fill_2 FILLER_36_134 ();
 sg13g2_fill_2 FILLER_36_150 ();
 sg13g2_fill_2 FILLER_36_166 ();
 sg13g2_fill_1 FILLER_36_168 ();
 sg13g2_fill_1 FILLER_36_225 ();
 sg13g2_fill_2 FILLER_36_236 ();
 sg13g2_fill_1 FILLER_36_238 ();
 sg13g2_decap_4 FILLER_36_248 ();
 sg13g2_fill_2 FILLER_36_261 ();
 sg13g2_fill_2 FILLER_36_271 ();
 sg13g2_fill_1 FILLER_36_273 ();
 sg13g2_fill_2 FILLER_36_283 ();
 sg13g2_fill_2 FILLER_36_298 ();
 sg13g2_fill_2 FILLER_36_304 ();
 sg13g2_fill_1 FILLER_36_309 ();
 sg13g2_decap_4 FILLER_36_313 ();
 sg13g2_fill_2 FILLER_36_317 ();
 sg13g2_decap_4 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_328 ();
 sg13g2_fill_2 FILLER_36_338 ();
 sg13g2_fill_1 FILLER_36_340 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_fill_2 FILLER_37_98 ();
 sg13g2_fill_1 FILLER_37_136 ();
 sg13g2_fill_2 FILLER_37_155 ();
 sg13g2_fill_1 FILLER_37_157 ();
 sg13g2_fill_2 FILLER_37_184 ();
 sg13g2_fill_1 FILLER_37_199 ();
 sg13g2_fill_1 FILLER_37_208 ();
 sg13g2_fill_2 FILLER_37_244 ();
 sg13g2_fill_1 FILLER_37_246 ();
 sg13g2_fill_1 FILLER_37_303 ();
 sg13g2_fill_1 FILLER_37_318 ();
 sg13g2_fill_1 FILLER_37_359 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_fill_2 FILLER_38_173 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_fill_1 FILLER_38_278 ();
 sg13g2_fill_2 FILLER_38_315 ();
 sg13g2_fill_1 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_343 ();
 sg13g2_fill_1 FILLER_38_348 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net12;
 assign uio_oe[1] = net13;
 assign uio_oe[2] = net14;
 assign uio_oe[3] = net15;
 assign uio_oe[4] = net16;
 assign uio_oe[5] = net17;
 assign uio_oe[6] = net166;
 assign uio_oe[7] = net167;
 assign uio_out[0] = net18;
 assign uio_out[1] = net19;
 assign uio_out[2] = net20;
 assign uio_out[3] = net21;
 assign uio_out[4] = net22;
 assign uio_out[5] = net23;
 assign uo_out[4] = net24;
 assign uo_out[5] = net25;
 assign uo_out[6] = net26;
 assign uo_out[7] = net27;
endmodule

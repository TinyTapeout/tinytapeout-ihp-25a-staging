module tt_um_rejunity_atari2600 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire \atari2600.address_bus_r[0] ;
 wire \atari2600.address_bus_r[10] ;
 wire \atari2600.address_bus_r[11] ;
 wire \atari2600.address_bus_r[12] ;
 wire \atari2600.address_bus_r[1] ;
 wire \atari2600.address_bus_r[2] ;
 wire \atari2600.address_bus_r[3] ;
 wire \atari2600.address_bus_r[4] ;
 wire \atari2600.address_bus_r[5] ;
 wire \atari2600.address_bus_r[6] ;
 wire \atari2600.address_bus_r[7] ;
 wire \atari2600.address_bus_r[8] ;
 wire \atari2600.address_bus_r[9] ;
 wire \atari2600.clk_counter[0] ;
 wire \atari2600.clk_counter[1] ;
 wire \atari2600.clk_counter[2] ;
 wire \atari2600.clk_counter[3] ;
 wire \atari2600.clk_counter[4] ;
 wire \atari2600.clk_counter[5] ;
 wire \atari2600.clk_counter[6] ;
 wire \atari2600.clk_counter[7] ;
 wire \atari2600.clk_counter[8] ;
 wire \atari2600.cpu.ABH[0] ;
 wire \atari2600.cpu.ABH[1] ;
 wire \atari2600.cpu.ABH[2] ;
 wire \atari2600.cpu.ABH[3] ;
 wire \atari2600.cpu.ABH[4] ;
 wire \atari2600.cpu.ABH[5] ;
 wire \atari2600.cpu.ABH[6] ;
 wire \atari2600.cpu.ABH[7] ;
 wire \atari2600.cpu.ABL[0] ;
 wire \atari2600.cpu.ABL[1] ;
 wire \atari2600.cpu.ABL[2] ;
 wire \atari2600.cpu.ABL[3] ;
 wire \atari2600.cpu.ABL[4] ;
 wire \atari2600.cpu.ABL[5] ;
 wire \atari2600.cpu.ABL[6] ;
 wire \atari2600.cpu.ABL[7] ;
 wire \atari2600.cpu.ADD[0] ;
 wire \atari2600.cpu.ADD[1] ;
 wire \atari2600.cpu.ADD[2] ;
 wire \atari2600.cpu.ADD[3] ;
 wire \atari2600.cpu.ADD[4] ;
 wire \atari2600.cpu.ADD[5] ;
 wire \atari2600.cpu.ADD[6] ;
 wire \atari2600.cpu.ADD[7] ;
 wire \atari2600.cpu.ALU.AI7 ;
 wire \atari2600.cpu.ALU.BI7 ;
 wire \atari2600.cpu.ALU.CO ;
 wire \atari2600.cpu.ALU.HC ;
 wire \atari2600.cpu.AXYS[0][0] ;
 wire \atari2600.cpu.AXYS[0][1] ;
 wire \atari2600.cpu.AXYS[0][2] ;
 wire \atari2600.cpu.AXYS[0][3] ;
 wire \atari2600.cpu.AXYS[0][4] ;
 wire \atari2600.cpu.AXYS[0][5] ;
 wire \atari2600.cpu.AXYS[0][6] ;
 wire \atari2600.cpu.AXYS[0][7] ;
 wire \atari2600.cpu.AXYS[1][0] ;
 wire \atari2600.cpu.AXYS[1][1] ;
 wire \atari2600.cpu.AXYS[1][2] ;
 wire \atari2600.cpu.AXYS[1][3] ;
 wire \atari2600.cpu.AXYS[1][4] ;
 wire \atari2600.cpu.AXYS[1][5] ;
 wire \atari2600.cpu.AXYS[1][6] ;
 wire \atari2600.cpu.AXYS[1][7] ;
 wire \atari2600.cpu.AXYS[2][0] ;
 wire \atari2600.cpu.AXYS[2][1] ;
 wire \atari2600.cpu.AXYS[2][2] ;
 wire \atari2600.cpu.AXYS[2][3] ;
 wire \atari2600.cpu.AXYS[2][4] ;
 wire \atari2600.cpu.AXYS[2][5] ;
 wire \atari2600.cpu.AXYS[2][6] ;
 wire \atari2600.cpu.AXYS[2][7] ;
 wire \atari2600.cpu.AXYS[3][0] ;
 wire \atari2600.cpu.AXYS[3][1] ;
 wire \atari2600.cpu.AXYS[3][2] ;
 wire \atari2600.cpu.AXYS[3][3] ;
 wire \atari2600.cpu.AXYS[3][4] ;
 wire \atari2600.cpu.AXYS[3][5] ;
 wire \atari2600.cpu.AXYS[3][6] ;
 wire \atari2600.cpu.AXYS[3][7] ;
 wire \atari2600.cpu.C ;
 wire \atari2600.cpu.D ;
 wire \atari2600.cpu.DIHOLD[0] ;
 wire \atari2600.cpu.DIHOLD[1] ;
 wire \atari2600.cpu.DIHOLD[2] ;
 wire \atari2600.cpu.DIHOLD[3] ;
 wire \atari2600.cpu.DIHOLD[4] ;
 wire \atari2600.cpu.DIHOLD[5] ;
 wire \atari2600.cpu.DIHOLD[6] ;
 wire \atari2600.cpu.DIHOLD[7] ;
 wire \atari2600.cpu.DIMUX[0] ;
 wire \atari2600.cpu.DIMUX[1] ;
 wire \atari2600.cpu.DIMUX[2] ;
 wire \atari2600.cpu.DIMUX[3] ;
 wire \atari2600.cpu.DIMUX[4] ;
 wire \atari2600.cpu.DIMUX[5] ;
 wire \atari2600.cpu.DIMUX[6] ;
 wire \atari2600.cpu.DIMUX[7] ;
 wire \atari2600.cpu.DI[0] ;
 wire \atari2600.cpu.DI[1] ;
 wire \atari2600.cpu.DI[2] ;
 wire \atari2600.cpu.DI[3] ;
 wire \atari2600.cpu.DI[4] ;
 wire \atari2600.cpu.DI[5] ;
 wire \atari2600.cpu.DI[6] ;
 wire \atari2600.cpu.DI[7] ;
 wire \atari2600.cpu.I ;
 wire \atari2600.cpu.IRHOLD[0] ;
 wire \atari2600.cpu.IRHOLD[1] ;
 wire \atari2600.cpu.IRHOLD[2] ;
 wire \atari2600.cpu.IRHOLD[3] ;
 wire \atari2600.cpu.IRHOLD[4] ;
 wire \atari2600.cpu.IRHOLD[5] ;
 wire \atari2600.cpu.IRHOLD[6] ;
 wire \atari2600.cpu.IRHOLD[7] ;
 wire \atari2600.cpu.IRHOLD_valid ;
 wire \atari2600.cpu.N ;
 wire \atari2600.cpu.PC[0] ;
 wire \atari2600.cpu.PC[10] ;
 wire \atari2600.cpu.PC[11] ;
 wire \atari2600.cpu.PC[12] ;
 wire \atari2600.cpu.PC[13] ;
 wire \atari2600.cpu.PC[14] ;
 wire \atari2600.cpu.PC[15] ;
 wire \atari2600.cpu.PC[1] ;
 wire \atari2600.cpu.PC[2] ;
 wire \atari2600.cpu.PC[3] ;
 wire \atari2600.cpu.PC[4] ;
 wire \atari2600.cpu.PC[5] ;
 wire \atari2600.cpu.PC[6] ;
 wire \atari2600.cpu.PC[7] ;
 wire \atari2600.cpu.PC[8] ;
 wire \atari2600.cpu.PC[9] ;
 wire \atari2600.cpu.V ;
 wire \atari2600.cpu.Z ;
 wire \atari2600.cpu.adc_bcd ;
 wire \atari2600.cpu.adc_sbc ;
 wire \atari2600.cpu.adj_bcd ;
 wire \atari2600.cpu.backwards ;
 wire \atari2600.cpu.bit_ins ;
 wire \atari2600.cpu.clc ;
 wire \atari2600.cpu.cld ;
 wire \atari2600.cpu.cli ;
 wire \atari2600.cpu.clv ;
 wire \atari2600.cpu.compare ;
 wire \atari2600.cpu.cond_code[0] ;
 wire \atari2600.cpu.cond_code[1] ;
 wire \atari2600.cpu.cond_code[2] ;
 wire \atari2600.cpu.dst_reg[0] ;
 wire \atari2600.cpu.dst_reg[1] ;
 wire \atari2600.cpu.inc ;
 wire \atari2600.cpu.index_y ;
 wire \atari2600.cpu.load_only ;
 wire \atari2600.cpu.load_reg ;
 wire \atari2600.cpu.op[0] ;
 wire \atari2600.cpu.op[1] ;
 wire \atari2600.cpu.op[2] ;
 wire \atari2600.cpu.op[3] ;
 wire \atari2600.cpu.php ;
 wire \atari2600.cpu.plp ;
 wire \atari2600.cpu.res ;
 wire \atari2600.cpu.rotate ;
 wire \atari2600.cpu.sec ;
 wire \atari2600.cpu.sed ;
 wire \atari2600.cpu.sei ;
 wire \atari2600.cpu.shift ;
 wire \atari2600.cpu.shift_right ;
 wire \atari2600.cpu.src_reg[0] ;
 wire \atari2600.cpu.src_reg[1] ;
 wire \atari2600.cpu.state[0] ;
 wire \atari2600.cpu.state[1] ;
 wire \atari2600.cpu.state[2] ;
 wire \atari2600.cpu.state[3] ;
 wire \atari2600.cpu.state[4] ;
 wire \atari2600.cpu.state[5] ;
 wire \atari2600.cpu.store ;
 wire \atari2600.cpu.write_back ;
 wire \atari2600.input_joystick_0[0] ;
 wire \atari2600.input_joystick_0[1] ;
 wire \atari2600.input_joystick_0[2] ;
 wire \atari2600.input_joystick_0[3] ;
 wire \atari2600.input_joystick_0[4] ;
 wire \atari2600.input_joystick_0[5] ;
 wire \atari2600.input_joystick_0[6] ;
 wire \atari2600.input_switches[0] ;
 wire \atari2600.input_switches[1] ;
 wire \atari2600.input_switches[2] ;
 wire \atari2600.input_switches[3] ;
 wire \atari2600.pia.dat_o[0] ;
 wire \atari2600.pia.dat_o[1] ;
 wire \atari2600.pia.dat_o[2] ;
 wire \atari2600.pia.dat_o[3] ;
 wire \atari2600.pia.dat_o[4] ;
 wire \atari2600.pia.dat_o[5] ;
 wire \atari2600.pia.dat_o[6] ;
 wire \atari2600.pia.dat_o[7] ;
 wire \atari2600.pia.diag[0] ;
 wire \atari2600.pia.diag[1] ;
 wire \atari2600.pia.diag[2] ;
 wire \atari2600.pia.diag[3] ;
 wire \atari2600.pia.diag[4] ;
 wire \atari2600.pia.diag[5] ;
 wire \atari2600.pia.diag[6] ;
 wire \atari2600.pia.diag[7] ;
 wire \atari2600.pia.instat[0] ;
 wire \atari2600.pia.instat[1] ;
 wire \atari2600.pia.interval[0] ;
 wire \atari2600.pia.interval[10] ;
 wire \atari2600.pia.interval[3] ;
 wire \atari2600.pia.interval[6] ;
 wire \atari2600.pia.reset_timer[0] ;
 wire \atari2600.pia.reset_timer[1] ;
 wire \atari2600.pia.reset_timer[2] ;
 wire \atari2600.pia.reset_timer[3] ;
 wire \atari2600.pia.reset_timer[4] ;
 wire \atari2600.pia.reset_timer[5] ;
 wire \atari2600.pia.reset_timer[6] ;
 wire \atari2600.pia.reset_timer[7] ;
 wire \atari2600.pia.swa_dir[0] ;
 wire \atari2600.pia.swa_dir[1] ;
 wire \atari2600.pia.swa_dir[2] ;
 wire \atari2600.pia.swa_dir[3] ;
 wire \atari2600.pia.swa_dir[4] ;
 wire \atari2600.pia.swa_dir[5] ;
 wire \atari2600.pia.swa_dir[6] ;
 wire \atari2600.pia.swa_dir[7] ;
 wire \atari2600.pia.swb_dir[2] ;
 wire \atari2600.pia.swb_dir[4] ;
 wire \atari2600.pia.swb_dir[5] ;
 wire \atari2600.pia.time_counter[0] ;
 wire \atari2600.pia.time_counter[10] ;
 wire \atari2600.pia.time_counter[11] ;
 wire \atari2600.pia.time_counter[12] ;
 wire \atari2600.pia.time_counter[13] ;
 wire \atari2600.pia.time_counter[14] ;
 wire \atari2600.pia.time_counter[15] ;
 wire \atari2600.pia.time_counter[16] ;
 wire \atari2600.pia.time_counter[17] ;
 wire \atari2600.pia.time_counter[18] ;
 wire \atari2600.pia.time_counter[19] ;
 wire \atari2600.pia.time_counter[1] ;
 wire \atari2600.pia.time_counter[20] ;
 wire \atari2600.pia.time_counter[21] ;
 wire \atari2600.pia.time_counter[22] ;
 wire \atari2600.pia.time_counter[23] ;
 wire \atari2600.pia.time_counter[2] ;
 wire \atari2600.pia.time_counter[3] ;
 wire \atari2600.pia.time_counter[4] ;
 wire \atari2600.pia.time_counter[5] ;
 wire \atari2600.pia.time_counter[6] ;
 wire \atari2600.pia.time_counter[7] ;
 wire \atari2600.pia.time_counter[8] ;
 wire \atari2600.pia.time_counter[9] ;
 wire \atari2600.pia.underflow ;
 wire \atari2600.ram[0][0] ;
 wire \atari2600.ram[0][1] ;
 wire \atari2600.ram[0][2] ;
 wire \atari2600.ram[0][3] ;
 wire \atari2600.ram[0][4] ;
 wire \atari2600.ram[0][5] ;
 wire \atari2600.ram[0][6] ;
 wire \atari2600.ram[0][7] ;
 wire \atari2600.ram[100][0] ;
 wire \atari2600.ram[100][1] ;
 wire \atari2600.ram[100][2] ;
 wire \atari2600.ram[100][3] ;
 wire \atari2600.ram[100][4] ;
 wire \atari2600.ram[100][5] ;
 wire \atari2600.ram[100][6] ;
 wire \atari2600.ram[100][7] ;
 wire \atari2600.ram[101][0] ;
 wire \atari2600.ram[101][1] ;
 wire \atari2600.ram[101][2] ;
 wire \atari2600.ram[101][3] ;
 wire \atari2600.ram[101][4] ;
 wire \atari2600.ram[101][5] ;
 wire \atari2600.ram[101][6] ;
 wire \atari2600.ram[101][7] ;
 wire \atari2600.ram[102][0] ;
 wire \atari2600.ram[102][1] ;
 wire \atari2600.ram[102][2] ;
 wire \atari2600.ram[102][3] ;
 wire \atari2600.ram[102][4] ;
 wire \atari2600.ram[102][5] ;
 wire \atari2600.ram[102][6] ;
 wire \atari2600.ram[102][7] ;
 wire \atari2600.ram[103][0] ;
 wire \atari2600.ram[103][1] ;
 wire \atari2600.ram[103][2] ;
 wire \atari2600.ram[103][3] ;
 wire \atari2600.ram[103][4] ;
 wire \atari2600.ram[103][5] ;
 wire \atari2600.ram[103][6] ;
 wire \atari2600.ram[103][7] ;
 wire \atari2600.ram[104][0] ;
 wire \atari2600.ram[104][1] ;
 wire \atari2600.ram[104][2] ;
 wire \atari2600.ram[104][3] ;
 wire \atari2600.ram[104][4] ;
 wire \atari2600.ram[104][5] ;
 wire \atari2600.ram[104][6] ;
 wire \atari2600.ram[104][7] ;
 wire \atari2600.ram[105][0] ;
 wire \atari2600.ram[105][1] ;
 wire \atari2600.ram[105][2] ;
 wire \atari2600.ram[105][3] ;
 wire \atari2600.ram[105][4] ;
 wire \atari2600.ram[105][5] ;
 wire \atari2600.ram[105][6] ;
 wire \atari2600.ram[105][7] ;
 wire \atari2600.ram[106][0] ;
 wire \atari2600.ram[106][1] ;
 wire \atari2600.ram[106][2] ;
 wire \atari2600.ram[106][3] ;
 wire \atari2600.ram[106][4] ;
 wire \atari2600.ram[106][5] ;
 wire \atari2600.ram[106][6] ;
 wire \atari2600.ram[106][7] ;
 wire \atari2600.ram[107][0] ;
 wire \atari2600.ram[107][1] ;
 wire \atari2600.ram[107][2] ;
 wire \atari2600.ram[107][3] ;
 wire \atari2600.ram[107][4] ;
 wire \atari2600.ram[107][5] ;
 wire \atari2600.ram[107][6] ;
 wire \atari2600.ram[107][7] ;
 wire \atari2600.ram[108][0] ;
 wire \atari2600.ram[108][1] ;
 wire \atari2600.ram[108][2] ;
 wire \atari2600.ram[108][3] ;
 wire \atari2600.ram[108][4] ;
 wire \atari2600.ram[108][5] ;
 wire \atari2600.ram[108][6] ;
 wire \atari2600.ram[108][7] ;
 wire \atari2600.ram[109][0] ;
 wire \atari2600.ram[109][1] ;
 wire \atari2600.ram[109][2] ;
 wire \atari2600.ram[109][3] ;
 wire \atari2600.ram[109][4] ;
 wire \atari2600.ram[109][5] ;
 wire \atari2600.ram[109][6] ;
 wire \atari2600.ram[109][7] ;
 wire \atari2600.ram[10][0] ;
 wire \atari2600.ram[10][1] ;
 wire \atari2600.ram[10][2] ;
 wire \atari2600.ram[10][3] ;
 wire \atari2600.ram[10][4] ;
 wire \atari2600.ram[10][5] ;
 wire \atari2600.ram[10][6] ;
 wire \atari2600.ram[10][7] ;
 wire \atari2600.ram[110][0] ;
 wire \atari2600.ram[110][1] ;
 wire \atari2600.ram[110][2] ;
 wire \atari2600.ram[110][3] ;
 wire \atari2600.ram[110][4] ;
 wire \atari2600.ram[110][5] ;
 wire \atari2600.ram[110][6] ;
 wire \atari2600.ram[110][7] ;
 wire \atari2600.ram[111][0] ;
 wire \atari2600.ram[111][1] ;
 wire \atari2600.ram[111][2] ;
 wire \atari2600.ram[111][3] ;
 wire \atari2600.ram[111][4] ;
 wire \atari2600.ram[111][5] ;
 wire \atari2600.ram[111][6] ;
 wire \atari2600.ram[111][7] ;
 wire \atari2600.ram[112][0] ;
 wire \atari2600.ram[112][1] ;
 wire \atari2600.ram[112][2] ;
 wire \atari2600.ram[112][3] ;
 wire \atari2600.ram[112][4] ;
 wire \atari2600.ram[112][5] ;
 wire \atari2600.ram[112][6] ;
 wire \atari2600.ram[112][7] ;
 wire \atari2600.ram[113][0] ;
 wire \atari2600.ram[113][1] ;
 wire \atari2600.ram[113][2] ;
 wire \atari2600.ram[113][3] ;
 wire \atari2600.ram[113][4] ;
 wire \atari2600.ram[113][5] ;
 wire \atari2600.ram[113][6] ;
 wire \atari2600.ram[113][7] ;
 wire \atari2600.ram[114][0] ;
 wire \atari2600.ram[114][1] ;
 wire \atari2600.ram[114][2] ;
 wire \atari2600.ram[114][3] ;
 wire \atari2600.ram[114][4] ;
 wire \atari2600.ram[114][5] ;
 wire \atari2600.ram[114][6] ;
 wire \atari2600.ram[114][7] ;
 wire \atari2600.ram[115][0] ;
 wire \atari2600.ram[115][1] ;
 wire \atari2600.ram[115][2] ;
 wire \atari2600.ram[115][3] ;
 wire \atari2600.ram[115][4] ;
 wire \atari2600.ram[115][5] ;
 wire \atari2600.ram[115][6] ;
 wire \atari2600.ram[115][7] ;
 wire \atari2600.ram[116][0] ;
 wire \atari2600.ram[116][1] ;
 wire \atari2600.ram[116][2] ;
 wire \atari2600.ram[116][3] ;
 wire \atari2600.ram[116][4] ;
 wire \atari2600.ram[116][5] ;
 wire \atari2600.ram[116][6] ;
 wire \atari2600.ram[116][7] ;
 wire \atari2600.ram[117][0] ;
 wire \atari2600.ram[117][1] ;
 wire \atari2600.ram[117][2] ;
 wire \atari2600.ram[117][3] ;
 wire \atari2600.ram[117][4] ;
 wire \atari2600.ram[117][5] ;
 wire \atari2600.ram[117][6] ;
 wire \atari2600.ram[117][7] ;
 wire \atari2600.ram[118][0] ;
 wire \atari2600.ram[118][1] ;
 wire \atari2600.ram[118][2] ;
 wire \atari2600.ram[118][3] ;
 wire \atari2600.ram[118][4] ;
 wire \atari2600.ram[118][5] ;
 wire \atari2600.ram[118][6] ;
 wire \atari2600.ram[118][7] ;
 wire \atari2600.ram[119][0] ;
 wire \atari2600.ram[119][1] ;
 wire \atari2600.ram[119][2] ;
 wire \atari2600.ram[119][3] ;
 wire \atari2600.ram[119][4] ;
 wire \atari2600.ram[119][5] ;
 wire \atari2600.ram[119][6] ;
 wire \atari2600.ram[119][7] ;
 wire \atari2600.ram[11][0] ;
 wire \atari2600.ram[11][1] ;
 wire \atari2600.ram[11][2] ;
 wire \atari2600.ram[11][3] ;
 wire \atari2600.ram[11][4] ;
 wire \atari2600.ram[11][5] ;
 wire \atari2600.ram[11][6] ;
 wire \atari2600.ram[11][7] ;
 wire \atari2600.ram[120][0] ;
 wire \atari2600.ram[120][1] ;
 wire \atari2600.ram[120][2] ;
 wire \atari2600.ram[120][3] ;
 wire \atari2600.ram[120][4] ;
 wire \atari2600.ram[120][5] ;
 wire \atari2600.ram[120][6] ;
 wire \atari2600.ram[120][7] ;
 wire \atari2600.ram[121][0] ;
 wire \atari2600.ram[121][1] ;
 wire \atari2600.ram[121][2] ;
 wire \atari2600.ram[121][3] ;
 wire \atari2600.ram[121][4] ;
 wire \atari2600.ram[121][5] ;
 wire \atari2600.ram[121][6] ;
 wire \atari2600.ram[121][7] ;
 wire \atari2600.ram[122][0] ;
 wire \atari2600.ram[122][1] ;
 wire \atari2600.ram[122][2] ;
 wire \atari2600.ram[122][3] ;
 wire \atari2600.ram[122][4] ;
 wire \atari2600.ram[122][5] ;
 wire \atari2600.ram[122][6] ;
 wire \atari2600.ram[122][7] ;
 wire \atari2600.ram[123][0] ;
 wire \atari2600.ram[123][1] ;
 wire \atari2600.ram[123][2] ;
 wire \atari2600.ram[123][3] ;
 wire \atari2600.ram[123][4] ;
 wire \atari2600.ram[123][5] ;
 wire \atari2600.ram[123][6] ;
 wire \atari2600.ram[123][7] ;
 wire \atari2600.ram[124][0] ;
 wire \atari2600.ram[124][1] ;
 wire \atari2600.ram[124][2] ;
 wire \atari2600.ram[124][3] ;
 wire \atari2600.ram[124][4] ;
 wire \atari2600.ram[124][5] ;
 wire \atari2600.ram[124][6] ;
 wire \atari2600.ram[124][7] ;
 wire \atari2600.ram[125][0] ;
 wire \atari2600.ram[125][1] ;
 wire \atari2600.ram[125][2] ;
 wire \atari2600.ram[125][3] ;
 wire \atari2600.ram[125][4] ;
 wire \atari2600.ram[125][5] ;
 wire \atari2600.ram[125][6] ;
 wire \atari2600.ram[125][7] ;
 wire \atari2600.ram[126][0] ;
 wire \atari2600.ram[126][1] ;
 wire \atari2600.ram[126][2] ;
 wire \atari2600.ram[126][3] ;
 wire \atari2600.ram[126][4] ;
 wire \atari2600.ram[126][5] ;
 wire \atari2600.ram[126][6] ;
 wire \atari2600.ram[126][7] ;
 wire \atari2600.ram[127][0] ;
 wire \atari2600.ram[127][1] ;
 wire \atari2600.ram[127][2] ;
 wire \atari2600.ram[127][3] ;
 wire \atari2600.ram[127][4] ;
 wire \atari2600.ram[127][5] ;
 wire \atari2600.ram[127][6] ;
 wire \atari2600.ram[127][7] ;
 wire \atari2600.ram[12][0] ;
 wire \atari2600.ram[12][1] ;
 wire \atari2600.ram[12][2] ;
 wire \atari2600.ram[12][3] ;
 wire \atari2600.ram[12][4] ;
 wire \atari2600.ram[12][5] ;
 wire \atari2600.ram[12][6] ;
 wire \atari2600.ram[12][7] ;
 wire \atari2600.ram[13][0] ;
 wire \atari2600.ram[13][1] ;
 wire \atari2600.ram[13][2] ;
 wire \atari2600.ram[13][3] ;
 wire \atari2600.ram[13][4] ;
 wire \atari2600.ram[13][5] ;
 wire \atari2600.ram[13][6] ;
 wire \atari2600.ram[13][7] ;
 wire \atari2600.ram[14][0] ;
 wire \atari2600.ram[14][1] ;
 wire \atari2600.ram[14][2] ;
 wire \atari2600.ram[14][3] ;
 wire \atari2600.ram[14][4] ;
 wire \atari2600.ram[14][5] ;
 wire \atari2600.ram[14][6] ;
 wire \atari2600.ram[14][7] ;
 wire \atari2600.ram[15][0] ;
 wire \atari2600.ram[15][1] ;
 wire \atari2600.ram[15][2] ;
 wire \atari2600.ram[15][3] ;
 wire \atari2600.ram[15][4] ;
 wire \atari2600.ram[15][5] ;
 wire \atari2600.ram[15][6] ;
 wire \atari2600.ram[15][7] ;
 wire \atari2600.ram[16][0] ;
 wire \atari2600.ram[16][1] ;
 wire \atari2600.ram[16][2] ;
 wire \atari2600.ram[16][3] ;
 wire \atari2600.ram[16][4] ;
 wire \atari2600.ram[16][5] ;
 wire \atari2600.ram[16][6] ;
 wire \atari2600.ram[16][7] ;
 wire \atari2600.ram[17][0] ;
 wire \atari2600.ram[17][1] ;
 wire \atari2600.ram[17][2] ;
 wire \atari2600.ram[17][3] ;
 wire \atari2600.ram[17][4] ;
 wire \atari2600.ram[17][5] ;
 wire \atari2600.ram[17][6] ;
 wire \atari2600.ram[17][7] ;
 wire \atari2600.ram[18][0] ;
 wire \atari2600.ram[18][1] ;
 wire \atari2600.ram[18][2] ;
 wire \atari2600.ram[18][3] ;
 wire \atari2600.ram[18][4] ;
 wire \atari2600.ram[18][5] ;
 wire \atari2600.ram[18][6] ;
 wire \atari2600.ram[18][7] ;
 wire \atari2600.ram[19][0] ;
 wire \atari2600.ram[19][1] ;
 wire \atari2600.ram[19][2] ;
 wire \atari2600.ram[19][3] ;
 wire \atari2600.ram[19][4] ;
 wire \atari2600.ram[19][5] ;
 wire \atari2600.ram[19][6] ;
 wire \atari2600.ram[19][7] ;
 wire \atari2600.ram[1][0] ;
 wire \atari2600.ram[1][1] ;
 wire \atari2600.ram[1][2] ;
 wire \atari2600.ram[1][3] ;
 wire \atari2600.ram[1][4] ;
 wire \atari2600.ram[1][5] ;
 wire \atari2600.ram[1][6] ;
 wire \atari2600.ram[1][7] ;
 wire \atari2600.ram[20][0] ;
 wire \atari2600.ram[20][1] ;
 wire \atari2600.ram[20][2] ;
 wire \atari2600.ram[20][3] ;
 wire \atari2600.ram[20][4] ;
 wire \atari2600.ram[20][5] ;
 wire \atari2600.ram[20][6] ;
 wire \atari2600.ram[20][7] ;
 wire \atari2600.ram[21][0] ;
 wire \atari2600.ram[21][1] ;
 wire \atari2600.ram[21][2] ;
 wire \atari2600.ram[21][3] ;
 wire \atari2600.ram[21][4] ;
 wire \atari2600.ram[21][5] ;
 wire \atari2600.ram[21][6] ;
 wire \atari2600.ram[21][7] ;
 wire \atari2600.ram[22][0] ;
 wire \atari2600.ram[22][1] ;
 wire \atari2600.ram[22][2] ;
 wire \atari2600.ram[22][3] ;
 wire \atari2600.ram[22][4] ;
 wire \atari2600.ram[22][5] ;
 wire \atari2600.ram[22][6] ;
 wire \atari2600.ram[22][7] ;
 wire \atari2600.ram[23][0] ;
 wire \atari2600.ram[23][1] ;
 wire \atari2600.ram[23][2] ;
 wire \atari2600.ram[23][3] ;
 wire \atari2600.ram[23][4] ;
 wire \atari2600.ram[23][5] ;
 wire \atari2600.ram[23][6] ;
 wire \atari2600.ram[23][7] ;
 wire \atari2600.ram[24][0] ;
 wire \atari2600.ram[24][1] ;
 wire \atari2600.ram[24][2] ;
 wire \atari2600.ram[24][3] ;
 wire \atari2600.ram[24][4] ;
 wire \atari2600.ram[24][5] ;
 wire \atari2600.ram[24][6] ;
 wire \atari2600.ram[24][7] ;
 wire \atari2600.ram[25][0] ;
 wire \atari2600.ram[25][1] ;
 wire \atari2600.ram[25][2] ;
 wire \atari2600.ram[25][3] ;
 wire \atari2600.ram[25][4] ;
 wire \atari2600.ram[25][5] ;
 wire \atari2600.ram[25][6] ;
 wire \atari2600.ram[25][7] ;
 wire \atari2600.ram[26][0] ;
 wire \atari2600.ram[26][1] ;
 wire \atari2600.ram[26][2] ;
 wire \atari2600.ram[26][3] ;
 wire \atari2600.ram[26][4] ;
 wire \atari2600.ram[26][5] ;
 wire \atari2600.ram[26][6] ;
 wire \atari2600.ram[26][7] ;
 wire \atari2600.ram[27][0] ;
 wire \atari2600.ram[27][1] ;
 wire \atari2600.ram[27][2] ;
 wire \atari2600.ram[27][3] ;
 wire \atari2600.ram[27][4] ;
 wire \atari2600.ram[27][5] ;
 wire \atari2600.ram[27][6] ;
 wire \atari2600.ram[27][7] ;
 wire \atari2600.ram[28][0] ;
 wire \atari2600.ram[28][1] ;
 wire \atari2600.ram[28][2] ;
 wire \atari2600.ram[28][3] ;
 wire \atari2600.ram[28][4] ;
 wire \atari2600.ram[28][5] ;
 wire \atari2600.ram[28][6] ;
 wire \atari2600.ram[28][7] ;
 wire \atari2600.ram[29][0] ;
 wire \atari2600.ram[29][1] ;
 wire \atari2600.ram[29][2] ;
 wire \atari2600.ram[29][3] ;
 wire \atari2600.ram[29][4] ;
 wire \atari2600.ram[29][5] ;
 wire \atari2600.ram[29][6] ;
 wire \atari2600.ram[29][7] ;
 wire \atari2600.ram[2][0] ;
 wire \atari2600.ram[2][1] ;
 wire \atari2600.ram[2][2] ;
 wire \atari2600.ram[2][3] ;
 wire \atari2600.ram[2][4] ;
 wire \atari2600.ram[2][5] ;
 wire \atari2600.ram[2][6] ;
 wire \atari2600.ram[2][7] ;
 wire \atari2600.ram[30][0] ;
 wire \atari2600.ram[30][1] ;
 wire \atari2600.ram[30][2] ;
 wire \atari2600.ram[30][3] ;
 wire \atari2600.ram[30][4] ;
 wire \atari2600.ram[30][5] ;
 wire \atari2600.ram[30][6] ;
 wire \atari2600.ram[30][7] ;
 wire \atari2600.ram[31][0] ;
 wire \atari2600.ram[31][1] ;
 wire \atari2600.ram[31][2] ;
 wire \atari2600.ram[31][3] ;
 wire \atari2600.ram[31][4] ;
 wire \atari2600.ram[31][5] ;
 wire \atari2600.ram[31][6] ;
 wire \atari2600.ram[31][7] ;
 wire \atari2600.ram[32][0] ;
 wire \atari2600.ram[32][1] ;
 wire \atari2600.ram[32][2] ;
 wire \atari2600.ram[32][3] ;
 wire \atari2600.ram[32][4] ;
 wire \atari2600.ram[32][5] ;
 wire \atari2600.ram[32][6] ;
 wire \atari2600.ram[32][7] ;
 wire \atari2600.ram[33][0] ;
 wire \atari2600.ram[33][1] ;
 wire \atari2600.ram[33][2] ;
 wire \atari2600.ram[33][3] ;
 wire \atari2600.ram[33][4] ;
 wire \atari2600.ram[33][5] ;
 wire \atari2600.ram[33][6] ;
 wire \atari2600.ram[33][7] ;
 wire \atari2600.ram[34][0] ;
 wire \atari2600.ram[34][1] ;
 wire \atari2600.ram[34][2] ;
 wire \atari2600.ram[34][3] ;
 wire \atari2600.ram[34][4] ;
 wire \atari2600.ram[34][5] ;
 wire \atari2600.ram[34][6] ;
 wire \atari2600.ram[34][7] ;
 wire \atari2600.ram[35][0] ;
 wire \atari2600.ram[35][1] ;
 wire \atari2600.ram[35][2] ;
 wire \atari2600.ram[35][3] ;
 wire \atari2600.ram[35][4] ;
 wire \atari2600.ram[35][5] ;
 wire \atari2600.ram[35][6] ;
 wire \atari2600.ram[35][7] ;
 wire \atari2600.ram[36][0] ;
 wire \atari2600.ram[36][1] ;
 wire \atari2600.ram[36][2] ;
 wire \atari2600.ram[36][3] ;
 wire \atari2600.ram[36][4] ;
 wire \atari2600.ram[36][5] ;
 wire \atari2600.ram[36][6] ;
 wire \atari2600.ram[36][7] ;
 wire \atari2600.ram[37][0] ;
 wire \atari2600.ram[37][1] ;
 wire \atari2600.ram[37][2] ;
 wire \atari2600.ram[37][3] ;
 wire \atari2600.ram[37][4] ;
 wire \atari2600.ram[37][5] ;
 wire \atari2600.ram[37][6] ;
 wire \atari2600.ram[37][7] ;
 wire \atari2600.ram[38][0] ;
 wire \atari2600.ram[38][1] ;
 wire \atari2600.ram[38][2] ;
 wire \atari2600.ram[38][3] ;
 wire \atari2600.ram[38][4] ;
 wire \atari2600.ram[38][5] ;
 wire \atari2600.ram[38][6] ;
 wire \atari2600.ram[38][7] ;
 wire \atari2600.ram[39][0] ;
 wire \atari2600.ram[39][1] ;
 wire \atari2600.ram[39][2] ;
 wire \atari2600.ram[39][3] ;
 wire \atari2600.ram[39][4] ;
 wire \atari2600.ram[39][5] ;
 wire \atari2600.ram[39][6] ;
 wire \atari2600.ram[39][7] ;
 wire \atari2600.ram[3][0] ;
 wire \atari2600.ram[3][1] ;
 wire \atari2600.ram[3][2] ;
 wire \atari2600.ram[3][3] ;
 wire \atari2600.ram[3][4] ;
 wire \atari2600.ram[3][5] ;
 wire \atari2600.ram[3][6] ;
 wire \atari2600.ram[3][7] ;
 wire \atari2600.ram[40][0] ;
 wire \atari2600.ram[40][1] ;
 wire \atari2600.ram[40][2] ;
 wire \atari2600.ram[40][3] ;
 wire \atari2600.ram[40][4] ;
 wire \atari2600.ram[40][5] ;
 wire \atari2600.ram[40][6] ;
 wire \atari2600.ram[40][7] ;
 wire \atari2600.ram[41][0] ;
 wire \atari2600.ram[41][1] ;
 wire \atari2600.ram[41][2] ;
 wire \atari2600.ram[41][3] ;
 wire \atari2600.ram[41][4] ;
 wire \atari2600.ram[41][5] ;
 wire \atari2600.ram[41][6] ;
 wire \atari2600.ram[41][7] ;
 wire \atari2600.ram[42][0] ;
 wire \atari2600.ram[42][1] ;
 wire \atari2600.ram[42][2] ;
 wire \atari2600.ram[42][3] ;
 wire \atari2600.ram[42][4] ;
 wire \atari2600.ram[42][5] ;
 wire \atari2600.ram[42][6] ;
 wire \atari2600.ram[42][7] ;
 wire \atari2600.ram[43][0] ;
 wire \atari2600.ram[43][1] ;
 wire \atari2600.ram[43][2] ;
 wire \atari2600.ram[43][3] ;
 wire \atari2600.ram[43][4] ;
 wire \atari2600.ram[43][5] ;
 wire \atari2600.ram[43][6] ;
 wire \atari2600.ram[43][7] ;
 wire \atari2600.ram[44][0] ;
 wire \atari2600.ram[44][1] ;
 wire \atari2600.ram[44][2] ;
 wire \atari2600.ram[44][3] ;
 wire \atari2600.ram[44][4] ;
 wire \atari2600.ram[44][5] ;
 wire \atari2600.ram[44][6] ;
 wire \atari2600.ram[44][7] ;
 wire \atari2600.ram[45][0] ;
 wire \atari2600.ram[45][1] ;
 wire \atari2600.ram[45][2] ;
 wire \atari2600.ram[45][3] ;
 wire \atari2600.ram[45][4] ;
 wire \atari2600.ram[45][5] ;
 wire \atari2600.ram[45][6] ;
 wire \atari2600.ram[45][7] ;
 wire \atari2600.ram[46][0] ;
 wire \atari2600.ram[46][1] ;
 wire \atari2600.ram[46][2] ;
 wire \atari2600.ram[46][3] ;
 wire \atari2600.ram[46][4] ;
 wire \atari2600.ram[46][5] ;
 wire \atari2600.ram[46][6] ;
 wire \atari2600.ram[46][7] ;
 wire \atari2600.ram[47][0] ;
 wire \atari2600.ram[47][1] ;
 wire \atari2600.ram[47][2] ;
 wire \atari2600.ram[47][3] ;
 wire \atari2600.ram[47][4] ;
 wire \atari2600.ram[47][5] ;
 wire \atari2600.ram[47][6] ;
 wire \atari2600.ram[47][7] ;
 wire \atari2600.ram[48][0] ;
 wire \atari2600.ram[48][1] ;
 wire \atari2600.ram[48][2] ;
 wire \atari2600.ram[48][3] ;
 wire \atari2600.ram[48][4] ;
 wire \atari2600.ram[48][5] ;
 wire \atari2600.ram[48][6] ;
 wire \atari2600.ram[48][7] ;
 wire \atari2600.ram[49][0] ;
 wire \atari2600.ram[49][1] ;
 wire \atari2600.ram[49][2] ;
 wire \atari2600.ram[49][3] ;
 wire \atari2600.ram[49][4] ;
 wire \atari2600.ram[49][5] ;
 wire \atari2600.ram[49][6] ;
 wire \atari2600.ram[49][7] ;
 wire \atari2600.ram[4][0] ;
 wire \atari2600.ram[4][1] ;
 wire \atari2600.ram[4][2] ;
 wire \atari2600.ram[4][3] ;
 wire \atari2600.ram[4][4] ;
 wire \atari2600.ram[4][5] ;
 wire \atari2600.ram[4][6] ;
 wire \atari2600.ram[4][7] ;
 wire \atari2600.ram[50][0] ;
 wire \atari2600.ram[50][1] ;
 wire \atari2600.ram[50][2] ;
 wire \atari2600.ram[50][3] ;
 wire \atari2600.ram[50][4] ;
 wire \atari2600.ram[50][5] ;
 wire \atari2600.ram[50][6] ;
 wire \atari2600.ram[50][7] ;
 wire \atari2600.ram[51][0] ;
 wire \atari2600.ram[51][1] ;
 wire \atari2600.ram[51][2] ;
 wire \atari2600.ram[51][3] ;
 wire \atari2600.ram[51][4] ;
 wire \atari2600.ram[51][5] ;
 wire \atari2600.ram[51][6] ;
 wire \atari2600.ram[51][7] ;
 wire \atari2600.ram[52][0] ;
 wire \atari2600.ram[52][1] ;
 wire \atari2600.ram[52][2] ;
 wire \atari2600.ram[52][3] ;
 wire \atari2600.ram[52][4] ;
 wire \atari2600.ram[52][5] ;
 wire \atari2600.ram[52][6] ;
 wire \atari2600.ram[52][7] ;
 wire \atari2600.ram[53][0] ;
 wire \atari2600.ram[53][1] ;
 wire \atari2600.ram[53][2] ;
 wire \atari2600.ram[53][3] ;
 wire \atari2600.ram[53][4] ;
 wire \atari2600.ram[53][5] ;
 wire \atari2600.ram[53][6] ;
 wire \atari2600.ram[53][7] ;
 wire \atari2600.ram[54][0] ;
 wire \atari2600.ram[54][1] ;
 wire \atari2600.ram[54][2] ;
 wire \atari2600.ram[54][3] ;
 wire \atari2600.ram[54][4] ;
 wire \atari2600.ram[54][5] ;
 wire \atari2600.ram[54][6] ;
 wire \atari2600.ram[54][7] ;
 wire \atari2600.ram[55][0] ;
 wire \atari2600.ram[55][1] ;
 wire \atari2600.ram[55][2] ;
 wire \atari2600.ram[55][3] ;
 wire \atari2600.ram[55][4] ;
 wire \atari2600.ram[55][5] ;
 wire \atari2600.ram[55][6] ;
 wire \atari2600.ram[55][7] ;
 wire \atari2600.ram[56][0] ;
 wire \atari2600.ram[56][1] ;
 wire \atari2600.ram[56][2] ;
 wire \atari2600.ram[56][3] ;
 wire \atari2600.ram[56][4] ;
 wire \atari2600.ram[56][5] ;
 wire \atari2600.ram[56][6] ;
 wire \atari2600.ram[56][7] ;
 wire \atari2600.ram[57][0] ;
 wire \atari2600.ram[57][1] ;
 wire \atari2600.ram[57][2] ;
 wire \atari2600.ram[57][3] ;
 wire \atari2600.ram[57][4] ;
 wire \atari2600.ram[57][5] ;
 wire \atari2600.ram[57][6] ;
 wire \atari2600.ram[57][7] ;
 wire \atari2600.ram[58][0] ;
 wire \atari2600.ram[58][1] ;
 wire \atari2600.ram[58][2] ;
 wire \atari2600.ram[58][3] ;
 wire \atari2600.ram[58][4] ;
 wire \atari2600.ram[58][5] ;
 wire \atari2600.ram[58][6] ;
 wire \atari2600.ram[58][7] ;
 wire \atari2600.ram[59][0] ;
 wire \atari2600.ram[59][1] ;
 wire \atari2600.ram[59][2] ;
 wire \atari2600.ram[59][3] ;
 wire \atari2600.ram[59][4] ;
 wire \atari2600.ram[59][5] ;
 wire \atari2600.ram[59][6] ;
 wire \atari2600.ram[59][7] ;
 wire \atari2600.ram[5][0] ;
 wire \atari2600.ram[5][1] ;
 wire \atari2600.ram[5][2] ;
 wire \atari2600.ram[5][3] ;
 wire \atari2600.ram[5][4] ;
 wire \atari2600.ram[5][5] ;
 wire \atari2600.ram[5][6] ;
 wire \atari2600.ram[5][7] ;
 wire \atari2600.ram[60][0] ;
 wire \atari2600.ram[60][1] ;
 wire \atari2600.ram[60][2] ;
 wire \atari2600.ram[60][3] ;
 wire \atari2600.ram[60][4] ;
 wire \atari2600.ram[60][5] ;
 wire \atari2600.ram[60][6] ;
 wire \atari2600.ram[60][7] ;
 wire \atari2600.ram[61][0] ;
 wire \atari2600.ram[61][1] ;
 wire \atari2600.ram[61][2] ;
 wire \atari2600.ram[61][3] ;
 wire \atari2600.ram[61][4] ;
 wire \atari2600.ram[61][5] ;
 wire \atari2600.ram[61][6] ;
 wire \atari2600.ram[61][7] ;
 wire \atari2600.ram[62][0] ;
 wire \atari2600.ram[62][1] ;
 wire \atari2600.ram[62][2] ;
 wire \atari2600.ram[62][3] ;
 wire \atari2600.ram[62][4] ;
 wire \atari2600.ram[62][5] ;
 wire \atari2600.ram[62][6] ;
 wire \atari2600.ram[62][7] ;
 wire \atari2600.ram[63][0] ;
 wire \atari2600.ram[63][1] ;
 wire \atari2600.ram[63][2] ;
 wire \atari2600.ram[63][3] ;
 wire \atari2600.ram[63][4] ;
 wire \atari2600.ram[63][5] ;
 wire \atari2600.ram[63][6] ;
 wire \atari2600.ram[63][7] ;
 wire \atari2600.ram[64][0] ;
 wire \atari2600.ram[64][1] ;
 wire \atari2600.ram[64][2] ;
 wire \atari2600.ram[64][3] ;
 wire \atari2600.ram[64][4] ;
 wire \atari2600.ram[64][5] ;
 wire \atari2600.ram[64][6] ;
 wire \atari2600.ram[64][7] ;
 wire \atari2600.ram[65][0] ;
 wire \atari2600.ram[65][1] ;
 wire \atari2600.ram[65][2] ;
 wire \atari2600.ram[65][3] ;
 wire \atari2600.ram[65][4] ;
 wire \atari2600.ram[65][5] ;
 wire \atari2600.ram[65][6] ;
 wire \atari2600.ram[65][7] ;
 wire \atari2600.ram[66][0] ;
 wire \atari2600.ram[66][1] ;
 wire \atari2600.ram[66][2] ;
 wire \atari2600.ram[66][3] ;
 wire \atari2600.ram[66][4] ;
 wire \atari2600.ram[66][5] ;
 wire \atari2600.ram[66][6] ;
 wire \atari2600.ram[66][7] ;
 wire \atari2600.ram[67][0] ;
 wire \atari2600.ram[67][1] ;
 wire \atari2600.ram[67][2] ;
 wire \atari2600.ram[67][3] ;
 wire \atari2600.ram[67][4] ;
 wire \atari2600.ram[67][5] ;
 wire \atari2600.ram[67][6] ;
 wire \atari2600.ram[67][7] ;
 wire \atari2600.ram[68][0] ;
 wire \atari2600.ram[68][1] ;
 wire \atari2600.ram[68][2] ;
 wire \atari2600.ram[68][3] ;
 wire \atari2600.ram[68][4] ;
 wire \atari2600.ram[68][5] ;
 wire \atari2600.ram[68][6] ;
 wire \atari2600.ram[68][7] ;
 wire \atari2600.ram[69][0] ;
 wire \atari2600.ram[69][1] ;
 wire \atari2600.ram[69][2] ;
 wire \atari2600.ram[69][3] ;
 wire \atari2600.ram[69][4] ;
 wire \atari2600.ram[69][5] ;
 wire \atari2600.ram[69][6] ;
 wire \atari2600.ram[69][7] ;
 wire \atari2600.ram[6][0] ;
 wire \atari2600.ram[6][1] ;
 wire \atari2600.ram[6][2] ;
 wire \atari2600.ram[6][3] ;
 wire \atari2600.ram[6][4] ;
 wire \atari2600.ram[6][5] ;
 wire \atari2600.ram[6][6] ;
 wire \atari2600.ram[6][7] ;
 wire \atari2600.ram[70][0] ;
 wire \atari2600.ram[70][1] ;
 wire \atari2600.ram[70][2] ;
 wire \atari2600.ram[70][3] ;
 wire \atari2600.ram[70][4] ;
 wire \atari2600.ram[70][5] ;
 wire \atari2600.ram[70][6] ;
 wire \atari2600.ram[70][7] ;
 wire \atari2600.ram[71][0] ;
 wire \atari2600.ram[71][1] ;
 wire \atari2600.ram[71][2] ;
 wire \atari2600.ram[71][3] ;
 wire \atari2600.ram[71][4] ;
 wire \atari2600.ram[71][5] ;
 wire \atari2600.ram[71][6] ;
 wire \atari2600.ram[71][7] ;
 wire \atari2600.ram[72][0] ;
 wire \atari2600.ram[72][1] ;
 wire \atari2600.ram[72][2] ;
 wire \atari2600.ram[72][3] ;
 wire \atari2600.ram[72][4] ;
 wire \atari2600.ram[72][5] ;
 wire \atari2600.ram[72][6] ;
 wire \atari2600.ram[72][7] ;
 wire \atari2600.ram[73][0] ;
 wire \atari2600.ram[73][1] ;
 wire \atari2600.ram[73][2] ;
 wire \atari2600.ram[73][3] ;
 wire \atari2600.ram[73][4] ;
 wire \atari2600.ram[73][5] ;
 wire \atari2600.ram[73][6] ;
 wire \atari2600.ram[73][7] ;
 wire \atari2600.ram[74][0] ;
 wire \atari2600.ram[74][1] ;
 wire \atari2600.ram[74][2] ;
 wire \atari2600.ram[74][3] ;
 wire \atari2600.ram[74][4] ;
 wire \atari2600.ram[74][5] ;
 wire \atari2600.ram[74][6] ;
 wire \atari2600.ram[74][7] ;
 wire \atari2600.ram[75][0] ;
 wire \atari2600.ram[75][1] ;
 wire \atari2600.ram[75][2] ;
 wire \atari2600.ram[75][3] ;
 wire \atari2600.ram[75][4] ;
 wire \atari2600.ram[75][5] ;
 wire \atari2600.ram[75][6] ;
 wire \atari2600.ram[75][7] ;
 wire \atari2600.ram[76][0] ;
 wire \atari2600.ram[76][1] ;
 wire \atari2600.ram[76][2] ;
 wire \atari2600.ram[76][3] ;
 wire \atari2600.ram[76][4] ;
 wire \atari2600.ram[76][5] ;
 wire \atari2600.ram[76][6] ;
 wire \atari2600.ram[76][7] ;
 wire \atari2600.ram[77][0] ;
 wire \atari2600.ram[77][1] ;
 wire \atari2600.ram[77][2] ;
 wire \atari2600.ram[77][3] ;
 wire \atari2600.ram[77][4] ;
 wire \atari2600.ram[77][5] ;
 wire \atari2600.ram[77][6] ;
 wire \atari2600.ram[77][7] ;
 wire \atari2600.ram[78][0] ;
 wire \atari2600.ram[78][1] ;
 wire \atari2600.ram[78][2] ;
 wire \atari2600.ram[78][3] ;
 wire \atari2600.ram[78][4] ;
 wire \atari2600.ram[78][5] ;
 wire \atari2600.ram[78][6] ;
 wire \atari2600.ram[78][7] ;
 wire \atari2600.ram[79][0] ;
 wire \atari2600.ram[79][1] ;
 wire \atari2600.ram[79][2] ;
 wire \atari2600.ram[79][3] ;
 wire \atari2600.ram[79][4] ;
 wire \atari2600.ram[79][5] ;
 wire \atari2600.ram[79][6] ;
 wire \atari2600.ram[79][7] ;
 wire \atari2600.ram[7][0] ;
 wire \atari2600.ram[7][1] ;
 wire \atari2600.ram[7][2] ;
 wire \atari2600.ram[7][3] ;
 wire \atari2600.ram[7][4] ;
 wire \atari2600.ram[7][5] ;
 wire \atari2600.ram[7][6] ;
 wire \atari2600.ram[7][7] ;
 wire \atari2600.ram[80][0] ;
 wire \atari2600.ram[80][1] ;
 wire \atari2600.ram[80][2] ;
 wire \atari2600.ram[80][3] ;
 wire \atari2600.ram[80][4] ;
 wire \atari2600.ram[80][5] ;
 wire \atari2600.ram[80][6] ;
 wire \atari2600.ram[80][7] ;
 wire \atari2600.ram[81][0] ;
 wire \atari2600.ram[81][1] ;
 wire \atari2600.ram[81][2] ;
 wire \atari2600.ram[81][3] ;
 wire \atari2600.ram[81][4] ;
 wire \atari2600.ram[81][5] ;
 wire \atari2600.ram[81][6] ;
 wire \atari2600.ram[81][7] ;
 wire \atari2600.ram[82][0] ;
 wire \atari2600.ram[82][1] ;
 wire \atari2600.ram[82][2] ;
 wire \atari2600.ram[82][3] ;
 wire \atari2600.ram[82][4] ;
 wire \atari2600.ram[82][5] ;
 wire \atari2600.ram[82][6] ;
 wire \atari2600.ram[82][7] ;
 wire \atari2600.ram[83][0] ;
 wire \atari2600.ram[83][1] ;
 wire \atari2600.ram[83][2] ;
 wire \atari2600.ram[83][3] ;
 wire \atari2600.ram[83][4] ;
 wire \atari2600.ram[83][5] ;
 wire \atari2600.ram[83][6] ;
 wire \atari2600.ram[83][7] ;
 wire \atari2600.ram[84][0] ;
 wire \atari2600.ram[84][1] ;
 wire \atari2600.ram[84][2] ;
 wire \atari2600.ram[84][3] ;
 wire \atari2600.ram[84][4] ;
 wire \atari2600.ram[84][5] ;
 wire \atari2600.ram[84][6] ;
 wire \atari2600.ram[84][7] ;
 wire \atari2600.ram[85][0] ;
 wire \atari2600.ram[85][1] ;
 wire \atari2600.ram[85][2] ;
 wire \atari2600.ram[85][3] ;
 wire \atari2600.ram[85][4] ;
 wire \atari2600.ram[85][5] ;
 wire \atari2600.ram[85][6] ;
 wire \atari2600.ram[85][7] ;
 wire \atari2600.ram[86][0] ;
 wire \atari2600.ram[86][1] ;
 wire \atari2600.ram[86][2] ;
 wire \atari2600.ram[86][3] ;
 wire \atari2600.ram[86][4] ;
 wire \atari2600.ram[86][5] ;
 wire \atari2600.ram[86][6] ;
 wire \atari2600.ram[86][7] ;
 wire \atari2600.ram[87][0] ;
 wire \atari2600.ram[87][1] ;
 wire \atari2600.ram[87][2] ;
 wire \atari2600.ram[87][3] ;
 wire \atari2600.ram[87][4] ;
 wire \atari2600.ram[87][5] ;
 wire \atari2600.ram[87][6] ;
 wire \atari2600.ram[87][7] ;
 wire \atari2600.ram[88][0] ;
 wire \atari2600.ram[88][1] ;
 wire \atari2600.ram[88][2] ;
 wire \atari2600.ram[88][3] ;
 wire \atari2600.ram[88][4] ;
 wire \atari2600.ram[88][5] ;
 wire \atari2600.ram[88][6] ;
 wire \atari2600.ram[88][7] ;
 wire \atari2600.ram[89][0] ;
 wire \atari2600.ram[89][1] ;
 wire \atari2600.ram[89][2] ;
 wire \atari2600.ram[89][3] ;
 wire \atari2600.ram[89][4] ;
 wire \atari2600.ram[89][5] ;
 wire \atari2600.ram[89][6] ;
 wire \atari2600.ram[89][7] ;
 wire \atari2600.ram[8][0] ;
 wire \atari2600.ram[8][1] ;
 wire \atari2600.ram[8][2] ;
 wire \atari2600.ram[8][3] ;
 wire \atari2600.ram[8][4] ;
 wire \atari2600.ram[8][5] ;
 wire \atari2600.ram[8][6] ;
 wire \atari2600.ram[8][7] ;
 wire \atari2600.ram[90][0] ;
 wire \atari2600.ram[90][1] ;
 wire \atari2600.ram[90][2] ;
 wire \atari2600.ram[90][3] ;
 wire \atari2600.ram[90][4] ;
 wire \atari2600.ram[90][5] ;
 wire \atari2600.ram[90][6] ;
 wire \atari2600.ram[90][7] ;
 wire \atari2600.ram[91][0] ;
 wire \atari2600.ram[91][1] ;
 wire \atari2600.ram[91][2] ;
 wire \atari2600.ram[91][3] ;
 wire \atari2600.ram[91][4] ;
 wire \atari2600.ram[91][5] ;
 wire \atari2600.ram[91][6] ;
 wire \atari2600.ram[91][7] ;
 wire \atari2600.ram[92][0] ;
 wire \atari2600.ram[92][1] ;
 wire \atari2600.ram[92][2] ;
 wire \atari2600.ram[92][3] ;
 wire \atari2600.ram[92][4] ;
 wire \atari2600.ram[92][5] ;
 wire \atari2600.ram[92][6] ;
 wire \atari2600.ram[92][7] ;
 wire \atari2600.ram[93][0] ;
 wire \atari2600.ram[93][1] ;
 wire \atari2600.ram[93][2] ;
 wire \atari2600.ram[93][3] ;
 wire \atari2600.ram[93][4] ;
 wire \atari2600.ram[93][5] ;
 wire \atari2600.ram[93][6] ;
 wire \atari2600.ram[93][7] ;
 wire \atari2600.ram[94][0] ;
 wire \atari2600.ram[94][1] ;
 wire \atari2600.ram[94][2] ;
 wire \atari2600.ram[94][3] ;
 wire \atari2600.ram[94][4] ;
 wire \atari2600.ram[94][5] ;
 wire \atari2600.ram[94][6] ;
 wire \atari2600.ram[94][7] ;
 wire \atari2600.ram[95][0] ;
 wire \atari2600.ram[95][1] ;
 wire \atari2600.ram[95][2] ;
 wire \atari2600.ram[95][3] ;
 wire \atari2600.ram[95][4] ;
 wire \atari2600.ram[95][5] ;
 wire \atari2600.ram[95][6] ;
 wire \atari2600.ram[95][7] ;
 wire \atari2600.ram[96][0] ;
 wire \atari2600.ram[96][1] ;
 wire \atari2600.ram[96][2] ;
 wire \atari2600.ram[96][3] ;
 wire \atari2600.ram[96][4] ;
 wire \atari2600.ram[96][5] ;
 wire \atari2600.ram[96][6] ;
 wire \atari2600.ram[96][7] ;
 wire \atari2600.ram[97][0] ;
 wire \atari2600.ram[97][1] ;
 wire \atari2600.ram[97][2] ;
 wire \atari2600.ram[97][3] ;
 wire \atari2600.ram[97][4] ;
 wire \atari2600.ram[97][5] ;
 wire \atari2600.ram[97][6] ;
 wire \atari2600.ram[97][7] ;
 wire \atari2600.ram[98][0] ;
 wire \atari2600.ram[98][1] ;
 wire \atari2600.ram[98][2] ;
 wire \atari2600.ram[98][3] ;
 wire \atari2600.ram[98][4] ;
 wire \atari2600.ram[98][5] ;
 wire \atari2600.ram[98][6] ;
 wire \atari2600.ram[98][7] ;
 wire \atari2600.ram[99][0] ;
 wire \atari2600.ram[99][1] ;
 wire \atari2600.ram[99][2] ;
 wire \atari2600.ram[99][3] ;
 wire \atari2600.ram[99][4] ;
 wire \atari2600.ram[99][5] ;
 wire \atari2600.ram[99][6] ;
 wire \atari2600.ram[99][7] ;
 wire \atari2600.ram[9][0] ;
 wire \atari2600.ram[9][1] ;
 wire \atari2600.ram[9][2] ;
 wire \atari2600.ram[9][3] ;
 wire \atari2600.ram[9][4] ;
 wire \atari2600.ram[9][5] ;
 wire \atari2600.ram[9][6] ;
 wire \atari2600.ram[9][7] ;
 wire \atari2600.ram_data[0] ;
 wire \atari2600.ram_data[1] ;
 wire \atari2600.ram_data[2] ;
 wire \atari2600.ram_data[3] ;
 wire \atari2600.ram_data[4] ;
 wire \atari2600.ram_data[5] ;
 wire \atari2600.ram_data[6] ;
 wire \atari2600.ram_data[7] ;
 wire \atari2600.rom_data[0] ;
 wire \atari2600.rom_data[1] ;
 wire \atari2600.rom_data[2] ;
 wire \atari2600.rom_data[3] ;
 wire \atari2600.rom_data[4] ;
 wire \atari2600.rom_data[5] ;
 wire \atari2600.rom_data[6] ;
 wire \atari2600.rom_data[7] ;
 wire \atari2600.stall_cpu ;
 wire \atari2600.tia.audc0[0] ;
 wire \atari2600.tia.audc0[1] ;
 wire \atari2600.tia.audc0[2] ;
 wire \atari2600.tia.audc0[3] ;
 wire \atari2600.tia.audc1[0] ;
 wire \atari2600.tia.audc1[1] ;
 wire \atari2600.tia.audc1[2] ;
 wire \atari2600.tia.audc1[3] ;
 wire \atari2600.tia.audf0[0] ;
 wire \atari2600.tia.audf0[1] ;
 wire \atari2600.tia.audf0[2] ;
 wire \atari2600.tia.audf0[3] ;
 wire \atari2600.tia.audf0[4] ;
 wire \atari2600.tia.audf1[0] ;
 wire \atari2600.tia.audf1[1] ;
 wire \atari2600.tia.audf1[2] ;
 wire \atari2600.tia.audf1[3] ;
 wire \atari2600.tia.audf1[4] ;
 wire \atari2600.tia.audio_l ;
 wire \atari2600.tia.audio_left_counter[0] ;
 wire \atari2600.tia.audio_left_counter[10] ;
 wire \atari2600.tia.audio_left_counter[11] ;
 wire \atari2600.tia.audio_left_counter[12] ;
 wire \atari2600.tia.audio_left_counter[13] ;
 wire \atari2600.tia.audio_left_counter[14] ;
 wire \atari2600.tia.audio_left_counter[15] ;
 wire \atari2600.tia.audio_left_counter[1] ;
 wire \atari2600.tia.audio_left_counter[2] ;
 wire \atari2600.tia.audio_left_counter[3] ;
 wire \atari2600.tia.audio_left_counter[4] ;
 wire \atari2600.tia.audio_left_counter[5] ;
 wire \atari2600.tia.audio_left_counter[6] ;
 wire \atari2600.tia.audio_left_counter[7] ;
 wire \atari2600.tia.audio_left_counter[8] ;
 wire \atari2600.tia.audio_left_counter[9] ;
 wire \atari2600.tia.audio_r ;
 wire \atari2600.tia.audio_right_counter[0] ;
 wire \atari2600.tia.audio_right_counter[10] ;
 wire \atari2600.tia.audio_right_counter[11] ;
 wire \atari2600.tia.audio_right_counter[12] ;
 wire \atari2600.tia.audio_right_counter[13] ;
 wire \atari2600.tia.audio_right_counter[14] ;
 wire \atari2600.tia.audio_right_counter[15] ;
 wire \atari2600.tia.audio_right_counter[1] ;
 wire \atari2600.tia.audio_right_counter[2] ;
 wire \atari2600.tia.audio_right_counter[3] ;
 wire \atari2600.tia.audio_right_counter[4] ;
 wire \atari2600.tia.audio_right_counter[5] ;
 wire \atari2600.tia.audio_right_counter[6] ;
 wire \atari2600.tia.audio_right_counter[7] ;
 wire \atari2600.tia.audio_right_counter[8] ;
 wire \atari2600.tia.audio_right_counter[9] ;
 wire \atari2600.tia.audv0[0] ;
 wire \atari2600.tia.audv0[1] ;
 wire \atari2600.tia.audv0[2] ;
 wire \atari2600.tia.audv0[3] ;
 wire \atari2600.tia.audv1[0] ;
 wire \atari2600.tia.audv1[1] ;
 wire \atari2600.tia.audv1[2] ;
 wire \atari2600.tia.audv1[3] ;
 wire \atari2600.tia.ball_w[0] ;
 wire \atari2600.tia.ball_w[1] ;
 wire \atari2600.tia.ball_w[2] ;
 wire \atari2600.tia.ball_w[3] ;
 wire \atari2600.tia.colubk[0] ;
 wire \atari2600.tia.colubk[1] ;
 wire \atari2600.tia.colubk[2] ;
 wire \atari2600.tia.colubk[3] ;
 wire \atari2600.tia.colubk[4] ;
 wire \atari2600.tia.colubk[5] ;
 wire \atari2600.tia.colubk[6] ;
 wire \atari2600.tia.colup0[0] ;
 wire \atari2600.tia.colup0[1] ;
 wire \atari2600.tia.colup0[2] ;
 wire \atari2600.tia.colup0[3] ;
 wire \atari2600.tia.colup0[4] ;
 wire \atari2600.tia.colup0[5] ;
 wire \atari2600.tia.colup0[6] ;
 wire \atari2600.tia.colup1[0] ;
 wire \atari2600.tia.colup1[1] ;
 wire \atari2600.tia.colup1[2] ;
 wire \atari2600.tia.colup1[3] ;
 wire \atari2600.tia.colup1[4] ;
 wire \atari2600.tia.colup1[5] ;
 wire \atari2600.tia.colup1[6] ;
 wire \atari2600.tia.colupf[0] ;
 wire \atari2600.tia.colupf[1] ;
 wire \atari2600.tia.colupf[2] ;
 wire \atari2600.tia.colupf[3] ;
 wire \atari2600.tia.colupf[4] ;
 wire \atari2600.tia.colupf[5] ;
 wire \atari2600.tia.colupf[6] ;
 wire \atari2600.tia.cx[0] ;
 wire \atari2600.tia.cx[10] ;
 wire \atari2600.tia.cx[11] ;
 wire \atari2600.tia.cx[12] ;
 wire \atari2600.tia.cx[13] ;
 wire \atari2600.tia.cx[14] ;
 wire \atari2600.tia.cx[1] ;
 wire \atari2600.tia.cx[2] ;
 wire \atari2600.tia.cx[3] ;
 wire \atari2600.tia.cx[4] ;
 wire \atari2600.tia.cx[5] ;
 wire \atari2600.tia.cx[6] ;
 wire \atari2600.tia.cx[7] ;
 wire \atari2600.tia.cx[8] ;
 wire \atari2600.tia.cx[9] ;
 wire \atari2600.tia.cx_clr ;
 wire \atari2600.tia.dat_o[6] ;
 wire \atari2600.tia.dat_o[7] ;
 wire \atari2600.tia.diag[100] ;
 wire \atari2600.tia.diag[101] ;
 wire \atari2600.tia.diag[102] ;
 wire \atari2600.tia.diag[103] ;
 wire \atari2600.tia.diag[104] ;
 wire \atari2600.tia.diag[105] ;
 wire \atari2600.tia.diag[106] ;
 wire \atari2600.tia.diag[107] ;
 wire \atari2600.tia.diag[108] ;
 wire \atari2600.tia.diag[109] ;
 wire \atari2600.tia.diag[110] ;
 wire \atari2600.tia.diag[111] ;
 wire \atari2600.tia.diag[32] ;
 wire \atari2600.tia.diag[33] ;
 wire \atari2600.tia.diag[34] ;
 wire \atari2600.tia.diag[35] ;
 wire \atari2600.tia.diag[36] ;
 wire \atari2600.tia.diag[37] ;
 wire \atari2600.tia.diag[38] ;
 wire \atari2600.tia.diag[39] ;
 wire \atari2600.tia.diag[40] ;
 wire \atari2600.tia.diag[41] ;
 wire \atari2600.tia.diag[42] ;
 wire \atari2600.tia.diag[43] ;
 wire \atari2600.tia.diag[44] ;
 wire \atari2600.tia.diag[45] ;
 wire \atari2600.tia.diag[46] ;
 wire \atari2600.tia.diag[47] ;
 wire \atari2600.tia.diag[48] ;
 wire \atari2600.tia.diag[49] ;
 wire \atari2600.tia.diag[50] ;
 wire \atari2600.tia.diag[51] ;
 wire \atari2600.tia.diag[52] ;
 wire \atari2600.tia.diag[53] ;
 wire \atari2600.tia.diag[54] ;
 wire \atari2600.tia.diag[55] ;
 wire \atari2600.tia.diag[56] ;
 wire \atari2600.tia.diag[57] ;
 wire \atari2600.tia.diag[58] ;
 wire \atari2600.tia.diag[59] ;
 wire \atari2600.tia.diag[60] ;
 wire \atari2600.tia.diag[61] ;
 wire \atari2600.tia.diag[62] ;
 wire \atari2600.tia.diag[63] ;
 wire \atari2600.tia.diag[64] ;
 wire \atari2600.tia.diag[65] ;
 wire \atari2600.tia.diag[66] ;
 wire \atari2600.tia.diag[67] ;
 wire \atari2600.tia.diag[68] ;
 wire \atari2600.tia.diag[69] ;
 wire \atari2600.tia.diag[70] ;
 wire \atari2600.tia.diag[71] ;
 wire \atari2600.tia.diag[76] ;
 wire \atari2600.tia.diag[77] ;
 wire \atari2600.tia.diag[78] ;
 wire \atari2600.tia.diag[79] ;
 wire \atari2600.tia.diag[80] ;
 wire \atari2600.tia.diag[81] ;
 wire \atari2600.tia.diag[82] ;
 wire \atari2600.tia.diag[83] ;
 wire \atari2600.tia.diag[84] ;
 wire \atari2600.tia.diag[85] ;
 wire \atari2600.tia.diag[86] ;
 wire \atari2600.tia.diag[87] ;
 wire \atari2600.tia.diag[88] ;
 wire \atari2600.tia.diag[89] ;
 wire \atari2600.tia.diag[90] ;
 wire \atari2600.tia.diag[91] ;
 wire \atari2600.tia.diag[92] ;
 wire \atari2600.tia.diag[93] ;
 wire \atari2600.tia.diag[94] ;
 wire \atari2600.tia.diag[95] ;
 wire \atari2600.tia.diag[96] ;
 wire \atari2600.tia.diag[97] ;
 wire \atari2600.tia.diag[98] ;
 wire \atari2600.tia.diag[99] ;
 wire \atari2600.tia.enabl ;
 wire \atari2600.tia.enam0 ;
 wire \atari2600.tia.enam1 ;
 wire \atari2600.tia.hmbl[0] ;
 wire \atari2600.tia.hmbl[1] ;
 wire \atari2600.tia.hmbl[2] ;
 wire \atari2600.tia.hmbl[3] ;
 wire \atari2600.tia.hmm0[0] ;
 wire \atari2600.tia.hmm0[1] ;
 wire \atari2600.tia.hmm0[2] ;
 wire \atari2600.tia.hmm0[3] ;
 wire \atari2600.tia.hmm1[0] ;
 wire \atari2600.tia.hmm1[1] ;
 wire \atari2600.tia.hmm1[2] ;
 wire \atari2600.tia.hmm1[3] ;
 wire \atari2600.tia.hmp0[0] ;
 wire \atari2600.tia.hmp0[1] ;
 wire \atari2600.tia.hmp0[2] ;
 wire \atari2600.tia.hmp0[3] ;
 wire \atari2600.tia.hmp1[0] ;
 wire \atari2600.tia.hmp1[1] ;
 wire \atari2600.tia.hmp1[2] ;
 wire \atari2600.tia.hmp1[3] ;
 wire \atari2600.tia.m0_w[0] ;
 wire \atari2600.tia.m0_w[1] ;
 wire \atari2600.tia.m0_w[2] ;
 wire \atari2600.tia.m0_w[3] ;
 wire \atari2600.tia.m1_w[0] ;
 wire \atari2600.tia.m1_w[1] ;
 wire \atari2600.tia.m1_w[2] ;
 wire \atari2600.tia.m1_w[3] ;
 wire \atari2600.tia.old_grp0[0] ;
 wire \atari2600.tia.old_grp0[1] ;
 wire \atari2600.tia.old_grp0[2] ;
 wire \atari2600.tia.old_grp0[3] ;
 wire \atari2600.tia.old_grp0[4] ;
 wire \atari2600.tia.old_grp0[5] ;
 wire \atari2600.tia.old_grp0[6] ;
 wire \atari2600.tia.old_grp0[7] ;
 wire \atari2600.tia.old_grp1[0] ;
 wire \atari2600.tia.old_grp1[1] ;
 wire \atari2600.tia.old_grp1[2] ;
 wire \atari2600.tia.old_grp1[3] ;
 wire \atari2600.tia.old_grp1[4] ;
 wire \atari2600.tia.old_grp1[5] ;
 wire \atari2600.tia.old_grp1[6] ;
 wire \atari2600.tia.old_grp1[7] ;
 wire \atari2600.tia.p0_copies[1] ;
 wire \atari2600.tia.p0_copies[2] ;
 wire \atari2600.tia.p0_scale[0] ;
 wire \atari2600.tia.p0_scale[1] ;
 wire \atari2600.tia.p0_spacing[4] ;
 wire \atari2600.tia.p0_spacing[5] ;
 wire \atari2600.tia.p0_spacing[6] ;
 wire \atari2600.tia.p0_w[3] ;
 wire \atari2600.tia.p0_w[4] ;
 wire \atari2600.tia.p0_w[5] ;
 wire \atari2600.tia.p1_copies[1] ;
 wire \atari2600.tia.p1_copies[2] ;
 wire \atari2600.tia.p1_scale[0] ;
 wire \atari2600.tia.p1_scale[1] ;
 wire \atari2600.tia.p1_spacing[4] ;
 wire \atari2600.tia.p1_spacing[5] ;
 wire \atari2600.tia.p1_spacing[6] ;
 wire \atari2600.tia.p1_w[3] ;
 wire \atari2600.tia.p1_w[4] ;
 wire \atari2600.tia.p1_w[5] ;
 wire \atari2600.tia.p4_l ;
 wire \atari2600.tia.p4_r ;
 wire \atari2600.tia.p5_l ;
 wire \atari2600.tia.p5_r ;
 wire \atari2600.tia.p9_l ;
 wire \atari2600.tia.p9_r ;
 wire \atari2600.tia.pf_priority ;
 wire \atari2600.tia.poly4_l.x[1] ;
 wire \atari2600.tia.poly4_l.x[2] ;
 wire \atari2600.tia.poly4_l.x[3] ;
 wire \atari2600.tia.poly4_r.x[1] ;
 wire \atari2600.tia.poly4_r.x[2] ;
 wire \atari2600.tia.poly4_r.x[3] ;
 wire \atari2600.tia.poly5_l.x[1] ;
 wire \atari2600.tia.poly5_l.x[2] ;
 wire \atari2600.tia.poly5_l.x[3] ;
 wire \atari2600.tia.poly5_l.x[4] ;
 wire \atari2600.tia.poly5_r.x[1] ;
 wire \atari2600.tia.poly5_r.x[2] ;
 wire \atari2600.tia.poly5_r.x[3] ;
 wire \atari2600.tia.poly5_r.x[4] ;
 wire \atari2600.tia.poly9_l.x[1] ;
 wire \atari2600.tia.poly9_l.x[2] ;
 wire \atari2600.tia.poly9_l.x[3] ;
 wire \atari2600.tia.poly9_l.x[4] ;
 wire \atari2600.tia.poly9_l.x[5] ;
 wire \atari2600.tia.poly9_l.x[6] ;
 wire \atari2600.tia.poly9_l.x[7] ;
 wire \atari2600.tia.poly9_l.x[8] ;
 wire \atari2600.tia.poly9_r.x[1] ;
 wire \atari2600.tia.poly9_r.x[2] ;
 wire \atari2600.tia.poly9_r.x[3] ;
 wire \atari2600.tia.poly9_r.x[4] ;
 wire \atari2600.tia.poly9_r.x[5] ;
 wire \atari2600.tia.poly9_r.x[6] ;
 wire \atari2600.tia.poly9_r.x[7] ;
 wire \atari2600.tia.poly9_r.x[8] ;
 wire \atari2600.tia.refp0 ;
 wire \atari2600.tia.refp1 ;
 wire \atari2600.tia.refpf ;
 wire \atari2600.tia.scorepf ;
 wire \atari2600.tia.vblank ;
 wire \atari2600.tia.vdelp0 ;
 wire \atari2600.tia.vdelp1 ;
 wire \atari2600.tia.vid_out[0] ;
 wire \atari2600.tia.vid_out[1] ;
 wire \atari2600.tia.vid_out[2] ;
 wire \atari2600.tia.vid_out[3] ;
 wire \atari2600.tia.vid_out[4] ;
 wire \atari2600.tia.vid_out[5] ;
 wire \atari2600.tia.vid_out[6] ;
 wire \atari2600.tia.vid_vsync ;
 wire \atari2600.tia.vid_xpos[0] ;
 wire \atari2600.tia.vid_xpos[1] ;
 wire \atari2600.tia.vid_xpos[2] ;
 wire \atari2600.tia.vid_xpos[3] ;
 wire \atari2600.tia.vid_xpos[4] ;
 wire \atari2600.tia.vid_xpos[5] ;
 wire \atari2600.tia.vid_xpos[6] ;
 wire \atari2600.tia.vid_xpos[7] ;
 wire \atari2600.tia.vid_ypos[0] ;
 wire \atari2600.tia.vid_ypos[1] ;
 wire \atari2600.tia.vid_ypos[2] ;
 wire \atari2600.tia.vid_ypos[3] ;
 wire \atari2600.tia.vid_ypos[4] ;
 wire \atari2600.tia.vid_ypos[5] ;
 wire \atari2600.tia.vid_ypos[6] ;
 wire \atari2600.tia.vid_ypos[7] ;
 wire \atari2600.tia.vid_ypos[8] ;
 wire audio_pwm;
 wire \audio_pwm_accumulator[0] ;
 wire \audio_pwm_accumulator[1] ;
 wire \audio_pwm_accumulator[2] ;
 wire \audio_pwm_accumulator[3] ;
 wire \audio_pwm_accumulator[4] ;
 wire \b_pwm_even[1] ;
 wire \b_pwm_even[2] ;
 wire \b_pwm_even[3] ;
 wire \b_pwm_even[4] ;
 wire \b_pwm_even[5] ;
 wire \b_pwm_even[6] ;
 wire \b_pwm_even[7] ;
 wire \b_pwm_even[8] ;
 wire \b_pwm_even[9] ;
 wire \b_pwm_odd[1] ;
 wire \b_pwm_odd[2] ;
 wire \b_pwm_odd[3] ;
 wire \b_pwm_odd[4] ;
 wire \b_pwm_odd[5] ;
 wire \b_pwm_odd[6] ;
 wire \b_pwm_odd[7] ;
 wire \b_pwm_odd[8] ;
 wire \b_pwm_odd[9] ;
 wire \flash_rom.addr[0] ;
 wire \flash_rom.addr[10] ;
 wire \flash_rom.addr[11] ;
 wire \flash_rom.addr[12] ;
 wire \flash_rom.addr[13] ;
 wire \flash_rom.addr[14] ;
 wire \flash_rom.addr[15] ;
 wire \flash_rom.addr[16] ;
 wire \flash_rom.addr[17] ;
 wire \flash_rom.addr[18] ;
 wire \flash_rom.addr[19] ;
 wire \flash_rom.addr[1] ;
 wire \flash_rom.addr[20] ;
 wire \flash_rom.addr[21] ;
 wire \flash_rom.addr[22] ;
 wire \flash_rom.addr[23] ;
 wire \flash_rom.addr[2] ;
 wire \flash_rom.addr[3] ;
 wire \flash_rom.addr[4] ;
 wire \flash_rom.addr[5] ;
 wire \flash_rom.addr[6] ;
 wire \flash_rom.addr[7] ;
 wire \flash_rom.addr[8] ;
 wire \flash_rom.addr[9] ;
 wire \flash_rom.data_ready ;
 wire \flash_rom.fsm_state[0] ;
 wire \flash_rom.fsm_state[1] ;
 wire \flash_rom.fsm_state[2] ;
 wire \flash_rom.nibbles_remaining[0] ;
 wire \flash_rom.nibbles_remaining[1] ;
 wire \flash_rom.nibbles_remaining[2] ;
 wire \flash_rom.spi_clk_out ;
 wire \flash_rom.spi_select ;
 wire \flash_rom.stall_read ;
 wire \frame_counter[0] ;
 wire \frame_counter[1] ;
 wire \frame_counter[2] ;
 wire \g_pwm_even[1] ;
 wire \g_pwm_even[2] ;
 wire \g_pwm_even[3] ;
 wire \g_pwm_even[4] ;
 wire \g_pwm_even[5] ;
 wire \g_pwm_even[6] ;
 wire \g_pwm_even[7] ;
 wire \g_pwm_even[8] ;
 wire \g_pwm_even[9] ;
 wire \g_pwm_odd[1] ;
 wire \g_pwm_odd[2] ;
 wire \g_pwm_odd[3] ;
 wire \g_pwm_odd[4] ;
 wire \g_pwm_odd[5] ;
 wire \g_pwm_odd[6] ;
 wire \g_pwm_odd[7] ;
 wire \g_pwm_odd[8] ;
 wire \g_pwm_odd[9] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vga.vpos[0] ;
 wire \hvsync_gen.vga.vpos[1] ;
 wire \hvsync_gen.vga.vpos[2] ;
 wire \hvsync_gen.vga.vpos[3] ;
 wire \hvsync_gen.vga.vpos[4] ;
 wire \hvsync_gen.vga.vpos[5] ;
 wire \hvsync_gen.vga.vpos[6] ;
 wire \hvsync_gen.vga.vpos[7] ;
 wire \hvsync_gen.vga.vpos[8] ;
 wire \hvsync_gen.vga.vpos[9] ;
 wire \hvsync_gen.vga.vsync ;
 wire \joypmod[2] ;
 wire \r_pwm_even[1] ;
 wire \r_pwm_even[2] ;
 wire \r_pwm_even[3] ;
 wire \r_pwm_even[4] ;
 wire \r_pwm_even[5] ;
 wire \r_pwm_even[6] ;
 wire \r_pwm_even[7] ;
 wire \r_pwm_even[8] ;
 wire \r_pwm_even[9] ;
 wire \r_pwm_odd[1] ;
 wire \r_pwm_odd[2] ;
 wire \r_pwm_odd[3] ;
 wire \r_pwm_odd[4] ;
 wire \r_pwm_odd[5] ;
 wire \r_pwm_odd[6] ;
 wire \r_pwm_odd[7] ;
 wire \r_pwm_odd[8] ;
 wire \r_pwm_odd[9] ;
 wire rom_data_pending;
 wire \rom_last_read_addr[0] ;
 wire \rom_last_read_addr[10] ;
 wire \rom_last_read_addr[11] ;
 wire \rom_last_read_addr[1] ;
 wire \rom_last_read_addr[2] ;
 wire \rom_last_read_addr[3] ;
 wire \rom_last_read_addr[4] ;
 wire \rom_last_read_addr[5] ;
 wire \rom_last_read_addr[6] ;
 wire \rom_last_read_addr[7] ;
 wire \rom_last_read_addr[8] ;
 wire \rom_last_read_addr[9] ;
 wire \rom_next_addr_in_queue[0] ;
 wire \rom_next_addr_in_queue[10] ;
 wire \rom_next_addr_in_queue[11] ;
 wire \rom_next_addr_in_queue[1] ;
 wire \rom_next_addr_in_queue[2] ;
 wire \rom_next_addr_in_queue[3] ;
 wire \rom_next_addr_in_queue[4] ;
 wire \rom_next_addr_in_queue[5] ;
 wire \rom_next_addr_in_queue[6] ;
 wire \rom_next_addr_in_queue[7] ;
 wire \rom_next_addr_in_queue[8] ;
 wire \rom_next_addr_in_queue[9] ;
 wire \scanline[0][0] ;
 wire \scanline[0][1] ;
 wire \scanline[0][2] ;
 wire \scanline[0][3] ;
 wire \scanline[0][4] ;
 wire \scanline[0][5] ;
 wire \scanline[0][6] ;
 wire \scanline[100][0] ;
 wire \scanline[100][1] ;
 wire \scanline[100][2] ;
 wire \scanline[100][3] ;
 wire \scanline[100][4] ;
 wire \scanline[100][5] ;
 wire \scanline[100][6] ;
 wire \scanline[101][0] ;
 wire \scanline[101][1] ;
 wire \scanline[101][2] ;
 wire \scanline[101][3] ;
 wire \scanline[101][4] ;
 wire \scanline[101][5] ;
 wire \scanline[101][6] ;
 wire \scanline[102][0] ;
 wire \scanline[102][1] ;
 wire \scanline[102][2] ;
 wire \scanline[102][3] ;
 wire \scanline[102][4] ;
 wire \scanline[102][5] ;
 wire \scanline[102][6] ;
 wire \scanline[103][0] ;
 wire \scanline[103][1] ;
 wire \scanline[103][2] ;
 wire \scanline[103][3] ;
 wire \scanline[103][4] ;
 wire \scanline[103][5] ;
 wire \scanline[103][6] ;
 wire \scanline[104][0] ;
 wire \scanline[104][1] ;
 wire \scanline[104][2] ;
 wire \scanline[104][3] ;
 wire \scanline[104][4] ;
 wire \scanline[104][5] ;
 wire \scanline[104][6] ;
 wire \scanline[105][0] ;
 wire \scanline[105][1] ;
 wire \scanline[105][2] ;
 wire \scanline[105][3] ;
 wire \scanline[105][4] ;
 wire \scanline[105][5] ;
 wire \scanline[105][6] ;
 wire \scanline[106][0] ;
 wire \scanline[106][1] ;
 wire \scanline[106][2] ;
 wire \scanline[106][3] ;
 wire \scanline[106][4] ;
 wire \scanline[106][5] ;
 wire \scanline[106][6] ;
 wire \scanline[107][0] ;
 wire \scanline[107][1] ;
 wire \scanline[107][2] ;
 wire \scanline[107][3] ;
 wire \scanline[107][4] ;
 wire \scanline[107][5] ;
 wire \scanline[107][6] ;
 wire \scanline[108][0] ;
 wire \scanline[108][1] ;
 wire \scanline[108][2] ;
 wire \scanline[108][3] ;
 wire \scanline[108][4] ;
 wire \scanline[108][5] ;
 wire \scanline[108][6] ;
 wire \scanline[109][0] ;
 wire \scanline[109][1] ;
 wire \scanline[109][2] ;
 wire \scanline[109][3] ;
 wire \scanline[109][4] ;
 wire \scanline[109][5] ;
 wire \scanline[109][6] ;
 wire \scanline[10][0] ;
 wire \scanline[10][1] ;
 wire \scanline[10][2] ;
 wire \scanline[10][3] ;
 wire \scanline[10][4] ;
 wire \scanline[10][5] ;
 wire \scanline[10][6] ;
 wire \scanline[110][0] ;
 wire \scanline[110][1] ;
 wire \scanline[110][2] ;
 wire \scanline[110][3] ;
 wire \scanline[110][4] ;
 wire \scanline[110][5] ;
 wire \scanline[110][6] ;
 wire \scanline[111][0] ;
 wire \scanline[111][1] ;
 wire \scanline[111][2] ;
 wire \scanline[111][3] ;
 wire \scanline[111][4] ;
 wire \scanline[111][5] ;
 wire \scanline[111][6] ;
 wire \scanline[112][0] ;
 wire \scanline[112][1] ;
 wire \scanline[112][2] ;
 wire \scanline[112][3] ;
 wire \scanline[112][4] ;
 wire \scanline[112][5] ;
 wire \scanline[112][6] ;
 wire \scanline[113][0] ;
 wire \scanline[113][1] ;
 wire \scanline[113][2] ;
 wire \scanline[113][3] ;
 wire \scanline[113][4] ;
 wire \scanline[113][5] ;
 wire \scanline[113][6] ;
 wire \scanline[114][0] ;
 wire \scanline[114][1] ;
 wire \scanline[114][2] ;
 wire \scanline[114][3] ;
 wire \scanline[114][4] ;
 wire \scanline[114][5] ;
 wire \scanline[114][6] ;
 wire \scanline[115][0] ;
 wire \scanline[115][1] ;
 wire \scanline[115][2] ;
 wire \scanline[115][3] ;
 wire \scanline[115][4] ;
 wire \scanline[115][5] ;
 wire \scanline[115][6] ;
 wire \scanline[116][0] ;
 wire \scanline[116][1] ;
 wire \scanline[116][2] ;
 wire \scanline[116][3] ;
 wire \scanline[116][4] ;
 wire \scanline[116][5] ;
 wire \scanline[116][6] ;
 wire \scanline[117][0] ;
 wire \scanline[117][1] ;
 wire \scanline[117][2] ;
 wire \scanline[117][3] ;
 wire \scanline[117][4] ;
 wire \scanline[117][5] ;
 wire \scanline[117][6] ;
 wire \scanline[118][0] ;
 wire \scanline[118][1] ;
 wire \scanline[118][2] ;
 wire \scanline[118][3] ;
 wire \scanline[118][4] ;
 wire \scanline[118][5] ;
 wire \scanline[118][6] ;
 wire \scanline[119][0] ;
 wire \scanline[119][1] ;
 wire \scanline[119][2] ;
 wire \scanline[119][3] ;
 wire \scanline[119][4] ;
 wire \scanline[119][5] ;
 wire \scanline[119][6] ;
 wire \scanline[11][0] ;
 wire \scanline[11][1] ;
 wire \scanline[11][2] ;
 wire \scanline[11][3] ;
 wire \scanline[11][4] ;
 wire \scanline[11][5] ;
 wire \scanline[11][6] ;
 wire \scanline[120][0] ;
 wire \scanline[120][1] ;
 wire \scanline[120][2] ;
 wire \scanline[120][3] ;
 wire \scanline[120][4] ;
 wire \scanline[120][5] ;
 wire \scanline[120][6] ;
 wire \scanline[121][0] ;
 wire \scanline[121][1] ;
 wire \scanline[121][2] ;
 wire \scanline[121][3] ;
 wire \scanline[121][4] ;
 wire \scanline[121][5] ;
 wire \scanline[121][6] ;
 wire \scanline[122][0] ;
 wire \scanline[122][1] ;
 wire \scanline[122][2] ;
 wire \scanline[122][3] ;
 wire \scanline[122][4] ;
 wire \scanline[122][5] ;
 wire \scanline[122][6] ;
 wire \scanline[123][0] ;
 wire \scanline[123][1] ;
 wire \scanline[123][2] ;
 wire \scanline[123][3] ;
 wire \scanline[123][4] ;
 wire \scanline[123][5] ;
 wire \scanline[123][6] ;
 wire \scanline[124][0] ;
 wire \scanline[124][1] ;
 wire \scanline[124][2] ;
 wire \scanline[124][3] ;
 wire \scanline[124][4] ;
 wire \scanline[124][5] ;
 wire \scanline[124][6] ;
 wire \scanline[125][0] ;
 wire \scanline[125][1] ;
 wire \scanline[125][2] ;
 wire \scanline[125][3] ;
 wire \scanline[125][4] ;
 wire \scanline[125][5] ;
 wire \scanline[125][6] ;
 wire \scanline[126][0] ;
 wire \scanline[126][1] ;
 wire \scanline[126][2] ;
 wire \scanline[126][3] ;
 wire \scanline[126][4] ;
 wire \scanline[126][5] ;
 wire \scanline[126][6] ;
 wire \scanline[127][0] ;
 wire \scanline[127][1] ;
 wire \scanline[127][2] ;
 wire \scanline[127][3] ;
 wire \scanline[127][4] ;
 wire \scanline[127][5] ;
 wire \scanline[127][6] ;
 wire \scanline[128][0] ;
 wire \scanline[128][1] ;
 wire \scanline[128][2] ;
 wire \scanline[128][3] ;
 wire \scanline[128][4] ;
 wire \scanline[128][5] ;
 wire \scanline[128][6] ;
 wire \scanline[129][0] ;
 wire \scanline[129][1] ;
 wire \scanline[129][2] ;
 wire \scanline[129][3] ;
 wire \scanline[129][4] ;
 wire \scanline[129][5] ;
 wire \scanline[129][6] ;
 wire \scanline[12][0] ;
 wire \scanline[12][1] ;
 wire \scanline[12][2] ;
 wire \scanline[12][3] ;
 wire \scanline[12][4] ;
 wire \scanline[12][5] ;
 wire \scanline[12][6] ;
 wire \scanline[130][0] ;
 wire \scanline[130][1] ;
 wire \scanline[130][2] ;
 wire \scanline[130][3] ;
 wire \scanline[130][4] ;
 wire \scanline[130][5] ;
 wire \scanline[130][6] ;
 wire \scanline[131][0] ;
 wire \scanline[131][1] ;
 wire \scanline[131][2] ;
 wire \scanline[131][3] ;
 wire \scanline[131][4] ;
 wire \scanline[131][5] ;
 wire \scanline[131][6] ;
 wire \scanline[132][0] ;
 wire \scanline[132][1] ;
 wire \scanline[132][2] ;
 wire \scanline[132][3] ;
 wire \scanline[132][4] ;
 wire \scanline[132][5] ;
 wire \scanline[132][6] ;
 wire \scanline[133][0] ;
 wire \scanline[133][1] ;
 wire \scanline[133][2] ;
 wire \scanline[133][3] ;
 wire \scanline[133][4] ;
 wire \scanline[133][5] ;
 wire \scanline[133][6] ;
 wire \scanline[134][0] ;
 wire \scanline[134][1] ;
 wire \scanline[134][2] ;
 wire \scanline[134][3] ;
 wire \scanline[134][4] ;
 wire \scanline[134][5] ;
 wire \scanline[134][6] ;
 wire \scanline[135][0] ;
 wire \scanline[135][1] ;
 wire \scanline[135][2] ;
 wire \scanline[135][3] ;
 wire \scanline[135][4] ;
 wire \scanline[135][5] ;
 wire \scanline[135][6] ;
 wire \scanline[136][0] ;
 wire \scanline[136][1] ;
 wire \scanline[136][2] ;
 wire \scanline[136][3] ;
 wire \scanline[136][4] ;
 wire \scanline[136][5] ;
 wire \scanline[136][6] ;
 wire \scanline[137][0] ;
 wire \scanline[137][1] ;
 wire \scanline[137][2] ;
 wire \scanline[137][3] ;
 wire \scanline[137][4] ;
 wire \scanline[137][5] ;
 wire \scanline[137][6] ;
 wire \scanline[138][0] ;
 wire \scanline[138][1] ;
 wire \scanline[138][2] ;
 wire \scanline[138][3] ;
 wire \scanline[138][4] ;
 wire \scanline[138][5] ;
 wire \scanline[138][6] ;
 wire \scanline[139][0] ;
 wire \scanline[139][1] ;
 wire \scanline[139][2] ;
 wire \scanline[139][3] ;
 wire \scanline[139][4] ;
 wire \scanline[139][5] ;
 wire \scanline[139][6] ;
 wire \scanline[13][0] ;
 wire \scanline[13][1] ;
 wire \scanline[13][2] ;
 wire \scanline[13][3] ;
 wire \scanline[13][4] ;
 wire \scanline[13][5] ;
 wire \scanline[13][6] ;
 wire \scanline[140][0] ;
 wire \scanline[140][1] ;
 wire \scanline[140][2] ;
 wire \scanline[140][3] ;
 wire \scanline[140][4] ;
 wire \scanline[140][5] ;
 wire \scanline[140][6] ;
 wire \scanline[141][0] ;
 wire \scanline[141][1] ;
 wire \scanline[141][2] ;
 wire \scanline[141][3] ;
 wire \scanline[141][4] ;
 wire \scanline[141][5] ;
 wire \scanline[141][6] ;
 wire \scanline[142][0] ;
 wire \scanline[142][1] ;
 wire \scanline[142][2] ;
 wire \scanline[142][3] ;
 wire \scanline[142][4] ;
 wire \scanline[142][5] ;
 wire \scanline[142][6] ;
 wire \scanline[143][0] ;
 wire \scanline[143][1] ;
 wire \scanline[143][2] ;
 wire \scanline[143][3] ;
 wire \scanline[143][4] ;
 wire \scanline[143][5] ;
 wire \scanline[143][6] ;
 wire \scanline[144][0] ;
 wire \scanline[144][1] ;
 wire \scanline[144][2] ;
 wire \scanline[144][3] ;
 wire \scanline[144][4] ;
 wire \scanline[144][5] ;
 wire \scanline[144][6] ;
 wire \scanline[145][0] ;
 wire \scanline[145][1] ;
 wire \scanline[145][2] ;
 wire \scanline[145][3] ;
 wire \scanline[145][4] ;
 wire \scanline[145][5] ;
 wire \scanline[145][6] ;
 wire \scanline[146][0] ;
 wire \scanline[146][1] ;
 wire \scanline[146][2] ;
 wire \scanline[146][3] ;
 wire \scanline[146][4] ;
 wire \scanline[146][5] ;
 wire \scanline[146][6] ;
 wire \scanline[147][0] ;
 wire \scanline[147][1] ;
 wire \scanline[147][2] ;
 wire \scanline[147][3] ;
 wire \scanline[147][4] ;
 wire \scanline[147][5] ;
 wire \scanline[147][6] ;
 wire \scanline[148][0] ;
 wire \scanline[148][1] ;
 wire \scanline[148][2] ;
 wire \scanline[148][3] ;
 wire \scanline[148][4] ;
 wire \scanline[148][5] ;
 wire \scanline[148][6] ;
 wire \scanline[149][0] ;
 wire \scanline[149][1] ;
 wire \scanline[149][2] ;
 wire \scanline[149][3] ;
 wire \scanline[149][4] ;
 wire \scanline[149][5] ;
 wire \scanline[149][6] ;
 wire \scanline[14][0] ;
 wire \scanline[14][1] ;
 wire \scanline[14][2] ;
 wire \scanline[14][3] ;
 wire \scanline[14][4] ;
 wire \scanline[14][5] ;
 wire \scanline[14][6] ;
 wire \scanline[150][0] ;
 wire \scanline[150][1] ;
 wire \scanline[150][2] ;
 wire \scanline[150][3] ;
 wire \scanline[150][4] ;
 wire \scanline[150][5] ;
 wire \scanline[150][6] ;
 wire \scanline[151][0] ;
 wire \scanline[151][1] ;
 wire \scanline[151][2] ;
 wire \scanline[151][3] ;
 wire \scanline[151][4] ;
 wire \scanline[151][5] ;
 wire \scanline[151][6] ;
 wire \scanline[152][0] ;
 wire \scanline[152][1] ;
 wire \scanline[152][2] ;
 wire \scanline[152][3] ;
 wire \scanline[152][4] ;
 wire \scanline[152][5] ;
 wire \scanline[152][6] ;
 wire \scanline[153][0] ;
 wire \scanline[153][1] ;
 wire \scanline[153][2] ;
 wire \scanline[153][3] ;
 wire \scanline[153][4] ;
 wire \scanline[153][5] ;
 wire \scanline[153][6] ;
 wire \scanline[154][0] ;
 wire \scanline[154][1] ;
 wire \scanline[154][2] ;
 wire \scanline[154][3] ;
 wire \scanline[154][4] ;
 wire \scanline[154][5] ;
 wire \scanline[154][6] ;
 wire \scanline[155][0] ;
 wire \scanline[155][1] ;
 wire \scanline[155][2] ;
 wire \scanline[155][3] ;
 wire \scanline[155][4] ;
 wire \scanline[155][5] ;
 wire \scanline[155][6] ;
 wire \scanline[156][0] ;
 wire \scanline[156][1] ;
 wire \scanline[156][2] ;
 wire \scanline[156][3] ;
 wire \scanline[156][4] ;
 wire \scanline[156][5] ;
 wire \scanline[156][6] ;
 wire \scanline[157][0] ;
 wire \scanline[157][1] ;
 wire \scanline[157][2] ;
 wire \scanline[157][3] ;
 wire \scanline[157][4] ;
 wire \scanline[157][5] ;
 wire \scanline[157][6] ;
 wire \scanline[158][0] ;
 wire \scanline[158][1] ;
 wire \scanline[158][2] ;
 wire \scanline[158][3] ;
 wire \scanline[158][4] ;
 wire \scanline[158][5] ;
 wire \scanline[158][6] ;
 wire \scanline[159][0] ;
 wire \scanline[159][1] ;
 wire \scanline[159][2] ;
 wire \scanline[159][3] ;
 wire \scanline[159][4] ;
 wire \scanline[159][5] ;
 wire \scanline[159][6] ;
 wire \scanline[15][0] ;
 wire \scanline[15][1] ;
 wire \scanline[15][2] ;
 wire \scanline[15][3] ;
 wire \scanline[15][4] ;
 wire \scanline[15][5] ;
 wire \scanline[15][6] ;
 wire \scanline[16][0] ;
 wire \scanline[16][1] ;
 wire \scanline[16][2] ;
 wire \scanline[16][3] ;
 wire \scanline[16][4] ;
 wire \scanline[16][5] ;
 wire \scanline[16][6] ;
 wire \scanline[17][0] ;
 wire \scanline[17][1] ;
 wire \scanline[17][2] ;
 wire \scanline[17][3] ;
 wire \scanline[17][4] ;
 wire \scanline[17][5] ;
 wire \scanline[17][6] ;
 wire \scanline[18][0] ;
 wire \scanline[18][1] ;
 wire \scanline[18][2] ;
 wire \scanline[18][3] ;
 wire \scanline[18][4] ;
 wire \scanline[18][5] ;
 wire \scanline[18][6] ;
 wire \scanline[19][0] ;
 wire \scanline[19][1] ;
 wire \scanline[19][2] ;
 wire \scanline[19][3] ;
 wire \scanline[19][4] ;
 wire \scanline[19][5] ;
 wire \scanline[19][6] ;
 wire \scanline[1][0] ;
 wire \scanline[1][1] ;
 wire \scanline[1][2] ;
 wire \scanline[1][3] ;
 wire \scanline[1][4] ;
 wire \scanline[1][5] ;
 wire \scanline[1][6] ;
 wire \scanline[20][0] ;
 wire \scanline[20][1] ;
 wire \scanline[20][2] ;
 wire \scanline[20][3] ;
 wire \scanline[20][4] ;
 wire \scanline[20][5] ;
 wire \scanline[20][6] ;
 wire \scanline[21][0] ;
 wire \scanline[21][1] ;
 wire \scanline[21][2] ;
 wire \scanline[21][3] ;
 wire \scanline[21][4] ;
 wire \scanline[21][5] ;
 wire \scanline[21][6] ;
 wire \scanline[22][0] ;
 wire \scanline[22][1] ;
 wire \scanline[22][2] ;
 wire \scanline[22][3] ;
 wire \scanline[22][4] ;
 wire \scanline[22][5] ;
 wire \scanline[22][6] ;
 wire \scanline[23][0] ;
 wire \scanline[23][1] ;
 wire \scanline[23][2] ;
 wire \scanline[23][3] ;
 wire \scanline[23][4] ;
 wire \scanline[23][5] ;
 wire \scanline[23][6] ;
 wire \scanline[24][0] ;
 wire \scanline[24][1] ;
 wire \scanline[24][2] ;
 wire \scanline[24][3] ;
 wire \scanline[24][4] ;
 wire \scanline[24][5] ;
 wire \scanline[24][6] ;
 wire \scanline[25][0] ;
 wire \scanline[25][1] ;
 wire \scanline[25][2] ;
 wire \scanline[25][3] ;
 wire \scanline[25][4] ;
 wire \scanline[25][5] ;
 wire \scanline[25][6] ;
 wire \scanline[26][0] ;
 wire \scanline[26][1] ;
 wire \scanline[26][2] ;
 wire \scanline[26][3] ;
 wire \scanline[26][4] ;
 wire \scanline[26][5] ;
 wire \scanline[26][6] ;
 wire \scanline[27][0] ;
 wire \scanline[27][1] ;
 wire \scanline[27][2] ;
 wire \scanline[27][3] ;
 wire \scanline[27][4] ;
 wire \scanline[27][5] ;
 wire \scanline[27][6] ;
 wire \scanline[28][0] ;
 wire \scanline[28][1] ;
 wire \scanline[28][2] ;
 wire \scanline[28][3] ;
 wire \scanline[28][4] ;
 wire \scanline[28][5] ;
 wire \scanline[28][6] ;
 wire \scanline[29][0] ;
 wire \scanline[29][1] ;
 wire \scanline[29][2] ;
 wire \scanline[29][3] ;
 wire \scanline[29][4] ;
 wire \scanline[29][5] ;
 wire \scanline[29][6] ;
 wire \scanline[2][0] ;
 wire \scanline[2][1] ;
 wire \scanline[2][2] ;
 wire \scanline[2][3] ;
 wire \scanline[2][4] ;
 wire \scanline[2][5] ;
 wire \scanline[2][6] ;
 wire \scanline[30][0] ;
 wire \scanline[30][1] ;
 wire \scanline[30][2] ;
 wire \scanline[30][3] ;
 wire \scanline[30][4] ;
 wire \scanline[30][5] ;
 wire \scanline[30][6] ;
 wire \scanline[31][0] ;
 wire \scanline[31][1] ;
 wire \scanline[31][2] ;
 wire \scanline[31][3] ;
 wire \scanline[31][4] ;
 wire \scanline[31][5] ;
 wire \scanline[31][6] ;
 wire \scanline[32][0] ;
 wire \scanline[32][1] ;
 wire \scanline[32][2] ;
 wire \scanline[32][3] ;
 wire \scanline[32][4] ;
 wire \scanline[32][5] ;
 wire \scanline[32][6] ;
 wire \scanline[33][0] ;
 wire \scanline[33][1] ;
 wire \scanline[33][2] ;
 wire \scanline[33][3] ;
 wire \scanline[33][4] ;
 wire \scanline[33][5] ;
 wire \scanline[33][6] ;
 wire \scanline[34][0] ;
 wire \scanline[34][1] ;
 wire \scanline[34][2] ;
 wire \scanline[34][3] ;
 wire \scanline[34][4] ;
 wire \scanline[34][5] ;
 wire \scanline[34][6] ;
 wire \scanline[35][0] ;
 wire \scanline[35][1] ;
 wire \scanline[35][2] ;
 wire \scanline[35][3] ;
 wire \scanline[35][4] ;
 wire \scanline[35][5] ;
 wire \scanline[35][6] ;
 wire \scanline[36][0] ;
 wire \scanline[36][1] ;
 wire \scanline[36][2] ;
 wire \scanline[36][3] ;
 wire \scanline[36][4] ;
 wire \scanline[36][5] ;
 wire \scanline[36][6] ;
 wire \scanline[37][0] ;
 wire \scanline[37][1] ;
 wire \scanline[37][2] ;
 wire \scanline[37][3] ;
 wire \scanline[37][4] ;
 wire \scanline[37][5] ;
 wire \scanline[37][6] ;
 wire \scanline[38][0] ;
 wire \scanline[38][1] ;
 wire \scanline[38][2] ;
 wire \scanline[38][3] ;
 wire \scanline[38][4] ;
 wire \scanline[38][5] ;
 wire \scanline[38][6] ;
 wire \scanline[39][0] ;
 wire \scanline[39][1] ;
 wire \scanline[39][2] ;
 wire \scanline[39][3] ;
 wire \scanline[39][4] ;
 wire \scanline[39][5] ;
 wire \scanline[39][6] ;
 wire \scanline[3][0] ;
 wire \scanline[3][1] ;
 wire \scanline[3][2] ;
 wire \scanline[3][3] ;
 wire \scanline[3][4] ;
 wire \scanline[3][5] ;
 wire \scanline[3][6] ;
 wire \scanline[40][0] ;
 wire \scanline[40][1] ;
 wire \scanline[40][2] ;
 wire \scanline[40][3] ;
 wire \scanline[40][4] ;
 wire \scanline[40][5] ;
 wire \scanline[40][6] ;
 wire \scanline[41][0] ;
 wire \scanline[41][1] ;
 wire \scanline[41][2] ;
 wire \scanline[41][3] ;
 wire \scanline[41][4] ;
 wire \scanline[41][5] ;
 wire \scanline[41][6] ;
 wire \scanline[42][0] ;
 wire \scanline[42][1] ;
 wire \scanline[42][2] ;
 wire \scanline[42][3] ;
 wire \scanline[42][4] ;
 wire \scanline[42][5] ;
 wire \scanline[42][6] ;
 wire \scanline[43][0] ;
 wire \scanline[43][1] ;
 wire \scanline[43][2] ;
 wire \scanline[43][3] ;
 wire \scanline[43][4] ;
 wire \scanline[43][5] ;
 wire \scanline[43][6] ;
 wire \scanline[44][0] ;
 wire \scanline[44][1] ;
 wire \scanline[44][2] ;
 wire \scanline[44][3] ;
 wire \scanline[44][4] ;
 wire \scanline[44][5] ;
 wire \scanline[44][6] ;
 wire \scanline[45][0] ;
 wire \scanline[45][1] ;
 wire \scanline[45][2] ;
 wire \scanline[45][3] ;
 wire \scanline[45][4] ;
 wire \scanline[45][5] ;
 wire \scanline[45][6] ;
 wire \scanline[46][0] ;
 wire \scanline[46][1] ;
 wire \scanline[46][2] ;
 wire \scanline[46][3] ;
 wire \scanline[46][4] ;
 wire \scanline[46][5] ;
 wire \scanline[46][6] ;
 wire \scanline[47][0] ;
 wire \scanline[47][1] ;
 wire \scanline[47][2] ;
 wire \scanline[47][3] ;
 wire \scanline[47][4] ;
 wire \scanline[47][5] ;
 wire \scanline[47][6] ;
 wire \scanline[48][0] ;
 wire \scanline[48][1] ;
 wire \scanline[48][2] ;
 wire \scanline[48][3] ;
 wire \scanline[48][4] ;
 wire \scanline[48][5] ;
 wire \scanline[48][6] ;
 wire \scanline[49][0] ;
 wire \scanline[49][1] ;
 wire \scanline[49][2] ;
 wire \scanline[49][3] ;
 wire \scanline[49][4] ;
 wire \scanline[49][5] ;
 wire \scanline[49][6] ;
 wire \scanline[4][0] ;
 wire \scanline[4][1] ;
 wire \scanline[4][2] ;
 wire \scanline[4][3] ;
 wire \scanline[4][4] ;
 wire \scanline[4][5] ;
 wire \scanline[4][6] ;
 wire \scanline[50][0] ;
 wire \scanline[50][1] ;
 wire \scanline[50][2] ;
 wire \scanline[50][3] ;
 wire \scanline[50][4] ;
 wire \scanline[50][5] ;
 wire \scanline[50][6] ;
 wire \scanline[51][0] ;
 wire \scanline[51][1] ;
 wire \scanline[51][2] ;
 wire \scanline[51][3] ;
 wire \scanline[51][4] ;
 wire \scanline[51][5] ;
 wire \scanline[51][6] ;
 wire \scanline[52][0] ;
 wire \scanline[52][1] ;
 wire \scanline[52][2] ;
 wire \scanline[52][3] ;
 wire \scanline[52][4] ;
 wire \scanline[52][5] ;
 wire \scanline[52][6] ;
 wire \scanline[53][0] ;
 wire \scanline[53][1] ;
 wire \scanline[53][2] ;
 wire \scanline[53][3] ;
 wire \scanline[53][4] ;
 wire \scanline[53][5] ;
 wire \scanline[53][6] ;
 wire \scanline[54][0] ;
 wire \scanline[54][1] ;
 wire \scanline[54][2] ;
 wire \scanline[54][3] ;
 wire \scanline[54][4] ;
 wire \scanline[54][5] ;
 wire \scanline[54][6] ;
 wire \scanline[55][0] ;
 wire \scanline[55][1] ;
 wire \scanline[55][2] ;
 wire \scanline[55][3] ;
 wire \scanline[55][4] ;
 wire \scanline[55][5] ;
 wire \scanline[55][6] ;
 wire \scanline[56][0] ;
 wire \scanline[56][1] ;
 wire \scanline[56][2] ;
 wire \scanline[56][3] ;
 wire \scanline[56][4] ;
 wire \scanline[56][5] ;
 wire \scanline[56][6] ;
 wire \scanline[57][0] ;
 wire \scanline[57][1] ;
 wire \scanline[57][2] ;
 wire \scanline[57][3] ;
 wire \scanline[57][4] ;
 wire \scanline[57][5] ;
 wire \scanline[57][6] ;
 wire \scanline[58][0] ;
 wire \scanline[58][1] ;
 wire \scanline[58][2] ;
 wire \scanline[58][3] ;
 wire \scanline[58][4] ;
 wire \scanline[58][5] ;
 wire \scanline[58][6] ;
 wire \scanline[59][0] ;
 wire \scanline[59][1] ;
 wire \scanline[59][2] ;
 wire \scanline[59][3] ;
 wire \scanline[59][4] ;
 wire \scanline[59][5] ;
 wire \scanline[59][6] ;
 wire \scanline[5][0] ;
 wire \scanline[5][1] ;
 wire \scanline[5][2] ;
 wire \scanline[5][3] ;
 wire \scanline[5][4] ;
 wire \scanline[5][5] ;
 wire \scanline[5][6] ;
 wire \scanline[60][0] ;
 wire \scanline[60][1] ;
 wire \scanline[60][2] ;
 wire \scanline[60][3] ;
 wire \scanline[60][4] ;
 wire \scanline[60][5] ;
 wire \scanline[60][6] ;
 wire \scanline[61][0] ;
 wire \scanline[61][1] ;
 wire \scanline[61][2] ;
 wire \scanline[61][3] ;
 wire \scanline[61][4] ;
 wire \scanline[61][5] ;
 wire \scanline[61][6] ;
 wire \scanline[62][0] ;
 wire \scanline[62][1] ;
 wire \scanline[62][2] ;
 wire \scanline[62][3] ;
 wire \scanline[62][4] ;
 wire \scanline[62][5] ;
 wire \scanline[62][6] ;
 wire \scanline[63][0] ;
 wire \scanline[63][1] ;
 wire \scanline[63][2] ;
 wire \scanline[63][3] ;
 wire \scanline[63][4] ;
 wire \scanline[63][5] ;
 wire \scanline[63][6] ;
 wire \scanline[64][0] ;
 wire \scanline[64][1] ;
 wire \scanline[64][2] ;
 wire \scanline[64][3] ;
 wire \scanline[64][4] ;
 wire \scanline[64][5] ;
 wire \scanline[64][6] ;
 wire \scanline[65][0] ;
 wire \scanline[65][1] ;
 wire \scanline[65][2] ;
 wire \scanline[65][3] ;
 wire \scanline[65][4] ;
 wire \scanline[65][5] ;
 wire \scanline[65][6] ;
 wire \scanline[66][0] ;
 wire \scanline[66][1] ;
 wire \scanline[66][2] ;
 wire \scanline[66][3] ;
 wire \scanline[66][4] ;
 wire \scanline[66][5] ;
 wire \scanline[66][6] ;
 wire \scanline[67][0] ;
 wire \scanline[67][1] ;
 wire \scanline[67][2] ;
 wire \scanline[67][3] ;
 wire \scanline[67][4] ;
 wire \scanline[67][5] ;
 wire \scanline[67][6] ;
 wire \scanline[68][0] ;
 wire \scanline[68][1] ;
 wire \scanline[68][2] ;
 wire \scanline[68][3] ;
 wire \scanline[68][4] ;
 wire \scanline[68][5] ;
 wire \scanline[68][6] ;
 wire \scanline[69][0] ;
 wire \scanline[69][1] ;
 wire \scanline[69][2] ;
 wire \scanline[69][3] ;
 wire \scanline[69][4] ;
 wire \scanline[69][5] ;
 wire \scanline[69][6] ;
 wire \scanline[6][0] ;
 wire \scanline[6][1] ;
 wire \scanline[6][2] ;
 wire \scanline[6][3] ;
 wire \scanline[6][4] ;
 wire \scanline[6][5] ;
 wire \scanline[6][6] ;
 wire \scanline[70][0] ;
 wire \scanline[70][1] ;
 wire \scanline[70][2] ;
 wire \scanline[70][3] ;
 wire \scanline[70][4] ;
 wire \scanline[70][5] ;
 wire \scanline[70][6] ;
 wire \scanline[71][0] ;
 wire \scanline[71][1] ;
 wire \scanline[71][2] ;
 wire \scanline[71][3] ;
 wire \scanline[71][4] ;
 wire \scanline[71][5] ;
 wire \scanline[71][6] ;
 wire \scanline[72][0] ;
 wire \scanline[72][1] ;
 wire \scanline[72][2] ;
 wire \scanline[72][3] ;
 wire \scanline[72][4] ;
 wire \scanline[72][5] ;
 wire \scanline[72][6] ;
 wire \scanline[73][0] ;
 wire \scanline[73][1] ;
 wire \scanline[73][2] ;
 wire \scanline[73][3] ;
 wire \scanline[73][4] ;
 wire \scanline[73][5] ;
 wire \scanline[73][6] ;
 wire \scanline[74][0] ;
 wire \scanline[74][1] ;
 wire \scanline[74][2] ;
 wire \scanline[74][3] ;
 wire \scanline[74][4] ;
 wire \scanline[74][5] ;
 wire \scanline[74][6] ;
 wire \scanline[75][0] ;
 wire \scanline[75][1] ;
 wire \scanline[75][2] ;
 wire \scanline[75][3] ;
 wire \scanline[75][4] ;
 wire \scanline[75][5] ;
 wire \scanline[75][6] ;
 wire \scanline[76][0] ;
 wire \scanline[76][1] ;
 wire \scanline[76][2] ;
 wire \scanline[76][3] ;
 wire \scanline[76][4] ;
 wire \scanline[76][5] ;
 wire \scanline[76][6] ;
 wire \scanline[77][0] ;
 wire \scanline[77][1] ;
 wire \scanline[77][2] ;
 wire \scanline[77][3] ;
 wire \scanline[77][4] ;
 wire \scanline[77][5] ;
 wire \scanline[77][6] ;
 wire \scanline[78][0] ;
 wire \scanline[78][1] ;
 wire \scanline[78][2] ;
 wire \scanline[78][3] ;
 wire \scanline[78][4] ;
 wire \scanline[78][5] ;
 wire \scanline[78][6] ;
 wire \scanline[79][0] ;
 wire \scanline[79][1] ;
 wire \scanline[79][2] ;
 wire \scanline[79][3] ;
 wire \scanline[79][4] ;
 wire \scanline[79][5] ;
 wire \scanline[79][6] ;
 wire \scanline[7][0] ;
 wire \scanline[7][1] ;
 wire \scanline[7][2] ;
 wire \scanline[7][3] ;
 wire \scanline[7][4] ;
 wire \scanline[7][5] ;
 wire \scanline[7][6] ;
 wire \scanline[80][0] ;
 wire \scanline[80][1] ;
 wire \scanline[80][2] ;
 wire \scanline[80][3] ;
 wire \scanline[80][4] ;
 wire \scanline[80][5] ;
 wire \scanline[80][6] ;
 wire \scanline[81][0] ;
 wire \scanline[81][1] ;
 wire \scanline[81][2] ;
 wire \scanline[81][3] ;
 wire \scanline[81][4] ;
 wire \scanline[81][5] ;
 wire \scanline[81][6] ;
 wire \scanline[82][0] ;
 wire \scanline[82][1] ;
 wire \scanline[82][2] ;
 wire \scanline[82][3] ;
 wire \scanline[82][4] ;
 wire \scanline[82][5] ;
 wire \scanline[82][6] ;
 wire \scanline[83][0] ;
 wire \scanline[83][1] ;
 wire \scanline[83][2] ;
 wire \scanline[83][3] ;
 wire \scanline[83][4] ;
 wire \scanline[83][5] ;
 wire \scanline[83][6] ;
 wire \scanline[84][0] ;
 wire \scanline[84][1] ;
 wire \scanline[84][2] ;
 wire \scanline[84][3] ;
 wire \scanline[84][4] ;
 wire \scanline[84][5] ;
 wire \scanline[84][6] ;
 wire \scanline[85][0] ;
 wire \scanline[85][1] ;
 wire \scanline[85][2] ;
 wire \scanline[85][3] ;
 wire \scanline[85][4] ;
 wire \scanline[85][5] ;
 wire \scanline[85][6] ;
 wire \scanline[86][0] ;
 wire \scanline[86][1] ;
 wire \scanline[86][2] ;
 wire \scanline[86][3] ;
 wire \scanline[86][4] ;
 wire \scanline[86][5] ;
 wire \scanline[86][6] ;
 wire \scanline[87][0] ;
 wire \scanline[87][1] ;
 wire \scanline[87][2] ;
 wire \scanline[87][3] ;
 wire \scanline[87][4] ;
 wire \scanline[87][5] ;
 wire \scanline[87][6] ;
 wire \scanline[88][0] ;
 wire \scanline[88][1] ;
 wire \scanline[88][2] ;
 wire \scanline[88][3] ;
 wire \scanline[88][4] ;
 wire \scanline[88][5] ;
 wire \scanline[88][6] ;
 wire \scanline[89][0] ;
 wire \scanline[89][1] ;
 wire \scanline[89][2] ;
 wire \scanline[89][3] ;
 wire \scanline[89][4] ;
 wire \scanline[89][5] ;
 wire \scanline[89][6] ;
 wire \scanline[8][0] ;
 wire \scanline[8][1] ;
 wire \scanline[8][2] ;
 wire \scanline[8][3] ;
 wire \scanline[8][4] ;
 wire \scanline[8][5] ;
 wire \scanline[8][6] ;
 wire \scanline[90][0] ;
 wire \scanline[90][1] ;
 wire \scanline[90][2] ;
 wire \scanline[90][3] ;
 wire \scanline[90][4] ;
 wire \scanline[90][5] ;
 wire \scanline[90][6] ;
 wire \scanline[91][0] ;
 wire \scanline[91][1] ;
 wire \scanline[91][2] ;
 wire \scanline[91][3] ;
 wire \scanline[91][4] ;
 wire \scanline[91][5] ;
 wire \scanline[91][6] ;
 wire \scanline[92][0] ;
 wire \scanline[92][1] ;
 wire \scanline[92][2] ;
 wire \scanline[92][3] ;
 wire \scanline[92][4] ;
 wire \scanline[92][5] ;
 wire \scanline[92][6] ;
 wire \scanline[93][0] ;
 wire \scanline[93][1] ;
 wire \scanline[93][2] ;
 wire \scanline[93][3] ;
 wire \scanline[93][4] ;
 wire \scanline[93][5] ;
 wire \scanline[93][6] ;
 wire \scanline[94][0] ;
 wire \scanline[94][1] ;
 wire \scanline[94][2] ;
 wire \scanline[94][3] ;
 wire \scanline[94][4] ;
 wire \scanline[94][5] ;
 wire \scanline[94][6] ;
 wire \scanline[95][0] ;
 wire \scanline[95][1] ;
 wire \scanline[95][2] ;
 wire \scanline[95][3] ;
 wire \scanline[95][4] ;
 wire \scanline[95][5] ;
 wire \scanline[95][6] ;
 wire \scanline[96][0] ;
 wire \scanline[96][1] ;
 wire \scanline[96][2] ;
 wire \scanline[96][3] ;
 wire \scanline[96][4] ;
 wire \scanline[96][5] ;
 wire \scanline[96][6] ;
 wire \scanline[97][0] ;
 wire \scanline[97][1] ;
 wire \scanline[97][2] ;
 wire \scanline[97][3] ;
 wire \scanline[97][4] ;
 wire \scanline[97][5] ;
 wire \scanline[97][6] ;
 wire \scanline[98][0] ;
 wire \scanline[98][1] ;
 wire \scanline[98][2] ;
 wire \scanline[98][3] ;
 wire \scanline[98][4] ;
 wire \scanline[98][5] ;
 wire \scanline[98][6] ;
 wire \scanline[99][0] ;
 wire \scanline[99][1] ;
 wire \scanline[99][2] ;
 wire \scanline[99][3] ;
 wire \scanline[99][4] ;
 wire \scanline[99][5] ;
 wire \scanline[99][6] ;
 wire \scanline[9][0] ;
 wire \scanline[9][1] ;
 wire \scanline[9][2] ;
 wire \scanline[9][3] ;
 wire \scanline[9][4] ;
 wire \scanline[9][5] ;
 wire \scanline[9][6] ;
 wire spi_data_ready_last;
 wire spi_restart;
 wire tia_vsync_last;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire clknet_leaf_0_clk;
 wire net4543;
 wire net4544;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net4570;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4625;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net4630;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4644;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net4997;
 wire net4998;
 wire net4999;
 wire net5000;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net5010;
 wire net5011;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5023;
 wire net5024;
 wire net5025;
 wire net5026;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5035;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5227;
 wire net5228;
 wire net5229;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net5260;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5278;
 wire net5279;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5346;
 wire net5347;
 wire net5348;
 wire net5349;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net5360;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net5386;
 wire net5387;
 wire net5388;
 wire net5389;
 wire net5390;
 wire net5391;
 wire net5392;
 wire net5393;
 wire net5394;
 wire net5395;
 wire net5396;
 wire net5397;
 wire net5398;
 wire net5399;
 wire net5400;
 wire net5401;
 wire net5402;
 wire net5403;
 wire net5404;
 wire net5405;
 wire net5406;
 wire net5407;
 wire net5408;
 wire net5409;
 wire net5410;
 wire net5411;
 wire net5412;
 wire net5413;
 wire net5414;
 wire net5415;
 wire net5416;
 wire net5417;
 wire net5418;
 wire net5419;
 wire net5420;
 wire net5421;
 wire net5422;
 wire net5423;
 wire net5424;
 wire net5425;
 wire net5426;
 wire net5427;
 wire net5428;
 wire net5429;
 wire net5430;
 wire net5431;
 wire net5432;
 wire net5433;
 wire net5434;
 wire net5435;
 wire net5436;
 wire net5437;
 wire net5438;
 wire net5439;
 wire net5440;
 wire net5441;
 wire net5442;
 wire net5443;
 wire net5444;
 wire net5445;
 wire net5446;
 wire net5447;
 wire net5448;
 wire net5449;
 wire net5450;
 wire net5451;
 wire net5452;
 wire net5453;
 wire net5454;
 wire net5455;
 wire net5456;
 wire net5457;
 wire net5458;
 wire net5459;
 wire net5460;
 wire net5461;
 wire net5462;
 wire net5463;
 wire net5464;
 wire net5465;
 wire net5466;
 wire net5467;
 wire net5468;
 wire net5469;
 wire net5470;
 wire net5471;
 wire net5472;
 wire net5473;
 wire net5474;
 wire net5475;
 wire net5476;
 wire net5477;
 wire net5478;
 wire net5479;
 wire net5480;
 wire net5481;
 wire net5482;
 wire net5483;
 wire net5484;
 wire net5485;
 wire net5486;
 wire net5487;
 wire net5488;
 wire net5489;
 wire net5490;
 wire net5491;
 wire net5492;
 wire net5493;
 wire net5494;
 wire net5495;
 wire net5496;
 wire net5497;
 wire net5498;
 wire net5499;
 wire net5500;
 wire net5501;
 wire net5502;
 wire net5503;
 wire net5504;
 wire net5505;
 wire net5506;
 wire net5507;
 wire net5508;
 wire net5509;
 wire net5510;
 wire net5511;
 wire net5512;
 wire net5513;
 wire net5514;
 wire net5515;
 wire net5516;
 wire net5517;
 wire net5518;
 wire net5519;
 wire net5520;
 wire net5521;
 wire net5522;
 wire net5523;
 wire net5524;
 wire net5525;
 wire net5526;
 wire net5527;
 wire net5528;
 wire net5529;
 wire net5530;
 wire net5531;
 wire net5532;
 wire net5533;
 wire net5534;
 wire net5535;
 wire net5536;
 wire net5537;
 wire net5538;
 wire net5539;
 wire net5540;
 wire net5541;
 wire net5542;
 wire net5543;
 wire net5544;
 wire net5545;
 wire net5546;
 wire net5547;
 wire net5548;
 wire net5549;
 wire net5550;
 wire net5551;
 wire net5552;
 wire net5553;
 wire net5554;
 wire net5555;
 wire net5556;
 wire net5557;
 wire net5558;
 wire net5559;
 wire net5560;
 wire net5561;
 wire net5562;
 wire net5563;
 wire net5564;
 wire net5565;
 wire net5566;
 wire net5567;
 wire net5568;
 wire net5569;
 wire net5570;
 wire net5571;
 wire net5572;
 wire net5573;
 wire net5574;
 wire net5575;
 wire net5576;
 wire net5577;
 wire net5578;
 wire net5579;
 wire net5580;
 wire net5581;
 wire net5582;
 wire net5583;
 wire net5584;
 wire net5585;
 wire net5586;
 wire net5587;
 wire net5588;
 wire net5589;
 wire net5590;
 wire net5591;
 wire net5592;
 wire net5593;
 wire net5594;
 wire net5595;
 wire net5596;
 wire net5597;
 wire net5598;
 wire net5599;
 wire net5600;
 wire net5601;
 wire net5602;
 wire net5603;
 wire net5604;
 wire net5605;
 wire net5606;
 wire net5607;
 wire net5608;
 wire net5609;
 wire net5610;
 wire net5611;
 wire net5612;
 wire net5613;
 wire net5614;
 wire net5615;
 wire net5616;
 wire net5617;
 wire net5618;
 wire net5619;
 wire net5620;
 wire net5621;
 wire net5622;
 wire net5623;
 wire net5624;
 wire net5625;
 wire net5626;
 wire net5627;
 wire net5628;
 wire net5629;
 wire net5630;
 wire net5631;
 wire net5632;
 wire net5633;
 wire net5634;
 wire net5635;
 wire net5636;
 wire net5637;
 wire net5638;
 wire net5639;
 wire net5640;
 wire net5641;
 wire net5642;
 wire net5643;
 wire net5644;
 wire net5645;
 wire net5646;
 wire net5647;
 wire net5648;
 wire net5649;
 wire net5650;
 wire net5651;
 wire net5652;
 wire net5653;
 wire net5654;
 wire net5655;
 wire net5656;
 wire net5657;
 wire net5658;
 wire net5659;
 wire net5660;
 wire net5661;
 wire net5662;
 wire net5663;
 wire net5664;
 wire net5665;
 wire net5666;
 wire net5667;
 wire net5668;
 wire net5669;
 wire net5670;
 wire net5671;
 wire net5672;
 wire net5673;
 wire net5674;
 wire net5675;
 wire net5676;
 wire net5677;
 wire net5678;
 wire net5679;
 wire net5680;
 wire net5681;
 wire net5682;
 wire net5683;
 wire net5684;
 wire net5685;
 wire net5686;
 wire net5687;
 wire net5688;
 wire net5689;
 wire net5690;
 wire net5691;
 wire net5692;
 wire net5693;
 wire net5694;
 wire net5695;
 wire net5696;
 wire net5697;
 wire net5698;
 wire net5699;
 wire net5700;
 wire net5701;
 wire net5702;
 wire net5703;
 wire net5704;
 wire net5705;
 wire net5706;
 wire net5707;
 wire net5708;
 wire net5709;
 wire net5710;
 wire net5711;
 wire net5712;
 wire net5713;
 wire net5714;
 wire net5715;
 wire net5716;
 wire net5717;
 wire net5718;
 wire net5719;
 wire net5720;
 wire net5721;
 wire net5722;
 wire net5723;
 wire net5724;
 wire net5725;
 wire net5726;
 wire net5727;
 wire net5728;
 wire net5729;
 wire net5730;
 wire net5731;
 wire net5732;
 wire net5733;
 wire net5734;
 wire net5735;
 wire net5736;
 wire net5737;
 wire net5738;
 wire net5739;
 wire net5740;
 wire net5741;
 wire net5742;
 wire net5743;
 wire net5744;
 wire net5745;
 wire net5746;
 wire net5747;
 wire net5748;
 wire net5749;
 wire net5750;
 wire net5751;
 wire net5752;
 wire net5753;
 wire net5754;
 wire net5755;
 wire net5756;
 wire net5757;
 wire net5758;
 wire net5759;
 wire net5760;
 wire net5761;
 wire net5762;
 wire net5763;
 wire net5764;
 wire net5765;
 wire net5766;
 wire net5767;
 wire net5768;
 wire net5769;
 wire net5770;
 wire net5771;
 wire net5772;
 wire net5773;
 wire net5774;
 wire net5775;
 wire net5776;
 wire net5777;
 wire net5778;
 wire net5779;
 wire net5780;
 wire net5781;
 wire net5782;
 wire net5783;
 wire net5784;
 wire net5785;
 wire net5786;
 wire net5787;
 wire net5788;
 wire net5789;
 wire net5790;
 wire net5791;
 wire net5792;
 wire net5793;
 wire net5794;
 wire net5795;
 wire net5796;
 wire net5797;
 wire net5798;
 wire net5799;
 wire net5800;
 wire net5801;
 wire net5802;
 wire net5803;
 wire net5804;
 wire net5805;
 wire net5806;
 wire net5807;
 wire net5808;
 wire net5809;
 wire net5810;
 wire net5811;
 wire net5812;
 wire net5813;
 wire net5814;
 wire net5815;
 wire net5816;
 wire net5817;
 wire net5818;
 wire net5819;
 wire net5820;
 wire net5821;
 wire net5822;
 wire net5823;
 wire net5824;
 wire net5825;
 wire net5826;
 wire net5827;
 wire net5828;
 wire net5829;
 wire net5830;
 wire net5831;
 wire net5832;
 wire net5833;
 wire net5834;
 wire net5835;
 wire net5836;
 wire net5837;
 wire net5838;
 wire net5839;
 wire net5840;
 wire net5841;
 wire net5842;
 wire net5843;
 wire net5844;
 wire net5845;
 wire net5846;
 wire net5847;
 wire net5848;
 wire net5849;
 wire net5850;
 wire net5851;
 wire net5852;
 wire net5853;
 wire net5854;
 wire net5855;
 wire net5856;
 wire net5857;
 wire net5858;
 wire net5859;
 wire net5860;
 wire net5861;
 wire net5862;
 wire net5863;
 wire net5864;
 wire net5865;
 wire net5866;
 wire net5867;
 wire net5868;
 wire net5869;
 wire net5870;
 wire net5871;
 wire net5872;
 wire net5873;
 wire net5874;
 wire net5875;
 wire net5876;
 wire net5877;
 wire net5878;
 wire net5879;
 wire net5880;
 wire net5881;
 wire net5882;
 wire net5883;
 wire net5884;
 wire net5885;
 wire net5886;
 wire net5887;
 wire net5888;
 wire net5889;
 wire net5890;
 wire net5891;
 wire net5892;
 wire net5893;
 wire net5894;
 wire net5895;
 wire net5896;
 wire net5897;
 wire net5898;
 wire net5899;
 wire net5900;
 wire net5901;
 wire net5902;
 wire net5903;
 wire net5904;
 wire net5905;
 wire net5906;
 wire net5907;
 wire net5908;
 wire net5909;
 wire net5910;
 wire net5911;
 wire net5912;
 wire net5913;
 wire net5914;
 wire net5915;
 wire net5916;
 wire net5917;
 wire net5918;
 wire net5919;
 wire net5920;
 wire net5921;
 wire net5922;
 wire net5923;
 wire net5924;
 wire net5925;
 wire net5926;
 wire net5927;
 wire net5928;
 wire net5929;
 wire net5930;
 wire net5931;
 wire net5932;
 wire net5933;
 wire net5934;
 wire net5935;
 wire net5936;
 wire net5937;
 wire net5938;
 wire net5939;
 wire net5940;
 wire net5941;
 wire net5942;
 wire net5943;
 wire net5944;
 wire net5945;
 wire net5946;
 wire net5947;
 wire net5948;
 wire net5949;
 wire net5950;
 wire net5951;
 wire net5952;
 wire net5953;
 wire net5954;
 wire net5955;
 wire net5956;
 wire net5957;
 wire net5958;
 wire net5959;
 wire net5960;
 wire net5961;
 wire net5962;
 wire net5963;
 wire net5964;
 wire net5965;
 wire net5966;
 wire net5967;
 wire net5968;
 wire net5969;
 wire net5970;
 wire net5971;
 wire net5972;
 wire net5973;
 wire net5974;
 wire net5975;
 wire net5976;
 wire net5977;
 wire net5978;
 wire net5979;
 wire net5980;
 wire net5981;
 wire net5982;
 wire net5983;
 wire net5984;
 wire net5985;
 wire net5986;
 wire net5987;
 wire net5988;
 wire net5989;
 wire net5990;
 wire net5991;
 wire net5992;
 wire net5993;
 wire net5994;
 wire net5995;
 wire net5996;
 wire net5997;
 wire net5998;
 wire net5999;
 wire net6000;
 wire net6001;
 wire net6002;
 wire net6003;
 wire net6004;
 wire net6005;
 wire net6006;
 wire net6007;
 wire net6008;
 wire net6009;
 wire net6010;
 wire net6011;
 wire net6012;
 wire net6013;
 wire net6014;
 wire net6015;
 wire net6016;
 wire net6017;
 wire net6018;
 wire net6019;
 wire net6020;
 wire net6021;
 wire net6022;
 wire net6023;
 wire net6024;
 wire net6025;
 wire net6026;
 wire net6027;
 wire net6028;
 wire net6029;
 wire net6030;
 wire net6031;
 wire net6032;
 wire net6033;
 wire net6034;
 wire net6035;
 wire net6036;
 wire net6037;
 wire net6038;
 wire net6039;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_leaf_313_clk;
 wire clknet_leaf_314_clk;
 wire clknet_leaf_315_clk;
 wire clknet_leaf_316_clk;
 wire clknet_leaf_317_clk;
 wire clknet_leaf_318_clk;
 wire clknet_leaf_319_clk;
 wire clknet_leaf_320_clk;
 wire clknet_leaf_321_clk;
 wire clknet_leaf_322_clk;
 wire clknet_leaf_323_clk;
 wire clknet_leaf_324_clk;
 wire clknet_leaf_325_clk;
 wire clknet_leaf_326_clk;
 wire clknet_leaf_327_clk;
 wire clknet_leaf_328_clk;
 wire clknet_leaf_329_clk;
 wire clknet_leaf_330_clk;
 wire clknet_leaf_331_clk;
 wire clknet_leaf_332_clk;
 wire clknet_leaf_333_clk;
 wire clknet_leaf_334_clk;
 wire clknet_leaf_335_clk;
 wire clknet_leaf_336_clk;
 wire clknet_leaf_337_clk;
 wire clknet_leaf_338_clk;
 wire clknet_leaf_339_clk;
 wire clknet_leaf_340_clk;
 wire clknet_leaf_341_clk;
 wire clknet_leaf_342_clk;
 wire clknet_leaf_343_clk;
 wire clknet_leaf_344_clk;
 wire clknet_leaf_345_clk;
 wire clknet_leaf_346_clk;
 wire clknet_leaf_347_clk;
 wire clknet_leaf_348_clk;
 wire clknet_leaf_349_clk;
 wire clknet_leaf_350_clk;
 wire clknet_leaf_351_clk;
 wire clknet_leaf_352_clk;
 wire clknet_leaf_353_clk;
 wire clknet_leaf_354_clk;
 wire clknet_leaf_355_clk;
 wire clknet_leaf_356_clk;
 wire clknet_leaf_357_clk;
 wire clknet_leaf_358_clk;
 wire clknet_leaf_359_clk;
 wire clknet_leaf_360_clk;
 wire clknet_leaf_361_clk;
 wire clknet_leaf_362_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4287;
 wire net4288;
 wire net4289;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4296;
 wire net4297;
 wire net4298;
 wire net4299;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4319;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net4340;
 wire net4341;
 wire net4342;
 wire net4343;
 wire net4344;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4348;
 wire net4349;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4353;
 wire net4354;
 wire net4355;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net4360;
 wire net4361;
 wire net4362;
 wire net4363;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4369;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net4380;
 wire net4381;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4388;
 wire net4389;
 wire net4390;
 wire net4391;
 wire net4392;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4397;
 wire net4398;
 wire net4399;
 wire net4400;
 wire net4401;
 wire net4402;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net4408;
 wire net4409;
 wire net4410;
 wire net4411;
 wire net4412;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4418;
 wire net4419;
 wire net4420;
 wire net4421;
 wire net4422;
 wire net4423;
 wire net4424;
 wire net4425;
 wire net4426;
 wire net4427;
 wire net4428;
 wire net4429;
 wire net4430;
 wire net4431;
 wire net4432;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net4440;
 wire net4441;
 wire net4442;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4446;
 wire net4447;
 wire net4448;
 wire net4449;
 wire net4450;
 wire net4451;
 wire net4452;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4456;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net4460;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4464;
 wire net4465;
 wire net4466;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net4470;
 wire net4471;
 wire net4472;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4476;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net4480;
 wire net4481;
 wire net4482;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4486;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4498;
 wire net4499;
 wire net4500;
 wire net4501;
 wire net4502;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4506;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4514;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4519;
 wire net4520;
 wire net4521;
 wire net4522;
 wire net4523;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4528;
 wire net4529;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4539;
 wire net4540;
 wire net4541;
 wire net4542;
 wire net6040;
 wire net6041;
 wire net6042;
 wire net6043;
 wire net6044;
 wire net6045;
 wire net6046;
 wire net6047;
 wire net6048;
 wire net6049;
 wire net6050;
 wire net6051;
 wire net6052;
 wire net6053;
 wire net6054;
 wire net6055;
 wire net6056;
 wire net6057;
 wire net6058;
 wire net6059;
 wire net6060;
 wire net6061;
 wire net6062;
 wire net6063;
 wire net6064;
 wire net6065;
 wire net6066;
 wire net6067;
 wire net6068;
 wire net6069;
 wire net6070;
 wire net6071;
 wire net6072;
 wire net6073;
 wire net6074;
 wire net6075;
 wire net6076;
 wire net6077;
 wire net6078;
 wire net6079;
 wire net6080;
 wire net6081;
 wire net6082;
 wire net6083;
 wire net6084;
 wire net6085;
 wire net6086;
 wire net6087;
 wire net6088;
 wire net6089;
 wire net6090;
 wire net6091;
 wire net6092;
 wire net6093;
 wire net6094;
 wire net6095;
 wire net6096;
 wire net6097;
 wire net6098;
 wire net6099;
 wire net6100;
 wire net6101;
 wire net6102;
 wire net6103;
 wire net6104;
 wire net6105;
 wire net6106;
 wire net6107;
 wire net6108;
 wire net6109;
 wire net6110;
 wire net6111;
 wire net6112;
 wire net6113;
 wire net6114;
 wire net6115;
 wire net6116;
 wire net6117;
 wire net6118;
 wire net6119;
 wire net6120;
 wire net6121;
 wire net6122;
 wire net6123;
 wire net6124;
 wire net6125;
 wire net6126;
 wire net6127;
 wire net6128;
 wire net6129;
 wire net6130;
 wire net6131;
 wire net6132;
 wire net6133;
 wire net6134;
 wire net6135;
 wire net6136;
 wire net6137;
 wire net6138;
 wire net6139;
 wire net6140;
 wire net6141;
 wire net6142;
 wire net6143;
 wire net6144;
 wire net6145;
 wire net6146;
 wire net6147;
 wire net6148;
 wire net6149;
 wire net6150;
 wire net6151;
 wire net6152;
 wire net6153;
 wire net6154;
 wire net6155;
 wire net6156;
 wire net6157;
 wire net6158;
 wire net6159;
 wire net6160;
 wire net6161;
 wire net6162;
 wire net6163;
 wire net6164;
 wire net6165;
 wire net6166;
 wire net6167;
 wire net6168;
 wire net6169;
 wire net6170;
 wire net6171;
 wire net6172;
 wire net6173;
 wire net6174;
 wire net6175;
 wire net6176;
 wire net6177;
 wire net6178;
 wire net6179;
 wire net6180;
 wire net6181;
 wire net6182;
 wire net6183;
 wire net6184;
 wire net6185;
 wire net6186;
 wire net6187;
 wire net6188;
 wire net6189;
 wire net6190;
 wire net6191;
 wire net6192;
 wire net6193;
 wire net6194;
 wire net6195;
 wire net6196;
 wire net6197;
 wire net6198;
 wire net6199;
 wire net6200;
 wire net6201;
 wire net6202;
 wire net6203;
 wire net6204;
 wire net6205;
 wire net6206;
 wire net6207;
 wire net6208;
 wire net6209;
 wire net6210;
 wire net6211;
 wire net6212;
 wire net6213;
 wire net6214;
 wire net6215;
 wire net6216;
 wire net6217;
 wire net6218;
 wire net6219;
 wire net6220;
 wire net6221;
 wire net6222;
 wire net6223;
 wire net6224;
 wire net6225;
 wire net6226;
 wire net6227;
 wire net6228;
 wire net6229;
 wire net6230;
 wire net6231;
 wire net6232;
 wire net6233;
 wire net6234;
 wire net6235;
 wire net6236;
 wire net6237;
 wire net6238;
 wire net6239;
 wire net6240;
 wire net6241;
 wire net6242;
 wire net6243;
 wire net6244;
 wire net6245;
 wire net6246;
 wire net6247;
 wire net6248;
 wire net6249;
 wire net6250;
 wire net6251;
 wire net6252;
 wire net6253;
 wire net6254;
 wire net6255;
 wire net6256;
 wire net6257;
 wire net6258;
 wire net6259;
 wire net6260;
 wire net6261;
 wire net6262;
 wire net6263;
 wire net6264;
 wire net6265;
 wire net6266;
 wire net6267;
 wire net6268;
 wire net6269;
 wire net6270;
 wire net6271;
 wire net6272;
 wire net6273;
 wire net6274;
 wire net6275;
 wire net6276;
 wire net6277;
 wire net6278;
 wire net6279;
 wire net6280;
 wire net6281;
 wire net6282;
 wire net6283;
 wire net6284;
 wire net6285;
 wire net6286;
 wire net6287;
 wire net6288;
 wire net6289;
 wire net6290;
 wire net6291;
 wire net6292;
 wire net6293;
 wire net6294;
 wire net6295;
 wire net6296;
 wire net6297;
 wire net6298;
 wire net6299;
 wire net6300;
 wire net6301;
 wire net6302;
 wire net6303;
 wire net6304;
 wire net6305;
 wire net6306;
 wire net6307;
 wire net6308;
 wire net6309;
 wire net6310;
 wire net6311;
 wire net6312;
 wire net6313;
 wire net6314;
 wire net6315;
 wire net6316;
 wire net6317;
 wire net6318;
 wire net6319;
 wire net6320;
 wire net6321;
 wire net6322;
 wire net6323;
 wire net6324;
 wire net6325;
 wire net6326;
 wire net6327;
 wire net6328;
 wire net6329;
 wire net6330;
 wire net6331;
 wire net6332;
 wire net6333;
 wire net6334;
 wire net6335;
 wire net6336;
 wire net6337;
 wire net6338;
 wire net6339;
 wire net6340;
 wire net6341;
 wire net6342;
 wire net6343;
 wire net6344;
 wire net6345;
 wire net6346;
 wire net6347;
 wire net6348;
 wire net6349;
 wire net6350;
 wire net6351;
 wire net6352;
 wire net6353;
 wire net6354;
 wire net6355;
 wire net6356;
 wire net6357;
 wire net6358;
 wire net6359;
 wire net6360;
 wire net6361;
 wire net6362;
 wire net6363;
 wire net6364;
 wire net6365;
 wire net6366;
 wire net6367;
 wire net6368;
 wire net6369;
 wire net6370;
 wire net6371;
 wire net6372;
 wire net6373;
 wire net6374;
 wire net6375;
 wire net6376;
 wire net6377;
 wire net6378;
 wire net6379;
 wire net6380;
 wire net6381;
 wire net6382;
 wire net6383;
 wire net6384;
 wire net6385;
 wire net6386;
 wire net6387;
 wire net6388;
 wire net6389;
 wire net6390;
 wire net6391;
 wire net6392;
 wire net6393;
 wire net6394;
 wire net6395;
 wire net6396;
 wire net6397;
 wire net6398;
 wire net6399;
 wire net6400;
 wire net6401;
 wire net6402;
 wire net6403;
 wire net6404;
 wire net6405;
 wire net6406;
 wire net6407;
 wire net6408;
 wire net6409;
 wire net6410;
 wire net6411;
 wire net6412;
 wire net6413;
 wire net6414;
 wire net6415;
 wire net6416;
 wire net6417;
 wire net6418;
 wire net6419;
 wire net6420;
 wire net6421;
 wire net6422;
 wire net6423;
 wire net6424;
 wire net6425;
 wire net6426;
 wire net6427;
 wire net6428;
 wire net6429;
 wire net6430;
 wire net6431;
 wire net6432;
 wire net6433;
 wire net6434;
 wire net6435;
 wire net6436;
 wire net6437;
 wire net6438;
 wire net6439;
 wire net6440;
 wire net6441;
 wire net6442;
 wire net6443;
 wire net6444;
 wire net6445;
 wire net6446;
 wire net6447;
 wire net6448;
 wire net6449;
 wire net6450;
 wire net6451;
 wire net6452;
 wire net6453;
 wire net6454;
 wire net6455;
 wire net6456;
 wire net6457;
 wire net6458;
 wire net6459;
 wire net6460;
 wire net6461;
 wire net6462;
 wire net6463;
 wire net6464;
 wire net6465;
 wire net6466;
 wire net6467;
 wire net6468;
 wire net6469;
 wire net6470;
 wire net6471;
 wire net6472;
 wire net6473;
 wire net6474;
 wire net6475;
 wire net6476;
 wire net6477;
 wire net6478;
 wire net6479;
 wire net6480;
 wire net6481;
 wire net6482;
 wire net6483;
 wire net6484;
 wire net6485;
 wire net6486;
 wire net6487;
 wire net6488;
 wire net6489;
 wire net6490;
 wire net6491;
 wire net6492;
 wire net6493;
 wire net6494;
 wire net6495;
 wire net6496;
 wire net6497;
 wire net6498;
 wire net6499;
 wire net6500;
 wire net6501;
 wire net6502;
 wire net6503;
 wire net6504;
 wire net6505;
 wire net6506;
 wire net6507;
 wire net6508;
 wire net6509;
 wire net6510;
 wire net6511;
 wire net6512;
 wire net6513;
 wire net6514;
 wire net6515;
 wire net6516;
 wire net6517;
 wire net6518;
 wire net6519;
 wire net6520;
 wire net6521;
 wire net6522;
 wire net6523;
 wire net6524;
 wire net6525;
 wire net6526;
 wire net6527;
 wire net6528;
 wire net6529;
 wire net6530;
 wire net6531;
 wire net6532;
 wire net6533;
 wire net6534;
 wire net6535;
 wire net6536;
 wire net6537;
 wire net6538;
 wire net6539;
 wire net6540;
 wire net6541;
 wire net6542;
 wire net6543;
 wire net6544;
 wire net6545;
 wire net6546;
 wire net6547;
 wire net6548;
 wire net6549;
 wire net6550;
 wire net6551;
 wire net6552;
 wire net6553;
 wire net6554;
 wire net6555;
 wire net6556;
 wire net6557;
 wire net6558;
 wire net6559;
 wire net6560;
 wire net6561;
 wire net6562;
 wire net6563;
 wire net6564;
 wire net6565;
 wire net6566;
 wire net6567;
 wire net6568;
 wire net6569;
 wire net6570;
 wire net6571;
 wire net6572;
 wire net6573;
 wire net6574;
 wire net6575;
 wire net6576;
 wire net6577;
 wire net6578;
 wire net6579;
 wire net6580;
 wire net6581;
 wire net6582;
 wire net6583;
 wire net6584;
 wire net6585;
 wire net6586;
 wire net6587;
 wire net6588;
 wire net6589;
 wire net6590;
 wire net6591;
 wire net6592;
 wire net6593;
 wire net6594;
 wire net6595;
 wire net6596;
 wire net6597;
 wire net6598;
 wire net6599;
 wire net6600;
 wire net6601;
 wire net6602;
 wire net6603;
 wire net6604;
 wire net6605;
 wire net6606;
 wire net6607;
 wire net6608;
 wire net6609;
 wire net6610;
 wire net6611;
 wire net6612;
 wire net6613;
 wire net6614;
 wire net6615;
 wire net6616;
 wire net6617;
 wire net6618;
 wire net6619;
 wire net6620;
 wire net6621;
 wire net6622;
 wire net6623;
 wire net6624;
 wire net6625;
 wire net6626;
 wire net6627;
 wire net6628;
 wire net6629;
 wire net6630;
 wire net6631;
 wire net6632;
 wire net6633;
 wire net6634;
 wire net6635;
 wire net6636;
 wire net6637;
 wire net6638;
 wire net6639;
 wire net6640;
 wire net6641;
 wire net6642;
 wire net6643;
 wire net6644;
 wire net6645;
 wire net6646;
 wire net6647;
 wire net6648;
 wire net6649;
 wire net6650;
 wire net6651;
 wire net6652;
 wire net6653;
 wire net6654;
 wire net6655;
 wire net6656;
 wire net6657;
 wire net6658;
 wire net6659;
 wire net6660;
 wire net6661;
 wire net6662;
 wire net6663;
 wire net6664;
 wire net6665;
 wire net6666;
 wire net6667;
 wire net6668;
 wire net6669;
 wire net6670;
 wire net6671;
 wire net6672;
 wire net6673;
 wire net6674;
 wire net6675;
 wire net6676;
 wire net6677;
 wire net6678;
 wire net6679;
 wire net6680;
 wire net6681;
 wire net6682;
 wire net6683;
 wire net6684;
 wire net6685;
 wire net6686;
 wire net6687;
 wire net6688;
 wire net6689;
 wire net6690;
 wire net6691;
 wire net6692;
 wire net6693;
 wire net6694;
 wire net6695;
 wire net6696;
 wire net6697;
 wire net6698;
 wire net6699;
 wire net6700;
 wire net6701;
 wire net6702;
 wire net6703;
 wire net6704;
 wire net6705;
 wire net6706;
 wire net6707;
 wire net6708;
 wire net6709;
 wire net6710;
 wire net6711;
 wire net6712;
 wire net6713;
 wire net6714;
 wire net6715;
 wire net6716;
 wire net6717;
 wire net6718;
 wire net6719;
 wire net6720;
 wire net6721;
 wire net6722;
 wire net6723;
 wire net6724;
 wire net6725;
 wire net6726;
 wire net6727;
 wire net6728;
 wire net6729;
 wire net6730;
 wire net6731;
 wire net6732;
 wire net6733;
 wire net6734;
 wire net6735;
 wire net6736;
 wire net6737;
 wire net6738;
 wire net6739;
 wire net6740;
 wire net6741;
 wire net6742;
 wire net6743;
 wire net6744;
 wire net6745;
 wire net6746;
 wire net6747;
 wire net6748;
 wire net6749;
 wire net6750;
 wire net6751;
 wire net6752;
 wire net6753;
 wire net6754;
 wire net6755;
 wire net6756;
 wire net6757;
 wire net6758;
 wire net6759;
 wire net6760;
 wire net6761;
 wire net6762;
 wire net6763;
 wire net6764;
 wire net6765;
 wire net6766;
 wire net6767;
 wire net6768;
 wire net6769;
 wire net6770;
 wire net6771;
 wire net6772;
 wire net6773;
 wire net6774;
 wire net6775;
 wire net6776;
 wire net6777;
 wire net6778;
 wire net6779;
 wire net6780;
 wire net6781;
 wire net6782;
 wire net6783;
 wire net6784;
 wire net6785;
 wire net6786;
 wire net6787;
 wire net6788;
 wire net6789;
 wire net6790;
 wire net6791;
 wire net6792;
 wire net6793;
 wire net6794;
 wire net6795;
 wire net6796;
 wire net6797;
 wire net6798;
 wire net6799;
 wire net6800;
 wire net6801;
 wire net6802;
 wire net6803;
 wire net6804;
 wire net6805;
 wire net6806;
 wire net6807;
 wire net6808;
 wire net6809;
 wire net6810;
 wire net6811;
 wire net6812;
 wire net6813;
 wire net6814;
 wire net6815;
 wire net6816;
 wire net6817;
 wire net6818;
 wire net6819;
 wire net6820;
 wire net6821;
 wire net6822;
 wire net6823;
 wire net6824;
 wire net6825;
 wire net6826;
 wire net6827;
 wire net6828;
 wire net6829;
 wire net6830;
 wire net6831;
 wire net6832;
 wire net6833;
 wire net6834;
 wire net6835;
 wire net6836;
 wire net6837;
 wire net6838;
 wire net6839;
 wire net6840;
 wire net6841;
 wire net6842;
 wire net6843;
 wire net6844;
 wire net6845;
 wire net6846;
 wire net6847;
 wire net6848;
 wire net6849;
 wire net6850;
 wire net6851;
 wire net6852;
 wire net6853;
 wire net6854;
 wire net6855;
 wire net6856;
 wire net6857;
 wire net6858;
 wire net6859;
 wire net6860;
 wire net6861;
 wire net6862;
 wire net6863;
 wire net6864;
 wire net6865;
 wire net6866;
 wire net6867;
 wire net6868;
 wire net6869;
 wire net6870;
 wire net6871;
 wire net6872;
 wire net6873;
 wire net6874;
 wire net6875;
 wire net6876;
 wire net6877;
 wire net6878;
 wire net6879;
 wire net6880;
 wire net6881;
 wire net6882;
 wire net6883;
 wire net6884;
 wire net6885;
 wire net6886;
 wire net6887;
 wire net6888;
 wire net6889;
 wire net6890;
 wire net6891;
 wire net6892;
 wire net6893;
 wire net6894;
 wire net6895;
 wire net6896;
 wire net6897;
 wire net6898;
 wire net6899;
 wire net6900;
 wire net6901;
 wire net6902;
 wire net6903;
 wire net6904;
 wire net6905;
 wire net6906;
 wire net6907;
 wire net6908;
 wire net6909;
 wire net6910;
 wire net6911;
 wire net6912;
 wire net6913;
 wire net6914;
 wire net6915;
 wire net6916;
 wire net6917;
 wire net6918;
 wire net6919;
 wire net6920;
 wire net6921;
 wire net6922;
 wire net6923;
 wire net6924;
 wire net6925;
 wire net6926;
 wire net6927;
 wire net6928;
 wire net6929;
 wire net6930;
 wire net6931;
 wire net6932;
 wire net6933;
 wire net6934;
 wire net6935;
 wire net6936;
 wire net6937;
 wire net6938;
 wire net6939;
 wire net6940;
 wire net6941;
 wire net6942;
 wire net6943;
 wire net6944;
 wire net6945;
 wire net6946;
 wire net6947;
 wire net6948;
 wire net6949;
 wire net6950;
 wire net6951;
 wire net6952;
 wire net6953;
 wire net6954;
 wire net6955;
 wire net6956;
 wire net6957;
 wire net6958;
 wire net6959;
 wire net6960;
 wire net6961;
 wire net6962;
 wire net6963;
 wire net6964;
 wire net6965;
 wire net6966;
 wire net6967;
 wire net6968;
 wire net6969;
 wire net6970;
 wire net6971;
 wire net6972;
 wire net6973;
 wire net6974;
 wire net6975;
 wire net6976;
 wire net6977;
 wire net6978;
 wire net6979;
 wire net6980;
 wire net6981;
 wire net6982;
 wire net6983;
 wire net6984;
 wire net6985;
 wire net6986;
 wire net6987;
 wire net6988;
 wire net6989;
 wire net6990;
 wire net6991;
 wire net6992;
 wire net6993;
 wire net6994;
 wire net6995;
 wire net6996;
 wire net6997;
 wire net6998;
 wire net6999;
 wire net7000;
 wire net7001;
 wire net7002;
 wire net7003;
 wire net7004;
 wire net7005;
 wire net7006;
 wire net7007;
 wire net7008;
 wire net7009;
 wire net7010;
 wire net7011;
 wire net7012;
 wire net7013;
 wire net7014;
 wire net7015;
 wire net7016;
 wire net7017;
 wire net7018;
 wire net7019;
 wire net7020;
 wire net7021;
 wire net7022;
 wire net7023;
 wire net7024;
 wire net7025;
 wire net7026;
 wire net7027;
 wire net7028;
 wire net7029;
 wire net7030;
 wire net7031;
 wire net7032;
 wire net7033;
 wire net7034;
 wire net7035;
 wire net7036;
 wire net7037;
 wire net7038;
 wire net7039;
 wire net7040;
 wire net7041;
 wire net7042;
 wire net7043;
 wire net7044;
 wire net7045;
 wire net7046;
 wire net7047;
 wire net7048;
 wire net7049;
 wire net7050;
 wire net7051;
 wire net7052;
 wire net7053;
 wire net7054;
 wire net7055;
 wire net7056;
 wire net7057;
 wire net7058;
 wire net7059;
 wire net7060;
 wire net7061;
 wire net7062;
 wire net7063;
 wire net7064;
 wire net7065;
 wire net7066;
 wire net7067;
 wire net7068;
 wire net7069;
 wire net7070;
 wire net7071;
 wire net7072;
 wire net7073;
 wire net7074;
 wire net7075;
 wire net7076;
 wire net7077;
 wire net7078;
 wire net7079;
 wire net7080;
 wire net7081;
 wire net7082;
 wire net7083;
 wire net7084;
 wire net7085;
 wire net7086;
 wire net7087;
 wire net7088;
 wire net7089;
 wire net7090;
 wire net7091;
 wire net7092;
 wire net7093;
 wire net7094;
 wire net7095;
 wire net7096;
 wire net7097;
 wire net7098;
 wire net7099;
 wire net7100;
 wire net7101;
 wire net7102;
 wire net7103;
 wire net7104;
 wire net7105;
 wire net7106;
 wire net7107;
 wire net7108;
 wire net7109;
 wire net7110;
 wire net7111;
 wire net7112;
 wire net7113;
 wire net7114;
 wire net7115;
 wire net7116;
 wire net7117;
 wire net7118;
 wire net7119;
 wire net7120;
 wire net7121;
 wire net7122;
 wire net7123;
 wire net7124;
 wire net7125;
 wire net7126;
 wire net7127;
 wire net7128;
 wire net7129;
 wire net7130;
 wire net7131;
 wire net7132;
 wire net7133;
 wire net7134;
 wire net7135;
 wire net7136;
 wire net7137;
 wire net7138;
 wire net7139;
 wire net7140;
 wire net7141;
 wire net7142;
 wire net7143;
 wire net7144;
 wire net7145;
 wire net7146;
 wire net7147;
 wire net7148;
 wire net7149;
 wire net7150;
 wire net7151;
 wire net7152;
 wire net7153;
 wire net7154;
 wire net7155;
 wire net7156;
 wire net7157;
 wire net7158;
 wire net7159;
 wire net7160;
 wire net7161;
 wire net7162;
 wire net7163;
 wire net7164;
 wire net7165;
 wire net7166;
 wire net7167;
 wire net7168;
 wire net7169;
 wire net7170;
 wire net7171;
 wire net7172;
 wire net7173;
 wire net7174;
 wire net7175;
 wire net7176;
 wire net7177;
 wire net7178;
 wire net7179;
 wire net7180;
 wire net7181;
 wire net7182;
 wire net7183;
 wire net7184;
 wire net7185;
 wire net7186;
 wire net7187;
 wire net7188;
 wire net7189;
 wire net7190;
 wire net7191;
 wire net7192;
 wire net7193;
 wire net7194;
 wire net7195;
 wire net7196;
 wire net7197;
 wire net7198;
 wire net7199;
 wire net7200;
 wire net7201;
 wire net7202;
 wire net7203;
 wire net7204;
 wire net7205;
 wire net7206;
 wire net7207;
 wire net7208;
 wire net7209;
 wire net7210;
 wire net7211;
 wire net7212;
 wire net7213;
 wire net7214;
 wire net7215;
 wire net7216;
 wire net7217;
 wire net7218;
 wire net7219;
 wire net7220;
 wire net7221;
 wire net7222;
 wire net7223;
 wire net7224;
 wire net7225;
 wire net7226;
 wire net7227;
 wire net7228;
 wire net7229;
 wire net7230;
 wire net7231;
 wire net7232;
 wire net7233;
 wire net7234;
 wire net7235;
 wire net7236;
 wire net7237;
 wire net7238;
 wire net7239;
 wire net7240;
 wire net7241;
 wire net7242;
 wire net7243;
 wire net7244;
 wire net7245;
 wire net7246;
 wire net7247;
 wire net7248;
 wire net7249;
 wire net7250;
 wire net7251;
 wire net7252;
 wire net7253;
 wire net7254;
 wire net7255;
 wire net7256;
 wire net7257;
 wire net7258;
 wire net7259;
 wire net7260;
 wire net7261;
 wire net7262;
 wire net7263;
 wire net7264;
 wire net7265;
 wire net7266;
 wire net7267;
 wire net7268;
 wire net7269;
 wire net7270;
 wire net7271;
 wire net7272;
 wire net7273;
 wire net7274;
 wire net7275;
 wire net7276;
 wire net7277;
 wire net7278;
 wire net7279;
 wire net7280;
 wire net7281;
 wire net7282;
 wire net7283;
 wire net7284;
 wire net7285;
 wire net7286;
 wire net7287;
 wire net7288;
 wire net7289;
 wire net7290;
 wire net7291;
 wire net7292;
 wire net7293;
 wire net7294;
 wire net7295;
 wire net7296;
 wire net7297;
 wire net7298;
 wire net7299;
 wire net7300;
 wire net7301;
 wire net7302;
 wire net7303;
 wire net7304;
 wire net7305;
 wire net7306;
 wire net7307;
 wire net7308;
 wire net7309;
 wire net7310;
 wire net7311;
 wire net7312;
 wire net7313;
 wire net7314;
 wire net7315;
 wire net7316;
 wire net7317;
 wire net7318;
 wire net7319;
 wire net7320;
 wire net7321;
 wire net7322;
 wire net7323;
 wire net7324;
 wire net7325;
 wire net7326;
 wire net7327;
 wire net7328;
 wire net7329;
 wire net7330;
 wire net7331;
 wire net7332;
 wire net7333;
 wire net7334;
 wire net7335;
 wire net7336;
 wire net7337;
 wire net7338;
 wire net7339;
 wire net7340;
 wire net7341;
 wire net7342;
 wire net7343;
 wire net7344;
 wire net7345;
 wire net7346;
 wire net7347;
 wire net7348;
 wire net7349;
 wire net7350;
 wire net7351;
 wire net7352;
 wire net7353;
 wire net7354;
 wire net7355;
 wire net7356;
 wire net7357;
 wire net7358;
 wire net7359;
 wire net7360;
 wire net7361;
 wire net7362;
 wire net7363;
 wire net7364;
 wire net7365;
 wire net7366;
 wire net7367;
 wire net7368;
 wire net7369;
 wire net7370;
 wire net7371;
 wire net7372;
 wire net7373;
 wire net7374;
 wire net7375;
 wire net7376;
 wire net7377;
 wire net7378;
 wire net7379;
 wire net7380;

 sg13g2_inv_1 _16142_ (.Y(_07920_),
    .A(net7178));
 sg13g2_inv_1 _16143_ (.Y(_07921_),
    .A(net5567));
 sg13g2_inv_1 _16144_ (.Y(_07922_),
    .A(net7174));
 sg13g2_inv_1 _16145_ (.Y(_07923_),
    .A(\atari2600.clk_counter[1] ));
 sg13g2_inv_1 _16146_ (.Y(_07924_),
    .A(\atari2600.clk_counter[0] ));
 sg13g2_inv_1 _16147_ (.Y(_07925_),
    .A(\atari2600.tia.diag[86] ));
 sg13g2_inv_1 _16148_ (.Y(_07926_),
    .A(\atari2600.tia.diag[82] ));
 sg13g2_inv_1 _16149_ (.Y(_07927_),
    .A(net2993));
 sg13g2_inv_1 _16150_ (.Y(_07928_),
    .A(net3659));
 sg13g2_inv_1 _16151_ (.Y(_07929_),
    .A(net2978));
 sg13g2_inv_1 _16152_ (.Y(_07930_),
    .A(\atari2600.tia.poly9_r.x[5] ));
 sg13g2_inv_1 _16153_ (.Y(_07931_),
    .A(\atari2600.tia.poly9_r.x[4] ));
 sg13g2_inv_1 _16154_ (.Y(_07932_),
    .A(\atari2600.tia.poly9_r.x[1] ));
 sg13g2_inv_1 _16155_ (.Y(_07933_),
    .A(net7016));
 sg13g2_inv_1 _16156_ (.Y(_07934_),
    .A(net3056));
 sg13g2_inv_1 _16157_ (.Y(_07935_),
    .A(\atari2600.tia.poly5_r.x[1] ));
 sg13g2_inv_1 _16158_ (.Y(_07936_),
    .A(net7001));
 sg13g2_inv_1 _16159_ (.Y(_07937_),
    .A(net6877));
 sg13g2_inv_1 _16160_ (.Y(_07938_),
    .A(net6818));
 sg13g2_inv_1 _16161_ (.Y(_07939_),
    .A(net4119));
 sg13g2_inv_1 _16162_ (.Y(_07940_),
    .A(net3753));
 sg13g2_inv_1 _16163_ (.Y(_07941_),
    .A(net3801));
 sg13g2_inv_1 _16164_ (.Y(_07942_),
    .A(net3913));
 sg13g2_inv_1 _16165_ (.Y(_07943_),
    .A(net3232));
 sg13g2_inv_1 _16166_ (.Y(_07944_),
    .A(net3505));
 sg13g2_inv_1 _16167_ (.Y(_07945_),
    .A(net3865));
 sg13g2_inv_2 _16168_ (.Y(_07946_),
    .A(net7311));
 sg13g2_inv_1 _16169_ (.Y(_07947_),
    .A(net5578));
 sg13g2_inv_1 _16170_ (.Y(_07948_),
    .A(net5579));
 sg13g2_inv_1 _16171_ (.Y(_07949_),
    .A(net5581));
 sg13g2_inv_1 _16172_ (.Y(_07950_),
    .A(net2950));
 sg13g2_inv_2 _16173_ (.Y(_07951_),
    .A(net7333));
 sg13g2_inv_1 _16174_ (.Y(_07952_),
    .A(net7263));
 sg13g2_inv_1 _16175_ (.Y(_07953_),
    .A(net7272));
 sg13g2_inv_1 _16176_ (.Y(_07954_),
    .A(net6979));
 sg13g2_inv_1 _16177_ (.Y(_07955_),
    .A(net4224));
 sg13g2_inv_1 _16178_ (.Y(_07956_),
    .A(net3893));
 sg13g2_inv_1 _16179_ (.Y(_07957_),
    .A(net3277));
 sg13g2_inv_1 _16180_ (.Y(_07958_),
    .A(net3379));
 sg13g2_inv_1 _16181_ (.Y(_07959_),
    .A(net3378));
 sg13g2_inv_1 _16182_ (.Y(_07960_),
    .A(net2988));
 sg13g2_inv_1 _16183_ (.Y(_07961_),
    .A(net2992));
 sg13g2_inv_1 _16184_ (.Y(_07962_),
    .A(net2936));
 sg13g2_inv_2 _16185_ (.Y(_07963_),
    .A(net7291));
 sg13g2_inv_2 _16186_ (.Y(_07964_),
    .A(net5583));
 sg13g2_inv_1 _16187_ (.Y(_07965_),
    .A(net7261));
 sg13g2_inv_1 _16188_ (.Y(_07966_),
    .A(net7268));
 sg13g2_inv_2 _16189_ (.Y(_07967_),
    .A(net7275));
 sg13g2_inv_1 _16190_ (.Y(_07968_),
    .A(\atari2600.tia.audc0[0] ));
 sg13g2_inv_1 _16191_ (.Y(_07969_),
    .A(net5584));
 sg13g2_inv_1 _16192_ (.Y(_07970_),
    .A(\atari2600.tia.hmbl[2] ));
 sg13g2_inv_1 _16193_ (.Y(_07971_),
    .A(\atari2600.tia.hmm1[3] ));
 sg13g2_inv_1 _16194_ (.Y(_07972_),
    .A(net5586));
 sg13g2_inv_1 _16195_ (.Y(_07973_),
    .A(\atari2600.tia.hmm0[1] ));
 sg13g2_inv_1 _16196_ (.Y(_07974_),
    .A(net5587));
 sg13g2_inv_1 _16197_ (.Y(_07975_),
    .A(\atari2600.tia.hmp1[2] ));
 sg13g2_inv_1 _16198_ (.Y(_07976_),
    .A(net5588));
 sg13g2_inv_1 _16199_ (.Y(_07977_),
    .A(\atari2600.tia.hmp0[2] ));
 sg13g2_inv_1 _16200_ (.Y(_07978_),
    .A(\atari2600.tia.diag[38] ));
 sg13g2_inv_1 _16201_ (.Y(_07979_),
    .A(\atari2600.tia.diag[37] ));
 sg13g2_inv_1 _16202_ (.Y(_07980_),
    .A(\atari2600.tia.diag[36] ));
 sg13g2_inv_1 _16203_ (.Y(_07981_),
    .A(\atari2600.tia.diag[35] ));
 sg13g2_inv_1 _16204_ (.Y(_07982_),
    .A(\atari2600.tia.diag[34] ));
 sg13g2_inv_1 _16205_ (.Y(_07983_),
    .A(\atari2600.tia.diag[33] ));
 sg13g2_inv_1 _16206_ (.Y(_07984_),
    .A(\atari2600.tia.diag[46] ));
 sg13g2_inv_1 _16207_ (.Y(_07985_),
    .A(\atari2600.tia.diag[45] ));
 sg13g2_inv_1 _16208_ (.Y(_07986_),
    .A(\atari2600.tia.diag[44] ));
 sg13g2_inv_2 _16209_ (.Y(_07987_),
    .A(net7166));
 sg13g2_inv_1 _16210_ (.Y(_07988_),
    .A(net7328));
 sg13g2_inv_1 _16211_ (.Y(_07989_),
    .A(net7350));
 sg13g2_inv_2 _16212_ (.Y(_07990_),
    .A(net7260));
 sg13g2_inv_1 _16213_ (.Y(_07991_),
    .A(\atari2600.tia.diag[50] ));
 sg13g2_inv_1 _16214_ (.Y(_07992_),
    .A(\atari2600.tia.diag[62] ));
 sg13g2_inv_2 _16215_ (.Y(_07993_),
    .A(\atari2600.tia.diag[61] ));
 sg13g2_inv_1 _16216_ (.Y(_07994_),
    .A(net5592));
 sg13g2_inv_2 _16217_ (.Y(_07995_),
    .A(\atari2600.tia.diag[70] ));
 sg13g2_inv_1 _16218_ (.Y(_07996_),
    .A(net5593));
 sg13g2_inv_1 _16219_ (.Y(_07997_),
    .A(net5594));
 sg13g2_inv_1 _16220_ (.Y(_07998_),
    .A(\atari2600.tia.diag[67] ));
 sg13g2_inv_2 _16221_ (.Y(_07999_),
    .A(\atari2600.tia.diag[65] ));
 sg13g2_inv_1 _16222_ (.Y(_08000_),
    .A(net3959));
 sg13g2_inv_1 _16223_ (.Y(_08001_),
    .A(net4088));
 sg13g2_inv_1 _16224_ (.Y(_08002_),
    .A(net4073));
 sg13g2_inv_1 _16225_ (.Y(_08003_),
    .A(net4278));
 sg13g2_inv_1 _16226_ (.Y(_08004_),
    .A(net6943));
 sg13g2_inv_1 _16227_ (.Y(_08005_),
    .A(net4163));
 sg13g2_inv_1 _16228_ (.Y(_08006_),
    .A(net4014));
 sg13g2_inv_1 _16229_ (.Y(_08007_),
    .A(net3369));
 sg13g2_inv_1 _16230_ (.Y(_08008_),
    .A(net3788));
 sg13g2_inv_1 _16231_ (.Y(_08009_),
    .A(net7321));
 sg13g2_inv_1 _16232_ (.Y(_08010_),
    .A(net7300));
 sg13g2_inv_1 _16233_ (.Y(_08011_),
    .A(\atari2600.tia.colupf[6] ));
 sg13g2_inv_1 _16234_ (.Y(_08012_),
    .A(\atari2600.tia.colupf[5] ));
 sg13g2_inv_1 _16235_ (.Y(_08013_),
    .A(\atari2600.tia.colupf[4] ));
 sg13g2_inv_1 _16236_ (.Y(_08014_),
    .A(\atari2600.tia.colupf[3] ));
 sg13g2_inv_1 _16237_ (.Y(_08015_),
    .A(\atari2600.tia.colupf[2] ));
 sg13g2_inv_1 _16238_ (.Y(_08016_),
    .A(\atari2600.tia.colupf[1] ));
 sg13g2_inv_1 _16239_ (.Y(_08017_),
    .A(\atari2600.tia.colupf[0] ));
 sg13g2_inv_1 _16240_ (.Y(_08018_),
    .A(net7005));
 sg13g2_inv_1 _16241_ (.Y(_08019_),
    .A(net7135));
 sg13g2_inv_1 _16242_ (.Y(_08020_),
    .A(\atari2600.tia.colup1[4] ));
 sg13g2_inv_1 _16243_ (.Y(_08021_),
    .A(\atari2600.tia.colup1[3] ));
 sg13g2_inv_1 _16244_ (.Y(_08022_),
    .A(net7024));
 sg13g2_inv_1 _16245_ (.Y(_08023_),
    .A(net7058));
 sg13g2_inv_1 _16246_ (.Y(_08024_),
    .A(net6958));
 sg13g2_inv_1 _16247_ (.Y(_08025_),
    .A(net7036));
 sg13g2_inv_1 _16248_ (.Y(_08026_),
    .A(\atari2600.tia.colup0[4] ));
 sg13g2_inv_1 _16249_ (.Y(_08027_),
    .A(\atari2600.tia.colup0[3] ));
 sg13g2_inv_1 _16250_ (.Y(_08028_),
    .A(net6164));
 sg13g2_inv_1 _16251_ (.Y(_08029_),
    .A(net4143));
 sg13g2_inv_1 _16252_ (.Y(_08030_),
    .A(net6905));
 sg13g2_inv_1 _16253_ (.Y(_08031_),
    .A(net7012));
 sg13g2_inv_1 _16254_ (.Y(_08032_),
    .A(\atari2600.tia.audio_right_counter[0] ));
 sg13g2_inv_1 _16255_ (.Y(_08033_),
    .A(\atari2600.tia.audio_left_counter[2] ));
 sg13g2_inv_1 _16256_ (.Y(_08034_),
    .A(net7153));
 sg13g2_inv_1 _16257_ (.Y(_08035_),
    .A(net4400));
 sg13g2_inv_1 _16258_ (.Y(_08036_),
    .A(\atari2600.tia.p0_w[4] ));
 sg13g2_inv_1 _16259_ (.Y(_08037_),
    .A(net5835));
 sg13g2_inv_1 _16260_ (.Y(_08038_),
    .A(net7196));
 sg13g2_inv_1 _16261_ (.Y(_08039_),
    .A(net6323));
 sg13g2_inv_1 _16262_ (.Y(_08040_),
    .A(net2995));
 sg13g2_inv_1 _16263_ (.Y(_08041_),
    .A(net6298));
 sg13g2_inv_1 _16264_ (.Y(_08042_),
    .A(net2895));
 sg13g2_inv_1 _16265_ (.Y(_08043_),
    .A(\atari2600.tia.vid_ypos[5] ));
 sg13g2_inv_2 _16266_ (.Y(_08044_),
    .A(\atari2600.tia.vid_ypos[4] ));
 sg13g2_inv_1 _16267_ (.Y(_08045_),
    .A(\atari2600.tia.vid_ypos[3] ));
 sg13g2_inv_1 _16268_ (.Y(_08046_),
    .A(\atari2600.tia.vid_ypos[2] ));
 sg13g2_inv_1 _16269_ (.Y(_08047_),
    .A(\hvsync_gen.vga.vpos[9] ));
 sg13g2_inv_1 _16270_ (.Y(_08048_),
    .A(\hvsync_gen.vga.vpos[8] ));
 sg13g2_inv_1 _16271_ (.Y(_08049_),
    .A(\hvsync_gen.vga.vpos[3] ));
 sg13g2_inv_1 _16272_ (.Y(_08050_),
    .A(_00078_));
 sg13g2_inv_1 _16273_ (.Y(_08051_),
    .A(net3858));
 sg13g2_inv_1 _16274_ (.Y(_08052_),
    .A(net4191));
 sg13g2_inv_1 _16275_ (.Y(_08053_),
    .A(net3305));
 sg13g2_inv_1 _16276_ (.Y(_08054_),
    .A(net6787));
 sg13g2_inv_1 _16277_ (.Y(_08055_),
    .A(_00081_));
 sg13g2_inv_1 _16278_ (.Y(_08056_),
    .A(net7003));
 sg13g2_inv_1 _16279_ (.Y(_08057_),
    .A(net5571));
 sg13g2_inv_1 _16280_ (.Y(_08058_),
    .A(_00082_));
 sg13g2_inv_1 _16281_ (.Y(_08059_),
    .A(net7197));
 sg13g2_inv_1 _16282_ (.Y(_08060_),
    .A(net3989));
 sg13g2_inv_1 _16283_ (.Y(_08061_),
    .A(\atari2600.cpu.ADD[1] ));
 sg13g2_inv_1 _16284_ (.Y(_08062_),
    .A(\atari2600.cpu.PC[1] ));
 sg13g2_inv_1 _16285_ (.Y(_08063_),
    .A(_00090_));
 sg13g2_inv_1 _16286_ (.Y(_08064_),
    .A(_00089_));
 sg13g2_inv_1 _16287_ (.Y(_08065_),
    .A(_00092_));
 sg13g2_inv_1 _16288_ (.Y(_08066_),
    .A(_00091_));
 sg13g2_inv_1 _16289_ (.Y(_08067_),
    .A(\atari2600.cpu.PC[0] ));
 sg13g2_inv_1 _16290_ (.Y(_08068_),
    .A(\atari2600.cpu.C ));
 sg13g2_inv_1 _16291_ (.Y(_08069_),
    .A(net7146));
 sg13g2_inv_2 _16292_ (.Y(_08070_),
    .A(\atari2600.cpu.ALU.CO ));
 sg13g2_inv_1 _16293_ (.Y(_08071_),
    .A(net7037));
 sg13g2_inv_1 _16294_ (.Y(_08072_),
    .A(net5568));
 sg13g2_inv_1 _16295_ (.Y(_08073_),
    .A(net7132));
 sg13g2_inv_1 _16296_ (.Y(_08074_),
    .A(_00097_));
 sg13g2_inv_1 _16297_ (.Y(_08075_),
    .A(net7137));
 sg13g2_inv_2 _16298_ (.Y(_08076_),
    .A(_00100_));
 sg13g2_inv_1 _16299_ (.Y(_08077_),
    .A(_00102_));
 sg13g2_inv_1 _16300_ (.Y(_08078_),
    .A(net6933));
 sg13g2_inv_1 _16301_ (.Y(_08079_),
    .A(net6723));
 sg13g2_inv_1 _16302_ (.Y(_08080_),
    .A(\atari2600.cpu.PC[7] ));
 sg13g2_inv_1 _16303_ (.Y(_08081_),
    .A(\atari2600.address_bus_r[7] ));
 sg13g2_inv_1 _16304_ (.Y(_08082_),
    .A(net6852));
 sg13g2_inv_1 _16305_ (.Y(_08083_),
    .A(net6984));
 sg13g2_inv_1 _16306_ (.Y(_08084_),
    .A(net7372));
 sg13g2_inv_1 _16307_ (.Y(_08085_),
    .A(net7053));
 sg13g2_inv_1 _16308_ (.Y(_08086_),
    .A(net6953));
 sg13g2_inv_1 _16309_ (.Y(_08087_),
    .A(net6767));
 sg13g2_inv_1 _16310_ (.Y(_08088_),
    .A(\rom_next_addr_in_queue[0] ));
 sg13g2_inv_1 _16311_ (.Y(_08089_),
    .A(net7209));
 sg13g2_inv_1 _16312_ (.Y(_08090_),
    .A(net7242));
 sg13g2_inv_1 _16313_ (.Y(_08091_),
    .A(net7136));
 sg13g2_inv_1 _16314_ (.Y(_08092_),
    .A(net7105));
 sg13g2_inv_1 _16315_ (.Y(_08093_),
    .A(net7086));
 sg13g2_inv_1 _16316_ (.Y(_08094_),
    .A(net7120));
 sg13g2_inv_1 _16317_ (.Y(_08095_),
    .A(net7223));
 sg13g2_inv_1 _16318_ (.Y(_08096_),
    .A(\atari2600.cpu.store ));
 sg13g2_inv_1 _16319_ (.Y(_08097_),
    .A(net6037));
 sg13g2_inv_1 _16320_ (.Y(_08098_),
    .A(_00107_));
 sg13g2_inv_1 _16321_ (.Y(_08099_),
    .A(_00106_));
 sg13g2_inv_1 _16322_ (.Y(_08100_),
    .A(_00112_));
 sg13g2_inv_1 _16323_ (.Y(_08101_),
    .A(_00118_));
 sg13g2_inv_1 _16324_ (.Y(_08102_),
    .A(_00119_));
 sg13g2_inv_1 _16325_ (.Y(_08103_),
    .A(_00122_));
 sg13g2_inv_1 _16326_ (.Y(_08104_),
    .A(_00128_));
 sg13g2_inv_2 _16327_ (.Y(_08105_),
    .A(_00134_));
 sg13g2_inv_1 _16328_ (.Y(_08106_),
    .A(net2892));
 sg13g2_inv_2 _16329_ (.Y(_08107_),
    .A(net5828));
 sg13g2_inv_4 _16330_ (.A(net5829),
    .Y(_08108_));
 sg13g2_inv_2 _16331_ (.Y(_08109_),
    .A(net5821));
 sg13g2_inv_2 _16332_ (.Y(_08110_),
    .A(net5823));
 sg13g2_inv_2 _16333_ (.Y(_08111_),
    .A(net5816));
 sg13g2_inv_1 _16334_ (.Y(_08112_),
    .A(net5811));
 sg13g2_inv_2 _16335_ (.Y(_08113_),
    .A(net5807));
 sg13g2_inv_2 _16336_ (.Y(_08114_),
    .A(net5802));
 sg13g2_inv_1 _16337_ (.Y(_08115_),
    .A(\atari2600.tia.p0_copies[1] ));
 sg13g2_inv_1 _16338_ (.Y(_08116_),
    .A(net3972));
 sg13g2_inv_4 _16339_ (.A(net5842),
    .Y(_08117_));
 sg13g2_inv_1 _16340_ (.Y(_08118_),
    .A(net5848));
 sg13g2_inv_2 _16341_ (.Y(_08119_),
    .A(net5841));
 sg13g2_inv_2 _16342_ (.Y(_08120_),
    .A(net5839));
 sg13g2_inv_1 _16343_ (.Y(_08121_),
    .A(\atari2600.cpu.PC[14] ));
 sg13g2_inv_1 _16344_ (.Y(_08122_),
    .A(_00149_));
 sg13g2_inv_1 _16345_ (.Y(_08123_),
    .A(\atari2600.cpu.PC[15] ));
 sg13g2_inv_1 _16346_ (.Y(_08124_),
    .A(_00150_));
 sg13g2_inv_1 _16347_ (.Y(_08125_),
    .A(net3065));
 sg13g2_inv_1 _16348_ (.Y(_08126_),
    .A(net3409));
 sg13g2_inv_1 _16349_ (.Y(_08127_),
    .A(\atari2600.cpu.cond_code[2] ));
 sg13g2_inv_1 _16350_ (.Y(_08128_),
    .A(net3034));
 sg13g2_inv_1 _16351_ (.Y(_08129_),
    .A(\scanline[40][4] ));
 sg13g2_inv_1 _16352_ (.Y(_08130_),
    .A(\b_pwm_even[1] ));
 sg13g2_nor2_1 _16353_ (.A(\atari2600.clk_counter[7] ),
    .B(\atari2600.clk_counter[6] ),
    .Y(_08131_));
 sg13g2_nor4_2 _16354_ (.A(\atari2600.clk_counter[5] ),
    .B(\atari2600.clk_counter[4] ),
    .C(\atari2600.clk_counter[3] ),
    .Y(_08132_),
    .D(\atari2600.clk_counter[2] ));
 sg13g2_nand3b_1 _16355_ (.B(_08131_),
    .C(_08132_),
    .Y(_08133_),
    .A_N(\atari2600.clk_counter[8] ));
 sg13g2_nor3_2 _16356_ (.A(\atari2600.clk_counter[1] ),
    .B(_07924_),
    .C(_08133_),
    .Y(_08134_));
 sg13g2_inv_1 _16357_ (.Y(_08135_),
    .A(_08134_));
 sg13g2_or2_1 _16358_ (.X(_08136_),
    .B(\atari2600.tia.vid_ypos[0] ),
    .A(\atari2600.tia.vid_ypos[1] ));
 sg13g2_o21ai_1 _16359_ (.B1(\atari2600.tia.vid_ypos[2] ),
    .Y(_08137_),
    .A1(\atari2600.tia.vid_ypos[1] ),
    .A2(\atari2600.tia.vid_ypos[0] ));
 sg13g2_and4_1 _16360_ (.A(\atari2600.tia.vid_ypos[5] ),
    .B(_08044_),
    .C(_08045_),
    .D(_08137_),
    .X(_08138_));
 sg13g2_nor2_1 _16361_ (.A(\atari2600.tia.vid_ypos[7] ),
    .B(\atari2600.tia.vid_ypos[6] ),
    .Y(_08139_));
 sg13g2_o21ai_1 _16362_ (.B1(_08139_),
    .Y(_08140_),
    .A1(_00077_),
    .A2(_08138_));
 sg13g2_a21oi_1 _16363_ (.A1(_08047_),
    .A2(_08140_),
    .Y(_08141_),
    .B1(\atari2600.tia.vid_ypos[8] ));
 sg13g2_nand2_1 _16364_ (.Y(_08142_),
    .A(\atari2600.tia.vid_ypos[7] ),
    .B(_08048_));
 sg13g2_nand2b_1 _16365_ (.Y(_08143_),
    .B(\hvsync_gen.vga.vpos[7] ),
    .A_N(\atari2600.tia.vid_ypos[6] ));
 sg13g2_o21ai_1 _16366_ (.B1(_08143_),
    .Y(_08144_),
    .A1(\atari2600.tia.vid_ypos[7] ),
    .A2(_08048_));
 sg13g2_nand2b_1 _16367_ (.Y(_08145_),
    .B(\hvsync_gen.vga.vpos[2] ),
    .A_N(\atari2600.tia.vid_ypos[1] ));
 sg13g2_nor2b_1 _16368_ (.A(\hvsync_gen.vga.vpos[1] ),
    .B_N(\atari2600.tia.vid_ypos[0] ),
    .Y(_08146_));
 sg13g2_nor2b_1 _16369_ (.A(\hvsync_gen.vga.vpos[2] ),
    .B_N(\atari2600.tia.vid_ypos[1] ),
    .Y(_08147_));
 sg13g2_a221oi_1 _16370_ (.B2(_08146_),
    .C1(_08147_),
    .B1(_08145_),
    .A1(\atari2600.tia.vid_ypos[2] ),
    .Y(_08148_),
    .A2(_08049_));
 sg13g2_a221oi_1 _16371_ (.B2(_08046_),
    .C1(_08148_),
    .B1(\hvsync_gen.vga.vpos[3] ),
    .A1(_08045_),
    .Y(_08149_),
    .A2(\hvsync_gen.vga.vpos[4] ));
 sg13g2_nand2b_1 _16372_ (.Y(_08150_),
    .B(\atari2600.tia.vid_ypos[3] ),
    .A_N(\hvsync_gen.vga.vpos[4] ));
 sg13g2_o21ai_1 _16373_ (.B1(_08150_),
    .Y(_08151_),
    .A1(_08044_),
    .A2(\hvsync_gen.vga.vpos[5] ));
 sg13g2_a22oi_1 _16374_ (.Y(_08152_),
    .B1(\hvsync_gen.vga.vpos[5] ),
    .B2(_08044_),
    .A2(\hvsync_gen.vga.vpos[6] ),
    .A1(_08043_));
 sg13g2_o21ai_1 _16375_ (.B1(_08152_),
    .Y(_08153_),
    .A1(_08149_),
    .A2(_08151_));
 sg13g2_nand2b_1 _16376_ (.Y(_08154_),
    .B(\atari2600.tia.vid_ypos[5] ),
    .A_N(\hvsync_gen.vga.vpos[6] ));
 sg13g2_nand2b_1 _16377_ (.Y(_08155_),
    .B(\atari2600.tia.vid_ypos[6] ),
    .A_N(\hvsync_gen.vga.vpos[7] ));
 sg13g2_and4_1 _16378_ (.A(_08142_),
    .B(_08143_),
    .C(_08154_),
    .D(_08155_),
    .X(_08156_));
 sg13g2_a221oi_1 _16379_ (.B2(_08156_),
    .C1(_08141_),
    .B1(_08153_),
    .A1(_08142_),
    .Y(_08157_),
    .A2(_08144_));
 sg13g2_nor2b_1 _16380_ (.A(\hvsync_gen.vga.vpos[9] ),
    .B_N(\atari2600.tia.vid_ypos[8] ),
    .Y(_08158_));
 sg13g2_a21o_1 _16381_ (.A2(_08134_),
    .A1(rom_data_pending),
    .B1(_08158_),
    .X(_08159_));
 sg13g2_or2_1 _16382_ (.X(_08160_),
    .B(_08159_),
    .A(_08157_));
 sg13g2_inv_1 _16383_ (.Y(_08161_),
    .A(net5385));
 sg13g2_nor2_1 _16384_ (.A(_08135_),
    .B(net5385),
    .Y(_08162_));
 sg13g2_nand2_2 _16385_ (.Y(_08163_),
    .A(_08134_),
    .B(_08161_));
 sg13g2_nor4_2 _16386_ (.A(\atari2600.stall_cpu ),
    .B(_08135_),
    .C(_08157_),
    .Y(_08164_),
    .D(_08159_));
 sg13g2_nand2b_2 _16387_ (.Y(_08165_),
    .B(net5353),
    .A_N(\atari2600.stall_cpu ));
 sg13g2_nor2b_1 _16388_ (.A(net5969),
    .B_N(net5971),
    .Y(_08166_));
 sg13g2_nand2b_1 _16389_ (.Y(_08167_),
    .B(net5972),
    .A_N(net5969));
 sg13g2_nor2b_1 _16390_ (.A(net5975),
    .B_N(net5974),
    .Y(_08168_));
 sg13g2_nand2b_2 _16391_ (.Y(_08169_),
    .B(net5974),
    .A_N(net5975));
 sg13g2_and2_1 _16392_ (.A(\atari2600.cpu.state[2] ),
    .B(\atari2600.cpu.state[3] ),
    .X(_08170_));
 sg13g2_nand2_2 _16393_ (.Y(_08171_),
    .A(\atari2600.cpu.state[2] ),
    .B(\atari2600.cpu.state[3] ));
 sg13g2_nand3_1 _16394_ (.B(_08168_),
    .C(net5548),
    .A(_08166_),
    .Y(_08172_));
 sg13g2_inv_1 _16395_ (.Y(_08173_),
    .A(_08172_));
 sg13g2_mux2_1 _16396_ (.A0(net7362),
    .A1(\atari2600.cpu.DI[5] ),
    .S(net5383),
    .X(\atari2600.cpu.DIMUX[5] ));
 sg13g2_nor2b_1 _16397_ (.A(net5573),
    .B_N(net5351),
    .Y(_08174_));
 sg13g2_a21o_2 _16398_ (.A2(\atari2600.cpu.IRHOLD[5] ),
    .A1(net5573),
    .B1(_08174_),
    .X(_08175_));
 sg13g2_a21oi_1 _16399_ (.A1(net5573),
    .A2(\atari2600.cpu.IRHOLD[5] ),
    .Y(_08176_),
    .B1(_08174_));
 sg13g2_and2_1 _16400_ (.A(net7202),
    .B(net5380),
    .X(_08177_));
 sg13g2_a21o_1 _16401_ (.A2(net5315),
    .A1(net7342),
    .B1(_08177_),
    .X(\atari2600.cpu.DIMUX[7] ));
 sg13g2_nand2b_1 _16402_ (.Y(_08178_),
    .B(net5576),
    .A_N(\atari2600.cpu.IRHOLD[7] ));
 sg13g2_o21ai_1 _16403_ (.B1(_08178_),
    .Y(_08179_),
    .A1(net5576),
    .A2(\atari2600.cpu.DIMUX[7] ));
 sg13g2_nor2b_1 _16404_ (.A(net5383),
    .B_N(\atari2600.cpu.DIHOLD[4] ),
    .Y(_08180_));
 sg13g2_a21oi_2 _16405_ (.B1(_08180_),
    .Y(_08181_),
    .A2(net5382),
    .A1(\atari2600.cpu.DI[4] ));
 sg13g2_inv_2 _16406_ (.Y(\atari2600.cpu.DIMUX[4] ),
    .A(_08181_));
 sg13g2_nor2_1 _16407_ (.A(net5573),
    .B(_08181_),
    .Y(_08182_));
 sg13g2_a21o_2 _16408_ (.A2(\atari2600.cpu.IRHOLD[4] ),
    .A1(net5574),
    .B1(_08182_),
    .X(_08183_));
 sg13g2_a21oi_2 _16409_ (.B1(_08182_),
    .Y(_08184_),
    .A2(\atari2600.cpu.IRHOLD[4] ),
    .A1(net5574));
 sg13g2_and2_2 _16410_ (.A(net5205),
    .B(_08184_),
    .X(_08185_));
 sg13g2_and2_1 _16411_ (.A(_08175_),
    .B(_08185_),
    .X(_08186_));
 sg13g2_mux2_2 _16412_ (.A0(_00087_),
    .A1(net7365),
    .S(net5380),
    .X(_08187_));
 sg13g2_inv_2 _16413_ (.Y(\atari2600.cpu.DIMUX[1] ),
    .A(_08187_));
 sg13g2_nor2_1 _16414_ (.A(net5574),
    .B(_08187_),
    .Y(_08188_));
 sg13g2_a21o_1 _16415_ (.A2(\atari2600.cpu.IRHOLD[1] ),
    .A1(net5574),
    .B1(_08188_),
    .X(_08189_));
 sg13g2_a21oi_2 _16416_ (.B1(_08188_),
    .Y(_08190_),
    .A2(\atari2600.cpu.IRHOLD[1] ),
    .A1(net5573));
 sg13g2_mux2_2 _16417_ (.A0(_00093_),
    .A1(net7347),
    .S(net5382),
    .X(_08191_));
 sg13g2_inv_2 _16418_ (.Y(\atari2600.cpu.DIMUX[0] ),
    .A(net7348));
 sg13g2_nor2_1 _16419_ (.A(net5573),
    .B(_08191_),
    .Y(_08192_));
 sg13g2_a21o_1 _16420_ (.A2(\atari2600.cpu.IRHOLD[0] ),
    .A1(net5573),
    .B1(_08192_),
    .X(_08193_));
 sg13g2_a21oi_2 _16421_ (.B1(_08192_),
    .Y(_08194_),
    .A2(\atari2600.cpu.IRHOLD[0] ),
    .A1(net5573));
 sg13g2_nor2b_1 _16422_ (.A(net5382),
    .B_N(\atari2600.cpu.DIHOLD[3] ),
    .Y(_08195_));
 sg13g2_a21oi_2 _16423_ (.B1(_08195_),
    .Y(_08196_),
    .A2(net5382),
    .A1(\atari2600.cpu.DI[3] ));
 sg13g2_inv_2 _16424_ (.Y(\atari2600.cpu.DIMUX[3] ),
    .A(_08196_));
 sg13g2_nor2_1 _16425_ (.A(net5575),
    .B(_08196_),
    .Y(_08197_));
 sg13g2_a21o_2 _16426_ (.A2(\atari2600.cpu.IRHOLD[3] ),
    .A1(net5575),
    .B1(_08197_),
    .X(_08198_));
 sg13g2_a21oi_2 _16427_ (.B1(_08197_),
    .Y(_08199_),
    .A2(\atari2600.cpu.IRHOLD[3] ),
    .A1(net5575));
 sg13g2_nor2b_1 _16428_ (.A(net5380),
    .B_N(\atari2600.cpu.DIHOLD[2] ),
    .Y(_08200_));
 sg13g2_a21oi_2 _16429_ (.B1(_08200_),
    .Y(_08201_),
    .A2(net5380),
    .A1(\atari2600.cpu.DI[2] ));
 sg13g2_inv_4 _16430_ (.A(_08201_),
    .Y(\atari2600.cpu.DIMUX[2] ));
 sg13g2_nor2_1 _16431_ (.A(net5575),
    .B(_08201_),
    .Y(_08202_));
 sg13g2_a21o_1 _16432_ (.A2(\atari2600.cpu.IRHOLD[2] ),
    .A1(net5575),
    .B1(_08202_),
    .X(_08203_));
 sg13g2_a21oi_2 _16433_ (.B1(_08202_),
    .Y(_08204_),
    .A2(net6917),
    .A1(net5575));
 sg13g2_nor2_2 _16434_ (.A(_08199_),
    .B(_08203_),
    .Y(_08205_));
 sg13g2_nand2_2 _16435_ (.Y(_08206_),
    .A(_08194_),
    .B(_08205_));
 sg13g2_nor2_1 _16436_ (.A(net5971),
    .B(net5970),
    .Y(_08207_));
 sg13g2_or2_1 _16437_ (.X(_08208_),
    .B(net5970),
    .A(net5971));
 sg13g2_nor2_1 _16438_ (.A(net5975),
    .B(net5974),
    .Y(_08209_));
 sg13g2_or2_1 _16439_ (.X(_08210_),
    .B(net5974),
    .A(net5975));
 sg13g2_nor3_2 _16440_ (.A(_08171_),
    .B(net5546),
    .C(_08210_),
    .Y(_08211_));
 sg13g2_nand3_1 _16441_ (.B(net5547),
    .C(net5544),
    .A(net5548),
    .Y(_08212_));
 sg13g2_nor2_1 _16442_ (.A(net5312),
    .B(_08212_),
    .Y(_08213_));
 sg13g2_nand2_1 _16443_ (.Y(_08214_),
    .A(net5363),
    .B(net5480));
 sg13g2_nand2_2 _16444_ (.Y(_08215_),
    .A(_08190_),
    .B(_08194_));
 sg13g2_nor2_2 _16445_ (.A(_08189_),
    .B(_08206_),
    .Y(_08216_));
 sg13g2_nand3_1 _16446_ (.B(_08194_),
    .C(_08205_),
    .A(_08190_),
    .Y(_08217_));
 sg13g2_nor2_1 _16447_ (.A(net5349),
    .B(_08217_),
    .Y(_08218_));
 sg13g2_nand2_1 _16448_ (.Y(_08219_),
    .A(net5271),
    .B(_08216_));
 sg13g2_a22oi_1 _16449_ (.Y(_08220_),
    .B1(_08186_),
    .B2(_08218_),
    .A2(_08173_),
    .A1(net5310));
 sg13g2_nor2_1 _16450_ (.A(_08183_),
    .B(net5350),
    .Y(_08221_));
 sg13g2_nor2_1 _16451_ (.A(_08189_),
    .B(_08194_),
    .Y(_08222_));
 sg13g2_nor2_2 _16452_ (.A(_08198_),
    .B(net5202),
    .Y(_08223_));
 sg13g2_nand3_1 _16453_ (.B(net5200),
    .C(_08223_),
    .A(_08221_),
    .Y(_08224_));
 sg13g2_nor2b_1 _16454_ (.A(net5971),
    .B_N(net5970),
    .Y(_08225_));
 sg13g2_nand2b_1 _16455_ (.Y(_08226_),
    .B(net5969),
    .A_N(net5971));
 sg13g2_nor2_2 _16456_ (.A(\atari2600.cpu.state[2] ),
    .B(net5973),
    .Y(_08227_));
 sg13g2_and2_1 _16457_ (.A(net5975),
    .B(net5974),
    .X(_08228_));
 sg13g2_nand2_1 _16458_ (.Y(_08229_),
    .A(net5975),
    .B(\atari2600.cpu.state[1] ));
 sg13g2_nand3_1 _16459_ (.B(net5540),
    .C(net5539),
    .A(net5543),
    .Y(_08230_));
 sg13g2_nor3_2 _16460_ (.A(_08169_),
    .B(_08171_),
    .C(net5541),
    .Y(_08231_));
 sg13g2_nand3_1 _16461_ (.B(net5548),
    .C(net5542),
    .A(net5549),
    .Y(_08232_));
 sg13g2_nor2_1 _16462_ (.A(net5368),
    .B(net5479),
    .Y(_08233_));
 sg13g2_a21oi_1 _16463_ (.A1(net5369),
    .A2(_08230_),
    .Y(_08234_),
    .B1(_08233_));
 sg13g2_nand3_1 _16464_ (.B(_08170_),
    .C(_08207_),
    .A(_08168_),
    .Y(_08235_));
 sg13g2_nor2_1 _16465_ (.A(net5375),
    .B(_08235_),
    .Y(_08236_));
 sg13g2_nor2_1 _16466_ (.A(_08234_),
    .B(_08236_),
    .Y(_08237_));
 sg13g2_nand3_1 _16467_ (.B(_08224_),
    .C(_08237_),
    .A(_08220_),
    .Y(_08238_));
 sg13g2_nor2b_2 _16468_ (.A(\atari2600.cpu.state[2] ),
    .B_N(net5973),
    .Y(_08239_));
 sg13g2_nand2b_2 _16469_ (.Y(_08240_),
    .B(net5973),
    .A_N(\atari2600.cpu.state[2] ));
 sg13g2_nor3_2 _16470_ (.A(_08167_),
    .B(_08210_),
    .C(_08240_),
    .Y(_08241_));
 sg13g2_nor3_2 _16471_ (.A(_08199_),
    .B(_08204_),
    .C(_08215_),
    .Y(_08242_));
 sg13g2_nor2b_1 _16472_ (.A(net5382),
    .B_N(\atari2600.cpu.DIHOLD[6] ),
    .Y(_08243_));
 sg13g2_a21oi_2 _16473_ (.B1(_08243_),
    .Y(_08244_),
    .A2(net5382),
    .A1(\atari2600.cpu.DI[6] ));
 sg13g2_inv_2 _16474_ (.Y(\atari2600.cpu.DIMUX[6] ),
    .A(_08244_));
 sg13g2_nor2_1 _16475_ (.A(net5576),
    .B(_08244_),
    .Y(_08245_));
 sg13g2_a21o_2 _16476_ (.A2(\atari2600.cpu.IRHOLD[6] ),
    .A1(net5576),
    .B1(_08245_),
    .X(_08246_));
 sg13g2_a21oi_2 _16477_ (.B1(_08245_),
    .Y(_08247_),
    .A2(\atari2600.cpu.IRHOLD[6] ),
    .A1(net5576));
 sg13g2_nor2_2 _16478_ (.A(net5274),
    .B(net5199),
    .Y(_08248_));
 sg13g2_and4_1 _16479_ (.A(_08185_),
    .B(net5272),
    .C(_08242_),
    .D(_08248_),
    .X(_08249_));
 sg13g2_a21oi_1 _16480_ (.A1(net5310),
    .A2(_08241_),
    .Y(_08250_),
    .B1(_08249_));
 sg13g2_nand3_1 _16481_ (.B(net5542),
    .C(_08239_),
    .A(net5549),
    .Y(_08251_));
 sg13g2_nor3_2 _16482_ (.A(_08198_),
    .B(net5202),
    .C(_08215_),
    .Y(_08252_));
 sg13g2_nand2_1 _16483_ (.Y(_08253_),
    .A(net5272),
    .B(_08252_));
 sg13g2_nand4_1 _16484_ (.B(net5272),
    .C(_08246_),
    .A(_08186_),
    .Y(_08254_),
    .D(_08252_));
 sg13g2_o21ai_1 _16485_ (.B1(_08254_),
    .Y(_08255_),
    .A1(net5378),
    .A2(_08251_));
 sg13g2_nor3_2 _16486_ (.A(net5550),
    .B(_08169_),
    .C(_08240_),
    .Y(_08256_));
 sg13g2_nand3_1 _16487_ (.B(net5549),
    .C(_08239_),
    .A(net5551),
    .Y(_08257_));
 sg13g2_nand2_1 _16488_ (.Y(_08258_),
    .A(net5310),
    .B(_08256_));
 sg13g2_nand2_2 _16489_ (.Y(_08259_),
    .A(_08186_),
    .B(net5199));
 sg13g2_o21ai_1 _16490_ (.B1(_08258_),
    .Y(_08260_),
    .A1(_08253_),
    .A2(_08259_));
 sg13g2_nor2_1 _16491_ (.A(_08255_),
    .B(_08260_),
    .Y(_08261_));
 sg13g2_nor2_1 _16492_ (.A(net5205),
    .B(_08193_),
    .Y(_08262_));
 sg13g2_a22oi_1 _16493_ (.Y(_08263_),
    .B1(_08223_),
    .B2(_08262_),
    .A2(net5200),
    .A1(_08205_));
 sg13g2_nor2b_1 _16494_ (.A(_08263_),
    .B_N(_08221_),
    .Y(_08264_));
 sg13g2_nand3_1 _16495_ (.B(net5544),
    .C(net5542),
    .A(_08170_),
    .Y(_08265_));
 sg13g2_nor2b_2 _16496_ (.A(net5974),
    .B_N(net5975),
    .Y(_08266_));
 sg13g2_nand2b_2 _16497_ (.Y(_08267_),
    .B(net5975),
    .A_N(net5974));
 sg13g2_nor2_1 _16498_ (.A(_08171_),
    .B(_08267_),
    .Y(_08268_));
 sg13g2_nand2_1 _16499_ (.Y(_08269_),
    .A(net5548),
    .B(_08266_));
 sg13g2_nor2_1 _16500_ (.A(net5971),
    .B(_08269_),
    .Y(_08270_));
 sg13g2_a21oi_1 _16501_ (.A1(net5970),
    .A2(_08270_),
    .Y(_08271_),
    .B1(net5374));
 sg13g2_a21oi_1 _16502_ (.A1(net5374),
    .A2(_08265_),
    .Y(_08272_),
    .B1(_08271_));
 sg13g2_nand3_1 _16503_ (.B(net5548),
    .C(net5544),
    .A(net5551),
    .Y(_08273_));
 sg13g2_a21oi_1 _16504_ (.A1(net5551),
    .A2(_08268_),
    .Y(_08274_),
    .B1(net5379));
 sg13g2_a21oi_1 _16505_ (.A1(net5370),
    .A2(_08273_),
    .Y(_08275_),
    .B1(_08274_));
 sg13g2_nor2_2 _16506_ (.A(net5546),
    .B(_08269_),
    .Y(_08276_));
 sg13g2_nor2b_1 _16507_ (.A(net5973),
    .B_N(\atari2600.cpu.state[2] ),
    .Y(_08277_));
 sg13g2_and2_1 _16508_ (.A(net5544),
    .B(net5538),
    .X(_08278_));
 sg13g2_nand2_2 _16509_ (.Y(_08279_),
    .A(net5544),
    .B(net5538));
 sg13g2_nor2_2 _16510_ (.A(net5545),
    .B(_08279_),
    .Y(_08280_));
 sg13g2_nand2_2 _16511_ (.Y(_08281_),
    .A(_08227_),
    .B(_08266_));
 sg13g2_and4_1 _16512_ (.A(net5971),
    .B(net5969),
    .C(net5540),
    .D(_08266_),
    .X(_08282_));
 sg13g2_nor2_2 _16513_ (.A(net5546),
    .B(_08281_),
    .Y(_08283_));
 sg13g2_nand2_1 _16514_ (.Y(_08284_),
    .A(net5548),
    .B(_08228_));
 sg13g2_nor2_1 _16515_ (.A(_08226_),
    .B(_08284_),
    .Y(_08285_));
 sg13g2_nand3_1 _16516_ (.B(net5543),
    .C(net5539),
    .A(net5548),
    .Y(_08286_));
 sg13g2_or4_2 _16517_ (.A(_08280_),
    .B(_08282_),
    .C(_08283_),
    .D(_08285_),
    .X(_08287_));
 sg13g2_o21ai_1 _16518_ (.B1(_08268_),
    .Y(_08288_),
    .A1(net5551),
    .A2(net5542));
 sg13g2_nand3_1 _16519_ (.B(net5540),
    .C(net5539),
    .A(net5547),
    .Y(_08289_));
 sg13g2_nor3_1 _16520_ (.A(\atari2600.cpu.ALU.CO ),
    .B(\atari2600.cpu.store ),
    .C(\atari2600.cpu.write_back ),
    .Y(_08290_));
 sg13g2_nor2b_1 _16521_ (.A(_08289_),
    .B_N(_08290_),
    .Y(_08291_));
 sg13g2_nand2_2 _16522_ (.Y(_08292_),
    .A(net5551),
    .B(_08278_));
 sg13g2_nor3_1 _16523_ (.A(\atari2600.cpu.ALU.CO ),
    .B(\atari2600.cpu.store ),
    .C(_08292_),
    .Y(_08293_));
 sg13g2_nand2_2 _16524_ (.Y(_08294_),
    .A(_08266_),
    .B(net5538));
 sg13g2_nand3_1 _16525_ (.B(_08266_),
    .C(_08277_),
    .A(_08166_),
    .Y(_08295_));
 sg13g2_nor3_1 _16526_ (.A(net5973),
    .B(net5550),
    .C(_08267_),
    .Y(_08296_));
 sg13g2_nor3_1 _16527_ (.A(_08291_),
    .B(_08293_),
    .C(_08296_),
    .Y(_08297_));
 sg13g2_nand3_1 _16528_ (.B(_08288_),
    .C(_08297_),
    .A(_08232_),
    .Y(_08298_));
 sg13g2_a21oi_1 _16529_ (.A1(_00141_),
    .A2(_08287_),
    .Y(_08299_),
    .B1(_08298_));
 sg13g2_nor2_1 _16530_ (.A(net5384),
    .B(_08276_),
    .Y(_08300_));
 sg13g2_a21oi_1 _16531_ (.A1(net5372),
    .A2(_08299_),
    .Y(_08301_),
    .B1(_08300_));
 sg13g2_or4_1 _16532_ (.A(_08264_),
    .B(_08272_),
    .C(_08275_),
    .D(_08301_),
    .X(_08302_));
 sg13g2_nor2_1 _16533_ (.A(_08198_),
    .B(_08204_),
    .Y(_08303_));
 sg13g2_a22oi_1 _16534_ (.Y(_08304_),
    .B1(_08303_),
    .B2(_08221_),
    .A2(_08285_),
    .A1(_08165_));
 sg13g2_nor2_2 _16535_ (.A(net5546),
    .B(_08284_),
    .Y(_08305_));
 sg13g2_nand2_1 _16536_ (.Y(_08306_),
    .A(net5377),
    .B(_08235_));
 sg13g2_o21ai_1 _16537_ (.B1(_08306_),
    .Y(_08307_),
    .A1(net5377),
    .A2(_08305_));
 sg13g2_nand2_1 _16538_ (.Y(_08308_),
    .A(_08304_),
    .B(_08307_));
 sg13g2_nand2_1 _16539_ (.Y(_08309_),
    .A(net5539),
    .B(_08239_));
 sg13g2_nor2_1 _16540_ (.A(net5545),
    .B(_08309_),
    .Y(_08310_));
 sg13g2_nand3_1 _16541_ (.B(net5539),
    .C(_08239_),
    .A(net5547),
    .Y(_08311_));
 sg13g2_nor2_1 _16542_ (.A(net5368),
    .B(_08310_),
    .Y(_08312_));
 sg13g2_nor3_2 _16543_ (.A(_08169_),
    .B(net5545),
    .C(_08240_),
    .Y(_08313_));
 sg13g2_nand3_1 _16544_ (.B(net5547),
    .C(_08239_),
    .A(net5549),
    .Y(_08314_));
 sg13g2_a21oi_1 _16545_ (.A1(net5368),
    .A2(net5475),
    .Y(_08315_),
    .B1(_08312_));
 sg13g2_nor2_2 _16546_ (.A(net5541),
    .B(_08309_),
    .Y(_08316_));
 sg13g2_nor2_1 _16547_ (.A(net5368),
    .B(_08316_),
    .Y(_08317_));
 sg13g2_a21oi_1 _16548_ (.A1(net5368),
    .A2(_08251_),
    .Y(_08318_),
    .B1(_08317_));
 sg13g2_nor2_1 _16549_ (.A(net5550),
    .B(_08309_),
    .Y(_08319_));
 sg13g2_nor2_1 _16550_ (.A(net5370),
    .B(_08319_),
    .Y(_08320_));
 sg13g2_a21oi_1 _16551_ (.A1(net5379),
    .A2(net5477),
    .Y(_08321_),
    .B1(_08320_));
 sg13g2_nor3_1 _16552_ (.A(_08315_),
    .B(_08318_),
    .C(_08321_),
    .Y(_08322_));
 sg13g2_nand3_1 _16553_ (.B(net5542),
    .C(_08239_),
    .A(net5544),
    .Y(_08323_));
 sg13g2_nor3_2 _16554_ (.A(net5541),
    .B(_08240_),
    .C(_08267_),
    .Y(_08324_));
 sg13g2_nor2_1 _16555_ (.A(net5374),
    .B(_08324_),
    .Y(_08325_));
 sg13g2_a21oi_2 _16556_ (.B1(_08325_),
    .Y(_08326_),
    .A2(_08323_),
    .A1(net5374));
 sg13g2_nor3_2 _16557_ (.A(net5550),
    .B(_08240_),
    .C(_08267_),
    .Y(_08327_));
 sg13g2_mux2_1 _16558_ (.A0(_08327_),
    .A1(_08241_),
    .S(net5378),
    .X(_08328_));
 sg13g2_nor3_2 _16559_ (.A(net5545),
    .B(_08240_),
    .C(_08267_),
    .Y(_08329_));
 sg13g2_nor2b_1 _16560_ (.A(net5369),
    .B_N(_08329_),
    .Y(_08330_));
 sg13g2_nand3_1 _16561_ (.B(net5544),
    .C(_08239_),
    .A(net5547),
    .Y(_08331_));
 sg13g2_nor2_2 _16562_ (.A(net5311),
    .B(_08331_),
    .Y(_08332_));
 sg13g2_nor4_2 _16563_ (.A(_08326_),
    .B(_08328_),
    .C(_08330_),
    .Y(_08333_),
    .D(_08332_));
 sg13g2_nand2_2 _16564_ (.Y(_08334_),
    .A(net5539),
    .B(net5538));
 sg13g2_nor2_2 _16565_ (.A(net5541),
    .B(_08334_),
    .Y(_08335_));
 sg13g2_nand3_1 _16566_ (.B(net5539),
    .C(net5538),
    .A(net5542),
    .Y(_08336_));
 sg13g2_nand2_1 _16567_ (.Y(_08337_),
    .A(net5369),
    .B(net5445));
 sg13g2_o21ai_1 _16568_ (.B1(_08337_),
    .Y(_08338_),
    .A1(net5375),
    .A2(_08323_));
 sg13g2_nor2_1 _16569_ (.A(net5311),
    .B(_08329_),
    .Y(_08339_));
 sg13g2_a21oi_1 _16570_ (.A1(net5310),
    .A2(net5475),
    .Y(_08340_),
    .B1(_08339_));
 sg13g2_nand3_1 _16571_ (.B(net5548),
    .C(_08228_),
    .A(net5551),
    .Y(_08341_));
 sg13g2_nor2b_1 _16572_ (.A(net5374),
    .B_N(_08341_),
    .Y(_08342_));
 sg13g2_a21oi_1 _16573_ (.A1(net5374),
    .A2(_08172_),
    .Y(_08343_),
    .B1(_08342_));
 sg13g2_nor3_1 _16574_ (.A(_08338_),
    .B(_08340_),
    .C(_08343_),
    .Y(_08344_));
 sg13g2_nand3_1 _16575_ (.B(_08333_),
    .C(_08344_),
    .A(_08322_),
    .Y(_08345_));
 sg13g2_nor3_1 _16576_ (.A(_08302_),
    .B(_08308_),
    .C(_08345_),
    .Y(_08346_));
 sg13g2_nand3_1 _16577_ (.B(_08261_),
    .C(_08346_),
    .A(_08250_),
    .Y(_08347_));
 sg13g2_and2_1 _16578_ (.A(net5549),
    .B(net5538),
    .X(_08348_));
 sg13g2_nand2_2 _16579_ (.Y(_08349_),
    .A(net5551),
    .B(_08348_));
 sg13g2_nand2_1 _16580_ (.Y(_08350_),
    .A(net5274),
    .B(_08185_));
 sg13g2_nand4_1 _16581_ (.B(_08185_),
    .C(_08242_),
    .A(net5274),
    .Y(_08351_),
    .D(_08246_));
 sg13g2_nor2_1 _16582_ (.A(_08212_),
    .B(_08351_),
    .Y(_08352_));
 sg13g2_nor4_1 _16583_ (.A(net5310),
    .B(_08310_),
    .C(_08327_),
    .D(_08352_),
    .Y(_08353_));
 sg13g2_a21oi_2 _16584_ (.B1(_08353_),
    .Y(_08354_),
    .A2(_08349_),
    .A1(net5310));
 sg13g2_inv_1 _16585_ (.Y(_08355_),
    .A(_08354_));
 sg13g2_nor2_1 _16586_ (.A(net5541),
    .B(_08294_),
    .Y(_08356_));
 sg13g2_nand3_1 _16587_ (.B(_08266_),
    .C(net5538),
    .A(net5543),
    .Y(_08357_));
 sg13g2_nand2_2 _16588_ (.Y(_08358_),
    .A(net5543),
    .B(_08348_));
 sg13g2_nand2_1 _16589_ (.Y(_08359_),
    .A(net5375),
    .B(_08356_));
 sg13g2_o21ai_1 _16590_ (.B1(_08359_),
    .Y(_08360_),
    .A1(net5375),
    .A2(_08358_));
 sg13g2_and2_1 _16591_ (.A(net5547),
    .B(_08348_),
    .X(_08361_));
 sg13g2_nand2_1 _16592_ (.Y(_08362_),
    .A(net5547),
    .B(_08348_));
 sg13g2_nor2_1 _16593_ (.A(net5545),
    .B(_08294_),
    .Y(_08363_));
 sg13g2_nand2_1 _16594_ (.Y(_08364_),
    .A(\atari2600.cpu.Z ),
    .B(\atari2600.cpu.cond_code[1] ));
 sg13g2_o21ai_1 _16595_ (.B1(_08364_),
    .Y(_08365_),
    .A1(_08068_),
    .A2(\atari2600.cpu.cond_code[1] ));
 sg13g2_nand2_1 _16596_ (.Y(_08366_),
    .A(\atari2600.cpu.cond_code[2] ),
    .B(_08365_));
 sg13g2_nor2b_1 _16597_ (.A(\atari2600.cpu.V ),
    .B_N(\atari2600.cpu.cond_code[1] ),
    .Y(_08367_));
 sg13g2_o21ai_1 _16598_ (.B1(_00058_),
    .Y(_08368_),
    .A1(_08122_),
    .A2(\atari2600.cpu.cond_code[1] ));
 sg13g2_o21ai_1 _16599_ (.B1(_08366_),
    .Y(_08369_),
    .A1(_08367_),
    .A2(_08368_));
 sg13g2_nor2_1 _16600_ (.A(_08127_),
    .B(_08365_),
    .Y(_08370_));
 sg13g2_a21oi_1 _16601_ (.A1(_00058_),
    .A2(_08367_),
    .Y(_08371_),
    .B1(_08370_));
 sg13g2_nor2_1 _16602_ (.A(\atari2600.cpu.cond_code[0] ),
    .B(_08371_),
    .Y(_08372_));
 sg13g2_o21ai_1 _16603_ (.B1(_00058_),
    .Y(_08373_),
    .A1(\atari2600.cpu.cond_code[1] ),
    .A2(\atari2600.cpu.cond_code[0] ));
 sg13g2_nor2_1 _16604_ (.A(\atari2600.cpu.N ),
    .B(\atari2600.cpu.cond_code[2] ),
    .Y(_08374_));
 sg13g2_a221oi_1 _16605_ (.B2(_08374_),
    .C1(_08372_),
    .B1(_08373_),
    .A1(\atari2600.cpu.cond_code[0] ),
    .Y(_08375_),
    .A2(_08369_));
 sg13g2_nand3b_1 _16606_ (.B(net5437),
    .C(net5363),
    .Y(_08376_),
    .A_N(_08375_));
 sg13g2_o21ai_1 _16607_ (.B1(_08376_),
    .Y(_08377_),
    .A1(net5372),
    .A2(net5440));
 sg13g2_nor4_2 _16608_ (.A(_08238_),
    .B(_08354_),
    .C(_08360_),
    .Y(_08378_),
    .D(_08377_));
 sg13g2_nand2_2 _16609_ (.Y(_08379_),
    .A(net5549),
    .B(net5540));
 sg13g2_nand3_1 _16610_ (.B(net5549),
    .C(_08227_),
    .A(net5551),
    .Y(_08380_));
 sg13g2_inv_1 _16611_ (.Y(_08381_),
    .A(_08380_));
 sg13g2_nor2_2 _16612_ (.A(net5203),
    .B(net5347),
    .Y(_08382_));
 sg13g2_nand3_1 _16613_ (.B(_08223_),
    .C(_08382_),
    .A(net5200),
    .Y(_08383_));
 sg13g2_o21ai_1 _16614_ (.B1(_08383_),
    .Y(_08384_),
    .A1(net5378),
    .A2(_08380_));
 sg13g2_nor2_1 _16615_ (.A(net5202),
    .B(net5200),
    .Y(_08385_));
 sg13g2_nor4_1 _16616_ (.A(net5203),
    .B(_08199_),
    .C(net5350),
    .D(_08385_),
    .Y(_08386_));
 sg13g2_nand3_1 _16617_ (.B(net5540),
    .C(_08266_),
    .A(net5542),
    .Y(_08387_));
 sg13g2_nand2_1 _16618_ (.Y(_08388_),
    .A(net5372),
    .B(_08387_));
 sg13g2_nor2_2 _16619_ (.A(net5541),
    .B(_08379_),
    .Y(_08389_));
 sg13g2_o21ai_1 _16620_ (.B1(_08388_),
    .Y(_08390_),
    .A1(net5368),
    .A2(net5436));
 sg13g2_nor2_1 _16621_ (.A(net5545),
    .B(_08379_),
    .Y(_08391_));
 sg13g2_nand3_1 _16622_ (.B(_08207_),
    .C(net5540),
    .A(net5549),
    .Y(_08392_));
 sg13g2_o21ai_1 _16623_ (.B1(_08390_),
    .Y(_08393_),
    .A1(_08339_),
    .A2(_08392_));
 sg13g2_nor4_1 _16624_ (.A(_08340_),
    .B(_08384_),
    .C(_08386_),
    .D(_08393_),
    .Y(_08394_));
 sg13g2_nand3_1 _16625_ (.B(_08378_),
    .C(_08394_),
    .A(_08261_),
    .Y(_08395_));
 sg13g2_inv_1 _16626_ (.Y(_08396_),
    .A(_08395_));
 sg13g2_nor3_1 _16627_ (.A(net5199),
    .B(_08253_),
    .C(_08350_),
    .Y(_08397_));
 sg13g2_a21oi_1 _16628_ (.A1(net5310),
    .A2(_08356_),
    .Y(_08398_),
    .B1(_08397_));
 sg13g2_a21oi_1 _16629_ (.A1(_08070_),
    .A2(_08096_),
    .Y(_08399_),
    .B1(_08292_));
 sg13g2_nor2_1 _16630_ (.A(net5379),
    .B(_08295_),
    .Y(_08400_));
 sg13g2_a21oi_1 _16631_ (.A1(net5371),
    .A2(_08399_),
    .Y(_08401_),
    .B1(_08400_));
 sg13g2_nand2_1 _16632_ (.Y(_08402_),
    .A(_08398_),
    .B(_08401_));
 sg13g2_nor2_1 _16633_ (.A(_08302_),
    .B(_08402_),
    .Y(_08403_));
 sg13g2_nor2_1 _16634_ (.A(net5373),
    .B(_08387_),
    .Y(_08404_));
 sg13g2_nor2_2 _16635_ (.A(_08217_),
    .B(_08350_),
    .Y(_08405_));
 sg13g2_a21oi_2 _16636_ (.B1(_08404_),
    .Y(_08406_),
    .A2(_08405_),
    .A1(net5272));
 sg13g2_nor2_1 _16637_ (.A(net5550),
    .B(_08334_),
    .Y(_08407_));
 sg13g2_nor2_1 _16638_ (.A(net5370),
    .B(_08407_),
    .Y(_08408_));
 sg13g2_a21oi_1 _16639_ (.A1(net5370),
    .A2(_08349_),
    .Y(_08409_),
    .B1(_08408_));
 sg13g2_nor2_1 _16640_ (.A(_08343_),
    .B(_08409_),
    .Y(_08410_));
 sg13g2_nand2_1 _16641_ (.Y(_08411_),
    .A(net5368),
    .B(_08358_));
 sg13g2_o21ai_1 _16642_ (.B1(_08411_),
    .Y(_08412_),
    .A1(net5368),
    .A2(net5445));
 sg13g2_nor2_1 _16643_ (.A(net5545),
    .B(_08334_),
    .Y(_08413_));
 sg13g2_nand3_1 _16644_ (.B(net5539),
    .C(net5538),
    .A(net5547),
    .Y(_08414_));
 sg13g2_xnor2_1 _16645_ (.Y(_08415_),
    .A(\atari2600.cpu.backwards ),
    .B(\atari2600.cpu.ALU.CO ));
 sg13g2_o21ai_1 _16646_ (.B1(net5372),
    .Y(_08416_),
    .A1(net5440),
    .A2(_08415_));
 sg13g2_o21ai_1 _16647_ (.B1(_08416_),
    .Y(_08417_),
    .A1(net5372),
    .A2(net5435));
 sg13g2_nand3_1 _16648_ (.B(_08412_),
    .C(_08417_),
    .A(_08410_),
    .Y(_08418_));
 sg13g2_or2_1 _16649_ (.X(_08419_),
    .B(_08418_),
    .A(_08308_));
 sg13g2_nor2_1 _16650_ (.A(net5371),
    .B(_08289_),
    .Y(_08420_));
 sg13g2_a21oi_1 _16651_ (.A1(net5371),
    .A2(_08391_),
    .Y(_08421_),
    .B1(_08420_));
 sg13g2_nand2_1 _16652_ (.Y(_08422_),
    .A(net5376),
    .B(_08380_));
 sg13g2_nor4_2 _16653_ (.A(\atari2600.cpu.state[2] ),
    .B(net5973),
    .C(net5550),
    .Y(_08423_),
    .D(_08229_));
 sg13g2_nand3_1 _16654_ (.B(_08227_),
    .C(_08228_),
    .A(_08166_),
    .Y(_08424_));
 sg13g2_o21ai_1 _16655_ (.B1(_08422_),
    .Y(_08425_),
    .A1(net5377),
    .A2(_08423_));
 sg13g2_nor2b_1 _16656_ (.A(_00141_),
    .B_N(_08287_),
    .Y(_08426_));
 sg13g2_nor2_1 _16657_ (.A(net5372),
    .B(_08230_),
    .Y(_08427_));
 sg13g2_a21oi_2 _16658_ (.B1(_08427_),
    .Y(_08428_),
    .A2(_08426_),
    .A1(net5372));
 sg13g2_nand4_1 _16659_ (.B(_08421_),
    .C(_08425_),
    .A(_08322_),
    .Y(_08429_),
    .D(_08428_));
 sg13g2_nor2_1 _16660_ (.A(_08419_),
    .B(_08429_),
    .Y(_08430_));
 sg13g2_nand2_2 _16661_ (.Y(_08431_),
    .A(net5544),
    .B(net5540));
 sg13g2_nand4_1 _16662_ (.B(net5969),
    .C(_08209_),
    .A(net5972),
    .Y(_08432_),
    .D(net5540));
 sg13g2_inv_1 _16663_ (.Y(_08433_),
    .A(_08432_));
 sg13g2_nor2_1 _16664_ (.A(net5376),
    .B(_08282_),
    .Y(_08434_));
 sg13g2_a21oi_1 _16665_ (.A1(net5376),
    .A2(_08432_),
    .Y(_08435_),
    .B1(_08434_));
 sg13g2_nor3_1 _16666_ (.A(net5376),
    .B(net5550),
    .C(_08281_),
    .Y(_08436_));
 sg13g2_nor2_1 _16667_ (.A(net5550),
    .B(_08431_),
    .Y(_08437_));
 sg13g2_and2_1 _16668_ (.A(net5377),
    .B(_08437_),
    .X(_08438_));
 sg13g2_nor3_1 _16669_ (.A(_08435_),
    .B(_08436_),
    .C(_08438_),
    .Y(_08439_));
 sg13g2_nor2_1 _16670_ (.A(net5546),
    .B(_08431_),
    .Y(_08440_));
 sg13g2_nand2b_1 _16671_ (.Y(_08441_),
    .B(net5376),
    .A_N(_08440_));
 sg13g2_o21ai_1 _16672_ (.B1(_08441_),
    .Y(_08442_),
    .A1(net5376),
    .A2(_08283_));
 sg13g2_nand4_1 _16673_ (.B(_08406_),
    .C(_08439_),
    .A(_08333_),
    .Y(_08443_),
    .D(_08442_));
 sg13g2_a221oi_1 _16674_ (.B2(_08252_),
    .C1(_08443_),
    .B1(_08382_),
    .A1(_08165_),
    .Y(_08444_),
    .A2(net5437));
 sg13g2_nand3_1 _16675_ (.B(_08430_),
    .C(_08444_),
    .A(_08403_),
    .Y(_00173_));
 sg13g2_nand2_1 _16676_ (.Y(_08445_),
    .A(net5203),
    .B(_08198_));
 sg13g2_nor2_2 _16677_ (.A(_08190_),
    .B(_08193_),
    .Y(_08446_));
 sg13g2_nand2_2 _16678_ (.Y(_08447_),
    .A(net5202),
    .B(_08446_));
 sg13g2_o21ai_1 _16679_ (.B1(net5202),
    .Y(_08448_),
    .A1(net5201),
    .A2(_08262_));
 sg13g2_a21oi_1 _16680_ (.A1(_08447_),
    .A2(_08448_),
    .Y(_08449_),
    .B1(_08445_));
 sg13g2_nor3_2 _16681_ (.A(_08204_),
    .B(_08215_),
    .C(_08259_),
    .Y(_08450_));
 sg13g2_a21oi_1 _16682_ (.A1(_08198_),
    .A2(_08450_),
    .Y(_08451_),
    .B1(_08449_));
 sg13g2_nor2_2 _16683_ (.A(net5541),
    .B(_08279_),
    .Y(_08452_));
 sg13g2_nand2_2 _16684_ (.Y(_08453_),
    .A(net5542),
    .B(_08278_));
 sg13g2_nand2_1 _16685_ (.Y(_08454_),
    .A(_08205_),
    .B(_08446_));
 sg13g2_a21oi_1 _16686_ (.A1(_08185_),
    .A2(_08190_),
    .Y(_08455_),
    .B1(_08206_));
 sg13g2_a22oi_1 _16687_ (.Y(_08456_),
    .B1(_08455_),
    .B2(_08213_),
    .A2(_08452_),
    .A1(net5310));
 sg13g2_nor2_1 _16688_ (.A(net5370),
    .B(_08292_),
    .Y(_08457_));
 sg13g2_a21oi_1 _16689_ (.A1(net5375),
    .A2(_08423_),
    .Y(_08458_),
    .B1(_08457_));
 sg13g2_o21ai_1 _16690_ (.B1(net5372),
    .Y(_08459_),
    .A1(_08289_),
    .A2(_08290_));
 sg13g2_o21ai_1 _16691_ (.B1(_08459_),
    .Y(_08460_),
    .A1(net5369),
    .A2(_08280_));
 sg13g2_nand3_1 _16692_ (.B(_08458_),
    .C(_08460_),
    .A(_08456_),
    .Y(_08461_));
 sg13g2_a22oi_1 _16693_ (.Y(_08462_),
    .B1(_08433_),
    .B2(_08165_),
    .A2(_08382_),
    .A1(_08303_));
 sg13g2_nor2b_1 _16694_ (.A(net5376),
    .B_N(_08437_),
    .Y(_08463_));
 sg13g2_a21oi_1 _16695_ (.A1(net5377),
    .A2(_08305_),
    .Y(_08464_),
    .B1(_08463_));
 sg13g2_nand2_1 _16696_ (.Y(_08465_),
    .A(_08462_),
    .B(_08464_));
 sg13g2_nor2_2 _16697_ (.A(net5541),
    .B(_08431_),
    .Y(_08466_));
 sg13g2_nor2_1 _16698_ (.A(net5374),
    .B(_08466_),
    .Y(_08467_));
 sg13g2_a21oi_1 _16699_ (.A1(net5375),
    .A2(_08341_),
    .Y(_08468_),
    .B1(_08467_));
 sg13g2_nor4_1 _16700_ (.A(net5972),
    .B(net5969),
    .C(net5376),
    .D(_08431_),
    .Y(_08469_));
 sg13g2_nor4_1 _16701_ (.A(_08461_),
    .B(_08465_),
    .C(_08468_),
    .D(_08469_),
    .Y(_08470_));
 sg13g2_o21ai_1 _16702_ (.B1(_08470_),
    .Y(_08471_),
    .A1(net5349),
    .A2(_08451_));
 sg13g2_nor3_1 _16703_ (.A(_08395_),
    .B(_00173_),
    .C(_08471_),
    .Y(_08472_));
 sg13g2_nand3_1 _16704_ (.B(_08242_),
    .C(_08246_),
    .A(_08185_),
    .Y(_08473_));
 sg13g2_o21ai_1 _16705_ (.B1(_08473_),
    .Y(_08474_),
    .A1(_08183_),
    .A2(_08263_));
 sg13g2_o21ai_1 _16706_ (.B1(_08252_),
    .Y(_08475_),
    .A1(net5205),
    .A2(_08183_));
 sg13g2_nand2b_1 _16707_ (.Y(_08476_),
    .B(_08445_),
    .A_N(_08385_));
 sg13g2_nand4_1 _16708_ (.B(_08451_),
    .C(_08475_),
    .A(_08206_),
    .Y(_08477_),
    .D(_08476_));
 sg13g2_o21ai_1 _16709_ (.B1(net5378),
    .Y(_08478_),
    .A1(_08474_),
    .A2(_08477_));
 sg13g2_and2_1 _16710_ (.A(net5480),
    .B(_08478_),
    .X(_08479_));
 sg13g2_nand2_1 _16711_ (.Y(_08480_),
    .A(net5370),
    .B(_08319_));
 sg13g2_o21ai_1 _16712_ (.B1(_08480_),
    .Y(_08481_),
    .A1(net5370),
    .A2(_08273_));
 sg13g2_nand2_1 _16713_ (.Y(_08482_),
    .A(net5444),
    .B(_08415_));
 sg13g2_nor2_1 _16714_ (.A(net5436),
    .B(_08452_),
    .Y(_08483_));
 sg13g2_nor3_1 _16715_ (.A(_08276_),
    .B(_08324_),
    .C(_08466_),
    .Y(_08484_));
 sg13g2_o21ai_1 _16716_ (.B1(_08483_),
    .Y(_08485_),
    .A1(net5970),
    .A2(_08334_));
 sg13g2_a21oi_1 _16717_ (.A1(net5437),
    .A2(_08375_),
    .Y(_08486_),
    .B1(_08485_));
 sg13g2_nand3_1 _16718_ (.B(_08484_),
    .C(_08486_),
    .A(_08482_),
    .Y(_08487_));
 sg13g2_nand2_1 _16719_ (.Y(_08488_),
    .A(net5370),
    .B(_08316_));
 sg13g2_o21ai_1 _16720_ (.B1(_08488_),
    .Y(_08489_),
    .A1(net5371),
    .A2(_08265_));
 sg13g2_a21o_1 _16721_ (.A2(_08487_),
    .A1(net5374),
    .B1(_08489_),
    .X(_08490_));
 sg13g2_nor4_1 _16722_ (.A(_08461_),
    .B(_08479_),
    .C(_08481_),
    .D(_08490_),
    .Y(_08491_));
 sg13g2_nor3_1 _16723_ (.A(_08238_),
    .B(_08347_),
    .C(_08472_),
    .Y(_00178_));
 sg13g2_nor2_1 _16724_ (.A(\flash_rom.fsm_state[2] ),
    .B(\flash_rom.fsm_state[0] ),
    .Y(_08492_));
 sg13g2_nor3_1 _16725_ (.A(net5567),
    .B(\flash_rom.fsm_state[1] ),
    .C(net2899),
    .Y(\flash_rom.spi_select ));
 sg13g2_nor3_1 _16726_ (.A(net7369),
    .B(\hvsync_gen.vga.vpos[7] ),
    .C(\hvsync_gen.vga.vpos[6] ),
    .Y(_08493_));
 sg13g2_nor4_1 _16727_ (.A(\hvsync_gen.vga.vpos[9] ),
    .B(\hvsync_gen.vga.vpos[5] ),
    .C(\hvsync_gen.vga.vpos[4] ),
    .D(\hvsync_gen.vga.vpos[1] ),
    .Y(_08494_));
 sg13g2_nand2_1 _16728_ (.Y(_08495_),
    .A(net7370),
    .B(_08494_));
 sg13g2_nor3_2 _16729_ (.A(net7236),
    .B(net7163),
    .C(net7371),
    .Y(_00013_));
 sg13g2_nand2_1 _16730_ (.Y(_08496_),
    .A(_08286_),
    .B(_08380_));
 sg13g2_nand2_2 _16731_ (.Y(_08497_),
    .A(net5477),
    .B(_08331_));
 sg13g2_nand2_1 _16732_ (.Y(_08498_),
    .A(_08251_),
    .B(_08357_));
 sg13g2_nor3_1 _16733_ (.A(net5436),
    .B(net5433),
    .C(_08498_),
    .Y(_08499_));
 sg13g2_or3_1 _16734_ (.A(net5436),
    .B(net5433),
    .C(_08498_),
    .X(_08500_));
 sg13g2_nand3_1 _16735_ (.B(_08323_),
    .C(_08341_),
    .A(_08265_),
    .Y(_08501_));
 sg13g2_nand3_1 _16736_ (.B(_08273_),
    .C(_08311_),
    .A(net5477),
    .Y(_08502_));
 sg13g2_nor2_2 _16737_ (.A(_08501_),
    .B(_08502_),
    .Y(_08503_));
 sg13g2_and4_1 _16738_ (.A(_08172_),
    .B(_08212_),
    .C(_08499_),
    .D(_08503_),
    .X(_08504_));
 sg13g2_nand4_1 _16739_ (.B(_08392_),
    .C(_08424_),
    .A(_08235_),
    .Y(_08505_),
    .D(_08432_));
 sg13g2_a221oi_1 _16740_ (.B2(_08055_),
    .C1(_08505_),
    .B1(_08504_),
    .A1(\atari2600.cpu.dst_reg[1] ),
    .Y(_08506_),
    .A2(net5480));
 sg13g2_nor2_1 _16741_ (.A(_00080_),
    .B(_08505_),
    .Y(_08507_));
 sg13g2_a22oi_1 _16742_ (.Y(_08508_),
    .B1(_08505_),
    .B2(\atari2600.cpu.index_y ),
    .A2(_08211_),
    .A1(\atari2600.cpu.dst_reg[0] ));
 sg13g2_nand4_1 _16743_ (.B(_08499_),
    .C(_08503_),
    .A(_08172_),
    .Y(_08509_),
    .D(_08508_));
 sg13g2_a21oi_2 _16744_ (.B1(_08509_),
    .Y(_08510_),
    .A2(_08507_),
    .A1(_08504_));
 sg13g2_and2_2 _16745_ (.A(_08506_),
    .B(_08510_),
    .X(_08511_));
 sg13g2_nor2_2 _16746_ (.A(_08506_),
    .B(_08510_),
    .Y(_08512_));
 sg13g2_a22oi_1 _16747_ (.Y(_08513_),
    .B1(_08512_),
    .B2(\atari2600.cpu.AXYS[3][3] ),
    .A2(_08511_),
    .A1(\atari2600.cpu.AXYS[0][3] ));
 sg13g2_nor2b_2 _16748_ (.A(_08510_),
    .B_N(_08506_),
    .Y(_08514_));
 sg13g2_nor2b_2 _16749_ (.A(_08506_),
    .B_N(_08510_),
    .Y(_08515_));
 sg13g2_a22oi_1 _16750_ (.Y(_08516_),
    .B1(_08515_),
    .B2(\atari2600.cpu.AXYS[2][3] ),
    .A2(_08514_),
    .A1(\atari2600.cpu.AXYS[1][3] ));
 sg13g2_nand2_2 _16751_ (.Y(_08517_),
    .A(_08513_),
    .B(_08516_));
 sg13g2_nor2_1 _16752_ (.A(_08305_),
    .B(_08335_),
    .Y(_08518_));
 sg13g2_or2_2 _16753_ (.X(_08519_),
    .B(_08329_),
    .A(_08319_));
 sg13g2_or4_1 _16754_ (.A(_08305_),
    .B(_08316_),
    .C(_08335_),
    .D(net5397),
    .X(_08520_));
 sg13g2_nand2_1 _16755_ (.Y(_08521_),
    .A(net5475),
    .B(_08358_));
 sg13g2_or2_1 _16756_ (.X(_08522_),
    .B(_08521_),
    .A(_08520_));
 sg13g2_nor4_2 _16757_ (.A(_08282_),
    .B(_08423_),
    .C(_08437_),
    .Y(_08523_),
    .D(_08501_));
 sg13g2_nor3_2 _16758_ (.A(_08324_),
    .B(_08327_),
    .C(_08407_),
    .Y(_08524_));
 sg13g2_nand2_2 _16759_ (.Y(_08525_),
    .A(_08289_),
    .B(_08292_));
 sg13g2_o21ai_1 _16760_ (.B1(_08524_),
    .Y(_08526_),
    .A1(net5970),
    .A2(_08281_));
 sg13g2_nor2_2 _16761_ (.A(_08525_),
    .B(_08526_),
    .Y(_08527_));
 sg13g2_or2_2 _16762_ (.X(_08528_),
    .B(_08526_),
    .A(_08525_));
 sg13g2_nand3b_1 _16763_ (.B(_08523_),
    .C(_08527_),
    .Y(_08529_),
    .A_N(net5361));
 sg13g2_nand2_2 _16764_ (.Y(_08530_),
    .A(_08230_),
    .B(_08453_));
 sg13g2_nand3b_1 _16765_ (.B(_08295_),
    .C(_08414_),
    .Y(_08531_),
    .A_N(_08280_));
 sg13g2_or3_1 _16766_ (.A(net5479),
    .B(_08530_),
    .C(net5396),
    .X(_08532_));
 sg13g2_nor4_1 _16767_ (.A(net5442),
    .B(net5434),
    .C(net5398),
    .D(_08532_),
    .Y(_08533_));
 sg13g2_nand2b_1 _16768_ (.Y(_08534_),
    .B(_08533_),
    .A_N(net5345));
 sg13g2_inv_2 _16769_ (.Y(_08535_),
    .A(net5307));
 sg13g2_nor2_1 _16770_ (.A(_00101_),
    .B(net5439),
    .Y(_08536_));
 sg13g2_a221oi_1 _16771_ (.B2(\atari2600.cpu.ABL[3] ),
    .C1(_08536_),
    .B1(net5392),
    .A1(\atari2600.cpu.ADD[3] ),
    .Y(_08537_),
    .A2(net5345));
 sg13g2_nand2_1 _16772_ (.Y(_08538_),
    .A(net5308),
    .B(_08537_));
 sg13g2_a221oi_1 _16773_ (.B2(_08517_),
    .C1(_08538_),
    .B1(net5398),
    .A1(\atari2600.cpu.DIMUX[3] ),
    .Y(_08539_),
    .A2(net5434));
 sg13g2_nor2_1 _16774_ (.A(\atari2600.cpu.PC[3] ),
    .B(net5308),
    .Y(_08540_));
 sg13g2_nor2_1 _16775_ (.A(_08539_),
    .B(_08540_),
    .Y(_08541_));
 sg13g2_nor2_1 _16776_ (.A(\atari2600.address_bus_r[3] ),
    .B(net5352),
    .Y(_08542_));
 sg13g2_o21ai_1 _16777_ (.B1(net5352),
    .Y(_08543_),
    .A1(_08539_),
    .A2(_08540_));
 sg13g2_nand2b_1 _16778_ (.Y(_08544_),
    .B(_08543_),
    .A_N(_08542_));
 sg13g2_nor2b_2 _16779_ (.A(_08542_),
    .B_N(_08543_),
    .Y(_08545_));
 sg13g2_mux4_1 _16780_ (.S0(_08510_),
    .A0(_00086_),
    .A1(_00085_),
    .A2(_00084_),
    .A3(_00083_),
    .S1(_08506_),
    .X(_08546_));
 sg13g2_nand2b_1 _16781_ (.Y(_08547_),
    .B(net5398),
    .A_N(_08546_));
 sg13g2_nor2_1 _16782_ (.A(_00097_),
    .B(net5439),
    .Y(_08548_));
 sg13g2_a221oi_1 _16783_ (.B2(\atari2600.cpu.ABL[1] ),
    .C1(_08548_),
    .B1(net5392),
    .A1(\atari2600.cpu.ADD[1] ),
    .Y(_08549_),
    .A2(net5345));
 sg13g2_nand2_1 _16784_ (.Y(_08550_),
    .A(net5307),
    .B(_08549_));
 sg13g2_a21oi_1 _16785_ (.A1(\atari2600.cpu.DIMUX[1] ),
    .A2(net5434),
    .Y(_08551_),
    .B1(_08550_));
 sg13g2_a22oi_1 _16786_ (.Y(_08552_),
    .B1(_08547_),
    .B2(_08551_),
    .A2(_08535_),
    .A1(_08062_));
 sg13g2_mux2_2 _16787_ (.A0(\atari2600.address_bus_r[1] ),
    .A1(_08552_),
    .S(net5353),
    .X(_08553_));
 sg13g2_inv_2 _16788_ (.Y(_08554_),
    .A(net5035));
 sg13g2_mux4_1 _16789_ (.S0(_08510_),
    .A0(_08065_),
    .A1(_08066_),
    .A2(_08063_),
    .A3(_08064_),
    .S1(_08506_),
    .X(_08555_));
 sg13g2_nand2_1 _16790_ (.Y(_08556_),
    .A(net5398),
    .B(_08555_));
 sg13g2_o21ai_1 _16791_ (.B1(\atari2600.cpu.ADD[0] ),
    .Y(_08557_),
    .A1(net5441),
    .A2(net5345));
 sg13g2_nand2_1 _16792_ (.Y(_08558_),
    .A(\atari2600.cpu.ABL[0] ),
    .B(net5392));
 sg13g2_nand3_1 _16793_ (.B(_08557_),
    .C(_08558_),
    .A(net5307),
    .Y(_08559_));
 sg13g2_a21oi_1 _16794_ (.A1(\atari2600.cpu.DIMUX[0] ),
    .A2(net5434),
    .Y(_08560_),
    .B1(_08559_));
 sg13g2_a22oi_1 _16795_ (.Y(_08561_),
    .B1(_08556_),
    .B2(_08560_),
    .A2(_08535_),
    .A1(_08067_));
 sg13g2_mux2_1 _16796_ (.A0(net7336),
    .A1(_08561_),
    .S(net5353),
    .X(_08562_));
 sg13g2_inv_4 _16797_ (.A(_08562_),
    .Y(_08563_));
 sg13g2_nor2_2 _16798_ (.A(net5035),
    .B(_08563_),
    .Y(_08564_));
 sg13g2_nand2_2 _16799_ (.Y(_08565_),
    .A(_08554_),
    .B(net5034));
 sg13g2_a22oi_1 _16800_ (.Y(_08566_),
    .B1(_08514_),
    .B2(\atari2600.cpu.AXYS[1][2] ),
    .A2(_08512_),
    .A1(\atari2600.cpu.AXYS[3][2] ));
 sg13g2_a22oi_1 _16801_ (.Y(_08567_),
    .B1(_08515_),
    .B2(\atari2600.cpu.AXYS[2][2] ),
    .A2(_08511_),
    .A1(\atari2600.cpu.AXYS[0][2] ));
 sg13g2_nand2_2 _16802_ (.Y(_08568_),
    .A(_08566_),
    .B(_08567_));
 sg13g2_nor2_1 _16803_ (.A(_00099_),
    .B(net5439),
    .Y(_08569_));
 sg13g2_a221oi_1 _16804_ (.B2(\atari2600.cpu.ABL[2] ),
    .C1(_08569_),
    .B1(net5392),
    .A1(net5571),
    .Y(_08570_),
    .A2(net5345));
 sg13g2_nand2_1 _16805_ (.Y(_08571_),
    .A(net5307),
    .B(_08570_));
 sg13g2_a221oi_1 _16806_ (.B2(_08568_),
    .C1(_08571_),
    .B1(net5398),
    .A1(\atari2600.cpu.DIMUX[2] ),
    .Y(_08572_),
    .A2(net5434));
 sg13g2_nor2_1 _16807_ (.A(\atari2600.cpu.PC[2] ),
    .B(net5307),
    .Y(_08573_));
 sg13g2_nor2_1 _16808_ (.A(_08572_),
    .B(_08573_),
    .Y(_08574_));
 sg13g2_nor2_1 _16809_ (.A(\atari2600.address_bus_r[2] ),
    .B(net5352),
    .Y(_08575_));
 sg13g2_o21ai_1 _16810_ (.B1(net5352),
    .Y(_08576_),
    .A1(_08572_),
    .A2(_08573_));
 sg13g2_nand2b_1 _16811_ (.Y(_08577_),
    .B(_08576_),
    .A_N(_08575_));
 sg13g2_nor2b_1 _16812_ (.A(_08575_),
    .B_N(_08576_),
    .Y(_08578_));
 sg13g2_nor2_1 _16813_ (.A(_08565_),
    .B(net5033),
    .Y(_08579_));
 sg13g2_nand2_2 _16814_ (.Y(_08580_),
    .A(net4915),
    .B(net5031));
 sg13g2_nor2_2 _16815_ (.A(_08545_),
    .B(net5032),
    .Y(_08581_));
 sg13g2_nand2_1 _16816_ (.Y(_08582_),
    .A(net5037),
    .B(net5030));
 sg13g2_nor2_2 _16817_ (.A(_08565_),
    .B(net5007),
    .Y(_08583_));
 sg13g2_nand2_1 _16818_ (.Y(_08584_),
    .A(net4911),
    .B(_08581_));
 sg13g2_nor4_2 _16819_ (.A(_08313_),
    .B(_08389_),
    .C(net5433),
    .Y(_08585_),
    .D(net5397));
 sg13g2_and2_2 _16820_ (.A(_08232_),
    .B(_08585_),
    .X(_08586_));
 sg13g2_nand2_2 _16821_ (.Y(_08587_),
    .A(_08232_),
    .B(_08585_));
 sg13g2_o21ai_1 _16822_ (.B1(\atari2600.cpu.store ),
    .Y(_08588_),
    .A1(_08287_),
    .A2(_08296_));
 sg13g2_o21ai_1 _16823_ (.B1(_08588_),
    .Y(_08589_),
    .A1(\atari2600.cpu.res ),
    .A2(_08586_));
 sg13g2_inv_1 _16824_ (.Y(_08590_),
    .A(_08589_));
 sg13g2_nand2_1 _16825_ (.Y(_08591_),
    .A(\atari2600.cpu.DIMUX[4] ),
    .B(_08528_));
 sg13g2_nand4_1 _16826_ (.B(_08232_),
    .C(net5440),
    .A(_08230_),
    .Y(_08592_),
    .D(_08453_));
 sg13g2_a22oi_1 _16827_ (.Y(_08593_),
    .B1(_08592_),
    .B2(\atari2600.cpu.ABH[4] ),
    .A2(net5396),
    .A1(\atari2600.cpu.ADD[4] ));
 sg13g2_nand3_1 _16828_ (.B(_08591_),
    .C(_08593_),
    .A(net5308),
    .Y(_08594_));
 sg13g2_o21ai_1 _16829_ (.B1(_08594_),
    .Y(_08595_),
    .A1(\atari2600.cpu.PC[12] ),
    .A2(net5308));
 sg13g2_nand2_2 _16830_ (.Y(_08596_),
    .A(net5352),
    .B(_08595_));
 sg13g2_a22oi_1 _16831_ (.Y(_08597_),
    .B1(_08512_),
    .B2(\atari2600.cpu.AXYS[3][7] ),
    .A2(_08511_),
    .A1(\atari2600.cpu.AXYS[0][7] ));
 sg13g2_a22oi_1 _16832_ (.Y(_08598_),
    .B1(_08515_),
    .B2(\atari2600.cpu.AXYS[2][7] ),
    .A2(_08514_),
    .A1(\atari2600.cpu.AXYS[1][7] ));
 sg13g2_nand2_2 _16833_ (.Y(_08599_),
    .A(_08597_),
    .B(_08598_));
 sg13g2_nor2_1 _16834_ (.A(_00104_),
    .B(net5439),
    .Y(_08600_));
 sg13g2_a221oi_1 _16835_ (.B2(\atari2600.cpu.ABL[7] ),
    .C1(_08600_),
    .B1(net5392),
    .A1(\atari2600.cpu.ADD[7] ),
    .Y(_08601_),
    .A2(net5345));
 sg13g2_nand2_1 _16836_ (.Y(_08602_),
    .A(net5308),
    .B(_08601_));
 sg13g2_a221oi_1 _16837_ (.B2(_08599_),
    .C1(_08602_),
    .B1(_08500_),
    .A1(net5273),
    .Y(_08603_),
    .A2(_08496_));
 sg13g2_a21oi_2 _16838_ (.B1(_08603_),
    .Y(_08604_),
    .A2(_08535_),
    .A1(_08080_));
 sg13g2_nor3_2 _16839_ (.A(_08590_),
    .B(_08596_),
    .C(_08604_),
    .Y(_08605_));
 sg13g2_inv_1 _16840_ (.Y(_08606_),
    .A(_08605_));
 sg13g2_a22oi_1 _16841_ (.Y(_08607_),
    .B1(_08514_),
    .B2(\atari2600.cpu.AXYS[1][5] ),
    .A2(_08512_),
    .A1(\atari2600.cpu.AXYS[3][5] ));
 sg13g2_a22oi_1 _16842_ (.Y(_08608_),
    .B1(_08515_),
    .B2(\atari2600.cpu.AXYS[2][5] ),
    .A2(_08511_),
    .A1(\atari2600.cpu.AXYS[0][5] ));
 sg13g2_nand2_2 _16843_ (.Y(_08609_),
    .A(_08607_),
    .B(_08608_));
 sg13g2_nor2_1 _16844_ (.A(_00100_),
    .B(net5439),
    .Y(_08610_));
 sg13g2_a221oi_1 _16845_ (.B2(\atari2600.cpu.ABL[5] ),
    .C1(_08610_),
    .B1(net5392),
    .A1(net5569),
    .Y(_08611_),
    .A2(net5345));
 sg13g2_nand2_1 _16846_ (.Y(_08612_),
    .A(net5308),
    .B(_08611_));
 sg13g2_a221oi_1 _16847_ (.B2(_08609_),
    .C1(_08612_),
    .B1(net5398),
    .A1(\atari2600.cpu.DIMUX[5] ),
    .Y(_08613_),
    .A2(net5434));
 sg13g2_a21oi_2 _16848_ (.B1(_08613_),
    .Y(_08614_),
    .A2(_08535_),
    .A1(_08073_));
 sg13g2_nor2_2 _16849_ (.A(net5316),
    .B(_08614_),
    .Y(_08615_));
 sg13g2_inv_1 _16850_ (.Y(_08616_),
    .A(_08615_));
 sg13g2_o21ai_1 _16851_ (.B1(_08616_),
    .Y(_08617_),
    .A1(\atari2600.address_bus_r[5] ),
    .A2(net5354));
 sg13g2_a22oi_1 _16852_ (.Y(_08618_),
    .B1(_08515_),
    .B2(\atari2600.cpu.AXYS[2][4] ),
    .A2(_08512_),
    .A1(\atari2600.cpu.AXYS[3][4] ));
 sg13g2_a22oi_1 _16853_ (.Y(_08619_),
    .B1(_08514_),
    .B2(\atari2600.cpu.AXYS[1][4] ),
    .A2(_08511_),
    .A1(\atari2600.cpu.AXYS[0][4] ));
 sg13g2_nand2_2 _16854_ (.Y(_08620_),
    .A(_08618_),
    .B(_08619_));
 sg13g2_o21ai_1 _16855_ (.B1(net5570),
    .Y(_08621_),
    .A1(net5441),
    .A2(_08529_));
 sg13g2_nand2_1 _16856_ (.Y(_08622_),
    .A(\atari2600.cpu.ABL[4] ),
    .B(net5392));
 sg13g2_nand3_1 _16857_ (.B(_08621_),
    .C(_08622_),
    .A(net5309),
    .Y(_08623_));
 sg13g2_a221oi_1 _16858_ (.B2(_08620_),
    .C1(_08623_),
    .B1(net5398),
    .A1(\atari2600.cpu.DIMUX[4] ),
    .Y(_08624_),
    .A2(net5434));
 sg13g2_nor2_1 _16859_ (.A(\atari2600.cpu.PC[4] ),
    .B(net5309),
    .Y(_08625_));
 sg13g2_nor2_1 _16860_ (.A(_08624_),
    .B(_08625_),
    .Y(_08626_));
 sg13g2_nor3_1 _16861_ (.A(net5316),
    .B(_08624_),
    .C(_08625_),
    .Y(_08627_));
 sg13g2_a21o_2 _16862_ (.A2(net5316),
    .A1(\atari2600.address_bus_r[4] ),
    .B1(_08627_),
    .X(_08628_));
 sg13g2_a21oi_1 _16863_ (.A1(net7226),
    .A2(net5316),
    .Y(_08629_),
    .B1(_08627_));
 sg13g2_nand2_1 _16864_ (.Y(_08630_),
    .A(net4876),
    .B(net5026));
 sg13g2_inv_4 _16865_ (.A(net4777),
    .Y(_08631_));
 sg13g2_nand2_2 _16866_ (.Y(_08632_),
    .A(_08605_),
    .B(_08631_));
 sg13g2_nor2_1 _16867_ (.A(_08584_),
    .B(_08632_),
    .Y(_08633_));
 sg13g2_nor2_2 _16868_ (.A(net5316),
    .B(_08604_),
    .Y(_08634_));
 sg13g2_nand3_1 _16869_ (.B(_08595_),
    .C(_08634_),
    .A(_08589_),
    .Y(_08635_));
 sg13g2_nor2_2 _16870_ (.A(net4778),
    .B(_08635_),
    .Y(_08636_));
 sg13g2_or2_2 _16871_ (.X(_08637_),
    .B(_08635_),
    .A(net4778));
 sg13g2_nor2_2 _16872_ (.A(net5984),
    .B(net4724),
    .Y(_08638_));
 sg13g2_nand2_1 _16873_ (.Y(_08639_),
    .A(net2958),
    .B(_08638_));
 sg13g2_a21oi_2 _16874_ (.B1(_08231_),
    .Y(_08640_),
    .A2(_08389_),
    .A1(_08075_));
 sg13g2_inv_1 _16875_ (.Y(_08641_),
    .A(_08640_));
 sg13g2_nand2_1 _16876_ (.Y(_08642_),
    .A(\atari2600.cpu.PC[0] ),
    .B(net5397));
 sg13g2_nand3_1 _16877_ (.B(\atari2600.cpu.php ),
    .C(net5436),
    .A(\atari2600.cpu.C ),
    .Y(_08643_));
 sg13g2_nand2b_1 _16878_ (.Y(_08644_),
    .B(_08313_),
    .A_N(_00095_));
 sg13g2_a22oi_1 _16879_ (.Y(_08645_),
    .B1(_08641_),
    .B2(\atari2600.cpu.ADD[0] ),
    .A2(net5433),
    .A1(\atari2600.cpu.PC[8] ));
 sg13g2_nand4_1 _16880_ (.B(_08643_),
    .C(_08644_),
    .A(_08642_),
    .Y(_08646_),
    .D(_08645_));
 sg13g2_and2_1 _16881_ (.A(_08555_),
    .B(_08586_),
    .X(_08647_));
 sg13g2_nor2_1 _16882_ (.A(_08646_),
    .B(_08647_),
    .Y(_08648_));
 sg13g2_or2_1 _16883_ (.X(_08649_),
    .B(_08647_),
    .A(_08646_));
 sg13g2_nor2_1 _16884_ (.A(_00099_),
    .B(_08640_),
    .Y(_08650_));
 sg13g2_a21oi_2 _16885_ (.B1(_08313_),
    .Y(_08651_),
    .A2(net5436),
    .A1(\atari2600.cpu.php ));
 sg13g2_a221oi_1 _16886_ (.B2(\atari2600.cpu.PC[2] ),
    .C1(_08650_),
    .B1(_08519_),
    .A1(\atari2600.cpu.PC[10] ),
    .Y(_08652_),
    .A2(_08497_));
 sg13g2_o21ai_1 _16887_ (.B1(_08652_),
    .Y(_08653_),
    .A1(_00098_),
    .A2(_08651_));
 sg13g2_nand2_1 _16888_ (.Y(_08654_),
    .A(_08568_),
    .B(_08586_));
 sg13g2_nor2b_1 _16889_ (.A(_08653_),
    .B_N(_08654_),
    .Y(_08655_));
 sg13g2_nand2b_2 _16890_ (.Y(_08656_),
    .B(_08654_),
    .A_N(_08653_));
 sg13g2_nor2_2 _16891_ (.A(net5265),
    .B(net5136),
    .Y(_08657_));
 sg13g2_xnor2_1 _16892_ (.Y(_08658_),
    .A(net5257),
    .B(net5136));
 sg13g2_inv_1 _16893_ (.Y(_08659_),
    .A(_08658_));
 sg13g2_nor2_1 _16894_ (.A(_00097_),
    .B(_08640_),
    .Y(_08660_));
 sg13g2_a221oi_1 _16895_ (.B2(\atari2600.cpu.PC[1] ),
    .C1(_08660_),
    .B1(_08519_),
    .A1(\atari2600.cpu.PC[9] ),
    .Y(_08661_),
    .A2(_08497_));
 sg13g2_o21ai_1 _16896_ (.B1(_08661_),
    .Y(_08662_),
    .A1(_00096_),
    .A2(_08651_));
 sg13g2_nor2_2 _16897_ (.A(_08546_),
    .B(_08587_),
    .Y(_08663_));
 sg13g2_nor2_2 _16898_ (.A(_08662_),
    .B(_08663_),
    .Y(_08664_));
 sg13g2_or2_1 _16899_ (.X(_08665_),
    .B(_08663_),
    .A(_08662_));
 sg13g2_nand2_2 _16900_ (.Y(_08666_),
    .A(net5265),
    .B(net5230));
 sg13g2_nor2_1 _16901_ (.A(net5129),
    .B(_08666_),
    .Y(_08667_));
 sg13g2_a21oi_1 _16902_ (.A1(_08658_),
    .A2(net5238),
    .Y(_08668_),
    .B1(_08667_));
 sg13g2_nor2_2 _16903_ (.A(net5988),
    .B(net5386),
    .Y(_08669_));
 sg13g2_nor3_1 _16904_ (.A(net5988),
    .B(_08135_),
    .C(net5385),
    .Y(_08670_));
 sg13g2_nand2_2 _16905_ (.Y(_08671_),
    .A(_08134_),
    .B(_08669_));
 sg13g2_nand2_1 _16906_ (.Y(_08672_),
    .A(net4724),
    .B(net5343));
 sg13g2_o21ai_1 _16907_ (.B1(_08639_),
    .Y(_00012_),
    .A1(_08668_),
    .A2(_08672_));
 sg13g2_nand2_1 _16908_ (.Y(_08673_),
    .A(net3723),
    .B(_08638_));
 sg13g2_nand2_1 _16909_ (.Y(_08674_),
    .A(_08658_),
    .B(net5230));
 sg13g2_o21ai_1 _16910_ (.B1(_08673_),
    .Y(_00011_),
    .A1(_08672_),
    .A2(_08674_));
 sg13g2_nor2_1 _16911_ (.A(net5035),
    .B(net5034),
    .Y(_08675_));
 sg13g2_nand2_2 _16912_ (.Y(_08676_),
    .A(_08554_),
    .B(_08563_));
 sg13g2_nand2_2 _16913_ (.Y(_08677_),
    .A(net5030),
    .B(net4975));
 sg13g2_nor2_1 _16914_ (.A(net5015),
    .B(_08676_),
    .Y(_08678_));
 sg13g2_nand2_2 _16915_ (.Y(_08679_),
    .A(_08581_),
    .B(net4992));
 sg13g2_nor2_2 _16916_ (.A(net4751),
    .B(_08679_),
    .Y(_08680_));
 sg13g2_nor2_2 _16917_ (.A(_08637_),
    .B(_08679_),
    .Y(_08681_));
 sg13g2_nor2_2 _16918_ (.A(net5984),
    .B(_08681_),
    .Y(_08682_));
 sg13g2_nand2_1 _16919_ (.Y(_08683_),
    .A(net2981),
    .B(_08682_));
 sg13g2_nand2_1 _16920_ (.Y(_08684_),
    .A(net5343),
    .B(_08681_));
 sg13g2_o21ai_1 _16921_ (.B1(_08683_),
    .Y(_00010_),
    .A1(_08668_),
    .A2(_08684_));
 sg13g2_nand2_1 _16922_ (.Y(_08685_),
    .A(net3130),
    .B(_08682_));
 sg13g2_o21ai_1 _16923_ (.B1(_08685_),
    .Y(_00009_),
    .A1(_08674_),
    .A2(_08684_));
 sg13g2_nor2_1 _16924_ (.A(net2892),
    .B(net5537),
    .Y(_00000_));
 sg13g2_nor2_2 _16925_ (.A(net5840),
    .B(_08120_),
    .Y(_08686_));
 sg13g2_nand2_1 _16926_ (.Y(_08687_),
    .A(net5552),
    .B(net5839));
 sg13g2_and2_1 _16927_ (.A(\hvsync_gen.hpos[4] ),
    .B(net5849),
    .X(_08688_));
 sg13g2_nand2_1 _16928_ (.Y(_08689_),
    .A(net5850),
    .B(net5849));
 sg13g2_nand3_1 _16929_ (.B(net5845),
    .C(net5531),
    .A(net5843),
    .Y(_08690_));
 sg13g2_a21oi_1 _16930_ (.A1(_08686_),
    .A2(_08690_),
    .Y(_08691_),
    .B1(net7366));
 sg13g2_nor2_1 _16931_ (.A(net5850),
    .B(net5849),
    .Y(_08692_));
 sg13g2_or2_1 _16932_ (.X(_08693_),
    .B(net5849),
    .A(net5850));
 sg13g2_nor2_2 _16933_ (.A(net5845),
    .B(net5516),
    .Y(_08694_));
 sg13g2_nor3_1 _16934_ (.A(net5846),
    .B(net5840),
    .C(net5516),
    .Y(_08695_));
 sg13g2_nor2_2 _16935_ (.A(net5843),
    .B(net5840),
    .Y(_08696_));
 sg13g2_nor2_1 _16936_ (.A(_08120_),
    .B(_08696_),
    .Y(_08697_));
 sg13g2_o21ai_1 _16937_ (.B1(net5839),
    .Y(_08698_),
    .A1(net5843),
    .A2(net5840));
 sg13g2_nor3_2 _16938_ (.A(_08691_),
    .B(_08695_),
    .C(net5512),
    .Y(_00047_));
 sg13g2_nand4_1 _16939_ (.B(net7039),
    .C(\hvsync_gen.vga.vpos[6] ),
    .A(\hvsync_gen.vga.vpos[8] ),
    .Y(_08699_),
    .D(\hvsync_gen.vga.vpos[5] ));
 sg13g2_nor2_1 _16940_ (.A(\atari2600.tia.vblank ),
    .B(\hvsync_gen.vga.vpos[9] ),
    .Y(_08700_));
 sg13g2_nand3_1 _16941_ (.B(_08699_),
    .C(_08700_),
    .A(_08698_),
    .Y(_08701_));
 sg13g2_xor2_1 _16942_ (.B(\hvsync_gen.vga.vpos[0] ),
    .A(\frame_counter[0] ),
    .X(_08702_));
 sg13g2_xnor2_1 _16943_ (.Y(_08703_),
    .A(\frame_counter[0] ),
    .B(\hvsync_gen.vga.vpos[0] ));
 sg13g2_nand2_1 _16944_ (.Y(_08704_),
    .A(\b_pwm_odd[8] ),
    .B(_08703_));
 sg13g2_nand2_1 _16945_ (.Y(_08705_),
    .A(\b_pwm_even[8] ),
    .B(_08702_));
 sg13g2_a21oi_2 _16946_ (.B1(_08701_),
    .Y(uo_out[6]),
    .A2(_08705_),
    .A1(_08704_));
 sg13g2_nand2_1 _16947_ (.Y(_08706_),
    .A(\b_pwm_odd[9] ),
    .B(_08703_));
 sg13g2_nand2_1 _16948_ (.Y(_08707_),
    .A(\b_pwm_even[9] ),
    .B(_08702_));
 sg13g2_a21oi_2 _16949_ (.B1(_08701_),
    .Y(uo_out[2]),
    .A2(_08707_),
    .A1(_08706_));
 sg13g2_nand2_1 _16950_ (.Y(_08708_),
    .A(\g_pwm_odd[8] ),
    .B(_08703_));
 sg13g2_nand2_1 _16951_ (.Y(_08709_),
    .A(\g_pwm_even[8] ),
    .B(_08702_));
 sg13g2_a21oi_2 _16952_ (.B1(_08701_),
    .Y(uo_out[5]),
    .A2(_08709_),
    .A1(_08708_));
 sg13g2_nand2_1 _16953_ (.Y(_08710_),
    .A(\g_pwm_odd[9] ),
    .B(_08703_));
 sg13g2_nand2_1 _16954_ (.Y(_08711_),
    .A(\g_pwm_even[9] ),
    .B(_08702_));
 sg13g2_a21oi_2 _16955_ (.B1(_08701_),
    .Y(uo_out[1]),
    .A2(_08711_),
    .A1(_08710_));
 sg13g2_nand2_1 _16956_ (.Y(_08712_),
    .A(\r_pwm_odd[8] ),
    .B(_08703_));
 sg13g2_nand2_1 _16957_ (.Y(_08713_),
    .A(\r_pwm_even[8] ),
    .B(_08702_));
 sg13g2_a21oi_2 _16958_ (.B1(_08701_),
    .Y(uo_out[4]),
    .A2(_08713_),
    .A1(_08712_));
 sg13g2_nand2_1 _16959_ (.Y(_08714_),
    .A(\r_pwm_odd[9] ),
    .B(_08703_));
 sg13g2_nand2_1 _16960_ (.Y(_08715_),
    .A(\r_pwm_even[9] ),
    .B(_08702_));
 sg13g2_a21oi_2 _16961_ (.B1(_08701_),
    .Y(uo_out[0]),
    .A2(_08715_),
    .A1(_08714_));
 sg13g2_a22oi_1 _16962_ (.Y(_08716_),
    .B1(_08512_),
    .B2(\atari2600.cpu.AXYS[3][6] ),
    .A2(_08511_),
    .A1(\atari2600.cpu.AXYS[0][6] ));
 sg13g2_a22oi_1 _16963_ (.Y(_08717_),
    .B1(_08515_),
    .B2(\atari2600.cpu.AXYS[2][6] ),
    .A2(_08514_),
    .A1(\atari2600.cpu.AXYS[1][6] ));
 sg13g2_nand2_2 _16964_ (.Y(_08718_),
    .A(_08716_),
    .B(_08717_));
 sg13g2_nor2_1 _16965_ (.A(_00103_),
    .B(net5439),
    .Y(_08719_));
 sg13g2_a221oi_1 _16966_ (.B2(\atari2600.cpu.ABL[6] ),
    .C1(_08719_),
    .B1(net5392),
    .A1(\atari2600.cpu.ADD[6] ),
    .Y(_08720_),
    .A2(net5345));
 sg13g2_nand2_1 _16967_ (.Y(_08721_),
    .A(net5308),
    .B(_08720_));
 sg13g2_a221oi_1 _16968_ (.B2(_08718_),
    .C1(_08721_),
    .B1(net5398),
    .A1(\atari2600.cpu.DIMUX[6] ),
    .Y(_08722_),
    .A2(net5434));
 sg13g2_nor2_1 _16969_ (.A(\atari2600.cpu.PC[6] ),
    .B(net5308),
    .Y(_08723_));
 sg13g2_nor2_1 _16970_ (.A(_08722_),
    .B(_08723_),
    .Y(_08724_));
 sg13g2_nor2_1 _16971_ (.A(\atari2600.address_bus_r[6] ),
    .B(net5352),
    .Y(_08725_));
 sg13g2_o21ai_1 _16972_ (.B1(net5352),
    .Y(_08726_),
    .A1(_08722_),
    .A2(_08723_));
 sg13g2_nand2b_1 _16973_ (.Y(_08727_),
    .B(_08726_),
    .A_N(_08725_));
 sg13g2_nor2b_1 _16974_ (.A(_08725_),
    .B_N(_08726_),
    .Y(_08728_));
 sg13g2_nand2b_1 _16975_ (.Y(_08729_),
    .B(net5028),
    .A_N(net4878));
 sg13g2_nand2_2 _16976_ (.Y(_08730_),
    .A(_08545_),
    .B(net5031));
 sg13g2_nor2_1 _16977_ (.A(_08554_),
    .B(_08563_),
    .Y(_08731_));
 sg13g2_nand2_2 _16978_ (.Y(_08732_),
    .A(net5035),
    .B(net5034));
 sg13g2_a22oi_1 _16979_ (.Y(_08733_),
    .B1(net4839),
    .B2(\atari2600.ram[63][0] ),
    .A2(net4969),
    .A1(\atari2600.ram[60][0] ));
 sg13g2_nor2_2 _16980_ (.A(_08554_),
    .B(net5034),
    .Y(_08734_));
 sg13g2_nand2_2 _16981_ (.Y(_08735_),
    .A(_08553_),
    .B(_08563_));
 sg13g2_a22oi_1 _16982_ (.Y(_08736_),
    .B1(net4793),
    .B2(\atari2600.ram[62][0] ),
    .A2(net4887),
    .A1(\atari2600.ram[61][0] ));
 sg13g2_a21oi_1 _16983_ (.A1(_08733_),
    .A2(_08736_),
    .Y(_08737_),
    .B1(net4953));
 sg13g2_a22oi_1 _16984_ (.Y(_08738_),
    .B1(net4855),
    .B2(\atari2600.ram[55][0] ),
    .A2(net4985),
    .A1(\atari2600.ram[52][0] ));
 sg13g2_a22oi_1 _16985_ (.Y(_08739_),
    .B1(net4810),
    .B2(\atari2600.ram[54][0] ),
    .A2(net4904),
    .A1(\atari2600.ram[53][0] ));
 sg13g2_a21oi_1 _16986_ (.A1(_08738_),
    .A2(_08739_),
    .Y(_08740_),
    .B1(net5012));
 sg13g2_nor2_2 _16987_ (.A(net5039),
    .B(net5031),
    .Y(_08741_));
 sg13g2_nand2_1 _16988_ (.Y(_08742_),
    .A(_08545_),
    .B(net5033));
 sg13g2_a22oi_1 _16989_ (.Y(_08743_),
    .B1(net4838),
    .B2(\atari2600.ram[59][0] ),
    .A2(net4968),
    .A1(\atari2600.ram[56][0] ));
 sg13g2_a22oi_1 _16990_ (.Y(_08744_),
    .B1(net4792),
    .B2(\atari2600.ram[58][0] ),
    .A2(net4886),
    .A1(\atari2600.ram[57][0] ));
 sg13g2_a21oi_2 _16991_ (.B1(net4940),
    .Y(_08745_),
    .A2(_08744_),
    .A1(_08743_));
 sg13g2_nor2_2 _16992_ (.A(net5036),
    .B(net5031),
    .Y(_08746_));
 sg13g2_nand2_1 _16993_ (.Y(_08747_),
    .A(net5039),
    .B(net5033));
 sg13g2_a22oi_1 _16994_ (.Y(_08748_),
    .B1(net4842),
    .B2(\atari2600.ram[51][0] ),
    .A2(net4972),
    .A1(\atari2600.ram[48][0] ));
 sg13g2_a22oi_1 _16995_ (.Y(_08749_),
    .B1(net4794),
    .B2(\atari2600.ram[50][0] ),
    .A2(net4888),
    .A1(\atari2600.ram[49][0] ));
 sg13g2_a21oi_1 _16996_ (.A1(_08748_),
    .A2(_08749_),
    .Y(_08750_),
    .B1(net4926));
 sg13g2_nor4_2 _16997_ (.A(_08737_),
    .B(_08740_),
    .C(_08745_),
    .Y(_08751_),
    .D(_08750_));
 sg13g2_nor2_1 _16998_ (.A(net4776),
    .B(_08751_),
    .Y(_08752_));
 sg13g2_and2_2 _16999_ (.A(net4879),
    .B(net5028),
    .X(_08753_));
 sg13g2_nand2_1 _17000_ (.Y(_08754_),
    .A(net4878),
    .B(net5028));
 sg13g2_a22oi_1 _17001_ (.Y(_08755_),
    .B1(net4851),
    .B2(\atari2600.ram[31][0] ),
    .A2(net4978),
    .A1(\atari2600.ram[28][0] ));
 sg13g2_a22oi_1 _17002_ (.Y(_08756_),
    .B1(net4806),
    .B2(\atari2600.ram[30][0] ),
    .A2(net4900),
    .A1(\atari2600.ram[29][0] ));
 sg13g2_a21oi_1 _17003_ (.A1(_08755_),
    .A2(_08756_),
    .Y(_08757_),
    .B1(net4952));
 sg13g2_a22oi_1 _17004_ (.Y(_08758_),
    .B1(net4841),
    .B2(\atari2600.ram[27][0] ),
    .A2(net4970),
    .A1(\atari2600.ram[24][0] ));
 sg13g2_a22oi_1 _17005_ (.Y(_08759_),
    .B1(net4794),
    .B2(\atari2600.ram[26][0] ),
    .A2(net4888),
    .A1(\atari2600.ram[25][0] ));
 sg13g2_a21oi_2 _17006_ (.B1(net4940),
    .Y(_08760_),
    .A2(_08759_),
    .A1(_08758_));
 sg13g2_a22oi_1 _17007_ (.Y(_08761_),
    .B1(net4848),
    .B2(\atari2600.ram[19][0] ),
    .A2(net4979),
    .A1(\atari2600.ram[16][0] ));
 sg13g2_a22oi_1 _17008_ (.Y(_08762_),
    .B1(net4802),
    .B2(\atari2600.ram[18][0] ),
    .A2(net4899),
    .A1(\atari2600.ram[17][0] ));
 sg13g2_a21oi_2 _17009_ (.B1(net4929),
    .Y(_08763_),
    .A2(_08762_),
    .A1(_08761_));
 sg13g2_a22oi_1 _17010_ (.Y(_08764_),
    .B1(net4847),
    .B2(\atari2600.ram[23][0] ),
    .A2(net4978),
    .A1(\atari2600.ram[20][0] ));
 sg13g2_a22oi_1 _17011_ (.Y(_08765_),
    .B1(net4802),
    .B2(\atari2600.ram[22][0] ),
    .A2(net4897),
    .A1(\atari2600.ram[21][0] ));
 sg13g2_a21oi_1 _17012_ (.A1(_08764_),
    .A2(_08765_),
    .Y(_08766_),
    .B1(net5008));
 sg13g2_nor4_2 _17013_ (.A(_08757_),
    .B(_08760_),
    .C(_08763_),
    .Y(_08767_),
    .D(_08766_));
 sg13g2_a22oi_1 _17014_ (.Y(_08768_),
    .B1(net4844),
    .B2(\atari2600.ram[3][0] ),
    .A2(net4974),
    .A1(\atari2600.ram[0][0] ));
 sg13g2_a22oi_1 _17015_ (.Y(_08769_),
    .B1(net4798),
    .B2(\atari2600.ram[2][0] ),
    .A2(net4892),
    .A1(\atari2600.ram[1][0] ));
 sg13g2_a21oi_2 _17016_ (.B1(net4927),
    .Y(_08770_),
    .A2(_08769_),
    .A1(_08768_));
 sg13g2_a22oi_1 _17017_ (.Y(_08771_),
    .B1(net4835),
    .B2(\atari2600.ram[15][0] ),
    .A2(net4965),
    .A1(\atari2600.ram[12][0] ));
 sg13g2_a22oi_1 _17018_ (.Y(_08772_),
    .B1(net4789),
    .B2(\atari2600.ram[14][0] ),
    .A2(net4883),
    .A1(\atari2600.ram[13][0] ));
 sg13g2_a21oi_2 _17019_ (.B1(net4950),
    .Y(_08773_),
    .A2(_08772_),
    .A1(_08771_));
 sg13g2_a22oi_1 _17020_ (.Y(_08774_),
    .B1(net4843),
    .B2(\atari2600.ram[7][0] ),
    .A2(net4973),
    .A1(\atari2600.ram[4][0] ));
 sg13g2_a22oi_1 _17021_ (.Y(_08775_),
    .B1(net4799),
    .B2(\atari2600.ram[6][0] ),
    .A2(net4893),
    .A1(\atari2600.ram[5][0] ));
 sg13g2_a21oi_1 _17022_ (.A1(_08774_),
    .A2(_08775_),
    .Y(_08776_),
    .B1(net5007));
 sg13g2_a22oi_1 _17023_ (.Y(_08777_),
    .B1(net4834),
    .B2(\atari2600.ram[11][0] ),
    .A2(net4964),
    .A1(\atari2600.ram[8][0] ));
 sg13g2_a22oi_1 _17024_ (.Y(_08778_),
    .B1(net4790),
    .B2(\atari2600.ram[10][0] ),
    .A2(net4892),
    .A1(\atari2600.ram[9][0] ));
 sg13g2_a21oi_1 _17025_ (.A1(_08777_),
    .A2(_08778_),
    .Y(_08779_),
    .B1(net4938));
 sg13g2_nor4_2 _17026_ (.A(_08770_),
    .B(_08773_),
    .C(_08776_),
    .Y(_08780_),
    .D(_08779_));
 sg13g2_nor2_1 _17027_ (.A(net4777),
    .B(_08780_),
    .Y(_08781_));
 sg13g2_nor2_2 _17028_ (.A(net4878),
    .B(net5028),
    .Y(_08782_));
 sg13g2_nand2b_1 _17029_ (.Y(_08783_),
    .B(net5025),
    .A_N(net4878));
 sg13g2_a22oi_1 _17030_ (.Y(_08784_),
    .B1(net4834),
    .B2(\atari2600.ram[43][0] ),
    .A2(net4964),
    .A1(\atari2600.ram[40][0] ));
 sg13g2_a22oi_1 _17031_ (.Y(_08785_),
    .B1(net4788),
    .B2(\atari2600.ram[42][0] ),
    .A2(net4884),
    .A1(\atari2600.ram[41][0] ));
 sg13g2_a21oi_1 _17032_ (.A1(_08784_),
    .A2(_08785_),
    .Y(_08786_),
    .B1(net4937));
 sg13g2_a22oi_1 _17033_ (.Y(_08787_),
    .B1(net4830),
    .B2(\atari2600.ram[39][0] ),
    .A2(net4960),
    .A1(\atari2600.ram[36][0] ));
 sg13g2_a22oi_1 _17034_ (.Y(_08788_),
    .B1(net4786),
    .B2(\atari2600.ram[38][0] ),
    .A2(net4882),
    .A1(\atari2600.ram[37][0] ));
 sg13g2_a21oi_2 _17035_ (.B1(net5006),
    .Y(_08789_),
    .A2(_08788_),
    .A1(_08787_));
 sg13g2_a22oi_1 _17036_ (.Y(_08790_),
    .B1(net4835),
    .B2(\atari2600.ram[47][0] ),
    .A2(net4965),
    .A1(\atari2600.ram[44][0] ));
 sg13g2_a22oi_1 _17037_ (.Y(_08791_),
    .B1(net4789),
    .B2(\atari2600.ram[46][0] ),
    .A2(net4883),
    .A1(\atari2600.ram[45][0] ));
 sg13g2_a21oi_1 _17038_ (.A1(_08790_),
    .A2(_08791_),
    .Y(_08792_),
    .B1(net4949));
 sg13g2_a22oi_1 _17039_ (.Y(_08793_),
    .B1(net4832),
    .B2(\atari2600.ram[35][0] ),
    .A2(net4962),
    .A1(\atari2600.ram[32][0] ));
 sg13g2_a22oi_1 _17040_ (.Y(_08794_),
    .B1(net4787),
    .B2(\atari2600.ram[34][0] ),
    .A2(net4881),
    .A1(\atari2600.ram[33][0] ));
 sg13g2_a21oi_2 _17041_ (.B1(net4925),
    .Y(_08795_),
    .A2(_08794_),
    .A1(_08793_));
 sg13g2_nor4_2 _17042_ (.A(_08786_),
    .B(_08789_),
    .C(_08792_),
    .Y(_08796_),
    .D(_08795_));
 sg13g2_nor2_1 _17043_ (.A(net4772),
    .B(_08796_),
    .Y(_08797_));
 sg13g2_o21ai_1 _17044_ (.B1(net5024),
    .Y(_08798_),
    .A1(net4773),
    .A2(_08767_));
 sg13g2_nor4_1 _17045_ (.A(_08752_),
    .B(_08781_),
    .C(_08797_),
    .D(_08798_),
    .Y(_08799_));
 sg13g2_a22oi_1 _17046_ (.Y(_08800_),
    .B1(net4859),
    .B2(\atari2600.ram[99][0] ),
    .A2(net4984),
    .A1(\atari2600.ram[96][0] ));
 sg13g2_a22oi_1 _17047_ (.Y(_08801_),
    .B1(net4813),
    .B2(\atari2600.ram[98][0] ),
    .A2(net4903),
    .A1(\atari2600.ram[97][0] ));
 sg13g2_a21oi_2 _17048_ (.B1(net4931),
    .Y(_08802_),
    .A2(_08801_),
    .A1(_08800_));
 sg13g2_a22oi_1 _17049_ (.Y(_08803_),
    .B1(net4861),
    .B2(\atari2600.ram[111][0] ),
    .A2(net4988),
    .A1(\atari2600.ram[108][0] ));
 sg13g2_a22oi_1 _17050_ (.Y(_08804_),
    .B1(net4812),
    .B2(\atari2600.ram[110][0] ),
    .A2(net4906),
    .A1(\atari2600.ram[109][0] ));
 sg13g2_a21oi_1 _17051_ (.A1(_08803_),
    .A2(_08804_),
    .Y(_08805_),
    .B1(net4956));
 sg13g2_a22oi_1 _17052_ (.Y(_08806_),
    .B1(net4855),
    .B2(\atari2600.ram[103][0] ),
    .A2(net4985),
    .A1(\atari2600.ram[100][0] ));
 sg13g2_a22oi_1 _17053_ (.Y(_08807_),
    .B1(net4809),
    .B2(\atari2600.ram[102][0] ),
    .A2(net4903),
    .A1(\atari2600.ram[101][0] ));
 sg13g2_a21oi_1 _17054_ (.A1(_08806_),
    .A2(_08807_),
    .Y(_08808_),
    .B1(net5012));
 sg13g2_a22oi_1 _17055_ (.Y(_08809_),
    .B1(net4859),
    .B2(\atari2600.ram[107][0] ),
    .A2(net4989),
    .A1(\atari2600.ram[104][0] ));
 sg13g2_a22oi_1 _17056_ (.Y(_08810_),
    .B1(net4813),
    .B2(\atari2600.ram[106][0] ),
    .A2(net4908),
    .A1(\atari2600.ram[105][0] ));
 sg13g2_a21oi_1 _17057_ (.A1(_08809_),
    .A2(_08810_),
    .Y(_08811_),
    .B1(net4943));
 sg13g2_nor4_2 _17058_ (.A(_08802_),
    .B(_08805_),
    .C(_08808_),
    .Y(_08812_),
    .D(_08811_));
 sg13g2_o21ai_1 _17059_ (.B1(net5020),
    .Y(_08813_),
    .A1(net4772),
    .A2(_08812_));
 sg13g2_a22oi_1 _17060_ (.Y(_08814_),
    .B1(net4857),
    .B2(\atari2600.ram[119][0] ),
    .A2(net4987),
    .A1(\atari2600.ram[116][0] ));
 sg13g2_a22oi_1 _17061_ (.Y(_08815_),
    .B1(net4796),
    .B2(\atari2600.ram[118][0] ),
    .A2(net4890),
    .A1(\atari2600.ram[117][0] ));
 sg13g2_a21oi_1 _17062_ (.A1(_08814_),
    .A2(_08815_),
    .Y(_08816_),
    .B1(net5013));
 sg13g2_a22oi_1 _17063_ (.Y(_08817_),
    .B1(net4863),
    .B2(\atari2600.ram[127][0] ),
    .A2(net4977),
    .A1(\atari2600.ram[124][0] ));
 sg13g2_a22oi_1 _17064_ (.Y(_08818_),
    .B1(net4818),
    .B2(\atari2600.ram[126][0] ),
    .A2(net4913),
    .A1(\atari2600.ram[125][0] ));
 sg13g2_a21oi_1 _17065_ (.A1(_08817_),
    .A2(_08818_),
    .Y(_08819_),
    .B1(net4956));
 sg13g2_a22oi_1 _17066_ (.Y(_08820_),
    .B1(net4853),
    .B2(\atari2600.ram[115][0] ),
    .A2(net4983),
    .A1(\atari2600.ram[112][0] ));
 sg13g2_a22oi_1 _17067_ (.Y(_08821_),
    .B1(net4808),
    .B2(\atari2600.ram[114][0] ),
    .A2(net4902),
    .A1(\atari2600.ram[113][0] ));
 sg13g2_a21oi_2 _17068_ (.B1(net4930),
    .Y(_08822_),
    .A2(_08821_),
    .A1(_08820_));
 sg13g2_a22oi_1 _17069_ (.Y(_08823_),
    .B1(net4858),
    .B2(\atari2600.ram[123][0] ),
    .A2(net4986),
    .A1(\atari2600.ram[120][0] ));
 sg13g2_a22oi_1 _17070_ (.Y(_08824_),
    .B1(net4817),
    .B2(\atari2600.ram[122][0] ),
    .A2(net4906),
    .A1(\atari2600.ram[121][0] ));
 sg13g2_a21oi_1 _17071_ (.A1(_08823_),
    .A2(_08824_),
    .Y(_08825_),
    .B1(net4944));
 sg13g2_nor4_1 _17072_ (.A(_08816_),
    .B(_08819_),
    .C(_08822_),
    .D(_08825_),
    .Y(_08826_));
 sg13g2_nor2_1 _17073_ (.A(_08729_),
    .B(_08826_),
    .Y(_08827_));
 sg13g2_a22oi_1 _17074_ (.Y(_08828_),
    .B1(net4870),
    .B2(\atari2600.ram[71][0] ),
    .A2(net5000),
    .A1(\atari2600.ram[68][0] ));
 sg13g2_a22oi_1 _17075_ (.Y(_08829_),
    .B1(net4826),
    .B2(\atari2600.ram[70][0] ),
    .A2(net4920),
    .A1(\atari2600.ram[69][0] ));
 sg13g2_a21oi_1 _17076_ (.A1(_08828_),
    .A2(_08829_),
    .Y(_08830_),
    .B1(net5015));
 sg13g2_a22oi_1 _17077_ (.Y(_08831_),
    .B1(net4869),
    .B2(\atari2600.ram[67][0] ),
    .A2(net5000),
    .A1(\atari2600.ram[64][0] ));
 sg13g2_a22oi_1 _17078_ (.Y(_08832_),
    .B1(net4825),
    .B2(\atari2600.ram[66][0] ),
    .A2(net4921),
    .A1(\atari2600.ram[65][0] ));
 sg13g2_a21oi_1 _17079_ (.A1(_08831_),
    .A2(_08832_),
    .Y(_08833_),
    .B1(net4934));
 sg13g2_a22oi_1 _17080_ (.Y(_08834_),
    .B1(net4872),
    .B2(\atari2600.ram[79][0] ),
    .A2(net5003),
    .A1(\atari2600.ram[76][0] ));
 sg13g2_a22oi_1 _17081_ (.Y(_08835_),
    .B1(net4827),
    .B2(\atari2600.ram[78][0] ),
    .A2(net4922),
    .A1(\atari2600.ram[77][0] ));
 sg13g2_a21oi_2 _17082_ (.B1(net4959),
    .Y(_08836_),
    .A2(_08835_),
    .A1(_08834_));
 sg13g2_a22oi_1 _17083_ (.Y(_08837_),
    .B1(net4871),
    .B2(\atari2600.ram[75][0] ),
    .A2(net5002),
    .A1(\atari2600.ram[72][0] ));
 sg13g2_a22oi_1 _17084_ (.Y(_08838_),
    .B1(net4827),
    .B2(\atari2600.ram[74][0] ),
    .A2(net4922),
    .A1(\atari2600.ram[73][0] ));
 sg13g2_a21oi_1 _17085_ (.A1(_08837_),
    .A2(_08838_),
    .Y(_08839_),
    .B1(net4946));
 sg13g2_nor4_2 _17086_ (.A(_08830_),
    .B(_08833_),
    .C(_08836_),
    .Y(_08840_),
    .D(_08839_));
 sg13g2_nor2_1 _17087_ (.A(net4779),
    .B(_08840_),
    .Y(_08841_));
 sg13g2_a22oi_1 _17088_ (.Y(_08842_),
    .B1(net4847),
    .B2(\atari2600.ram[87][0] ),
    .A2(net4977),
    .A1(\atari2600.ram[84][0] ));
 sg13g2_a22oi_1 _17089_ (.Y(_08843_),
    .B1(net4803),
    .B2(\atari2600.ram[86][0] ),
    .A2(net4898),
    .A1(\atari2600.ram[85][0] ));
 sg13g2_a21oi_1 _17090_ (.A1(_08842_),
    .A2(_08843_),
    .Y(_08844_),
    .B1(net5009));
 sg13g2_a22oi_1 _17091_ (.Y(_08845_),
    .B1(net4867),
    .B2(\atari2600.ram[95][0] ),
    .A2(net4997),
    .A1(\atari2600.ram[92][0] ));
 sg13g2_a22oi_1 _17092_ (.Y(_08846_),
    .B1(net4822),
    .B2(\atari2600.ram[94][0] ),
    .A2(net4917),
    .A1(\atari2600.ram[93][0] ));
 sg13g2_a21oi_2 _17093_ (.B1(net4957),
    .Y(_08847_),
    .A2(_08846_),
    .A1(_08845_));
 sg13g2_a22oi_1 _17094_ (.Y(_08848_),
    .B1(net4864),
    .B2(\atari2600.ram[83][0] ),
    .A2(net4995),
    .A1(\atari2600.ram[80][0] ));
 sg13g2_a22oi_1 _17095_ (.Y(_08849_),
    .B1(net4820),
    .B2(\atari2600.ram[82][0] ),
    .A2(net4915),
    .A1(\atari2600.ram[81][0] ));
 sg13g2_a21oi_1 _17096_ (.A1(_08848_),
    .A2(_08849_),
    .Y(_08850_),
    .B1(net4934));
 sg13g2_a22oi_1 _17097_ (.Y(_08851_),
    .B1(net4850),
    .B2(\atari2600.ram[91][0] ),
    .A2(net4980),
    .A1(\atari2600.ram[88][0] ));
 sg13g2_a22oi_1 _17098_ (.Y(_08852_),
    .B1(net4821),
    .B2(\atari2600.ram[90][0] ),
    .A2(net4916),
    .A1(\atari2600.ram[89][0] ));
 sg13g2_a21oi_2 _17099_ (.B1(net4942),
    .Y(_08853_),
    .A2(_08852_),
    .A1(_08851_));
 sg13g2_nor4_2 _17100_ (.A(_08844_),
    .B(_08847_),
    .C(_08850_),
    .Y(_08854_),
    .D(_08853_));
 sg13g2_nor2_1 _17101_ (.A(net4775),
    .B(_08854_),
    .Y(_08855_));
 sg13g2_nor4_2 _17102_ (.A(_08813_),
    .B(_08827_),
    .C(_08841_),
    .Y(_08856_),
    .D(_08855_));
 sg13g2_nor2_2 _17103_ (.A(_08799_),
    .B(_08856_),
    .Y(_00001_));
 sg13g2_a22oi_1 _17104_ (.Y(_08857_),
    .B1(net4983),
    .B2(\atari2600.ram[52][1] ),
    .A2(net4902),
    .A1(\atari2600.ram[53][1] ));
 sg13g2_a22oi_1 _17105_ (.Y(_08858_),
    .B1(net4792),
    .B2(\atari2600.ram[54][1] ),
    .A2(net4853),
    .A1(\atari2600.ram[55][1] ));
 sg13g2_a21oi_2 _17106_ (.B1(net5012),
    .Y(_08859_),
    .A2(_08858_),
    .A1(_08857_));
 sg13g2_a22oi_1 _17107_ (.Y(_08860_),
    .B1(net4840),
    .B2(\atari2600.ram[51][1] ),
    .A2(net4970),
    .A1(\atari2600.ram[48][1] ));
 sg13g2_a22oi_1 _17108_ (.Y(_08861_),
    .B1(net4795),
    .B2(\atari2600.ram[50][1] ),
    .A2(net4889),
    .A1(\atari2600.ram[49][1] ));
 sg13g2_a21oi_2 _17109_ (.B1(net4936),
    .Y(_08862_),
    .A2(_08861_),
    .A1(_08860_));
 sg13g2_a22oi_1 _17110_ (.Y(_08863_),
    .B1(net4839),
    .B2(\atari2600.ram[63][1] ),
    .A2(net4969),
    .A1(\atari2600.ram[60][1] ));
 sg13g2_a22oi_1 _17111_ (.Y(_08864_),
    .B1(net4791),
    .B2(\atari2600.ram[62][1] ),
    .A2(net4887),
    .A1(\atari2600.ram[61][1] ));
 sg13g2_a21oi_1 _17112_ (.A1(_08863_),
    .A2(_08864_),
    .Y(_08865_),
    .B1(net4951));
 sg13g2_a22oi_1 _17113_ (.Y(_08866_),
    .B1(net4837),
    .B2(\atari2600.ram[59][1] ),
    .A2(net4967),
    .A1(\atari2600.ram[56][1] ));
 sg13g2_a22oi_1 _17114_ (.Y(_08867_),
    .B1(net4791),
    .B2(\atari2600.ram[58][1] ),
    .A2(net4885),
    .A1(\atari2600.ram[57][1] ));
 sg13g2_a21oi_1 _17115_ (.A1(_08866_),
    .A2(_08867_),
    .Y(_08868_),
    .B1(net4937));
 sg13g2_nor2_1 _17116_ (.A(net5025),
    .B(_08865_),
    .Y(_08869_));
 sg13g2_nor3_2 _17117_ (.A(_08859_),
    .B(_08862_),
    .C(_08868_),
    .Y(_08870_));
 sg13g2_a22oi_1 _17118_ (.Y(_08871_),
    .B1(net4839),
    .B2(\atari2600.ram[43][1] ),
    .A2(net4969),
    .A1(\atari2600.ram[40][1] ));
 sg13g2_a22oi_1 _17119_ (.Y(_08872_),
    .B1(net4793),
    .B2(\atari2600.ram[42][1] ),
    .A2(net4882),
    .A1(\atari2600.ram[41][1] ));
 sg13g2_a21oi_1 _17120_ (.A1(_08871_),
    .A2(_08872_),
    .Y(_08873_),
    .B1(net4937));
 sg13g2_a22oi_1 _17121_ (.Y(_08874_),
    .B1(net4833),
    .B2(\atari2600.ram[47][1] ),
    .A2(net4963),
    .A1(\atari2600.ram[44][1] ));
 sg13g2_a22oi_1 _17122_ (.Y(_08875_),
    .B1(net4788),
    .B2(\atari2600.ram[46][1] ),
    .A2(net4882),
    .A1(\atari2600.ram[45][1] ));
 sg13g2_a21o_1 _17123_ (.A2(_08875_),
    .A1(_08874_),
    .B1(net4949),
    .X(_08876_));
 sg13g2_a22oi_1 _17124_ (.Y(_08877_),
    .B1(net4837),
    .B2(\atari2600.ram[35][1] ),
    .A2(net4967),
    .A1(\atari2600.ram[32][1] ));
 sg13g2_a22oi_1 _17125_ (.Y(_08878_),
    .B1(net4791),
    .B2(\atari2600.ram[34][1] ),
    .A2(net4885),
    .A1(\atari2600.ram[33][1] ));
 sg13g2_a21oi_1 _17126_ (.A1(_08877_),
    .A2(_08878_),
    .Y(_08879_),
    .B1(net4925));
 sg13g2_a22oi_1 _17127_ (.Y(_08880_),
    .B1(net4960),
    .B2(\atari2600.ram[36][1] ),
    .A2(net4880),
    .A1(\atari2600.ram[37][1] ));
 sg13g2_a22oi_1 _17128_ (.Y(_08881_),
    .B1(net4785),
    .B2(\atari2600.ram[38][1] ),
    .A2(net4830),
    .A1(\atari2600.ram[39][1] ));
 sg13g2_a21oi_2 _17129_ (.B1(net5006),
    .Y(_08882_),
    .A2(_08881_),
    .A1(_08880_));
 sg13g2_nor4_1 _17130_ (.A(net5027),
    .B(_08873_),
    .C(_08879_),
    .D(_08882_),
    .Y(_08883_));
 sg13g2_a221oi_1 _17131_ (.B2(_08883_),
    .C1(net4876),
    .B1(_08876_),
    .A1(_08869_),
    .Y(_08884_),
    .A2(_08870_));
 sg13g2_a22oi_1 _17132_ (.Y(_08885_),
    .B1(net4836),
    .B2(\atari2600.ram[11][1] ),
    .A2(net4966),
    .A1(\atari2600.ram[8][1] ));
 sg13g2_a22oi_1 _17133_ (.Y(_08886_),
    .B1(net4790),
    .B2(\atari2600.ram[10][1] ),
    .A2(net4884),
    .A1(\atari2600.ram[9][1] ));
 sg13g2_a21oi_2 _17134_ (.B1(net4938),
    .Y(_08887_),
    .A2(_08886_),
    .A1(_08885_));
 sg13g2_a22oi_1 _17135_ (.Y(_08888_),
    .B1(net4835),
    .B2(\atari2600.ram[15][1] ),
    .A2(net4965),
    .A1(\atari2600.ram[12][1] ));
 sg13g2_a22oi_1 _17136_ (.Y(_08889_),
    .B1(net4789),
    .B2(\atari2600.ram[14][1] ),
    .A2(net4883),
    .A1(\atari2600.ram[13][1] ));
 sg13g2_a21oi_2 _17137_ (.B1(net4950),
    .Y(_08890_),
    .A2(_08889_),
    .A1(_08888_));
 sg13g2_a22oi_1 _17138_ (.Y(_08891_),
    .B1(net4844),
    .B2(\atari2600.ram[3][1] ),
    .A2(net4974),
    .A1(\atari2600.ram[0][1] ));
 sg13g2_a22oi_1 _17139_ (.Y(_08892_),
    .B1(net4798),
    .B2(\atari2600.ram[2][1] ),
    .A2(net4894),
    .A1(\atari2600.ram[1][1] ));
 sg13g2_a21oi_2 _17140_ (.B1(net4927),
    .Y(_08893_),
    .A2(_08892_),
    .A1(_08891_));
 sg13g2_a22oi_1 _17141_ (.Y(_08894_),
    .B1(net4843),
    .B2(\atari2600.ram[7][1] ),
    .A2(net4973),
    .A1(\atari2600.ram[4][1] ));
 sg13g2_a22oi_1 _17142_ (.Y(_08895_),
    .B1(net4799),
    .B2(\atari2600.ram[6][1] ),
    .A2(net4893),
    .A1(\atari2600.ram[5][1] ));
 sg13g2_a21oi_1 _17143_ (.A1(_08894_),
    .A2(_08895_),
    .Y(_08896_),
    .B1(net5010));
 sg13g2_nor4_2 _17144_ (.A(_08887_),
    .B(_08890_),
    .C(_08893_),
    .Y(_08897_),
    .D(_08896_));
 sg13g2_a22oi_1 _17145_ (.Y(_08898_),
    .B1(net4848),
    .B2(\atari2600.ram[23][1] ),
    .A2(net4979),
    .A1(\atari2600.ram[20][1] ));
 sg13g2_a22oi_1 _17146_ (.Y(_08899_),
    .B1(net4802),
    .B2(\atari2600.ram[22][1] ),
    .A2(net4897),
    .A1(\atari2600.ram[21][1] ));
 sg13g2_a21oi_1 _17147_ (.A1(_08898_),
    .A2(_08899_),
    .Y(_08900_),
    .B1(net5008));
 sg13g2_a22oi_1 _17148_ (.Y(_08901_),
    .B1(net4849),
    .B2(\atari2600.ram[19][1] ),
    .A2(net4975),
    .A1(\atari2600.ram[16][1] ));
 sg13g2_a22oi_1 _17149_ (.Y(_08902_),
    .B1(net4800),
    .B2(\atari2600.ram[18][1] ),
    .A2(net4895),
    .A1(\atari2600.ram[17][1] ));
 sg13g2_a21oi_2 _17150_ (.B1(net4928),
    .Y(_08903_),
    .A2(_08902_),
    .A1(_08901_));
 sg13g2_a22oi_1 _17151_ (.Y(_08904_),
    .B1(net4846),
    .B2(\atari2600.ram[27][1] ),
    .A2(net4976),
    .A1(\atari2600.ram[24][1] ));
 sg13g2_a22oi_1 _17152_ (.Y(_08905_),
    .B1(net4801),
    .B2(\atari2600.ram[26][1] ),
    .A2(net4896),
    .A1(\atari2600.ram[25][1] ));
 sg13g2_a21oi_2 _17153_ (.B1(net4941),
    .Y(_08906_),
    .A2(_08905_),
    .A1(_08904_));
 sg13g2_a22oi_1 _17154_ (.Y(_08907_),
    .B1(net4851),
    .B2(\atari2600.ram[31][1] ),
    .A2(net4981),
    .A1(\atari2600.ram[28][1] ));
 sg13g2_a22oi_1 _17155_ (.Y(_08908_),
    .B1(net4804),
    .B2(\atari2600.ram[30][1] ),
    .A2(net4899),
    .A1(\atari2600.ram[29][1] ));
 sg13g2_a21oi_1 _17156_ (.A1(_08907_),
    .A2(_08908_),
    .Y(_08909_),
    .B1(net4952));
 sg13g2_nor4_2 _17157_ (.A(_08900_),
    .B(_08903_),
    .C(_08906_),
    .Y(_08910_),
    .D(_08909_));
 sg13g2_nor2_1 _17158_ (.A(net4773),
    .B(_08910_),
    .Y(_08911_));
 sg13g2_o21ai_1 _17159_ (.B1(net5023),
    .Y(_08912_),
    .A1(net4780),
    .A2(_08897_));
 sg13g2_nor3_1 _17160_ (.A(_08884_),
    .B(_08911_),
    .C(_08912_),
    .Y(_08913_));
 sg13g2_a22oi_1 _17161_ (.Y(_08914_),
    .B1(net4856),
    .B2(\atari2600.ram[123][1] ),
    .A2(net4988),
    .A1(\atari2600.ram[120][1] ));
 sg13g2_a22oi_1 _17162_ (.Y(_08915_),
    .B1(net4809),
    .B2(\atari2600.ram[122][1] ),
    .A2(net4905),
    .A1(\atari2600.ram[121][1] ));
 sg13g2_a21oi_1 _17163_ (.A1(_08914_),
    .A2(_08915_),
    .Y(_08916_),
    .B1(net4943));
 sg13g2_a22oi_1 _17164_ (.Y(_08917_),
    .B1(net4865),
    .B2(\atari2600.ram[127][1] ),
    .A2(net4999),
    .A1(\atari2600.ram[124][1] ));
 sg13g2_a22oi_1 _17165_ (.Y(_08918_),
    .B1(net4819),
    .B2(\atari2600.ram[126][1] ),
    .A2(net4914),
    .A1(\atari2600.ram[125][1] ));
 sg13g2_a21oi_1 _17166_ (.A1(_08917_),
    .A2(_08918_),
    .Y(_08919_),
    .B1(net4958));
 sg13g2_a22oi_1 _17167_ (.Y(_08920_),
    .B1(net4986),
    .B2(\atari2600.ram[116][1] ),
    .A2(net4907),
    .A1(\atari2600.ram[117][1] ));
 sg13g2_a22oi_1 _17168_ (.Y(_08921_),
    .B1(net4812),
    .B2(\atari2600.ram[118][1] ),
    .A2(net4857),
    .A1(\atari2600.ram[119][1] ));
 sg13g2_a21oi_1 _17169_ (.A1(_08920_),
    .A2(_08921_),
    .Y(_08922_),
    .B1(net5013));
 sg13g2_a22oi_1 _17170_ (.Y(_08923_),
    .B1(net4854),
    .B2(\atari2600.ram[115][1] ),
    .A2(net4984),
    .A1(\atari2600.ram[112][1] ));
 sg13g2_a22oi_1 _17171_ (.Y(_08924_),
    .B1(net4810),
    .B2(\atari2600.ram[114][1] ),
    .A2(net4904),
    .A1(\atari2600.ram[113][1] ));
 sg13g2_a21oi_1 _17172_ (.A1(_08923_),
    .A2(_08924_),
    .Y(_08925_),
    .B1(net4930));
 sg13g2_nor2_1 _17173_ (.A(net5026),
    .B(_08919_),
    .Y(_08926_));
 sg13g2_nor3_1 _17174_ (.A(_08916_),
    .B(_08922_),
    .C(_08925_),
    .Y(_08927_));
 sg13g2_a22oi_1 _17175_ (.Y(_08928_),
    .B1(net4854),
    .B2(\atari2600.ram[99][1] ),
    .A2(net4984),
    .A1(\atari2600.ram[96][1] ));
 sg13g2_a22oi_1 _17176_ (.Y(_08929_),
    .B1(net4809),
    .B2(\atari2600.ram[98][1] ),
    .A2(net4903),
    .A1(\atari2600.ram[97][1] ));
 sg13g2_a21oi_1 _17177_ (.A1(_08928_),
    .A2(_08929_),
    .Y(_08930_),
    .B1(net4931));
 sg13g2_a22oi_1 _17178_ (.Y(_08931_),
    .B1(net4856),
    .B2(\atari2600.ram[111][1] ),
    .A2(net4987),
    .A1(\atari2600.ram[108][1] ));
 sg13g2_a22oi_1 _17179_ (.Y(_08932_),
    .B1(net4811),
    .B2(\atari2600.ram[110][1] ),
    .A2(net4905),
    .A1(\atari2600.ram[109][1] ));
 sg13g2_a21o_1 _17180_ (.A2(_08932_),
    .A1(_08931_),
    .B1(net4956),
    .X(_08933_));
 sg13g2_a22oi_1 _17181_ (.Y(_08934_),
    .B1(net4985),
    .B2(\atari2600.ram[100][1] ),
    .A2(net4903),
    .A1(\atari2600.ram[101][1] ));
 sg13g2_a22oi_1 _17182_ (.Y(_08935_),
    .B1(net4809),
    .B2(\atari2600.ram[102][1] ),
    .A2(net4854),
    .A1(\atari2600.ram[103][1] ));
 sg13g2_a21oi_1 _17183_ (.A1(_08934_),
    .A2(_08935_),
    .Y(_08936_),
    .B1(net5012));
 sg13g2_a22oi_1 _17184_ (.Y(_08937_),
    .B1(net4860),
    .B2(\atari2600.ram[107][1] ),
    .A2(net4990),
    .A1(\atari2600.ram[104][1] ));
 sg13g2_a22oi_1 _17185_ (.Y(_08938_),
    .B1(net4815),
    .B2(\atari2600.ram[106][1] ),
    .A2(net4909),
    .A1(\atari2600.ram[105][1] ));
 sg13g2_a21oi_2 _17186_ (.B1(net4946),
    .Y(_08939_),
    .A2(_08938_),
    .A1(_08937_));
 sg13g2_nor4_2 _17187_ (.A(net5028),
    .B(_08930_),
    .C(_08936_),
    .Y(_08940_),
    .D(_08939_));
 sg13g2_a221oi_1 _17188_ (.B2(_08940_),
    .C1(net4879),
    .B1(_08933_),
    .A1(_08926_),
    .Y(_08941_),
    .A2(_08927_));
 sg13g2_a22oi_1 _17189_ (.Y(_08942_),
    .B1(net4871),
    .B2(\atari2600.ram[79][1] ),
    .A2(net5002),
    .A1(\atari2600.ram[76][1] ));
 sg13g2_a22oi_1 _17190_ (.Y(_08943_),
    .B1(net4827),
    .B2(\atari2600.ram[78][1] ),
    .A2(net4922),
    .A1(\atari2600.ram[77][1] ));
 sg13g2_a21oi_2 _17191_ (.B1(net4959),
    .Y(_08944_),
    .A2(_08943_),
    .A1(_08942_));
 sg13g2_a22oi_1 _17192_ (.Y(_08945_),
    .B1(net4869),
    .B2(\atari2600.ram[67][1] ),
    .A2(net5001),
    .A1(\atari2600.ram[64][1] ));
 sg13g2_a22oi_1 _17193_ (.Y(_08946_),
    .B1(net4818),
    .B2(\atari2600.ram[66][1] ),
    .A2(net4913),
    .A1(\atari2600.ram[65][1] ));
 sg13g2_a21oi_1 _17194_ (.A1(_08945_),
    .A2(_08946_),
    .Y(_08947_),
    .B1(net4933));
 sg13g2_a22oi_1 _17195_ (.Y(_08948_),
    .B1(net4871),
    .B2(\atari2600.ram[75][1] ),
    .A2(net5002),
    .A1(\atari2600.ram[72][1] ));
 sg13g2_a22oi_1 _17196_ (.Y(_08949_),
    .B1(net4827),
    .B2(\atari2600.ram[74][1] ),
    .A2(net4922),
    .A1(\atari2600.ram[73][1] ));
 sg13g2_a21oi_1 _17197_ (.A1(_08948_),
    .A2(_08949_),
    .Y(_08950_),
    .B1(net4945));
 sg13g2_a22oi_1 _17198_ (.Y(_08951_),
    .B1(net4869),
    .B2(\atari2600.ram[71][1] ),
    .A2(net5000),
    .A1(\atari2600.ram[68][1] ));
 sg13g2_a22oi_1 _17199_ (.Y(_08952_),
    .B1(net4825),
    .B2(\atari2600.ram[70][1] ),
    .A2(net4920),
    .A1(\atari2600.ram[69][1] ));
 sg13g2_a21oi_1 _17200_ (.A1(_08951_),
    .A2(_08952_),
    .Y(_08953_),
    .B1(net5015));
 sg13g2_nor4_1 _17201_ (.A(_08944_),
    .B(_08947_),
    .C(_08950_),
    .D(_08953_),
    .Y(_08954_));
 sg13g2_nor2_1 _17202_ (.A(net4778),
    .B(_08954_),
    .Y(_08955_));
 sg13g2_a22oi_1 _17203_ (.Y(_08956_),
    .B1(net4850),
    .B2(\atari2600.ram[91][1] ),
    .A2(net4981),
    .A1(\atari2600.ram[88][1] ));
 sg13g2_a22oi_1 _17204_ (.Y(_08957_),
    .B1(net4821),
    .B2(\atari2600.ram[90][1] ),
    .A2(net4916),
    .A1(\atari2600.ram[89][1] ));
 sg13g2_a21oi_2 _17205_ (.B1(net4942),
    .Y(_08958_),
    .A2(_08957_),
    .A1(_08956_));
 sg13g2_a22oi_1 _17206_ (.Y(_08959_),
    .B1(net4867),
    .B2(\atari2600.ram[95][1] ),
    .A2(net4997),
    .A1(\atari2600.ram[92][1] ));
 sg13g2_a22oi_1 _17207_ (.Y(_08960_),
    .B1(net4822),
    .B2(\atari2600.ram[94][1] ),
    .A2(net4917),
    .A1(\atari2600.ram[93][1] ));
 sg13g2_a21oi_2 _17208_ (.B1(net4957),
    .Y(_08961_),
    .A2(_08960_),
    .A1(_08959_));
 sg13g2_a22oi_1 _17209_ (.Y(_08962_),
    .B1(net4864),
    .B2(\atari2600.ram[83][1] ),
    .A2(net4995),
    .A1(\atari2600.ram[80][1] ));
 sg13g2_a22oi_1 _17210_ (.Y(_08963_),
    .B1(net4820),
    .B2(\atari2600.ram[82][1] ),
    .A2(net4915),
    .A1(\atari2600.ram[81][1] ));
 sg13g2_a21oi_1 _17211_ (.A1(_08962_),
    .A2(_08963_),
    .Y(_08964_),
    .B1(net4934));
 sg13g2_a22oi_1 _17212_ (.Y(_08965_),
    .B1(net4847),
    .B2(\atari2600.ram[87][1] ),
    .A2(net4977),
    .A1(\atari2600.ram[84][1] ));
 sg13g2_a22oi_1 _17213_ (.Y(_08966_),
    .B1(net4803),
    .B2(\atari2600.ram[86][1] ),
    .A2(net4898),
    .A1(\atari2600.ram[85][1] ));
 sg13g2_a21oi_2 _17214_ (.B1(net5009),
    .Y(_08967_),
    .A2(_08966_),
    .A1(_08965_));
 sg13g2_nor4_2 _17215_ (.A(_08958_),
    .B(_08961_),
    .C(_08964_),
    .Y(_08968_),
    .D(_08967_));
 sg13g2_o21ai_1 _17216_ (.B1(net5020),
    .Y(_08969_),
    .A1(net4774),
    .A2(_08968_));
 sg13g2_nor3_2 _17217_ (.A(_08941_),
    .B(_08955_),
    .C(_08969_),
    .Y(_08970_));
 sg13g2_nor2_2 _17218_ (.A(_08913_),
    .B(_08970_),
    .Y(_00002_));
 sg13g2_a22oi_1 _17219_ (.Y(_08971_),
    .B1(net4837),
    .B2(\atari2600.ram[63][2] ),
    .A2(net4967),
    .A1(\atari2600.ram[60][2] ));
 sg13g2_a22oi_1 _17220_ (.Y(_08972_),
    .B1(net4791),
    .B2(\atari2600.ram[62][2] ),
    .A2(net4885),
    .A1(\atari2600.ram[61][2] ));
 sg13g2_a21oi_1 _17221_ (.A1(_08971_),
    .A2(_08972_),
    .Y(_08973_),
    .B1(net4951));
 sg13g2_a22oi_1 _17222_ (.Y(_08974_),
    .B1(net4837),
    .B2(\atari2600.ram[59][2] ),
    .A2(net4967),
    .A1(\atari2600.ram[56][2] ));
 sg13g2_a22oi_1 _17223_ (.Y(_08975_),
    .B1(net4791),
    .B2(\atari2600.ram[58][2] ),
    .A2(net4885),
    .A1(\atari2600.ram[57][2] ));
 sg13g2_a21oi_1 _17224_ (.A1(_08974_),
    .A2(_08975_),
    .Y(_08976_),
    .B1(net4937));
 sg13g2_a22oi_1 _17225_ (.Y(_08977_),
    .B1(net4840),
    .B2(\atari2600.ram[51][2] ),
    .A2(net4970),
    .A1(\atari2600.ram[48][2] ));
 sg13g2_a22oi_1 _17226_ (.Y(_08978_),
    .B1(net4795),
    .B2(\atari2600.ram[50][2] ),
    .A2(net4889),
    .A1(\atari2600.ram[49][2] ));
 sg13g2_a21oi_1 _17227_ (.A1(_08977_),
    .A2(_08978_),
    .Y(_08979_),
    .B1(net4926));
 sg13g2_a22oi_1 _17228_ (.Y(_08980_),
    .B1(net4983),
    .B2(\atari2600.ram[52][2] ),
    .A2(net4902),
    .A1(\atari2600.ram[53][2] ));
 sg13g2_a22oi_1 _17229_ (.Y(_08981_),
    .B1(net4808),
    .B2(\atari2600.ram[54][2] ),
    .A2(net4853),
    .A1(\atari2600.ram[55][2] ));
 sg13g2_a21oi_2 _17230_ (.B1(net5012),
    .Y(_08982_),
    .A2(_08981_),
    .A1(_08980_));
 sg13g2_nor2_1 _17231_ (.A(net5025),
    .B(_08979_),
    .Y(_08983_));
 sg13g2_nor3_2 _17232_ (.A(_08973_),
    .B(_08976_),
    .C(_08982_),
    .Y(_08984_));
 sg13g2_a22oi_1 _17233_ (.Y(_08985_),
    .B1(net4830),
    .B2(\atari2600.ram[47][2] ),
    .A2(net4960),
    .A1(\atari2600.ram[44][2] ));
 sg13g2_a22oi_1 _17234_ (.Y(_08986_),
    .B1(net4786),
    .B2(\atari2600.ram[46][2] ),
    .A2(net4883),
    .A1(\atari2600.ram[45][2] ));
 sg13g2_a21oi_1 _17235_ (.A1(_08985_),
    .A2(_08986_),
    .Y(_08987_),
    .B1(net4949));
 sg13g2_a22oi_1 _17236_ (.Y(_08988_),
    .B1(net4832),
    .B2(\atari2600.ram[35][2] ),
    .A2(net4962),
    .A1(\atari2600.ram[32][2] ));
 sg13g2_a22oi_1 _17237_ (.Y(_08989_),
    .B1(net4787),
    .B2(\atari2600.ram[34][2] ),
    .A2(net4881),
    .A1(\atari2600.ram[33][2] ));
 sg13g2_a21oi_1 _17238_ (.A1(_08988_),
    .A2(_08989_),
    .Y(_08990_),
    .B1(net4925));
 sg13g2_a22oi_1 _17239_ (.Y(_08991_),
    .B1(net4840),
    .B2(\atari2600.ram[43][2] ),
    .A2(net4970),
    .A1(\atari2600.ram[40][2] ));
 sg13g2_a22oi_1 _17240_ (.Y(_08992_),
    .B1(net4795),
    .B2(\atari2600.ram[42][2] ),
    .A2(net4889),
    .A1(\atari2600.ram[41][2] ));
 sg13g2_a21o_1 _17241_ (.A2(_08992_),
    .A1(_08991_),
    .B1(net4938),
    .X(_08993_));
 sg13g2_a22oi_1 _17242_ (.Y(_08994_),
    .B1(net4960),
    .B2(\atari2600.ram[36][2] ),
    .A2(net4880),
    .A1(\atari2600.ram[37][2] ));
 sg13g2_a22oi_1 _17243_ (.Y(_08995_),
    .B1(net4785),
    .B2(\atari2600.ram[38][2] ),
    .A2(net4830),
    .A1(\atari2600.ram[39][2] ));
 sg13g2_a21oi_1 _17244_ (.A1(_08994_),
    .A2(_08995_),
    .Y(_08996_),
    .B1(net5006));
 sg13g2_nor4_2 _17245_ (.A(net5027),
    .B(_08987_),
    .C(_08990_),
    .Y(_08997_),
    .D(_08996_));
 sg13g2_a221oi_1 _17246_ (.B2(_08997_),
    .C1(net4876),
    .B1(_08993_),
    .A1(_08983_),
    .Y(_08998_),
    .A2(_08984_));
 sg13g2_a22oi_1 _17247_ (.Y(_08999_),
    .B1(net4845),
    .B2(\atari2600.ram[19][2] ),
    .A2(net4975),
    .A1(\atari2600.ram[16][2] ));
 sg13g2_a22oi_1 _17248_ (.Y(_09000_),
    .B1(net4800),
    .B2(\atari2600.ram[18][2] ),
    .A2(net4895),
    .A1(\atari2600.ram[17][2] ));
 sg13g2_a21oi_2 _17249_ (.B1(net4928),
    .Y(_09001_),
    .A2(_09000_),
    .A1(_08999_));
 sg13g2_a22oi_1 _17250_ (.Y(_09002_),
    .B1(net4849),
    .B2(\atari2600.ram[31][2] ),
    .A2(net4980),
    .A1(\atari2600.ram[28][2] ));
 sg13g2_a22oi_1 _17251_ (.Y(_09003_),
    .B1(net4802),
    .B2(\atari2600.ram[30][2] ),
    .A2(net4897),
    .A1(\atari2600.ram[29][2] ));
 sg13g2_a21oi_1 _17252_ (.A1(_09002_),
    .A2(_09003_),
    .Y(_09004_),
    .B1(net4952));
 sg13g2_a22oi_1 _17253_ (.Y(_09005_),
    .B1(net4840),
    .B2(\atari2600.ram[27][2] ),
    .A2(net4970),
    .A1(\atari2600.ram[24][2] ));
 sg13g2_a22oi_1 _17254_ (.Y(_09006_),
    .B1(net4795),
    .B2(\atari2600.ram[26][2] ),
    .A2(net4889),
    .A1(\atari2600.ram[25][2] ));
 sg13g2_a21oi_2 _17255_ (.B1(net4939),
    .Y(_09007_),
    .A2(_09006_),
    .A1(_09005_));
 sg13g2_a22oi_1 _17256_ (.Y(_09008_),
    .B1(net4845),
    .B2(\atari2600.ram[23][2] ),
    .A2(net4975),
    .A1(\atari2600.ram[20][2] ));
 sg13g2_a22oi_1 _17257_ (.Y(_09009_),
    .B1(net4800),
    .B2(\atari2600.ram[22][2] ),
    .A2(net4895),
    .A1(\atari2600.ram[21][2] ));
 sg13g2_a21oi_1 _17258_ (.A1(_09008_),
    .A2(_09009_),
    .Y(_09010_),
    .B1(net5010));
 sg13g2_nor4_2 _17259_ (.A(_09001_),
    .B(_09004_),
    .C(_09007_),
    .Y(_09011_),
    .D(_09010_));
 sg13g2_nor2_1 _17260_ (.A(net4773),
    .B(_09011_),
    .Y(_09012_));
 sg13g2_a22oi_1 _17261_ (.Y(_09013_),
    .B1(net4844),
    .B2(\atari2600.ram[3][2] ),
    .A2(net4974),
    .A1(\atari2600.ram[0][2] ));
 sg13g2_a22oi_1 _17262_ (.Y(_09014_),
    .B1(net4807),
    .B2(\atari2600.ram[2][2] ),
    .A2(net4901),
    .A1(\atari2600.ram[1][2] ));
 sg13g2_a21oi_1 _17263_ (.A1(_09013_),
    .A2(_09014_),
    .Y(_09015_),
    .B1(net4927));
 sg13g2_a22oi_1 _17264_ (.Y(_09016_),
    .B1(net4835),
    .B2(\atari2600.ram[15][2] ),
    .A2(net4965),
    .A1(\atari2600.ram[12][2] ));
 sg13g2_a22oi_1 _17265_ (.Y(_09017_),
    .B1(net4789),
    .B2(\atari2600.ram[14][2] ),
    .A2(net4883),
    .A1(\atari2600.ram[13][2] ));
 sg13g2_a21oi_1 _17266_ (.A1(_09016_),
    .A2(_09017_),
    .Y(_09018_),
    .B1(net4950));
 sg13g2_a22oi_1 _17267_ (.Y(_09019_),
    .B1(net4834),
    .B2(\atari2600.ram[11][2] ),
    .A2(net4964),
    .A1(\atari2600.ram[8][2] ));
 sg13g2_a22oi_1 _17268_ (.Y(_09020_),
    .B1(net4798),
    .B2(\atari2600.ram[10][2] ),
    .A2(net4892),
    .A1(\atari2600.ram[9][2] ));
 sg13g2_a21oi_1 _17269_ (.A1(_09019_),
    .A2(_09020_),
    .Y(_09021_),
    .B1(net4941));
 sg13g2_a22oi_1 _17270_ (.Y(_09022_),
    .B1(net4843),
    .B2(\atari2600.ram[7][2] ),
    .A2(net4973),
    .A1(\atari2600.ram[4][2] ));
 sg13g2_a22oi_1 _17271_ (.Y(_09023_),
    .B1(net4799),
    .B2(\atari2600.ram[6][2] ),
    .A2(net4893),
    .A1(\atari2600.ram[5][2] ));
 sg13g2_a21oi_1 _17272_ (.A1(_09022_),
    .A2(_09023_),
    .Y(_09024_),
    .B1(net5007));
 sg13g2_nor4_1 _17273_ (.A(_09015_),
    .B(_09018_),
    .C(_09021_),
    .D(_09024_),
    .Y(_09025_));
 sg13g2_o21ai_1 _17274_ (.B1(net5023),
    .Y(_09026_),
    .A1(net4777),
    .A2(_09025_));
 sg13g2_nor3_1 _17275_ (.A(_08998_),
    .B(_09012_),
    .C(_09026_),
    .Y(_09027_));
 sg13g2_a22oi_1 _17276_ (.Y(_09028_),
    .B1(net4857),
    .B2(\atari2600.ram[119][2] ),
    .A2(net4987),
    .A1(\atari2600.ram[116][2] ));
 sg13g2_a22oi_1 _17277_ (.Y(_09029_),
    .B1(net4812),
    .B2(\atari2600.ram[118][2] ),
    .A2(net4907),
    .A1(\atari2600.ram[117][2] ));
 sg13g2_a21oi_1 _17278_ (.A1(_09028_),
    .A2(_09029_),
    .Y(_09030_),
    .B1(net5016));
 sg13g2_a22oi_1 _17279_ (.Y(_09031_),
    .B1(net4851),
    .B2(\atari2600.ram[127][2] ),
    .A2(net4977),
    .A1(\atari2600.ram[124][2] ));
 sg13g2_a22oi_1 _17280_ (.Y(_09032_),
    .B1(net4818),
    .B2(\atari2600.ram[126][2] ),
    .A2(net4913),
    .A1(\atari2600.ram[125][2] ));
 sg13g2_a21oi_1 _17281_ (.A1(_09031_),
    .A2(_09032_),
    .Y(_09033_),
    .B1(net4958));
 sg13g2_a22oi_1 _17282_ (.Y(_09034_),
    .B1(net4858),
    .B2(\atari2600.ram[123][2] ),
    .A2(net4986),
    .A1(\atari2600.ram[120][2] ));
 sg13g2_a22oi_1 _17283_ (.Y(_09035_),
    .B1(net4811),
    .B2(\atari2600.ram[122][2] ),
    .A2(net4906),
    .A1(\atari2600.ram[121][2] ));
 sg13g2_a21oi_1 _17284_ (.A1(_09034_),
    .A2(_09035_),
    .Y(_09036_),
    .B1(net4944));
 sg13g2_a22oi_1 _17285_ (.Y(_09037_),
    .B1(net4853),
    .B2(\atari2600.ram[115][2] ),
    .A2(net4983),
    .A1(\atari2600.ram[112][2] ));
 sg13g2_a22oi_1 _17286_ (.Y(_09038_),
    .B1(net4808),
    .B2(\atari2600.ram[114][2] ),
    .A2(net4902),
    .A1(\atari2600.ram[113][2] ));
 sg13g2_a21oi_2 _17287_ (.B1(net4930),
    .Y(_09039_),
    .A2(_09038_),
    .A1(_09037_));
 sg13g2_nor4_1 _17288_ (.A(_09030_),
    .B(_09033_),
    .C(_09036_),
    .D(_09039_),
    .Y(_09040_));
 sg13g2_nor2_1 _17289_ (.A(_08729_),
    .B(_09040_),
    .Y(_09041_));
 sg13g2_a22oi_1 _17290_ (.Y(_09042_),
    .B1(net4867),
    .B2(\atari2600.ram[83][2] ),
    .A2(net4997),
    .A1(\atari2600.ram[80][2] ));
 sg13g2_a22oi_1 _17291_ (.Y(_09043_),
    .B1(net4820),
    .B2(\atari2600.ram[82][2] ),
    .A2(net4915),
    .A1(\atari2600.ram[81][2] ));
 sg13g2_a21oi_1 _17292_ (.A1(_09042_),
    .A2(_09043_),
    .Y(_09044_),
    .B1(net4934));
 sg13g2_a22oi_1 _17293_ (.Y(_09045_),
    .B1(net4864),
    .B2(\atari2600.ram[87][2] ),
    .A2(net4995),
    .A1(\atari2600.ram[84][2] ));
 sg13g2_a22oi_1 _17294_ (.Y(_09046_),
    .B1(net4820),
    .B2(\atari2600.ram[86][2] ),
    .A2(net4915),
    .A1(\atari2600.ram[85][2] ));
 sg13g2_a21oi_1 _17295_ (.A1(_09045_),
    .A2(_09046_),
    .Y(_09047_),
    .B1(net5016));
 sg13g2_a22oi_1 _17296_ (.Y(_09048_),
    .B1(net4850),
    .B2(\atari2600.ram[91][2] ),
    .A2(net4980),
    .A1(\atari2600.ram[88][2] ));
 sg13g2_a22oi_1 _17297_ (.Y(_09049_),
    .B1(net4804),
    .B2(\atari2600.ram[90][2] ),
    .A2(net4899),
    .A1(\atari2600.ram[89][2] ));
 sg13g2_a21oi_2 _17298_ (.B1(net4942),
    .Y(_09050_),
    .A2(_09049_),
    .A1(_09048_));
 sg13g2_a22oi_1 _17299_ (.Y(_09051_),
    .B1(net4867),
    .B2(\atari2600.ram[95][2] ),
    .A2(net4997),
    .A1(\atari2600.ram[92][2] ));
 sg13g2_a22oi_1 _17300_ (.Y(_09052_),
    .B1(net4822),
    .B2(\atari2600.ram[94][2] ),
    .A2(net4917),
    .A1(\atari2600.ram[93][2] ));
 sg13g2_a21oi_2 _17301_ (.B1(net4957),
    .Y(_09053_),
    .A2(_09052_),
    .A1(_09051_));
 sg13g2_nor4_2 _17302_ (.A(_09044_),
    .B(_09047_),
    .C(_09050_),
    .Y(_09054_),
    .D(_09053_));
 sg13g2_a22oi_1 _17303_ (.Y(_09055_),
    .B1(net4870),
    .B2(\atari2600.ram[67][2] ),
    .A2(net5000),
    .A1(\atari2600.ram[64][2] ));
 sg13g2_a22oi_1 _17304_ (.Y(_09056_),
    .B1(net4826),
    .B2(\atari2600.ram[66][2] ),
    .A2(net4921),
    .A1(\atari2600.ram[65][2] ));
 sg13g2_a21oi_1 _17305_ (.A1(_09055_),
    .A2(_09056_),
    .Y(_09057_),
    .B1(net4934));
 sg13g2_a22oi_1 _17306_ (.Y(_09058_),
    .B1(net4871),
    .B2(\atari2600.ram[75][2] ),
    .A2(net5002),
    .A1(\atari2600.ram[72][2] ));
 sg13g2_a22oi_1 _17307_ (.Y(_09059_),
    .B1(net4828),
    .B2(\atari2600.ram[74][2] ),
    .A2(net4923),
    .A1(\atari2600.ram[73][2] ));
 sg13g2_a21oi_1 _17308_ (.A1(_09058_),
    .A2(_09059_),
    .Y(_09060_),
    .B1(net4945));
 sg13g2_a22oi_1 _17309_ (.Y(_09061_),
    .B1(net4870),
    .B2(\atari2600.ram[71][2] ),
    .A2(net5001),
    .A1(\atari2600.ram[68][2] ));
 sg13g2_a22oi_1 _17310_ (.Y(_09062_),
    .B1(net4826),
    .B2(\atari2600.ram[70][2] ),
    .A2(net4921),
    .A1(\atari2600.ram[69][2] ));
 sg13g2_a21oi_1 _17311_ (.A1(_09061_),
    .A2(_09062_),
    .Y(_09063_),
    .B1(net5016));
 sg13g2_a22oi_1 _17312_ (.Y(_09064_),
    .B1(net4872),
    .B2(\atari2600.ram[79][2] ),
    .A2(net5003),
    .A1(\atari2600.ram[76][2] ));
 sg13g2_a22oi_1 _17313_ (.Y(_09065_),
    .B1(net4827),
    .B2(\atari2600.ram[78][2] ),
    .A2(net4922),
    .A1(\atari2600.ram[77][2] ));
 sg13g2_a21oi_2 _17314_ (.B1(net4959),
    .Y(_09066_),
    .A2(_09065_),
    .A1(_09064_));
 sg13g2_nor4_2 _17315_ (.A(_09057_),
    .B(_09060_),
    .C(_09063_),
    .Y(_09067_),
    .D(_09066_));
 sg13g2_nor2_1 _17316_ (.A(net4779),
    .B(_09067_),
    .Y(_09068_));
 sg13g2_a22oi_1 _17317_ (.Y(_09069_),
    .B1(net4860),
    .B2(\atari2600.ram[103][2] ),
    .A2(net4990),
    .A1(\atari2600.ram[100][2] ));
 sg13g2_a22oi_1 _17318_ (.Y(_09070_),
    .B1(net4814),
    .B2(\atari2600.ram[102][2] ),
    .A2(net4909),
    .A1(\atari2600.ram[101][2] ));
 sg13g2_a21oi_1 _17319_ (.A1(_09069_),
    .A2(_09070_),
    .Y(_09071_),
    .B1(net5014));
 sg13g2_a22oi_1 _17320_ (.Y(_09072_),
    .B1(net4861),
    .B2(\atari2600.ram[111][2] ),
    .A2(net4991),
    .A1(\atari2600.ram[108][2] ));
 sg13g2_a22oi_1 _17321_ (.Y(_09073_),
    .B1(net4816),
    .B2(\atari2600.ram[110][2] ),
    .A2(net4910),
    .A1(\atari2600.ram[109][2] ));
 sg13g2_a21oi_2 _17322_ (.B1(net4954),
    .Y(_09074_),
    .A2(_09073_),
    .A1(_09072_));
 sg13g2_a22oi_1 _17323_ (.Y(_09075_),
    .B1(net4859),
    .B2(\atari2600.ram[99][2] ),
    .A2(net4989),
    .A1(\atari2600.ram[96][2] ));
 sg13g2_a22oi_1 _17324_ (.Y(_09076_),
    .B1(net4813),
    .B2(\atari2600.ram[98][2] ),
    .A2(net4908),
    .A1(\atari2600.ram[97][2] ));
 sg13g2_a21oi_2 _17325_ (.B1(net4932),
    .Y(_09077_),
    .A2(_09076_),
    .A1(_09075_));
 sg13g2_a22oi_1 _17326_ (.Y(_09078_),
    .B1(net4859),
    .B2(\atari2600.ram[107][2] ),
    .A2(net4989),
    .A1(\atari2600.ram[104][2] ));
 sg13g2_a22oi_1 _17327_ (.Y(_09079_),
    .B1(net4813),
    .B2(\atari2600.ram[106][2] ),
    .A2(net4908),
    .A1(\atari2600.ram[105][2] ));
 sg13g2_a21oi_1 _17328_ (.A1(_09078_),
    .A2(_09079_),
    .Y(_09080_),
    .B1(net4946));
 sg13g2_nor4_2 _17329_ (.A(_09071_),
    .B(_09074_),
    .C(_09077_),
    .Y(_09081_),
    .D(_09080_));
 sg13g2_nor2_2 _17330_ (.A(net4771),
    .B(_09081_),
    .Y(_09082_));
 sg13g2_o21ai_1 _17331_ (.B1(net5022),
    .Y(_09083_),
    .A1(net4774),
    .A2(_09054_));
 sg13g2_nor4_2 _17332_ (.A(_09041_),
    .B(_09068_),
    .C(_09082_),
    .Y(_09084_),
    .D(_09083_));
 sg13g2_nor2_2 _17333_ (.A(_09027_),
    .B(_09084_),
    .Y(_00003_));
 sg13g2_a22oi_1 _17334_ (.Y(_09085_),
    .B1(net4840),
    .B2(\atari2600.ram[51][3] ),
    .A2(net4970),
    .A1(\atari2600.ram[48][3] ));
 sg13g2_a22oi_1 _17335_ (.Y(_09086_),
    .B1(net4795),
    .B2(\atari2600.ram[50][3] ),
    .A2(net4889),
    .A1(\atari2600.ram[49][3] ));
 sg13g2_a21oi_1 _17336_ (.A1(_09085_),
    .A2(_09086_),
    .Y(_09087_),
    .B1(net4926));
 sg13g2_a22oi_1 _17337_ (.Y(_09088_),
    .B1(net4838),
    .B2(\atari2600.ram[59][3] ),
    .A2(net4967),
    .A1(\atari2600.ram[56][3] ));
 sg13g2_a22oi_1 _17338_ (.Y(_09089_),
    .B1(net4792),
    .B2(\atari2600.ram[58][3] ),
    .A2(net4885),
    .A1(\atari2600.ram[57][3] ));
 sg13g2_a21oi_1 _17339_ (.A1(_09088_),
    .A2(_09089_),
    .Y(_09090_),
    .B1(net4940));
 sg13g2_a22oi_1 _17340_ (.Y(_09091_),
    .B1(net4837),
    .B2(\atari2600.ram[63][3] ),
    .A2(net4969),
    .A1(\atari2600.ram[60][3] ));
 sg13g2_a22oi_1 _17341_ (.Y(_09092_),
    .B1(net4793),
    .B2(\atari2600.ram[62][3] ),
    .A2(net4887),
    .A1(\atari2600.ram[61][3] ));
 sg13g2_a21oi_1 _17342_ (.A1(_09091_),
    .A2(_09092_),
    .Y(_09093_),
    .B1(net4951));
 sg13g2_a22oi_1 _17343_ (.Y(_09094_),
    .B1(net4983),
    .B2(\atari2600.ram[52][3] ),
    .A2(net4904),
    .A1(\atari2600.ram[53][3] ));
 sg13g2_a22oi_1 _17344_ (.Y(_09095_),
    .B1(net4808),
    .B2(\atari2600.ram[54][3] ),
    .A2(net4853),
    .A1(\atari2600.ram[55][3] ));
 sg13g2_a21oi_1 _17345_ (.A1(_09094_),
    .A2(_09095_),
    .Y(_09096_),
    .B1(net5011));
 sg13g2_nor2_1 _17346_ (.A(net5025),
    .B(_09093_),
    .Y(_09097_));
 sg13g2_nor3_1 _17347_ (.A(_09087_),
    .B(_09090_),
    .C(_09096_),
    .Y(_09098_));
 sg13g2_a22oi_1 _17348_ (.Y(_09099_),
    .B1(net4837),
    .B2(\atari2600.ram[43][3] ),
    .A2(net4967),
    .A1(\atari2600.ram[40][3] ));
 sg13g2_a22oi_1 _17349_ (.Y(_09100_),
    .B1(net4791),
    .B2(\atari2600.ram[42][3] ),
    .A2(net4885),
    .A1(\atari2600.ram[41][3] ));
 sg13g2_a21o_1 _17350_ (.A2(_09100_),
    .A1(_09099_),
    .B1(net4939),
    .X(_09101_));
 sg13g2_a22oi_1 _17351_ (.Y(_09102_),
    .B1(net4960),
    .B2(\atari2600.ram[36][3] ),
    .A2(net4880),
    .A1(\atari2600.ram[37][3] ));
 sg13g2_a22oi_1 _17352_ (.Y(_09103_),
    .B1(net4785),
    .B2(\atari2600.ram[38][3] ),
    .A2(net4830),
    .A1(\atari2600.ram[39][3] ));
 sg13g2_a21oi_1 _17353_ (.A1(_09102_),
    .A2(_09103_),
    .Y(_09104_),
    .B1(net5006));
 sg13g2_a22oi_1 _17354_ (.Y(_09105_),
    .B1(net4831),
    .B2(\atari2600.ram[47][3] ),
    .A2(net4961),
    .A1(\atari2600.ram[44][3] ));
 sg13g2_a22oi_1 _17355_ (.Y(_09106_),
    .B1(net4786),
    .B2(\atari2600.ram[46][3] ),
    .A2(net4882),
    .A1(\atari2600.ram[45][3] ));
 sg13g2_a21oi_1 _17356_ (.A1(_09105_),
    .A2(_09106_),
    .Y(_09107_),
    .B1(net4949));
 sg13g2_a22oi_1 _17357_ (.Y(_09108_),
    .B1(net4832),
    .B2(\atari2600.ram[35][3] ),
    .A2(net4962),
    .A1(\atari2600.ram[32][3] ));
 sg13g2_a22oi_1 _17358_ (.Y(_09109_),
    .B1(net4787),
    .B2(\atari2600.ram[34][3] ),
    .A2(net4881),
    .A1(\atari2600.ram[33][3] ));
 sg13g2_a21oi_2 _17359_ (.B1(net4925),
    .Y(_09110_),
    .A2(_09109_),
    .A1(_09108_));
 sg13g2_nor4_2 _17360_ (.A(net5027),
    .B(_09104_),
    .C(_09107_),
    .Y(_09111_),
    .D(_09110_));
 sg13g2_a221oi_1 _17361_ (.B2(_09111_),
    .C1(net4876),
    .B1(_09101_),
    .A1(_09097_),
    .Y(_09112_),
    .A2(_09098_));
 sg13g2_a22oi_1 _17362_ (.Y(_09113_),
    .B1(net4844),
    .B2(\atari2600.ram[3][3] ),
    .A2(net4974),
    .A1(\atari2600.ram[0][3] ));
 sg13g2_a22oi_1 _17363_ (.Y(_09114_),
    .B1(net4798),
    .B2(\atari2600.ram[2][3] ),
    .A2(net4894),
    .A1(\atari2600.ram[1][3] ));
 sg13g2_a21oi_1 _17364_ (.A1(_09113_),
    .A2(_09114_),
    .Y(_09115_),
    .B1(net4927));
 sg13g2_a22oi_1 _17365_ (.Y(_09116_),
    .B1(net4836),
    .B2(\atari2600.ram[11][3] ),
    .A2(net4966),
    .A1(\atari2600.ram[8][3] ));
 sg13g2_a22oi_1 _17366_ (.Y(_09117_),
    .B1(net4790),
    .B2(\atari2600.ram[10][3] ),
    .A2(net4884),
    .A1(\atari2600.ram[9][3] ));
 sg13g2_a21oi_2 _17367_ (.B1(net4938),
    .Y(_09118_),
    .A2(_09117_),
    .A1(_09116_));
 sg13g2_a22oi_1 _17368_ (.Y(_09119_),
    .B1(net4835),
    .B2(\atari2600.ram[15][3] ),
    .A2(net4965),
    .A1(\atari2600.ram[12][3] ));
 sg13g2_a22oi_1 _17369_ (.Y(_09120_),
    .B1(net4789),
    .B2(\atari2600.ram[14][3] ),
    .A2(net4883),
    .A1(\atari2600.ram[13][3] ));
 sg13g2_a21oi_2 _17370_ (.B1(net4950),
    .Y(_09121_),
    .A2(_09120_),
    .A1(_09119_));
 sg13g2_a22oi_1 _17371_ (.Y(_09122_),
    .B1(net4843),
    .B2(\atari2600.ram[7][3] ),
    .A2(net4973),
    .A1(\atari2600.ram[4][3] ));
 sg13g2_a22oi_1 _17372_ (.Y(_09123_),
    .B1(net4799),
    .B2(\atari2600.ram[6][3] ),
    .A2(net4893),
    .A1(\atari2600.ram[5][3] ));
 sg13g2_a21oi_1 _17373_ (.A1(_09122_),
    .A2(_09123_),
    .Y(_09124_),
    .B1(net5007));
 sg13g2_nor4_2 _17374_ (.A(_09115_),
    .B(_09118_),
    .C(_09121_),
    .Y(_09125_),
    .D(_09124_));
 sg13g2_nor2_1 _17375_ (.A(net4777),
    .B(_09125_),
    .Y(_09126_));
 sg13g2_a22oi_1 _17376_ (.Y(_09127_),
    .B1(net4846),
    .B2(\atari2600.ram[27][3] ),
    .A2(net4976),
    .A1(\atari2600.ram[24][3] ));
 sg13g2_a22oi_1 _17377_ (.Y(_09128_),
    .B1(net4806),
    .B2(\atari2600.ram[26][3] ),
    .A2(net4900),
    .A1(\atari2600.ram[25][3] ));
 sg13g2_a21oi_2 _17378_ (.B1(net4941),
    .Y(_09129_),
    .A2(_09128_),
    .A1(_09127_));
 sg13g2_a22oi_1 _17379_ (.Y(_09130_),
    .B1(net4848),
    .B2(\atari2600.ram[19][3] ),
    .A2(net4979),
    .A1(\atari2600.ram[16][3] ));
 sg13g2_a22oi_1 _17380_ (.Y(_09131_),
    .B1(net4802),
    .B2(\atari2600.ram[18][3] ),
    .A2(net4897),
    .A1(\atari2600.ram[17][3] ));
 sg13g2_a21oi_1 _17381_ (.A1(_09130_),
    .A2(_09131_),
    .Y(_09132_),
    .B1(net4928));
 sg13g2_a22oi_1 _17382_ (.Y(_09133_),
    .B1(net4848),
    .B2(\atari2600.ram[23][3] ),
    .A2(net4979),
    .A1(\atari2600.ram[20][3] ));
 sg13g2_a22oi_1 _17383_ (.Y(_09134_),
    .B1(net4802),
    .B2(\atari2600.ram[22][3] ),
    .A2(net4897),
    .A1(\atari2600.ram[21][3] ));
 sg13g2_a21oi_1 _17384_ (.A1(_09133_),
    .A2(_09134_),
    .Y(_09135_),
    .B1(net5008));
 sg13g2_a22oi_1 _17385_ (.Y(_09136_),
    .B1(net4848),
    .B2(\atari2600.ram[31][3] ),
    .A2(net4979),
    .A1(\atari2600.ram[28][3] ));
 sg13g2_a22oi_1 _17386_ (.Y(_09137_),
    .B1(net4803),
    .B2(\atari2600.ram[30][3] ),
    .A2(net4898),
    .A1(\atari2600.ram[29][3] ));
 sg13g2_a21oi_1 _17387_ (.A1(_09136_),
    .A2(_09137_),
    .Y(_09138_),
    .B1(net4952));
 sg13g2_nor4_2 _17388_ (.A(_09129_),
    .B(_09132_),
    .C(_09135_),
    .Y(_09139_),
    .D(_09138_));
 sg13g2_o21ai_1 _17389_ (.B1(net5023),
    .Y(_09140_),
    .A1(net4773),
    .A2(_09139_));
 sg13g2_nor3_1 _17390_ (.A(_09112_),
    .B(_09126_),
    .C(_09140_),
    .Y(_09141_));
 sg13g2_a22oi_1 _17391_ (.Y(_09142_),
    .B1(net4847),
    .B2(\atari2600.ram[87][3] ),
    .A2(net4977),
    .A1(\atari2600.ram[84][3] ));
 sg13g2_a22oi_1 _17392_ (.Y(_09143_),
    .B1(net4803),
    .B2(\atari2600.ram[86][3] ),
    .A2(net4898),
    .A1(\atari2600.ram[85][3] ));
 sg13g2_a21oi_2 _17393_ (.B1(net5008),
    .Y(_09144_),
    .A2(_09143_),
    .A1(_09142_));
 sg13g2_a22oi_1 _17394_ (.Y(_09145_),
    .B1(net4850),
    .B2(\atari2600.ram[91][3] ),
    .A2(net4980),
    .A1(\atari2600.ram[88][3] ));
 sg13g2_a22oi_1 _17395_ (.Y(_09146_),
    .B1(net4821),
    .B2(\atari2600.ram[90][3] ),
    .A2(net4916),
    .A1(\atari2600.ram[89][3] ));
 sg13g2_a21oi_2 _17396_ (.B1(net4942),
    .Y(_09147_),
    .A2(_09146_),
    .A1(_09145_));
 sg13g2_a22oi_1 _17397_ (.Y(_09148_),
    .B1(net4868),
    .B2(\atari2600.ram[95][3] ),
    .A2(net4997),
    .A1(\atari2600.ram[92][3] ));
 sg13g2_a22oi_1 _17398_ (.Y(_09149_),
    .B1(net4823),
    .B2(\atari2600.ram[94][3] ),
    .A2(net4918),
    .A1(\atari2600.ram[93][3] ));
 sg13g2_a21oi_1 _17399_ (.A1(_09148_),
    .A2(_09149_),
    .Y(_09150_),
    .B1(net4957));
 sg13g2_a22oi_1 _17400_ (.Y(_09151_),
    .B1(net4866),
    .B2(\atari2600.ram[83][3] ),
    .A2(net4996),
    .A1(\atari2600.ram[80][3] ));
 sg13g2_a22oi_1 _17401_ (.Y(_09152_),
    .B1(net4823),
    .B2(\atari2600.ram[82][3] ),
    .A2(net4918),
    .A1(\atari2600.ram[81][3] ));
 sg13g2_a21oi_1 _17402_ (.A1(_09151_),
    .A2(_09152_),
    .Y(_09153_),
    .B1(net4933));
 sg13g2_nor4_2 _17403_ (.A(_09144_),
    .B(_09147_),
    .C(_09150_),
    .Y(_09154_),
    .D(_09153_));
 sg13g2_nor2_1 _17404_ (.A(net4774),
    .B(_09154_),
    .Y(_09155_));
 sg13g2_a22oi_1 _17405_ (.Y(_09156_),
    .B1(net4865),
    .B2(\atari2600.ram[71][3] ),
    .A2(net4996),
    .A1(\atari2600.ram[68][3] ));
 sg13g2_a22oi_1 _17406_ (.Y(_09157_),
    .B1(net4819),
    .B2(\atari2600.ram[70][3] ),
    .A2(net4914),
    .A1(\atari2600.ram[69][3] ));
 sg13g2_a21oi_2 _17407_ (.B1(net5016),
    .Y(_09158_),
    .A2(_09157_),
    .A1(_09156_));
 sg13g2_a22oi_1 _17408_ (.Y(_09159_),
    .B1(net4865),
    .B2(\atari2600.ram[67][3] ),
    .A2(net4996),
    .A1(\atari2600.ram[64][3] ));
 sg13g2_a22oi_1 _17409_ (.Y(_09160_),
    .B1(net4818),
    .B2(\atari2600.ram[66][3] ),
    .A2(net4913),
    .A1(\atari2600.ram[65][3] ));
 sg13g2_a21oi_1 _17410_ (.A1(_09159_),
    .A2(_09160_),
    .Y(_09161_),
    .B1(net4933));
 sg13g2_a22oi_1 _17411_ (.Y(_09162_),
    .B1(net4872),
    .B2(\atari2600.ram[79][3] ),
    .A2(net4998),
    .A1(\atari2600.ram[76][3] ));
 sg13g2_a22oi_1 _17412_ (.Y(_09163_),
    .B1(net4822),
    .B2(\atari2600.ram[78][3] ),
    .A2(net4917),
    .A1(\atari2600.ram[77][3] ));
 sg13g2_a21oi_2 _17413_ (.B1(net4958),
    .Y(_09164_),
    .A2(_09163_),
    .A1(_09162_));
 sg13g2_a22oi_1 _17414_ (.Y(_09165_),
    .B1(net4868),
    .B2(\atari2600.ram[75][3] ),
    .A2(net4998),
    .A1(\atari2600.ram[72][3] ));
 sg13g2_a22oi_1 _17415_ (.Y(_09166_),
    .B1(net4823),
    .B2(\atari2600.ram[74][3] ),
    .A2(net4918),
    .A1(\atari2600.ram[73][3] ));
 sg13g2_a21oi_1 _17416_ (.A1(_09165_),
    .A2(_09166_),
    .Y(_09167_),
    .B1(net4945));
 sg13g2_nor4_2 _17417_ (.A(_09158_),
    .B(_09161_),
    .C(_09164_),
    .Y(_09168_),
    .D(_09167_));
 sg13g2_a22oi_1 _17418_ (.Y(_09169_),
    .B1(net4842),
    .B2(\atari2600.ram[119][3] ),
    .A2(net4972),
    .A1(\atari2600.ram[116][3] ));
 sg13g2_a22oi_1 _17419_ (.Y(_09170_),
    .B1(net4794),
    .B2(\atari2600.ram[118][3] ),
    .A2(net4888),
    .A1(\atari2600.ram[117][3] ));
 sg13g2_a21oi_1 _17420_ (.A1(_09169_),
    .A2(_09170_),
    .Y(_09171_),
    .B1(net5009));
 sg13g2_a22oi_1 _17421_ (.Y(_09172_),
    .B1(net4863),
    .B2(\atari2600.ram[127][3] ),
    .A2(net4994),
    .A1(\atari2600.ram[124][3] ));
 sg13g2_a22oi_1 _17422_ (.Y(_09173_),
    .B1(net4818),
    .B2(\atari2600.ram[126][3] ),
    .A2(net4913),
    .A1(\atari2600.ram[125][3] ));
 sg13g2_a21oi_1 _17423_ (.A1(_09172_),
    .A2(_09173_),
    .Y(_09174_),
    .B1(net4958));
 sg13g2_a22oi_1 _17424_ (.Y(_09175_),
    .B1(net4853),
    .B2(\atari2600.ram[115][3] ),
    .A2(net4983),
    .A1(\atari2600.ram[112][3] ));
 sg13g2_a22oi_1 _17425_ (.Y(_09176_),
    .B1(net4808),
    .B2(\atari2600.ram[114][3] ),
    .A2(net4902),
    .A1(\atari2600.ram[113][3] ));
 sg13g2_a21oi_2 _17426_ (.B1(net4930),
    .Y(_09177_),
    .A2(_09176_),
    .A1(_09175_));
 sg13g2_a22oi_1 _17427_ (.Y(_09178_),
    .B1(net4863),
    .B2(\atari2600.ram[123][3] ),
    .A2(net4994),
    .A1(\atari2600.ram[120][3] ));
 sg13g2_a22oi_1 _17428_ (.Y(_09179_),
    .B1(net4811),
    .B2(\atari2600.ram[122][3] ),
    .A2(net4906),
    .A1(\atari2600.ram[121][3] ));
 sg13g2_a21oi_1 _17429_ (.A1(_09178_),
    .A2(_09179_),
    .Y(_09180_),
    .B1(net4943));
 sg13g2_nor4_1 _17430_ (.A(_09171_),
    .B(_09174_),
    .C(_09177_),
    .D(_09180_),
    .Y(_09181_));
 sg13g2_nor2_1 _17431_ (.A(_08729_),
    .B(_09181_),
    .Y(_09182_));
 sg13g2_a22oi_1 _17432_ (.Y(_09183_),
    .B1(net4859),
    .B2(\atari2600.ram[107][3] ),
    .A2(net4989),
    .A1(\atari2600.ram[104][3] ));
 sg13g2_a22oi_1 _17433_ (.Y(_09184_),
    .B1(net4814),
    .B2(\atari2600.ram[106][3] ),
    .A2(net4910),
    .A1(\atari2600.ram[105][3] ));
 sg13g2_a21oi_1 _17434_ (.A1(_09183_),
    .A2(_09184_),
    .Y(_09185_),
    .B1(net4946));
 sg13g2_a22oi_1 _17435_ (.Y(_09186_),
    .B1(net4859),
    .B2(\atari2600.ram[99][3] ),
    .A2(net4989),
    .A1(\atari2600.ram[96][3] ));
 sg13g2_a22oi_1 _17436_ (.Y(_09187_),
    .B1(net4813),
    .B2(\atari2600.ram[98][3] ),
    .A2(net4908),
    .A1(\atari2600.ram[97][3] ));
 sg13g2_a21oi_2 _17437_ (.B1(net4932),
    .Y(_09188_),
    .A2(_09187_),
    .A1(_09186_));
 sg13g2_a22oi_1 _17438_ (.Y(_09189_),
    .B1(net4861),
    .B2(\atari2600.ram[103][3] ),
    .A2(net4991),
    .A1(\atari2600.ram[100][3] ));
 sg13g2_a22oi_1 _17439_ (.Y(_09190_),
    .B1(net4816),
    .B2(\atari2600.ram[102][3] ),
    .A2(net4910),
    .A1(\atari2600.ram[101][3] ));
 sg13g2_a21oi_1 _17440_ (.A1(_09189_),
    .A2(_09190_),
    .Y(_09191_),
    .B1(net5014));
 sg13g2_a22oi_1 _17441_ (.Y(_09192_),
    .B1(net4861),
    .B2(\atari2600.ram[111][3] ),
    .A2(net4991),
    .A1(\atari2600.ram[108][3] ));
 sg13g2_a22oi_1 _17442_ (.Y(_09193_),
    .B1(net4816),
    .B2(\atari2600.ram[110][3] ),
    .A2(net4910),
    .A1(\atari2600.ram[109][3] ));
 sg13g2_a21oi_1 _17443_ (.A1(_09192_),
    .A2(_09193_),
    .Y(_09194_),
    .B1(net4954));
 sg13g2_nor4_2 _17444_ (.A(_09185_),
    .B(_09188_),
    .C(_09191_),
    .Y(_09195_),
    .D(_09194_));
 sg13g2_nor2_2 _17445_ (.A(net4771),
    .B(_09195_),
    .Y(_09196_));
 sg13g2_o21ai_1 _17446_ (.B1(net5020),
    .Y(_09197_),
    .A1(net4778),
    .A2(_09168_));
 sg13g2_nor4_2 _17447_ (.A(_09155_),
    .B(_09182_),
    .C(_09196_),
    .Y(_09198_),
    .D(_09197_));
 sg13g2_nor2_2 _17448_ (.A(_09141_),
    .B(_09198_),
    .Y(_00004_));
 sg13g2_a22oi_1 _17449_ (.Y(_09199_),
    .B1(net4967),
    .B2(\atari2600.ram[56][4] ),
    .A2(net4885),
    .A1(\atari2600.ram[57][4] ));
 sg13g2_a22oi_1 _17450_ (.Y(_09200_),
    .B1(net4791),
    .B2(\atari2600.ram[58][4] ),
    .A2(net4837),
    .A1(\atari2600.ram[59][4] ));
 sg13g2_a21oi_1 _17451_ (.A1(_09199_),
    .A2(_09200_),
    .Y(_09201_),
    .B1(net4937));
 sg13g2_a22oi_1 _17452_ (.Y(_09202_),
    .B1(net4840),
    .B2(\atari2600.ram[51][4] ),
    .A2(net4970),
    .A1(\atari2600.ram[48][4] ));
 sg13g2_a22oi_1 _17453_ (.Y(_09203_),
    .B1(net4795),
    .B2(\atari2600.ram[50][4] ),
    .A2(net4889),
    .A1(\atari2600.ram[49][4] ));
 sg13g2_a21oi_1 _17454_ (.A1(_09202_),
    .A2(_09203_),
    .Y(_09204_),
    .B1(net4926));
 sg13g2_a22oi_1 _17455_ (.Y(_09205_),
    .B1(net4855),
    .B2(\atari2600.ram[55][4] ),
    .A2(net4968),
    .A1(\atari2600.ram[52][4] ));
 sg13g2_a22oi_1 _17456_ (.Y(_09206_),
    .B1(net4808),
    .B2(\atari2600.ram[54][4] ),
    .A2(net4902),
    .A1(\atari2600.ram[53][4] ));
 sg13g2_a21oi_2 _17457_ (.B1(net5012),
    .Y(_09207_),
    .A2(_09206_),
    .A1(_09205_));
 sg13g2_a22oi_1 _17458_ (.Y(_09208_),
    .B1(net4838),
    .B2(\atari2600.ram[63][4] ),
    .A2(net4969),
    .A1(\atari2600.ram[60][4] ));
 sg13g2_a22oi_1 _17459_ (.Y(_09209_),
    .B1(net4793),
    .B2(\atari2600.ram[62][4] ),
    .A2(net4887),
    .A1(\atari2600.ram[61][4] ));
 sg13g2_a21oi_1 _17460_ (.A1(_09208_),
    .A2(_09209_),
    .Y(_09210_),
    .B1(net4951));
 sg13g2_nor2_1 _17461_ (.A(net5025),
    .B(_09207_),
    .Y(_09211_));
 sg13g2_nor3_1 _17462_ (.A(_09201_),
    .B(_09204_),
    .C(_09210_),
    .Y(_09212_));
 sg13g2_a22oi_1 _17463_ (.Y(_09213_),
    .B1(net4831),
    .B2(\atari2600.ram[47][4] ),
    .A2(net4961),
    .A1(\atari2600.ram[44][4] ));
 sg13g2_a22oi_1 _17464_ (.Y(_09214_),
    .B1(net4785),
    .B2(\atari2600.ram[46][4] ),
    .A2(net4880),
    .A1(\atari2600.ram[45][4] ));
 sg13g2_a21oi_1 _17465_ (.A1(_09213_),
    .A2(_09214_),
    .Y(_09215_),
    .B1(net4949));
 sg13g2_a22oi_1 _17466_ (.Y(_09216_),
    .B1(net4837),
    .B2(\atari2600.ram[35][4] ),
    .A2(net4967),
    .A1(\atari2600.ram[32][4] ));
 sg13g2_a22oi_1 _17467_ (.Y(_09217_),
    .B1(net4791),
    .B2(\atari2600.ram[34][4] ),
    .A2(net4885),
    .A1(\atari2600.ram[33][4] ));
 sg13g2_a21o_1 _17468_ (.A2(_09217_),
    .A1(_09216_),
    .B1(net4925),
    .X(_09218_));
 sg13g2_a22oi_1 _17469_ (.Y(_09219_),
    .B1(net4833),
    .B2(\atari2600.ram[43][4] ),
    .A2(net4963),
    .A1(\atari2600.ram[40][4] ));
 sg13g2_a22oi_1 _17470_ (.Y(_09220_),
    .B1(net4787),
    .B2(\atari2600.ram[42][4] ),
    .A2(net4881),
    .A1(\atari2600.ram[41][4] ));
 sg13g2_a21oi_1 _17471_ (.A1(_09219_),
    .A2(_09220_),
    .Y(_09221_),
    .B1(net4937));
 sg13g2_a22oi_1 _17472_ (.Y(_09222_),
    .B1(net4960),
    .B2(\atari2600.ram[36][4] ),
    .A2(net4880),
    .A1(\atari2600.ram[37][4] ));
 sg13g2_a22oi_1 _17473_ (.Y(_09223_),
    .B1(net4785),
    .B2(\atari2600.ram[38][4] ),
    .A2(net4830),
    .A1(\atari2600.ram[39][4] ));
 sg13g2_a21oi_1 _17474_ (.A1(_09222_),
    .A2(_09223_),
    .Y(_09224_),
    .B1(net5006));
 sg13g2_nor4_2 _17475_ (.A(net5027),
    .B(_09215_),
    .C(_09221_),
    .Y(_09225_),
    .D(_09224_));
 sg13g2_a221oi_1 _17476_ (.B2(_09225_),
    .C1(net4876),
    .B1(_09218_),
    .A1(_09211_),
    .Y(_09226_),
    .A2(_09212_));
 sg13g2_a22oi_1 _17477_ (.Y(_09227_),
    .B1(net4848),
    .B2(\atari2600.ram[31][4] ),
    .A2(net4979),
    .A1(\atari2600.ram[28][4] ));
 sg13g2_a22oi_1 _17478_ (.Y(_09228_),
    .B1(net4803),
    .B2(\atari2600.ram[30][4] ),
    .A2(net4898),
    .A1(\atari2600.ram[29][4] ));
 sg13g2_a21oi_1 _17479_ (.A1(_09227_),
    .A2(_09228_),
    .Y(_09229_),
    .B1(net4952));
 sg13g2_a22oi_1 _17480_ (.Y(_09230_),
    .B1(net4846),
    .B2(\atari2600.ram[27][4] ),
    .A2(net4976),
    .A1(\atari2600.ram[24][4] ));
 sg13g2_a22oi_1 _17481_ (.Y(_09231_),
    .B1(net4801),
    .B2(\atari2600.ram[26][4] ),
    .A2(net4896),
    .A1(\atari2600.ram[25][4] ));
 sg13g2_a21oi_2 _17482_ (.B1(net4941),
    .Y(_09232_),
    .A2(_09231_),
    .A1(_09230_));
 sg13g2_a22oi_1 _17483_ (.Y(_09233_),
    .B1(net4848),
    .B2(\atari2600.ram[19][4] ),
    .A2(net4979),
    .A1(\atari2600.ram[16][4] ));
 sg13g2_a22oi_1 _17484_ (.Y(_09234_),
    .B1(net4802),
    .B2(\atari2600.ram[18][4] ),
    .A2(net4897),
    .A1(\atari2600.ram[17][4] ));
 sg13g2_a21oi_2 _17485_ (.B1(net4928),
    .Y(_09235_),
    .A2(_09234_),
    .A1(_09233_));
 sg13g2_a22oi_1 _17486_ (.Y(_09236_),
    .B1(net4848),
    .B2(\atari2600.ram[23][4] ),
    .A2(net4979),
    .A1(\atari2600.ram[20][4] ));
 sg13g2_a22oi_1 _17487_ (.Y(_09237_),
    .B1(net4802),
    .B2(\atari2600.ram[22][4] ),
    .A2(net4897),
    .A1(\atari2600.ram[21][4] ));
 sg13g2_a21oi_1 _17488_ (.A1(_09236_),
    .A2(_09237_),
    .Y(_09238_),
    .B1(net5008));
 sg13g2_nor4_2 _17489_ (.A(_09229_),
    .B(_09232_),
    .C(_09235_),
    .Y(_09239_),
    .D(_09238_));
 sg13g2_a22oi_1 _17490_ (.Y(_09240_),
    .B1(net4844),
    .B2(\atari2600.ram[3][4] ),
    .A2(net4974),
    .A1(\atari2600.ram[0][4] ));
 sg13g2_a22oi_1 _17491_ (.Y(_09241_),
    .B1(net4807),
    .B2(\atari2600.ram[2][4] ),
    .A2(net4901),
    .A1(\atari2600.ram[1][4] ));
 sg13g2_a21oi_1 _17492_ (.A1(_09240_),
    .A2(_09241_),
    .Y(_09242_),
    .B1(net4927));
 sg13g2_a22oi_1 _17493_ (.Y(_09243_),
    .B1(net4834),
    .B2(\atari2600.ram[11][4] ),
    .A2(net4964),
    .A1(\atari2600.ram[8][4] ));
 sg13g2_a22oi_1 _17494_ (.Y(_09244_),
    .B1(net4798),
    .B2(\atari2600.ram[10][4] ),
    .A2(net4892),
    .A1(\atari2600.ram[9][4] ));
 sg13g2_a21oi_1 _17495_ (.A1(_09243_),
    .A2(_09244_),
    .Y(_09245_),
    .B1(net4941));
 sg13g2_a22oi_1 _17496_ (.Y(_09246_),
    .B1(net4834),
    .B2(\atari2600.ram[15][4] ),
    .A2(net4966),
    .A1(\atari2600.ram[12][4] ));
 sg13g2_a22oi_1 _17497_ (.Y(_09247_),
    .B1(net4798),
    .B2(\atari2600.ram[14][4] ),
    .A2(net4892),
    .A1(\atari2600.ram[13][4] ));
 sg13g2_a21oi_1 _17498_ (.A1(_09246_),
    .A2(_09247_),
    .Y(_09248_),
    .B1(net4950));
 sg13g2_a22oi_1 _17499_ (.Y(_09249_),
    .B1(net4843),
    .B2(\atari2600.ram[7][4] ),
    .A2(net4973),
    .A1(\atari2600.ram[4][4] ));
 sg13g2_a22oi_1 _17500_ (.Y(_09250_),
    .B1(net4799),
    .B2(\atari2600.ram[6][4] ),
    .A2(net4893),
    .A1(\atari2600.ram[5][4] ));
 sg13g2_a21oi_1 _17501_ (.A1(_09249_),
    .A2(_09250_),
    .Y(_09251_),
    .B1(net5007));
 sg13g2_nor4_1 _17502_ (.A(_09242_),
    .B(_09245_),
    .C(_09248_),
    .D(_09251_),
    .Y(_09252_));
 sg13g2_nor2_1 _17503_ (.A(net4777),
    .B(_09252_),
    .Y(_09253_));
 sg13g2_o21ai_1 _17504_ (.B1(net5023),
    .Y(_09254_),
    .A1(net4773),
    .A2(_09239_));
 sg13g2_nor3_1 _17505_ (.A(_09226_),
    .B(_09253_),
    .C(_09254_),
    .Y(_09255_));
 sg13g2_a22oi_1 _17506_ (.Y(_09256_),
    .B1(net4863),
    .B2(\atari2600.ram[127][4] ),
    .A2(net4994),
    .A1(\atari2600.ram[124][4] ));
 sg13g2_a22oi_1 _17507_ (.Y(_09257_),
    .B1(net4819),
    .B2(\atari2600.ram[126][4] ),
    .A2(net4914),
    .A1(\atari2600.ram[125][4] ));
 sg13g2_a21oi_1 _17508_ (.A1(_09256_),
    .A2(_09257_),
    .Y(_09258_),
    .B1(net4958));
 sg13g2_a22oi_1 _17509_ (.Y(_09259_),
    .B1(net4857),
    .B2(\atari2600.ram[119][4] ),
    .A2(net4987),
    .A1(\atari2600.ram[116][4] ));
 sg13g2_a22oi_1 _17510_ (.Y(_09260_),
    .B1(net4812),
    .B2(\atari2600.ram[118][4] ),
    .A2(net4907),
    .A1(\atari2600.ram[117][4] ));
 sg13g2_a21oi_1 _17511_ (.A1(_09259_),
    .A2(_09260_),
    .Y(_09261_),
    .B1(net5016));
 sg13g2_a22oi_1 _17512_ (.Y(_09262_),
    .B1(net4854),
    .B2(\atari2600.ram[115][4] ),
    .A2(net4984),
    .A1(\atari2600.ram[112][4] ));
 sg13g2_a22oi_1 _17513_ (.Y(_09263_),
    .B1(net4809),
    .B2(\atari2600.ram[114][4] ),
    .A2(net4903),
    .A1(\atari2600.ram[113][4] ));
 sg13g2_a21oi_2 _17514_ (.B1(net4930),
    .Y(_09264_),
    .A2(_09263_),
    .A1(_09262_));
 sg13g2_a22oi_1 _17515_ (.Y(_09265_),
    .B1(net4856),
    .B2(\atari2600.ram[123][4] ),
    .A2(net4987),
    .A1(\atari2600.ram[120][4] ));
 sg13g2_a22oi_1 _17516_ (.Y(_09266_),
    .B1(net4811),
    .B2(\atari2600.ram[122][4] ),
    .A2(net4905),
    .A1(\atari2600.ram[121][4] ));
 sg13g2_a21oi_1 _17517_ (.A1(_09265_),
    .A2(_09266_),
    .Y(_09267_),
    .B1(net4943));
 sg13g2_nor4_1 _17518_ (.A(_09258_),
    .B(_09261_),
    .C(_09264_),
    .D(_09267_),
    .Y(_09268_));
 sg13g2_o21ai_1 _17519_ (.B1(net5020),
    .Y(_09269_),
    .A1(net4776),
    .A2(_09268_));
 sg13g2_a22oi_1 _17520_ (.Y(_09270_),
    .B1(net4871),
    .B2(\atari2600.ram[75][4] ),
    .A2(net5002),
    .A1(\atari2600.ram[72][4] ));
 sg13g2_a22oi_1 _17521_ (.Y(_09271_),
    .B1(net4827),
    .B2(\atari2600.ram[74][4] ),
    .A2(net4922),
    .A1(\atari2600.ram[73][4] ));
 sg13g2_a21oi_2 _17522_ (.B1(net4945),
    .Y(_09272_),
    .A2(_09271_),
    .A1(_09270_));
 sg13g2_a22oi_1 _17523_ (.Y(_09273_),
    .B1(net4869),
    .B2(\atari2600.ram[71][4] ),
    .A2(net5000),
    .A1(\atari2600.ram[68][4] ));
 sg13g2_a22oi_1 _17524_ (.Y(_09274_),
    .B1(net4825),
    .B2(\atari2600.ram[70][4] ),
    .A2(net4920),
    .A1(\atari2600.ram[69][4] ));
 sg13g2_a21oi_1 _17525_ (.A1(_09273_),
    .A2(_09274_),
    .Y(_09275_),
    .B1(net5015));
 sg13g2_a22oi_1 _17526_ (.Y(_09276_),
    .B1(net4871),
    .B2(\atari2600.ram[79][4] ),
    .A2(net5003),
    .A1(\atari2600.ram[76][4] ));
 sg13g2_a22oi_1 _17527_ (.Y(_09277_),
    .B1(net4827),
    .B2(\atari2600.ram[78][4] ),
    .A2(net4922),
    .A1(\atari2600.ram[77][4] ));
 sg13g2_a21oi_2 _17528_ (.B1(net4959),
    .Y(_09278_),
    .A2(_09277_),
    .A1(_09276_));
 sg13g2_a22oi_1 _17529_ (.Y(_09279_),
    .B1(net4869),
    .B2(\atari2600.ram[67][4] ),
    .A2(net5000),
    .A1(\atari2600.ram[64][4] ));
 sg13g2_a22oi_1 _17530_ (.Y(_09280_),
    .B1(net4825),
    .B2(\atari2600.ram[66][4] ),
    .A2(net4920),
    .A1(\atari2600.ram[65][4] ));
 sg13g2_a21oi_1 _17531_ (.A1(_09279_),
    .A2(_09280_),
    .Y(_09281_),
    .B1(net4935));
 sg13g2_nor4_2 _17532_ (.A(_09272_),
    .B(_09275_),
    .C(_09278_),
    .Y(_09282_),
    .D(_09281_));
 sg13g2_nor2_1 _17533_ (.A(net4778),
    .B(_09282_),
    .Y(_09283_));
 sg13g2_a22oi_1 _17534_ (.Y(_09284_),
    .B1(net4863),
    .B2(\atari2600.ram[87][4] ),
    .A2(net4994),
    .A1(\atari2600.ram[84][4] ));
 sg13g2_a22oi_1 _17535_ (.Y(_09285_),
    .B1(net4820),
    .B2(\atari2600.ram[86][4] ),
    .A2(net4915),
    .A1(\atari2600.ram[85][4] ));
 sg13g2_a21oi_1 _17536_ (.A1(_09284_),
    .A2(_09285_),
    .Y(_09286_),
    .B1(net5016));
 sg13g2_a22oi_1 _17537_ (.Y(_09287_),
    .B1(net4865),
    .B2(\atari2600.ram[83][4] ),
    .A2(net4996),
    .A1(\atari2600.ram[80][4] ));
 sg13g2_a22oi_1 _17538_ (.Y(_09288_),
    .B1(net4823),
    .B2(\atari2600.ram[82][4] ),
    .A2(net4918),
    .A1(\atari2600.ram[81][4] ));
 sg13g2_a21oi_1 _17539_ (.A1(_09287_),
    .A2(_09288_),
    .Y(_09289_),
    .B1(net4933));
 sg13g2_a22oi_1 _17540_ (.Y(_09290_),
    .B1(net4867),
    .B2(\atari2600.ram[91][4] ),
    .A2(net4998),
    .A1(\atari2600.ram[88][4] ));
 sg13g2_a22oi_1 _17541_ (.Y(_09291_),
    .B1(net4821),
    .B2(\atari2600.ram[90][4] ),
    .A2(net4916),
    .A1(\atari2600.ram[89][4] ));
 sg13g2_a21oi_2 _17542_ (.B1(net4942),
    .Y(_09292_),
    .A2(_09291_),
    .A1(_09290_));
 sg13g2_a22oi_1 _17543_ (.Y(_09293_),
    .B1(net4868),
    .B2(\atari2600.ram[95][4] ),
    .A2(net4998),
    .A1(\atari2600.ram[92][4] ));
 sg13g2_a22oi_1 _17544_ (.Y(_09294_),
    .B1(net4822),
    .B2(\atari2600.ram[94][4] ),
    .A2(net4917),
    .A1(\atari2600.ram[93][4] ));
 sg13g2_a21oi_2 _17545_ (.B1(net4958),
    .Y(_09295_),
    .A2(_09294_),
    .A1(_09293_));
 sg13g2_nor4_1 _17546_ (.A(_09286_),
    .B(_09289_),
    .C(_09292_),
    .D(_09295_),
    .Y(_09296_));
 sg13g2_nor2_1 _17547_ (.A(net4775),
    .B(_09296_),
    .Y(_09297_));
 sg13g2_a22oi_1 _17548_ (.Y(_09298_),
    .B1(net4860),
    .B2(\atari2600.ram[107][4] ),
    .A2(net4990),
    .A1(\atari2600.ram[104][4] ));
 sg13g2_a22oi_1 _17549_ (.Y(_09299_),
    .B1(net4815),
    .B2(\atari2600.ram[106][4] ),
    .A2(net4909),
    .A1(\atari2600.ram[105][4] ));
 sg13g2_a21oi_1 _17550_ (.A1(_09298_),
    .A2(_09299_),
    .Y(_09300_),
    .B1(net4944));
 sg13g2_a22oi_1 _17551_ (.Y(_09301_),
    .B1(net4862),
    .B2(\atari2600.ram[111][4] ),
    .A2(net4991),
    .A1(\atari2600.ram[108][4] ));
 sg13g2_a22oi_1 _17552_ (.Y(_09302_),
    .B1(net4816),
    .B2(\atari2600.ram[110][4] ),
    .A2(net4910),
    .A1(\atari2600.ram[109][4] ));
 sg13g2_a21oi_2 _17553_ (.B1(net4954),
    .Y(_09303_),
    .A2(_09302_),
    .A1(_09301_));
 sg13g2_a22oi_1 _17554_ (.Y(_09304_),
    .B1(net4860),
    .B2(\atari2600.ram[99][4] ),
    .A2(net4990),
    .A1(\atari2600.ram[96][4] ));
 sg13g2_a22oi_1 _17555_ (.Y(_09305_),
    .B1(net4815),
    .B2(\atari2600.ram[98][4] ),
    .A2(net4909),
    .A1(\atari2600.ram[97][4] ));
 sg13g2_a21oi_1 _17556_ (.A1(_09304_),
    .A2(_09305_),
    .Y(_09306_),
    .B1(net4932));
 sg13g2_a22oi_1 _17557_ (.Y(_09307_),
    .B1(net4861),
    .B2(\atari2600.ram[103][4] ),
    .A2(net4991),
    .A1(\atari2600.ram[100][4] ));
 sg13g2_a22oi_1 _17558_ (.Y(_09308_),
    .B1(net4814),
    .B2(\atari2600.ram[102][4] ),
    .A2(net4910),
    .A1(\atari2600.ram[101][4] ));
 sg13g2_a21oi_1 _17559_ (.A1(_09307_),
    .A2(_09308_),
    .Y(_09309_),
    .B1(net5014));
 sg13g2_nor4_2 _17560_ (.A(_09300_),
    .B(_09303_),
    .C(_09306_),
    .Y(_09310_),
    .D(_09309_));
 sg13g2_nor2_1 _17561_ (.A(_08783_),
    .B(_09310_),
    .Y(_09311_));
 sg13g2_nor4_2 _17562_ (.A(_09269_),
    .B(_09283_),
    .C(_09297_),
    .Y(_09312_),
    .D(_09311_));
 sg13g2_nor2_2 _17563_ (.A(_09255_),
    .B(_09312_),
    .Y(_00005_));
 sg13g2_a22oi_1 _17564_ (.Y(_09313_),
    .B1(net4856),
    .B2(\atari2600.ram[123][5] ),
    .A2(net4988),
    .A1(\atari2600.ram[120][5] ));
 sg13g2_a22oi_1 _17565_ (.Y(_09314_),
    .B1(net4811),
    .B2(\atari2600.ram[122][5] ),
    .A2(net4905),
    .A1(\atari2600.ram[121][5] ));
 sg13g2_a21oi_1 _17566_ (.A1(_09313_),
    .A2(_09314_),
    .Y(_09315_),
    .B1(net4943));
 sg13g2_a22oi_1 _17567_ (.Y(_09316_),
    .B1(net4986),
    .B2(\atari2600.ram[116][5] ),
    .A2(net4907),
    .A1(\atari2600.ram[117][5] ));
 sg13g2_a22oi_1 _17568_ (.Y(_09317_),
    .B1(net4812),
    .B2(\atari2600.ram[118][5] ),
    .A2(net4857),
    .A1(\atari2600.ram[119][5] ));
 sg13g2_a21oi_1 _17569_ (.A1(_09316_),
    .A2(_09317_),
    .Y(_09318_),
    .B1(net5013));
 sg13g2_a22oi_1 _17570_ (.Y(_09319_),
    .B1(net4865),
    .B2(\atari2600.ram[127][5] ),
    .A2(net4999),
    .A1(\atari2600.ram[124][5] ));
 sg13g2_a22oi_1 _17571_ (.Y(_09320_),
    .B1(net4819),
    .B2(\atari2600.ram[126][5] ),
    .A2(net4914),
    .A1(\atari2600.ram[125][5] ));
 sg13g2_a21oi_2 _17572_ (.B1(net4956),
    .Y(_09321_),
    .A2(_09320_),
    .A1(_09319_));
 sg13g2_a22oi_1 _17573_ (.Y(_09322_),
    .B1(net4854),
    .B2(\atari2600.ram[115][5] ),
    .A2(net4984),
    .A1(\atari2600.ram[112][5] ));
 sg13g2_a22oi_1 _17574_ (.Y(_09323_),
    .B1(net4810),
    .B2(\atari2600.ram[114][5] ),
    .A2(net4903),
    .A1(\atari2600.ram[113][5] ));
 sg13g2_a21oi_1 _17575_ (.A1(_09322_),
    .A2(_09323_),
    .Y(_09324_),
    .B1(net4930));
 sg13g2_nor2_1 _17576_ (.A(net5025),
    .B(_09321_),
    .Y(_09325_));
 sg13g2_nor3_1 _17577_ (.A(_09315_),
    .B(_09318_),
    .C(_09324_),
    .Y(_09326_));
 sg13g2_a22oi_1 _17578_ (.Y(_09327_),
    .B1(net4856),
    .B2(\atari2600.ram[111][5] ),
    .A2(net4987),
    .A1(\atari2600.ram[108][5] ));
 sg13g2_a22oi_1 _17579_ (.Y(_09328_),
    .B1(net4811),
    .B2(\atari2600.ram[110][5] ),
    .A2(net4905),
    .A1(\atari2600.ram[109][5] ));
 sg13g2_a21oi_1 _17580_ (.A1(_09327_),
    .A2(_09328_),
    .Y(_09329_),
    .B1(net4956));
 sg13g2_a22oi_1 _17581_ (.Y(_09330_),
    .B1(net4854),
    .B2(\atari2600.ram[99][5] ),
    .A2(net4984),
    .A1(\atari2600.ram[96][5] ));
 sg13g2_a22oi_1 _17582_ (.Y(_09331_),
    .B1(net4809),
    .B2(\atari2600.ram[98][5] ),
    .A2(net4903),
    .A1(\atari2600.ram[97][5] ));
 sg13g2_a21o_2 _17583_ (.A2(_09331_),
    .A1(_09330_),
    .B1(net4931),
    .X(_09332_));
 sg13g2_a22oi_1 _17584_ (.Y(_09333_),
    .B1(net4988),
    .B2(\atari2600.ram[100][5] ),
    .A2(net4905),
    .A1(\atari2600.ram[101][5] ));
 sg13g2_a22oi_1 _17585_ (.Y(_09334_),
    .B1(net4809),
    .B2(\atari2600.ram[102][5] ),
    .A2(net4856),
    .A1(\atari2600.ram[103][5] ));
 sg13g2_a21oi_1 _17586_ (.A1(_09333_),
    .A2(_09334_),
    .Y(_09335_),
    .B1(net5013));
 sg13g2_a22oi_1 _17587_ (.Y(_09336_),
    .B1(net4854),
    .B2(\atari2600.ram[107][5] ),
    .A2(net4984),
    .A1(\atari2600.ram[104][5] ));
 sg13g2_a22oi_1 _17588_ (.Y(_09337_),
    .B1(net4813),
    .B2(\atari2600.ram[106][5] ),
    .A2(net4908),
    .A1(\atari2600.ram[105][5] ));
 sg13g2_a21oi_2 _17589_ (.B1(net4943),
    .Y(_09338_),
    .A2(_09337_),
    .A1(_09336_));
 sg13g2_nor4_2 _17590_ (.A(net5027),
    .B(_09329_),
    .C(_09335_),
    .Y(_09339_),
    .D(_09338_));
 sg13g2_a221oi_1 _17591_ (.B2(_09339_),
    .C1(net4879),
    .B1(_09332_),
    .A1(_09325_),
    .Y(_09340_),
    .A2(_09326_));
 sg13g2_a22oi_1 _17592_ (.Y(_09341_),
    .B1(net4847),
    .B2(\atari2600.ram[87][5] ),
    .A2(net4977),
    .A1(\atari2600.ram[84][5] ));
 sg13g2_a22oi_1 _17593_ (.Y(_09342_),
    .B1(net4803),
    .B2(\atari2600.ram[86][5] ),
    .A2(net4898),
    .A1(\atari2600.ram[85][5] ));
 sg13g2_a21oi_2 _17594_ (.B1(net5009),
    .Y(_09343_),
    .A2(_09342_),
    .A1(_09341_));
 sg13g2_a22oi_1 _17595_ (.Y(_09344_),
    .B1(net4868),
    .B2(\atari2600.ram[95][5] ),
    .A2(net4997),
    .A1(\atari2600.ram[92][5] ));
 sg13g2_a22oi_1 _17596_ (.Y(_09345_),
    .B1(net4822),
    .B2(\atari2600.ram[94][5] ),
    .A2(net4917),
    .A1(\atari2600.ram[93][5] ));
 sg13g2_a21oi_2 _17597_ (.B1(net4957),
    .Y(_09346_),
    .A2(_09345_),
    .A1(_09344_));
 sg13g2_a22oi_1 _17598_ (.Y(_09347_),
    .B1(net4864),
    .B2(\atari2600.ram[83][5] ),
    .A2(net4995),
    .A1(\atari2600.ram[80][5] ));
 sg13g2_a22oi_1 _17599_ (.Y(_09348_),
    .B1(net4821),
    .B2(\atari2600.ram[82][5] ),
    .A2(net4916),
    .A1(\atari2600.ram[81][5] ));
 sg13g2_a21oi_1 _17600_ (.A1(_09347_),
    .A2(_09348_),
    .Y(_09349_),
    .B1(net4933));
 sg13g2_a22oi_1 _17601_ (.Y(_09350_),
    .B1(net4867),
    .B2(\atari2600.ram[91][5] ),
    .A2(net4997),
    .A1(\atari2600.ram[88][5] ));
 sg13g2_a22oi_1 _17602_ (.Y(_09351_),
    .B1(net4820),
    .B2(\atari2600.ram[90][5] ),
    .A2(net4915),
    .A1(\atari2600.ram[89][5] ));
 sg13g2_a21oi_2 _17603_ (.B1(net4942),
    .Y(_09352_),
    .A2(_09351_),
    .A1(_09350_));
 sg13g2_nor4_2 _17604_ (.A(_09343_),
    .B(_09346_),
    .C(_09349_),
    .Y(_09353_),
    .D(_09352_));
 sg13g2_a22oi_1 _17605_ (.Y(_09354_),
    .B1(net4869),
    .B2(\atari2600.ram[71][5] ),
    .A2(net5000),
    .A1(\atari2600.ram[68][5] ));
 sg13g2_a22oi_1 _17606_ (.Y(_09355_),
    .B1(net4825),
    .B2(\atari2600.ram[70][5] ),
    .A2(net4920),
    .A1(\atari2600.ram[69][5] ));
 sg13g2_a21oi_2 _17607_ (.B1(net5015),
    .Y(_09356_),
    .A2(_09355_),
    .A1(_09354_));
 sg13g2_a22oi_1 _17608_ (.Y(_09357_),
    .B1(net4868),
    .B2(\atari2600.ram[75][5] ),
    .A2(net4998),
    .A1(\atari2600.ram[72][5] ));
 sg13g2_a22oi_1 _17609_ (.Y(_09358_),
    .B1(net4823),
    .B2(\atari2600.ram[74][5] ),
    .A2(net4918),
    .A1(\atari2600.ram[73][5] ));
 sg13g2_a21oi_1 _17610_ (.A1(_09357_),
    .A2(_09358_),
    .Y(_09359_),
    .B1(net4945));
 sg13g2_a22oi_1 _17611_ (.Y(_09360_),
    .B1(net4871),
    .B2(\atari2600.ram[79][5] ),
    .A2(net5002),
    .A1(\atari2600.ram[76][5] ));
 sg13g2_a22oi_1 _17612_ (.Y(_09361_),
    .B1(net4822),
    .B2(\atari2600.ram[78][5] ),
    .A2(net4917),
    .A1(\atari2600.ram[77][5] ));
 sg13g2_a21oi_2 _17613_ (.B1(net4957),
    .Y(_09362_),
    .A2(_09361_),
    .A1(_09360_));
 sg13g2_a22oi_1 _17614_ (.Y(_09363_),
    .B1(net4865),
    .B2(\atari2600.ram[67][5] ),
    .A2(net4996),
    .A1(\atari2600.ram[64][5] ));
 sg13g2_a22oi_1 _17615_ (.Y(_09364_),
    .B1(net4818),
    .B2(\atari2600.ram[66][5] ),
    .A2(net4913),
    .A1(\atari2600.ram[65][5] ));
 sg13g2_a21oi_1 _17616_ (.A1(_09363_),
    .A2(_09364_),
    .Y(_09365_),
    .B1(net4933));
 sg13g2_nor4_1 _17617_ (.A(_09356_),
    .B(_09359_),
    .C(_09362_),
    .D(_09365_),
    .Y(_09366_));
 sg13g2_nor2_1 _17618_ (.A(net4778),
    .B(_09366_),
    .Y(_09367_));
 sg13g2_o21ai_1 _17619_ (.B1(net5020),
    .Y(_09368_),
    .A1(net4775),
    .A2(_09353_));
 sg13g2_nor3_2 _17620_ (.A(_09340_),
    .B(_09367_),
    .C(_09368_),
    .Y(_09369_));
 sg13g2_a22oi_1 _17621_ (.Y(_09370_),
    .B1(net4844),
    .B2(\atari2600.ram[3][5] ),
    .A2(net4974),
    .A1(\atari2600.ram[0][5] ));
 sg13g2_a22oi_1 _17622_ (.Y(_09371_),
    .B1(net4800),
    .B2(\atari2600.ram[2][5] ),
    .A2(net4894),
    .A1(\atari2600.ram[1][5] ));
 sg13g2_a21oi_1 _17623_ (.A1(_09370_),
    .A2(_09371_),
    .Y(_09372_),
    .B1(net4927));
 sg13g2_a22oi_1 _17624_ (.Y(_09373_),
    .B1(net4835),
    .B2(\atari2600.ram[15][5] ),
    .A2(net4965),
    .A1(\atari2600.ram[12][5] ));
 sg13g2_a22oi_1 _17625_ (.Y(_09374_),
    .B1(net4789),
    .B2(\atari2600.ram[14][5] ),
    .A2(net4883),
    .A1(\atari2600.ram[13][5] ));
 sg13g2_a21oi_1 _17626_ (.A1(_09373_),
    .A2(_09374_),
    .Y(_09375_),
    .B1(net4950));
 sg13g2_a22oi_1 _17627_ (.Y(_09376_),
    .B1(net4834),
    .B2(\atari2600.ram[11][5] ),
    .A2(net4964),
    .A1(\atari2600.ram[8][5] ));
 sg13g2_a22oi_1 _17628_ (.Y(_09377_),
    .B1(net4789),
    .B2(\atari2600.ram[10][5] ),
    .A2(net4884),
    .A1(\atari2600.ram[9][5] ));
 sg13g2_a21oi_1 _17629_ (.A1(_09376_),
    .A2(_09377_),
    .Y(_09378_),
    .B1(net4938));
 sg13g2_a22oi_1 _17630_ (.Y(_09379_),
    .B1(net4843),
    .B2(\atari2600.ram[7][5] ),
    .A2(net4973),
    .A1(\atari2600.ram[4][5] ));
 sg13g2_a22oi_1 _17631_ (.Y(_09380_),
    .B1(net4799),
    .B2(\atari2600.ram[6][5] ),
    .A2(net4893),
    .A1(\atari2600.ram[5][5] ));
 sg13g2_a21oi_1 _17632_ (.A1(_09379_),
    .A2(_09380_),
    .Y(_09381_),
    .B1(net5007));
 sg13g2_nor4_1 _17633_ (.A(_09372_),
    .B(_09375_),
    .C(_09378_),
    .D(_09381_),
    .Y(_09382_));
 sg13g2_nor2_1 _17634_ (.A(net4777),
    .B(_09382_),
    .Y(_09383_));
 sg13g2_a22oi_1 _17635_ (.Y(_09384_),
    .B1(net4839),
    .B2(\atari2600.ram[63][5] ),
    .A2(net4968),
    .A1(\atari2600.ram[60][5] ));
 sg13g2_a22oi_1 _17636_ (.Y(_09385_),
    .B1(net4793),
    .B2(\atari2600.ram[62][5] ),
    .A2(net4886),
    .A1(\atari2600.ram[61][5] ));
 sg13g2_a21oi_1 _17637_ (.A1(_09384_),
    .A2(_09385_),
    .Y(_09386_),
    .B1(net4953));
 sg13g2_a22oi_1 _17638_ (.Y(_09387_),
    .B1(net4838),
    .B2(\atari2600.ram[59][5] ),
    .A2(net4968),
    .A1(\atari2600.ram[56][5] ));
 sg13g2_a22oi_1 _17639_ (.Y(_09388_),
    .B1(net4792),
    .B2(\atari2600.ram[58][5] ),
    .A2(net4886),
    .A1(\atari2600.ram[57][5] ));
 sg13g2_a21oi_2 _17640_ (.B1(net4940),
    .Y(_09389_),
    .A2(_09388_),
    .A1(_09387_));
 sg13g2_a22oi_1 _17641_ (.Y(_09390_),
    .B1(net4841),
    .B2(\atari2600.ram[51][5] ),
    .A2(net4972),
    .A1(\atari2600.ram[48][5] ));
 sg13g2_a22oi_1 _17642_ (.Y(_09391_),
    .B1(net4794),
    .B2(\atari2600.ram[50][5] ),
    .A2(net4888),
    .A1(\atari2600.ram[49][5] ));
 sg13g2_a21oi_1 _17643_ (.A1(_09390_),
    .A2(_09391_),
    .Y(_09392_),
    .B1(net4926));
 sg13g2_a22oi_1 _17644_ (.Y(_09393_),
    .B1(net4857),
    .B2(\atari2600.ram[55][5] ),
    .A2(net4986),
    .A1(\atari2600.ram[52][5] ));
 sg13g2_a22oi_1 _17645_ (.Y(_09394_),
    .B1(net4810),
    .B2(\atari2600.ram[54][5] ),
    .A2(net4904),
    .A1(\atari2600.ram[53][5] ));
 sg13g2_a21oi_1 _17646_ (.A1(_09393_),
    .A2(_09394_),
    .Y(_09395_),
    .B1(net5012));
 sg13g2_nor4_2 _17647_ (.A(_09386_),
    .B(_09389_),
    .C(_09392_),
    .Y(_09396_),
    .D(_09395_));
 sg13g2_nor2_2 _17648_ (.A(net4776),
    .B(_09396_),
    .Y(_09397_));
 sg13g2_a22oi_1 _17649_ (.Y(_09398_),
    .B1(net4831),
    .B2(\atari2600.ram[39][5] ),
    .A2(net4961),
    .A1(\atari2600.ram[36][5] ));
 sg13g2_a22oi_1 _17650_ (.Y(_09399_),
    .B1(net4786),
    .B2(\atari2600.ram[38][5] ),
    .A2(net4882),
    .A1(\atari2600.ram[37][5] ));
 sg13g2_a21oi_2 _17651_ (.B1(net5006),
    .Y(_09400_),
    .A2(_09399_),
    .A1(_09398_));
 sg13g2_a22oi_1 _17652_ (.Y(_09401_),
    .B1(net4834),
    .B2(\atari2600.ram[43][5] ),
    .A2(net4964),
    .A1(\atari2600.ram[40][5] ));
 sg13g2_a22oi_1 _17653_ (.Y(_09402_),
    .B1(net4790),
    .B2(\atari2600.ram[42][5] ),
    .A2(net4884),
    .A1(\atari2600.ram[41][5] ));
 sg13g2_a21oi_1 _17654_ (.A1(_09401_),
    .A2(_09402_),
    .Y(_09403_),
    .B1(net4938));
 sg13g2_a22oi_1 _17655_ (.Y(_09404_),
    .B1(net4835),
    .B2(\atari2600.ram[47][5] ),
    .A2(net4965),
    .A1(\atari2600.ram[44][5] ));
 sg13g2_a22oi_1 _17656_ (.Y(_09405_),
    .B1(net4789),
    .B2(\atari2600.ram[46][5] ),
    .A2(net4883),
    .A1(\atari2600.ram[45][5] ));
 sg13g2_a21oi_1 _17657_ (.A1(_09404_),
    .A2(_09405_),
    .Y(_09406_),
    .B1(net4949));
 sg13g2_a22oi_1 _17658_ (.Y(_09407_),
    .B1(net4832),
    .B2(\atari2600.ram[35][5] ),
    .A2(net4962),
    .A1(\atari2600.ram[32][5] ));
 sg13g2_a22oi_1 _17659_ (.Y(_09408_),
    .B1(net4787),
    .B2(\atari2600.ram[34][5] ),
    .A2(net4881),
    .A1(\atari2600.ram[33][5] ));
 sg13g2_a21oi_2 _17660_ (.B1(net4925),
    .Y(_09409_),
    .A2(_09408_),
    .A1(_09407_));
 sg13g2_nor4_2 _17661_ (.A(_09400_),
    .B(_09403_),
    .C(_09406_),
    .Y(_09410_),
    .D(_09409_));
 sg13g2_a22oi_1 _17662_ (.Y(_09411_),
    .B1(net4847),
    .B2(\atari2600.ram[31][5] ),
    .A2(net4978),
    .A1(\atari2600.ram[28][5] ));
 sg13g2_a22oi_1 _17663_ (.Y(_09412_),
    .B1(net4806),
    .B2(\atari2600.ram[30][5] ),
    .A2(net4900),
    .A1(\atari2600.ram[29][5] ));
 sg13g2_a21oi_1 _17664_ (.A1(_09411_),
    .A2(_09412_),
    .Y(_09413_),
    .B1(net4952));
 sg13g2_a22oi_1 _17665_ (.Y(_09414_),
    .B1(net4845),
    .B2(\atari2600.ram[19][5] ),
    .A2(net4975),
    .A1(\atari2600.ram[16][5] ));
 sg13g2_a22oi_1 _17666_ (.Y(_09415_),
    .B1(net4800),
    .B2(\atari2600.ram[18][5] ),
    .A2(net4895),
    .A1(\atari2600.ram[17][5] ));
 sg13g2_a21oi_2 _17667_ (.B1(net4928),
    .Y(_09416_),
    .A2(_09415_),
    .A1(_09414_));
 sg13g2_a22oi_1 _17668_ (.Y(_09417_),
    .B1(net4846),
    .B2(\atari2600.ram[23][5] ),
    .A2(net4976),
    .A1(\atari2600.ram[20][5] ));
 sg13g2_a22oi_1 _17669_ (.Y(_09418_),
    .B1(net4801),
    .B2(\atari2600.ram[22][5] ),
    .A2(net4896),
    .A1(\atari2600.ram[21][5] ));
 sg13g2_a21oi_1 _17670_ (.A1(_09417_),
    .A2(_09418_),
    .Y(_09419_),
    .B1(net5008));
 sg13g2_a22oi_1 _17671_ (.Y(_09420_),
    .B1(net4841),
    .B2(\atari2600.ram[27][5] ),
    .A2(net4971),
    .A1(\atari2600.ram[24][5] ));
 sg13g2_a22oi_1 _17672_ (.Y(_09421_),
    .B1(net4795),
    .B2(\atari2600.ram[26][5] ),
    .A2(net4889),
    .A1(\atari2600.ram[25][5] ));
 sg13g2_a21oi_2 _17673_ (.B1(net4939),
    .Y(_09422_),
    .A2(_09421_),
    .A1(_09420_));
 sg13g2_nor4_1 _17674_ (.A(_09413_),
    .B(_09416_),
    .C(_09419_),
    .D(_09422_),
    .Y(_09423_));
 sg13g2_nor2_1 _17675_ (.A(net4774),
    .B(_09423_),
    .Y(_09424_));
 sg13g2_o21ai_1 _17676_ (.B1(net5023),
    .Y(_09425_),
    .A1(net4772),
    .A2(_09410_));
 sg13g2_nor4_2 _17677_ (.A(_09383_),
    .B(_09397_),
    .C(_09424_),
    .Y(_09426_),
    .D(_09425_));
 sg13g2_nor2_2 _17678_ (.A(_09369_),
    .B(_09426_),
    .Y(_00006_));
 sg13g2_a22oi_1 _17679_ (.Y(_09427_),
    .B1(net4856),
    .B2(\atari2600.ram[123][6] ),
    .A2(net4986),
    .A1(\atari2600.ram[120][6] ));
 sg13g2_a22oi_1 _17680_ (.Y(_09428_),
    .B1(net4811),
    .B2(\atari2600.ram[122][6] ),
    .A2(net4905),
    .A1(\atari2600.ram[121][6] ));
 sg13g2_a21oi_1 _17681_ (.A1(_09427_),
    .A2(_09428_),
    .Y(_09429_),
    .B1(net4943));
 sg13g2_a22oi_1 _17682_ (.Y(_09430_),
    .B1(net4857),
    .B2(\atari2600.ram[119][6] ),
    .A2(net4986),
    .A1(\atari2600.ram[116][6] ));
 sg13g2_a22oi_1 _17683_ (.Y(_09431_),
    .B1(net4812),
    .B2(\atari2600.ram[118][6] ),
    .A2(net4907),
    .A1(\atari2600.ram[117][6] ));
 sg13g2_a21oi_1 _17684_ (.A1(_09430_),
    .A2(_09431_),
    .Y(_09432_),
    .B1(net5013));
 sg13g2_a22oi_1 _17685_ (.Y(_09433_),
    .B1(net4853),
    .B2(\atari2600.ram[115][6] ),
    .A2(net4983),
    .A1(\atari2600.ram[112][6] ));
 sg13g2_a22oi_1 _17686_ (.Y(_09434_),
    .B1(net4808),
    .B2(\atari2600.ram[114][6] ),
    .A2(net4902),
    .A1(\atari2600.ram[113][6] ));
 sg13g2_a21oi_2 _17687_ (.B1(net4930),
    .Y(_09435_),
    .A2(_09434_),
    .A1(_09433_));
 sg13g2_a22oi_1 _17688_ (.Y(_09436_),
    .B1(net4863),
    .B2(\atari2600.ram[127][6] ),
    .A2(net4994),
    .A1(\atari2600.ram[124][6] ));
 sg13g2_a22oi_1 _17689_ (.Y(_09437_),
    .B1(net4818),
    .B2(\atari2600.ram[126][6] ),
    .A2(net4913),
    .A1(\atari2600.ram[125][6] ));
 sg13g2_a21oi_1 _17690_ (.A1(_09436_),
    .A2(_09437_),
    .Y(_09438_),
    .B1(net4956));
 sg13g2_nor4_1 _17691_ (.A(_09429_),
    .B(_09432_),
    .C(_09435_),
    .D(_09438_),
    .Y(_09439_));
 sg13g2_o21ai_1 _17692_ (.B1(net5021),
    .Y(_09440_),
    .A1(net4776),
    .A2(_09439_));
 sg13g2_a22oi_1 _17693_ (.Y(_09441_),
    .B1(net4861),
    .B2(\atari2600.ram[103][6] ),
    .A2(net4991),
    .A1(\atari2600.ram[100][6] ));
 sg13g2_a22oi_1 _17694_ (.Y(_09442_),
    .B1(net4816),
    .B2(\atari2600.ram[102][6] ),
    .A2(net4910),
    .A1(\atari2600.ram[101][6] ));
 sg13g2_a21oi_1 _17695_ (.A1(_09441_),
    .A2(_09442_),
    .Y(_09443_),
    .B1(net5014));
 sg13g2_a22oi_1 _17696_ (.Y(_09444_),
    .B1(net4861),
    .B2(\atari2600.ram[111][6] ),
    .A2(net4991),
    .A1(\atari2600.ram[108][6] ));
 sg13g2_a22oi_1 _17697_ (.Y(_09445_),
    .B1(net4816),
    .B2(\atari2600.ram[110][6] ),
    .A2(net4911),
    .A1(\atari2600.ram[109][6] ));
 sg13g2_a21oi_1 _17698_ (.A1(_09444_),
    .A2(_09445_),
    .Y(_09446_),
    .B1(net4954));
 sg13g2_a22oi_1 _17699_ (.Y(_09447_),
    .B1(net4859),
    .B2(\atari2600.ram[107][6] ),
    .A2(net4989),
    .A1(\atari2600.ram[104][6] ));
 sg13g2_a22oi_1 _17700_ (.Y(_09448_),
    .B1(net4814),
    .B2(\atari2600.ram[106][6] ),
    .A2(net4908),
    .A1(\atari2600.ram[105][6] ));
 sg13g2_a21oi_1 _17701_ (.A1(_09447_),
    .A2(_09448_),
    .Y(_09449_),
    .B1(net4944));
 sg13g2_a22oi_1 _17702_ (.Y(_09450_),
    .B1(net4860),
    .B2(\atari2600.ram[99][6] ),
    .A2(net4989),
    .A1(\atari2600.ram[96][6] ));
 sg13g2_a22oi_1 _17703_ (.Y(_09451_),
    .B1(net4813),
    .B2(\atari2600.ram[98][6] ),
    .A2(net4908),
    .A1(\atari2600.ram[97][6] ));
 sg13g2_a21oi_2 _17704_ (.B1(net4932),
    .Y(_09452_),
    .A2(_09451_),
    .A1(_09450_));
 sg13g2_nor4_2 _17705_ (.A(_09443_),
    .B(_09446_),
    .C(_09449_),
    .Y(_09453_),
    .D(_09452_));
 sg13g2_nor2_2 _17706_ (.A(net4772),
    .B(_09453_),
    .Y(_09454_));
 sg13g2_a22oi_1 _17707_ (.Y(_09455_),
    .B1(net4873),
    .B2(\atari2600.ram[79][6] ),
    .A2(net5002),
    .A1(\atari2600.ram[76][6] ));
 sg13g2_a22oi_1 _17708_ (.Y(_09456_),
    .B1(net4828),
    .B2(\atari2600.ram[78][6] ),
    .A2(net4923),
    .A1(\atari2600.ram[77][6] ));
 sg13g2_a21oi_2 _17709_ (.B1(net4959),
    .Y(_09457_),
    .A2(_09456_),
    .A1(_09455_));
 sg13g2_a22oi_1 _17710_ (.Y(_09458_),
    .B1(net4870),
    .B2(\atari2600.ram[71][6] ),
    .A2(net5001),
    .A1(\atari2600.ram[68][6] ));
 sg13g2_a22oi_1 _17711_ (.Y(_09459_),
    .B1(net4826),
    .B2(\atari2600.ram[70][6] ),
    .A2(net4921),
    .A1(\atari2600.ram[69][6] ));
 sg13g2_a21oi_1 _17712_ (.A1(_09458_),
    .A2(_09459_),
    .Y(_09460_),
    .B1(net5015));
 sg13g2_a22oi_1 _17713_ (.Y(_09461_),
    .B1(net4870),
    .B2(\atari2600.ram[67][6] ),
    .A2(net5001),
    .A1(\atari2600.ram[64][6] ));
 sg13g2_a22oi_1 _17714_ (.Y(_09462_),
    .B1(net4825),
    .B2(\atari2600.ram[66][6] ),
    .A2(net4920),
    .A1(\atari2600.ram[65][6] ));
 sg13g2_a21oi_1 _17715_ (.A1(_09461_),
    .A2(_09462_),
    .Y(_09463_),
    .B1(net4934));
 sg13g2_a22oi_1 _17716_ (.Y(_09464_),
    .B1(net4873),
    .B2(\atari2600.ram[75][6] ),
    .A2(net5004),
    .A1(\atari2600.ram[72][6] ));
 sg13g2_a22oi_1 _17717_ (.Y(_09465_),
    .B1(net4828),
    .B2(\atari2600.ram[74][6] ),
    .A2(net4923),
    .A1(\atari2600.ram[73][6] ));
 sg13g2_a21oi_2 _17718_ (.B1(net4945),
    .Y(_09466_),
    .A2(_09465_),
    .A1(_09464_));
 sg13g2_nor4_2 _17719_ (.A(_09457_),
    .B(_09460_),
    .C(_09463_),
    .Y(_09467_),
    .D(_09466_));
 sg13g2_nor2_1 _17720_ (.A(net4779),
    .B(_09467_),
    .Y(_09468_));
 sg13g2_a22oi_1 _17721_ (.Y(_09469_),
    .B1(net4865),
    .B2(\atari2600.ram[83][6] ),
    .A2(net4996),
    .A1(\atari2600.ram[80][6] ));
 sg13g2_a22oi_1 _17722_ (.Y(_09470_),
    .B1(net4823),
    .B2(\atari2600.ram[82][6] ),
    .A2(net4918),
    .A1(\atari2600.ram[81][6] ));
 sg13g2_a21oi_1 _17723_ (.A1(_09469_),
    .A2(_09470_),
    .Y(_09471_),
    .B1(net4933));
 sg13g2_a22oi_1 _17724_ (.Y(_09472_),
    .B1(net4863),
    .B2(\atari2600.ram[87][6] ),
    .A2(net4994),
    .A1(\atari2600.ram[84][6] ));
 sg13g2_a22oi_1 _17725_ (.Y(_09473_),
    .B1(net4820),
    .B2(\atari2600.ram[86][6] ),
    .A2(net4915),
    .A1(\atari2600.ram[85][6] ));
 sg13g2_a21oi_1 _17726_ (.A1(_09472_),
    .A2(_09473_),
    .Y(_09474_),
    .B1(net5016));
 sg13g2_a22oi_1 _17727_ (.Y(_09475_),
    .B1(net4867),
    .B2(\atari2600.ram[95][6] ),
    .A2(net4997),
    .A1(\atari2600.ram[92][6] ));
 sg13g2_a22oi_1 _17728_ (.Y(_09476_),
    .B1(net4822),
    .B2(\atari2600.ram[94][6] ),
    .A2(net4917),
    .A1(\atari2600.ram[93][6] ));
 sg13g2_a21oi_2 _17729_ (.B1(net4957),
    .Y(_09477_),
    .A2(_09476_),
    .A1(_09475_));
 sg13g2_a22oi_1 _17730_ (.Y(_09478_),
    .B1(net4850),
    .B2(\atari2600.ram[91][6] ),
    .A2(net4980),
    .A1(\atari2600.ram[88][6] ));
 sg13g2_a22oi_1 _17731_ (.Y(_09479_),
    .B1(net4804),
    .B2(\atari2600.ram[90][6] ),
    .A2(net4898),
    .A1(\atari2600.ram[89][6] ));
 sg13g2_a21oi_2 _17732_ (.B1(net4941),
    .Y(_09480_),
    .A2(_09479_),
    .A1(_09478_));
 sg13g2_nor4_2 _17733_ (.A(_09471_),
    .B(_09474_),
    .C(_09477_),
    .Y(_09481_),
    .D(_09480_));
 sg13g2_nor2_1 _17734_ (.A(net4774),
    .B(_09481_),
    .Y(_09482_));
 sg13g2_nor4_2 _17735_ (.A(_09440_),
    .B(_09454_),
    .C(_09468_),
    .Y(_09483_),
    .D(_09482_));
 sg13g2_a22oi_1 _17736_ (.Y(_09484_),
    .B1(net4830),
    .B2(\atari2600.ram[39][6] ),
    .A2(net4960),
    .A1(\atari2600.ram[36][6] ));
 sg13g2_a22oi_1 _17737_ (.Y(_09485_),
    .B1(net4785),
    .B2(\atari2600.ram[38][6] ),
    .A2(net4880),
    .A1(\atari2600.ram[37][6] ));
 sg13g2_a21oi_2 _17738_ (.B1(net5006),
    .Y(_09486_),
    .A2(_09485_),
    .A1(_09484_));
 sg13g2_a22oi_1 _17739_ (.Y(_09487_),
    .B1(net4832),
    .B2(\atari2600.ram[47][6] ),
    .A2(net4962),
    .A1(\atari2600.ram[44][6] ));
 sg13g2_a22oi_1 _17740_ (.Y(_09488_),
    .B1(net4790),
    .B2(\atari2600.ram[46][6] ),
    .A2(net4884),
    .A1(\atari2600.ram[45][6] ));
 sg13g2_a21oi_1 _17741_ (.A1(_09487_),
    .A2(_09488_),
    .Y(_09489_),
    .B1(net4949));
 sg13g2_a22oi_1 _17742_ (.Y(_09490_),
    .B1(net4832),
    .B2(\atari2600.ram[43][6] ),
    .A2(net4962),
    .A1(\atari2600.ram[40][6] ));
 sg13g2_a22oi_1 _17743_ (.Y(_09491_),
    .B1(net4787),
    .B2(\atari2600.ram[42][6] ),
    .A2(net4881),
    .A1(\atari2600.ram[41][6] ));
 sg13g2_a21oi_1 _17744_ (.A1(_09490_),
    .A2(_09491_),
    .Y(_09492_),
    .B1(net4937));
 sg13g2_a22oi_1 _17745_ (.Y(_09493_),
    .B1(net4832),
    .B2(\atari2600.ram[35][6] ),
    .A2(net4962),
    .A1(\atari2600.ram[32][6] ));
 sg13g2_a22oi_1 _17746_ (.Y(_09494_),
    .B1(net4787),
    .B2(\atari2600.ram[34][6] ),
    .A2(net4881),
    .A1(\atari2600.ram[33][6] ));
 sg13g2_a21oi_1 _17747_ (.A1(_09493_),
    .A2(_09494_),
    .Y(_09495_),
    .B1(net4925));
 sg13g2_nor4_2 _17748_ (.A(_09486_),
    .B(_09489_),
    .C(_09492_),
    .Y(_09496_),
    .D(_09495_));
 sg13g2_nor2_1 _17749_ (.A(net4772),
    .B(_09496_),
    .Y(_09497_));
 sg13g2_a22oi_1 _17750_ (.Y(_09498_),
    .B1(net4846),
    .B2(\atari2600.ram[23][6] ),
    .A2(net4976),
    .A1(\atari2600.ram[20][6] ));
 sg13g2_a22oi_1 _17751_ (.Y(_09499_),
    .B1(net4801),
    .B2(\atari2600.ram[22][6] ),
    .A2(net4896),
    .A1(\atari2600.ram[21][6] ));
 sg13g2_a21oi_1 _17752_ (.A1(_09498_),
    .A2(_09499_),
    .Y(_09500_),
    .B1(net5009));
 sg13g2_a22oi_1 _17753_ (.Y(_09501_),
    .B1(net4841),
    .B2(\atari2600.ram[27][6] ),
    .A2(net4971),
    .A1(\atari2600.ram[24][6] ));
 sg13g2_a22oi_1 _17754_ (.Y(_09502_),
    .B1(net4794),
    .B2(\atari2600.ram[26][6] ),
    .A2(net4888),
    .A1(\atari2600.ram[25][6] ));
 sg13g2_a21oi_1 _17755_ (.A1(_09501_),
    .A2(_09502_),
    .Y(_09503_),
    .B1(net4938));
 sg13g2_a22oi_1 _17756_ (.Y(_09504_),
    .B1(net4846),
    .B2(\atari2600.ram[31][6] ),
    .A2(net4976),
    .A1(\atari2600.ram[28][6] ));
 sg13g2_a22oi_1 _17757_ (.Y(_09505_),
    .B1(net4801),
    .B2(\atari2600.ram[30][6] ),
    .A2(net4896),
    .A1(\atari2600.ram[29][6] ));
 sg13g2_a21oi_1 _17758_ (.A1(_09504_),
    .A2(_09505_),
    .Y(_09506_),
    .B1(net4952));
 sg13g2_a22oi_1 _17759_ (.Y(_09507_),
    .B1(net4849),
    .B2(\atari2600.ram[19][6] ),
    .A2(net4980),
    .A1(\atari2600.ram[16][6] ));
 sg13g2_a22oi_1 _17760_ (.Y(_09508_),
    .B1(net4800),
    .B2(\atari2600.ram[18][6] ),
    .A2(net4895),
    .A1(\atari2600.ram[17][6] ));
 sg13g2_a21oi_2 _17761_ (.B1(net4928),
    .Y(_09509_),
    .A2(_09508_),
    .A1(_09507_));
 sg13g2_nor4_1 _17762_ (.A(_09500_),
    .B(_09503_),
    .C(_09506_),
    .D(_09509_),
    .Y(_09510_));
 sg13g2_nor2_1 _17763_ (.A(net4773),
    .B(_09510_),
    .Y(_09511_));
 sg13g2_a22oi_1 _17764_ (.Y(_09512_),
    .B1(net4843),
    .B2(\atari2600.ram[7][6] ),
    .A2(net4973),
    .A1(\atari2600.ram[4][6] ));
 sg13g2_a22oi_1 _17765_ (.Y(_09513_),
    .B1(net4799),
    .B2(\atari2600.ram[6][6] ),
    .A2(net4893),
    .A1(\atari2600.ram[5][6] ));
 sg13g2_a21oi_1 _17766_ (.A1(_09512_),
    .A2(_09513_),
    .Y(_09514_),
    .B1(net5007));
 sg13g2_a22oi_1 _17767_ (.Y(_09515_),
    .B1(net4836),
    .B2(\atari2600.ram[15][6] ),
    .A2(net4964),
    .A1(\atari2600.ram[12][6] ));
 sg13g2_a22oi_1 _17768_ (.Y(_09516_),
    .B1(net4790),
    .B2(\atari2600.ram[14][6] ),
    .A2(net4892),
    .A1(\atari2600.ram[13][6] ));
 sg13g2_a21oi_1 _17769_ (.A1(_09515_),
    .A2(_09516_),
    .Y(_09517_),
    .B1(net4950));
 sg13g2_a22oi_1 _17770_ (.Y(_09518_),
    .B1(net4840),
    .B2(\atari2600.ram[11][6] ),
    .A2(net4971),
    .A1(\atari2600.ram[8][6] ));
 sg13g2_a22oi_1 _17771_ (.Y(_09519_),
    .B1(net4801),
    .B2(\atari2600.ram[10][6] ),
    .A2(net4896),
    .A1(\atari2600.ram[9][6] ));
 sg13g2_a21oi_1 _17772_ (.A1(_09518_),
    .A2(_09519_),
    .Y(_09520_),
    .B1(net4941));
 sg13g2_a22oi_1 _17773_ (.Y(_09521_),
    .B1(net4844),
    .B2(\atari2600.ram[3][6] ),
    .A2(net4974),
    .A1(\atari2600.ram[0][6] ));
 sg13g2_a22oi_1 _17774_ (.Y(_09522_),
    .B1(net4798),
    .B2(\atari2600.ram[2][6] ),
    .A2(net4892),
    .A1(\atari2600.ram[1][6] ));
 sg13g2_a21oi_1 _17775_ (.A1(_09521_),
    .A2(_09522_),
    .Y(_09523_),
    .B1(net4927));
 sg13g2_nor4_1 _17776_ (.A(_09514_),
    .B(_09517_),
    .C(_09520_),
    .D(_09523_),
    .Y(_09524_));
 sg13g2_a22oi_1 _17777_ (.Y(_09525_),
    .B1(net4838),
    .B2(\atari2600.ram[59][6] ),
    .A2(net4968),
    .A1(\atari2600.ram[56][6] ));
 sg13g2_a22oi_1 _17778_ (.Y(_09526_),
    .B1(net4792),
    .B2(\atari2600.ram[58][6] ),
    .A2(net4886),
    .A1(\atari2600.ram[57][6] ));
 sg13g2_a21oi_2 _17779_ (.B1(net4940),
    .Y(_09527_),
    .A2(_09526_),
    .A1(_09525_));
 sg13g2_a22oi_1 _17780_ (.Y(_09528_),
    .B1(net4841),
    .B2(\atari2600.ram[51][6] ),
    .A2(net4972),
    .A1(\atari2600.ram[48][6] ));
 sg13g2_a22oi_1 _17781_ (.Y(_09529_),
    .B1(net4794),
    .B2(\atari2600.ram[50][6] ),
    .A2(net4888),
    .A1(\atari2600.ram[49][6] ));
 sg13g2_a21oi_1 _17782_ (.A1(_09528_),
    .A2(_09529_),
    .Y(_09530_),
    .B1(net4926));
 sg13g2_a22oi_1 _17783_ (.Y(_09531_),
    .B1(net4838),
    .B2(\atari2600.ram[63][6] ),
    .A2(net4968),
    .A1(\atari2600.ram[60][6] ));
 sg13g2_a22oi_1 _17784_ (.Y(_09532_),
    .B1(net4793),
    .B2(\atari2600.ram[62][6] ),
    .A2(net4886),
    .A1(\atari2600.ram[61][6] ));
 sg13g2_a21oi_1 _17785_ (.A1(_09531_),
    .A2(_09532_),
    .Y(_09533_),
    .B1(net4951));
 sg13g2_a22oi_1 _17786_ (.Y(_09534_),
    .B1(net4842),
    .B2(\atari2600.ram[55][6] ),
    .A2(net4972),
    .A1(\atari2600.ram[52][6] ));
 sg13g2_a22oi_1 _17787_ (.Y(_09535_),
    .B1(net4792),
    .B2(\atari2600.ram[54][6] ),
    .A2(net4886),
    .A1(\atari2600.ram[53][6] ));
 sg13g2_a21oi_1 _17788_ (.A1(_09534_),
    .A2(_09535_),
    .Y(_09536_),
    .B1(net5011));
 sg13g2_nor4_2 _17789_ (.A(_09527_),
    .B(_09530_),
    .C(_09533_),
    .Y(_09537_),
    .D(_09536_));
 sg13g2_nor2_1 _17790_ (.A(net4776),
    .B(_09537_),
    .Y(_09538_));
 sg13g2_o21ai_1 _17791_ (.B1(net5023),
    .Y(_09539_),
    .A1(net4777),
    .A2(_09524_));
 sg13g2_nor4_1 _17792_ (.A(_09497_),
    .B(_09511_),
    .C(_09538_),
    .D(_09539_),
    .Y(_09540_));
 sg13g2_nor2_2 _17793_ (.A(_09483_),
    .B(_09540_),
    .Y(_00007_));
 sg13g2_a22oi_1 _17794_ (.Y(_09541_),
    .B1(net4869),
    .B2(\atari2600.ram[71][7] ),
    .A2(net5000),
    .A1(\atari2600.ram[68][7] ));
 sg13g2_a22oi_1 _17795_ (.Y(_09542_),
    .B1(net4825),
    .B2(\atari2600.ram[70][7] ),
    .A2(net4920),
    .A1(\atari2600.ram[69][7] ));
 sg13g2_a21oi_1 _17796_ (.A1(_09541_),
    .A2(_09542_),
    .Y(_09543_),
    .B1(net5015));
 sg13g2_a22oi_1 _17797_ (.Y(_09544_),
    .B1(net4869),
    .B2(\atari2600.ram[67][7] ),
    .A2(net5001),
    .A1(\atari2600.ram[64][7] ));
 sg13g2_a22oi_1 _17798_ (.Y(_09545_),
    .B1(net4825),
    .B2(\atari2600.ram[66][7] ),
    .A2(net4920),
    .A1(\atari2600.ram[65][7] ));
 sg13g2_a21oi_1 _17799_ (.A1(_09544_),
    .A2(_09545_),
    .Y(_09546_),
    .B1(net4935));
 sg13g2_a22oi_1 _17800_ (.Y(_09547_),
    .B1(net4871),
    .B2(\atari2600.ram[75][7] ),
    .A2(net5002),
    .A1(\atari2600.ram[72][7] ));
 sg13g2_a22oi_1 _17801_ (.Y(_09548_),
    .B1(net4827),
    .B2(\atari2600.ram[74][7] ),
    .A2(net4922),
    .A1(\atari2600.ram[73][7] ));
 sg13g2_a21oi_2 _17802_ (.B1(net4945),
    .Y(_09549_),
    .A2(_09548_),
    .A1(_09547_));
 sg13g2_a22oi_1 _17803_ (.Y(_09550_),
    .B1(net4872),
    .B2(\atari2600.ram[79][7] ),
    .A2(net5003),
    .A1(\atari2600.ram[76][7] ));
 sg13g2_a22oi_1 _17804_ (.Y(_09551_),
    .B1(net4828),
    .B2(\atari2600.ram[78][7] ),
    .A2(net4923),
    .A1(\atari2600.ram[77][7] ));
 sg13g2_a21oi_2 _17805_ (.B1(net4959),
    .Y(_09552_),
    .A2(_09551_),
    .A1(_09550_));
 sg13g2_nor4_2 _17806_ (.A(_09543_),
    .B(_09546_),
    .C(_09549_),
    .Y(_09553_),
    .D(_09552_));
 sg13g2_nor2_1 _17807_ (.A(net4779),
    .B(_09553_),
    .Y(_09554_));
 sg13g2_a22oi_1 _17808_ (.Y(_09555_),
    .B1(net4861),
    .B2(\atari2600.ram[111][7] ),
    .A2(net4991),
    .A1(\atari2600.ram[108][7] ));
 sg13g2_a22oi_1 _17809_ (.Y(_09556_),
    .B1(net4816),
    .B2(\atari2600.ram[110][7] ),
    .A2(net4910),
    .A1(\atari2600.ram[109][7] ));
 sg13g2_a21oi_2 _17810_ (.B1(net4955),
    .Y(_09557_),
    .A2(_09556_),
    .A1(_09555_));
 sg13g2_a22oi_1 _17811_ (.Y(_09558_),
    .B1(net4859),
    .B2(\atari2600.ram[103][7] ),
    .A2(net4989),
    .A1(\atari2600.ram[100][7] ));
 sg13g2_a22oi_1 _17812_ (.Y(_09559_),
    .B1(net4814),
    .B2(\atari2600.ram[102][7] ),
    .A2(net4909),
    .A1(\atari2600.ram[101][7] ));
 sg13g2_a21oi_1 _17813_ (.A1(_09558_),
    .A2(_09559_),
    .Y(_09560_),
    .B1(net5014));
 sg13g2_a22oi_1 _17814_ (.Y(_09561_),
    .B1(net4860),
    .B2(\atari2600.ram[99][7] ),
    .A2(net4990),
    .A1(\atari2600.ram[96][7] ));
 sg13g2_a22oi_1 _17815_ (.Y(_09562_),
    .B1(net4813),
    .B2(\atari2600.ram[98][7] ),
    .A2(net4908),
    .A1(\atari2600.ram[97][7] ));
 sg13g2_a21oi_2 _17816_ (.B1(net4932),
    .Y(_09563_),
    .A2(_09562_),
    .A1(_09561_));
 sg13g2_a22oi_1 _17817_ (.Y(_09564_),
    .B1(net4860),
    .B2(\atari2600.ram[107][7] ),
    .A2(net4990),
    .A1(\atari2600.ram[104][7] ));
 sg13g2_a22oi_1 _17818_ (.Y(_09565_),
    .B1(net4815),
    .B2(\atari2600.ram[106][7] ),
    .A2(net4909),
    .A1(\atari2600.ram[105][7] ));
 sg13g2_a21oi_1 _17819_ (.A1(_09564_),
    .A2(_09565_),
    .Y(_09566_),
    .B1(net4944));
 sg13g2_nor4_2 _17820_ (.A(_09557_),
    .B(_09560_),
    .C(_09563_),
    .Y(_09567_),
    .D(_09566_));
 sg13g2_nor2_1 _17821_ (.A(net4772),
    .B(_09567_),
    .Y(_09568_));
 sg13g2_a22oi_1 _17822_ (.Y(_09569_),
    .B1(net4867),
    .B2(\atari2600.ram[95][7] ),
    .A2(net4998),
    .A1(\atari2600.ram[92][7] ));
 sg13g2_a22oi_1 _17823_ (.Y(_09570_),
    .B1(net4823),
    .B2(\atari2600.ram[94][7] ),
    .A2(net4918),
    .A1(\atari2600.ram[93][7] ));
 sg13g2_a21oi_1 _17824_ (.A1(_09569_),
    .A2(_09570_),
    .Y(_09571_),
    .B1(net4957));
 sg13g2_a22oi_1 _17825_ (.Y(_09572_),
    .B1(net4847),
    .B2(\atari2600.ram[87][7] ),
    .A2(net4977),
    .A1(\atari2600.ram[84][7] ));
 sg13g2_a22oi_1 _17826_ (.Y(_09573_),
    .B1(net4803),
    .B2(\atari2600.ram[86][7] ),
    .A2(net4898),
    .A1(\atari2600.ram[85][7] ));
 sg13g2_a21oi_2 _17827_ (.B1(net5008),
    .Y(_09574_),
    .A2(_09573_),
    .A1(_09572_));
 sg13g2_a22oi_1 _17828_ (.Y(_09575_),
    .B1(net4850),
    .B2(\atari2600.ram[91][7] ),
    .A2(net4981),
    .A1(\atari2600.ram[88][7] ));
 sg13g2_a22oi_1 _17829_ (.Y(_09576_),
    .B1(net4804),
    .B2(\atari2600.ram[90][7] ),
    .A2(net4899),
    .A1(\atari2600.ram[89][7] ));
 sg13g2_a21oi_2 _17830_ (.B1(net4941),
    .Y(_09577_),
    .A2(_09576_),
    .A1(_09575_));
 sg13g2_a22oi_1 _17831_ (.Y(_09578_),
    .B1(net4863),
    .B2(\atari2600.ram[83][7] ),
    .A2(net4994),
    .A1(\atari2600.ram[80][7] ));
 sg13g2_a22oi_1 _17832_ (.Y(_09579_),
    .B1(net4820),
    .B2(\atari2600.ram[82][7] ),
    .A2(net4916),
    .A1(\atari2600.ram[81][7] ));
 sg13g2_a21oi_1 _17833_ (.A1(_09578_),
    .A2(_09579_),
    .Y(_09580_),
    .B1(net4933));
 sg13g2_nor4_2 _17834_ (.A(_09571_),
    .B(_09574_),
    .C(_09577_),
    .Y(_09581_),
    .D(_09580_));
 sg13g2_a22oi_1 _17835_ (.Y(_09582_),
    .B1(net4865),
    .B2(\atari2600.ram[127][7] ),
    .A2(net4994),
    .A1(\atari2600.ram[124][7] ));
 sg13g2_a22oi_1 _17836_ (.Y(_09583_),
    .B1(net4818),
    .B2(\atari2600.ram[126][7] ),
    .A2(net4913),
    .A1(\atari2600.ram[125][7] ));
 sg13g2_a21oi_2 _17837_ (.B1(net4958),
    .Y(_09584_),
    .A2(_09583_),
    .A1(_09582_));
 sg13g2_a22oi_1 _17838_ (.Y(_09585_),
    .B1(net4854),
    .B2(\atari2600.ram[115][7] ),
    .A2(net4984),
    .A1(\atari2600.ram[112][7] ));
 sg13g2_a22oi_1 _17839_ (.Y(_09586_),
    .B1(net4809),
    .B2(\atari2600.ram[114][7] ),
    .A2(net4903),
    .A1(\atari2600.ram[113][7] ));
 sg13g2_a21oi_2 _17840_ (.B1(net4930),
    .Y(_09587_),
    .A2(_09586_),
    .A1(_09585_));
 sg13g2_a22oi_1 _17841_ (.Y(_09588_),
    .B1(net4856),
    .B2(\atari2600.ram[123][7] ),
    .A2(net4987),
    .A1(\atari2600.ram[120][7] ));
 sg13g2_a22oi_1 _17842_ (.Y(_09589_),
    .B1(net4811),
    .B2(\atari2600.ram[122][7] ),
    .A2(net4905),
    .A1(\atari2600.ram[121][7] ));
 sg13g2_a21oi_1 _17843_ (.A1(_09588_),
    .A2(_09589_),
    .Y(_09590_),
    .B1(net4943));
 sg13g2_a22oi_1 _17844_ (.Y(_09591_),
    .B1(net4857),
    .B2(\atari2600.ram[119][7] ),
    .A2(net4986),
    .A1(\atari2600.ram[116][7] ));
 sg13g2_a22oi_1 _17845_ (.Y(_09592_),
    .B1(net4812),
    .B2(\atari2600.ram[118][7] ),
    .A2(net4907),
    .A1(\atari2600.ram[117][7] ));
 sg13g2_a21oi_1 _17846_ (.A1(_09591_),
    .A2(_09592_),
    .Y(_09593_),
    .B1(net5013));
 sg13g2_nor4_2 _17847_ (.A(_09584_),
    .B(_09587_),
    .C(_09590_),
    .Y(_09594_),
    .D(_09593_));
 sg13g2_nor2_1 _17848_ (.A(net4776),
    .B(_09594_),
    .Y(_09595_));
 sg13g2_o21ai_1 _17849_ (.B1(net5020),
    .Y(_09596_),
    .A1(net4774),
    .A2(_09581_));
 sg13g2_nor4_2 _17850_ (.A(_09554_),
    .B(_09568_),
    .C(_09595_),
    .Y(_09597_),
    .D(_09596_));
 sg13g2_a22oi_1 _17851_ (.Y(_09598_),
    .B1(net4840),
    .B2(\atari2600.ram[11][7] ),
    .A2(net4970),
    .A1(\atari2600.ram[8][7] ));
 sg13g2_a22oi_1 _17852_ (.Y(_09599_),
    .B1(net4795),
    .B2(\atari2600.ram[10][7] ),
    .A2(net4889),
    .A1(\atari2600.ram[9][7] ));
 sg13g2_a21oi_1 _17853_ (.A1(_09598_),
    .A2(_09599_),
    .Y(_09600_),
    .B1(net4938));
 sg13g2_a22oi_1 _17854_ (.Y(_09601_),
    .B1(net4834),
    .B2(\atari2600.ram[15][7] ),
    .A2(net4964),
    .A1(\atari2600.ram[12][7] ));
 sg13g2_a22oi_1 _17855_ (.Y(_09602_),
    .B1(net4790),
    .B2(\atari2600.ram[14][7] ),
    .A2(net4884),
    .A1(\atari2600.ram[13][7] ));
 sg13g2_a21oi_1 _17856_ (.A1(_09601_),
    .A2(_09602_),
    .Y(_09603_),
    .B1(net4950));
 sg13g2_a22oi_1 _17857_ (.Y(_09604_),
    .B1(net4844),
    .B2(\atari2600.ram[3][7] ),
    .A2(net4974),
    .A1(\atari2600.ram[0][7] ));
 sg13g2_a22oi_1 _17858_ (.Y(_09605_),
    .B1(net4798),
    .B2(\atari2600.ram[2][7] ),
    .A2(net4892),
    .A1(\atari2600.ram[1][7] ));
 sg13g2_a21oi_1 _17859_ (.A1(_09604_),
    .A2(_09605_),
    .Y(_09606_),
    .B1(net4927));
 sg13g2_a22oi_1 _17860_ (.Y(_09607_),
    .B1(net4843),
    .B2(\atari2600.ram[7][7] ),
    .A2(net4973),
    .A1(\atari2600.ram[4][7] ));
 sg13g2_a22oi_1 _17861_ (.Y(_09608_),
    .B1(net4799),
    .B2(\atari2600.ram[6][7] ),
    .A2(net4893),
    .A1(\atari2600.ram[5][7] ));
 sg13g2_a21oi_2 _17862_ (.B1(net5007),
    .Y(_09609_),
    .A2(_09608_),
    .A1(_09607_));
 sg13g2_nor4_1 _17863_ (.A(_09600_),
    .B(_09603_),
    .C(_09606_),
    .D(_09609_),
    .Y(_09610_));
 sg13g2_nor2_1 _17864_ (.A(net4777),
    .B(_09610_),
    .Y(_09611_));
 sg13g2_a22oi_1 _17865_ (.Y(_09612_),
    .B1(net4841),
    .B2(\atari2600.ram[51][7] ),
    .A2(net4972),
    .A1(\atari2600.ram[48][7] ));
 sg13g2_a22oi_1 _17866_ (.Y(_09613_),
    .B1(net4794),
    .B2(\atari2600.ram[50][7] ),
    .A2(net4888),
    .A1(\atari2600.ram[49][7] ));
 sg13g2_a21oi_2 _17867_ (.B1(net4926),
    .Y(_09614_),
    .A2(_09613_),
    .A1(_09612_));
 sg13g2_a22oi_1 _17868_ (.Y(_09615_),
    .B1(net4838),
    .B2(\atari2600.ram[59][7] ),
    .A2(net4968),
    .A1(\atari2600.ram[56][7] ));
 sg13g2_a22oi_1 _17869_ (.Y(_09616_),
    .B1(net4792),
    .B2(\atari2600.ram[58][7] ),
    .A2(net4886),
    .A1(\atari2600.ram[57][7] ));
 sg13g2_a21oi_1 _17870_ (.A1(_09615_),
    .A2(_09616_),
    .Y(_09617_),
    .B1(net4940));
 sg13g2_a22oi_1 _17871_ (.Y(_09618_),
    .B1(net4853),
    .B2(\atari2600.ram[55][7] ),
    .A2(net4983),
    .A1(\atari2600.ram[52][7] ));
 sg13g2_a22oi_1 _17872_ (.Y(_09619_),
    .B1(net4808),
    .B2(\atari2600.ram[54][7] ),
    .A2(net4902),
    .A1(\atari2600.ram[53][7] ));
 sg13g2_a21oi_2 _17873_ (.B1(net5012),
    .Y(_09620_),
    .A2(_09619_),
    .A1(_09618_));
 sg13g2_a22oi_1 _17874_ (.Y(_09621_),
    .B1(net4838),
    .B2(\atari2600.ram[63][7] ),
    .A2(net4968),
    .A1(\atari2600.ram[60][7] ));
 sg13g2_a22oi_1 _17875_ (.Y(_09622_),
    .B1(net4792),
    .B2(\atari2600.ram[62][7] ),
    .A2(net4886),
    .A1(\atari2600.ram[61][7] ));
 sg13g2_a21oi_1 _17876_ (.A1(_09621_),
    .A2(_09622_),
    .Y(_09623_),
    .B1(net4951));
 sg13g2_nor4_2 _17877_ (.A(_09614_),
    .B(_09617_),
    .C(_09620_),
    .Y(_09624_),
    .D(_09623_));
 sg13g2_nor2_1 _17878_ (.A(net4776),
    .B(_09624_),
    .Y(_09625_));
 sg13g2_a22oi_1 _17879_ (.Y(_09626_),
    .B1(net4832),
    .B2(\atari2600.ram[35][7] ),
    .A2(net4962),
    .A1(\atari2600.ram[32][7] ));
 sg13g2_a22oi_1 _17880_ (.Y(_09627_),
    .B1(net4787),
    .B2(\atari2600.ram[34][7] ),
    .A2(net4881),
    .A1(\atari2600.ram[33][7] ));
 sg13g2_a21oi_1 _17881_ (.A1(_09626_),
    .A2(_09627_),
    .Y(_09628_),
    .B1(net4925));
 sg13g2_a22oi_1 _17882_ (.Y(_09629_),
    .B1(net4830),
    .B2(\atari2600.ram[39][7] ),
    .A2(net4960),
    .A1(\atari2600.ram[36][7] ));
 sg13g2_a22oi_1 _17883_ (.Y(_09630_),
    .B1(net4785),
    .B2(\atari2600.ram[38][7] ),
    .A2(net4880),
    .A1(\atari2600.ram[37][7] ));
 sg13g2_a21oi_2 _17884_ (.B1(net5006),
    .Y(_09631_),
    .A2(_09630_),
    .A1(_09629_));
 sg13g2_a22oi_1 _17885_ (.Y(_09632_),
    .B1(net4831),
    .B2(\atari2600.ram[47][7] ),
    .A2(net4961),
    .A1(\atari2600.ram[44][7] ));
 sg13g2_a22oi_1 _17886_ (.Y(_09633_),
    .B1(net4785),
    .B2(\atari2600.ram[46][7] ),
    .A2(net4880),
    .A1(\atari2600.ram[45][7] ));
 sg13g2_a21oi_2 _17887_ (.B1(net4949),
    .Y(_09634_),
    .A2(_09633_),
    .A1(_09632_));
 sg13g2_a22oi_1 _17888_ (.Y(_09635_),
    .B1(net4833),
    .B2(\atari2600.ram[43][7] ),
    .A2(net4963),
    .A1(\atari2600.ram[40][7] ));
 sg13g2_a22oi_1 _17889_ (.Y(_09636_),
    .B1(net4788),
    .B2(\atari2600.ram[42][7] ),
    .A2(net4882),
    .A1(\atari2600.ram[41][7] ));
 sg13g2_a21oi_1 _17890_ (.A1(_09635_),
    .A2(_09636_),
    .Y(_09637_),
    .B1(net4937));
 sg13g2_nor4_2 _17891_ (.A(_09628_),
    .B(_09631_),
    .C(_09634_),
    .Y(_09638_),
    .D(_09637_));
 sg13g2_nor2_1 _17892_ (.A(net4772),
    .B(_09638_),
    .Y(_09639_));
 sg13g2_a22oi_1 _17893_ (.Y(_09640_),
    .B1(net4846),
    .B2(\atari2600.ram[31][7] ),
    .A2(net4976),
    .A1(\atari2600.ram[28][7] ));
 sg13g2_a22oi_1 _17894_ (.Y(_09641_),
    .B1(net4801),
    .B2(\atari2600.ram[30][7] ),
    .A2(net4896),
    .A1(\atari2600.ram[29][7] ));
 sg13g2_a21oi_1 _17895_ (.A1(_09640_),
    .A2(_09641_),
    .Y(_09642_),
    .B1(net4953));
 sg13g2_a22oi_1 _17896_ (.Y(_09643_),
    .B1(net4846),
    .B2(\atari2600.ram[23][7] ),
    .A2(net4976),
    .A1(\atari2600.ram[20][7] ));
 sg13g2_a22oi_1 _17897_ (.Y(_09644_),
    .B1(net4801),
    .B2(\atari2600.ram[22][7] ),
    .A2(net4896),
    .A1(\atari2600.ram[21][7] ));
 sg13g2_a21oi_1 _17898_ (.A1(_09643_),
    .A2(_09644_),
    .Y(_09645_),
    .B1(net5008));
 sg13g2_a22oi_1 _17899_ (.Y(_09646_),
    .B1(net4841),
    .B2(\atari2600.ram[27][7] ),
    .A2(net4971),
    .A1(\atari2600.ram[24][7] ));
 sg13g2_a22oi_1 _17900_ (.Y(_09647_),
    .B1(net4794),
    .B2(\atari2600.ram[26][7] ),
    .A2(net4888),
    .A1(\atari2600.ram[25][7] ));
 sg13g2_a21oi_2 _17901_ (.B1(net4940),
    .Y(_09648_),
    .A2(_09647_),
    .A1(_09646_));
 sg13g2_a22oi_1 _17902_ (.Y(_09649_),
    .B1(net4849),
    .B2(\atari2600.ram[19][7] ),
    .A2(net4980),
    .A1(\atari2600.ram[16][7] ));
 sg13g2_a22oi_1 _17903_ (.Y(_09650_),
    .B1(net4805),
    .B2(\atari2600.ram[18][7] ),
    .A2(net4897),
    .A1(\atari2600.ram[17][7] ));
 sg13g2_a21oi_2 _17904_ (.B1(net4929),
    .Y(_09651_),
    .A2(_09650_),
    .A1(_09649_));
 sg13g2_nor4_2 _17905_ (.A(_09642_),
    .B(_09645_),
    .C(_09648_),
    .Y(_09652_),
    .D(_09651_));
 sg13g2_o21ai_1 _17906_ (.B1(net5023),
    .Y(_09653_),
    .A1(net4773),
    .A2(_09652_));
 sg13g2_nor4_1 _17907_ (.A(_09611_),
    .B(_09625_),
    .C(_09639_),
    .D(_09653_),
    .Y(_09654_));
 sg13g2_nor2_2 _17908_ (.A(_09597_),
    .B(_09654_),
    .Y(_00008_));
 sg13g2_nor2_1 _17909_ (.A(\atari2600.clk_counter[1] ),
    .B(net7122),
    .Y(_09655_));
 sg13g2_nand4_1 _17910_ (.B(_08131_),
    .C(_08132_),
    .A(_00142_),
    .Y(_09656_),
    .D(_09655_));
 sg13g2_o21ai_1 _17911_ (.B1(_09656_),
    .Y(_09657_),
    .A1(_07923_),
    .A2(_08133_));
 sg13g2_nand2_2 _17912_ (.Y(_09658_),
    .A(_08669_),
    .B(_09657_));
 sg13g2_inv_2 _17913_ (.Y(_09659_),
    .A(_09658_));
 sg13g2_a21oi_1 _17914_ (.A1(net7379),
    .A2(_09659_),
    .Y(_09660_),
    .B1(net5988));
 sg13g2_nand2_1 _17915_ (.Y(_09661_),
    .A(net3014),
    .B(net5197));
 sg13g2_nand2b_1 _17916_ (.Y(_09662_),
    .B(net5825),
    .A_N(\atari2600.tia.diag[57] ));
 sg13g2_nor2b_1 _17917_ (.A(net5825),
    .B_N(\atari2600.tia.diag[57] ),
    .Y(_09663_));
 sg13g2_xor2_1 _17918_ (.B(net5825),
    .A(\atari2600.tia.diag[57] ),
    .X(_09664_));
 sg13g2_nor2b_1 _17919_ (.A(net5829),
    .B_N(\atari2600.tia.diag[56] ),
    .Y(_09665_));
 sg13g2_o21ai_1 _17920_ (.B1(_09662_),
    .Y(_09666_),
    .A1(_09664_),
    .A2(_09665_));
 sg13g2_nor2_1 _17921_ (.A(\atari2600.tia.diag[58] ),
    .B(net5561),
    .Y(_09667_));
 sg13g2_nand2_1 _17922_ (.Y(_09668_),
    .A(\atari2600.tia.diag[58] ),
    .B(net5561));
 sg13g2_nand2b_1 _17923_ (.Y(_09669_),
    .B(_09668_),
    .A_N(_09667_));
 sg13g2_xnor2_1 _17924_ (.Y(_09670_),
    .A(_09666_),
    .B(_09669_));
 sg13g2_xor2_1 _17925_ (.B(net5820),
    .A(net5592),
    .X(_09671_));
 sg13g2_a21oi_2 _17926_ (.B1(_09667_),
    .Y(_09672_),
    .A2(_09668_),
    .A1(_09666_));
 sg13g2_nor2_1 _17927_ (.A(_09671_),
    .B(_09672_),
    .Y(_09673_));
 sg13g2_xnor2_1 _17928_ (.Y(_09674_),
    .A(_09671_),
    .B(_09672_));
 sg13g2_nor2_1 _17929_ (.A(net5837),
    .B(_09670_),
    .Y(_09675_));
 sg13g2_a21oi_1 _17930_ (.A1(net5837),
    .A2(_09674_),
    .Y(_09676_),
    .B1(_09675_));
 sg13g2_nor2_1 _17931_ (.A(net5590),
    .B(net5560),
    .Y(_09677_));
 sg13g2_xnor2_1 _17932_ (.Y(_09678_),
    .A(net5590),
    .B(net5818));
 sg13g2_a21oi_2 _17933_ (.B1(_09673_),
    .Y(_09679_),
    .A2(net5820),
    .A1(_07994_));
 sg13g2_inv_1 _17934_ (.Y(_09680_),
    .A(_09679_));
 sg13g2_xnor2_1 _17935_ (.Y(_09681_),
    .A(_09678_),
    .B(_09679_));
 sg13g2_xor2_1 _17936_ (.B(net5812),
    .A(\atari2600.tia.diag[61] ),
    .X(_09682_));
 sg13g2_a21oi_2 _17937_ (.B1(_09677_),
    .Y(_09683_),
    .A2(_09680_),
    .A1(_09678_));
 sg13g2_nor2_1 _17938_ (.A(_09682_),
    .B(_09683_),
    .Y(_09684_));
 sg13g2_xnor2_1 _17939_ (.Y(_09685_),
    .A(_09682_),
    .B(_09683_));
 sg13g2_nand2_1 _17940_ (.Y(_09686_),
    .A(net5838),
    .B(_09685_));
 sg13g2_o21ai_1 _17941_ (.B1(_09686_),
    .Y(_09687_),
    .A1(net5838),
    .A2(_09681_));
 sg13g2_nor2_1 _17942_ (.A(net5836),
    .B(_09676_),
    .Y(_09688_));
 sg13g2_a21oi_2 _17943_ (.B1(_09688_),
    .Y(_09689_),
    .A2(_09687_),
    .A1(net5836));
 sg13g2_xor2_1 _17944_ (.B(_09689_),
    .A(_00159_),
    .X(_09690_));
 sg13g2_xnor2_1 _17945_ (.Y(_09691_),
    .A(_09664_),
    .B(_09665_));
 sg13g2_nor2_1 _17946_ (.A(net5837),
    .B(_09674_),
    .Y(_09692_));
 sg13g2_a21oi_1 _17947_ (.A1(net5838),
    .A2(_09681_),
    .Y(_09693_),
    .B1(_09692_));
 sg13g2_or2_1 _17948_ (.X(_09694_),
    .B(_09691_),
    .A(net5837));
 sg13g2_a21oi_1 _17949_ (.A1(net5837),
    .A2(_09670_),
    .Y(_09695_),
    .B1(net5836));
 sg13g2_a22oi_1 _17950_ (.Y(_09696_),
    .B1(_09694_),
    .B2(_09695_),
    .A2(_09693_),
    .A1(net5836));
 sg13g2_xnor2_1 _17951_ (.Y(_09697_),
    .A(_00159_),
    .B(_09696_));
 sg13g2_nand2b_1 _17952_ (.Y(_09698_),
    .B(net5829),
    .A_N(\atari2600.tia.diag[56] ));
 sg13g2_nand2b_1 _17953_ (.Y(_09699_),
    .B(_09698_),
    .A_N(_09665_));
 sg13g2_or2_1 _17954_ (.X(_09700_),
    .B(_09699_),
    .A(net5837));
 sg13g2_a21oi_1 _17955_ (.A1(net5837),
    .A2(_09691_),
    .Y(_09701_),
    .B1(net5836));
 sg13g2_a22oi_1 _17956_ (.Y(_09702_),
    .B1(_09700_),
    .B2(_09701_),
    .A2(_09676_),
    .A1(net5836));
 sg13g2_xnor2_1 _17957_ (.Y(_09703_),
    .A(_00159_),
    .B(_09702_));
 sg13g2_mux4_1 _17958_ (.S0(_09697_),
    .A0(\atari2600.tia.diag[98] ),
    .A1(\atari2600.tia.diag[96] ),
    .A2(\atari2600.tia.old_grp1[2] ),
    .A3(\atari2600.tia.old_grp1[0] ),
    .S1(\atari2600.tia.vdelp1 ),
    .X(_09704_));
 sg13g2_mux4_1 _17959_ (.S0(_09697_),
    .A0(\atari2600.tia.diag[99] ),
    .A1(\atari2600.tia.diag[97] ),
    .A2(\atari2600.tia.old_grp1[3] ),
    .A3(\atari2600.tia.old_grp1[1] ),
    .S1(\atari2600.tia.vdelp1 ),
    .X(_09705_));
 sg13g2_mux2_1 _17960_ (.A0(_09704_),
    .A1(_09705_),
    .S(_09703_),
    .X(_09706_));
 sg13g2_nor2_1 _17961_ (.A(_09690_),
    .B(_09706_),
    .Y(_09707_));
 sg13g2_mux4_1 _17962_ (.S0(_09697_),
    .A0(\atari2600.tia.diag[102] ),
    .A1(\atari2600.tia.diag[100] ),
    .A2(\atari2600.tia.old_grp1[6] ),
    .A3(\atari2600.tia.old_grp1[4] ),
    .S1(\atari2600.tia.vdelp1 ),
    .X(_09708_));
 sg13g2_mux4_1 _17963_ (.S0(_09697_),
    .A0(\atari2600.tia.diag[103] ),
    .A1(\atari2600.tia.diag[101] ),
    .A2(\atari2600.tia.old_grp1[7] ),
    .A3(\atari2600.tia.old_grp1[5] ),
    .S1(\atari2600.tia.vdelp1 ),
    .X(_09709_));
 sg13g2_mux2_1 _17964_ (.A0(_09708_),
    .A1(_09709_),
    .S(_09703_),
    .X(_09710_));
 sg13g2_nor2b_1 _17965_ (.A(_09710_),
    .B_N(_09690_),
    .Y(_09711_));
 sg13g2_xnor2_1 _17966_ (.Y(_09712_),
    .A(\atari2600.tia.diag[63] ),
    .B(net5800));
 sg13g2_nor2_1 _17967_ (.A(net5589),
    .B(net5558),
    .Y(_09713_));
 sg13g2_xnor2_1 _17968_ (.Y(_09714_),
    .A(net5589),
    .B(net5804));
 sg13g2_a21oi_1 _17969_ (.A1(_07993_),
    .A2(net5812),
    .Y(_09715_),
    .B1(_09684_));
 sg13g2_nor2b_1 _17970_ (.A(_09715_),
    .B_N(_09714_),
    .Y(_09716_));
 sg13g2_o21ai_1 _17971_ (.B1(_09712_),
    .Y(_09717_),
    .A1(_09713_),
    .A2(_09716_));
 sg13g2_o21ai_1 _17972_ (.B1(_09717_),
    .Y(_09718_),
    .A1(\atari2600.tia.diag[63] ),
    .A2(net5557));
 sg13g2_nand2_1 _17973_ (.Y(_09719_),
    .A(\atari2600.tia.diag[61] ),
    .B(\atari2600.tia.p1_w[5] ));
 sg13g2_xor2_1 _17974_ (.B(\atari2600.tia.p1_w[5] ),
    .A(\atari2600.tia.diag[61] ),
    .X(_09720_));
 sg13g2_nand2_1 _17975_ (.Y(_09721_),
    .A(net5591),
    .B(\atari2600.tia.p1_w[4] ));
 sg13g2_nand2_1 _17976_ (.Y(_09722_),
    .A(\atari2600.tia.diag[59] ),
    .B(\atari2600.tia.p1_w[3] ));
 sg13g2_nor2_1 _17977_ (.A(net5591),
    .B(\atari2600.tia.p1_w[4] ),
    .Y(_09723_));
 sg13g2_xor2_1 _17978_ (.B(\atari2600.tia.p1_w[4] ),
    .A(net5591),
    .X(_09724_));
 sg13g2_o21ai_1 _17979_ (.B1(_09721_),
    .Y(_09725_),
    .A1(_09722_),
    .A2(_09723_));
 sg13g2_nand2_1 _17980_ (.Y(_09726_),
    .A(_09720_),
    .B(_09725_));
 sg13g2_nand2_1 _17981_ (.Y(_09727_),
    .A(_09719_),
    .B(_09726_));
 sg13g2_xnor2_1 _17982_ (.Y(_09728_),
    .A(net5589),
    .B(_09727_));
 sg13g2_inv_1 _17983_ (.Y(_09729_),
    .A(_09728_));
 sg13g2_nand2_1 _17984_ (.Y(_09730_),
    .A(net5806),
    .B(_09728_));
 sg13g2_xnor2_1 _17985_ (.Y(_09731_),
    .A(_09720_),
    .B(_09725_));
 sg13g2_xor2_1 _17986_ (.B(\atari2600.tia.p1_w[3] ),
    .A(net5592),
    .X(_09732_));
 sg13g2_a21o_1 _17987_ (.A2(_09732_),
    .A1(_00152_),
    .B1(_09672_),
    .X(_09733_));
 sg13g2_o21ai_1 _17988_ (.B1(_09733_),
    .Y(_09734_),
    .A1(net5819),
    .A2(_09732_));
 sg13g2_xnor2_1 _17989_ (.Y(_09735_),
    .A(_09722_),
    .B(_09724_));
 sg13g2_nor2_1 _17990_ (.A(net5814),
    .B(_09735_),
    .Y(_09736_));
 sg13g2_nor2_1 _17991_ (.A(_09734_),
    .B(_09736_),
    .Y(_09737_));
 sg13g2_and2_1 _17992_ (.A(net5814),
    .B(_09735_),
    .X(_09738_));
 sg13g2_nor2_1 _17993_ (.A(_09737_),
    .B(_09738_),
    .Y(_09739_));
 sg13g2_xnor2_1 _17994_ (.Y(_09740_),
    .A(net5809),
    .B(_09731_));
 sg13g2_a22oi_1 _17995_ (.Y(_09741_),
    .B1(_09739_),
    .B2(_09740_),
    .A2(_09731_),
    .A1(net5811));
 sg13g2_xor2_1 _17996_ (.B(_09728_),
    .A(net5803),
    .X(_09742_));
 sg13g2_o21ai_1 _17997_ (.B1(_09730_),
    .Y(_09743_),
    .A1(_09741_),
    .A2(_09742_));
 sg13g2_nand3_1 _17998_ (.B(_09720_),
    .C(_09725_),
    .A(net5589),
    .Y(_09744_));
 sg13g2_o21ai_1 _17999_ (.B1(_09744_),
    .Y(_09745_),
    .A1(_00155_),
    .A2(_09719_));
 sg13g2_xnor2_1 _18000_ (.Y(_09746_),
    .A(\atari2600.tia.diag[63] ),
    .B(_09745_));
 sg13g2_xor2_1 _18001_ (.B(_09745_),
    .A(_09712_),
    .X(_09747_));
 sg13g2_a22oi_1 _18002_ (.Y(_09748_),
    .B1(_09747_),
    .B2(_09743_),
    .A2(_09746_),
    .A1(_08124_));
 sg13g2_and2_1 _18003_ (.A(_09718_),
    .B(_09748_),
    .X(_09749_));
 sg13g2_nor2_1 _18004_ (.A(\atari2600.tia.p1_spacing[6] ),
    .B(net5558),
    .Y(_09750_));
 sg13g2_nand2_1 _18005_ (.Y(_09751_),
    .A(\atari2600.tia.p1_spacing[4] ),
    .B(net5560));
 sg13g2_xnor2_1 _18006_ (.Y(_09752_),
    .A(\atari2600.tia.p1_spacing[5] ),
    .B(net5811));
 sg13g2_nand2_1 _18007_ (.Y(_09753_),
    .A(_09751_),
    .B(_09752_));
 sg13g2_o21ai_1 _18008_ (.B1(_09753_),
    .Y(_09754_),
    .A1(\atari2600.tia.p1_spacing[5] ),
    .A2(net5559));
 sg13g2_xnor2_1 _18009_ (.Y(_09755_),
    .A(\atari2600.tia.p1_spacing[6] ),
    .B(net5805));
 sg13g2_a21oi_1 _18010_ (.A1(_09754_),
    .A2(_09755_),
    .Y(_09756_),
    .B1(_09750_));
 sg13g2_xnor2_1 _18011_ (.Y(_09757_),
    .A(_00150_),
    .B(_09756_));
 sg13g2_nand2_1 _18012_ (.Y(_09758_),
    .A(_00158_),
    .B(_09757_));
 sg13g2_xnor2_1 _18013_ (.Y(_09759_),
    .A(_09754_),
    .B(_09755_));
 sg13g2_inv_1 _18014_ (.Y(_09760_),
    .A(_09759_));
 sg13g2_nor2_1 _18015_ (.A(net5589),
    .B(_09759_),
    .Y(_09761_));
 sg13g2_xor2_1 _18016_ (.B(_09752_),
    .A(_09751_),
    .X(_09762_));
 sg13g2_xnor2_1 _18017_ (.Y(_09763_),
    .A(\atari2600.tia.p1_spacing[4] ),
    .B(net5816));
 sg13g2_o21ai_1 _18018_ (.B1(_09679_),
    .Y(_09764_),
    .A1(net5590),
    .A2(_09763_));
 sg13g2_nand2_1 _18019_ (.Y(_09765_),
    .A(net5591),
    .B(_09763_));
 sg13g2_o21ai_1 _18020_ (.B1(_09765_),
    .Y(_09766_),
    .A1(_00157_),
    .A2(_09762_));
 sg13g2_a21oi_1 _18021_ (.A1(_00157_),
    .A2(_09762_),
    .Y(_09767_),
    .B1(_09766_));
 sg13g2_a22oi_1 _18022_ (.Y(_09768_),
    .B1(_09764_),
    .B2(_09767_),
    .A2(_09762_),
    .A1(_07993_));
 sg13g2_xor2_1 _18023_ (.B(_09759_),
    .A(_00155_),
    .X(_09769_));
 sg13g2_nor2_1 _18024_ (.A(_09768_),
    .B(_09769_),
    .Y(_09770_));
 sg13g2_xnor2_1 _18025_ (.Y(_09771_),
    .A(\atari2600.tia.diag[63] ),
    .B(_09757_));
 sg13g2_o21ai_1 _18026_ (.B1(_09771_),
    .Y(_09772_),
    .A1(_09761_),
    .A2(_09770_));
 sg13g2_nor2_1 _18027_ (.A(_09731_),
    .B(_09762_),
    .Y(_09773_));
 sg13g2_nor2_1 _18028_ (.A(_09735_),
    .B(_09763_),
    .Y(_09774_));
 sg13g2_a21oi_1 _18029_ (.A1(_09735_),
    .A2(_09763_),
    .Y(_09775_),
    .B1(_09773_));
 sg13g2_o21ai_1 _18030_ (.B1(_09775_),
    .Y(_09776_),
    .A1(_09734_),
    .A2(_09774_));
 sg13g2_a22oi_1 _18031_ (.Y(_09777_),
    .B1(_09762_),
    .B2(_09731_),
    .A2(_09760_),
    .A1(_09728_));
 sg13g2_a22oi_1 _18032_ (.Y(_09778_),
    .B1(_09776_),
    .B2(_09777_),
    .A2(_09759_),
    .A1(_09729_));
 sg13g2_o21ai_1 _18033_ (.B1(_09778_),
    .Y(_09779_),
    .A1(_09746_),
    .A2(_09757_));
 sg13g2_o21ai_1 _18034_ (.B1(_09779_),
    .Y(_09780_),
    .A1(\atari2600.tia.p1_copies[2] ),
    .A2(\atari2600.tia.p1_copies[1] ));
 sg13g2_a221oi_1 _18035_ (.B2(_09772_),
    .C1(_09780_),
    .B1(_09758_),
    .A1(_09746_),
    .Y(_09781_),
    .A2(_09757_));
 sg13g2_nand2b_1 _18036_ (.Y(_09782_),
    .B(net5806),
    .A_N(\atari2600.tia.p1_spacing[5] ));
 sg13g2_xor2_1 _18037_ (.B(net5806),
    .A(\atari2600.tia.p1_spacing[5] ),
    .X(_09783_));
 sg13g2_nor2_1 _18038_ (.A(_07920_),
    .B(net5811),
    .Y(_09784_));
 sg13g2_o21ai_1 _18039_ (.B1(_09782_),
    .Y(_09785_),
    .A1(_09783_),
    .A2(_09784_));
 sg13g2_xor2_1 _18040_ (.B(net5800),
    .A(\atari2600.tia.p1_spacing[6] ),
    .X(_09786_));
 sg13g2_xnor2_1 _18041_ (.Y(_09787_),
    .A(_09785_),
    .B(_09786_));
 sg13g2_nand2_1 _18042_ (.Y(_09788_),
    .A(_00158_),
    .B(_09787_));
 sg13g2_xor2_1 _18043_ (.B(_09784_),
    .A(_09783_),
    .X(_09789_));
 sg13g2_xnor2_1 _18044_ (.Y(_09790_),
    .A(_09783_),
    .B(_09784_));
 sg13g2_xor2_1 _18045_ (.B(net5811),
    .A(\atari2600.tia.p1_spacing[4] ),
    .X(_09791_));
 sg13g2_nand2_1 _18046_ (.Y(_09792_),
    .A(_00157_),
    .B(_09791_));
 sg13g2_xnor2_1 _18047_ (.Y(_09793_),
    .A(_07993_),
    .B(_09791_));
 sg13g2_o21ai_1 _18048_ (.B1(_09792_),
    .Y(_09794_),
    .A1(_09683_),
    .A2(_09793_));
 sg13g2_xnor2_1 _18049_ (.Y(_09795_),
    .A(_00155_),
    .B(_09790_));
 sg13g2_a22oi_1 _18050_ (.Y(_09796_),
    .B1(_09794_),
    .B2(_09795_),
    .A2(_09789_),
    .A1(_07992_));
 sg13g2_xor2_1 _18051_ (.B(_09787_),
    .A(\atari2600.tia.diag[63] ),
    .X(_09797_));
 sg13g2_o21ai_1 _18052_ (.B1(_09788_),
    .Y(_09798_),
    .A1(_09796_),
    .A2(_09797_));
 sg13g2_xnor2_1 _18053_ (.Y(_09799_),
    .A(net5819),
    .B(_09732_));
 sg13g2_a221oi_1 _18054_ (.B2(_09698_),
    .C1(_09663_),
    .B1(_09662_),
    .A1(\atari2600.tia.diag[58] ),
    .Y(_09800_),
    .A2(net5561));
 sg13g2_nor3_1 _18055_ (.A(_09667_),
    .B(_09799_),
    .C(_09800_),
    .Y(_09801_));
 sg13g2_a21oi_1 _18056_ (.A1(net5563),
    .A2(_09732_),
    .Y(_09802_),
    .B1(_09801_));
 sg13g2_nor4_2 _18057_ (.A(_09664_),
    .B(_09669_),
    .C(_09699_),
    .Y(_09803_),
    .D(_09799_));
 sg13g2_nor3_1 _18058_ (.A(_09736_),
    .B(_09802_),
    .C(_09803_),
    .Y(_09804_));
 sg13g2_nor2_1 _18059_ (.A(_09731_),
    .B(_09791_),
    .Y(_09805_));
 sg13g2_nor3_1 _18060_ (.A(_09738_),
    .B(_09804_),
    .C(_09805_),
    .Y(_09806_));
 sg13g2_a221oi_1 _18061_ (.B2(_09731_),
    .C1(_09806_),
    .B1(_09791_),
    .A1(_09728_),
    .Y(_09807_),
    .A2(_09789_));
 sg13g2_a21oi_1 _18062_ (.A1(_09729_),
    .A2(_09790_),
    .Y(_09808_),
    .B1(_09807_));
 sg13g2_o21ai_1 _18063_ (.B1(_09808_),
    .Y(_09809_),
    .A1(_09746_),
    .A2(_09787_));
 sg13g2_nand3_1 _18064_ (.B(_09798_),
    .C(_09809_),
    .A(\atari2600.tia.p1_copies[1] ),
    .Y(_09810_));
 sg13g2_a21oi_1 _18065_ (.A1(_09746_),
    .A2(_09787_),
    .Y(_09811_),
    .B1(_09810_));
 sg13g2_nor3_2 _18066_ (.A(_09749_),
    .B(_09781_),
    .C(_09811_),
    .Y(_09812_));
 sg13g2_or3_1 _18067_ (.A(_09712_),
    .B(_09713_),
    .C(_09716_),
    .X(_09813_));
 sg13g2_nand3_1 _18068_ (.B(_09717_),
    .C(_09813_),
    .A(net5838),
    .Y(_09814_));
 sg13g2_xnor2_1 _18069_ (.Y(_09815_),
    .A(_09714_),
    .B(_09715_));
 sg13g2_o21ai_1 _18070_ (.B1(net5836),
    .Y(_09816_),
    .A1(net5838),
    .A2(_09685_));
 sg13g2_nor2_1 _18071_ (.A(_09815_),
    .B(_09816_),
    .Y(_09817_));
 sg13g2_nor2b_1 _18072_ (.A(net5836),
    .B_N(_09693_),
    .Y(_09818_));
 sg13g2_a22oi_1 _18073_ (.Y(_09819_),
    .B1(_09818_),
    .B2(_09687_),
    .A2(_09817_),
    .A1(_09814_));
 sg13g2_or4_2 _18074_ (.A(_09707_),
    .B(_09711_),
    .C(_09812_),
    .D(_09819_),
    .X(_09820_));
 sg13g2_inv_1 _18075_ (.Y(_09821_),
    .A(net4770));
 sg13g2_nor2_1 _18076_ (.A(\atari2600.tia.vid_ypos[3] ),
    .B(_08137_),
    .Y(_09822_));
 sg13g2_nor2_1 _18077_ (.A(\atari2600.tia.vid_ypos[5] ),
    .B(\atari2600.tia.vid_ypos[4] ),
    .Y(_09823_));
 sg13g2_nand3_1 _18078_ (.B(_08139_),
    .C(_09823_),
    .A(_00144_),
    .Y(_09824_));
 sg13g2_o21ai_1 _18079_ (.B1(\atari2600.tia.vid_ypos[8] ),
    .Y(_09825_),
    .A1(_09822_),
    .A2(_09824_));
 sg13g2_nor2b_2 _18080_ (.A(_09658_),
    .B_N(_09825_),
    .Y(_09826_));
 sg13g2_nand2_2 _18081_ (.Y(_09827_),
    .A(_09659_),
    .B(_09825_));
 sg13g2_xor2_1 _18082_ (.B(net5820),
    .A(net5595),
    .X(_09828_));
 sg13g2_nor2_1 _18083_ (.A(net5596),
    .B(net5561),
    .Y(_09829_));
 sg13g2_xor2_1 _18084_ (.B(net5823),
    .A(net5596),
    .X(_09830_));
 sg13g2_nand2_1 _18085_ (.Y(_09831_),
    .A(_07999_),
    .B(net5825));
 sg13g2_nor2_1 _18086_ (.A(_07999_),
    .B(net5825),
    .Y(_09832_));
 sg13g2_xor2_1 _18087_ (.B(net5825),
    .A(\atari2600.tia.diag[65] ),
    .X(_09833_));
 sg13g2_nor2b_1 _18088_ (.A(net5829),
    .B_N(\atari2600.tia.diag[64] ),
    .Y(_09834_));
 sg13g2_nor2_1 _18089_ (.A(_09833_),
    .B(_09834_),
    .Y(_09835_));
 sg13g2_a21oi_1 _18090_ (.A1(_07999_),
    .A2(net5825),
    .Y(_09836_),
    .B1(_09835_));
 sg13g2_nor2_1 _18091_ (.A(_09830_),
    .B(_09836_),
    .Y(_09837_));
 sg13g2_nor2_2 _18092_ (.A(_09829_),
    .B(_09837_),
    .Y(_09838_));
 sg13g2_nor2_1 _18093_ (.A(_09828_),
    .B(_09838_),
    .Y(_09839_));
 sg13g2_a21oi_2 _18094_ (.B1(_09839_),
    .Y(_09840_),
    .A2(net5820),
    .A1(_07998_));
 sg13g2_xnor2_1 _18095_ (.Y(_09841_),
    .A(\atari2600.tia.diag[68] ),
    .B(net5818));
 sg13g2_nor2b_1 _18096_ (.A(_09840_),
    .B_N(_09841_),
    .Y(_09842_));
 sg13g2_xnor2_1 _18097_ (.Y(_09843_),
    .A(_09840_),
    .B(_09841_));
 sg13g2_a21oi_2 _18098_ (.B1(_09842_),
    .Y(_09844_),
    .A2(net5818),
    .A1(_07997_));
 sg13g2_xnor2_1 _18099_ (.Y(_09845_),
    .A(net5593),
    .B(net5810));
 sg13g2_nor2b_1 _18100_ (.A(_09844_),
    .B_N(_09845_),
    .Y(_09846_));
 sg13g2_xor2_1 _18101_ (.B(_09845_),
    .A(_09844_),
    .X(_09847_));
 sg13g2_nor2_1 _18102_ (.A(_08037_),
    .B(_09847_),
    .Y(_09848_));
 sg13g2_a21oi_1 _18103_ (.A1(_08037_),
    .A2(_09843_),
    .Y(_09849_),
    .B1(_09848_));
 sg13g2_xnor2_1 _18104_ (.Y(_09850_),
    .A(_09830_),
    .B(_09836_));
 sg13g2_inv_1 _18105_ (.Y(_09851_),
    .A(_09850_));
 sg13g2_xor2_1 _18106_ (.B(_09838_),
    .A(_09828_),
    .X(_09852_));
 sg13g2_nand2_1 _18107_ (.Y(_09853_),
    .A(net5835),
    .B(_09852_));
 sg13g2_o21ai_1 _18108_ (.B1(_09853_),
    .Y(_09854_),
    .A1(net5835),
    .A2(_09850_));
 sg13g2_nor2_1 _18109_ (.A(net5834),
    .B(_09854_),
    .Y(_09855_));
 sg13g2_a21oi_1 _18110_ (.A1(net5834),
    .A2(_09849_),
    .Y(_09856_),
    .B1(_09855_));
 sg13g2_nand2_1 _18111_ (.Y(_09857_),
    .A(_00163_),
    .B(_09856_));
 sg13g2_or2_1 _18112_ (.X(_09858_),
    .B(_09856_),
    .A(_00163_));
 sg13g2_nand2_1 _18113_ (.Y(_09859_),
    .A(_09857_),
    .B(_09858_));
 sg13g2_xnor2_1 _18114_ (.Y(_09860_),
    .A(_09833_),
    .B(_09834_));
 sg13g2_nand2_1 _18115_ (.Y(_09861_),
    .A(net5835),
    .B(_09860_));
 sg13g2_nand2b_1 _18116_ (.Y(_09862_),
    .B(net5829),
    .A_N(\atari2600.tia.diag[64] ));
 sg13g2_nor2b_1 _18117_ (.A(_09834_),
    .B_N(_09862_),
    .Y(_09863_));
 sg13g2_a21oi_1 _18118_ (.A1(_08037_),
    .A2(_09863_),
    .Y(_09864_),
    .B1(net5834));
 sg13g2_a22oi_1 _18119_ (.Y(_09865_),
    .B1(_09861_),
    .B2(_09864_),
    .A2(_09854_),
    .A1(net5834));
 sg13g2_xnor2_1 _18120_ (.Y(_09866_),
    .A(_00163_),
    .B(_09865_));
 sg13g2_and2_1 _18121_ (.A(_08037_),
    .B(_09852_),
    .X(_09867_));
 sg13g2_a21oi_1 _18122_ (.A1(\atari2600.tia.p0_scale[0] ),
    .A2(_09843_),
    .Y(_09868_),
    .B1(_09867_));
 sg13g2_nand2b_1 _18123_ (.Y(_09869_),
    .B(_08037_),
    .A_N(_09860_));
 sg13g2_a21oi_1 _18124_ (.A1(net5835),
    .A2(_09851_),
    .Y(_09870_),
    .B1(net5834));
 sg13g2_a22oi_1 _18125_ (.Y(_09871_),
    .B1(_09869_),
    .B2(_09870_),
    .A2(_09868_),
    .A1(net5834));
 sg13g2_xor2_1 _18126_ (.B(_09871_),
    .A(_00163_),
    .X(_09872_));
 sg13g2_mux4_1 _18127_ (.S0(\atari2600.tia.vdelp0 ),
    .A0(\atari2600.tia.diag[104] ),
    .A1(\atari2600.tia.old_grp0[0] ),
    .A2(\atari2600.tia.diag[106] ),
    .A3(\atari2600.tia.old_grp0[2] ),
    .S1(_09872_),
    .X(_09873_));
 sg13g2_mux4_1 _18128_ (.S0(\atari2600.tia.vdelp0 ),
    .A0(\atari2600.tia.diag[105] ),
    .A1(\atari2600.tia.old_grp0[1] ),
    .A2(\atari2600.tia.diag[107] ),
    .A3(\atari2600.tia.old_grp0[3] ),
    .S1(_09872_),
    .X(_09874_));
 sg13g2_nor2b_1 _18129_ (.A(_09866_),
    .B_N(_09873_),
    .Y(_09875_));
 sg13g2_a221oi_1 _18130_ (.B2(_09874_),
    .C1(_09875_),
    .B1(_09866_),
    .A1(_09857_),
    .Y(_09876_),
    .A2(_09858_));
 sg13g2_mux4_1 _18131_ (.S0(\atari2600.tia.vdelp0 ),
    .A0(\atari2600.tia.diag[110] ),
    .A1(\atari2600.tia.old_grp0[6] ),
    .A2(\atari2600.tia.diag[111] ),
    .A3(\atari2600.tia.old_grp0[7] ),
    .S1(_09866_),
    .X(_09877_));
 sg13g2_mux4_1 _18132_ (.S0(\atari2600.tia.vdelp0 ),
    .A0(\atari2600.tia.diag[108] ),
    .A1(\atari2600.tia.old_grp0[4] ),
    .A2(\atari2600.tia.diag[109] ),
    .A3(\atari2600.tia.old_grp0[5] ),
    .S1(_09866_),
    .X(_09878_));
 sg13g2_mux2_1 _18133_ (.A0(_09878_),
    .A1(_09877_),
    .S(_09872_),
    .X(_09879_));
 sg13g2_xor2_1 _18134_ (.B(net5802),
    .A(\atari2600.tia.diag[71] ),
    .X(_09880_));
 sg13g2_xnor2_1 _18135_ (.Y(_09881_),
    .A(\atari2600.tia.diag[70] ),
    .B(net5804));
 sg13g2_a21oi_1 _18136_ (.A1(_07996_),
    .A2(net5810),
    .Y(_09882_),
    .B1(_09846_));
 sg13g2_nor2b_1 _18137_ (.A(_09882_),
    .B_N(_09881_),
    .Y(_09883_));
 sg13g2_a21oi_1 _18138_ (.A1(_07995_),
    .A2(net5804),
    .Y(_09884_),
    .B1(_09883_));
 sg13g2_or2_1 _18139_ (.X(_09885_),
    .B(_09884_),
    .A(_09880_));
 sg13g2_o21ai_1 _18140_ (.B1(_09885_),
    .Y(_09886_),
    .A1(\atari2600.tia.diag[71] ),
    .A2(net5557));
 sg13g2_nand2_1 _18141_ (.Y(_09887_),
    .A(\atari2600.tia.diag[69] ),
    .B(\atari2600.tia.p0_w[5] ));
 sg13g2_xor2_1 _18142_ (.B(\atari2600.tia.p0_w[5] ),
    .A(\atari2600.tia.diag[69] ),
    .X(_09888_));
 sg13g2_nand2_1 _18143_ (.Y(_09889_),
    .A(net5595),
    .B(\atari2600.tia.p0_w[3] ));
 sg13g2_xor2_1 _18144_ (.B(\atari2600.tia.p0_w[4] ),
    .A(\atari2600.tia.diag[68] ),
    .X(_09890_));
 sg13g2_nand2b_1 _18145_ (.Y(_09891_),
    .B(_09890_),
    .A_N(_09889_));
 sg13g2_o21ai_1 _18146_ (.B1(_09891_),
    .Y(_09892_),
    .A1(_07997_),
    .A2(_08036_));
 sg13g2_nand2_1 _18147_ (.Y(_09893_),
    .A(_09888_),
    .B(_09892_));
 sg13g2_nand2_1 _18148_ (.Y(_09894_),
    .A(_09887_),
    .B(_09893_));
 sg13g2_xnor2_1 _18149_ (.Y(_09895_),
    .A(\atari2600.tia.diag[70] ),
    .B(_09894_));
 sg13g2_xor2_1 _18150_ (.B(_09892_),
    .A(_09888_),
    .X(_09896_));
 sg13g2_nand2b_1 _18151_ (.Y(_09897_),
    .B(net5810),
    .A_N(_09896_));
 sg13g2_xnor2_1 _18152_ (.Y(_09898_),
    .A(_09889_),
    .B(_09890_));
 sg13g2_nor2_1 _18153_ (.A(net5814),
    .B(_09898_),
    .Y(_09899_));
 sg13g2_xor2_1 _18154_ (.B(\atari2600.tia.p0_w[3] ),
    .A(net5595),
    .X(_09900_));
 sg13g2_nand2_1 _18155_ (.Y(_09901_),
    .A(net5819),
    .B(_09900_));
 sg13g2_o21ai_1 _18156_ (.B1(_09838_),
    .Y(_09902_),
    .A1(net5819),
    .A2(_09900_));
 sg13g2_nand2_1 _18157_ (.Y(_09903_),
    .A(_09901_),
    .B(_09902_));
 sg13g2_a21oi_1 _18158_ (.A1(_09901_),
    .A2(_09902_),
    .Y(_09904_),
    .B1(_09899_));
 sg13g2_a22oi_1 _18159_ (.Y(_09905_),
    .B1(_09898_),
    .B2(net5814),
    .A2(_09896_),
    .A1(net5809));
 sg13g2_o21ai_1 _18160_ (.B1(_09905_),
    .Y(_09906_),
    .A1(net5809),
    .A2(_09896_));
 sg13g2_o21ai_1 _18161_ (.B1(_09897_),
    .Y(_09907_),
    .A1(_09904_),
    .A2(_09906_));
 sg13g2_xnor2_1 _18162_ (.Y(_09908_),
    .A(net5803),
    .B(_09895_));
 sg13g2_a22oi_1 _18163_ (.Y(_09909_),
    .B1(_09907_),
    .B2(_09908_),
    .A2(_09895_),
    .A1(net5804));
 sg13g2_nand3_1 _18164_ (.B(_09888_),
    .C(_09892_),
    .A(\atari2600.tia.diag[70] ),
    .Y(_09910_));
 sg13g2_o21ai_1 _18165_ (.B1(_09910_),
    .Y(_09911_),
    .A1(_00160_),
    .A2(_09887_));
 sg13g2_xnor2_1 _18166_ (.Y(_09912_),
    .A(\atari2600.tia.diag[71] ),
    .B(_09911_));
 sg13g2_xor2_1 _18167_ (.B(_09911_),
    .A(_09880_),
    .X(_09913_));
 sg13g2_nor2_1 _18168_ (.A(_09909_),
    .B(_09913_),
    .Y(_09914_));
 sg13g2_a21oi_1 _18169_ (.A1(_08124_),
    .A2(_09912_),
    .Y(_09915_),
    .B1(_09914_));
 sg13g2_nand2b_1 _18170_ (.Y(_09916_),
    .B(net5805),
    .A_N(\atari2600.tia.p0_spacing[5] ));
 sg13g2_xor2_1 _18171_ (.B(net5805),
    .A(\atari2600.tia.p0_spacing[5] ),
    .X(_09917_));
 sg13g2_nor2_1 _18172_ (.A(_08038_),
    .B(net5813),
    .Y(_09918_));
 sg13g2_o21ai_1 _18173_ (.B1(_09916_),
    .Y(_09919_),
    .A1(_09917_),
    .A2(_09918_));
 sg13g2_xor2_1 _18174_ (.B(net5802),
    .A(\atari2600.tia.p0_spacing[6] ),
    .X(_09920_));
 sg13g2_xnor2_1 _18175_ (.Y(_09921_),
    .A(_09919_),
    .B(_09920_));
 sg13g2_xnor2_1 _18176_ (.Y(_09922_),
    .A(_09917_),
    .B(_09918_));
 sg13g2_xnor2_1 _18177_ (.Y(_09923_),
    .A(\atari2600.tia.p0_spacing[4] ),
    .B(net5810));
 sg13g2_nand2b_1 _18178_ (.Y(_09924_),
    .B(_00161_),
    .A_N(_09923_));
 sg13g2_xnor2_1 _18179_ (.Y(_09925_),
    .A(net5593),
    .B(_09923_));
 sg13g2_o21ai_1 _18180_ (.B1(_09924_),
    .Y(_09926_),
    .A1(_09844_),
    .A2(_09925_));
 sg13g2_xnor2_1 _18181_ (.Y(_09927_),
    .A(_00160_),
    .B(_09922_));
 sg13g2_nand2_1 _18182_ (.Y(_09928_),
    .A(_09926_),
    .B(_09927_));
 sg13g2_o21ai_1 _18183_ (.B1(_09928_),
    .Y(_09929_),
    .A1(\atari2600.tia.diag[70] ),
    .A2(_09922_));
 sg13g2_xnor2_1 _18184_ (.Y(_09930_),
    .A(\atari2600.tia.diag[71] ),
    .B(_09921_));
 sg13g2_a22oi_1 _18185_ (.Y(_09931_),
    .B1(_09929_),
    .B2(_09930_),
    .A2(_09921_),
    .A1(_00162_));
 sg13g2_and2_1 _18186_ (.A(net5563),
    .B(_09900_),
    .X(_09932_));
 sg13g2_xnor2_1 _18187_ (.Y(_09933_),
    .A(net5819),
    .B(_09900_));
 sg13g2_a221oi_1 _18188_ (.B2(_09862_),
    .C1(_09832_),
    .B1(_09831_),
    .A1(net5596),
    .Y(_09934_),
    .A2(net5561));
 sg13g2_nor3_1 _18189_ (.A(_09829_),
    .B(_09933_),
    .C(_09934_),
    .Y(_09935_));
 sg13g2_nor3_1 _18190_ (.A(_09830_),
    .B(_09833_),
    .C(_09933_),
    .Y(_09936_));
 sg13g2_a21oi_1 _18191_ (.A1(_09863_),
    .A2(_09936_),
    .Y(_09937_),
    .B1(_09899_));
 sg13g2_o21ai_1 _18192_ (.B1(_09937_),
    .Y(_09938_),
    .A1(_09932_),
    .A2(_09935_));
 sg13g2_a22oi_1 _18193_ (.Y(_09939_),
    .B1(_09923_),
    .B2(_09896_),
    .A2(_09898_),
    .A1(net5814));
 sg13g2_nand2b_1 _18194_ (.Y(_09940_),
    .B(_09895_),
    .A_N(_09922_));
 sg13g2_o21ai_1 _18195_ (.B1(_09940_),
    .Y(_09941_),
    .A1(_09896_),
    .A2(_09923_));
 sg13g2_a21oi_1 _18196_ (.A1(_09938_),
    .A2(_09939_),
    .Y(_09942_),
    .B1(_09941_));
 sg13g2_nand2b_1 _18197_ (.Y(_09943_),
    .B(_09922_),
    .A_N(_09895_));
 sg13g2_o21ai_1 _18198_ (.B1(_09943_),
    .Y(_09944_),
    .A1(_09912_),
    .A2(_09921_));
 sg13g2_nand2_1 _18199_ (.Y(_09945_),
    .A(_09912_),
    .B(_09921_));
 sg13g2_o21ai_1 _18200_ (.B1(_09945_),
    .Y(_09946_),
    .A1(_09942_),
    .A2(_09944_));
 sg13g2_nor3_1 _18201_ (.A(_08115_),
    .B(_09931_),
    .C(_09946_),
    .Y(_09947_));
 sg13g2_nor2_1 _18202_ (.A(\atari2600.tia.p0_spacing[6] ),
    .B(net5558),
    .Y(_09948_));
 sg13g2_nand2_1 _18203_ (.Y(_09949_),
    .A(\atari2600.tia.p0_spacing[4] ),
    .B(net5560));
 sg13g2_xnor2_1 _18204_ (.Y(_09950_),
    .A(\atari2600.tia.p0_spacing[5] ),
    .B(net5813));
 sg13g2_nand2_1 _18205_ (.Y(_09951_),
    .A(_09949_),
    .B(_09950_));
 sg13g2_o21ai_1 _18206_ (.B1(_09951_),
    .Y(_09952_),
    .A1(\atari2600.tia.p0_spacing[5] ),
    .A2(net5559));
 sg13g2_xnor2_1 _18207_ (.Y(_09953_),
    .A(\atari2600.tia.p0_spacing[6] ),
    .B(net5805));
 sg13g2_a21oi_1 _18208_ (.A1(_09952_),
    .A2(_09953_),
    .Y(_09954_),
    .B1(_09948_));
 sg13g2_xnor2_1 _18209_ (.Y(_09955_),
    .A(_00150_),
    .B(_09954_));
 sg13g2_nand2_1 _18210_ (.Y(_09956_),
    .A(_00162_),
    .B(_09955_));
 sg13g2_xor2_1 _18211_ (.B(_09953_),
    .A(_09952_),
    .X(_09957_));
 sg13g2_xnor2_1 _18212_ (.Y(_09958_),
    .A(_09949_),
    .B(_09950_));
 sg13g2_xnor2_1 _18213_ (.Y(_09959_),
    .A(\atari2600.tia.p0_spacing[4] ),
    .B(net5818));
 sg13g2_o21ai_1 _18214_ (.B1(_09840_),
    .Y(_09960_),
    .A1(\atari2600.tia.diag[68] ),
    .A2(_09959_));
 sg13g2_nand2_1 _18215_ (.Y(_09961_),
    .A(net5594),
    .B(_09959_));
 sg13g2_xnor2_1 _18216_ (.Y(_09962_),
    .A(_00161_),
    .B(_09958_));
 sg13g2_nand3_1 _18217_ (.B(_09961_),
    .C(_09962_),
    .A(_09960_),
    .Y(_09963_));
 sg13g2_o21ai_1 _18218_ (.B1(_09963_),
    .Y(_09964_),
    .A1(net5593),
    .A2(_09958_));
 sg13g2_xor2_1 _18219_ (.B(_09957_),
    .A(_00160_),
    .X(_09965_));
 sg13g2_a22oi_1 _18220_ (.Y(_09966_),
    .B1(_09964_),
    .B2(_09965_),
    .A2(_09957_),
    .A1(_07995_));
 sg13g2_xor2_1 _18221_ (.B(_09955_),
    .A(\atari2600.tia.diag[71] ),
    .X(_09967_));
 sg13g2_o21ai_1 _18222_ (.B1(_09956_),
    .Y(_09968_),
    .A1(_09966_),
    .A2(_09967_));
 sg13g2_o21ai_1 _18223_ (.B1(_09903_),
    .Y(_09969_),
    .A1(_09898_),
    .A2(_09959_));
 sg13g2_a22oi_1 _18224_ (.Y(_09970_),
    .B1(_09959_),
    .B2(_09898_),
    .A2(_09958_),
    .A1(_09896_));
 sg13g2_nor2_1 _18225_ (.A(_09896_),
    .B(_09958_),
    .Y(_09971_));
 sg13g2_a221oi_1 _18226_ (.B2(_09970_),
    .C1(_09971_),
    .B1(_09969_),
    .A1(_09895_),
    .Y(_09972_),
    .A2(_09957_));
 sg13g2_nor2_1 _18227_ (.A(_09895_),
    .B(_09957_),
    .Y(_09973_));
 sg13g2_nor2_1 _18228_ (.A(_09972_),
    .B(_09973_),
    .Y(_09974_));
 sg13g2_o21ai_1 _18229_ (.B1(_09974_),
    .Y(_09975_),
    .A1(_09912_),
    .A2(_09955_));
 sg13g2_o21ai_1 _18230_ (.B1(_09975_),
    .Y(_09976_),
    .A1(\atari2600.tia.p0_copies[2] ),
    .A2(\atari2600.tia.p0_copies[1] ));
 sg13g2_a21oi_1 _18231_ (.A1(_09912_),
    .A2(_09955_),
    .Y(_09977_),
    .B1(_09976_));
 sg13g2_a221oi_1 _18232_ (.B2(_09977_),
    .C1(_09947_),
    .B1(_09968_),
    .A1(_09886_),
    .Y(_09978_),
    .A2(_09915_));
 sg13g2_nand2_1 _18233_ (.Y(_09979_),
    .A(net5835),
    .B(_09885_));
 sg13g2_a21oi_1 _18234_ (.A1(_09880_),
    .A2(_09884_),
    .Y(_09980_),
    .B1(_09979_));
 sg13g2_xor2_1 _18235_ (.B(_09882_),
    .A(_09881_),
    .X(_09981_));
 sg13g2_o21ai_1 _18236_ (.B1(_09981_),
    .Y(_09982_),
    .A1(net5835),
    .A2(_09847_));
 sg13g2_o21ai_1 _18237_ (.B1(\atari2600.tia.p0_scale[1] ),
    .Y(_09983_),
    .A1(_09980_),
    .A2(_09982_));
 sg13g2_a21oi_1 _18238_ (.A1(_09849_),
    .A2(_09868_),
    .Y(_09984_),
    .B1(net5834));
 sg13g2_o21ai_1 _18239_ (.B1(_09983_),
    .Y(_09985_),
    .A1(_09859_),
    .A2(_09879_));
 sg13g2_nor4_1 _18240_ (.A(_09876_),
    .B(_09978_),
    .C(_09984_),
    .D(_09985_),
    .Y(_09986_));
 sg13g2_nand2_2 _18241_ (.Y(_09987_),
    .A(net5216),
    .B(net4584));
 sg13g2_inv_1 _18242_ (.Y(_09988_),
    .A(_09987_));
 sg13g2_o21ai_1 _18243_ (.B1(_09661_),
    .Y(_00021_),
    .A1(net4770),
    .A2(_09987_));
 sg13g2_nand2_1 _18244_ (.Y(_09989_),
    .A(\atari2600.tia.diag[43] ),
    .B(\atari2600.tia.m1_w[3] ));
 sg13g2_and2_1 _18245_ (.A(\atari2600.tia.diag[42] ),
    .B(\atari2600.tia.m1_w[2] ),
    .X(_09990_));
 sg13g2_xor2_1 _18246_ (.B(\atari2600.tia.m1_w[2] ),
    .A(\atari2600.tia.diag[42] ),
    .X(_09991_));
 sg13g2_nand2_1 _18247_ (.Y(_09992_),
    .A(\atari2600.tia.diag[41] ),
    .B(\atari2600.tia.m1_w[1] ));
 sg13g2_xnor2_1 _18248_ (.Y(_09993_),
    .A(\atari2600.tia.diag[41] ),
    .B(\atari2600.tia.m1_w[1] ));
 sg13g2_nand2_1 _18249_ (.Y(_09994_),
    .A(\atari2600.tia.diag[40] ),
    .B(\atari2600.tia.m1_w[0] ));
 sg13g2_o21ai_1 _18250_ (.B1(_09992_),
    .Y(_09995_),
    .A1(_09993_),
    .A2(_09994_));
 sg13g2_a21o_1 _18251_ (.A2(_09995_),
    .A1(_09991_),
    .B1(_09990_),
    .X(_09996_));
 sg13g2_xor2_1 _18252_ (.B(\atari2600.tia.m1_w[3] ),
    .A(\atari2600.tia.diag[43] ),
    .X(_09997_));
 sg13g2_nand2_1 _18253_ (.Y(_09998_),
    .A(_09996_),
    .B(_09997_));
 sg13g2_nand2_1 _18254_ (.Y(_09999_),
    .A(_09989_),
    .B(_09998_));
 sg13g2_a21oi_2 _18255_ (.B1(_07986_),
    .Y(_10000_),
    .A2(_09998_),
    .A1(_09989_));
 sg13g2_nand3_1 _18256_ (.B(\atari2600.tia.diag[45] ),
    .C(_10000_),
    .A(\atari2600.tia.diag[46] ),
    .Y(_10001_));
 sg13g2_xor2_1 _18257_ (.B(_10001_),
    .A(\atari2600.tia.diag[47] ),
    .X(_10002_));
 sg13g2_nor2_1 _18258_ (.A(net5801),
    .B(_10002_),
    .Y(_10003_));
 sg13g2_a21o_1 _18259_ (.A2(_10000_),
    .A1(\atari2600.tia.diag[45] ),
    .B1(\atari2600.tia.diag[46] ),
    .X(_10004_));
 sg13g2_nand2_1 _18260_ (.Y(_10005_),
    .A(_10001_),
    .B(_10004_));
 sg13g2_xnor2_1 _18261_ (.Y(_10006_),
    .A(\atari2600.tia.diag[45] ),
    .B(_10000_));
 sg13g2_nor2_1 _18262_ (.A(net5812),
    .B(_10006_),
    .Y(_10007_));
 sg13g2_xnor2_1 _18263_ (.Y(_10008_),
    .A(\atari2600.tia.diag[40] ),
    .B(\atari2600.tia.m1_w[0] ));
 sg13g2_xnor2_1 _18264_ (.Y(_10009_),
    .A(_09996_),
    .B(_09997_));
 sg13g2_nand2_1 _18265_ (.Y(_10010_),
    .A(net5820),
    .B(_10009_));
 sg13g2_nand2b_1 _18266_ (.Y(_10011_),
    .B(net5563),
    .A_N(_10009_));
 sg13g2_xnor2_1 _18267_ (.Y(_10012_),
    .A(_09991_),
    .B(_09995_));
 sg13g2_xnor2_1 _18268_ (.Y(_10013_),
    .A(_00151_),
    .B(_10012_));
 sg13g2_nand3_1 _18269_ (.B(_10011_),
    .C(_10013_),
    .A(_10010_),
    .Y(_10014_));
 sg13g2_inv_1 _18270_ (.Y(_10015_),
    .A(_10014_));
 sg13g2_xnor2_1 _18271_ (.Y(_10016_),
    .A(_09993_),
    .B(_09994_));
 sg13g2_xor2_1 _18272_ (.B(_10016_),
    .A(_00164_),
    .X(_10017_));
 sg13g2_xnor2_1 _18273_ (.Y(_10018_),
    .A(_07986_),
    .B(_09999_));
 sg13g2_nand2_1 _18274_ (.Y(_10019_),
    .A(net5815),
    .B(_10018_));
 sg13g2_inv_1 _18275_ (.Y(_10020_),
    .A(_10019_));
 sg13g2_o21ai_1 _18276_ (.B1(_10011_),
    .Y(_10021_),
    .A1(net5823),
    .A2(_10012_));
 sg13g2_a21o_1 _18277_ (.A2(_10008_),
    .A1(net5831),
    .B1(_10017_),
    .X(_10022_));
 sg13g2_o21ai_1 _18278_ (.B1(_10022_),
    .Y(_10023_),
    .A1(net5828),
    .A2(_10016_));
 sg13g2_a221oi_1 _18279_ (.B2(_10015_),
    .C1(_10020_),
    .B1(_10023_),
    .A1(_10010_),
    .Y(_10024_),
    .A2(_10021_));
 sg13g2_xor2_1 _18280_ (.B(_10006_),
    .A(net5809),
    .X(_10025_));
 sg13g2_nor2_1 _18281_ (.A(net5815),
    .B(_10018_),
    .Y(_10026_));
 sg13g2_nor3_1 _18282_ (.A(_10024_),
    .B(_10025_),
    .C(_10026_),
    .Y(_10027_));
 sg13g2_xnor2_1 _18283_ (.Y(_10028_),
    .A(net5803),
    .B(_10005_));
 sg13g2_o21ai_1 _18284_ (.B1(_10028_),
    .Y(_10029_),
    .A1(_10007_),
    .A2(_10027_));
 sg13g2_o21ai_1 _18285_ (.B1(_10029_),
    .Y(_10030_),
    .A1(net5808),
    .A2(_10005_));
 sg13g2_xor2_1 _18286_ (.B(_10008_),
    .A(_00165_),
    .X(_10031_));
 sg13g2_nor2_1 _18287_ (.A(_10014_),
    .B(_10026_),
    .Y(_10032_));
 sg13g2_nor2_1 _18288_ (.A(_10025_),
    .B(_10031_),
    .Y(_10033_));
 sg13g2_nor2_1 _18289_ (.A(_10017_),
    .B(_10020_),
    .Y(_10034_));
 sg13g2_nand4_1 _18290_ (.B(_10032_),
    .C(_10033_),
    .A(_10028_),
    .Y(_10035_),
    .D(_10034_));
 sg13g2_a21oi_1 _18291_ (.A1(_10030_),
    .A2(_10035_),
    .Y(_10036_),
    .B1(_10003_));
 sg13g2_nor2_1 _18292_ (.A(\atari2600.tia.diag[47] ),
    .B(_08114_),
    .Y(_10037_));
 sg13g2_nor2_1 _18293_ (.A(\atari2600.tia.diag[42] ),
    .B(net5562),
    .Y(_10038_));
 sg13g2_nor2_1 _18294_ (.A(\atari2600.tia.diag[41] ),
    .B(_08107_),
    .Y(_10039_));
 sg13g2_a22oi_1 _18295_ (.Y(_10040_),
    .B1(_08108_),
    .B2(\atari2600.tia.diag[40] ),
    .A2(_08107_),
    .A1(\atari2600.tia.diag[41] ));
 sg13g2_or3_1 _18296_ (.A(_10038_),
    .B(_10039_),
    .C(_10040_),
    .X(_10041_));
 sg13g2_a22oi_1 _18297_ (.Y(_10042_),
    .B1(net5561),
    .B2(\atari2600.tia.diag[42] ),
    .A2(net5563),
    .A1(\atari2600.tia.diag[43] ));
 sg13g2_nor2_1 _18298_ (.A(\atari2600.tia.diag[43] ),
    .B(net5563),
    .Y(_10043_));
 sg13g2_a221oi_1 _18299_ (.B2(_10042_),
    .C1(_10043_),
    .B1(_10041_),
    .A1(_07986_),
    .Y(_10044_),
    .A2(net5817));
 sg13g2_a221oi_1 _18300_ (.B2(\atari2600.tia.diag[45] ),
    .C1(_10044_),
    .B1(_08112_),
    .A1(\atari2600.tia.diag[44] ),
    .Y(_10045_),
    .A2(_08111_));
 sg13g2_a221oi_1 _18301_ (.B2(_07984_),
    .C1(_10045_),
    .B1(net5808),
    .A1(_07985_),
    .Y(_10046_),
    .A2(net5812));
 sg13g2_a21oi_1 _18302_ (.A1(\atari2600.tia.diag[46] ),
    .A2(_08113_),
    .Y(_10047_),
    .B1(_10046_));
 sg13g2_o21ai_1 _18303_ (.B1(\atari2600.tia.enam1 ),
    .Y(_10048_),
    .A1(_10037_),
    .A2(_10047_));
 sg13g2_a21oi_1 _18304_ (.A1(net5801),
    .A2(_10002_),
    .Y(_10049_),
    .B1(_10048_));
 sg13g2_nand2b_1 _18305_ (.Y(_10050_),
    .B(_10049_),
    .A_N(_10036_));
 sg13g2_a21oi_2 _18306_ (.B1(_10050_),
    .Y(_10051_),
    .A2(_08114_),
    .A1(\atari2600.tia.diag[47] ));
 sg13g2_inv_2 _18307_ (.Y(_10052_),
    .A(net4768));
 sg13g2_nand2_1 _18308_ (.Y(_10053_),
    .A(\atari2600.tia.diag[51] ),
    .B(\atari2600.tia.m0_w[3] ));
 sg13g2_and2_1 _18309_ (.A(\atari2600.tia.diag[50] ),
    .B(\atari2600.tia.m0_w[2] ),
    .X(_10054_));
 sg13g2_xor2_1 _18310_ (.B(\atari2600.tia.m0_w[2] ),
    .A(\atari2600.tia.diag[50] ),
    .X(_10055_));
 sg13g2_nand2_1 _18311_ (.Y(_10056_),
    .A(\atari2600.tia.diag[49] ),
    .B(\atari2600.tia.m0_w[1] ));
 sg13g2_nor2_1 _18312_ (.A(\atari2600.tia.diag[49] ),
    .B(\atari2600.tia.m0_w[1] ),
    .Y(_10057_));
 sg13g2_xor2_1 _18313_ (.B(\atari2600.tia.m0_w[1] ),
    .A(\atari2600.tia.diag[49] ),
    .X(_10058_));
 sg13g2_nand2_1 _18314_ (.Y(_10059_),
    .A(\atari2600.tia.diag[48] ),
    .B(\atari2600.tia.m0_w[0] ));
 sg13g2_o21ai_1 _18315_ (.B1(_10056_),
    .Y(_10060_),
    .A1(_10057_),
    .A2(_10059_));
 sg13g2_a21o_1 _18316_ (.A2(_10060_),
    .A1(_10055_),
    .B1(_10054_),
    .X(_10061_));
 sg13g2_xor2_1 _18317_ (.B(\atari2600.tia.m0_w[3] ),
    .A(\atari2600.tia.diag[51] ),
    .X(_10062_));
 sg13g2_nand2_1 _18318_ (.Y(_10063_),
    .A(_10061_),
    .B(_10062_));
 sg13g2_a21oi_2 _18319_ (.B1(_07990_),
    .Y(_10064_),
    .A2(_10063_),
    .A1(_10053_));
 sg13g2_nand3_1 _18320_ (.B(\atari2600.tia.diag[53] ),
    .C(_10064_),
    .A(\atari2600.tia.diag[54] ),
    .Y(_10065_));
 sg13g2_xnor2_1 _18321_ (.Y(_10066_),
    .A(_07987_),
    .B(_10065_));
 sg13g2_a21o_1 _18322_ (.A2(_10064_),
    .A1(\atari2600.tia.diag[53] ),
    .B1(\atari2600.tia.diag[54] ),
    .X(_10067_));
 sg13g2_nand2_1 _18323_ (.Y(_10068_),
    .A(_10065_),
    .B(_10067_));
 sg13g2_nor2_1 _18324_ (.A(net5804),
    .B(_10068_),
    .Y(_10069_));
 sg13g2_xnor2_1 _18325_ (.Y(_10070_),
    .A(\atari2600.tia.diag[53] ),
    .B(_10064_));
 sg13g2_nand3_1 _18326_ (.B(_10053_),
    .C(_10063_),
    .A(_07990_),
    .Y(_10071_));
 sg13g2_nor2b_1 _18327_ (.A(_10064_),
    .B_N(_10071_),
    .Y(_10072_));
 sg13g2_and2_1 _18328_ (.A(net5814),
    .B(_10072_),
    .X(_10073_));
 sg13g2_xnor2_1 _18329_ (.Y(_10074_),
    .A(_10061_),
    .B(_10062_));
 sg13g2_nand2_1 _18330_ (.Y(_10075_),
    .A(net5820),
    .B(_10074_));
 sg13g2_o21ai_1 _18331_ (.B1(_10075_),
    .Y(_10076_),
    .A1(net5814),
    .A2(_10072_));
 sg13g2_inv_1 _18332_ (.Y(_10077_),
    .A(_10076_));
 sg13g2_xnor2_1 _18333_ (.Y(_10078_),
    .A(_10058_),
    .B(_10059_));
 sg13g2_xnor2_1 _18334_ (.Y(_10079_),
    .A(\atari2600.tia.diag[48] ),
    .B(\atari2600.tia.m0_w[0] ));
 sg13g2_xnor2_1 _18335_ (.Y(_10080_),
    .A(_00164_),
    .B(_10078_));
 sg13g2_a21oi_1 _18336_ (.A1(net5829),
    .A2(_10079_),
    .Y(_10081_),
    .B1(_10080_));
 sg13g2_a21oi_1 _18337_ (.A1(_08107_),
    .A2(_10078_),
    .Y(_10082_),
    .B1(_10081_));
 sg13g2_xnor2_1 _18338_ (.Y(_10083_),
    .A(_10055_),
    .B(_10060_));
 sg13g2_xnor2_1 _18339_ (.Y(_10084_),
    .A(_00151_),
    .B(_10083_));
 sg13g2_nor2b_1 _18340_ (.A(_10082_),
    .B_N(_10084_),
    .Y(_10085_));
 sg13g2_nor2_1 _18341_ (.A(net5823),
    .B(_10083_),
    .Y(_10086_));
 sg13g2_nor2_1 _18342_ (.A(net5820),
    .B(_10074_),
    .Y(_10087_));
 sg13g2_nor3_1 _18343_ (.A(_10085_),
    .B(_10086_),
    .C(_10087_),
    .Y(_10088_));
 sg13g2_nor2_1 _18344_ (.A(_10076_),
    .B(_10088_),
    .Y(_10089_));
 sg13g2_xnor2_1 _18345_ (.Y(_10090_),
    .A(net5809),
    .B(_10070_));
 sg13g2_o21ai_1 _18346_ (.B1(_10090_),
    .Y(_10091_),
    .A1(_10073_),
    .A2(_10089_));
 sg13g2_o21ai_1 _18347_ (.B1(_10091_),
    .Y(_10092_),
    .A1(net5810),
    .A2(_10070_));
 sg13g2_xnor2_1 _18348_ (.Y(_10093_),
    .A(net5803),
    .B(_10068_));
 sg13g2_a21oi_1 _18349_ (.A1(_10092_),
    .A2(_10093_),
    .Y(_10094_),
    .B1(_10069_));
 sg13g2_xor2_1 _18350_ (.B(_10079_),
    .A(_00165_),
    .X(_10095_));
 sg13g2_nor4_1 _18351_ (.A(_10073_),
    .B(_10080_),
    .C(_10087_),
    .D(_10095_),
    .Y(_10096_));
 sg13g2_and4_1 _18352_ (.A(_10077_),
    .B(_10084_),
    .C(_10090_),
    .D(_10096_),
    .X(_10097_));
 sg13g2_a21o_1 _18353_ (.A2(_10097_),
    .A1(_10093_),
    .B1(_10094_),
    .X(_10098_));
 sg13g2_o21ai_1 _18354_ (.B1(_10098_),
    .Y(_10099_),
    .A1(net5800),
    .A2(_10066_));
 sg13g2_nand2_1 _18355_ (.Y(_10100_),
    .A(net5800),
    .B(_10066_));
 sg13g2_nand2_1 _18356_ (.Y(_10101_),
    .A(_07987_),
    .B(net5800));
 sg13g2_nand2_1 _18357_ (.Y(_10102_),
    .A(_07990_),
    .B(net5818));
 sg13g2_nand2b_1 _18358_ (.Y(_10103_),
    .B(net5825),
    .A_N(\atari2600.tia.diag[49] ));
 sg13g2_nand3_1 _18359_ (.B(_08108_),
    .C(_10103_),
    .A(\atari2600.tia.diag[48] ),
    .Y(_10104_));
 sg13g2_a22oi_1 _18360_ (.Y(_10105_),
    .B1(net5561),
    .B2(\atari2600.tia.diag[50] ),
    .A2(_08107_),
    .A1(\atari2600.tia.diag[49] ));
 sg13g2_a22oi_1 _18361_ (.Y(_10106_),
    .B1(_10104_),
    .B2(_10105_),
    .A2(net5823),
    .A1(_07991_));
 sg13g2_o21ai_1 _18362_ (.B1(_10106_),
    .Y(_10107_),
    .A1(\atari2600.tia.diag[51] ),
    .A2(net5563));
 sg13g2_a22oi_1 _18363_ (.Y(_10108_),
    .B1(net5560),
    .B2(\atari2600.tia.diag[52] ),
    .A2(net5563),
    .A1(\atari2600.tia.diag[51] ));
 sg13g2_nand2_1 _18364_ (.Y(_10109_),
    .A(_10107_),
    .B(_10108_));
 sg13g2_a22oi_1 _18365_ (.Y(_10110_),
    .B1(_10102_),
    .B2(_10109_),
    .A2(net5559),
    .A1(\atari2600.tia.diag[53] ));
 sg13g2_a221oi_1 _18366_ (.B2(_07988_),
    .C1(_10110_),
    .B1(net5804),
    .A1(_07989_),
    .Y(_10111_),
    .A2(net5810));
 sg13g2_nand2_1 _18367_ (.Y(_10112_),
    .A(\atari2600.tia.diag[54] ),
    .B(net5558));
 sg13g2_o21ai_1 _18368_ (.B1(_10112_),
    .Y(_10113_),
    .A1(_07987_),
    .A2(net5800));
 sg13g2_o21ai_1 _18369_ (.B1(_10101_),
    .Y(_10114_),
    .A1(_10111_),
    .A2(_10113_));
 sg13g2_nand4_1 _18370_ (.B(_10099_),
    .C(_10100_),
    .A(net7380),
    .Y(_10115_),
    .D(_10114_));
 sg13g2_or2_1 _18371_ (.X(_10116_),
    .B(net4784),
    .A(_09827_));
 sg13g2_inv_1 _18372_ (.Y(_10117_),
    .A(_10116_));
 sg13g2_a22oi_1 _18373_ (.Y(_10118_),
    .B1(net4768),
    .B2(_10117_),
    .A2(net5197),
    .A1(net3955));
 sg13g2_inv_1 _18374_ (.Y(_00015_),
    .A(_10118_));
 sg13g2_nand2_1 _18375_ (.Y(_10119_),
    .A(\atari2600.tia.diag[35] ),
    .B(\atari2600.tia.ball_w[3] ));
 sg13g2_xor2_1 _18376_ (.B(\atari2600.tia.ball_w[2] ),
    .A(\atari2600.tia.diag[34] ),
    .X(_10120_));
 sg13g2_nand2_1 _18377_ (.Y(_10121_),
    .A(\atari2600.tia.diag[33] ),
    .B(\atari2600.tia.ball_w[1] ));
 sg13g2_xnor2_1 _18378_ (.Y(_10122_),
    .A(\atari2600.tia.diag[33] ),
    .B(\atari2600.tia.ball_w[1] ));
 sg13g2_nand2_1 _18379_ (.Y(_10123_),
    .A(\atari2600.tia.diag[32] ),
    .B(\atari2600.tia.ball_w[0] ));
 sg13g2_o21ai_1 _18380_ (.B1(_10121_),
    .Y(_10124_),
    .A1(_10122_),
    .A2(_10123_));
 sg13g2_nand2_1 _18381_ (.Y(_10125_),
    .A(_10120_),
    .B(_10124_));
 sg13g2_o21ai_1 _18382_ (.B1(_10125_),
    .Y(_10126_),
    .A1(_07982_),
    .A2(_08035_));
 sg13g2_xor2_1 _18383_ (.B(\atari2600.tia.ball_w[3] ),
    .A(\atari2600.tia.diag[35] ),
    .X(_10127_));
 sg13g2_nand2_1 _18384_ (.Y(_10128_),
    .A(_10126_),
    .B(_10127_));
 sg13g2_nand2_1 _18385_ (.Y(_10129_),
    .A(_10119_),
    .B(_10128_));
 sg13g2_a21oi_2 _18386_ (.B1(_07980_),
    .Y(_10130_),
    .A2(_10128_),
    .A1(_10119_));
 sg13g2_nand3_1 _18387_ (.B(\atari2600.tia.diag[37] ),
    .C(_10130_),
    .A(\atari2600.tia.diag[38] ),
    .Y(_10131_));
 sg13g2_xor2_1 _18388_ (.B(_10131_),
    .A(\atari2600.tia.diag[39] ),
    .X(_10132_));
 sg13g2_nor2_1 _18389_ (.A(net5801),
    .B(_10132_),
    .Y(_10133_));
 sg13g2_a21o_1 _18390_ (.A2(_10130_),
    .A1(\atari2600.tia.diag[37] ),
    .B1(\atari2600.tia.diag[38] ),
    .X(_10134_));
 sg13g2_nand2_1 _18391_ (.Y(_10135_),
    .A(_10131_),
    .B(_10134_));
 sg13g2_nand3_1 _18392_ (.B(_10131_),
    .C(_10134_),
    .A(net5558),
    .Y(_10136_));
 sg13g2_xnor2_1 _18393_ (.Y(_10137_),
    .A(\atari2600.tia.diag[37] ),
    .B(_10130_));
 sg13g2_nor2_1 _18394_ (.A(net5812),
    .B(_10137_),
    .Y(_10138_));
 sg13g2_xor2_1 _18395_ (.B(_10137_),
    .A(net5809),
    .X(_10139_));
 sg13g2_xnor2_1 _18396_ (.Y(_10140_),
    .A(_10122_),
    .B(_10123_));
 sg13g2_xnor2_1 _18397_ (.Y(_10141_),
    .A(\atari2600.tia.diag[32] ),
    .B(\atari2600.tia.ball_w[0] ));
 sg13g2_xor2_1 _18398_ (.B(_10140_),
    .A(_00164_),
    .X(_10142_));
 sg13g2_a21o_1 _18399_ (.A2(_10141_),
    .A1(net5830),
    .B1(_10142_),
    .X(_10143_));
 sg13g2_o21ai_1 _18400_ (.B1(_10143_),
    .Y(_10144_),
    .A1(net5826),
    .A2(_10140_));
 sg13g2_xnor2_1 _18401_ (.Y(_10145_),
    .A(_07980_),
    .B(_10129_));
 sg13g2_nor2_1 _18402_ (.A(net5814),
    .B(_10145_),
    .Y(_10146_));
 sg13g2_xnor2_1 _18403_ (.Y(_10147_),
    .A(_10126_),
    .B(_10127_));
 sg13g2_nand2_1 _18404_ (.Y(_10148_),
    .A(\atari2600.tia.vid_xpos[3] ),
    .B(_10147_));
 sg13g2_xor2_1 _18405_ (.B(_10124_),
    .A(_10120_),
    .X(_10149_));
 sg13g2_xnor2_1 _18406_ (.Y(_10150_),
    .A(_00151_),
    .B(_10149_));
 sg13g2_xnor2_1 _18407_ (.Y(_10151_),
    .A(\atari2600.tia.vid_xpos[3] ),
    .B(_10147_));
 sg13g2_nor3_1 _18408_ (.A(_10146_),
    .B(_10150_),
    .C(_10151_),
    .Y(_10152_));
 sg13g2_nand2_1 _18409_ (.Y(_10153_),
    .A(net5815),
    .B(_10145_));
 sg13g2_nand2_1 _18410_ (.Y(_10154_),
    .A(net5562),
    .B(_10149_));
 sg13g2_o21ai_1 _18411_ (.B1(_10154_),
    .Y(_10155_),
    .A1(net5822),
    .A2(_10147_));
 sg13g2_nand2_1 _18412_ (.Y(_10156_),
    .A(_10148_),
    .B(_10155_));
 sg13g2_o21ai_1 _18413_ (.B1(_10153_),
    .Y(_10157_),
    .A1(_10146_),
    .A2(_10156_));
 sg13g2_a21oi_1 _18414_ (.A1(_10144_),
    .A2(_10152_),
    .Y(_10158_),
    .B1(_10157_));
 sg13g2_nor2_1 _18415_ (.A(_10139_),
    .B(_10158_),
    .Y(_10159_));
 sg13g2_xnor2_1 _18416_ (.Y(_10160_),
    .A(net5803),
    .B(_10135_));
 sg13g2_o21ai_1 _18417_ (.B1(_10160_),
    .Y(_10161_),
    .A1(_10138_),
    .A2(_10159_));
 sg13g2_xor2_1 _18418_ (.B(_10141_),
    .A(_00165_),
    .X(_10162_));
 sg13g2_nor2_1 _18419_ (.A(_10142_),
    .B(_10162_),
    .Y(_10163_));
 sg13g2_nand3_1 _18420_ (.B(_10153_),
    .C(_10163_),
    .A(_10152_),
    .Y(_10164_));
 sg13g2_nor2_1 _18421_ (.A(_10139_),
    .B(_10164_),
    .Y(_10165_));
 sg13g2_a22oi_1 _18422_ (.Y(_10166_),
    .B1(_10165_),
    .B2(_10160_),
    .A2(_10161_),
    .A1(_10136_));
 sg13g2_or2_1 _18423_ (.X(_10167_),
    .B(_10166_),
    .A(_10133_));
 sg13g2_a22oi_1 _18424_ (.Y(_10168_),
    .B1(_08108_),
    .B2(\atari2600.tia.diag[32] ),
    .A2(_08107_),
    .A1(\atari2600.tia.diag[33] ));
 sg13g2_a221oi_1 _18425_ (.B2(_07982_),
    .C1(_10168_),
    .B1(net5823),
    .A1(_07983_),
    .Y(_10169_),
    .A2(net5826));
 sg13g2_a221oi_1 _18426_ (.B2(\atari2600.tia.diag[34] ),
    .C1(_10169_),
    .B1(net5562),
    .A1(\atari2600.tia.diag[35] ),
    .Y(_10170_),
    .A2(net5564));
 sg13g2_a221oi_1 _18427_ (.B2(_07980_),
    .C1(_10170_),
    .B1(net5817),
    .A1(_07981_),
    .Y(_10171_),
    .A2(net5822));
 sg13g2_a21oi_1 _18428_ (.A1(\atari2600.tia.diag[36] ),
    .A2(net5560),
    .Y(_10172_),
    .B1(_10171_));
 sg13g2_a21oi_1 _18429_ (.A1(_07979_),
    .A2(net5812),
    .Y(_10173_),
    .B1(_10172_));
 sg13g2_nand2_1 _18430_ (.Y(_10174_),
    .A(_07978_),
    .B(net5808));
 sg13g2_a221oi_1 _18431_ (.B2(\atari2600.tia.diag[38] ),
    .C1(_10173_),
    .B1(net5558),
    .A1(\atari2600.tia.diag[37] ),
    .Y(_10175_),
    .A2(net5559));
 sg13g2_o21ai_1 _18432_ (.B1(_10174_),
    .Y(_10176_),
    .A1(\atari2600.tia.diag[39] ),
    .A2(net5557));
 sg13g2_nand2_1 _18433_ (.Y(_10177_),
    .A(\atari2600.tia.diag[39] ),
    .B(net5557));
 sg13g2_o21ai_1 _18434_ (.B1(\atari2600.tia.enabl ),
    .Y(_10178_),
    .A1(_10175_),
    .A2(_10176_));
 sg13g2_a21oi_1 _18435_ (.A1(net5801),
    .A2(_10132_),
    .Y(_10179_),
    .B1(_10178_));
 sg13g2_nand3_1 _18436_ (.B(_10177_),
    .C(_10179_),
    .A(_10167_),
    .Y(_10180_));
 sg13g2_nor2_2 _18437_ (.A(net5816),
    .B(net5811),
    .Y(_10181_));
 sg13g2_nand2_2 _18438_ (.Y(_10182_),
    .A(net5560),
    .B(net5559));
 sg13g2_a21oi_2 _18439_ (.B1(net5801),
    .Y(_10183_),
    .A2(_10182_),
    .A1(net5806));
 sg13g2_nor2_2 _18440_ (.A(net5806),
    .B(net5557),
    .Y(_10184_));
 sg13g2_a21oi_1 _18441_ (.A1(_08010_),
    .A2(net5816),
    .Y(_10185_),
    .B1(net5811));
 sg13g2_mux2_1 _18442_ (.A0(net5806),
    .A1(_10184_),
    .S(_10185_),
    .X(_10186_));
 sg13g2_a21o_2 _18443_ (.A2(_10183_),
    .A1(_00154_),
    .B1(_10186_),
    .X(_10187_));
 sg13g2_nand2_1 _18444_ (.Y(_10188_),
    .A(_00151_),
    .B(_10183_));
 sg13g2_xor2_1 _18445_ (.B(net5823),
    .A(\atari2600.tia.refpf ),
    .X(_10189_));
 sg13g2_o21ai_1 _18446_ (.B1(_10188_),
    .Y(_10190_),
    .A1(_10183_),
    .A2(_10189_));
 sg13g2_nor2_2 _18447_ (.A(net5807),
    .B(net5802),
    .Y(_10191_));
 sg13g2_nor2_1 _18448_ (.A(net5816),
    .B(_10183_),
    .Y(_10192_));
 sg13g2_a21oi_2 _18449_ (.B1(_10192_),
    .Y(_10193_),
    .A2(_10191_),
    .A1(net5816));
 sg13g2_xor2_1 _18450_ (.B(net5820),
    .A(\atari2600.tia.refpf ),
    .X(_10194_));
 sg13g2_nand2_1 _18451_ (.Y(_10195_),
    .A(net5819),
    .B(_10183_));
 sg13g2_o21ai_1 _18452_ (.B1(_10195_),
    .Y(_10196_),
    .A1(_10183_),
    .A2(_10194_));
 sg13g2_or2_1 _18453_ (.X(_10197_),
    .B(_10183_),
    .A(\atari2600.tia.refpf ));
 sg13g2_nand2_2 _18454_ (.Y(_10198_),
    .A(net5817),
    .B(net5813));
 sg13g2_inv_4 _18455_ (.A(_10198_),
    .Y(_10199_));
 sg13g2_nor2_2 _18456_ (.A(net5560),
    .B(net5813),
    .Y(_10200_));
 sg13g2_nor2_2 _18457_ (.A(net5816),
    .B(net5559),
    .Y(_10201_));
 sg13g2_nor3_1 _18458_ (.A(_10181_),
    .B(_10197_),
    .C(_10199_),
    .Y(_10202_));
 sg13g2_a21oi_2 _18459_ (.B1(_10202_),
    .Y(_10203_),
    .A2(_10197_),
    .A1(net5809));
 sg13g2_mux2_1 _18460_ (.A0(\atari2600.tia.diag[81] ),
    .A1(\atari2600.tia.diag[80] ),
    .S(net5390),
    .X(_10204_));
 sg13g2_a21oi_1 _18461_ (.A1(_07928_),
    .A2(net5391),
    .Y(_10205_),
    .B1(net5389));
 sg13g2_o21ai_1 _18462_ (.B1(_10205_),
    .Y(_10206_),
    .A1(\atari2600.tia.diag[79] ),
    .A2(net5390));
 sg13g2_mux2_1 _18463_ (.A0(\atari2600.tia.diag[77] ),
    .A1(\atari2600.tia.diag[76] ),
    .S(net5390),
    .X(_10207_));
 sg13g2_a21o_1 _18464_ (.A2(_10182_),
    .A1(net5806),
    .B1(_00150_),
    .X(_10208_));
 sg13g2_a21oi_1 _18465_ (.A1(net5557),
    .A2(_00150_),
    .Y(_10209_),
    .B1(\atari2600.tia.refpf ));
 sg13g2_o21ai_1 _18466_ (.B1(net5802),
    .Y(_10210_),
    .A1(net5813),
    .A2(net5805));
 sg13g2_a21oi_2 _18467_ (.B1(net5557),
    .Y(_10211_),
    .A2(net5558),
    .A1(net5559));
 sg13g2_mux2_1 _18468_ (.A0(\atari2600.tia.diag[85] ),
    .A1(\atari2600.tia.diag[84] ),
    .S(net5390),
    .X(_10212_));
 sg13g2_nand2_1 _18469_ (.Y(_10213_),
    .A(net5389),
    .B(_10212_));
 sg13g2_a21oi_1 _18470_ (.A1(_07925_),
    .A2(net5390),
    .Y(_10214_),
    .B1(net5389));
 sg13g2_o21ai_1 _18471_ (.B1(_10214_),
    .Y(_10215_),
    .A1(\atari2600.tia.diag[87] ),
    .A2(net5391));
 sg13g2_and2_1 _18472_ (.A(_10193_),
    .B(_10215_),
    .X(_10216_));
 sg13g2_mux2_1 _18473_ (.A0(\atari2600.tia.diag[91] ),
    .A1(\atari2600.tia.diag[90] ),
    .S(net5390),
    .X(_10217_));
 sg13g2_nand2b_1 _18474_ (.Y(_10218_),
    .B(_10217_),
    .A_N(net5389));
 sg13g2_mux2_1 _18475_ (.A0(\atari2600.tia.diag[89] ),
    .A1(\atari2600.tia.diag[88] ),
    .S(net5391),
    .X(_10219_));
 sg13g2_a21oi_1 _18476_ (.A1(net5389),
    .A2(_10219_),
    .Y(_10220_),
    .B1(_10193_));
 sg13g2_a22oi_1 _18477_ (.Y(_10221_),
    .B1(_10218_),
    .B2(_10220_),
    .A2(_10216_),
    .A1(_10213_));
 sg13g2_nand2_1 _18478_ (.Y(_10222_),
    .A(_10187_),
    .B(_10221_));
 sg13g2_nand2_1 _18479_ (.Y(_10223_),
    .A(_10187_),
    .B(_10193_));
 sg13g2_a21oi_1 _18480_ (.A1(net5389),
    .A2(_10207_),
    .Y(_10224_),
    .B1(_10223_));
 sg13g2_a21oi_1 _18481_ (.A1(_07926_),
    .A2(net5390),
    .Y(_10225_),
    .B1(net5389));
 sg13g2_o21ai_1 _18482_ (.B1(_10225_),
    .Y(_10226_),
    .A1(\atari2600.tia.diag[83] ),
    .A2(net5391));
 sg13g2_a21oi_1 _18483_ (.A1(net5389),
    .A2(_10204_),
    .Y(_10227_),
    .B1(_10193_));
 sg13g2_a22oi_1 _18484_ (.Y(_10228_),
    .B1(_10226_),
    .B2(_10227_),
    .A2(_10224_),
    .A1(_10206_));
 sg13g2_mux4_1 _18485_ (.S0(net5390),
    .A0(\atari2600.tia.diag[95] ),
    .A1(\atari2600.tia.diag[94] ),
    .A2(\atari2600.tia.diag[93] ),
    .A3(\atari2600.tia.diag[92] ),
    .S1(_10196_),
    .X(_10229_));
 sg13g2_a21oi_1 _18486_ (.A1(_10193_),
    .A2(_10229_),
    .Y(_10230_),
    .B1(_10187_));
 sg13g2_a21oi_1 _18487_ (.A1(\atari2600.tia.refpf ),
    .A2(net5474),
    .Y(_10231_),
    .B1(_10230_));
 sg13g2_o21ai_1 _18488_ (.B1(_10231_),
    .Y(_10232_),
    .A1(_10203_),
    .A2(_10228_));
 sg13g2_a221oi_1 _18489_ (.B2(_10203_),
    .C1(_10232_),
    .B1(_10222_),
    .A1(_10208_),
    .Y(_10233_),
    .A2(_10209_));
 sg13g2_nand2_2 _18490_ (.Y(_10234_),
    .A(net5216),
    .B(_10233_));
 sg13g2_inv_1 _18491_ (.Y(_10235_),
    .A(_10234_));
 sg13g2_nand2_1 _18492_ (.Y(_10236_),
    .A(net2918),
    .B(net5197));
 sg13g2_o21ai_1 _18493_ (.B1(_10236_),
    .Y(_00022_),
    .A1(net4766),
    .A2(_10234_));
 sg13g2_nor3_1 _18494_ (.A(_09827_),
    .B(_10052_),
    .C(net4766),
    .Y(_10237_));
 sg13g2_a21o_1 _18495_ (.A2(net5198),
    .A1(net3808),
    .B1(_10237_),
    .X(_00023_));
 sg13g2_a22oi_1 _18496_ (.Y(_10238_),
    .B1(net4768),
    .B2(_10235_),
    .A2(net5197),
    .A1(net2985));
 sg13g2_inv_1 _18497_ (.Y(_00024_),
    .A(_10238_));
 sg13g2_nand2_1 _18498_ (.Y(_10239_),
    .A(net2962),
    .B(net5197));
 sg13g2_o21ai_1 _18499_ (.B1(_10239_),
    .Y(_00025_),
    .A1(_10116_),
    .A2(net4766));
 sg13g2_nand2_1 _18500_ (.Y(_10240_),
    .A(net2933),
    .B(net5197));
 sg13g2_o21ai_1 _18501_ (.B1(_10240_),
    .Y(_00026_),
    .A1(net4784),
    .A2(_10234_));
 sg13g2_nand2_1 _18502_ (.Y(_10241_),
    .A(net2929),
    .B(net5198));
 sg13g2_nand2_2 _18503_ (.Y(_10242_),
    .A(_09821_),
    .B(net5216));
 sg13g2_inv_1 _18504_ (.Y(_10243_),
    .A(_10242_));
 sg13g2_o21ai_1 _18505_ (.B1(_10241_),
    .Y(_00027_),
    .A1(net4766),
    .A2(_10242_));
 sg13g2_nand2_1 _18506_ (.Y(_10244_),
    .A(net2976),
    .B(net5198));
 sg13g2_o21ai_1 _18507_ (.B1(_10244_),
    .Y(_00028_),
    .A1(net4770),
    .A2(_10234_));
 sg13g2_nand2_1 _18508_ (.Y(_10245_),
    .A(net3025),
    .B(net5197));
 sg13g2_o21ai_1 _18509_ (.B1(_10245_),
    .Y(_00029_),
    .A1(_09987_),
    .A2(net4766));
 sg13g2_a22oi_1 _18510_ (.Y(_10246_),
    .B1(net4584),
    .B2(_10235_),
    .A2(net5197),
    .A1(net3037));
 sg13g2_inv_1 _18511_ (.Y(_00016_),
    .A(_10246_));
 sg13g2_a22oi_1 _18512_ (.Y(_10247_),
    .B1(net4768),
    .B2(_10243_),
    .A2(net5198),
    .A1(net3704));
 sg13g2_inv_1 _18513_ (.Y(_00017_),
    .A(_10247_));
 sg13g2_a22oi_1 _18514_ (.Y(_10248_),
    .B1(_09988_),
    .B2(net4768),
    .A2(net5198),
    .A1(net3222));
 sg13g2_inv_1 _18515_ (.Y(_00018_),
    .A(_10248_));
 sg13g2_nand2_1 _18516_ (.Y(_10249_),
    .A(net2991),
    .B(net5198));
 sg13g2_o21ai_1 _18517_ (.B1(_10249_),
    .Y(_00019_),
    .A1(_09987_),
    .A2(net4784));
 sg13g2_nand2_1 _18518_ (.Y(_10250_),
    .A(net2953),
    .B(net5198));
 sg13g2_o21ai_1 _18519_ (.B1(net2954),
    .Y(_00020_),
    .A1(net4784),
    .A2(_10242_));
 sg13g2_nor2_1 _18520_ (.A(net5029),
    .B(_08676_),
    .Y(_10251_));
 sg13g2_nand2_2 _18521_ (.Y(_10252_),
    .A(net5032),
    .B(net4977));
 sg13g2_nand2_2 _18522_ (.Y(_10253_),
    .A(net5039),
    .B(net5026));
 sg13g2_nand4_1 _18523_ (.B(_08605_),
    .C(_08615_),
    .A(net5039),
    .Y(_10254_),
    .D(net5025));
 sg13g2_nor2_1 _18524_ (.A(_10252_),
    .B(_10253_),
    .Y(_10255_));
 sg13g2_nand4_1 _18525_ (.B(_08615_),
    .C(net5224),
    .A(_08605_),
    .Y(_10256_),
    .D(_10255_));
 sg13g2_or2_2 _18526_ (.X(_10257_),
    .B(_10256_),
    .A(\atari2600.tia.vid_vsync ));
 sg13g2_nand2_2 _18527_ (.Y(_10258_),
    .A(net6034),
    .B(net4750));
 sg13g2_nand2_2 _18528_ (.Y(_10259_),
    .A(net5564),
    .B(_08110_));
 sg13g2_and2_2 _18529_ (.A(net5826),
    .B(net5830),
    .X(_10260_));
 sg13g2_nand2_2 _18530_ (.Y(_10261_),
    .A(net5826),
    .B(net5830));
 sg13g2_nand4_1 _18531_ (.B(net5562),
    .C(net5560),
    .A(net5563),
    .Y(_10262_),
    .D(_10261_));
 sg13g2_and4_2 _18532_ (.A(net5810),
    .B(net5804),
    .C(net5800),
    .D(_10262_),
    .X(_10263_));
 sg13g2_nand4_1 _18533_ (.B(net5804),
    .C(net5800),
    .A(net5810),
    .Y(_10264_),
    .D(_10262_));
 sg13g2_nor2_2 _18534_ (.A(_09827_),
    .B(_10263_),
    .Y(_10265_));
 sg13g2_nor2_2 _18535_ (.A(_09658_),
    .B(_10265_),
    .Y(_10266_));
 sg13g2_or2_1 _18536_ (.X(_10267_),
    .B(_10266_),
    .A(net2897));
 sg13g2_nand3_1 _18537_ (.B(net5216),
    .C(_10263_),
    .A(net2897),
    .Y(_10268_));
 sg13g2_o21ai_1 _18538_ (.B1(_10268_),
    .Y(_00038_),
    .A1(_10258_),
    .A2(_10267_));
 sg13g2_nand2_1 _18539_ (.Y(_10269_),
    .A(\atari2600.tia.vid_ypos[1] ),
    .B(\atari2600.tia.vid_ypos[0] ));
 sg13g2_nand3_1 _18540_ (.B(_09826_),
    .C(_10269_),
    .A(_08136_),
    .Y(_10270_));
 sg13g2_a21oi_1 _18541_ (.A1(_10266_),
    .A2(_10270_),
    .Y(_10271_),
    .B1(net2908));
 sg13g2_nand3_1 _18542_ (.B(net4750),
    .C(_10271_),
    .A(net6035),
    .Y(_10272_));
 sg13g2_o21ai_1 _18543_ (.B1(_10272_),
    .Y(_00039_),
    .A1(_10264_),
    .A2(_10270_));
 sg13g2_nand3_1 _18544_ (.B(\atari2600.tia.vid_ypos[1] ),
    .C(\atari2600.tia.vid_ypos[0] ),
    .A(\atari2600.tia.vid_ypos[2] ),
    .Y(_10273_));
 sg13g2_nand2_1 _18545_ (.Y(_10274_),
    .A(_08046_),
    .B(_10269_));
 sg13g2_nand3_1 _18546_ (.B(_10273_),
    .C(_10274_),
    .A(_09826_),
    .Y(_10275_));
 sg13g2_a21oi_1 _18547_ (.A1(_10266_),
    .A2(_10275_),
    .Y(_10276_),
    .B1(net3280));
 sg13g2_nand3_1 _18548_ (.B(net4750),
    .C(_10276_),
    .A(net6034),
    .Y(_10277_));
 sg13g2_o21ai_1 _18549_ (.B1(_10277_),
    .Y(_00040_),
    .A1(_10264_),
    .A2(_10275_));
 sg13g2_nor2_1 _18550_ (.A(net3280),
    .B(_10269_),
    .Y(_10278_));
 sg13g2_xnor2_1 _18551_ (.Y(_10279_),
    .A(\atari2600.tia.vid_ypos[3] ),
    .B(_10278_));
 sg13g2_a21oi_1 _18552_ (.A1(_10263_),
    .A2(_10279_),
    .Y(_10280_),
    .B1(_09827_));
 sg13g2_nor2_1 _18553_ (.A(_09658_),
    .B(_10280_),
    .Y(_10281_));
 sg13g2_nor3_1 _18554_ (.A(net6398),
    .B(_10258_),
    .C(_10281_),
    .Y(_10282_));
 sg13g2_a21o_1 _18555_ (.A2(_10280_),
    .A1(_10263_),
    .B1(_10282_),
    .X(_00041_));
 sg13g2_or2_1 _18556_ (.X(_10283_),
    .B(_10273_),
    .A(_08045_));
 sg13g2_a21oi_1 _18557_ (.A1(_08044_),
    .A2(_10283_),
    .Y(_10284_),
    .B1(_09827_));
 sg13g2_o21ai_1 _18558_ (.B1(_10284_),
    .Y(_10285_),
    .A1(_08044_),
    .A2(_10283_));
 sg13g2_a21oi_1 _18559_ (.A1(_10266_),
    .A2(_10285_),
    .Y(_10286_),
    .B1(net6756));
 sg13g2_nand3_1 _18560_ (.B(net4750),
    .C(_10286_),
    .A(net6034),
    .Y(_10287_));
 sg13g2_o21ai_1 _18561_ (.B1(_10287_),
    .Y(_00042_),
    .A1(_10264_),
    .A2(_10285_));
 sg13g2_nor3_1 _18562_ (.A(\atari2600.tia.vid_ypos[5] ),
    .B(_00051_),
    .C(_10283_),
    .Y(_10288_));
 sg13g2_o21ai_1 _18563_ (.B1(\atari2600.tia.vid_ypos[5] ),
    .Y(_10289_),
    .A1(_00051_),
    .A2(_10283_));
 sg13g2_nand2_1 _18564_ (.Y(_10290_),
    .A(_10263_),
    .B(_10289_));
 sg13g2_o21ai_1 _18565_ (.B1(net5216),
    .Y(_10291_),
    .A1(_10288_),
    .A2(_10290_));
 sg13g2_and2_1 _18566_ (.A(_09659_),
    .B(_10291_),
    .X(_10292_));
 sg13g2_or3_1 _18567_ (.A(net3679),
    .B(_10258_),
    .C(_10292_),
    .X(_10293_));
 sg13g2_o21ai_1 _18568_ (.B1(_10293_),
    .Y(_00043_),
    .A1(_10264_),
    .A2(_10291_));
 sg13g2_or3_2 _18569_ (.A(_08043_),
    .B(_08044_),
    .C(_10283_),
    .X(_10294_));
 sg13g2_a21oi_1 _18570_ (.A1(\atari2600.tia.vid_ypos[6] ),
    .A2(_10294_),
    .Y(_10295_),
    .B1(_10264_));
 sg13g2_o21ai_1 _18571_ (.B1(_10295_),
    .Y(_10296_),
    .A1(\atari2600.tia.vid_ypos[6] ),
    .A2(_10294_));
 sg13g2_nand3_1 _18572_ (.B(_10263_),
    .C(_10296_),
    .A(net5216),
    .Y(_10297_));
 sg13g2_a21oi_1 _18573_ (.A1(_09825_),
    .A2(_10296_),
    .Y(_10298_),
    .B1(_09658_));
 sg13g2_or2_1 _18574_ (.X(_10299_),
    .B(_10298_),
    .A(net6882));
 sg13g2_o21ai_1 _18575_ (.B1(_10297_),
    .Y(_00044_),
    .A1(_10258_),
    .A2(_10299_));
 sg13g2_nor3_1 _18576_ (.A(\atari2600.tia.vid_ypos[7] ),
    .B(_00052_),
    .C(_10294_),
    .Y(_10300_));
 sg13g2_o21ai_1 _18577_ (.B1(\atari2600.tia.vid_ypos[7] ),
    .Y(_10301_),
    .A1(_00052_),
    .A2(_10294_));
 sg13g2_nand2_1 _18578_ (.Y(_10302_),
    .A(_10263_),
    .B(_10301_));
 sg13g2_o21ai_1 _18579_ (.B1(net5216),
    .Y(_10303_),
    .A1(_10300_),
    .A2(_10302_));
 sg13g2_and2_1 _18580_ (.A(_09659_),
    .B(_10303_),
    .X(_10304_));
 sg13g2_or3_1 _18581_ (.A(net2930),
    .B(_10258_),
    .C(_10304_),
    .X(_10305_));
 sg13g2_o21ai_1 _18582_ (.B1(_10305_),
    .Y(_00045_),
    .A1(_10264_),
    .A2(_10303_));
 sg13g2_nand2_1 _18583_ (.Y(_10306_),
    .A(\atari2600.tia.vid_ypos[7] ),
    .B(\atari2600.tia.vid_ypos[6] ));
 sg13g2_nor3_1 _18584_ (.A(\atari2600.tia.vid_ypos[8] ),
    .B(_10294_),
    .C(_10306_),
    .Y(_10307_));
 sg13g2_o21ai_1 _18585_ (.B1(\atari2600.tia.vid_ypos[8] ),
    .Y(_10308_),
    .A1(_10294_),
    .A2(_10306_));
 sg13g2_nand2_1 _18586_ (.Y(_10309_),
    .A(_10263_),
    .B(_10308_));
 sg13g2_o21ai_1 _18587_ (.B1(net5216),
    .Y(_10310_),
    .A1(_10307_),
    .A2(_10309_));
 sg13g2_and2_1 _18588_ (.A(_09659_),
    .B(_10310_),
    .X(_10311_));
 sg13g2_or3_1 _18589_ (.A(net7035),
    .B(_10258_),
    .C(_10311_),
    .X(_10312_));
 sg13g2_o21ai_1 _18590_ (.B1(_10312_),
    .Y(_00046_),
    .A1(_10264_),
    .A2(_10310_));
 sg13g2_nand2_2 _18591_ (.Y(_10313_),
    .A(net6032),
    .B(_09827_));
 sg13g2_nor2_1 _18592_ (.A(net7368),
    .B(_10313_),
    .Y(_10314_));
 sg13g2_a22oi_1 _18593_ (.Y(_10315_),
    .B1(_10314_),
    .B2(net4749),
    .A2(net5113),
    .A1(_08108_));
 sg13g2_inv_1 _18594_ (.Y(_00030_),
    .A(_10315_));
 sg13g2_nor2b_2 _18595_ (.A(net5830),
    .B_N(net5826),
    .Y(_10316_));
 sg13g2_nand2_2 _18596_ (.Y(_10317_),
    .A(net5826),
    .B(_08108_));
 sg13g2_nor2_2 _18597_ (.A(net5826),
    .B(_08108_),
    .Y(_10318_));
 sg13g2_nand2b_2 _18598_ (.Y(_10319_),
    .B(net5830),
    .A_N(net5826));
 sg13g2_o21ai_1 _18599_ (.B1(net5113),
    .Y(_10320_),
    .A1(_10316_),
    .A2(_10318_));
 sg13g2_nor2_1 _18600_ (.A(net7359),
    .B(_10313_),
    .Y(_10321_));
 sg13g2_nand2_1 _18601_ (.Y(_10322_),
    .A(net4749),
    .B(_10321_));
 sg13g2_nand2_1 _18602_ (.Y(_00031_),
    .A(_10320_),
    .B(_10322_));
 sg13g2_nor2_1 _18603_ (.A(_00151_),
    .B(_10313_),
    .Y(_10323_));
 sg13g2_nand2_1 _18604_ (.Y(_10324_),
    .A(net4749),
    .B(_10323_));
 sg13g2_nor2_1 _18605_ (.A(_00151_),
    .B(_10261_),
    .Y(_10325_));
 sg13g2_nand2_1 _18606_ (.Y(_10326_),
    .A(_00151_),
    .B(_10261_));
 sg13g2_nand2_1 _18607_ (.Y(_10327_),
    .A(net5113),
    .B(_10326_));
 sg13g2_o21ai_1 _18608_ (.B1(_10324_),
    .Y(_00032_),
    .A1(_10325_),
    .A2(_10327_));
 sg13g2_xnor2_1 _18609_ (.Y(_10328_),
    .A(net5819),
    .B(_10325_));
 sg13g2_nor2_1 _18610_ (.A(net5819),
    .B(_10313_),
    .Y(_10329_));
 sg13g2_a22oi_1 _18611_ (.Y(_10330_),
    .B1(_10329_),
    .B2(net4749),
    .A2(_10328_),
    .A1(net5113));
 sg13g2_inv_1 _18612_ (.Y(_00033_),
    .A(_10330_));
 sg13g2_nor2_1 _18613_ (.A(net5815),
    .B(_10313_),
    .Y(_10331_));
 sg13g2_nand2_1 _18614_ (.Y(_10332_),
    .A(net5824),
    .B(_10260_));
 sg13g2_nand2_1 _18615_ (.Y(_10333_),
    .A(net5822),
    .B(net5824));
 sg13g2_or2_2 _18616_ (.X(_10334_),
    .B(_10333_),
    .A(_10261_));
 sg13g2_nor2_1 _18617_ (.A(net5815),
    .B(net5472),
    .Y(_10335_));
 sg13g2_xor2_1 _18618_ (.B(net5472),
    .A(net5815),
    .X(_10336_));
 sg13g2_a22oi_1 _18619_ (.Y(_10337_),
    .B1(_10336_),
    .B2(net5113),
    .A2(_10331_),
    .A1(net4749));
 sg13g2_inv_1 _18620_ (.Y(_00034_),
    .A(_10337_));
 sg13g2_xnor2_1 _18621_ (.Y(_10338_),
    .A(net7066),
    .B(_10335_));
 sg13g2_nor2_1 _18622_ (.A(net7066),
    .B(_10313_),
    .Y(_10339_));
 sg13g2_a22oi_1 _18623_ (.Y(_10340_),
    .B1(_10339_),
    .B2(net4749),
    .A2(_10338_),
    .A1(net5113));
 sg13g2_inv_1 _18624_ (.Y(_00035_),
    .A(_10340_));
 sg13g2_nor2_1 _18625_ (.A(net5803),
    .B(_10313_),
    .Y(_10341_));
 sg13g2_nor3_1 _18626_ (.A(net7320),
    .B(_10198_),
    .C(net5472),
    .Y(_10342_));
 sg13g2_o21ai_1 _18627_ (.B1(net7320),
    .Y(_10343_),
    .A1(_10198_),
    .A2(net5472));
 sg13g2_nor2b_1 _18628_ (.A(_10342_),
    .B_N(_10343_),
    .Y(_10344_));
 sg13g2_a22oi_1 _18629_ (.Y(_10345_),
    .B1(_10344_),
    .B2(net5113),
    .A2(_10341_),
    .A1(net4749));
 sg13g2_inv_1 _18630_ (.Y(_00036_),
    .A(_10345_));
 sg13g2_xnor2_1 _18631_ (.Y(_10346_),
    .A(_00150_),
    .B(_10342_));
 sg13g2_nor2_1 _18632_ (.A(net7373),
    .B(_10313_),
    .Y(_10347_));
 sg13g2_a22oi_1 _18633_ (.Y(_10348_),
    .B1(_10347_),
    .B2(net4749),
    .A2(_10346_),
    .A1(net5113));
 sg13g2_inv_1 _18634_ (.Y(_00037_),
    .A(_10348_));
 sg13g2_nor2b_1 _18635_ (.A(\flash_rom.fsm_state[0] ),
    .B_N(\flash_rom.fsm_state[1] ),
    .Y(_10349_));
 sg13g2_nand2_1 _18636_ (.Y(_10350_),
    .A(_07921_),
    .B(\flash_rom.fsm_state[1] ));
 sg13g2_nor2_2 _18637_ (.A(\flash_rom.fsm_state[0] ),
    .B(_10350_),
    .Y(_10351_));
 sg13g2_nor2b_2 _18638_ (.A(\flash_rom.fsm_state[1] ),
    .B_N(\flash_rom.fsm_state[0] ),
    .Y(_10352_));
 sg13g2_nand2_1 _18639_ (.Y(_10353_),
    .A(_00102_),
    .B(_10352_));
 sg13g2_o21ai_1 _18640_ (.B1(\flash_rom.nibbles_remaining[2] ),
    .Y(_10354_),
    .A1(\flash_rom.nibbles_remaining[1] ),
    .A2(\flash_rom.nibbles_remaining[0] ));
 sg13g2_a21oi_1 _18641_ (.A1(\flash_rom.nibbles_remaining[1] ),
    .A2(_07922_),
    .Y(_10355_),
    .B1(\flash_rom.nibbles_remaining[2] ));
 sg13g2_nor2_1 _18642_ (.A(_10353_),
    .B(_10355_),
    .Y(_10356_));
 sg13g2_a22oi_1 _18643_ (.Y(uio_out[1]),
    .B1(_10354_),
    .B2(_10356_),
    .A2(_10351_),
    .A1(_08034_));
 sg13g2_and2_1 _18644_ (.A(\flash_rom.addr[21] ),
    .B(_10351_),
    .X(uio_out[2]));
 sg13g2_and2_1 _18645_ (.A(\flash_rom.addr[22] ),
    .B(_10351_),
    .X(uio_out[4]));
 sg13g2_and2_1 _18646_ (.A(\flash_rom.addr[23] ),
    .B(_10351_),
    .X(uio_out[5]));
 sg13g2_nand2_1 _18647_ (.Y(_00174_),
    .A(_08396_),
    .B(_08430_));
 sg13g2_a221oi_1 _18648_ (.B2(_08252_),
    .C1(_08419_),
    .B1(_08382_),
    .A1(net5315),
    .Y(_10357_),
    .A2(net5437));
 sg13g2_nand4_1 _18649_ (.B(_08403_),
    .C(_08491_),
    .A(_08378_),
    .Y(_00175_),
    .D(_10357_));
 sg13g2_and2_1 _18650_ (.A(_08401_),
    .B(_08425_),
    .X(_10358_));
 sg13g2_nor4_1 _18651_ (.A(_08275_),
    .B(_08321_),
    .C(_08328_),
    .D(_08481_),
    .Y(_10359_));
 sg13g2_and2_1 _18652_ (.A(_08410_),
    .B(_10359_),
    .X(_10360_));
 sg13g2_nand4_1 _18653_ (.B(_08458_),
    .C(_10358_),
    .A(_08439_),
    .Y(_10361_),
    .D(_10360_));
 sg13g2_nor4_1 _18654_ (.A(_08260_),
    .B(_08384_),
    .C(_08465_),
    .D(_10361_),
    .Y(_10362_));
 sg13g2_nand4_1 _18655_ (.B(_08250_),
    .C(_08355_),
    .A(_08220_),
    .Y(_00176_),
    .D(_10362_));
 sg13g2_nand2_1 _18656_ (.Y(_10363_),
    .A(_08412_),
    .B(_08428_));
 sg13g2_nor3_1 _18657_ (.A(_08234_),
    .B(_08272_),
    .C(_08326_),
    .Y(_10364_));
 sg13g2_nor4_1 _18658_ (.A(_08338_),
    .B(_08360_),
    .C(_08468_),
    .D(_08489_),
    .Y(_10365_));
 sg13g2_nand3_1 _18659_ (.B(_10364_),
    .C(_10365_),
    .A(_08390_),
    .Y(_10366_));
 sg13g2_nor4_1 _18660_ (.A(_08318_),
    .B(_08435_),
    .C(_10363_),
    .D(_10366_),
    .Y(_10367_));
 sg13g2_nand3_1 _18661_ (.B(_08462_),
    .C(_10367_),
    .A(_08304_),
    .Y(_10368_));
 sg13g2_nor2_1 _18662_ (.A(_08255_),
    .B(_10368_),
    .Y(_10369_));
 sg13g2_nand4_1 _18663_ (.B(_08406_),
    .C(_08456_),
    .A(_08398_),
    .Y(_00177_),
    .D(_10369_));
 sg13g2_and2_1 _18664_ (.A(net6733),
    .B(\atari2600.cpu.adc_sbc ),
    .X(_00014_));
 sg13g2_nor2_2 _18665_ (.A(net5822),
    .B(net5562),
    .Y(_10370_));
 sg13g2_nand2_2 _18666_ (.Y(_10371_),
    .A(net5564),
    .B(net5824));
 sg13g2_nor2_2 _18667_ (.A(_10319_),
    .B(_10371_),
    .Y(_10372_));
 sg13g2_nand2_2 _18668_ (.Y(_10373_),
    .A(_10318_),
    .B(_10370_));
 sg13g2_nor2_2 _18669_ (.A(net5558),
    .B(net5801),
    .Y(_10374_));
 sg13g2_nand2_2 _18670_ (.Y(_10375_),
    .A(net5806),
    .B(net5557));
 sg13g2_nor2_2 _18671_ (.A(_10182_),
    .B(_10375_),
    .Y(_10376_));
 sg13g2_nand2_2 _18672_ (.Y(_10377_),
    .A(_10181_),
    .B(_10374_));
 sg13g2_nand2_2 _18673_ (.Y(_10378_),
    .A(_10372_),
    .B(net5432));
 sg13g2_mux2_1 _18674_ (.A0(net5773),
    .A1(net6590),
    .S(_10378_),
    .X(_00179_));
 sg13g2_mux2_1 _18675_ (.A0(net5745),
    .A1(net4476),
    .S(_10378_),
    .X(_00180_));
 sg13g2_mux2_1 _18676_ (.A0(net5717),
    .A1(net6192),
    .S(_10378_),
    .X(_00181_));
 sg13g2_mux2_1 _18677_ (.A0(net5689),
    .A1(net6605),
    .S(_10378_),
    .X(_00182_));
 sg13g2_mux2_1 _18678_ (.A0(net5658),
    .A1(net6630),
    .S(_10378_),
    .X(_00183_));
 sg13g2_mux2_1 _18679_ (.A0(net5628),
    .A1(net4538),
    .S(_10378_),
    .X(_00184_));
 sg13g2_mux2_1 _18680_ (.A0(net5601),
    .A1(net6064),
    .S(_10378_),
    .X(_00185_));
 sg13g2_nor2_2 _18681_ (.A(net5564),
    .B(net5824),
    .Y(_10379_));
 sg13g2_nand2_2 _18682_ (.Y(_10380_),
    .A(net5822),
    .B(net5562));
 sg13g2_nor2_2 _18683_ (.A(_10317_),
    .B(_10380_),
    .Y(_10381_));
 sg13g2_nand2_2 _18684_ (.Y(_10382_),
    .A(_10316_),
    .B(_10379_));
 sg13g2_and2_2 _18685_ (.A(_10184_),
    .B(_10200_),
    .X(_10383_));
 sg13g2_nand2_2 _18686_ (.Y(_10384_),
    .A(_10184_),
    .B(_10200_));
 sg13g2_nor2_2 _18687_ (.A(_10382_),
    .B(net5430),
    .Y(_10385_));
 sg13g2_mux2_1 _18688_ (.A0(net3308),
    .A1(net5776),
    .S(_10385_),
    .X(_00186_));
 sg13g2_mux2_1 _18689_ (.A0(net3850),
    .A1(net5750),
    .S(_10385_),
    .X(_00187_));
 sg13g2_mux2_1 _18690_ (.A0(net3293),
    .A1(net5720),
    .S(_10385_),
    .X(_00188_));
 sg13g2_mux2_1 _18691_ (.A0(net3560),
    .A1(net5691),
    .S(_10385_),
    .X(_00189_));
 sg13g2_mux2_1 _18692_ (.A0(net3751),
    .A1(net5662),
    .S(_10385_),
    .X(_00190_));
 sg13g2_mux2_1 _18693_ (.A0(net3873),
    .A1(net5636),
    .S(_10385_),
    .X(_00191_));
 sg13g2_mux2_1 _18694_ (.A0(net3867),
    .A1(net5604),
    .S(_10385_),
    .X(_00192_));
 sg13g2_xnor2_1 _18695_ (.Y(_10386_),
    .A(\rom_last_read_addr[2] ),
    .B(net5032));
 sg13g2_a22oi_1 _18696_ (.Y(_10387_),
    .B1(_08592_),
    .B2(\atari2600.cpu.ABH[2] ),
    .A2(net5396),
    .A1(net5571));
 sg13g2_o21ai_1 _18697_ (.B1(_10387_),
    .Y(_10388_),
    .A1(_08201_),
    .A2(_08527_));
 sg13g2_mux2_2 _18698_ (.A0(\atari2600.cpu.PC[10] ),
    .A1(_10388_),
    .S(net5309),
    .X(_10389_));
 sg13g2_mux2_2 _18699_ (.A0(net7195),
    .A1(_10389_),
    .S(net5353),
    .X(_10390_));
 sg13g2_xnor2_1 _18700_ (.Y(_10391_),
    .A(\rom_last_read_addr[10] ),
    .B(_10390_));
 sg13g2_o21ai_1 _18701_ (.B1(_10391_),
    .Y(_10392_),
    .A1(\rom_last_read_addr[5] ),
    .A2(net4877));
 sg13g2_xnor2_1 _18702_ (.Y(_10393_),
    .A(\rom_last_read_addr[1] ),
    .B(net5035));
 sg13g2_a22oi_1 _18703_ (.Y(_10394_),
    .B1(_08592_),
    .B2(\atari2600.cpu.ABH[0] ),
    .A2(net5396),
    .A1(net5572));
 sg13g2_o21ai_1 _18704_ (.B1(_10394_),
    .Y(_10395_),
    .A1(_08191_),
    .A2(_08527_));
 sg13g2_mux2_2 _18705_ (.A0(\atari2600.cpu.PC[8] ),
    .A1(_10395_),
    .S(net5307),
    .X(_10396_));
 sg13g2_mux2_2 _18706_ (.A0(net7335),
    .A1(_10396_),
    .S(net5353),
    .X(_10397_));
 sg13g2_inv_1 _18707_ (.Y(_10398_),
    .A(_10397_));
 sg13g2_a22oi_1 _18708_ (.Y(_10399_),
    .B1(_08592_),
    .B2(\atari2600.cpu.ABH[1] ),
    .A2(net5396),
    .A1(\atari2600.cpu.ADD[1] ));
 sg13g2_o21ai_1 _18709_ (.B1(_10399_),
    .Y(_10400_),
    .A1(_08187_),
    .A2(_08527_));
 sg13g2_mux2_1 _18710_ (.A0(\atari2600.cpu.PC[9] ),
    .A1(_10400_),
    .S(net5307),
    .X(_10401_));
 sg13g2_nor2_2 _18711_ (.A(net5316),
    .B(_10401_),
    .Y(_10402_));
 sg13g2_a21oi_2 _18712_ (.B1(_10402_),
    .Y(_10403_),
    .A2(net5316),
    .A1(_08084_));
 sg13g2_inv_1 _18713_ (.Y(_10404_),
    .A(_10403_));
 sg13g2_a22oi_1 _18714_ (.Y(_10405_),
    .B1(_10404_),
    .B2(\rom_last_read_addr[9] ),
    .A2(_10398_),
    .A1(\rom_last_read_addr[8] ));
 sg13g2_a22oi_1 _18715_ (.Y(_10406_),
    .B1(_10403_),
    .B2(_08085_),
    .A2(_10397_),
    .A1(_08083_));
 sg13g2_nand3_1 _18716_ (.B(_10405_),
    .C(_10406_),
    .A(_10393_),
    .Y(_10407_));
 sg13g2_xnor2_1 _18717_ (.Y(_10408_),
    .A(\rom_last_read_addr[6] ),
    .B(net5024));
 sg13g2_a22oi_1 _18718_ (.Y(_10409_),
    .B1(_08592_),
    .B2(\atari2600.cpu.ABH[3] ),
    .A2(net5396),
    .A1(\atari2600.cpu.ADD[3] ));
 sg13g2_o21ai_1 _18719_ (.B1(_10409_),
    .Y(_10410_),
    .A1(_08196_),
    .A2(_08527_));
 sg13g2_mux2_2 _18720_ (.A0(\atari2600.cpu.PC[11] ),
    .A1(_10410_),
    .S(net5307),
    .X(_10411_));
 sg13g2_mux2_2 _18721_ (.A0(net7185),
    .A1(_10411_),
    .S(net5353),
    .X(_10412_));
 sg13g2_xnor2_1 _18722_ (.Y(_10413_),
    .A(\rom_last_read_addr[11] ),
    .B(_10412_));
 sg13g2_o21ai_1 _18723_ (.B1(_10413_),
    .Y(_10414_),
    .A1(\rom_last_read_addr[3] ),
    .A2(net5037));
 sg13g2_nor2_1 _18724_ (.A(_10408_),
    .B(_10414_),
    .Y(_10415_));
 sg13g2_a22oi_1 _18725_ (.Y(_10416_),
    .B1(net5026),
    .B2(\rom_last_read_addr[4] ),
    .A2(net4877),
    .A1(\rom_last_read_addr[5] ));
 sg13g2_a21oi_2 _18726_ (.B1(_08634_),
    .Y(_10417_),
    .A2(net5316),
    .A1(_08081_));
 sg13g2_xnor2_1 _18727_ (.Y(_10418_),
    .A(\rom_last_read_addr[7] ),
    .B(_10417_));
 sg13g2_nand2b_1 _18728_ (.Y(_10419_),
    .B(net5034),
    .A_N(\rom_last_read_addr[0] ));
 sg13g2_o21ai_1 _18729_ (.B1(_10419_),
    .Y(_10420_),
    .A1(\rom_last_read_addr[4] ),
    .A2(net5026));
 sg13g2_a221oi_1 _18730_ (.B2(\rom_last_read_addr[0] ),
    .C1(_10420_),
    .B1(_08563_),
    .A1(\rom_last_read_addr[3] ),
    .Y(_10421_),
    .A2(net5037));
 sg13g2_nand4_1 _18731_ (.B(_10416_),
    .C(_10418_),
    .A(_10415_),
    .Y(_10422_),
    .D(_10421_));
 sg13g2_nor4_1 _18732_ (.A(_10386_),
    .B(_10392_),
    .C(_10407_),
    .D(_10422_),
    .Y(_10423_));
 sg13g2_o21ai_1 _18733_ (.B1(_08596_),
    .Y(_10424_),
    .A1(\atari2600.address_bus_r[12] ),
    .A2(net5353));
 sg13g2_inv_1 _18734_ (.Y(_10425_),
    .A(net4781));
 sg13g2_xnor2_1 _18735_ (.Y(_10426_),
    .A(\rom_next_addr_in_queue[7] ),
    .B(_10417_));
 sg13g2_xnor2_1 _18736_ (.Y(_10427_),
    .A(_08092_),
    .B(net5027));
 sg13g2_xnor2_1 _18737_ (.Y(_10428_),
    .A(_00105_),
    .B(net5034));
 sg13g2_xnor2_1 _18738_ (.Y(_10429_),
    .A(\rom_next_addr_in_queue[9] ),
    .B(_10403_));
 sg13g2_xnor2_1 _18739_ (.Y(_10430_),
    .A(\rom_next_addr_in_queue[8] ),
    .B(_10397_));
 sg13g2_xnor2_1 _18740_ (.Y(_10431_),
    .A(_08095_),
    .B(_10412_));
 sg13g2_xnor2_1 _18741_ (.Y(_10432_),
    .A(\rom_next_addr_in_queue[10] ),
    .B(_10390_));
 sg13g2_xnor2_1 _18742_ (.Y(_10433_),
    .A(_08089_),
    .B(net5035));
 sg13g2_nor3_1 _18743_ (.A(_10427_),
    .B(_10431_),
    .C(_10433_),
    .Y(_10434_));
 sg13g2_xnor2_1 _18744_ (.Y(_10435_),
    .A(\rom_next_addr_in_queue[6] ),
    .B(net5024));
 sg13g2_nor2_1 _18745_ (.A(_10428_),
    .B(_10435_),
    .Y(_10436_));
 sg13g2_a22oi_1 _18746_ (.Y(_10437_),
    .B1(net5029),
    .B2(_08090_),
    .A2(net5036),
    .A1(_08091_));
 sg13g2_nand4_1 _18747_ (.B(_10434_),
    .C(_10436_),
    .A(_10429_),
    .Y(_10438_),
    .D(_10437_));
 sg13g2_a22oi_1 _18748_ (.Y(_10439_),
    .B1(net4877),
    .B2(\rom_next_addr_in_queue[5] ),
    .A2(net5037),
    .A1(\rom_next_addr_in_queue[3] ));
 sg13g2_o21ai_1 _18749_ (.B1(_10439_),
    .Y(_10440_),
    .A1(\rom_next_addr_in_queue[5] ),
    .A2(net4877));
 sg13g2_a21oi_1 _18750_ (.A1(\rom_next_addr_in_queue[2] ),
    .A2(net5032),
    .Y(_10441_),
    .B1(_10440_));
 sg13g2_nand4_1 _18751_ (.B(_10430_),
    .C(_10432_),
    .A(_10426_),
    .Y(_10442_),
    .D(_10441_));
 sg13g2_nor2_1 _18752_ (.A(_10438_),
    .B(_10442_),
    .Y(_10443_));
 sg13g2_or4_1 _18753_ (.A(net5315),
    .B(_10423_),
    .C(_10424_),
    .D(_10443_),
    .X(_10444_));
 sg13g2_nor2b_1 _18754_ (.A(spi_restart),
    .B_N(_10444_),
    .Y(_10445_));
 sg13g2_nor2b_1 _18755_ (.A(_10445_),
    .B_N(net5537),
    .Y(_10446_));
 sg13g2_nor3_1 _18756_ (.A(\flash_rom.fsm_state[0] ),
    .B(_00137_),
    .C(_10350_),
    .Y(_10447_));
 sg13g2_nand2b_1 _18757_ (.Y(_10448_),
    .B(_10351_),
    .A_N(_00137_));
 sg13g2_nor2_2 _18758_ (.A(net4566),
    .B(net5426),
    .Y(_10449_));
 sg13g2_a22oi_1 _18759_ (.Y(_10450_),
    .B1(_10449_),
    .B2(net2967),
    .A2(net4566),
    .A1(net5034));
 sg13g2_inv_1 _18760_ (.Y(_00193_),
    .A(_10450_));
 sg13g2_a22oi_1 _18761_ (.Y(_10451_),
    .B1(_10449_),
    .B2(net2911),
    .A2(net4566),
    .A1(net5035));
 sg13g2_inv_1 _18762_ (.Y(_00194_),
    .A(_10451_));
 sg13g2_a22oi_1 _18763_ (.Y(_10452_),
    .B1(_10449_),
    .B2(net2925),
    .A2(net4564),
    .A1(net5029));
 sg13g2_inv_1 _18764_ (.Y(_00195_),
    .A(_10452_));
 sg13g2_a22oi_1 _18765_ (.Y(_10453_),
    .B1(_10449_),
    .B2(net2920),
    .A2(net4564),
    .A1(net5036));
 sg13g2_inv_1 _18766_ (.Y(_00196_),
    .A(_10453_));
 sg13g2_nand2_1 _18767_ (.Y(_10454_),
    .A(net5027),
    .B(net4568));
 sg13g2_or2_1 _18768_ (.X(_10455_),
    .B(net5426),
    .A(net7110));
 sg13g2_o21ai_1 _18769_ (.B1(_10455_),
    .Y(_10456_),
    .A1(net2967),
    .A2(net5393));
 sg13g2_o21ai_1 _18770_ (.B1(_10454_),
    .Y(_00197_),
    .A1(net4566),
    .A2(_10456_));
 sg13g2_nand2b_1 _18771_ (.Y(_10457_),
    .B(net4568),
    .A_N(net4877));
 sg13g2_or2_1 _18772_ (.X(_10458_),
    .B(net5426),
    .A(net7220));
 sg13g2_o21ai_1 _18773_ (.B1(_10458_),
    .Y(_10459_),
    .A1(net2911),
    .A2(net5393));
 sg13g2_o21ai_1 _18774_ (.B1(_10457_),
    .Y(_00198_),
    .A1(net4566),
    .A2(_10459_));
 sg13g2_nand2_1 _18775_ (.Y(_10460_),
    .A(net5022),
    .B(net4564));
 sg13g2_or2_1 _18776_ (.X(_10461_),
    .B(net5426),
    .A(net7175));
 sg13g2_o21ai_1 _18777_ (.B1(_10461_),
    .Y(_10462_),
    .A1(net2925),
    .A2(net5393));
 sg13g2_o21ai_1 _18778_ (.B1(_10460_),
    .Y(_00199_),
    .A1(net4564),
    .A2(_10462_));
 sg13g2_nand2_1 _18779_ (.Y(_10463_),
    .A(_10417_),
    .B(net4564));
 sg13g2_or2_1 _18780_ (.X(_10464_),
    .B(net5426),
    .A(net7140));
 sg13g2_o21ai_1 _18781_ (.B1(_10464_),
    .Y(_10465_),
    .A1(net2920),
    .A2(net5393));
 sg13g2_o21ai_1 _18782_ (.B1(_10463_),
    .Y(_00200_),
    .A1(net4565),
    .A2(_10465_));
 sg13g2_nand2_1 _18783_ (.Y(_10466_),
    .A(_10397_),
    .B(net4565));
 sg13g2_or2_1 _18784_ (.X(_10467_),
    .B(net5426),
    .A(\flash_rom.addr[8] ));
 sg13g2_o21ai_1 _18785_ (.B1(_10467_),
    .Y(_10468_),
    .A1(net7110),
    .A2(net5393));
 sg13g2_o21ai_1 _18786_ (.B1(_10466_),
    .Y(_00201_),
    .A1(net4569),
    .A2(net7111));
 sg13g2_nand2_1 _18787_ (.Y(_10469_),
    .A(_10403_),
    .B(net4566));
 sg13g2_or2_1 _18788_ (.X(_10470_),
    .B(net5427),
    .A(net3021));
 sg13g2_o21ai_1 _18789_ (.B1(_10470_),
    .Y(_10471_),
    .A1(net7220),
    .A2(net5393));
 sg13g2_o21ai_1 _18790_ (.B1(_10469_),
    .Y(_00202_),
    .A1(net4569),
    .A2(_10471_));
 sg13g2_nand2_1 _18791_ (.Y(_10472_),
    .A(_10390_),
    .B(net4564));
 sg13g2_or2_1 _18792_ (.X(_10473_),
    .B(net5426),
    .A(net4066));
 sg13g2_o21ai_1 _18793_ (.B1(_10473_),
    .Y(_10474_),
    .A1(net7175),
    .A2(net5393));
 sg13g2_o21ai_1 _18794_ (.B1(_10472_),
    .Y(_00203_),
    .A1(net4564),
    .A2(_10474_));
 sg13g2_nand2_1 _18795_ (.Y(_10475_),
    .A(_10412_),
    .B(net4565));
 sg13g2_or2_1 _18796_ (.X(_10476_),
    .B(net5426),
    .A(net3846));
 sg13g2_o21ai_1 _18797_ (.B1(_10476_),
    .Y(_10477_),
    .A1(net7140),
    .A2(net5393));
 sg13g2_o21ai_1 _18798_ (.B1(_10475_),
    .Y(_00204_),
    .A1(net4565),
    .A2(_10477_));
 sg13g2_nor2_2 _18799_ (.A(_10261_),
    .B(_10380_),
    .Y(_10478_));
 sg13g2_nand2_2 _18800_ (.Y(_10479_),
    .A(_10260_),
    .B(_10379_));
 sg13g2_nor3_2 _18801_ (.A(net5807),
    .B(net5801),
    .C(_10198_),
    .Y(_10480_));
 sg13g2_nand2_2 _18802_ (.Y(_10481_),
    .A(_10191_),
    .B(_10199_));
 sg13g2_nor2_2 _18803_ (.A(_10479_),
    .B(net5425),
    .Y(_10482_));
 sg13g2_mux2_1 _18804_ (.A0(net3612),
    .A1(net5790),
    .S(_10482_),
    .X(_00205_));
 sg13g2_mux2_1 _18805_ (.A0(net3401),
    .A1(net5756),
    .S(_10482_),
    .X(_00206_));
 sg13g2_mux2_1 _18806_ (.A0(net3619),
    .A1(net5723),
    .S(_10482_),
    .X(_00207_));
 sg13g2_mux2_1 _18807_ (.A0(net3536),
    .A1(net5694),
    .S(_10482_),
    .X(_00208_));
 sg13g2_mux2_1 _18808_ (.A0(net3831),
    .A1(net5665),
    .S(_10482_),
    .X(_00209_));
 sg13g2_mux2_1 _18809_ (.A0(net3658),
    .A1(net5640),
    .S(_10482_),
    .X(_00210_));
 sg13g2_mux2_1 _18810_ (.A0(net3311),
    .A1(net5614),
    .S(_10482_),
    .X(_00211_));
 sg13g2_nor2_1 _18811_ (.A(net4165),
    .B(net5394),
    .Y(_10483_));
 sg13g2_nor2_1 _18812_ (.A(net4221),
    .B(net5428),
    .Y(_10484_));
 sg13g2_nor3_1 _18813_ (.A(net4571),
    .B(_10483_),
    .C(_10484_),
    .Y(_00212_));
 sg13g2_nor2_1 _18814_ (.A(\flash_rom.addr[13] ),
    .B(net5394),
    .Y(_10485_));
 sg13g2_nor2_1 _18815_ (.A(net4009),
    .B(net5428),
    .Y(_10486_));
 sg13g2_nor3_1 _18816_ (.A(net4571),
    .B(_10485_),
    .C(_10486_),
    .Y(_00213_));
 sg13g2_nor2_1 _18817_ (.A(net3646),
    .B(net5394),
    .Y(_10487_));
 sg13g2_nor2_1 _18818_ (.A(\flash_rom.addr[18] ),
    .B(net5428),
    .Y(_10488_));
 sg13g2_nor3_1 _18819_ (.A(net4570),
    .B(_10487_),
    .C(_10488_),
    .Y(_00214_));
 sg13g2_nor2_1 _18820_ (.A(net3952),
    .B(net5394),
    .Y(_10489_));
 sg13g2_nor2_1 _18821_ (.A(net3707),
    .B(net5428),
    .Y(_10490_));
 sg13g2_nor3_1 _18822_ (.A(net4570),
    .B(_10489_),
    .C(_10490_),
    .Y(_00215_));
 sg13g2_nor2_1 _18823_ (.A(net4009),
    .B(net5395),
    .Y(_10491_));
 sg13g2_nor2_1 _18824_ (.A(net4215),
    .B(net5429),
    .Y(_10492_));
 sg13g2_nor3_1 _18825_ (.A(net4570),
    .B(_10491_),
    .C(net4216),
    .Y(_00216_));
 sg13g2_nor2_1 _18826_ (.A(\flash_rom.addr[18] ),
    .B(net5395),
    .Y(_10493_));
 sg13g2_nor2_1 _18827_ (.A(net3710),
    .B(net5428),
    .Y(_10494_));
 sg13g2_nor3_1 _18828_ (.A(net4570),
    .B(_10493_),
    .C(_10494_),
    .Y(_00217_));
 sg13g2_nor2_1 _18829_ (.A(net3707),
    .B(net5394),
    .Y(_10495_));
 sg13g2_nor2_1 _18830_ (.A(\flash_rom.addr[23] ),
    .B(net5428),
    .Y(_10496_));
 sg13g2_nor3_1 _18831_ (.A(net4571),
    .B(_10495_),
    .C(_10496_),
    .Y(_00218_));
 sg13g2_nor3_2 _18832_ (.A(net5827),
    .B(net5831),
    .C(_10259_),
    .Y(_10497_));
 sg13g2_and2_1 _18833_ (.A(_10191_),
    .B(_10201_),
    .X(_10498_));
 sg13g2_nand2_2 _18834_ (.Y(_10499_),
    .A(_10191_),
    .B(_10201_));
 sg13g2_nand2_2 _18835_ (.Y(_10500_),
    .A(net5424),
    .B(net5423));
 sg13g2_mux2_1 _18836_ (.A0(net5789),
    .A1(net6264),
    .S(_10500_),
    .X(_00219_));
 sg13g2_mux2_1 _18837_ (.A0(net5755),
    .A1(net6965),
    .S(_10500_),
    .X(_00220_));
 sg13g2_mux2_1 _18838_ (.A0(net5723),
    .A1(net6507),
    .S(_10500_),
    .X(_00221_));
 sg13g2_mux2_1 _18839_ (.A0(net5694),
    .A1(net6140),
    .S(_10500_),
    .X(_00222_));
 sg13g2_mux2_1 _18840_ (.A0(net5665),
    .A1(net6371),
    .S(_10500_),
    .X(_00223_));
 sg13g2_mux2_1 _18841_ (.A0(net5640),
    .A1(net6740),
    .S(_10500_),
    .X(_00224_));
 sg13g2_mux2_1 _18842_ (.A0(net5608),
    .A1(net6451),
    .S(_10500_),
    .X(_00225_));
 sg13g2_and2_1 _18843_ (.A(_10191_),
    .B(_10200_),
    .X(_10501_));
 sg13g2_nand2_2 _18844_ (.Y(_10502_),
    .A(_10191_),
    .B(_10200_));
 sg13g2_nor2_2 _18845_ (.A(net5473),
    .B(_10502_),
    .Y(_10503_));
 sg13g2_mux2_1 _18846_ (.A0(net3555),
    .A1(net5784),
    .S(_10503_),
    .X(_00226_));
 sg13g2_mux2_1 _18847_ (.A0(net3561),
    .A1(net5763),
    .S(_10503_),
    .X(_00227_));
 sg13g2_mux2_1 _18848_ (.A0(net3842),
    .A1(net5730),
    .S(_10503_),
    .X(_00228_));
 sg13g2_mux2_1 _18849_ (.A0(net3578),
    .A1(net5703),
    .S(_10503_),
    .X(_00229_));
 sg13g2_mux2_1 _18850_ (.A0(net3937),
    .A1(net5675),
    .S(_10503_),
    .X(_00230_));
 sg13g2_mux2_1 _18851_ (.A0(net3450),
    .A1(net5642),
    .S(_10503_),
    .X(_00231_));
 sg13g2_mux2_1 _18852_ (.A0(net3843),
    .A1(net5617),
    .S(_10503_),
    .X(_00232_));
 sg13g2_nand3_1 _18853_ (.B(net5823),
    .C(_10316_),
    .A(net5822),
    .Y(_10504_));
 sg13g2_nor2_2 _18854_ (.A(_10502_),
    .B(_10504_),
    .Y(_10505_));
 sg13g2_mux2_1 _18855_ (.A0(net3919),
    .A1(net5787),
    .S(_10505_),
    .X(_00233_));
 sg13g2_mux2_1 _18856_ (.A0(net3460),
    .A1(net5763),
    .S(_10505_),
    .X(_00234_));
 sg13g2_mux2_1 _18857_ (.A0(net3690),
    .A1(net5730),
    .S(_10505_),
    .X(_00235_));
 sg13g2_mux2_1 _18858_ (.A0(net3303),
    .A1(net5703),
    .S(_10505_),
    .X(_00236_));
 sg13g2_mux2_1 _18859_ (.A0(net3187),
    .A1(net5675),
    .S(_10505_),
    .X(_00237_));
 sg13g2_mux2_1 _18860_ (.A0(net3664),
    .A1(net5642),
    .S(_10505_),
    .X(_00238_));
 sg13g2_mux2_1 _18861_ (.A0(net3641),
    .A1(net5616),
    .S(_10505_),
    .X(_00239_));
 sg13g2_and2_1 _18862_ (.A(_10181_),
    .B(_10191_),
    .X(_10506_));
 sg13g2_nor2_2 _18863_ (.A(_10259_),
    .B(_10317_),
    .Y(_10507_));
 sg13g2_nand2_2 _18864_ (.Y(_10508_),
    .A(net5470),
    .B(_10507_));
 sg13g2_mux2_1 _18865_ (.A0(net5787),
    .A1(net6529),
    .S(_10508_),
    .X(_00240_));
 sg13g2_mux2_1 _18866_ (.A0(net5754),
    .A1(net6436),
    .S(_10508_),
    .X(_00241_));
 sg13g2_mux2_1 _18867_ (.A0(net5725),
    .A1(net6728),
    .S(_10508_),
    .X(_00242_));
 sg13g2_mux2_1 _18868_ (.A0(net5705),
    .A1(net6750),
    .S(_10508_),
    .X(_00243_));
 sg13g2_mux2_1 _18869_ (.A0(net5668),
    .A1(net6762),
    .S(_10508_),
    .X(_00244_));
 sg13g2_mux2_1 _18870_ (.A0(net5641),
    .A1(net6565),
    .S(_10508_),
    .X(_00245_));
 sg13g2_mux2_1 _18871_ (.A0(net5609),
    .A1(net4502),
    .S(_10508_),
    .X(_00246_));
 sg13g2_nor3_2 _18872_ (.A(net5827),
    .B(net5830),
    .C(_10333_),
    .Y(_10509_));
 sg13g2_nand2_2 _18873_ (.Y(_10510_),
    .A(net5420),
    .B(net5468));
 sg13g2_mux2_1 _18874_ (.A0(net5788),
    .A1(net4246),
    .S(_10510_),
    .X(_00247_));
 sg13g2_mux2_1 _18875_ (.A0(net5763),
    .A1(net6559),
    .S(_10510_),
    .X(_00248_));
 sg13g2_mux2_1 _18876_ (.A0(net5730),
    .A1(net6386),
    .S(_10510_),
    .X(_00249_));
 sg13g2_mux2_1 _18877_ (.A0(net5702),
    .A1(net6211),
    .S(_10510_),
    .X(_00250_));
 sg13g2_mux2_1 _18878_ (.A0(net5675),
    .A1(net6440),
    .S(_10510_),
    .X(_00251_));
 sg13g2_mux2_1 _18879_ (.A0(net5642),
    .A1(net4399),
    .S(_10510_),
    .X(_00252_));
 sg13g2_mux2_1 _18880_ (.A0(net5616),
    .A1(net4407),
    .S(_10510_),
    .X(_00253_));
 sg13g2_nand2_2 _18881_ (.Y(_10511_),
    .A(_10478_),
    .B(net5420));
 sg13g2_mux2_1 _18882_ (.A0(net5784),
    .A1(net6506),
    .S(_10511_),
    .X(_00254_));
 sg13g2_mux2_1 _18883_ (.A0(net5761),
    .A1(net6870),
    .S(_10511_),
    .X(_00255_));
 sg13g2_mux2_1 _18884_ (.A0(net5730),
    .A1(net6573),
    .S(_10511_),
    .X(_00256_));
 sg13g2_mux2_1 _18885_ (.A0(net5702),
    .A1(net6480),
    .S(_10511_),
    .X(_00257_));
 sg13g2_mux2_1 _18886_ (.A0(net5675),
    .A1(net6925),
    .S(_10511_),
    .X(_00258_));
 sg13g2_mux2_1 _18887_ (.A0(net5642),
    .A1(net6887),
    .S(_10511_),
    .X(_00259_));
 sg13g2_mux2_1 _18888_ (.A0(net5616),
    .A1(net6845),
    .S(_10511_),
    .X(_00260_));
 sg13g2_nand2_2 _18889_ (.Y(_10512_),
    .A(_10381_),
    .B(net5420));
 sg13g2_mux2_1 _18890_ (.A0(net5784),
    .A1(net6592),
    .S(_10512_),
    .X(_00261_));
 sg13g2_mux2_1 _18891_ (.A0(net5761),
    .A1(net6183),
    .S(_10512_),
    .X(_00262_));
 sg13g2_mux2_1 _18892_ (.A0(net5730),
    .A1(net6695),
    .S(_10512_),
    .X(_00263_));
 sg13g2_mux2_1 _18893_ (.A0(net5702),
    .A1(net6093),
    .S(_10512_),
    .X(_00264_));
 sg13g2_mux2_1 _18894_ (.A0(net5675),
    .A1(net6577),
    .S(_10512_),
    .X(_00265_));
 sg13g2_mux2_1 _18895_ (.A0(net5642),
    .A1(net6675),
    .S(_10512_),
    .X(_00266_));
 sg13g2_mux2_1 _18896_ (.A0(net5616),
    .A1(net6856),
    .S(_10512_),
    .X(_00267_));
 sg13g2_nor2_2 _18897_ (.A(_10319_),
    .B(_10380_),
    .Y(_02995_));
 sg13g2_nand2_2 _18898_ (.Y(_02996_),
    .A(_10318_),
    .B(_10379_));
 sg13g2_nand2_2 _18899_ (.Y(_02997_),
    .A(net5420),
    .B(_02995_));
 sg13g2_mux2_1 _18900_ (.A0(net5785),
    .A1(net4506),
    .S(_02997_),
    .X(_00268_));
 sg13g2_mux2_1 _18901_ (.A0(net5761),
    .A1(net4289),
    .S(_02997_),
    .X(_00269_));
 sg13g2_mux2_1 _18902_ (.A0(net5730),
    .A1(net4510),
    .S(_02997_),
    .X(_00270_));
 sg13g2_mux2_1 _18903_ (.A0(net5702),
    .A1(net6450),
    .S(_02997_),
    .X(_00271_));
 sg13g2_mux2_1 _18904_ (.A0(net5675),
    .A1(net6923),
    .S(_02997_),
    .X(_00272_));
 sg13g2_mux2_1 _18905_ (.A0(net5642),
    .A1(net4282),
    .S(_02997_),
    .X(_00273_));
 sg13g2_mux2_1 _18906_ (.A0(net5616),
    .A1(net6300),
    .S(_02997_),
    .X(_00274_));
 sg13g2_or2_2 _18907_ (.X(_02998_),
    .B(_10333_),
    .A(_10319_));
 sg13g2_nor2_2 _18908_ (.A(_10481_),
    .B(_02998_),
    .Y(_02999_));
 sg13g2_mux2_1 _18909_ (.A0(net3521),
    .A1(net5790),
    .S(_02999_),
    .X(_00275_));
 sg13g2_mux2_1 _18910_ (.A0(net3296),
    .A1(net5756),
    .S(_02999_),
    .X(_00276_));
 sg13g2_mux2_1 _18911_ (.A0(net3417),
    .A1(net5727),
    .S(_02999_),
    .X(_00277_));
 sg13g2_mux2_1 _18912_ (.A0(net3392),
    .A1(net5698),
    .S(_02999_),
    .X(_00278_));
 sg13g2_mux2_1 _18913_ (.A0(net3821),
    .A1(net5670),
    .S(_02999_),
    .X(_00279_));
 sg13g2_mux2_1 _18914_ (.A0(net3531),
    .A1(net5646),
    .S(_02999_),
    .X(_00280_));
 sg13g2_mux2_1 _18915_ (.A0(net3290),
    .A1(net5613),
    .S(_02999_),
    .X(_00281_));
 sg13g2_nand2_2 _18916_ (.Y(_03000_),
    .A(_10480_),
    .B(_10509_));
 sg13g2_mux2_1 _18917_ (.A0(net5790),
    .A1(net6713),
    .S(_03000_),
    .X(_00282_));
 sg13g2_mux2_1 _18918_ (.A0(net5756),
    .A1(net6157),
    .S(_03000_),
    .X(_00283_));
 sg13g2_mux2_1 _18919_ (.A0(net5727),
    .A1(net6727),
    .S(_03000_),
    .X(_00284_));
 sg13g2_mux2_1 _18920_ (.A0(net5698),
    .A1(net6866),
    .S(_03000_),
    .X(_00285_));
 sg13g2_mux2_1 _18921_ (.A0(net5673),
    .A1(net6390),
    .S(_03000_),
    .X(_00286_));
 sg13g2_mux2_1 _18922_ (.A0(net5646),
    .A1(net6101),
    .S(_03000_),
    .X(_00287_));
 sg13g2_mux2_1 _18923_ (.A0(net5613),
    .A1(net4372),
    .S(_03000_),
    .X(_00288_));
 sg13g2_nand2_1 _18924_ (.Y(_03001_),
    .A(net4878),
    .B(net5021));
 sg13g2_nand2_2 _18925_ (.Y(_03002_),
    .A(net5039),
    .B(net5028));
 sg13g2_nor2_2 _18926_ (.A(_03001_),
    .B(_03002_),
    .Y(_03003_));
 sg13g2_inv_1 _18927_ (.Y(_03004_),
    .A(_03003_));
 sg13g2_nand2_1 _18928_ (.Y(_03005_),
    .A(_08553_),
    .B(net5029));
 sg13g2_and2_1 _18929_ (.A(_10417_),
    .B(net4781),
    .X(_03006_));
 sg13g2_and3_2 _18930_ (.X(_03007_),
    .A(_08589_),
    .B(_10402_),
    .C(_03006_));
 sg13g2_nand3_1 _18931_ (.B(_10402_),
    .C(_03006_),
    .A(_08589_),
    .Y(_03008_));
 sg13g2_nor3_2 _18932_ (.A(net5032),
    .B(net4948),
    .C(_03008_),
    .Y(_03009_));
 sg13g2_nand2_2 _18933_ (.Y(_03010_),
    .A(_03003_),
    .B(_03009_));
 sg13g2_mux2_1 _18934_ (.A0(net5251),
    .A1(net4332),
    .S(_03010_),
    .X(_00289_));
 sg13g2_mux2_1 _18935_ (.A0(net5224),
    .A1(net6217),
    .S(_03010_),
    .X(_00290_));
 sg13g2_mux2_1 _18936_ (.A0(net5123),
    .A1(net6473),
    .S(_03010_),
    .X(_00291_));
 sg13g2_nor2_1 _18937_ (.A(_00101_),
    .B(_08640_),
    .Y(_03011_));
 sg13g2_a221oi_1 _18938_ (.B2(\atari2600.cpu.PC[3] ),
    .C1(_03011_),
    .B1(_08519_),
    .A1(\atari2600.cpu.PC[11] ),
    .Y(_03012_),
    .A2(_08497_));
 sg13g2_o21ai_1 _18939_ (.B1(_03012_),
    .Y(_03013_),
    .A1(_00147_),
    .A2(_08651_));
 sg13g2_nand2_1 _18940_ (.Y(_03014_),
    .A(_08517_),
    .B(_08586_));
 sg13g2_nor2b_2 _18941_ (.A(_03013_),
    .B_N(_03014_),
    .Y(_03015_));
 sg13g2_nand2b_2 _18942_ (.Y(_03016_),
    .B(_03014_),
    .A_N(_03013_));
 sg13g2_mux2_1 _18943_ (.A0(net5094),
    .A1(net6046),
    .S(_03010_),
    .X(_00292_));
 sg13g2_nand3_1 _18944_ (.B(_08618_),
    .C(_08619_),
    .A(_08586_),
    .Y(_03017_));
 sg13g2_o21ai_1 _18945_ (.B1(net5570),
    .Y(_03018_),
    .A1(net5479),
    .A2(net5436));
 sg13g2_a22oi_1 _18946_ (.Y(_03019_),
    .B1(net5397),
    .B2(\atari2600.cpu.PC[4] ),
    .A2(net5433),
    .A1(\atari2600.cpu.PC[12] ));
 sg13g2_nand4_1 _18947_ (.B(_08651_),
    .C(_03018_),
    .A(_08587_),
    .Y(_03020_),
    .D(_03019_));
 sg13g2_and2_1 _18948_ (.A(_03017_),
    .B(_03020_),
    .X(_03021_));
 sg13g2_nand2_2 _18949_ (.Y(_03022_),
    .A(_03017_),
    .B(_03020_));
 sg13g2_mux2_1 _18950_ (.A0(net5190),
    .A1(net4444),
    .S(_03010_),
    .X(_00293_));
 sg13g2_nand3_1 _18951_ (.B(_08607_),
    .C(_08608_),
    .A(_08586_),
    .Y(_03023_));
 sg13g2_a22oi_1 _18952_ (.Y(_03024_),
    .B1(net5436),
    .B2(\atari2600.cpu.ADD[5] ),
    .A2(net5479),
    .A1(_08076_));
 sg13g2_a22oi_1 _18953_ (.Y(_03025_),
    .B1(net5397),
    .B2(\atari2600.cpu.PC[5] ),
    .A2(net5433),
    .A1(\atari2600.cpu.PC[13] ));
 sg13g2_nand4_1 _18954_ (.B(_08651_),
    .C(_03024_),
    .A(_08587_),
    .Y(_03026_),
    .D(_03025_));
 sg13g2_and2_1 _18955_ (.A(_03023_),
    .B(_03026_),
    .X(_03027_));
 sg13g2_nand2_1 _18956_ (.Y(_03028_),
    .A(_03023_),
    .B(_03026_));
 sg13g2_mux2_1 _18957_ (.A0(net5163),
    .A1(net4383),
    .S(_03010_),
    .X(_00294_));
 sg13g2_nor2_1 _18958_ (.A(_00103_),
    .B(_08640_),
    .Y(_03029_));
 sg13g2_a221oi_1 _18959_ (.B2(\atari2600.cpu.PC[6] ),
    .C1(_03029_),
    .B1(net5397),
    .A1(\atari2600.cpu.PC[14] ),
    .Y(_03030_),
    .A2(net5433));
 sg13g2_o21ai_1 _18960_ (.B1(_03030_),
    .Y(_03031_),
    .A1(_00148_),
    .A2(_08651_));
 sg13g2_nand2_1 _18961_ (.Y(_03032_),
    .A(_08586_),
    .B(_08718_));
 sg13g2_nor2b_2 _18962_ (.A(_03031_),
    .B_N(_03032_),
    .Y(_03033_));
 sg13g2_nand2b_2 _18963_ (.Y(_03034_),
    .B(_03032_),
    .A_N(_03031_));
 sg13g2_mux2_1 _18964_ (.A0(net5071),
    .A1(net6678),
    .S(_03010_),
    .X(_00295_));
 sg13g2_nor2_1 _18965_ (.A(_00104_),
    .B(_08640_),
    .Y(_03035_));
 sg13g2_a221oi_1 _18966_ (.B2(\atari2600.cpu.PC[7] ),
    .C1(_03035_),
    .B1(net5397),
    .A1(\atari2600.cpu.PC[15] ),
    .Y(_03036_),
    .A2(net5433));
 sg13g2_o21ai_1 _18967_ (.B1(_03036_),
    .Y(_03037_),
    .A1(_00149_),
    .A2(_08651_));
 sg13g2_nand2_1 _18968_ (.Y(_03038_),
    .A(_08586_),
    .B(_08599_));
 sg13g2_nor2b_2 _18969_ (.A(_03037_),
    .B_N(_03038_),
    .Y(_03039_));
 sg13g2_nand2b_2 _18970_ (.Y(_03040_),
    .B(_03038_),
    .A_N(_03037_));
 sg13g2_mux2_1 _18971_ (.A0(net5045),
    .A1(net6129),
    .S(_03010_),
    .X(_00296_));
 sg13g2_nor3_2 _18972_ (.A(net5039),
    .B(net5021),
    .C(net4773),
    .Y(_03041_));
 sg13g2_inv_1 _18973_ (.Y(_03042_),
    .A(_03041_));
 sg13g2_nor2_2 _18974_ (.A(net5031),
    .B(_08732_),
    .Y(_03043_));
 sg13g2_and2_1 _18975_ (.A(_03007_),
    .B(_03043_),
    .X(_03044_));
 sg13g2_nand2_2 _18976_ (.Y(_03045_),
    .A(_03041_),
    .B(net4746));
 sg13g2_mux2_1 _18977_ (.A0(net5248),
    .A1(net4460),
    .S(_03045_),
    .X(_00297_));
 sg13g2_mux2_1 _18978_ (.A0(net5222),
    .A1(net6414),
    .S(_03045_),
    .X(_00298_));
 sg13g2_mux2_1 _18979_ (.A0(net5118),
    .A1(net4275),
    .S(_03045_),
    .X(_00299_));
 sg13g2_mux2_1 _18980_ (.A0(net5094),
    .A1(net6239),
    .S(_03045_),
    .X(_00300_));
 sg13g2_mux2_1 _18981_ (.A0(net5190),
    .A1(net4441),
    .S(_03045_),
    .X(_00301_));
 sg13g2_mux2_1 _18982_ (.A0(net5159),
    .A1(net6564),
    .S(_03045_),
    .X(_00302_));
 sg13g2_mux2_1 _18983_ (.A0(net5066),
    .A1(net6752),
    .S(_03045_),
    .X(_00303_));
 sg13g2_mux2_1 _18984_ (.A0(net5044),
    .A1(net6106),
    .S(_03045_),
    .X(_00304_));
 sg13g2_nor2_2 _18985_ (.A(net5472),
    .B(net5430),
    .Y(_03046_));
 sg13g2_mux2_1 _18986_ (.A0(net3449),
    .A1(net5779),
    .S(_03046_),
    .X(_00305_));
 sg13g2_mux2_1 _18987_ (.A0(net3991),
    .A1(net5749),
    .S(_03046_),
    .X(_00306_));
 sg13g2_mux2_1 _18988_ (.A0(net3586),
    .A1(net5719),
    .S(_03046_),
    .X(_00307_));
 sg13g2_mux2_1 _18989_ (.A0(net3390),
    .A1(net5686),
    .S(_03046_),
    .X(_00308_));
 sg13g2_mux2_1 _18990_ (.A0(net3204),
    .A1(net5656),
    .S(_03046_),
    .X(_00309_));
 sg13g2_mux2_1 _18991_ (.A0(net3614),
    .A1(net5635),
    .S(_03046_),
    .X(_00310_));
 sg13g2_mux2_1 _18992_ (.A0(net3609),
    .A1(net5599),
    .S(_03046_),
    .X(_00311_));
 sg13g2_nand2_2 _18993_ (.Y(_03047_),
    .A(net5036),
    .B(net5020));
 sg13g2_nor2_2 _18994_ (.A(net4775),
    .B(_03047_),
    .Y(_03048_));
 sg13g2_nand3_1 _18995_ (.B(net4803),
    .C(_03007_),
    .A(net5033),
    .Y(_03049_));
 sg13g2_nor3_2 _18996_ (.A(net4775),
    .B(_03047_),
    .C(net4744),
    .Y(_03050_));
 sg13g2_nor2_1 _18997_ (.A(net3851),
    .B(net4722),
    .Y(_03051_));
 sg13g2_a21oi_1 _18998_ (.A1(net5261),
    .A2(net4722),
    .Y(_00312_),
    .B1(_03051_));
 sg13g2_nor2_1 _18999_ (.A(net3611),
    .B(net4722),
    .Y(_03052_));
 sg13g2_a21oi_1 _19000_ (.A1(net5236),
    .A2(net4722),
    .Y(_00313_),
    .B1(_03052_));
 sg13g2_nor2_1 _19001_ (.A(net3637),
    .B(net4722),
    .Y(_03053_));
 sg13g2_a21oi_1 _19002_ (.A1(net5133),
    .A2(net4722),
    .Y(_00314_),
    .B1(_03053_));
 sg13g2_nor2_1 _19003_ (.A(net3020),
    .B(net4722),
    .Y(_03054_));
 sg13g2_a21oi_1 _19004_ (.A1(net5109),
    .A2(net4722),
    .Y(_00315_),
    .B1(_03054_));
 sg13g2_nor2_1 _19005_ (.A(net3087),
    .B(net4721),
    .Y(_03055_));
 sg13g2_a21oi_1 _19006_ (.A1(net5177),
    .A2(net4721),
    .Y(_00316_),
    .B1(_03055_));
 sg13g2_nor2_1 _19007_ (.A(net3477),
    .B(net4721),
    .Y(_03056_));
 sg13g2_a21oi_1 _19008_ (.A1(net5148),
    .A2(net4721),
    .Y(_00317_),
    .B1(_03056_));
 sg13g2_nor2_1 _19009_ (.A(net3900),
    .B(net4721),
    .Y(_03057_));
 sg13g2_a21oi_1 _19010_ (.A1(net5081),
    .A2(net4721),
    .Y(_00318_),
    .B1(_03057_));
 sg13g2_nor2_1 _19011_ (.A(net3161),
    .B(net4721),
    .Y(_03058_));
 sg13g2_a21oi_1 _19012_ (.A1(net5057),
    .A2(net4721),
    .Y(_00319_),
    .B1(_03058_));
 sg13g2_nor2_2 _19013_ (.A(_10253_),
    .B(_03001_),
    .Y(_03059_));
 sg13g2_inv_1 _19014_ (.Y(_03060_),
    .A(_03059_));
 sg13g2_nand3_1 _19015_ (.B(net4819),
    .C(_03007_),
    .A(net5031),
    .Y(_03061_));
 sg13g2_nor2_1 _19016_ (.A(_03060_),
    .B(net4742),
    .Y(_03062_));
 sg13g2_nor2_1 _19017_ (.A(net3089),
    .B(net4720),
    .Y(_03063_));
 sg13g2_a21oi_1 _19018_ (.A1(net5268),
    .A2(net4720),
    .Y(_00320_),
    .B1(_03063_));
 sg13g2_nor2_1 _19019_ (.A(net3309),
    .B(net4719),
    .Y(_03064_));
 sg13g2_a21oi_1 _19020_ (.A1(net5242),
    .A2(net4719),
    .Y(_00321_),
    .B1(_03064_));
 sg13g2_nor2_1 _19021_ (.A(net3471),
    .B(net4720),
    .Y(_03065_));
 sg13g2_a21oi_1 _19022_ (.A1(net5139),
    .A2(net4720),
    .Y(_00322_),
    .B1(_03065_));
 sg13g2_nor2_1 _19023_ (.A(net3986),
    .B(net4719),
    .Y(_03066_));
 sg13g2_a21oi_1 _19024_ (.A1(net5110),
    .A2(net4719),
    .Y(_00323_),
    .B1(_03066_));
 sg13g2_nor2_1 _19025_ (.A(net3099),
    .B(net4719),
    .Y(_03067_));
 sg13g2_a21oi_1 _19026_ (.A1(net5183),
    .A2(net4719),
    .Y(_00324_),
    .B1(_03067_));
 sg13g2_nor2_1 _19027_ (.A(net3074),
    .B(net4719),
    .Y(_03068_));
 sg13g2_a21oi_1 _19028_ (.A1(net5154),
    .A2(net4719),
    .Y(_00325_),
    .B1(_03068_));
 sg13g2_nor2_1 _19029_ (.A(net3642),
    .B(net4720),
    .Y(_03069_));
 sg13g2_a21oi_1 _19030_ (.A1(net5084),
    .A2(net4720),
    .Y(_00326_),
    .B1(_03069_));
 sg13g2_nor2_1 _19031_ (.A(net3120),
    .B(net4720),
    .Y(_03070_));
 sg13g2_a21oi_1 _19032_ (.A1(net5062),
    .A2(net4720),
    .Y(_00327_),
    .B1(_03070_));
 sg13g2_nor2_2 _19033_ (.A(_10373_),
    .B(net5430),
    .Y(_03071_));
 sg13g2_mux2_1 _19034_ (.A0(net4094),
    .A1(net5778),
    .S(_03071_),
    .X(_00328_));
 sg13g2_mux2_1 _19035_ (.A0(net3398),
    .A1(net5750),
    .S(_03071_),
    .X(_00329_));
 sg13g2_mux2_1 _19036_ (.A0(net3223),
    .A1(net5719),
    .S(_03071_),
    .X(_00330_));
 sg13g2_mux2_1 _19037_ (.A0(net3911),
    .A1(net5687),
    .S(_03071_),
    .X(_00331_));
 sg13g2_mux2_1 _19038_ (.A0(net3816),
    .A1(net5662),
    .S(_03071_),
    .X(_00332_));
 sg13g2_mux2_1 _19039_ (.A0(net3716),
    .A1(net5634),
    .S(_03071_),
    .X(_00333_));
 sg13g2_mux2_1 _19040_ (.A0(net3814),
    .A1(net5605),
    .S(_03071_),
    .X(_00334_));
 sg13g2_and2_1 _19041_ (.A(_10181_),
    .B(_10184_),
    .X(_03072_));
 sg13g2_nand2_2 _19042_ (.Y(_03073_),
    .A(_10478_),
    .B(net5417));
 sg13g2_mux2_1 _19043_ (.A0(net5771),
    .A1(net6808),
    .S(_03073_),
    .X(_00335_));
 sg13g2_mux2_1 _19044_ (.A0(net5742),
    .A1(net6591),
    .S(_03073_),
    .X(_00336_));
 sg13g2_mux2_1 _19045_ (.A0(net5713),
    .A1(net6949),
    .S(_03073_),
    .X(_00337_));
 sg13g2_mux2_1 _19046_ (.A0(net5685),
    .A1(net6500),
    .S(_03073_),
    .X(_00338_));
 sg13g2_mux2_1 _19047_ (.A0(net5656),
    .A1(net6079),
    .S(_03073_),
    .X(_00339_));
 sg13g2_mux2_1 _19048_ (.A0(net5626),
    .A1(net6753),
    .S(_03073_),
    .X(_00340_));
 sg13g2_mux2_1 _19049_ (.A0(net5598),
    .A1(net6425),
    .S(_03073_),
    .X(_00341_));
 sg13g2_nor2_2 _19050_ (.A(_10259_),
    .B(_10319_),
    .Y(_03074_));
 sg13g2_nand2_2 _19051_ (.Y(_03075_),
    .A(_03072_),
    .B(net5416));
 sg13g2_mux2_1 _19052_ (.A0(net5775),
    .A1(net6803),
    .S(_03075_),
    .X(_00342_));
 sg13g2_mux2_1 _19053_ (.A0(net5746),
    .A1(net4373),
    .S(_03075_),
    .X(_00343_));
 sg13g2_mux2_1 _19054_ (.A0(net5716),
    .A1(net6963),
    .S(_03075_),
    .X(_00344_));
 sg13g2_mux2_1 _19055_ (.A0(net5688),
    .A1(net4311),
    .S(_03075_),
    .X(_00345_));
 sg13g2_mux2_1 _19056_ (.A0(net5661),
    .A1(net6524),
    .S(_03075_),
    .X(_00346_));
 sg13g2_mux2_1 _19057_ (.A0(net5631),
    .A1(net6202),
    .S(_03075_),
    .X(_00347_));
 sg13g2_mux2_1 _19058_ (.A0(net5606),
    .A1(net6313),
    .S(_03075_),
    .X(_00348_));
 sg13g2_nor2_2 _19059_ (.A(_10261_),
    .B(_10371_),
    .Y(_03076_));
 sg13g2_nand2_2 _19060_ (.Y(_03077_),
    .A(_10260_),
    .B(_10370_));
 sg13g2_nor2_2 _19061_ (.A(_10198_),
    .B(_10375_),
    .Y(_03078_));
 sg13g2_nand2_2 _19062_ (.Y(_03079_),
    .A(_10199_),
    .B(_10374_));
 sg13g2_nor2_2 _19063_ (.A(_03077_),
    .B(_03079_),
    .Y(_03080_));
 sg13g2_mux2_1 _19064_ (.A0(net3334),
    .A1(net5797),
    .S(_03080_),
    .X(_00349_));
 sg13g2_mux2_1 _19065_ (.A0(net3315),
    .A1(net5767),
    .S(_03080_),
    .X(_00350_));
 sg13g2_mux2_1 _19066_ (.A0(net3402),
    .A1(net5737),
    .S(_03080_),
    .X(_00351_));
 sg13g2_mux2_1 _19067_ (.A0(net3177),
    .A1(net5707),
    .S(_03080_),
    .X(_00352_));
 sg13g2_mux2_1 _19068_ (.A0(net3601),
    .A1(net5680),
    .S(_03080_),
    .X(_00353_));
 sg13g2_mux2_1 _19069_ (.A0(net3229),
    .A1(net5652),
    .S(_03080_),
    .X(_00354_));
 sg13g2_mux2_1 _19070_ (.A0(net3131),
    .A1(net5621),
    .S(_03080_),
    .X(_00355_));
 sg13g2_nor3_2 _19071_ (.A(net5816),
    .B(net5559),
    .C(_10375_),
    .Y(_03081_));
 sg13g2_nand2_2 _19072_ (.Y(_03082_),
    .A(_10201_),
    .B(_10374_));
 sg13g2_nor2_2 _19073_ (.A(_02998_),
    .B(net5414),
    .Y(_03083_));
 sg13g2_mux2_1 _19074_ (.A0(net3157),
    .A1(net5793),
    .S(_03083_),
    .X(_00356_));
 sg13g2_mux2_1 _19075_ (.A0(net3400),
    .A1(net5758),
    .S(_03083_),
    .X(_00357_));
 sg13g2_mux2_1 _19076_ (.A0(net3235),
    .A1(net5728),
    .S(_03083_),
    .X(_00358_));
 sg13g2_mux2_1 _19077_ (.A0(net3746),
    .A1(net5701),
    .S(_03083_),
    .X(_00359_));
 sg13g2_mux2_1 _19078_ (.A0(net3335),
    .A1(net5670),
    .S(_03083_),
    .X(_00360_));
 sg13g2_mux2_1 _19079_ (.A0(net3575),
    .A1(net5647),
    .S(_03083_),
    .X(_00361_));
 sg13g2_mux2_1 _19080_ (.A0(net3607),
    .A1(net5612),
    .S(_03083_),
    .X(_00362_));
 sg13g2_nor2_2 _19081_ (.A(_10504_),
    .B(net5415),
    .Y(_03084_));
 sg13g2_mux2_1 _19082_ (.A0(net3299),
    .A1(net5795),
    .S(_03084_),
    .X(_00363_));
 sg13g2_mux2_1 _19083_ (.A0(net3973),
    .A1(net5766),
    .S(_03084_),
    .X(_00364_));
 sg13g2_mux2_1 _19084_ (.A0(net3483),
    .A1(net5737),
    .S(_03084_),
    .X(_00365_));
 sg13g2_mux2_1 _19085_ (.A0(net3255),
    .A1(net5708),
    .S(_03084_),
    .X(_00366_));
 sg13g2_mux2_1 _19086_ (.A0(net3689),
    .A1(net5680),
    .S(_03084_),
    .X(_00367_));
 sg13g2_mux2_1 _19087_ (.A0(net3381),
    .A1(net5651),
    .S(_03084_),
    .X(_00368_));
 sg13g2_mux2_1 _19088_ (.A0(net3163),
    .A1(net5622),
    .S(_03084_),
    .X(_00369_));
 sg13g2_nor2_2 _19089_ (.A(net5467),
    .B(net5415),
    .Y(_03085_));
 sg13g2_mux2_1 _19090_ (.A0(net3699),
    .A1(net5795),
    .S(_03085_),
    .X(_00370_));
 sg13g2_mux2_1 _19091_ (.A0(net4104),
    .A1(net5766),
    .S(_03085_),
    .X(_00371_));
 sg13g2_mux2_1 _19092_ (.A0(net3725),
    .A1(net5737),
    .S(_03085_),
    .X(_00372_));
 sg13g2_mux2_1 _19093_ (.A0(net3246),
    .A1(net5708),
    .S(_03085_),
    .X(_00373_));
 sg13g2_mux2_1 _19094_ (.A0(net3216),
    .A1(net5680),
    .S(_03085_),
    .X(_00374_));
 sg13g2_mux2_1 _19095_ (.A0(net3387),
    .A1(net5650),
    .S(_03085_),
    .X(_00375_));
 sg13g2_mux2_1 _19096_ (.A0(net3736),
    .A1(net5622),
    .S(_03085_),
    .X(_00376_));
 sg13g2_and2_2 _19097_ (.A(_10509_),
    .B(_03078_),
    .X(_03086_));
 sg13g2_mux2_1 _19098_ (.A0(net3728),
    .A1(net5795),
    .S(_03086_),
    .X(_00377_));
 sg13g2_mux2_1 _19099_ (.A0(net2969),
    .A1(net5766),
    .S(_03086_),
    .X(_00378_));
 sg13g2_mux2_1 _19100_ (.A0(net3458),
    .A1(net5735),
    .S(_03086_),
    .X(_00379_));
 sg13g2_mux2_1 _19101_ (.A0(net3665),
    .A1(net5709),
    .S(_03086_),
    .X(_00380_));
 sg13g2_mux2_1 _19102_ (.A0(net3629),
    .A1(net5680),
    .S(_03086_),
    .X(_00381_));
 sg13g2_mux2_1 _19103_ (.A0(net3434),
    .A1(net5651),
    .S(_03086_),
    .X(_00382_));
 sg13g2_mux2_1 _19104_ (.A0(net3116),
    .A1(net5622),
    .S(_03086_),
    .X(_00383_));
 sg13g2_nor2_2 _19105_ (.A(net4778),
    .B(_03047_),
    .Y(_03087_));
 sg13g2_or2_1 _19106_ (.X(_03088_),
    .B(_03047_),
    .A(net4778));
 sg13g2_nand2_2 _19107_ (.Y(_03089_),
    .A(_03007_),
    .B(_03087_));
 sg13g2_nor2_2 _19108_ (.A(_10252_),
    .B(_03008_),
    .Y(_03090_));
 sg13g2_and2_1 _19109_ (.A(_03087_),
    .B(net4740),
    .X(_03091_));
 sg13g2_nor2_1 _19110_ (.A(net3722),
    .B(net4718),
    .Y(_03092_));
 sg13g2_a21oi_1 _19111_ (.A1(net5266),
    .A2(net4718),
    .Y(_00384_),
    .B1(_03092_));
 sg13g2_nor2_1 _19112_ (.A(net3005),
    .B(net4718),
    .Y(_03093_));
 sg13g2_a21oi_1 _19113_ (.A1(net5242),
    .A2(net4718),
    .Y(_00385_),
    .B1(_03093_));
 sg13g2_nor2_1 _19114_ (.A(net2986),
    .B(net4718),
    .Y(_03094_));
 sg13g2_a21oi_1 _19115_ (.A1(net5138),
    .A2(net4718),
    .Y(_00386_),
    .B1(_03094_));
 sg13g2_nor2_1 _19116_ (.A(net3097),
    .B(net4717),
    .Y(_03095_));
 sg13g2_a21oi_1 _19117_ (.A1(net5108),
    .A2(net4717),
    .Y(_00387_),
    .B1(_03095_));
 sg13g2_nor2_1 _19118_ (.A(net3105),
    .B(net4717),
    .Y(_03096_));
 sg13g2_a21oi_1 _19119_ (.A1(net5181),
    .A2(net4717),
    .Y(_00388_),
    .B1(_03096_));
 sg13g2_nor2_1 _19120_ (.A(net3553),
    .B(net4717),
    .Y(_03097_));
 sg13g2_a21oi_1 _19121_ (.A1(net5153),
    .A2(net4717),
    .Y(_00389_),
    .B1(_03097_));
 sg13g2_nor2_1 _19122_ (.A(net3694),
    .B(net4718),
    .Y(_03098_));
 sg13g2_a21oi_1 _19123_ (.A1(net5084),
    .A2(net4718),
    .Y(_00390_),
    .B1(_03098_));
 sg13g2_nor2_1 _19124_ (.A(net3010),
    .B(net4717),
    .Y(_03099_));
 sg13g2_a21oi_1 _19125_ (.A1(net5060),
    .A2(net4717),
    .Y(_00391_),
    .B1(_03099_));
 sg13g2_nor2_2 _19126_ (.A(_10259_),
    .B(_10261_),
    .Y(_03100_));
 sg13g2_nand3_1 _19127_ (.B(net5562),
    .C(_10260_),
    .A(net5564),
    .Y(_03101_));
 sg13g2_nor2_2 _19128_ (.A(net5414),
    .B(_03101_),
    .Y(_03102_));
 sg13g2_mux2_1 _19129_ (.A0(net3512),
    .A1(net5791),
    .S(_03102_),
    .X(_00392_));
 sg13g2_mux2_1 _19130_ (.A0(net3624),
    .A1(net5759),
    .S(_03102_),
    .X(_00393_));
 sg13g2_mux2_1 _19131_ (.A0(net3540),
    .A1(net5735),
    .S(_03102_),
    .X(_00394_));
 sg13g2_mux2_1 _19132_ (.A0(net3950),
    .A1(net5706),
    .S(_03102_),
    .X(_00395_));
 sg13g2_mux2_1 _19133_ (.A0(net3748),
    .A1(net5670),
    .S(_03102_),
    .X(_00396_));
 sg13g2_mux2_1 _19134_ (.A0(net3548),
    .A1(net5646),
    .S(_03102_),
    .X(_00397_));
 sg13g2_mux2_1 _19135_ (.A0(net3767),
    .A1(net5622),
    .S(_03102_),
    .X(_00398_));
 sg13g2_nand2_2 _19136_ (.Y(_03103_),
    .A(_10372_),
    .B(net5470));
 sg13g2_mux2_1 _19137_ (.A0(net5785),
    .A1(net6280),
    .S(_03103_),
    .X(_00399_));
 sg13g2_mux2_1 _19138_ (.A0(net5753),
    .A1(net6617),
    .S(_03103_),
    .X(_00400_));
 sg13g2_mux2_1 _19139_ (.A0(net5724),
    .A1(net6698),
    .S(_03103_),
    .X(_00401_));
 sg13g2_mux2_1 _19140_ (.A0(net5695),
    .A1(net6111),
    .S(_03103_),
    .X(_00402_));
 sg13g2_mux2_1 _19141_ (.A0(net5668),
    .A1(net6304),
    .S(_03103_),
    .X(_00403_));
 sg13g2_mux2_1 _19142_ (.A0(net5639),
    .A1(net6052),
    .S(_03103_),
    .X(_00404_));
 sg13g2_mux2_1 _19143_ (.A0(net5609),
    .A1(net6896),
    .S(_03103_),
    .X(_00405_));
 sg13g2_nor3_2 _19144_ (.A(_08111_),
    .B(net5811),
    .C(_10375_),
    .Y(_03104_));
 sg13g2_nand2_2 _19145_ (.Y(_03105_),
    .A(_10200_),
    .B(_10374_));
 sg13g2_nor2_2 _19146_ (.A(_02996_),
    .B(_03105_),
    .Y(_03106_));
 sg13g2_mux2_1 _19147_ (.A0(net3673),
    .A1(net5787),
    .S(_03106_),
    .X(_00406_));
 sg13g2_mux2_1 _19148_ (.A0(net3388),
    .A1(net5762),
    .S(_03106_),
    .X(_00407_));
 sg13g2_mux2_1 _19149_ (.A0(net3276),
    .A1(net5731),
    .S(_03106_),
    .X(_00408_));
 sg13g2_mux2_1 _19150_ (.A0(net3183),
    .A1(net5705),
    .S(_03106_),
    .X(_00409_));
 sg13g2_mux2_1 _19151_ (.A0(net3170),
    .A1(net5676),
    .S(_03106_),
    .X(_00410_));
 sg13g2_mux2_1 _19152_ (.A0(net3813),
    .A1(net5645),
    .S(_03106_),
    .X(_00411_));
 sg13g2_mux2_1 _19153_ (.A0(net3418),
    .A1(net5617),
    .S(_03106_),
    .X(_00412_));
 sg13g2_nor2_2 _19154_ (.A(_10382_),
    .B(net5425),
    .Y(_03107_));
 sg13g2_mux2_1 _19155_ (.A0(net3310),
    .A1(net5790),
    .S(_03107_),
    .X(_00413_));
 sg13g2_mux2_1 _19156_ (.A0(net3499),
    .A1(net5756),
    .S(_03107_),
    .X(_00414_));
 sg13g2_mux2_1 _19157_ (.A0(net3493),
    .A1(net5723),
    .S(_03107_),
    .X(_00415_));
 sg13g2_mux2_1 _19158_ (.A0(net3681),
    .A1(net5694),
    .S(_03107_),
    .X(_00416_));
 sg13g2_mux2_1 _19159_ (.A0(net3516),
    .A1(net5665),
    .S(_03107_),
    .X(_00417_));
 sg13g2_mux2_1 _19160_ (.A0(net4015),
    .A1(net5640),
    .S(_03107_),
    .X(_00418_));
 sg13g2_mux2_1 _19161_ (.A0(net3740),
    .A1(net5608),
    .S(_03107_),
    .X(_00419_));
 sg13g2_nor2_2 _19162_ (.A(net5472),
    .B(_10377_),
    .Y(_03108_));
 sg13g2_mux2_1 _19163_ (.A0(net3526),
    .A1(net5771),
    .S(_03108_),
    .X(_00420_));
 sg13g2_mux2_1 _19164_ (.A0(net3441),
    .A1(net5742),
    .S(_03108_),
    .X(_00421_));
 sg13g2_mux2_1 _19165_ (.A0(net3709),
    .A1(net5713),
    .S(_03108_),
    .X(_00422_));
 sg13g2_mux2_1 _19166_ (.A0(net3468),
    .A1(net5684),
    .S(_03108_),
    .X(_00423_));
 sg13g2_mux2_1 _19167_ (.A0(net3545),
    .A1(net5655),
    .S(_03108_),
    .X(_00424_));
 sg13g2_mux2_1 _19168_ (.A0(net3544),
    .A1(net5626),
    .S(_03108_),
    .X(_00425_));
 sg13g2_mux2_1 _19169_ (.A0(net3809),
    .A1(net5597),
    .S(_03108_),
    .X(_00426_));
 sg13g2_nor2_2 _19170_ (.A(_10479_),
    .B(net5415),
    .Y(_03109_));
 sg13g2_mux2_1 _19171_ (.A0(net3270),
    .A1(net5798),
    .S(_03109_),
    .X(_00427_));
 sg13g2_mux2_1 _19172_ (.A0(net3470),
    .A1(net5767),
    .S(_03109_),
    .X(_00428_));
 sg13g2_mux2_1 _19173_ (.A0(net3902),
    .A1(net5739),
    .S(_03109_),
    .X(_00429_));
 sg13g2_mux2_1 _19174_ (.A0(net3429),
    .A1(net5709),
    .S(_03109_),
    .X(_00430_));
 sg13g2_mux2_1 _19175_ (.A0(net3583),
    .A1(net5681),
    .S(_03109_),
    .X(_00431_));
 sg13g2_mux2_1 _19176_ (.A0(net3922),
    .A1(net5652),
    .S(_03109_),
    .X(_00432_));
 sg13g2_mux2_1 _19177_ (.A0(net3180),
    .A1(net5623),
    .S(_03109_),
    .X(_00433_));
 sg13g2_nor2_2 _19178_ (.A(net5430),
    .B(_02996_),
    .Y(_03110_));
 sg13g2_mux2_1 _19179_ (.A0(net3494),
    .A1(net5776),
    .S(_03110_),
    .X(_00434_));
 sg13g2_mux2_1 _19180_ (.A0(net3631),
    .A1(net5749),
    .S(_03110_),
    .X(_00435_));
 sg13g2_mux2_1 _19181_ (.A0(net3495),
    .A1(net5720),
    .S(_03110_),
    .X(_00436_));
 sg13g2_mux2_1 _19182_ (.A0(net3737),
    .A1(net5692),
    .S(_03110_),
    .X(_00437_));
 sg13g2_mux2_1 _19183_ (.A0(net3476),
    .A1(net5662),
    .S(_03110_),
    .X(_00438_));
 sg13g2_mux2_1 _19184_ (.A0(net3938),
    .A1(net5636),
    .S(_03110_),
    .X(_00439_));
 sg13g2_mux2_1 _19185_ (.A0(net3403),
    .A1(net5604),
    .S(_03110_),
    .X(_00440_));
 sg13g2_nor2_2 _19186_ (.A(_10382_),
    .B(net5415),
    .Y(_03111_));
 sg13g2_mux2_1 _19187_ (.A0(net3550),
    .A1(net5798),
    .S(_03111_),
    .X(_00441_));
 sg13g2_mux2_1 _19188_ (.A0(net3885),
    .A1(net5767),
    .S(_03111_),
    .X(_00442_));
 sg13g2_mux2_1 _19189_ (.A0(net3357),
    .A1(net5739),
    .S(_03111_),
    .X(_00443_));
 sg13g2_mux2_1 _19190_ (.A0(net3446),
    .A1(net5709),
    .S(_03111_),
    .X(_00444_));
 sg13g2_mux2_1 _19191_ (.A0(net3832),
    .A1(net5681),
    .S(_03111_),
    .X(_00445_));
 sg13g2_mux2_1 _19192_ (.A0(net3940),
    .A1(net5653),
    .S(_03111_),
    .X(_00446_));
 sg13g2_mux2_1 _19193_ (.A0(net3345),
    .A1(net5623),
    .S(_03111_),
    .X(_00447_));
 sg13g2_nor2_2 _19194_ (.A(_02996_),
    .B(net5415),
    .Y(_03112_));
 sg13g2_mux2_1 _19195_ (.A0(net3127),
    .A1(net5798),
    .S(_03112_),
    .X(_00448_));
 sg13g2_mux2_1 _19196_ (.A0(net3206),
    .A1(net5766),
    .S(_03112_),
    .X(_00449_));
 sg13g2_mux2_1 _19197_ (.A0(net3672),
    .A1(net5738),
    .S(_03112_),
    .X(_00450_));
 sg13g2_mux2_1 _19198_ (.A0(net3273),
    .A1(net5709),
    .S(_03112_),
    .X(_00451_));
 sg13g2_mux2_1 _19199_ (.A0(net3768),
    .A1(net5681),
    .S(_03112_),
    .X(_00452_));
 sg13g2_mux2_1 _19200_ (.A0(net3944),
    .A1(net5653),
    .S(_03112_),
    .X(_00453_));
 sg13g2_mux2_1 _19201_ (.A0(net3563),
    .A1(net5621),
    .S(_03112_),
    .X(_00454_));
 sg13g2_nor3_2 _19202_ (.A(net5827),
    .B(net5830),
    .C(_10380_),
    .Y(_03113_));
 sg13g2_nand2_2 _19203_ (.Y(_03114_),
    .A(_03078_),
    .B(net5412));
 sg13g2_mux2_1 _19204_ (.A0(net5798),
    .A1(net4134),
    .S(_03114_),
    .X(_00455_));
 sg13g2_mux2_1 _19205_ (.A0(net5766),
    .A1(net6195),
    .S(_03114_),
    .X(_00456_));
 sg13g2_mux2_1 _19206_ (.A0(net5739),
    .A1(net6201),
    .S(_03114_),
    .X(_00457_));
 sg13g2_mux2_1 _19207_ (.A0(net5708),
    .A1(net4359),
    .S(_03114_),
    .X(_00458_));
 sg13g2_mux2_1 _19208_ (.A0(net5681),
    .A1(net4199),
    .S(_03114_),
    .X(_00459_));
 sg13g2_mux2_1 _19209_ (.A0(net5652),
    .A1(net6432),
    .S(_03114_),
    .X(_00460_));
 sg13g2_mux2_1 _19210_ (.A0(net5621),
    .A1(net6071),
    .S(_03114_),
    .X(_00461_));
 sg13g2_nand2_2 _19211_ (.Y(_03115_),
    .A(_10383_),
    .B(net5412));
 sg13g2_mux2_1 _19212_ (.A0(net5776),
    .A1(net6652),
    .S(_03115_),
    .X(_00462_));
 sg13g2_mux2_1 _19213_ (.A0(net5749),
    .A1(net6312),
    .S(_03115_),
    .X(_00463_));
 sg13g2_mux2_1 _19214_ (.A0(net5719),
    .A1(net4519),
    .S(_03115_),
    .X(_00464_));
 sg13g2_mux2_1 _19215_ (.A0(net5691),
    .A1(net6548),
    .S(_03115_),
    .X(_00465_));
 sg13g2_mux2_1 _19216_ (.A0(net5662),
    .A1(net6136),
    .S(_03115_),
    .X(_00466_));
 sg13g2_mux2_1 _19217_ (.A0(net5636),
    .A1(net6585),
    .S(_03115_),
    .X(_00467_));
 sg13g2_mux2_1 _19218_ (.A0(net5604),
    .A1(net6165),
    .S(_03115_),
    .X(_00468_));
 sg13g2_nand2_2 _19219_ (.Y(_03116_),
    .A(_10478_),
    .B(net5469));
 sg13g2_mux2_1 _19220_ (.A0(net5782),
    .A1(net6621),
    .S(_03116_),
    .X(_00469_));
 sg13g2_mux2_1 _19221_ (.A0(net5753),
    .A1(net6811),
    .S(_03116_),
    .X(_00470_));
 sg13g2_mux2_1 _19222_ (.A0(net5724),
    .A1(net6786),
    .S(_03116_),
    .X(_00471_));
 sg13g2_mux2_1 _19223_ (.A0(net5695),
    .A1(net4467),
    .S(_03116_),
    .X(_00472_));
 sg13g2_mux2_1 _19224_ (.A0(net5667),
    .A1(net6936),
    .S(_03116_),
    .X(_00473_));
 sg13g2_mux2_1 _19225_ (.A0(net5639),
    .A1(net6799),
    .S(_03116_),
    .X(_00474_));
 sg13g2_mux2_1 _19226_ (.A0(net5609),
    .A1(net6777),
    .S(_03116_),
    .X(_00475_));
 sg13g2_nor2_2 _19227_ (.A(net5430),
    .B(_03077_),
    .Y(_03117_));
 sg13g2_mux2_1 _19228_ (.A0(net3705),
    .A1(net5778),
    .S(_03117_),
    .X(_00476_));
 sg13g2_mux2_1 _19229_ (.A0(net3617),
    .A1(net5750),
    .S(_03117_),
    .X(_00477_));
 sg13g2_mux2_1 _19230_ (.A0(net3656),
    .A1(net5719),
    .S(_03117_),
    .X(_00478_));
 sg13g2_mux2_1 _19231_ (.A0(net3549),
    .A1(net5692),
    .S(_03117_),
    .X(_00479_));
 sg13g2_mux2_1 _19232_ (.A0(net3205),
    .A1(net5662),
    .S(_03117_),
    .X(_00480_));
 sg13g2_mux2_1 _19233_ (.A0(net3558),
    .A1(net5636),
    .S(_03117_),
    .X(_00481_));
 sg13g2_mux2_1 _19234_ (.A0(net3350),
    .A1(net5604),
    .S(_03117_),
    .X(_00482_));
 sg13g2_nor2_2 _19235_ (.A(_10317_),
    .B(_10371_),
    .Y(_03118_));
 sg13g2_nand2_2 _19236_ (.Y(_03119_),
    .A(_10316_),
    .B(_10370_));
 sg13g2_nor2_2 _19237_ (.A(_03079_),
    .B(_03119_),
    .Y(_03120_));
 sg13g2_mux2_1 _19238_ (.A0(net3212),
    .A1(net5797),
    .S(_03120_),
    .X(_00483_));
 sg13g2_mux2_1 _19239_ (.A0(net3254),
    .A1(net5767),
    .S(_03120_),
    .X(_00484_));
 sg13g2_mux2_1 _19240_ (.A0(net3790),
    .A1(net5736),
    .S(_03120_),
    .X(_00485_));
 sg13g2_mux2_1 _19241_ (.A0(net3405),
    .A1(net5706),
    .S(_03120_),
    .X(_00486_));
 sg13g2_mux2_1 _19242_ (.A0(net3490),
    .A1(net5680),
    .S(_03120_),
    .X(_00487_));
 sg13g2_mux2_1 _19243_ (.A0(net3436),
    .A1(net5652),
    .S(_03120_),
    .X(_00488_));
 sg13g2_mux2_1 _19244_ (.A0(net3215),
    .A1(net5621),
    .S(_03120_),
    .X(_00489_));
 sg13g2_nor2_2 _19245_ (.A(net5430),
    .B(_03119_),
    .Y(_03121_));
 sg13g2_mux2_1 _19246_ (.A0(net3758),
    .A1(net5778),
    .S(_03121_),
    .X(_00490_));
 sg13g2_mux2_1 _19247_ (.A0(net3925),
    .A1(net5750),
    .S(_03121_),
    .X(_00491_));
 sg13g2_mux2_1 _19248_ (.A0(net3834),
    .A1(net5719),
    .S(_03121_),
    .X(_00492_));
 sg13g2_mux2_1 _19249_ (.A0(net3541),
    .A1(net5691),
    .S(_03121_),
    .X(_00493_));
 sg13g2_mux2_1 _19250_ (.A0(net3661),
    .A1(net5662),
    .S(_03121_),
    .X(_00494_));
 sg13g2_mux2_1 _19251_ (.A0(net3841),
    .A1(net5634),
    .S(_03121_),
    .X(_00495_));
 sg13g2_mux2_1 _19252_ (.A0(net3608),
    .A1(net5605),
    .S(_03121_),
    .X(_00496_));
 sg13g2_nor2_2 _19253_ (.A(_10373_),
    .B(net5415),
    .Y(_03122_));
 sg13g2_mux2_1 _19254_ (.A0(net3603),
    .A1(net5797),
    .S(_03122_),
    .X(_00497_));
 sg13g2_mux2_1 _19255_ (.A0(net3683),
    .A1(net5767),
    .S(_03122_),
    .X(_00498_));
 sg13g2_mux2_1 _19256_ (.A0(net3997),
    .A1(net5736),
    .S(_03122_),
    .X(_00499_));
 sg13g2_mux2_1 _19257_ (.A0(net3543),
    .A1(net5707),
    .S(_03122_),
    .X(_00500_));
 sg13g2_mux2_1 _19258_ (.A0(net3141),
    .A1(net5680),
    .S(_03122_),
    .X(_00501_));
 sg13g2_mux2_1 _19259_ (.A0(net3327),
    .A1(net5652),
    .S(_03122_),
    .X(_00502_));
 sg13g2_mux2_1 _19260_ (.A0(net3510),
    .A1(net5621),
    .S(_03122_),
    .X(_00503_));
 sg13g2_nor2b_2 _19261_ (.A(net5471),
    .B_N(net5470),
    .Y(_03123_));
 sg13g2_mux2_1 _19262_ (.A0(net3917),
    .A1(net5783),
    .S(_03123_),
    .X(_00504_));
 sg13g2_mux2_1 _19263_ (.A0(net3667),
    .A1(net5754),
    .S(_03123_),
    .X(_00505_));
 sg13g2_mux2_1 _19264_ (.A0(net3261),
    .A1(net5725),
    .S(_03123_),
    .X(_00506_));
 sg13g2_mux2_1 _19265_ (.A0(net3384),
    .A1(net5696),
    .S(_03123_),
    .X(_00507_));
 sg13g2_mux2_1 _19266_ (.A0(net3745),
    .A1(net5668),
    .S(_03123_),
    .X(_00508_));
 sg13g2_mux2_1 _19267_ (.A0(net3437),
    .A1(net5641),
    .S(_03123_),
    .X(_00509_));
 sg13g2_mux2_1 _19268_ (.A0(net3696),
    .A1(net5610),
    .S(_03123_),
    .X(_00510_));
 sg13g2_nor3_2 _19269_ (.A(net5827),
    .B(net5830),
    .C(_10371_),
    .Y(_03124_));
 sg13g2_nand2_2 _19270_ (.Y(_03125_),
    .A(_03078_),
    .B(net5411));
 sg13g2_mux2_1 _19271_ (.A0(net5797),
    .A1(net4435),
    .S(_03125_),
    .X(_00511_));
 sg13g2_mux2_1 _19272_ (.A0(net5767),
    .A1(net6361),
    .S(_03125_),
    .X(_00512_));
 sg13g2_mux2_1 _19273_ (.A0(net5736),
    .A1(net4323),
    .S(_03125_),
    .X(_00513_));
 sg13g2_mux2_1 _19274_ (.A0(net5707),
    .A1(net6168),
    .S(_03125_),
    .X(_00514_));
 sg13g2_mux2_1 _19275_ (.A0(net5680),
    .A1(net4189),
    .S(_03125_),
    .X(_00515_));
 sg13g2_mux2_1 _19276_ (.A0(net5652),
    .A1(net6528),
    .S(_03125_),
    .X(_00516_));
 sg13g2_mux2_1 _19277_ (.A0(net5621),
    .A1(net6612),
    .S(_03125_),
    .X(_00517_));
 sg13g2_nand2_2 _19278_ (.Y(_03126_),
    .A(_10383_),
    .B(net5411));
 sg13g2_mux2_1 _19279_ (.A0(net5778),
    .A1(net6293),
    .S(_03126_),
    .X(_00518_));
 sg13g2_mux2_1 _19280_ (.A0(net5744),
    .A1(net6751),
    .S(_03126_),
    .X(_00519_));
 sg13g2_mux2_1 _19281_ (.A0(net5719),
    .A1(net4433),
    .S(_03126_),
    .X(_00520_));
 sg13g2_mux2_1 _19282_ (.A0(net5687),
    .A1(net6956),
    .S(_03126_),
    .X(_00521_));
 sg13g2_mux2_1 _19283_ (.A0(net5662),
    .A1(net6267),
    .S(_03126_),
    .X(_00522_));
 sg13g2_mux2_1 _19284_ (.A0(net5634),
    .A1(net6944),
    .S(_03126_),
    .X(_00523_));
 sg13g2_mux2_1 _19285_ (.A0(net5605),
    .A1(net4430),
    .S(_03126_),
    .X(_00524_));
 sg13g2_nor2_2 _19286_ (.A(net5415),
    .B(_03101_),
    .Y(_03127_));
 sg13g2_mux2_1 _19287_ (.A0(net3484),
    .A1(net5794),
    .S(_03127_),
    .X(_00525_));
 sg13g2_mux2_1 _19288_ (.A0(net3682),
    .A1(net5768),
    .S(_03127_),
    .X(_00526_));
 sg13g2_mux2_1 _19289_ (.A0(net3594),
    .A1(net5738),
    .S(_03127_),
    .X(_00527_));
 sg13g2_mux2_1 _19290_ (.A0(net3507),
    .A1(net5708),
    .S(_03127_),
    .X(_00528_));
 sg13g2_mux2_1 _19291_ (.A0(net3427),
    .A1(net5681),
    .S(_03127_),
    .X(_00529_));
 sg13g2_mux2_1 _19292_ (.A0(net3478),
    .A1(net5652),
    .S(_03127_),
    .X(_00530_));
 sg13g2_mux2_1 _19293_ (.A0(net3391),
    .A1(net5624),
    .S(_03127_),
    .X(_00531_));
 sg13g2_nor2_2 _19294_ (.A(net5430),
    .B(_03101_),
    .Y(_03128_));
 sg13g2_mux2_1 _19295_ (.A0(net3248),
    .A1(net5776),
    .S(_03128_),
    .X(_00532_));
 sg13g2_mux2_1 _19296_ (.A0(net3827),
    .A1(net5750),
    .S(_03128_),
    .X(_00533_));
 sg13g2_mux2_1 _19297_ (.A0(net4061),
    .A1(net5718),
    .S(_03128_),
    .X(_00534_));
 sg13g2_mux2_1 _19298_ (.A0(net3924),
    .A1(net5691),
    .S(_03128_),
    .X(_00535_));
 sg13g2_mux2_1 _19299_ (.A0(net3368),
    .A1(net5661),
    .S(_03128_),
    .X(_00536_));
 sg13g2_mux2_1 _19300_ (.A0(net3595),
    .A1(net5631),
    .S(_03128_),
    .X(_00537_));
 sg13g2_mux2_1 _19301_ (.A0(net3538),
    .A1(net5605),
    .S(_03128_),
    .X(_00538_));
 sg13g2_and2_2 _19302_ (.A(_10507_),
    .B(_03078_),
    .X(_03129_));
 sg13g2_mux2_1 _19303_ (.A0(net3363),
    .A1(net5794),
    .S(_03129_),
    .X(_00539_));
 sg13g2_mux2_1 _19304_ (.A0(net3598),
    .A1(net5768),
    .S(_03129_),
    .X(_00540_));
 sg13g2_mux2_1 _19305_ (.A0(net3234),
    .A1(net5738),
    .S(_03129_),
    .X(_00541_));
 sg13g2_mux2_1 _19306_ (.A0(net3634),
    .A1(net5708),
    .S(_03129_),
    .X(_00542_));
 sg13g2_mux2_1 _19307_ (.A0(net3613),
    .A1(net5681),
    .S(_03129_),
    .X(_00543_));
 sg13g2_mux2_1 _19308_ (.A0(net3258),
    .A1(net5650),
    .S(_03129_),
    .X(_00544_));
 sg13g2_mux2_1 _19309_ (.A0(net3625),
    .A1(net5624),
    .S(_03129_),
    .X(_00545_));
 sg13g2_nand2_2 _19310_ (.Y(_03130_),
    .A(_10383_),
    .B(net5419));
 sg13g2_mux2_1 _19311_ (.A0(net5776),
    .A1(net6895),
    .S(_03130_),
    .X(_00546_));
 sg13g2_mux2_1 _19312_ (.A0(net5750),
    .A1(net6485),
    .S(_03130_),
    .X(_00547_));
 sg13g2_mux2_1 _19313_ (.A0(net5718),
    .A1(net6551),
    .S(_03130_),
    .X(_00548_));
 sg13g2_mux2_1 _19314_ (.A0(net5691),
    .A1(net6294),
    .S(_03130_),
    .X(_00549_));
 sg13g2_mux2_1 _19315_ (.A0(net5661),
    .A1(net6894),
    .S(_03130_),
    .X(_00550_));
 sg13g2_mux2_1 _19316_ (.A0(net5631),
    .A1(net6462),
    .S(_03130_),
    .X(_00551_));
 sg13g2_mux2_1 _19317_ (.A0(net5604),
    .A1(net6463),
    .S(_03130_),
    .X(_00552_));
 sg13g2_and2_2 _19318_ (.A(_03074_),
    .B(_03078_),
    .X(_03131_));
 sg13g2_mux2_1 _19319_ (.A0(net3481),
    .A1(net5795),
    .S(_03131_),
    .X(_00553_));
 sg13g2_mux2_1 _19320_ (.A0(net3600),
    .A1(net5768),
    .S(_03131_),
    .X(_00554_));
 sg13g2_mux2_1 _19321_ (.A0(net3285),
    .A1(net5738),
    .S(_03131_),
    .X(_00555_));
 sg13g2_mux2_1 _19322_ (.A0(net4029),
    .A1(net5708),
    .S(_03131_),
    .X(_00556_));
 sg13g2_mux2_1 _19323_ (.A0(net3592),
    .A1(net5681),
    .S(_03131_),
    .X(_00557_));
 sg13g2_mux2_1 _19324_ (.A0(net3567),
    .A1(net5650),
    .S(_03131_),
    .X(_00558_));
 sg13g2_mux2_1 _19325_ (.A0(net3620),
    .A1(net5624),
    .S(_03131_),
    .X(_00559_));
 sg13g2_nand2_2 _19326_ (.Y(_03132_),
    .A(_10383_),
    .B(net5416));
 sg13g2_mux2_1 _19327_ (.A0(net5776),
    .A1(net6964),
    .S(_03132_),
    .X(_00560_));
 sg13g2_mux2_1 _19328_ (.A0(net5749),
    .A1(net4512),
    .S(_03132_),
    .X(_00561_));
 sg13g2_mux2_1 _19329_ (.A0(net5718),
    .A1(net6334),
    .S(_03132_),
    .X(_00562_));
 sg13g2_mux2_1 _19330_ (.A0(net5691),
    .A1(net4471),
    .S(_03132_),
    .X(_00563_));
 sg13g2_mux2_1 _19331_ (.A0(net5661),
    .A1(net6608),
    .S(_03132_),
    .X(_00564_));
 sg13g2_mux2_1 _19332_ (.A0(net5631),
    .A1(net6396),
    .S(_03132_),
    .X(_00565_));
 sg13g2_mux2_1 _19333_ (.A0(net5604),
    .A1(net6861),
    .S(_03132_),
    .X(_00566_));
 sg13g2_nand2_2 _19334_ (.Y(_03133_),
    .A(_10497_),
    .B(_03078_));
 sg13g2_nor2_1 _19335_ (.A(net5795),
    .B(_03133_),
    .Y(_03134_));
 sg13g2_a21oi_1 _19336_ (.A1(_08128_),
    .A2(_03133_),
    .Y(_00567_),
    .B1(_03134_));
 sg13g2_mux2_1 _19337_ (.A0(net5768),
    .A1(net6912),
    .S(_03133_),
    .X(_00568_));
 sg13g2_mux2_1 _19338_ (.A0(net5739),
    .A1(net6873),
    .S(_03133_),
    .X(_00569_));
 sg13g2_mux2_1 _19339_ (.A0(net5708),
    .A1(net6647),
    .S(_03133_),
    .X(_00570_));
 sg13g2_mux2_1 _19340_ (.A0(net5681),
    .A1(net6444),
    .S(_03133_),
    .X(_00571_));
 sg13g2_mux2_1 _19341_ (.A0(net5650),
    .A1(net6796),
    .S(_03133_),
    .X(_00572_));
 sg13g2_mux2_1 _19342_ (.A0(net5624),
    .A1(net6699),
    .S(_03133_),
    .X(_00573_));
 sg13g2_nand2_2 _19343_ (.Y(_03135_),
    .A(_10383_),
    .B(net5424));
 sg13g2_mux2_1 _19344_ (.A0(net5776),
    .A1(net4374),
    .S(_03135_),
    .X(_00574_));
 sg13g2_mux2_1 _19345_ (.A0(net5749),
    .A1(net4416),
    .S(_03135_),
    .X(_00575_));
 sg13g2_mux2_1 _19346_ (.A0(net5715),
    .A1(net6683),
    .S(_03135_),
    .X(_00576_));
 sg13g2_mux2_1 _19347_ (.A0(net5691),
    .A1(net4434),
    .S(_03135_),
    .X(_00577_));
 sg13g2_mux2_1 _19348_ (.A0(net5661),
    .A1(net4307),
    .S(_03135_),
    .X(_00578_));
 sg13g2_mux2_1 _19349_ (.A0(net5631),
    .A1(net6163),
    .S(_03135_),
    .X(_00579_));
 sg13g2_mux2_1 _19350_ (.A0(net5604),
    .A1(net6648),
    .S(_03135_),
    .X(_00580_));
 sg13g2_nor2_2 _19351_ (.A(net5473),
    .B(net5414),
    .Y(_03136_));
 sg13g2_mux2_1 _19352_ (.A0(net3828),
    .A1(net5793),
    .S(_03136_),
    .X(_00581_));
 sg13g2_mux2_1 _19353_ (.A0(net3227),
    .A1(net5758),
    .S(_03136_),
    .X(_00582_));
 sg13g2_mux2_1 _19354_ (.A0(net3236),
    .A1(net5728),
    .S(_03136_),
    .X(_00583_));
 sg13g2_mux2_1 _19355_ (.A0(net3424),
    .A1(net5701),
    .S(_03136_),
    .X(_00584_));
 sg13g2_mux2_1 _19356_ (.A0(net3574),
    .A1(net5671),
    .S(_03136_),
    .X(_00585_));
 sg13g2_mux2_1 _19357_ (.A0(net3432),
    .A1(net5646),
    .S(_03136_),
    .X(_00586_));
 sg13g2_mux2_1 _19358_ (.A0(net4002),
    .A1(net5612),
    .S(_03136_),
    .X(_00587_));
 sg13g2_nand2_2 _19359_ (.Y(_03137_),
    .A(net5420),
    .B(_03076_));
 sg13g2_mux2_1 _19360_ (.A0(net5784),
    .A1(net6131),
    .S(_03137_),
    .X(_00588_));
 sg13g2_mux2_1 _19361_ (.A0(net5761),
    .A1(net6532),
    .S(_03137_),
    .X(_00589_));
 sg13g2_mux2_1 _19362_ (.A0(net5732),
    .A1(net6541),
    .S(_03137_),
    .X(_00590_));
 sg13g2_mux2_1 _19363_ (.A0(net5703),
    .A1(net6486),
    .S(_03137_),
    .X(_00591_));
 sg13g2_mux2_1 _19364_ (.A0(net5677),
    .A1(net6609),
    .S(_03137_),
    .X(_00592_));
 sg13g2_mux2_1 _19365_ (.A0(net5643),
    .A1(net6545),
    .S(_03137_),
    .X(_00593_));
 sg13g2_mux2_1 _19366_ (.A0(net5618),
    .A1(net6932),
    .S(_03137_),
    .X(_00594_));
 sg13g2_nand2_2 _19367_ (.Y(_03138_),
    .A(net5420),
    .B(_03118_));
 sg13g2_mux2_1 _19368_ (.A0(net5784),
    .A1(net6674),
    .S(_03138_),
    .X(_00595_));
 sg13g2_mux2_1 _19369_ (.A0(net5761),
    .A1(net6880),
    .S(_03138_),
    .X(_00596_));
 sg13g2_mux2_1 _19370_ (.A0(net5732),
    .A1(net6772),
    .S(_03138_),
    .X(_00597_));
 sg13g2_mux2_1 _19371_ (.A0(net5702),
    .A1(net6216),
    .S(_03138_),
    .X(_00598_));
 sg13g2_mux2_1 _19372_ (.A0(net5677),
    .A1(net6955),
    .S(_03138_),
    .X(_00599_));
 sg13g2_mux2_1 _19373_ (.A0(net5643),
    .A1(net6693),
    .S(_03138_),
    .X(_00600_));
 sg13g2_mux2_1 _19374_ (.A0(net5618),
    .A1(net6194),
    .S(_03138_),
    .X(_00601_));
 sg13g2_nand2_2 _19375_ (.Y(_03139_),
    .A(_10372_),
    .B(net5420));
 sg13g2_mux2_1 _19376_ (.A0(net5784),
    .A1(net4329),
    .S(_03139_),
    .X(_00602_));
 sg13g2_mux2_1 _19377_ (.A0(net5761),
    .A1(net6731),
    .S(_03139_),
    .X(_00603_));
 sg13g2_mux2_1 _19378_ (.A0(net5732),
    .A1(net4330),
    .S(_03139_),
    .X(_00604_));
 sg13g2_mux2_1 _19379_ (.A0(net5702),
    .A1(net6246),
    .S(_03139_),
    .X(_00605_));
 sg13g2_mux2_1 _19380_ (.A0(net5677),
    .A1(net6909),
    .S(_03139_),
    .X(_00606_));
 sg13g2_mux2_1 _19381_ (.A0(net5643),
    .A1(net4469),
    .S(_03139_),
    .X(_00607_));
 sg13g2_mux2_1 _19382_ (.A0(net5618),
    .A1(net6639),
    .S(_03139_),
    .X(_00608_));
 sg13g2_nand2_2 _19383_ (.Y(_03140_),
    .A(net5420),
    .B(net5411));
 sg13g2_mux2_1 _19384_ (.A0(net5785),
    .A1(net6292),
    .S(_03140_),
    .X(_00609_));
 sg13g2_mux2_1 _19385_ (.A0(net5761),
    .A1(net6043),
    .S(_03140_),
    .X(_00610_));
 sg13g2_mux2_1 _19386_ (.A0(net5732),
    .A1(net6152),
    .S(_03140_),
    .X(_00611_));
 sg13g2_mux2_1 _19387_ (.A0(net5702),
    .A1(net4352),
    .S(_03140_),
    .X(_00612_));
 sg13g2_mux2_1 _19388_ (.A0(net5677),
    .A1(net6763),
    .S(_03140_),
    .X(_00613_));
 sg13g2_mux2_1 _19389_ (.A0(net5643),
    .A1(net6277),
    .S(_03140_),
    .X(_00614_));
 sg13g2_mux2_1 _19390_ (.A0(net5618),
    .A1(net6443),
    .S(_03140_),
    .X(_00615_));
 sg13g2_nand2_2 _19391_ (.Y(_03141_),
    .A(net5470),
    .B(_03074_));
 sg13g2_mux2_1 _19392_ (.A0(net5787),
    .A1(net6847),
    .S(_03141_),
    .X(_00616_));
 sg13g2_mux2_1 _19393_ (.A0(net5754),
    .A1(net6317),
    .S(_03141_),
    .X(_00617_));
 sg13g2_mux2_1 _19394_ (.A0(net5725),
    .A1(net6834),
    .S(_03141_),
    .X(_00618_));
 sg13g2_mux2_1 _19395_ (.A0(net5705),
    .A1(net6587),
    .S(_03141_),
    .X(_00619_));
 sg13g2_mux2_1 _19396_ (.A0(net5668),
    .A1(net6349),
    .S(_03141_),
    .X(_00620_));
 sg13g2_mux2_1 _19397_ (.A0(net5641),
    .A1(net6908),
    .S(_03141_),
    .X(_00621_));
 sg13g2_mux2_1 _19398_ (.A0(net5613),
    .A1(net7051),
    .S(_03141_),
    .X(_00622_));
 sg13g2_nand2_2 _19399_ (.Y(_03142_),
    .A(net5421),
    .B(_03113_));
 sg13g2_mux2_1 _19400_ (.A0(net5785),
    .A1(net6081),
    .S(_03142_),
    .X(_00623_));
 sg13g2_mux2_1 _19401_ (.A0(net5761),
    .A1(net4516),
    .S(_03142_),
    .X(_00624_));
 sg13g2_mux2_1 _19402_ (.A0(net5730),
    .A1(net6305),
    .S(_03142_),
    .X(_00625_));
 sg13g2_mux2_1 _19403_ (.A0(net5705),
    .A1(net4458),
    .S(_03142_),
    .X(_00626_));
 sg13g2_mux2_1 _19404_ (.A0(net5675),
    .A1(net6668),
    .S(_03142_),
    .X(_00627_));
 sg13g2_mux2_1 _19405_ (.A0(net5642),
    .A1(net6245),
    .S(_03142_),
    .X(_00628_));
 sg13g2_mux2_1 _19406_ (.A0(net5616),
    .A1(net6780),
    .S(_03142_),
    .X(_00629_));
 sg13g2_nand2_2 _19407_ (.Y(_03143_),
    .A(net5421),
    .B(net5419));
 sg13g2_mux2_1 _19408_ (.A0(net5784),
    .A1(net6604),
    .S(_03143_),
    .X(_00630_));
 sg13g2_mux2_1 _19409_ (.A0(net5763),
    .A1(net6231),
    .S(_03143_),
    .X(_00631_));
 sg13g2_mux2_1 _19410_ (.A0(net5732),
    .A1(net6402),
    .S(_03143_),
    .X(_00632_));
 sg13g2_mux2_1 _19411_ (.A0(net5703),
    .A1(net6839),
    .S(_03143_),
    .X(_00633_));
 sg13g2_mux2_1 _19412_ (.A0(net5677),
    .A1(net6212),
    .S(_03143_),
    .X(_00634_));
 sg13g2_mux2_1 _19413_ (.A0(net5643),
    .A1(net4257),
    .S(_03143_),
    .X(_00635_));
 sg13g2_mux2_1 _19414_ (.A0(net5618),
    .A1(net6798),
    .S(_03143_),
    .X(_00636_));
 sg13g2_nand2_2 _19415_ (.Y(_03144_),
    .A(net5421),
    .B(net5416));
 sg13g2_mux2_1 _19416_ (.A0(net5786),
    .A1(net6654),
    .S(_03144_),
    .X(_00637_));
 sg13g2_mux2_1 _19417_ (.A0(net5763),
    .A1(net4244),
    .S(_03144_),
    .X(_00638_));
 sg13g2_mux2_1 _19418_ (.A0(net5732),
    .A1(net6739),
    .S(_03144_),
    .X(_00639_));
 sg13g2_mux2_1 _19419_ (.A0(net5703),
    .A1(net4481),
    .S(_03144_),
    .X(_00640_));
 sg13g2_mux2_1 _19420_ (.A0(net5677),
    .A1(net6375),
    .S(_03144_),
    .X(_00641_));
 sg13g2_mux2_1 _19421_ (.A0(net5643),
    .A1(net6084),
    .S(_03144_),
    .X(_00642_));
 sg13g2_mux2_1 _19422_ (.A0(net5618),
    .A1(net6629),
    .S(_03144_),
    .X(_00643_));
 sg13g2_nand2_2 _19423_ (.Y(_03145_),
    .A(_10497_),
    .B(net5421));
 sg13g2_mux2_1 _19424_ (.A0(net5786),
    .A1(net6187),
    .S(_03145_),
    .X(_00644_));
 sg13g2_mux2_1 _19425_ (.A0(net5763),
    .A1(net6248),
    .S(_03145_),
    .X(_00645_));
 sg13g2_mux2_1 _19426_ (.A0(net5732),
    .A1(net6350),
    .S(_03145_),
    .X(_00646_));
 sg13g2_mux2_1 _19427_ (.A0(net5703),
    .A1(net6415),
    .S(_03145_),
    .X(_00647_));
 sg13g2_mux2_1 _19428_ (.A0(net5677),
    .A1(net6525),
    .S(_03145_),
    .X(_00648_));
 sg13g2_mux2_1 _19429_ (.A0(net5643),
    .A1(net4466),
    .S(_03145_),
    .X(_00649_));
 sg13g2_mux2_1 _19430_ (.A0(net5618),
    .A1(net6077),
    .S(_03145_),
    .X(_00650_));
 sg13g2_nor2b_2 _19431_ (.A(net5473),
    .B_N(net5470),
    .Y(_03146_));
 sg13g2_mux2_1 _19432_ (.A0(net3265),
    .A1(net5783),
    .S(_03146_),
    .X(_00651_));
 sg13g2_mux2_1 _19433_ (.A0(net3192),
    .A1(net5754),
    .S(_03146_),
    .X(_00652_));
 sg13g2_mux2_1 _19434_ (.A0(net3312),
    .A1(net5725),
    .S(_03146_),
    .X(_00653_));
 sg13g2_mux2_1 _19435_ (.A0(net3691),
    .A1(net5696),
    .S(_03146_),
    .X(_00654_));
 sg13g2_mux2_1 _19436_ (.A0(net3636),
    .A1(net5667),
    .S(_03146_),
    .X(_00655_));
 sg13g2_mux2_1 _19437_ (.A0(net3278),
    .A1(net5641),
    .S(_03146_),
    .X(_00656_));
 sg13g2_mux2_1 _19438_ (.A0(net3616),
    .A1(net5610),
    .S(_03146_),
    .X(_00657_));
 sg13g2_nor2_2 _19439_ (.A(_10384_),
    .B(net5471),
    .Y(_03147_));
 sg13g2_mux2_1 _19440_ (.A0(net3393),
    .A1(net5779),
    .S(_03147_),
    .X(_00658_));
 sg13g2_mux2_1 _19441_ (.A0(net3453),
    .A1(net5749),
    .S(_03147_),
    .X(_00659_));
 sg13g2_mux2_1 _19442_ (.A0(net3140),
    .A1(net5719),
    .S(_03147_),
    .X(_00660_));
 sg13g2_mux2_1 _19443_ (.A0(net3935),
    .A1(net5686),
    .S(_03147_),
    .X(_00661_));
 sg13g2_mux2_1 _19444_ (.A0(net3214),
    .A1(net5656),
    .S(_03147_),
    .X(_00662_));
 sg13g2_mux2_1 _19445_ (.A0(net3741),
    .A1(net5635),
    .S(_03147_),
    .X(_00663_));
 sg13g2_mux2_1 _19446_ (.A0(net3948),
    .A1(net5599),
    .S(_03147_),
    .X(_00664_));
 sg13g2_nor2_2 _19447_ (.A(_10384_),
    .B(net5467),
    .Y(_03148_));
 sg13g2_mux2_1 _19448_ (.A0(net3523),
    .A1(net5779),
    .S(_03148_),
    .X(_00665_));
 sg13g2_mux2_1 _19449_ (.A0(net3864),
    .A1(net5749),
    .S(_03148_),
    .X(_00666_));
 sg13g2_mux2_1 _19450_ (.A0(net3451),
    .A1(net5719),
    .S(_03148_),
    .X(_00667_));
 sg13g2_mux2_1 _19451_ (.A0(net4036),
    .A1(net5686),
    .S(_03148_),
    .X(_00668_));
 sg13g2_mux2_1 _19452_ (.A0(net3770),
    .A1(net5683),
    .S(_03148_),
    .X(_00669_));
 sg13g2_mux2_1 _19453_ (.A0(net3302),
    .A1(net5635),
    .S(_03148_),
    .X(_00670_));
 sg13g2_mux2_1 _19454_ (.A0(net3731),
    .A1(net5599),
    .S(_03148_),
    .X(_00671_));
 sg13g2_nand2_2 _19455_ (.Y(_03149_),
    .A(_10383_),
    .B(net5468));
 sg13g2_mux2_1 _19456_ (.A0(net5779),
    .A1(net6616),
    .S(_03149_),
    .X(_00672_));
 sg13g2_mux2_1 _19457_ (.A0(net5744),
    .A1(net6230),
    .S(_03149_),
    .X(_00673_));
 sg13g2_mux2_1 _19458_ (.A0(net5714),
    .A1(net6959),
    .S(_03149_),
    .X(_00674_));
 sg13g2_mux2_1 _19459_ (.A0(net5686),
    .A1(net6784),
    .S(_03149_),
    .X(_00675_));
 sg13g2_mux2_1 _19460_ (.A0(net5656),
    .A1(net6632),
    .S(_03149_),
    .X(_00676_));
 sg13g2_mux2_1 _19461_ (.A0(net5635),
    .A1(net6287),
    .S(_03149_),
    .X(_00677_));
 sg13g2_mux2_1 _19462_ (.A0(net5599),
    .A1(net6840),
    .S(_03149_),
    .X(_00678_));
 sg13g2_nor2_2 _19463_ (.A(net5430),
    .B(_10479_),
    .Y(_03150_));
 sg13g2_mux2_1 _19464_ (.A0(net3301),
    .A1(net5776),
    .S(_03150_),
    .X(_00679_));
 sg13g2_mux2_1 _19465_ (.A0(net3779),
    .A1(net5749),
    .S(_03150_),
    .X(_00680_));
 sg13g2_mux2_1 _19466_ (.A0(net3337),
    .A1(net5720),
    .S(_03150_),
    .X(_00681_));
 sg13g2_mux2_1 _19467_ (.A0(net3514),
    .A1(net5691),
    .S(_03150_),
    .X(_00682_));
 sg13g2_mux2_1 _19468_ (.A0(net3645),
    .A1(net5662),
    .S(_03150_),
    .X(_00683_));
 sg13g2_mux2_1 _19469_ (.A0(net3719),
    .A1(net5636),
    .S(_03150_),
    .X(_00684_));
 sg13g2_mux2_1 _19470_ (.A0(net3389),
    .A1(net5604),
    .S(_03150_),
    .X(_00685_));
 sg13g2_nand2_2 _19471_ (.Y(_03151_),
    .A(net5431),
    .B(net5412));
 sg13g2_mux2_1 _19472_ (.A0(net5774),
    .A1(net6579),
    .S(_03151_),
    .X(_00686_));
 sg13g2_mux2_1 _19473_ (.A0(net5745),
    .A1(net6452),
    .S(_03151_),
    .X(_00687_));
 sg13g2_mux2_1 _19474_ (.A0(net5716),
    .A1(net6380),
    .S(_03151_),
    .X(_00688_));
 sg13g2_mux2_1 _19475_ (.A0(net5690),
    .A1(net6725),
    .S(_03151_),
    .X(_00689_));
 sg13g2_mux2_1 _19476_ (.A0(net5655),
    .A1(net6806),
    .S(_03151_),
    .X(_00690_));
 sg13g2_mux2_1 _19477_ (.A0(net5629),
    .A1(net6384),
    .S(_03151_),
    .X(_00691_));
 sg13g2_mux2_1 _19478_ (.A0(net5597),
    .A1(net6190),
    .S(_03151_),
    .X(_00692_));
 sg13g2_nand2_2 _19479_ (.Y(_03152_),
    .A(net5431),
    .B(_10381_));
 sg13g2_mux2_1 _19480_ (.A0(net5774),
    .A1(net6301),
    .S(_03152_),
    .X(_00693_));
 sg13g2_mux2_1 _19481_ (.A0(net5745),
    .A1(net4527),
    .S(_03152_),
    .X(_00694_));
 sg13g2_mux2_1 _19482_ (.A0(net5716),
    .A1(net6362),
    .S(_03152_),
    .X(_00695_));
 sg13g2_mux2_1 _19483_ (.A0(net5690),
    .A1(net4305),
    .S(_03152_),
    .X(_00696_));
 sg13g2_mux2_1 _19484_ (.A0(net5661),
    .A1(net6489),
    .S(_03152_),
    .X(_00697_));
 sg13g2_mux2_1 _19485_ (.A0(net5628),
    .A1(net6557),
    .S(_03152_),
    .X(_00698_));
 sg13g2_mux2_1 _19486_ (.A0(net5600),
    .A1(net6272),
    .S(_03152_),
    .X(_00699_));
 sg13g2_nand2_2 _19487_ (.Y(_03153_),
    .A(net5416),
    .B(_03104_));
 sg13g2_mux2_1 _19488_ (.A0(net5786),
    .A1(net6182),
    .S(_03153_),
    .X(_00700_));
 sg13g2_mux2_1 _19489_ (.A0(net5764),
    .A1(net6498),
    .S(_03153_),
    .X(_00701_));
 sg13g2_mux2_1 _19490_ (.A0(net5733),
    .A1(net6147),
    .S(_03153_),
    .X(_00702_));
 sg13g2_mux2_1 _19491_ (.A0(net5704),
    .A1(net6732),
    .S(_03153_),
    .X(_00703_));
 sg13g2_mux2_1 _19492_ (.A0(net5678),
    .A1(net6705),
    .S(_03153_),
    .X(_00704_));
 sg13g2_mux2_1 _19493_ (.A0(net5644),
    .A1(net4301),
    .S(_03153_),
    .X(_00705_));
 sg13g2_mux2_1 _19494_ (.A0(net5619),
    .A1(net4308),
    .S(_03153_),
    .X(_00706_));
 sg13g2_nand2_2 _19495_ (.Y(_03154_),
    .A(net5432),
    .B(_03076_));
 sg13g2_mux2_1 _19496_ (.A0(net5774),
    .A1(net6857),
    .S(_03154_),
    .X(_00707_));
 sg13g2_mux2_1 _19497_ (.A0(net5747),
    .A1(net6379),
    .S(_03154_),
    .X(_00708_));
 sg13g2_mux2_1 _19498_ (.A0(net5717),
    .A1(net6123),
    .S(_03154_),
    .X(_00709_));
 sg13g2_mux2_1 _19499_ (.A0(net5689),
    .A1(net6742),
    .S(_03154_),
    .X(_00710_));
 sg13g2_mux2_1 _19500_ (.A0(net5659),
    .A1(net6184),
    .S(_03154_),
    .X(_00711_));
 sg13g2_mux2_1 _19501_ (.A0(net5628),
    .A1(net6316),
    .S(_03154_),
    .X(_00712_));
 sg13g2_mux2_1 _19502_ (.A0(net5601),
    .A1(net6711),
    .S(_03154_),
    .X(_00713_));
 sg13g2_nand2_2 _19503_ (.Y(_03155_),
    .A(net5431),
    .B(net5468));
 sg13g2_mux2_1 _19504_ (.A0(net5771),
    .A1(net4293),
    .S(_03155_),
    .X(_00714_));
 sg13g2_mux2_1 _19505_ (.A0(net5742),
    .A1(net4164),
    .S(_03155_),
    .X(_00715_));
 sg13g2_mux2_1 _19506_ (.A0(net5713),
    .A1(net6531),
    .S(_03155_),
    .X(_00716_));
 sg13g2_mux2_1 _19507_ (.A0(net5684),
    .A1(net6644),
    .S(_03155_),
    .X(_00717_));
 sg13g2_mux2_1 _19508_ (.A0(net5655),
    .A1(net4267),
    .S(_03155_),
    .X(_00718_));
 sg13g2_mux2_1 _19509_ (.A0(net5626),
    .A1(net6623),
    .S(_03155_),
    .X(_00719_));
 sg13g2_mux2_1 _19510_ (.A0(net5597),
    .A1(net6930),
    .S(_03155_),
    .X(_00720_));
 sg13g2_nand2_2 _19511_ (.Y(_03156_),
    .A(_10480_),
    .B(net5416));
 sg13g2_mux2_1 _19512_ (.A0(net5791),
    .A1(net6254),
    .S(_03156_),
    .X(_00721_));
 sg13g2_mux2_1 _19513_ (.A0(net5751),
    .A1(net6738),
    .S(_03156_),
    .X(_00722_));
 sg13g2_mux2_1 _19514_ (.A0(net5720),
    .A1(net6950),
    .S(_03156_),
    .X(_00723_));
 sg13g2_mux2_1 _19515_ (.A0(net5699),
    .A1(net6788),
    .S(_03156_),
    .X(_00724_));
 sg13g2_mux2_1 _19516_ (.A0(net5663),
    .A1(net6603),
    .S(_03156_),
    .X(_00725_));
 sg13g2_mux2_1 _19517_ (.A0(net5637),
    .A1(net6416),
    .S(_03156_),
    .X(_00726_));
 sg13g2_mux2_1 _19518_ (.A0(net5605),
    .A1(net6405),
    .S(_03156_),
    .X(_00727_));
 sg13g2_nand2_2 _19519_ (.Y(_03157_),
    .A(net5422),
    .B(_03076_));
 sg13g2_mux2_1 _19520_ (.A0(net5781),
    .A1(net6726),
    .S(_03157_),
    .X(_00728_));
 sg13g2_mux2_1 _19521_ (.A0(net5752),
    .A1(net6058),
    .S(_03157_),
    .X(_00729_));
 sg13g2_mux2_1 _19522_ (.A0(net5722),
    .A1(net6829),
    .S(_03157_),
    .X(_00730_));
 sg13g2_mux2_1 _19523_ (.A0(net5693),
    .A1(net6156),
    .S(_03157_),
    .X(_00731_));
 sg13g2_mux2_1 _19524_ (.A0(net5665),
    .A1(net6493),
    .S(_03157_),
    .X(_00732_));
 sg13g2_mux2_1 _19525_ (.A0(net5638),
    .A1(net4530),
    .S(_03157_),
    .X(_00733_));
 sg13g2_mux2_1 _19526_ (.A0(net5607),
    .A1(net6701),
    .S(_03157_),
    .X(_00734_));
 sg13g2_nor3_2 _19527_ (.A(net5036),
    .B(net5021),
    .C(net4774),
    .Y(_03158_));
 sg13g2_nor2_2 _19528_ (.A(_08580_),
    .B(_03008_),
    .Y(_03159_));
 sg13g2_nand2_2 _19529_ (.Y(_03160_),
    .A(net4763),
    .B(net4737));
 sg13g2_mux2_1 _19530_ (.A0(net5253),
    .A1(net6454),
    .S(_03160_),
    .X(_00735_));
 sg13g2_mux2_1 _19531_ (.A0(net5223),
    .A1(net6844),
    .S(_03160_),
    .X(_00736_));
 sg13g2_mux2_1 _19532_ (.A0(net5119),
    .A1(net4085),
    .S(_03160_),
    .X(_00737_));
 sg13g2_mux2_1 _19533_ (.A0(net5096),
    .A1(net4363),
    .S(_03160_),
    .X(_00738_));
 sg13g2_mux2_1 _19534_ (.A0(net5189),
    .A1(net4290),
    .S(_03160_),
    .X(_00739_));
 sg13g2_mux2_1 _19535_ (.A0(net5164),
    .A1(net4080),
    .S(_03160_),
    .X(_00740_));
 sg13g2_mux2_1 _19536_ (.A0(net5069),
    .A1(net4037),
    .S(_03160_),
    .X(_00741_));
 sg13g2_mux2_1 _19537_ (.A0(net5046),
    .A1(net6935),
    .S(_03160_),
    .X(_00742_));
 sg13g2_nor2_2 _19538_ (.A(_10502_),
    .B(net5467),
    .Y(_03161_));
 sg13g2_mux2_1 _19539_ (.A0(net3386),
    .A1(net5784),
    .S(_03161_),
    .X(_00743_));
 sg13g2_mux2_1 _19540_ (.A0(net3347),
    .A1(net5763),
    .S(_03161_),
    .X(_00744_));
 sg13g2_mux2_1 _19541_ (.A0(net3135),
    .A1(net5730),
    .S(_03161_),
    .X(_00745_));
 sg13g2_mux2_1 _19542_ (.A0(net3356),
    .A1(net5702),
    .S(_03161_),
    .X(_00746_));
 sg13g2_mux2_1 _19543_ (.A0(net3399),
    .A1(net5675),
    .S(_03161_),
    .X(_00747_));
 sg13g2_mux2_1 _19544_ (.A0(net3194),
    .A1(net5642),
    .S(_03161_),
    .X(_00748_));
 sg13g2_mux2_1 _19545_ (.A0(net3338),
    .A1(net5616),
    .S(_03161_),
    .X(_00749_));
 sg13g2_nand2_2 _19546_ (.Y(_03162_),
    .A(net5421),
    .B(_03100_));
 sg13g2_mux2_1 _19547_ (.A0(net5786),
    .A1(net6848),
    .S(_03162_),
    .X(_00750_));
 sg13g2_mux2_1 _19548_ (.A0(net5763),
    .A1(net6460),
    .S(_03162_),
    .X(_00751_));
 sg13g2_mux2_1 _19549_ (.A0(net5732),
    .A1(net6850),
    .S(_03162_),
    .X(_00752_));
 sg13g2_mux2_1 _19550_ (.A0(net5703),
    .A1(net4487),
    .S(_03162_),
    .X(_00753_));
 sg13g2_mux2_1 _19551_ (.A0(net5677),
    .A1(net6755),
    .S(_03162_),
    .X(_00754_));
 sg13g2_mux2_1 _19552_ (.A0(net5643),
    .A1(net6810),
    .S(_03162_),
    .X(_00755_));
 sg13g2_mux2_1 _19553_ (.A0(net5618),
    .A1(net6353),
    .S(_03162_),
    .X(_00756_));
 sg13g2_nor2_2 _19554_ (.A(net4780),
    .B(net5022),
    .Y(_03163_));
 sg13g2_nand2_2 _19555_ (.Y(_03164_),
    .A(_08631_),
    .B(net5023));
 sg13g2_nor2_2 _19556_ (.A(net5038),
    .B(_03164_),
    .Y(_03165_));
 sg13g2_nand2_2 _19557_ (.Y(_03166_),
    .A(net4895),
    .B(net5032));
 sg13g2_nor2_1 _19558_ (.A(_03008_),
    .B(_03166_),
    .Y(_03167_));
 sg13g2_nand2_2 _19559_ (.Y(_03168_),
    .A(_03165_),
    .B(net4735));
 sg13g2_mux2_1 _19560_ (.A0(net5254),
    .A1(net4271),
    .S(_03168_),
    .X(_00757_));
 sg13g2_mux2_1 _19561_ (.A0(net5222),
    .A1(net4115),
    .S(_03168_),
    .X(_00758_));
 sg13g2_mux2_1 _19562_ (.A0(net5118),
    .A1(net6472),
    .S(_03168_),
    .X(_00759_));
 sg13g2_mux2_1 _19563_ (.A0(net5090),
    .A1(net4158),
    .S(_03168_),
    .X(_00760_));
 sg13g2_mux2_1 _19564_ (.A0(net5188),
    .A1(net4192),
    .S(_03168_),
    .X(_00761_));
 sg13g2_mux2_1 _19565_ (.A0(net5162),
    .A1(net6918),
    .S(_03168_),
    .X(_00762_));
 sg13g2_mux2_1 _19566_ (.A0(net5069),
    .A1(net4150),
    .S(_03168_),
    .X(_00763_));
 sg13g2_mux2_1 _19567_ (.A0(net5047),
    .A1(net4484),
    .S(_03168_),
    .X(_00764_));
 sg13g2_nor2_2 _19568_ (.A(net5425),
    .B(_02996_),
    .Y(_03169_));
 sg13g2_mux2_1 _19569_ (.A0(net3376),
    .A1(net5790),
    .S(_03169_),
    .X(_00765_));
 sg13g2_mux2_1 _19570_ (.A0(net3693),
    .A1(net5756),
    .S(_03169_),
    .X(_00766_));
 sg13g2_mux2_1 _19571_ (.A0(net3515),
    .A1(net5722),
    .S(_03169_),
    .X(_00767_));
 sg13g2_mux2_1 _19572_ (.A0(net3422),
    .A1(net5694),
    .S(_03169_),
    .X(_00768_));
 sg13g2_mux2_1 _19573_ (.A0(net3717),
    .A1(net5666),
    .S(_03169_),
    .X(_00769_));
 sg13g2_mux2_1 _19574_ (.A0(net3903),
    .A1(net5640),
    .S(_03169_),
    .X(_00770_));
 sg13g2_mux2_1 _19575_ (.A0(net3190),
    .A1(net5614),
    .S(_03169_),
    .X(_00771_));
 sg13g2_nor2_2 _19576_ (.A(net5471),
    .B(net5414),
    .Y(_03170_));
 sg13g2_mux2_1 _19577_ (.A0(net3714),
    .A1(net5792),
    .S(_03170_),
    .X(_00772_));
 sg13g2_mux2_1 _19578_ (.A0(net3283),
    .A1(net5758),
    .S(_03170_),
    .X(_00773_));
 sg13g2_mux2_1 _19579_ (.A0(net3442),
    .A1(net5729),
    .S(_03170_),
    .X(_00774_));
 sg13g2_mux2_1 _19580_ (.A0(net3200),
    .A1(net5700),
    .S(_03170_),
    .X(_00775_));
 sg13g2_mux2_1 _19581_ (.A0(net3067),
    .A1(net5671),
    .S(_03170_),
    .X(_00776_));
 sg13g2_mux2_1 _19582_ (.A0(net3323),
    .A1(net5647),
    .S(_03170_),
    .X(_00777_));
 sg13g2_mux2_1 _19583_ (.A0(net3818),
    .A1(net5612),
    .S(_03170_),
    .X(_00778_));
 sg13g2_nor2b_2 _19584_ (.A(net5472),
    .B_N(net5418),
    .Y(_03171_));
 sg13g2_mux2_1 _19585_ (.A0(net3591),
    .A1(net5772),
    .S(_03171_),
    .X(_00779_));
 sg13g2_mux2_1 _19586_ (.A0(net3726),
    .A1(net5743),
    .S(_03171_),
    .X(_00780_));
 sg13g2_mux2_1 _19587_ (.A0(net3866),
    .A1(net5714),
    .S(_03171_),
    .X(_00781_));
 sg13g2_mux2_1 _19588_ (.A0(net3964),
    .A1(net5686),
    .S(_03171_),
    .X(_00782_));
 sg13g2_mux2_1 _19589_ (.A0(net3440),
    .A1(net5657),
    .S(_03171_),
    .X(_00783_));
 sg13g2_mux2_1 _19590_ (.A0(net3776),
    .A1(net5634),
    .S(_03171_),
    .X(_00784_));
 sg13g2_mux2_1 _19591_ (.A0(net3220),
    .A1(net5598),
    .S(_03171_),
    .X(_00785_));
 sg13g2_nand2_2 _19592_ (.Y(_03172_),
    .A(_10381_),
    .B(net5469));
 sg13g2_mux2_1 _19593_ (.A0(net5782),
    .A1(net6602),
    .S(_03172_),
    .X(_00786_));
 sg13g2_mux2_1 _19594_ (.A0(net5753),
    .A1(net6383),
    .S(_03172_),
    .X(_00787_));
 sg13g2_mux2_1 _19595_ (.A0(net5724),
    .A1(net6938),
    .S(_03172_),
    .X(_00788_));
 sg13g2_mux2_1 _19596_ (.A0(net5695),
    .A1(net4535),
    .S(_03172_),
    .X(_00789_));
 sg13g2_mux2_1 _19597_ (.A0(net5667),
    .A1(net4355),
    .S(_03172_),
    .X(_00790_));
 sg13g2_mux2_1 _19598_ (.A0(net5639),
    .A1(net6510),
    .S(_03172_),
    .X(_00791_));
 sg13g2_mux2_1 _19599_ (.A0(net5607),
    .A1(net6263),
    .S(_03172_),
    .X(_00792_));
 sg13g2_nand2_2 _19600_ (.Y(_03173_),
    .A(net5468),
    .B(_03081_));
 sg13g2_mux2_1 _19601_ (.A0(net5792),
    .A1(net6469),
    .S(_03173_),
    .X(_00793_));
 sg13g2_mux2_1 _19602_ (.A0(net5757),
    .A1(net6359),
    .S(_03173_),
    .X(_00794_));
 sg13g2_mux2_1 _19603_ (.A0(net5727),
    .A1(net6435),
    .S(_03173_),
    .X(_00795_));
 sg13g2_mux2_1 _19604_ (.A0(net5700),
    .A1(net6491),
    .S(_03173_),
    .X(_00796_));
 sg13g2_mux2_1 _19605_ (.A0(net5670),
    .A1(net4485),
    .S(_03173_),
    .X(_00797_));
 sg13g2_mux2_1 _19606_ (.A0(net5647),
    .A1(net6710),
    .S(_03173_),
    .X(_00798_));
 sg13g2_mux2_1 _19607_ (.A0(net5612),
    .A1(net4348),
    .S(_03173_),
    .X(_00799_));
 sg13g2_nor2b_2 _19608_ (.A(net5471),
    .B_N(net5418),
    .Y(_03174_));
 sg13g2_mux2_1 _19609_ (.A0(net3419),
    .A1(net5772),
    .S(_03174_),
    .X(_00800_));
 sg13g2_mux2_1 _19610_ (.A0(net3367),
    .A1(net5743),
    .S(_03174_),
    .X(_00801_));
 sg13g2_mux2_1 _19611_ (.A0(net3739),
    .A1(net5714),
    .S(_03174_),
    .X(_00802_));
 sg13g2_mux2_1 _19612_ (.A0(net3721),
    .A1(net5686),
    .S(_03174_),
    .X(_00803_));
 sg13g2_mux2_1 _19613_ (.A0(net3678),
    .A1(net5657),
    .S(_03174_),
    .X(_00804_));
 sg13g2_mux2_1 _19614_ (.A0(net3904),
    .A1(net5634),
    .S(_03174_),
    .X(_00805_));
 sg13g2_mux2_1 _19615_ (.A0(net3638),
    .A1(net5598),
    .S(_03174_),
    .X(_00806_));
 sg13g2_nor2_2 _19616_ (.A(_10479_),
    .B(_03082_),
    .Y(_03175_));
 sg13g2_mux2_1 _19617_ (.A0(net3929),
    .A1(net5797),
    .S(_03175_),
    .X(_00807_));
 sg13g2_mux2_1 _19618_ (.A0(net3826),
    .A1(net5758),
    .S(_03175_),
    .X(_00808_));
 sg13g2_mux2_1 _19619_ (.A0(net3260),
    .A1(net5736),
    .S(_03175_),
    .X(_00809_));
 sg13g2_mux2_1 _19620_ (.A0(net3349),
    .A1(net5707),
    .S(_03175_),
    .X(_00810_));
 sg13g2_mux2_1 _19621_ (.A0(net3522),
    .A1(net5672),
    .S(_03175_),
    .X(_00811_));
 sg13g2_mux2_1 _19622_ (.A0(net3546),
    .A1(net5649),
    .S(_03175_),
    .X(_00812_));
 sg13g2_mux2_1 _19623_ (.A0(net3702),
    .A1(net5621),
    .S(_03175_),
    .X(_00813_));
 sg13g2_nor2_2 _19624_ (.A(_10382_),
    .B(net5414),
    .Y(_03176_));
 sg13g2_mux2_1 _19625_ (.A0(net3727),
    .A1(net5797),
    .S(_03176_),
    .X(_00814_));
 sg13g2_mux2_1 _19626_ (.A0(net3936),
    .A1(net5758),
    .S(_03176_),
    .X(_00815_));
 sg13g2_mux2_1 _19627_ (.A0(net3750),
    .A1(net5736),
    .S(_03176_),
    .X(_00816_));
 sg13g2_mux2_1 _19628_ (.A0(net3263),
    .A1(net5707),
    .S(_03176_),
    .X(_00817_));
 sg13g2_mux2_1 _19629_ (.A0(net3999),
    .A1(net5672),
    .S(_03176_),
    .X(_00818_));
 sg13g2_mux2_1 _19630_ (.A0(net3962),
    .A1(net5649),
    .S(_03176_),
    .X(_00819_));
 sg13g2_mux2_1 _19631_ (.A0(net3352),
    .A1(net5621),
    .S(_03176_),
    .X(_00820_));
 sg13g2_nor2b_2 _19632_ (.A(net5467),
    .B_N(net5418),
    .Y(_03177_));
 sg13g2_mux2_1 _19633_ (.A0(net3799),
    .A1(net5772),
    .S(_03177_),
    .X(_00821_));
 sg13g2_mux2_1 _19634_ (.A0(net3535),
    .A1(net5743),
    .S(_03177_),
    .X(_00822_));
 sg13g2_mux2_1 _19635_ (.A0(net3224),
    .A1(net5714),
    .S(_03177_),
    .X(_00823_));
 sg13g2_mux2_1 _19636_ (.A0(net3534),
    .A1(net5686),
    .S(_03177_),
    .X(_00824_));
 sg13g2_mux2_1 _19637_ (.A0(net3373),
    .A1(net5657),
    .S(_03177_),
    .X(_00825_));
 sg13g2_mux2_1 _19638_ (.A0(net3321),
    .A1(net5634),
    .S(_03177_),
    .X(_00826_));
 sg13g2_mux2_1 _19639_ (.A0(net3509),
    .A1(net5598),
    .S(_03177_),
    .X(_00827_));
 sg13g2_nor2_2 _19640_ (.A(_02996_),
    .B(net5414),
    .Y(_03178_));
 sg13g2_mux2_1 _19641_ (.A0(net3502),
    .A1(net5797),
    .S(_03178_),
    .X(_00828_));
 sg13g2_mux2_1 _19642_ (.A0(net3250),
    .A1(net5758),
    .S(_03178_),
    .X(_00829_));
 sg13g2_mux2_1 _19643_ (.A0(net3333),
    .A1(net5736),
    .S(_03178_),
    .X(_00830_));
 sg13g2_mux2_1 _19644_ (.A0(net3346),
    .A1(net5707),
    .S(_03178_),
    .X(_00831_));
 sg13g2_mux2_1 _19645_ (.A0(net3589),
    .A1(net5672),
    .S(_03178_),
    .X(_00832_));
 sg13g2_mux2_1 _19646_ (.A0(net3184),
    .A1(net5649),
    .S(_03178_),
    .X(_00833_));
 sg13g2_mux2_1 _19647_ (.A0(net3564),
    .A1(net5612),
    .S(_03178_),
    .X(_00834_));
 sg13g2_nand2_2 _19648_ (.Y(_03179_),
    .A(_03081_),
    .B(net5412));
 sg13g2_mux2_1 _19649_ (.A0(net5797),
    .A1(net6886),
    .S(_03179_),
    .X(_00835_));
 sg13g2_mux2_1 _19650_ (.A0(net5758),
    .A1(net6413),
    .S(_03179_),
    .X(_00836_));
 sg13g2_mux2_1 _19651_ (.A0(net5736),
    .A1(net6367),
    .S(_03179_),
    .X(_00837_));
 sg13g2_mux2_1 _19652_ (.A0(net5707),
    .A1(net6247),
    .S(_03179_),
    .X(_00838_));
 sg13g2_mux2_1 _19653_ (.A0(net5672),
    .A1(net6864),
    .S(_03179_),
    .X(_00839_));
 sg13g2_mux2_1 _19654_ (.A0(net5649),
    .A1(net6518),
    .S(_03179_),
    .X(_00840_));
 sg13g2_mux2_1 _19655_ (.A0(net5612),
    .A1(net6215),
    .S(_03179_),
    .X(_00841_));
 sg13g2_nand2_2 _19656_ (.Y(_03180_),
    .A(net5468),
    .B(net5418));
 sg13g2_mux2_1 _19657_ (.A0(net5772),
    .A1(net6233),
    .S(_03180_),
    .X(_00842_));
 sg13g2_mux2_1 _19658_ (.A0(net5743),
    .A1(net4366),
    .S(_03180_),
    .X(_00843_));
 sg13g2_mux2_1 _19659_ (.A0(net5714),
    .A1(net6542),
    .S(_03180_),
    .X(_00844_));
 sg13g2_mux2_1 _19660_ (.A0(net5686),
    .A1(net6539),
    .S(_03180_),
    .X(_00845_));
 sg13g2_mux2_1 _19661_ (.A0(net5657),
    .A1(net4368),
    .S(_03180_),
    .X(_00846_));
 sg13g2_mux2_1 _19662_ (.A0(net5634),
    .A1(net6915),
    .S(_03180_),
    .X(_00847_));
 sg13g2_mux2_1 _19663_ (.A0(net5599),
    .A1(net6879),
    .S(_03180_),
    .X(_00848_));
 sg13g2_nor2_2 _19664_ (.A(_03077_),
    .B(net5414),
    .Y(_03181_));
 sg13g2_mux2_1 _19665_ (.A0(net3945),
    .A1(net5793),
    .S(_03181_),
    .X(_00849_));
 sg13g2_mux2_1 _19666_ (.A0(net3783),
    .A1(net5760),
    .S(_03181_),
    .X(_00850_));
 sg13g2_mux2_1 _19667_ (.A0(net4223),
    .A1(net5729),
    .S(_03181_),
    .X(_00851_));
 sg13g2_mux2_1 _19668_ (.A0(net3852),
    .A1(net5700),
    .S(_03181_),
    .X(_00852_));
 sg13g2_mux2_1 _19669_ (.A0(net3584),
    .A1(net5672),
    .S(_03181_),
    .X(_00853_));
 sg13g2_mux2_1 _19670_ (.A0(net3643),
    .A1(net5648),
    .S(_03181_),
    .X(_00854_));
 sg13g2_mux2_1 _19671_ (.A0(net3517),
    .A1(net5615),
    .S(_03181_),
    .X(_00855_));
 sg13g2_nor2_2 _19672_ (.A(net5414),
    .B(_03119_),
    .Y(_03182_));
 sg13g2_mux2_1 _19673_ (.A0(net3504),
    .A1(net5792),
    .S(_03182_),
    .X(_00856_));
 sg13g2_mux2_1 _19674_ (.A0(net3435),
    .A1(net5759),
    .S(_03182_),
    .X(_00857_));
 sg13g2_mux2_1 _19675_ (.A0(net3712),
    .A1(net5729),
    .S(_03182_),
    .X(_00858_));
 sg13g2_mux2_1 _19676_ (.A0(net3297),
    .A1(net5700),
    .S(_03182_),
    .X(_00859_));
 sg13g2_mux2_1 _19677_ (.A0(net3894),
    .A1(net5672),
    .S(_03182_),
    .X(_00860_));
 sg13g2_mux2_1 _19678_ (.A0(net3189),
    .A1(net5648),
    .S(_03182_),
    .X(_00861_));
 sg13g2_mux2_1 _19679_ (.A0(net3695),
    .A1(net5615),
    .S(_03182_),
    .X(_00862_));
 sg13g2_nor4_2 _19680_ (.A(net5807),
    .B(net5801),
    .C(_10182_),
    .Y(_03183_),
    .D(net5467));
 sg13g2_mux2_1 _19681_ (.A0(net3980),
    .A1(net5783),
    .S(_03183_),
    .X(_00863_));
 sg13g2_mux2_1 _19682_ (.A0(net3622),
    .A1(net5754),
    .S(_03183_),
    .X(_00864_));
 sg13g2_mux2_1 _19683_ (.A0(net3486),
    .A1(net5725),
    .S(_03183_),
    .X(_00865_));
 sg13g2_mux2_1 _19684_ (.A0(net3559),
    .A1(net5696),
    .S(_03183_),
    .X(_00866_));
 sg13g2_mux2_1 _19685_ (.A0(net3374),
    .A1(net5667),
    .S(_03183_),
    .X(_00867_));
 sg13g2_mux2_1 _19686_ (.A0(net3547),
    .A1(net5640),
    .S(_03183_),
    .X(_00868_));
 sg13g2_mux2_1 _19687_ (.A0(net3570),
    .A1(net5610),
    .S(_03183_),
    .X(_00869_));
 sg13g2_nor2_2 _19688_ (.A(_10373_),
    .B(_03082_),
    .Y(_03184_));
 sg13g2_mux2_1 _19689_ (.A0(net3599),
    .A1(net5793),
    .S(_03184_),
    .X(_00870_));
 sg13g2_mux2_1 _19690_ (.A0(net3585),
    .A1(net5758),
    .S(_03184_),
    .X(_00871_));
 sg13g2_mux2_1 _19691_ (.A0(net3881),
    .A1(net5728),
    .S(_03184_),
    .X(_00872_));
 sg13g2_mux2_1 _19692_ (.A0(net3178),
    .A1(net5700),
    .S(_03184_),
    .X(_00873_));
 sg13g2_mux2_1 _19693_ (.A0(net3211),
    .A1(net5672),
    .S(_03184_),
    .X(_00874_));
 sg13g2_mux2_1 _19694_ (.A0(net3569),
    .A1(net5648),
    .S(_03184_),
    .X(_00875_));
 sg13g2_mux2_1 _19695_ (.A0(net3307),
    .A1(net5612),
    .S(_03184_),
    .X(_00876_));
 sg13g2_nand2_2 _19696_ (.Y(_03185_),
    .A(_03081_),
    .B(net5411));
 sg13g2_mux2_1 _19697_ (.A0(net5792),
    .A1(net6364),
    .S(_03185_),
    .X(_00877_));
 sg13g2_mux2_1 _19698_ (.A0(net5760),
    .A1(net6867),
    .S(_03185_),
    .X(_00878_));
 sg13g2_mux2_1 _19699_ (.A0(net5728),
    .A1(net6357),
    .S(_03185_),
    .X(_00879_));
 sg13g2_mux2_1 _19700_ (.A0(net5700),
    .A1(net4380),
    .S(_03185_),
    .X(_00880_));
 sg13g2_mux2_1 _19701_ (.A0(net5670),
    .A1(net4319),
    .S(_03185_),
    .X(_00881_));
 sg13g2_mux2_1 _19702_ (.A0(net5648),
    .A1(net6766),
    .S(_03185_),
    .X(_00882_));
 sg13g2_mux2_1 _19703_ (.A0(net5612),
    .A1(net6262),
    .S(_03185_),
    .X(_00883_));
 sg13g2_nand2_2 _19704_ (.Y(_03186_),
    .A(_10381_),
    .B(net5417));
 sg13g2_mux2_1 _19705_ (.A0(net5771),
    .A1(net4302),
    .S(_03186_),
    .X(_00884_));
 sg13g2_mux2_1 _19706_ (.A0(net5742),
    .A1(net6417),
    .S(_03186_),
    .X(_00885_));
 sg13g2_mux2_1 _19707_ (.A0(net5713),
    .A1(net6800),
    .S(_03186_),
    .X(_00886_));
 sg13g2_mux2_1 _19708_ (.A0(net5684),
    .A1(net6794),
    .S(_03186_),
    .X(_00887_));
 sg13g2_mux2_1 _19709_ (.A0(net5655),
    .A1(net6613),
    .S(_03186_),
    .X(_00888_));
 sg13g2_mux2_1 _19710_ (.A0(net5626),
    .A1(net6514),
    .S(_03186_),
    .X(_00889_));
 sg13g2_mux2_1 _19711_ (.A0(net5598),
    .A1(net6197),
    .S(_03186_),
    .X(_00890_));
 sg13g2_nand2_2 _19712_ (.Y(_03187_),
    .A(net5424),
    .B(net5470));
 sg13g2_mux2_1 _19713_ (.A0(net5787),
    .A1(net6107),
    .S(_03187_),
    .X(_00891_));
 sg13g2_mux2_1 _19714_ (.A0(net5754),
    .A1(net6704),
    .S(_03187_),
    .X(_00892_));
 sg13g2_mux2_1 _19715_ (.A0(net5725),
    .A1(net6382),
    .S(_03187_),
    .X(_00893_));
 sg13g2_mux2_1 _19716_ (.A0(net5705),
    .A1(net6428),
    .S(_03187_),
    .X(_00894_));
 sg13g2_mux2_1 _19717_ (.A0(net5668),
    .A1(net6831),
    .S(_03187_),
    .X(_00895_));
 sg13g2_mux2_1 _19718_ (.A0(net5639),
    .A1(net6242),
    .S(_03187_),
    .X(_00896_));
 sg13g2_mux2_1 _19719_ (.A0(net5609),
    .A1(net6530),
    .S(_03187_),
    .X(_00897_));
 sg13g2_nand2_2 _19720_ (.Y(_03188_),
    .A(net5419),
    .B(_03081_));
 sg13g2_mux2_1 _19721_ (.A0(net5791),
    .A1(net6775),
    .S(_03188_),
    .X(_00898_));
 sg13g2_mux2_1 _19722_ (.A0(net5759),
    .A1(net6689),
    .S(_03188_),
    .X(_00899_));
 sg13g2_mux2_1 _19723_ (.A0(net5735),
    .A1(net6718),
    .S(_03188_),
    .X(_00900_));
 sg13g2_mux2_1 _19724_ (.A0(net5706),
    .A1(net6720),
    .S(_03188_),
    .X(_00901_));
 sg13g2_mux2_1 _19725_ (.A0(net5671),
    .A1(net6661),
    .S(_03188_),
    .X(_00902_));
 sg13g2_mux2_1 _19726_ (.A0(net5646),
    .A1(net6746),
    .S(_03188_),
    .X(_00903_));
 sg13g2_mux2_1 _19727_ (.A0(net5613),
    .A1(net4404),
    .S(_03188_),
    .X(_00904_));
 sg13g2_nand2_2 _19728_ (.Y(_03189_),
    .A(_02995_),
    .B(net5417));
 sg13g2_mux2_1 _19729_ (.A0(net5771),
    .A1(net4262),
    .S(_03189_),
    .X(_00905_));
 sg13g2_mux2_1 _19730_ (.A0(net5742),
    .A1(net4439),
    .S(_03189_),
    .X(_00906_));
 sg13g2_mux2_1 _19731_ (.A0(net5713),
    .A1(net6226),
    .S(_03189_),
    .X(_00907_));
 sg13g2_mux2_1 _19732_ (.A0(net5684),
    .A1(net4232),
    .S(_03189_),
    .X(_00908_));
 sg13g2_mux2_1 _19733_ (.A0(net5655),
    .A1(net4397),
    .S(_03189_),
    .X(_00909_));
 sg13g2_mux2_1 _19734_ (.A0(net5626),
    .A1(net6910),
    .S(_03189_),
    .X(_00910_));
 sg13g2_mux2_1 _19735_ (.A0(net5597),
    .A1(net6449),
    .S(_03189_),
    .X(_00911_));
 sg13g2_nand2_2 _19736_ (.Y(_03190_),
    .A(net5416),
    .B(_03081_));
 sg13g2_mux2_1 _19737_ (.A0(net5793),
    .A1(net4288),
    .S(_03190_),
    .X(_00912_));
 sg13g2_mux2_1 _19738_ (.A0(net5759),
    .A1(net6688),
    .S(_03190_),
    .X(_00913_));
 sg13g2_mux2_1 _19739_ (.A0(net5736),
    .A1(net6488),
    .S(_03190_),
    .X(_00914_));
 sg13g2_mux2_1 _19740_ (.A0(net5706),
    .A1(net6562),
    .S(_03190_),
    .X(_00915_));
 sg13g2_mux2_1 _19741_ (.A0(net5671),
    .A1(net6789),
    .S(_03190_),
    .X(_00916_));
 sg13g2_mux2_1 _19742_ (.A0(net5646),
    .A1(net6624),
    .S(_03190_),
    .X(_00917_));
 sg13g2_mux2_1 _19743_ (.A0(net5613),
    .A1(net6278),
    .S(_03190_),
    .X(_00918_));
 sg13g2_nand2_2 _19744_ (.Y(_03191_),
    .A(net5424),
    .B(_03081_));
 sg13g2_mux2_1 _19745_ (.A0(net5790),
    .A1(net4478),
    .S(_03191_),
    .X(_00919_));
 sg13g2_mux2_1 _19746_ (.A0(net5759),
    .A1(net6074),
    .S(_03191_),
    .X(_00920_));
 sg13g2_mux2_1 _19747_ (.A0(net5735),
    .A1(net4511),
    .S(_03191_),
    .X(_00921_));
 sg13g2_mux2_1 _19748_ (.A0(net5706),
    .A1(net6232),
    .S(_03191_),
    .X(_00922_));
 sg13g2_mux2_1 _19749_ (.A0(net5670),
    .A1(net6911),
    .S(_03191_),
    .X(_00923_));
 sg13g2_mux2_1 _19750_ (.A0(net5646),
    .A1(net6783),
    .S(_03191_),
    .X(_00924_));
 sg13g2_mux2_1 _19751_ (.A0(net5613),
    .A1(net6830),
    .S(_03191_),
    .X(_00925_));
 sg13g2_nand2_2 _19752_ (.Y(_03192_),
    .A(net5417),
    .B(net5412));
 sg13g2_mux2_1 _19753_ (.A0(net5771),
    .A1(net4280),
    .S(_03192_),
    .X(_00926_));
 sg13g2_mux2_1 _19754_ (.A0(net5742),
    .A1(net6407),
    .S(_03192_),
    .X(_00927_));
 sg13g2_mux2_1 _19755_ (.A0(net5713),
    .A1(net6637),
    .S(_03192_),
    .X(_00928_));
 sg13g2_mux2_1 _19756_ (.A0(net5684),
    .A1(net6188),
    .S(_03192_),
    .X(_00929_));
 sg13g2_mux2_1 _19757_ (.A0(net5655),
    .A1(net6663),
    .S(_03192_),
    .X(_00930_));
 sg13g2_mux2_1 _19758_ (.A0(net5626),
    .A1(net6995),
    .S(_03192_),
    .X(_00931_));
 sg13g2_mux2_1 _19759_ (.A0(net5597),
    .A1(net6892),
    .S(_03192_),
    .X(_00932_));
 sg13g2_nor2_2 _19760_ (.A(net5473),
    .B(net5413),
    .Y(_03193_));
 sg13g2_mux2_1 _19761_ (.A0(net3342),
    .A1(net5794),
    .S(_03193_),
    .X(_00933_));
 sg13g2_mux2_1 _19762_ (.A0(net3154),
    .A1(net5769),
    .S(_03193_),
    .X(_00934_));
 sg13g2_mux2_1 _19763_ (.A0(net3606),
    .A1(net5738),
    .S(_03193_),
    .X(_00935_));
 sg13g2_mux2_1 _19764_ (.A0(net3284),
    .A1(net5710),
    .S(_03193_),
    .X(_00936_));
 sg13g2_mux2_1 _19765_ (.A0(net3150),
    .A1(net5678),
    .S(_03193_),
    .X(_00937_));
 sg13g2_mux2_1 _19766_ (.A0(net3433),
    .A1(net5650),
    .S(_03193_),
    .X(_00938_));
 sg13g2_mux2_1 _19767_ (.A0(net3877),
    .A1(net5623),
    .S(_03193_),
    .X(_00939_));
 sg13g2_nor2_2 _19768_ (.A(net5471),
    .B(net5413),
    .Y(_03194_));
 sg13g2_mux2_1 _19769_ (.A0(net3577),
    .A1(net5794),
    .S(_03194_),
    .X(_00940_));
 sg13g2_mux2_1 _19770_ (.A0(net3670),
    .A1(net5769),
    .S(_03194_),
    .X(_00941_));
 sg13g2_mux2_1 _19771_ (.A0(net3420),
    .A1(net5738),
    .S(_03194_),
    .X(_00942_));
 sg13g2_mux2_1 _19772_ (.A0(net3774),
    .A1(net5710),
    .S(_03194_),
    .X(_00943_));
 sg13g2_mux2_1 _19773_ (.A0(net3341),
    .A1(net5678),
    .S(_03194_),
    .X(_00944_));
 sg13g2_mux2_1 _19774_ (.A0(net3618),
    .A1(net5650),
    .S(_03194_),
    .X(_00945_));
 sg13g2_mux2_1 _19775_ (.A0(net3860),
    .A1(net5623),
    .S(_03194_),
    .X(_00946_));
 sg13g2_nand2_2 _19776_ (.Y(_03195_),
    .A(net5418),
    .B(_03076_));
 sg13g2_mux2_1 _19777_ (.A0(net5772),
    .A1(net6805),
    .S(_03195_),
    .X(_00947_));
 sg13g2_mux2_1 _19778_ (.A0(net5746),
    .A1(net6307),
    .S(_03195_),
    .X(_00948_));
 sg13g2_mux2_1 _19779_ (.A0(net5715),
    .A1(net6116),
    .S(_03195_),
    .X(_00949_));
 sg13g2_mux2_1 _19780_ (.A0(net5684),
    .A1(net6977),
    .S(_03195_),
    .X(_00950_));
 sg13g2_mux2_1 _19781_ (.A0(net5656),
    .A1(net6656),
    .S(_03195_),
    .X(_00951_));
 sg13g2_mux2_1 _19782_ (.A0(net5627),
    .A1(net6869),
    .S(_03195_),
    .X(_00952_));
 sg13g2_mux2_1 _19783_ (.A0(net5600),
    .A1(net6191),
    .S(_03195_),
    .X(_00953_));
 sg13g2_nor2_2 _19784_ (.A(net5467),
    .B(net5413),
    .Y(_03196_));
 sg13g2_mux2_1 _19785_ (.A0(net3316),
    .A1(net5794),
    .S(_03196_),
    .X(_00954_));
 sg13g2_mux2_1 _19786_ (.A0(net3287),
    .A1(net5768),
    .S(_03196_),
    .X(_00955_));
 sg13g2_mux2_1 _19787_ (.A0(net3836),
    .A1(net5738),
    .S(_03196_),
    .X(_00956_));
 sg13g2_mux2_1 _19788_ (.A0(net3527),
    .A1(net5710),
    .S(_03196_),
    .X(_00957_));
 sg13g2_mux2_1 _19789_ (.A0(net3395),
    .A1(net5678),
    .S(_03196_),
    .X(_00958_));
 sg13g2_mux2_1 _19790_ (.A0(net3789),
    .A1(net5650),
    .S(_03196_),
    .X(_00959_));
 sg13g2_mux2_1 _19791_ (.A0(net3686),
    .A1(net5623),
    .S(_03196_),
    .X(_00960_));
 sg13g2_nand2_2 _19792_ (.Y(_03197_),
    .A(net5468),
    .B(_03104_));
 sg13g2_mux2_1 _19793_ (.A0(net5794),
    .A1(net6802),
    .S(_03197_),
    .X(_00961_));
 sg13g2_mux2_1 _19794_ (.A0(net5768),
    .A1(net6053),
    .S(_03197_),
    .X(_00962_));
 sg13g2_mux2_1 _19795_ (.A0(net5738),
    .A1(net6483),
    .S(_03197_),
    .X(_00963_));
 sg13g2_mux2_1 _19796_ (.A0(net5710),
    .A1(net6177),
    .S(_03197_),
    .X(_00964_));
 sg13g2_mux2_1 _19797_ (.A0(net5678),
    .A1(net6730),
    .S(_03197_),
    .X(_00965_));
 sg13g2_mux2_1 _19798_ (.A0(net5650),
    .A1(net6234),
    .S(_03197_),
    .X(_00966_));
 sg13g2_mux2_1 _19799_ (.A0(net5623),
    .A1(net6642),
    .S(_03197_),
    .X(_00967_));
 sg13g2_nand2_2 _19800_ (.Y(_03198_),
    .A(net5417),
    .B(_03118_));
 sg13g2_mux2_1 _19801_ (.A0(net5772),
    .A1(net6080),
    .S(_03198_),
    .X(_00968_));
 sg13g2_mux2_1 _19802_ (.A0(net5743),
    .A1(net6801),
    .S(_03198_),
    .X(_00969_));
 sg13g2_mux2_1 _19803_ (.A0(net5715),
    .A1(net6366),
    .S(_03198_),
    .X(_00970_));
 sg13g2_mux2_1 _19804_ (.A0(net5685),
    .A1(net6907),
    .S(_03198_),
    .X(_00971_));
 sg13g2_mux2_1 _19805_ (.A0(net5656),
    .A1(net6826),
    .S(_03198_),
    .X(_00972_));
 sg13g2_mux2_1 _19806_ (.A0(net5627),
    .A1(net6774),
    .S(_03198_),
    .X(_00973_));
 sg13g2_mux2_1 _19807_ (.A0(net5600),
    .A1(net6236),
    .S(_03198_),
    .X(_00974_));
 sg13g2_nor2_2 _19808_ (.A(_10479_),
    .B(_03105_),
    .Y(_03199_));
 sg13g2_mux2_1 _19809_ (.A0(net4032),
    .A1(net5786),
    .S(_03199_),
    .X(_00975_));
 sg13g2_mux2_1 _19810_ (.A0(net3394),
    .A1(net5762),
    .S(_03199_),
    .X(_00976_));
 sg13g2_mux2_1 _19811_ (.A0(net3562),
    .A1(net5733),
    .S(_03199_),
    .X(_00977_));
 sg13g2_mux2_1 _19812_ (.A0(net3198),
    .A1(net5705),
    .S(_03199_),
    .X(_00978_));
 sg13g2_mux2_1 _19813_ (.A0(net3463),
    .A1(net5676),
    .S(_03199_),
    .X(_00979_));
 sg13g2_mux2_1 _19814_ (.A0(net3910),
    .A1(net5644),
    .S(_03199_),
    .X(_00980_));
 sg13g2_mux2_1 _19815_ (.A0(net3443),
    .A1(net5617),
    .S(_03199_),
    .X(_00981_));
 sg13g2_nor2_2 _19816_ (.A(_10382_),
    .B(net5413),
    .Y(_03200_));
 sg13g2_mux2_1 _19817_ (.A0(net3518),
    .A1(net5787),
    .S(_03200_),
    .X(_00982_));
 sg13g2_mux2_1 _19818_ (.A0(net3121),
    .A1(net5762),
    .S(_03200_),
    .X(_00983_));
 sg13g2_mux2_1 _19819_ (.A0(net3459),
    .A1(net5731),
    .S(_03200_),
    .X(_00984_));
 sg13g2_mux2_1 _19820_ (.A0(net3674),
    .A1(net5704),
    .S(_03200_),
    .X(_00985_));
 sg13g2_mux2_1 _19821_ (.A0(net3375),
    .A1(net5676),
    .S(_03200_),
    .X(_00986_));
 sg13g2_mux2_1 _19822_ (.A0(net3196),
    .A1(net5645),
    .S(_03200_),
    .X(_00987_));
 sg13g2_mux2_1 _19823_ (.A0(net3590),
    .A1(net5617),
    .S(_03200_),
    .X(_00988_));
 sg13g2_nand2_2 _19824_ (.Y(_03201_),
    .A(_10372_),
    .B(net5417));
 sg13g2_mux2_1 _19825_ (.A0(net5772),
    .A1(net6042),
    .S(_03201_),
    .X(_00989_));
 sg13g2_mux2_1 _19826_ (.A0(net5746),
    .A1(net6570),
    .S(_03201_),
    .X(_00990_));
 sg13g2_mux2_1 _19827_ (.A0(net5715),
    .A1(net6373),
    .S(_03201_),
    .X(_00991_));
 sg13g2_mux2_1 _19828_ (.A0(net5685),
    .A1(net6041),
    .S(_03201_),
    .X(_00992_));
 sg13g2_mux2_1 _19829_ (.A0(net5656),
    .A1(net6047),
    .S(_03201_),
    .X(_00993_));
 sg13g2_mux2_1 _19830_ (.A0(net5627),
    .A1(net4406),
    .S(_03201_),
    .X(_00994_));
 sg13g2_mux2_1 _19831_ (.A0(net5598),
    .A1(net6412),
    .S(_03201_),
    .X(_00995_));
 sg13g2_nand2_2 _19832_ (.Y(_03202_),
    .A(net5469),
    .B(net5412));
 sg13g2_mux2_1 _19833_ (.A0(net5782),
    .A1(net6352),
    .S(_03202_),
    .X(_00996_));
 sg13g2_mux2_1 _19834_ (.A0(net5753),
    .A1(net6328),
    .S(_03202_),
    .X(_00997_));
 sg13g2_mux2_1 _19835_ (.A0(net5724),
    .A1(net4339),
    .S(_03202_),
    .X(_00998_));
 sg13g2_mux2_1 _19836_ (.A0(net5695),
    .A1(net6684),
    .S(_03202_),
    .X(_00999_));
 sg13g2_mux2_1 _19837_ (.A0(net5667),
    .A1(net6303),
    .S(_03202_),
    .X(_01000_));
 sg13g2_mux2_1 _19838_ (.A0(net5638),
    .A1(net4520),
    .S(_03202_),
    .X(_01001_));
 sg13g2_mux2_1 _19839_ (.A0(net5607),
    .A1(net6200),
    .S(_03202_),
    .X(_01002_));
 sg13g2_nand2_2 _19840_ (.Y(_03203_),
    .A(_03104_),
    .B(net5412));
 sg13g2_mux2_1 _19841_ (.A0(net5787),
    .A1(net6779),
    .S(_03203_),
    .X(_01003_));
 sg13g2_mux2_1 _19842_ (.A0(net5762),
    .A1(net6290),
    .S(_03203_),
    .X(_01004_));
 sg13g2_mux2_1 _19843_ (.A0(net5731),
    .A1(net6594),
    .S(_03203_),
    .X(_01005_));
 sg13g2_mux2_1 _19844_ (.A0(net5704),
    .A1(net6208),
    .S(_03203_),
    .X(_01006_));
 sg13g2_mux2_1 _19845_ (.A0(net5676),
    .A1(net6261),
    .S(_03203_),
    .X(_01007_));
 sg13g2_mux2_1 _19846_ (.A0(net5644),
    .A1(net6902),
    .S(_03203_),
    .X(_01008_));
 sg13g2_mux2_1 _19847_ (.A0(net5617),
    .A1(net6271),
    .S(_03203_),
    .X(_01009_));
 sg13g2_nand2_2 _19848_ (.Y(_03204_),
    .A(net5417),
    .B(net5411));
 sg13g2_mux2_1 _19849_ (.A0(net5772),
    .A1(net6134),
    .S(_03204_),
    .X(_01010_));
 sg13g2_mux2_1 _19850_ (.A0(net5746),
    .A1(net6099),
    .S(_03204_),
    .X(_01011_));
 sg13g2_mux2_1 _19851_ (.A0(net5715),
    .A1(net6338),
    .S(_03204_),
    .X(_01012_));
 sg13g2_mux2_1 _19852_ (.A0(net5685),
    .A1(net6387),
    .S(_03204_),
    .X(_01013_));
 sg13g2_mux2_1 _19853_ (.A0(net5657),
    .A1(net6758),
    .S(_03204_),
    .X(_01014_));
 sg13g2_mux2_1 _19854_ (.A0(net5627),
    .A1(net6411),
    .S(_03204_),
    .X(_01015_));
 sg13g2_mux2_1 _19855_ (.A0(net5600),
    .A1(net6461),
    .S(_03204_),
    .X(_01016_));
 sg13g2_nor2_2 _19856_ (.A(_03077_),
    .B(net5413),
    .Y(_03205_));
 sg13g2_mux2_1 _19857_ (.A0(net3792),
    .A1(net5794),
    .S(_03205_),
    .X(_01017_));
 sg13g2_mux2_1 _19858_ (.A0(net3675),
    .A1(net5766),
    .S(_03205_),
    .X(_01018_));
 sg13g2_mux2_1 _19859_ (.A0(net3213),
    .A1(net5735),
    .S(_03205_),
    .X(_01019_));
 sg13g2_mux2_1 _19860_ (.A0(net3498),
    .A1(net5710),
    .S(_03205_),
    .X(_01020_));
 sg13g2_mux2_1 _19861_ (.A0(net3542),
    .A1(net5676),
    .S(_03205_),
    .X(_01021_));
 sg13g2_mux2_1 _19862_ (.A0(net3503),
    .A1(net5651),
    .S(_03205_),
    .X(_01022_));
 sg13g2_mux2_1 _19863_ (.A0(net3457),
    .A1(net5622),
    .S(_03205_),
    .X(_01023_));
 sg13g2_nor2_2 _19864_ (.A(net5413),
    .B(_03119_),
    .Y(_03206_));
 sg13g2_mux2_1 _19865_ (.A0(net3360),
    .A1(net5796),
    .S(_03206_),
    .X(_01024_));
 sg13g2_mux2_1 _19866_ (.A0(net3225),
    .A1(net5766),
    .S(_03206_),
    .X(_01025_));
 sg13g2_mux2_1 _19867_ (.A0(net3552),
    .A1(net5735),
    .S(_03206_),
    .X(_01026_));
 sg13g2_mux2_1 _19868_ (.A0(net3587),
    .A1(net5706),
    .S(_03206_),
    .X(_01027_));
 sg13g2_mux2_1 _19869_ (.A0(net3520),
    .A1(net5676),
    .S(_03206_),
    .X(_01028_));
 sg13g2_mux2_1 _19870_ (.A0(net3209),
    .A1(net5651),
    .S(_03206_),
    .X(_01029_));
 sg13g2_mux2_1 _19871_ (.A0(net3444),
    .A1(net5622),
    .S(_03206_),
    .X(_01030_));
 sg13g2_nand2_2 _19872_ (.Y(_03207_),
    .A(net5418),
    .B(_03100_));
 sg13g2_mux2_1 _19873_ (.A0(net5775),
    .A1(net6087),
    .S(_03207_),
    .X(_01031_));
 sg13g2_mux2_1 _19874_ (.A0(net5745),
    .A1(net6286),
    .S(_03207_),
    .X(_01032_));
 sg13g2_mux2_1 _19875_ (.A0(net5715),
    .A1(net6326),
    .S(_03207_),
    .X(_01033_));
 sg13g2_mux2_1 _19876_ (.A0(net5688),
    .A1(net6646),
    .S(_03207_),
    .X(_01034_));
 sg13g2_mux2_1 _19877_ (.A0(net5659),
    .A1(net6797),
    .S(_03207_),
    .X(_01035_));
 sg13g2_mux2_1 _19878_ (.A0(net5631),
    .A1(net4528),
    .S(_03207_),
    .X(_01036_));
 sg13g2_mux2_1 _19879_ (.A0(net5600),
    .A1(net6871),
    .S(_03207_),
    .X(_01037_));
 sg13g2_nor2_2 _19880_ (.A(_10373_),
    .B(net5413),
    .Y(_03208_));
 sg13g2_mux2_1 _19881_ (.A0(net3651),
    .A1(net5796),
    .S(_03208_),
    .X(_01038_));
 sg13g2_mux2_1 _19882_ (.A0(net3896),
    .A1(net5759),
    .S(_03208_),
    .X(_01039_));
 sg13g2_mux2_1 _19883_ (.A0(net3181),
    .A1(net5735),
    .S(_03208_),
    .X(_01040_));
 sg13g2_mux2_1 _19884_ (.A0(net3862),
    .A1(net5706),
    .S(_03208_),
    .X(_01041_));
 sg13g2_mux2_1 _19885_ (.A0(net3445),
    .A1(net5669),
    .S(_03208_),
    .X(_01042_));
 sg13g2_mux2_1 _19886_ (.A0(net3358),
    .A1(net5651),
    .S(_03208_),
    .X(_01043_));
 sg13g2_mux2_1 _19887_ (.A0(net3791),
    .A1(net5622),
    .S(_03208_),
    .X(_01044_));
 sg13g2_nand2_2 _19888_ (.Y(_03209_),
    .A(_03104_),
    .B(net5411));
 sg13g2_mux2_1 _19889_ (.A0(net5796),
    .A1(net6900),
    .S(_03209_),
    .X(_01045_));
 sg13g2_mux2_1 _19890_ (.A0(net5759),
    .A1(net6327),
    .S(_03209_),
    .X(_01046_));
 sg13g2_mux2_1 _19891_ (.A0(net5735),
    .A1(net4337),
    .S(_03209_),
    .X(_01047_));
 sg13g2_mux2_1 _19892_ (.A0(net5706),
    .A1(net6770),
    .S(_03209_),
    .X(_01048_));
 sg13g2_mux2_1 _19893_ (.A0(net5669),
    .A1(net6653),
    .S(_03209_),
    .X(_01049_));
 sg13g2_mux2_1 _19894_ (.A0(net5651),
    .A1(net6255),
    .S(_03209_),
    .X(_01050_));
 sg13g2_mux2_1 _19895_ (.A0(net5616),
    .A1(net6315),
    .S(_03209_),
    .X(_01051_));
 sg13g2_nand2_2 _19896_ (.Y(_03210_),
    .A(net5419),
    .B(net5418));
 sg13g2_mux2_1 _19897_ (.A0(net5775),
    .A1(net6706),
    .S(_03210_),
    .X(_01052_));
 sg13g2_mux2_1 _19898_ (.A0(net5745),
    .A1(net6662),
    .S(_03210_),
    .X(_01053_));
 sg13g2_mux2_1 _19899_ (.A0(net5715),
    .A1(net6238),
    .S(_03210_),
    .X(_01054_));
 sg13g2_mux2_1 _19900_ (.A0(net5688),
    .A1(net3961),
    .S(_03210_),
    .X(_01055_));
 sg13g2_mux2_1 _19901_ (.A0(net5660),
    .A1(net6781),
    .S(_03210_),
    .X(_01056_));
 sg13g2_mux2_1 _19902_ (.A0(net5631),
    .A1(net6744),
    .S(_03210_),
    .X(_01057_));
 sg13g2_mux2_1 _19903_ (.A0(net5600),
    .A1(net4382),
    .S(_03210_),
    .X(_01058_));
 sg13g2_nor2_2 _19904_ (.A(_03101_),
    .B(net5413),
    .Y(_03211_));
 sg13g2_mux2_1 _19905_ (.A0(net3718),
    .A1(net5786),
    .S(_03211_),
    .X(_01059_));
 sg13g2_mux2_1 _19906_ (.A0(net3769),
    .A1(net5764),
    .S(_03211_),
    .X(_01060_));
 sg13g2_mux2_1 _19907_ (.A0(net3266),
    .A1(net5733),
    .S(_03211_),
    .X(_01061_));
 sg13g2_mux2_1 _19908_ (.A0(net3413),
    .A1(net5704),
    .S(_03211_),
    .X(_01062_));
 sg13g2_mux2_1 _19909_ (.A0(net3519),
    .A1(net5678),
    .S(_03211_),
    .X(_01063_));
 sg13g2_mux2_1 _19910_ (.A0(net3784),
    .A1(net5644),
    .S(_03211_),
    .X(_01064_));
 sg13g2_mux2_1 _19911_ (.A0(net3956),
    .A1(net5619),
    .S(_03211_),
    .X(_01065_));
 sg13g2_nand2_2 _19912_ (.Y(_03212_),
    .A(net5419),
    .B(_03104_));
 sg13g2_mux2_1 _19913_ (.A0(net5786),
    .A1(net4505),
    .S(_03212_),
    .X(_01066_));
 sg13g2_mux2_1 _19914_ (.A0(net5764),
    .A1(net6448),
    .S(_03212_),
    .X(_01067_));
 sg13g2_mux2_1 _19915_ (.A0(net5733),
    .A1(net6567),
    .S(_03212_),
    .X(_01068_));
 sg13g2_mux2_1 _19916_ (.A0(net5704),
    .A1(net6137),
    .S(_03212_),
    .X(_01069_));
 sg13g2_mux2_1 _19917_ (.A0(net5678),
    .A1(net6476),
    .S(_03212_),
    .X(_01070_));
 sg13g2_mux2_1 _19918_ (.A0(net5644),
    .A1(net6249),
    .S(_03212_),
    .X(_01071_));
 sg13g2_mux2_1 _19919_ (.A0(net5619),
    .A1(net6898),
    .S(_03212_),
    .X(_01072_));
 sg13g2_nand2_2 _19920_ (.Y(_03213_),
    .A(net5470),
    .B(net5468));
 sg13g2_mux2_1 _19921_ (.A0(net5783),
    .A1(net6186),
    .S(_03213_),
    .X(_01073_));
 sg13g2_mux2_1 _19922_ (.A0(net5754),
    .A1(net6161),
    .S(_03213_),
    .X(_01074_));
 sg13g2_mux2_1 _19923_ (.A0(net5725),
    .A1(net6759),
    .S(_03213_),
    .X(_01075_));
 sg13g2_mux2_1 _19924_ (.A0(net5696),
    .A1(net6291),
    .S(_03213_),
    .X(_01076_));
 sg13g2_mux2_1 _19925_ (.A0(net5667),
    .A1(net4344),
    .S(_03213_),
    .X(_01077_));
 sg13g2_mux2_1 _19926_ (.A0(net5640),
    .A1(net6159),
    .S(_03213_),
    .X(_01078_));
 sg13g2_mux2_1 _19927_ (.A0(net5610),
    .A1(net6068),
    .S(_03213_),
    .X(_01079_));
 sg13g2_nand2_2 _19928_ (.Y(_03214_),
    .A(net5469),
    .B(_03076_));
 sg13g2_mux2_1 _19929_ (.A0(net5785),
    .A1(net6497),
    .S(_03214_),
    .X(_01080_));
 sg13g2_mux2_1 _19930_ (.A0(net5753),
    .A1(net6645),
    .S(_03214_),
    .X(_01081_));
 sg13g2_mux2_1 _19931_ (.A0(net5724),
    .A1(net6760),
    .S(_03214_),
    .X(_01082_));
 sg13g2_mux2_1 _19932_ (.A0(net5695),
    .A1(net6533),
    .S(_03214_),
    .X(_01083_));
 sg13g2_mux2_1 _19933_ (.A0(net5669),
    .A1(net4303),
    .S(_03214_),
    .X(_01084_));
 sg13g2_mux2_1 _19934_ (.A0(net5639),
    .A1(net6824),
    .S(_03214_),
    .X(_01085_));
 sg13g2_mux2_1 _19935_ (.A0(net5609),
    .A1(net6927),
    .S(_03214_),
    .X(_01086_));
 sg13g2_nor2_2 _19936_ (.A(_10377_),
    .B(net5471),
    .Y(_03215_));
 sg13g2_mux2_1 _19937_ (.A0(net3475),
    .A1(net5771),
    .S(_03215_),
    .X(_01087_));
 sg13g2_mux2_1 _19938_ (.A0(net3362),
    .A1(net5742),
    .S(_03215_),
    .X(_01088_));
 sg13g2_mux2_1 _19939_ (.A0(net3482),
    .A1(net5713),
    .S(_03215_),
    .X(_01089_));
 sg13g2_mux2_1 _19940_ (.A0(net3148),
    .A1(net5684),
    .S(_03215_),
    .X(_01090_));
 sg13g2_mux2_1 _19941_ (.A0(net3469),
    .A1(net5655),
    .S(_03215_),
    .X(_01091_));
 sg13g2_mux2_1 _19942_ (.A0(net3524),
    .A1(net5626),
    .S(_03215_),
    .X(_01092_));
 sg13g2_mux2_1 _19943_ (.A0(net3954),
    .A1(net5597),
    .S(_03215_),
    .X(_01093_));
 sg13g2_nand2_2 _19944_ (.Y(_03216_),
    .A(net5431),
    .B(_10478_));
 sg13g2_mux2_1 _19945_ (.A0(net5774),
    .A1(net6520),
    .S(_03216_),
    .X(_01094_));
 sg13g2_mux2_1 _19946_ (.A0(net5745),
    .A1(net6627),
    .S(_03216_),
    .X(_01095_));
 sg13g2_mux2_1 _19947_ (.A0(net5716),
    .A1(net6397),
    .S(_03216_),
    .X(_01096_));
 sg13g2_mux2_1 _19948_ (.A0(net5690),
    .A1(net6650),
    .S(_03216_),
    .X(_01097_));
 sg13g2_mux2_1 _19949_ (.A0(net5661),
    .A1(net6833),
    .S(_03216_),
    .X(_01098_));
 sg13g2_mux2_1 _19950_ (.A0(net5628),
    .A1(net6088),
    .S(_03216_),
    .X(_01099_));
 sg13g2_mux2_1 _19951_ (.A0(net5600),
    .A1(net6754),
    .S(_03216_),
    .X(_01100_));
 sg13g2_nor2_2 _19952_ (.A(_10377_),
    .B(net5467),
    .Y(_03217_));
 sg13g2_mux2_1 _19953_ (.A0(net3803),
    .A1(net5771),
    .S(_03217_),
    .X(_01101_));
 sg13g2_mux2_1 _19954_ (.A0(net3438),
    .A1(net5742),
    .S(_03217_),
    .X(_01102_));
 sg13g2_mux2_1 _19955_ (.A0(net3306),
    .A1(net5713),
    .S(_03217_),
    .X(_01103_));
 sg13g2_mux2_1 _19956_ (.A0(net3537),
    .A1(net5684),
    .S(_03217_),
    .X(_01104_));
 sg13g2_mux2_1 _19957_ (.A0(net3949),
    .A1(net5655),
    .S(_03217_),
    .X(_01105_));
 sg13g2_mux2_1 _19958_ (.A0(net3396),
    .A1(net5626),
    .S(_03217_),
    .X(_01106_));
 sg13g2_mux2_1 _19959_ (.A0(net3274),
    .A1(net5597),
    .S(_03217_),
    .X(_01107_));
 sg13g2_nand2_2 _19960_ (.Y(_03218_),
    .A(net5432),
    .B(_03118_));
 sg13g2_mux2_1 _19961_ (.A0(net5773),
    .A1(net4490),
    .S(_03218_),
    .X(_01108_));
 sg13g2_mux2_1 _19962_ (.A0(net5747),
    .A1(net4360),
    .S(_03218_),
    .X(_01109_));
 sg13g2_mux2_1 _19963_ (.A0(net5717),
    .A1(net6258),
    .S(_03218_),
    .X(_01110_));
 sg13g2_mux2_1 _19964_ (.A0(net5689),
    .A1(net6595),
    .S(_03218_),
    .X(_01111_));
 sg13g2_mux2_1 _19965_ (.A0(net5658),
    .A1(net6376),
    .S(_03218_),
    .X(_01112_));
 sg13g2_mux2_1 _19966_ (.A0(net5628),
    .A1(net6543),
    .S(_03218_),
    .X(_01113_));
 sg13g2_mux2_1 _19967_ (.A0(net5601),
    .A1(net4172),
    .S(_03218_),
    .X(_01114_));
 sg13g2_nand2_2 _19968_ (.Y(_03219_),
    .A(net5431),
    .B(_02995_));
 sg13g2_mux2_1 _19969_ (.A0(net5773),
    .A1(net6589),
    .S(_03219_),
    .X(_01115_));
 sg13g2_mux2_1 _19970_ (.A0(net5745),
    .A1(net6511),
    .S(_03219_),
    .X(_01116_));
 sg13g2_mux2_1 _19971_ (.A0(net5716),
    .A1(net6199),
    .S(_03219_),
    .X(_01117_));
 sg13g2_mux2_1 _19972_ (.A0(net5690),
    .A1(net6968),
    .S(_03219_),
    .X(_01118_));
 sg13g2_mux2_1 _19973_ (.A0(net5661),
    .A1(net6406),
    .S(_03219_),
    .X(_01119_));
 sg13g2_mux2_1 _19974_ (.A0(net5629),
    .A1(net6481),
    .S(_03219_),
    .X(_01120_));
 sg13g2_mux2_1 _19975_ (.A0(net5597),
    .A1(net6561),
    .S(_03219_),
    .X(_01121_));
 sg13g2_nand2_1 _19976_ (.Y(_03220_),
    .A(net3122),
    .B(net5999));
 sg13g2_a21oi_1 _19977_ (.A1(_10444_),
    .A2(_03220_),
    .Y(_01122_),
    .B1(net5537));
 sg13g2_nor2_1 _19978_ (.A(net7027),
    .B(rom_data_pending),
    .Y(_03221_));
 sg13g2_nor3_1 _19979_ (.A(_08106_),
    .B(net5315),
    .C(_10424_),
    .Y(_03222_));
 sg13g2_a21oi_1 _19980_ (.A1(_10443_),
    .A2(_03222_),
    .Y(_01123_),
    .B1(net7028));
 sg13g2_and2_2 _19981_ (.A(\hvsync_gen.hpos[0] ),
    .B(net7179),
    .X(_03223_));
 sg13g2_nand3_1 _19982_ (.B(net5925),
    .C(_03223_),
    .A(net5871),
    .Y(_03224_));
 sg13g2_or2_2 _19983_ (.X(_03225_),
    .B(net5845),
    .A(net5843));
 sg13g2_or2_2 _19984_ (.X(_03226_),
    .B(net5509),
    .A(net5552));
 sg13g2_nor2b_1 _19985_ (.A(net5849),
    .B_N(net5850),
    .Y(_03227_));
 sg13g2_nand2b_1 _19986_ (.Y(_03228_),
    .B(net5850),
    .A_N(net5849));
 sg13g2_or4_2 _19987_ (.A(_08120_),
    .B(_03224_),
    .C(_03226_),
    .D(net5498),
    .X(_03229_));
 sg13g2_and2_2 _19988_ (.A(net6037),
    .B(_03229_),
    .X(_03230_));
 sg13g2_nand2_2 _19989_ (.Y(_03231_),
    .A(net6037),
    .B(_03229_));
 sg13g2_and2_1 _19990_ (.A(net2891),
    .B(_03230_),
    .X(_01124_));
 sg13g2_nor2_2 _19991_ (.A(\hvsync_gen.hpos[0] ),
    .B(net7179),
    .Y(_03232_));
 sg13g2_nor3_1 _19992_ (.A(net5991),
    .B(_03223_),
    .C(_03232_),
    .Y(_01125_));
 sg13g2_nor2_1 _19993_ (.A(_08106_),
    .B(spi_data_ready_last),
    .Y(_03233_));
 sg13g2_nand2b_1 _19994_ (.Y(_03234_),
    .B(\flash_rom.data_ready ),
    .A_N(spi_data_ready_last));
 sg13g2_nand3_1 _19995_ (.B(net4568),
    .C(net5496),
    .A(net5034),
    .Y(_03235_));
 sg13g2_nor3_1 _19996_ (.A(net5978),
    .B(net4568),
    .C(net5464),
    .Y(_03236_));
 sg13g2_nand3b_1 _19997_ (.B(net5496),
    .C(net5999),
    .Y(_03237_),
    .A_N(net4567));
 sg13g2_nand2_1 _19998_ (.Y(_03238_),
    .A(\rom_next_addr_in_queue[0] ),
    .B(net5465));
 sg13g2_nand3_1 _19999_ (.B(net4557),
    .C(_03238_),
    .A(_03235_),
    .Y(_03239_));
 sg13g2_o21ai_1 _20000_ (.B1(_03239_),
    .Y(_03240_),
    .A1(net7213),
    .A2(_03237_));
 sg13g2_inv_1 _20001_ (.Y(_01126_),
    .A(net7214));
 sg13g2_a21oi_1 _20002_ (.A1(net5035),
    .A2(net4567),
    .Y(_03241_),
    .B1(net5465));
 sg13g2_a21oi_1 _20003_ (.A1(_08089_),
    .A2(net5465),
    .Y(_03242_),
    .B1(_03241_));
 sg13g2_a21o_1 _20004_ (.A2(net4561),
    .A1(net6983),
    .B1(_03242_),
    .X(_01127_));
 sg13g2_nand3_1 _20005_ (.B(net4567),
    .C(net5496),
    .A(net5029),
    .Y(_03243_));
 sg13g2_a21oi_1 _20006_ (.A1(\rom_next_addr_in_queue[2] ),
    .A2(net5464),
    .Y(_03244_),
    .B1(net4561));
 sg13g2_a22oi_1 _20007_ (.Y(_01128_),
    .B1(_03243_),
    .B2(_03244_),
    .A2(net4562),
    .A1(_08078_));
 sg13g2_and3_1 _20008_ (.X(_03245_),
    .A(net5036),
    .B(net4568),
    .C(net5496));
 sg13g2_a21oi_1 _20009_ (.A1(\rom_next_addr_in_queue[3] ),
    .A2(net5465),
    .Y(_03246_),
    .B1(_03245_));
 sg13g2_nor2_1 _20010_ (.A(net6618),
    .B(net4557),
    .Y(_03247_));
 sg13g2_a21oi_1 _20011_ (.A1(net4557),
    .A2(_03246_),
    .Y(_01129_),
    .B1(_03247_));
 sg13g2_nor2_1 _20012_ (.A(_10454_),
    .B(net5464),
    .Y(_03248_));
 sg13g2_a21oi_1 _20013_ (.A1(\rom_next_addr_in_queue[4] ),
    .A2(net5464),
    .Y(_03249_),
    .B1(_03248_));
 sg13g2_nor2_1 _20014_ (.A(net3974),
    .B(net4556),
    .Y(_03250_));
 sg13g2_a21oi_1 _20015_ (.A1(net4556),
    .A2(_03249_),
    .Y(_01130_),
    .B1(_03250_));
 sg13g2_nor2_1 _20016_ (.A(_10457_),
    .B(net5464),
    .Y(_03251_));
 sg13g2_a21oi_1 _20017_ (.A1(\rom_next_addr_in_queue[5] ),
    .A2(net5464),
    .Y(_03252_),
    .B1(_03251_));
 sg13g2_nor2_1 _20018_ (.A(net3977),
    .B(net4556),
    .Y(_03253_));
 sg13g2_a21oi_1 _20019_ (.A1(net4556),
    .A2(_03252_),
    .Y(_01131_),
    .B1(_03253_));
 sg13g2_nand3_1 _20020_ (.B(net4567),
    .C(net5495),
    .A(net5022),
    .Y(_03254_));
 sg13g2_a21oi_1 _20021_ (.A1(\rom_next_addr_in_queue[6] ),
    .A2(net5466),
    .Y(_03255_),
    .B1(net4563));
 sg13g2_a22oi_1 _20022_ (.Y(_01132_),
    .B1(_03254_),
    .B2(_03255_),
    .A2(net4563),
    .A1(_08079_));
 sg13g2_nand3_1 _20023_ (.B(net4567),
    .C(net5495),
    .A(_10417_),
    .Y(_03256_));
 sg13g2_a21oi_1 _20024_ (.A1(\rom_next_addr_in_queue[7] ),
    .A2(net5463),
    .Y(_03257_),
    .B1(net4559));
 sg13g2_a22oi_1 _20025_ (.Y(_01133_),
    .B1(_03256_),
    .B2(_03257_),
    .A2(net4559),
    .A1(_08082_));
 sg13g2_nand3_1 _20026_ (.B(net4567),
    .C(net5495),
    .A(_10397_),
    .Y(_03258_));
 sg13g2_a21oi_1 _20027_ (.A1(\rom_next_addr_in_queue[8] ),
    .A2(net5463),
    .Y(_03259_),
    .B1(net4558));
 sg13g2_a22oi_1 _20028_ (.Y(_01134_),
    .B1(_03258_),
    .B2(_03259_),
    .A2(net4559),
    .A1(_08083_));
 sg13g2_nand3_1 _20029_ (.B(net4567),
    .C(net5495),
    .A(_10403_),
    .Y(_03260_));
 sg13g2_a21oi_1 _20030_ (.A1(\rom_next_addr_in_queue[9] ),
    .A2(net5463),
    .Y(_03261_),
    .B1(net4560));
 sg13g2_a22oi_1 _20031_ (.Y(_01135_),
    .B1(_03260_),
    .B2(_03261_),
    .A2(net4560),
    .A1(_08085_));
 sg13g2_nand3_1 _20032_ (.B(net4564),
    .C(net5495),
    .A(_10390_),
    .Y(_03262_));
 sg13g2_a21oi_1 _20033_ (.A1(\rom_next_addr_in_queue[10] ),
    .A2(net5463),
    .Y(_03263_),
    .B1(net4558));
 sg13g2_a22oi_1 _20034_ (.Y(_01136_),
    .B1(_03262_),
    .B2(_03263_),
    .A2(net4558),
    .A1(_08086_));
 sg13g2_nand3_1 _20035_ (.B(net4567),
    .C(net5495),
    .A(_10412_),
    .Y(_03264_));
 sg13g2_a21oi_1 _20036_ (.A1(\rom_next_addr_in_queue[11] ),
    .A2(net5463),
    .Y(_03265_),
    .B1(net4558));
 sg13g2_a22oi_1 _20037_ (.Y(_01137_),
    .B1(_03264_),
    .B2(_03265_),
    .A2(net4559),
    .A1(_08087_));
 sg13g2_a21oi_1 _20038_ (.A1(net7018),
    .A2(net5465),
    .Y(_03266_),
    .B1(net4561));
 sg13g2_a22oi_1 _20039_ (.Y(_01138_),
    .B1(_03266_),
    .B2(_03235_),
    .A2(net4561),
    .A1(_08088_));
 sg13g2_o21ai_1 _20040_ (.B1(net4557),
    .Y(_03267_),
    .A1(net7209),
    .A2(_03238_));
 sg13g2_a21oi_1 _20041_ (.A1(_03238_),
    .A2(_03242_),
    .Y(_03268_),
    .B1(net7210));
 sg13g2_a21oi_1 _20042_ (.A1(_08089_),
    .A2(net4561),
    .Y(_01139_),
    .B1(net7211));
 sg13g2_nor3_1 _20043_ (.A(_08088_),
    .B(_08089_),
    .C(_08090_),
    .Y(_03269_));
 sg13g2_a21oi_1 _20044_ (.A1(\rom_next_addr_in_queue[0] ),
    .A2(net7209),
    .Y(_03270_),
    .B1(net7242));
 sg13g2_nor3_1 _20045_ (.A(net5496),
    .B(_03269_),
    .C(_03270_),
    .Y(_03271_));
 sg13g2_nor2_1 _20046_ (.A(net4561),
    .B(_03271_),
    .Y(_03272_));
 sg13g2_a22oi_1 _20047_ (.Y(_01140_),
    .B1(_03243_),
    .B2(_03272_),
    .A2(net4561),
    .A1(_08090_));
 sg13g2_and2_1 _20048_ (.A(\rom_next_addr_in_queue[3] ),
    .B(_03269_),
    .X(_03273_));
 sg13g2_nor2_1 _20049_ (.A(net7136),
    .B(_03269_),
    .Y(_03274_));
 sg13g2_nor3_1 _20050_ (.A(net5496),
    .B(_03273_),
    .C(_03274_),
    .Y(_03275_));
 sg13g2_nor3_1 _20051_ (.A(net4562),
    .B(_03245_),
    .C(_03275_),
    .Y(_03276_));
 sg13g2_a21oi_1 _20052_ (.A1(_08091_),
    .A2(net4562),
    .Y(_01141_),
    .B1(_03276_));
 sg13g2_and2_1 _20053_ (.A(\rom_next_addr_in_queue[4] ),
    .B(_03273_),
    .X(_03277_));
 sg13g2_o21ai_1 _20054_ (.B1(net5464),
    .Y(_03278_),
    .A1(net7105),
    .A2(_03273_));
 sg13g2_o21ai_1 _20055_ (.B1(net4557),
    .Y(_03279_),
    .A1(_03277_),
    .A2(_03278_));
 sg13g2_nor2_1 _20056_ (.A(_03248_),
    .B(_03279_),
    .Y(_03280_));
 sg13g2_a21oi_1 _20057_ (.A1(_08092_),
    .A2(net4561),
    .Y(_01142_),
    .B1(_03280_));
 sg13g2_and2_1 _20058_ (.A(\rom_next_addr_in_queue[5] ),
    .B(_03277_),
    .X(_03281_));
 sg13g2_o21ai_1 _20059_ (.B1(net5464),
    .Y(_03282_),
    .A1(\rom_next_addr_in_queue[5] ),
    .A2(_03277_));
 sg13g2_o21ai_1 _20060_ (.B1(net4557),
    .Y(_03283_),
    .A1(_03281_),
    .A2(_03282_));
 sg13g2_nor2_1 _20061_ (.A(_03251_),
    .B(_03283_),
    .Y(_03284_));
 sg13g2_a21oi_1 _20062_ (.A1(_08093_),
    .A2(net4562),
    .Y(_01143_),
    .B1(_03284_));
 sg13g2_and2_1 _20063_ (.A(\rom_next_addr_in_queue[6] ),
    .B(_03281_),
    .X(_03285_));
 sg13g2_o21ai_1 _20064_ (.B1(net5466),
    .Y(_03286_),
    .A1(\rom_next_addr_in_queue[6] ),
    .A2(_03281_));
 sg13g2_o21ai_1 _20065_ (.B1(_03254_),
    .Y(_03287_),
    .A1(_03285_),
    .A2(_03286_));
 sg13g2_mux2_1 _20066_ (.A0(net7119),
    .A1(_03287_),
    .S(net4557),
    .X(_01144_));
 sg13g2_and2_1 _20067_ (.A(\rom_next_addr_in_queue[7] ),
    .B(_03285_),
    .X(_03288_));
 sg13g2_o21ai_1 _20068_ (.B1(net5463),
    .Y(_03289_),
    .A1(\rom_next_addr_in_queue[7] ),
    .A2(_03285_));
 sg13g2_o21ai_1 _20069_ (.B1(_03256_),
    .Y(_03290_),
    .A1(_03288_),
    .A2(_03289_));
 sg13g2_mux2_1 _20070_ (.A0(net7128),
    .A1(_03290_),
    .S(net4556),
    .X(_01145_));
 sg13g2_and2_1 _20071_ (.A(\rom_next_addr_in_queue[8] ),
    .B(_03288_),
    .X(_03291_));
 sg13g2_o21ai_1 _20072_ (.B1(net5463),
    .Y(_03292_),
    .A1(\rom_next_addr_in_queue[8] ),
    .A2(_03288_));
 sg13g2_o21ai_1 _20073_ (.B1(_03258_),
    .Y(_03293_),
    .A1(_03291_),
    .A2(_03292_));
 sg13g2_mux2_1 _20074_ (.A0(net7151),
    .A1(_03293_),
    .S(net4556),
    .X(_01146_));
 sg13g2_a21oi_1 _20075_ (.A1(\rom_next_addr_in_queue[9] ),
    .A2(_03291_),
    .Y(_03294_),
    .B1(net5495));
 sg13g2_o21ai_1 _20076_ (.B1(_03294_),
    .Y(_03295_),
    .A1(\rom_next_addr_in_queue[9] ),
    .A2(_03291_));
 sg13g2_nand3_1 _20077_ (.B(_03260_),
    .C(_03295_),
    .A(net4556),
    .Y(_03296_));
 sg13g2_o21ai_1 _20078_ (.B1(_03296_),
    .Y(_03297_),
    .A1(net7294),
    .A2(net4556));
 sg13g2_inv_1 _20079_ (.Y(_01147_),
    .A(_03297_));
 sg13g2_nand3_1 _20080_ (.B(net7120),
    .C(_03291_),
    .A(\rom_next_addr_in_queue[9] ),
    .Y(_03298_));
 sg13g2_a21oi_1 _20081_ (.A1(\rom_next_addr_in_queue[9] ),
    .A2(_03291_),
    .Y(_03299_),
    .B1(net7120));
 sg13g2_nor2_1 _20082_ (.A(net5495),
    .B(_03299_),
    .Y(_03300_));
 sg13g2_a21oi_1 _20083_ (.A1(_03298_),
    .A2(_03300_),
    .Y(_03301_),
    .B1(net4558));
 sg13g2_a22oi_1 _20084_ (.Y(_01148_),
    .B1(_03262_),
    .B2(_03301_),
    .A2(net4558),
    .A1(_08094_));
 sg13g2_xnor2_1 _20085_ (.Y(_03302_),
    .A(net7223),
    .B(_03298_));
 sg13g2_a21oi_1 _20086_ (.A1(net5463),
    .A2(_03302_),
    .Y(_03303_),
    .B1(net4558));
 sg13g2_a22oi_1 _20087_ (.Y(_01149_),
    .B1(_03264_),
    .B2(_03303_),
    .A2(net4558),
    .A1(_08095_));
 sg13g2_a21oi_1 _20088_ (.A1(net3379),
    .A2(net5832),
    .Y(_03304_),
    .B1(\audio_pwm_accumulator[0] ));
 sg13g2_nand3_1 _20089_ (.B(net5832),
    .C(\audio_pwm_accumulator[0] ),
    .A(net3379),
    .Y(_03305_));
 sg13g2_nand2b_1 _20090_ (.Y(_03306_),
    .B(_03305_),
    .A_N(_03304_));
 sg13g2_nand2_1 _20091_ (.Y(_03307_),
    .A(net2936),
    .B(net7012));
 sg13g2_o21ai_1 _20092_ (.B1(net6022),
    .Y(_03308_),
    .A1(_03306_),
    .A2(_03307_));
 sg13g2_a21oi_1 _20093_ (.A1(_03306_),
    .A2(_03307_),
    .Y(_01150_),
    .B1(_03308_));
 sg13g2_o21ai_1 _20094_ (.B1(_03305_),
    .Y(_03309_),
    .A1(_03304_),
    .A2(_03307_));
 sg13g2_nand2_1 _20095_ (.Y(_03310_),
    .A(\atari2600.tia.audv0[1] ),
    .B(\atari2600.tia.audio_l ));
 sg13g2_nand3_1 _20096_ (.B(net5833),
    .C(\audio_pwm_accumulator[1] ),
    .A(\atari2600.tia.audv1[1] ),
    .Y(_03311_));
 sg13g2_a21o_1 _20097_ (.A2(net5833),
    .A1(\atari2600.tia.audv1[1] ),
    .B1(\audio_pwm_accumulator[1] ),
    .X(_03312_));
 sg13g2_nand2_1 _20098_ (.Y(_03313_),
    .A(_03311_),
    .B(_03312_));
 sg13g2_xor2_1 _20099_ (.B(_03313_),
    .A(_03310_),
    .X(_03314_));
 sg13g2_or2_1 _20100_ (.X(_03315_),
    .B(_03314_),
    .A(_03309_));
 sg13g2_nand2_1 _20101_ (.Y(_03316_),
    .A(_03309_),
    .B(_03314_));
 sg13g2_and3_1 _20102_ (.X(_01151_),
    .A(net6022),
    .B(_03315_),
    .C(_03316_));
 sg13g2_nand2_1 _20103_ (.Y(_03317_),
    .A(\atari2600.tia.audv0[2] ),
    .B(\atari2600.tia.audio_l ));
 sg13g2_and3_1 _20104_ (.X(_03318_),
    .A(\atari2600.tia.audv1[2] ),
    .B(net5832),
    .C(\audio_pwm_accumulator[2] ));
 sg13g2_nand3_1 _20105_ (.B(net5832),
    .C(\audio_pwm_accumulator[2] ),
    .A(\atari2600.tia.audv1[2] ),
    .Y(_03319_));
 sg13g2_a21oi_1 _20106_ (.A1(\atari2600.tia.audv1[2] ),
    .A2(net5832),
    .Y(_03320_),
    .B1(\audio_pwm_accumulator[2] ));
 sg13g2_nor2_1 _20107_ (.A(_03318_),
    .B(_03320_),
    .Y(_03321_));
 sg13g2_xnor2_1 _20108_ (.Y(_03322_),
    .A(_03317_),
    .B(_03321_));
 sg13g2_o21ai_1 _20109_ (.B1(_03311_),
    .Y(_03323_),
    .A1(_03310_),
    .A2(_03313_));
 sg13g2_nand2_1 _20110_ (.Y(_03324_),
    .A(_03322_),
    .B(_03323_));
 sg13g2_xnor2_1 _20111_ (.Y(_03325_),
    .A(_03322_),
    .B(_03323_));
 sg13g2_or2_1 _20112_ (.X(_03326_),
    .B(_03325_),
    .A(_03316_));
 sg13g2_nand2_1 _20113_ (.Y(_03327_),
    .A(net6023),
    .B(_03326_));
 sg13g2_a21oi_1 _20114_ (.A1(_03316_),
    .A2(_03325_),
    .Y(_01152_),
    .B1(_03327_));
 sg13g2_nand2_1 _20115_ (.Y(_03328_),
    .A(_03324_),
    .B(_03326_));
 sg13g2_nand2_1 _20116_ (.Y(_03329_),
    .A(\atari2600.tia.audv0[3] ),
    .B(\atari2600.tia.audio_l ));
 sg13g2_and3_1 _20117_ (.X(_03330_),
    .A(\atari2600.tia.audv1[3] ),
    .B(net5832),
    .C(\audio_pwm_accumulator[3] ));
 sg13g2_nand3_1 _20118_ (.B(net5832),
    .C(\audio_pwm_accumulator[3] ),
    .A(\atari2600.tia.audv1[3] ),
    .Y(_03331_));
 sg13g2_a21oi_1 _20119_ (.A1(\atari2600.tia.audv1[3] ),
    .A2(net5832),
    .Y(_03332_),
    .B1(\audio_pwm_accumulator[3] ));
 sg13g2_nor2_1 _20120_ (.A(_03330_),
    .B(_03332_),
    .Y(_03333_));
 sg13g2_xnor2_1 _20121_ (.Y(_03334_),
    .A(_03329_),
    .B(_03333_));
 sg13g2_o21ai_1 _20122_ (.B1(_03319_),
    .Y(_03335_),
    .A1(_03317_),
    .A2(_03320_));
 sg13g2_nand2_1 _20123_ (.Y(_03336_),
    .A(_03334_),
    .B(_03335_));
 sg13g2_xor2_1 _20124_ (.B(_03335_),
    .A(_03334_),
    .X(_03337_));
 sg13g2_nand2_1 _20125_ (.Y(_03338_),
    .A(_03328_),
    .B(_03337_));
 sg13g2_o21ai_1 _20126_ (.B1(net6022),
    .Y(_03339_),
    .A1(_03328_),
    .A2(_03337_));
 sg13g2_nor2b_1 _20127_ (.A(_03339_),
    .B_N(_03338_),
    .Y(_01153_));
 sg13g2_o21ai_1 _20128_ (.B1(_03331_),
    .Y(_03340_),
    .A1(_03329_),
    .A2(_03332_));
 sg13g2_nand2_1 _20129_ (.Y(_03341_),
    .A(net7360),
    .B(_03340_));
 sg13g2_xnor2_1 _20130_ (.Y(_03342_),
    .A(net7360),
    .B(_03340_));
 sg13g2_nand3_1 _20131_ (.B(_03338_),
    .C(_03342_),
    .A(_03336_),
    .Y(_03343_));
 sg13g2_a21o_1 _20132_ (.A2(_03338_),
    .A1(_03336_),
    .B1(_03342_),
    .X(_03344_));
 sg13g2_and3_1 _20133_ (.X(_01154_),
    .A(net6023),
    .B(_03343_),
    .C(_03344_));
 sg13g2_a21oi_2 _20134_ (.B1(net5987),
    .Y(_01155_),
    .A2(_03344_),
    .A1(_03341_));
 sg13g2_xnor2_1 _20135_ (.Y(_03345_),
    .A(\frame_counter[2] ),
    .B(net7179));
 sg13g2_xnor2_1 _20136_ (.Y(_03346_),
    .A(\frame_counter[1] ),
    .B(\hvsync_gen.hpos[0] ));
 sg13g2_nand2_1 _20137_ (.Y(_03347_),
    .A(_03345_),
    .B(_03346_));
 sg13g2_nor3_2 _20138_ (.A(net5871),
    .B(net5928),
    .C(net5839),
    .Y(_03348_));
 sg13g2_and4_2 _20139_ (.A(_08694_),
    .B(_08696_),
    .C(_03232_),
    .D(_03348_),
    .X(_03349_));
 sg13g2_nand4_1 _20140_ (.B(_08696_),
    .C(_03232_),
    .A(_08694_),
    .Y(_03350_),
    .D(_03348_));
 sg13g2_and3_1 _20141_ (.X(_01156_),
    .A(net2901),
    .B(net5456),
    .C(net5403));
 sg13g2_nor2_1 _20142_ (.A(net5843),
    .B(_08687_),
    .Y(_03351_));
 sg13g2_mux4_1 _20143_ (.S0(net5923),
    .A0(\scanline[156][5] ),
    .A1(\scanline[157][5] ),
    .A2(\scanline[158][5] ),
    .A3(\scanline[159][5] ),
    .S1(net5868),
    .X(_03352_));
 sg13g2_o21ai_1 _20144_ (.B1(net5844),
    .Y(_03353_),
    .A1(net5526),
    .A2(_03352_));
 sg13g2_mux4_1 _20145_ (.S0(net5910),
    .A0(\scanline[144][5] ),
    .A1(\scanline[145][5] ),
    .A2(\scanline[146][5] ),
    .A3(\scanline[147][5] ),
    .S1(net5854),
    .X(_03354_));
 sg13g2_nor2_1 _20146_ (.A(net5515),
    .B(_03354_),
    .Y(_03355_));
 sg13g2_nor2b_1 _20147_ (.A(net5850),
    .B_N(net5849),
    .Y(_03356_));
 sg13g2_nand2b_1 _20148_ (.Y(_03357_),
    .B(net5849),
    .A_N(net5850));
 sg13g2_mux4_1 _20149_ (.S0(net5922),
    .A0(\scanline[152][5] ),
    .A1(\scanline[153][5] ),
    .A2(\scanline[154][5] ),
    .A3(\scanline[155][5] ),
    .S1(net5866),
    .X(_03358_));
 sg13g2_nor2_1 _20150_ (.A(net5484),
    .B(_03358_),
    .Y(_03359_));
 sg13g2_mux4_1 _20151_ (.S0(net5924),
    .A0(\scanline[148][5] ),
    .A1(\scanline[149][5] ),
    .A2(\scanline[150][5] ),
    .A3(\scanline[151][5] ),
    .S1(net5867),
    .X(_03360_));
 sg13g2_nor2_1 _20152_ (.A(net5498),
    .B(_03360_),
    .Y(_03361_));
 sg13g2_nor4_1 _20153_ (.A(_03353_),
    .B(_03355_),
    .C(_03359_),
    .D(_03361_),
    .Y(_03362_));
 sg13g2_mux4_1 _20154_ (.S0(net5910),
    .A0(\scanline[128][5] ),
    .A1(\scanline[129][5] ),
    .A2(\scanline[130][5] ),
    .A3(\scanline[131][5] ),
    .S1(net5854),
    .X(_03363_));
 sg13g2_nor2_1 _20155_ (.A(net5514),
    .B(_03363_),
    .Y(_03364_));
 sg13g2_mux4_1 _20156_ (.S0(net5910),
    .A0(\scanline[136][5] ),
    .A1(\scanline[137][5] ),
    .A2(\scanline[138][5] ),
    .A3(\scanline[139][5] ),
    .S1(net5854),
    .X(_03365_));
 sg13g2_nor2_1 _20157_ (.A(net5483),
    .B(_03365_),
    .Y(_03366_));
 sg13g2_mux4_1 _20158_ (.S0(net5923),
    .A0(\scanline[140][5] ),
    .A1(\scanline[141][5] ),
    .A2(\scanline[142][5] ),
    .A3(\scanline[143][5] ),
    .S1(net5868),
    .X(_03367_));
 sg13g2_nor2_1 _20159_ (.A(net5525),
    .B(_03367_),
    .Y(_03368_));
 sg13g2_mux4_1 _20160_ (.S0(net5909),
    .A0(\scanline[132][5] ),
    .A1(\scanline[133][5] ),
    .A2(\scanline[134][5] ),
    .A3(\scanline[135][5] ),
    .S1(net5853),
    .X(_03369_));
 sg13g2_o21ai_1 _20161_ (.B1(net5553),
    .Y(_03370_),
    .A1(net5497),
    .A2(_03369_));
 sg13g2_nor4_2 _20162_ (.A(_03364_),
    .B(_03366_),
    .C(_03368_),
    .Y(_03371_),
    .D(_03370_));
 sg13g2_or2_1 _20163_ (.X(_03372_),
    .B(_03371_),
    .A(_03362_));
 sg13g2_mux4_1 _20164_ (.S0(net5954),
    .A0(\scanline[100][5] ),
    .A1(\scanline[101][5] ),
    .A2(\scanline[102][5] ),
    .A3(\scanline[103][5] ),
    .S1(net5895),
    .X(_03373_));
 sg13g2_mux4_1 _20165_ (.S0(net5955),
    .A0(\scanline[104][5] ),
    .A1(\scanline[105][5] ),
    .A2(\scanline[106][5] ),
    .A3(\scanline[107][5] ),
    .S1(net5896),
    .X(_03374_));
 sg13g2_mux4_1 _20166_ (.S0(net5949),
    .A0(\scanline[108][5] ),
    .A1(\scanline[109][5] ),
    .A2(\scanline[110][5] ),
    .A3(\scanline[111][5] ),
    .S1(net5891),
    .X(_03375_));
 sg13g2_mux4_1 _20167_ (.S0(net5952),
    .A0(\scanline[96][5] ),
    .A1(\scanline[97][5] ),
    .A2(\scanline[98][5] ),
    .A3(\scanline[99][5] ),
    .S1(net5893),
    .X(_03376_));
 sg13g2_a22oi_1 _20168_ (.Y(_03377_),
    .B1(_03374_),
    .B2(net5493),
    .A2(_03373_),
    .A1(net5502));
 sg13g2_a221oi_1 _20169_ (.B2(net5519),
    .C1(net5847),
    .B1(_03376_),
    .A1(net5535),
    .Y(_03378_),
    .A2(_03375_));
 sg13g2_nand2_1 _20170_ (.Y(_03379_),
    .A(_03377_),
    .B(_03378_));
 sg13g2_mux4_1 _20171_ (.S0(net5964),
    .A0(\scanline[116][5] ),
    .A1(\scanline[117][5] ),
    .A2(\scanline[118][5] ),
    .A3(\scanline[119][5] ),
    .S1(net5903),
    .X(_03380_));
 sg13g2_a21oi_1 _20172_ (.A1(net5507),
    .A2(_03380_),
    .Y(_03381_),
    .B1(net5555));
 sg13g2_mux4_1 _20173_ (.S0(net5966),
    .A0(\scanline[120][5] ),
    .A1(\scanline[121][5] ),
    .A2(\scanline[122][5] ),
    .A3(\scanline[123][5] ),
    .S1(net5904),
    .X(_03382_));
 sg13g2_nor2b_1 _20174_ (.A(net5961),
    .B_N(\scanline[126][5] ),
    .Y(_03383_));
 sg13g2_a21oi_1 _20175_ (.A1(net5961),
    .A2(\scanline[127][5] ),
    .Y(_03384_),
    .B1(_03383_));
 sg13g2_nand2b_1 _20176_ (.Y(_03385_),
    .B(\scanline[124][5] ),
    .A_N(net5961));
 sg13g2_a21oi_1 _20177_ (.A1(net5961),
    .A2(\scanline[125][5] ),
    .Y(_03386_),
    .B1(net5900));
 sg13g2_a221oi_1 _20178_ (.B2(_03386_),
    .C1(net5528),
    .B1(_03385_),
    .A1(net5900),
    .Y(_03387_),
    .A2(_03384_));
 sg13g2_mux4_1 _20179_ (.S0(net5962),
    .A0(\scanline[112][5] ),
    .A1(\scanline[113][5] ),
    .A2(\scanline[114][5] ),
    .A3(\scanline[115][5] ),
    .S1(net5900),
    .X(_03388_));
 sg13g2_a221oi_1 _20180_ (.B2(net5524),
    .C1(_03387_),
    .B1(_03388_),
    .A1(net5492),
    .Y(_03389_),
    .A2(_03382_));
 sg13g2_a21oi_2 _20181_ (.B1(_08117_),
    .Y(_03390_),
    .A2(_03389_),
    .A1(_03381_));
 sg13g2_nand2_2 _20182_ (.Y(_03391_),
    .A(_03379_),
    .B(_03390_));
 sg13g2_nor2_1 _20183_ (.A(net5842),
    .B(net5554),
    .Y(_03392_));
 sg13g2_nand2_2 _20184_ (.Y(_03393_),
    .A(_08117_),
    .B(net5847));
 sg13g2_mux4_1 _20185_ (.S0(net5963),
    .A0(\scanline[92][5] ),
    .A1(\scanline[93][5] ),
    .A2(\scanline[94][5] ),
    .A3(\scanline[95][5] ),
    .S1(net5901),
    .X(_03394_));
 sg13g2_mux4_1 _20186_ (.S0(net5960),
    .A0(\scanline[84][5] ),
    .A1(\scanline[85][5] ),
    .A2(\scanline[86][5] ),
    .A3(\scanline[87][5] ),
    .S1(net5899),
    .X(_03395_));
 sg13g2_a22oi_1 _20187_ (.Y(_03396_),
    .B1(_03395_),
    .B2(net5506),
    .A2(_03394_),
    .A1(net5534));
 sg13g2_mux4_1 _20188_ (.S0(net5944),
    .A0(\scanline[80][5] ),
    .A1(\scanline[81][5] ),
    .A2(\scanline[82][5] ),
    .A3(\scanline[83][5] ),
    .S1(net5887),
    .X(_03397_));
 sg13g2_mux4_1 _20189_ (.S0(net5942),
    .A0(\scanline[88][5] ),
    .A1(\scanline[89][5] ),
    .A2(\scanline[90][5] ),
    .A3(\scanline[91][5] ),
    .S1(net5886),
    .X(_03398_));
 sg13g2_a22oi_1 _20190_ (.Y(_03399_),
    .B1(_03398_),
    .B2(net5494),
    .A2(_03397_),
    .A1(net5520));
 sg13g2_a21oi_2 _20191_ (.B1(_03393_),
    .Y(_03400_),
    .A2(_03399_),
    .A1(_03396_));
 sg13g2_mux4_1 _20192_ (.S0(net5908),
    .A0(\scanline[76][5] ),
    .A1(\scanline[77][5] ),
    .A2(\scanline[78][5] ),
    .A3(\scanline[79][5] ),
    .S1(net5852),
    .X(_03401_));
 sg13g2_mux4_1 _20193_ (.S0(net5907),
    .A0(\scanline[72][5] ),
    .A1(\scanline[73][5] ),
    .A2(\scanline[74][5] ),
    .A3(\scanline[75][5] ),
    .S1(net5851),
    .X(_03402_));
 sg13g2_mux4_1 _20194_ (.S0(net5913),
    .A0(\scanline[68][5] ),
    .A1(\scanline[69][5] ),
    .A2(\scanline[70][5] ),
    .A3(\scanline[71][5] ),
    .S1(net5857),
    .X(_03403_));
 sg13g2_mux4_1 _20195_ (.S0(net5914),
    .A0(\scanline[64][5] ),
    .A1(\scanline[65][5] ),
    .A2(\scanline[66][5] ),
    .A3(\scanline[67][5] ),
    .S1(net5858),
    .X(_03404_));
 sg13g2_a22oi_1 _20196_ (.Y(_03405_),
    .B1(_03404_),
    .B2(net5517),
    .A2(_03402_),
    .A1(net5486));
 sg13g2_a22oi_1 _20197_ (.Y(_03406_),
    .B1(_03403_),
    .B2(net5500),
    .A2(_03401_),
    .A1(net5529));
 sg13g2_a21oi_2 _20198_ (.B1(net5509),
    .Y(_03407_),
    .A2(_03406_),
    .A1(_03405_));
 sg13g2_nor3_1 _20199_ (.A(net5552),
    .B(_03400_),
    .C(_03407_),
    .Y(_03408_));
 sg13g2_nand2b_1 _20200_ (.Y(_03409_),
    .B(\scanline[36][5] ),
    .A_N(net5916));
 sg13g2_a21oi_1 _20201_ (.A1(net5916),
    .A2(\scanline[37][5] ),
    .Y(_03410_),
    .B1(net5860));
 sg13g2_nor2b_1 _20202_ (.A(net5915),
    .B_N(\scanline[38][5] ),
    .Y(_03411_));
 sg13g2_a21oi_1 _20203_ (.A1(net5915),
    .A2(\scanline[39][5] ),
    .Y(_03412_),
    .B1(_03411_));
 sg13g2_a221oi_1 _20204_ (.B2(net5859),
    .C1(net5499),
    .B1(_03412_),
    .A1(_03409_),
    .Y(_03413_),
    .A2(_03410_));
 sg13g2_mux4_1 _20205_ (.S0(net5919),
    .A0(\scanline[32][5] ),
    .A1(\scanline[33][5] ),
    .A2(\scanline[34][5] ),
    .A3(\scanline[35][5] ),
    .S1(net5862),
    .X(_03414_));
 sg13g2_mux4_1 _20206_ (.S0(net5915),
    .A0(\scanline[40][5] ),
    .A1(\scanline[41][5] ),
    .A2(\scanline[42][5] ),
    .A3(\scanline[43][5] ),
    .S1(net5859),
    .X(_03415_));
 sg13g2_mux4_1 _20207_ (.S0(net5919),
    .A0(\scanline[44][5] ),
    .A1(\scanline[45][5] ),
    .A2(\scanline[46][5] ),
    .A3(\scanline[47][5] ),
    .S1(net5862),
    .X(_03416_));
 sg13g2_a21oi_1 _20208_ (.A1(net5518),
    .A2(_03414_),
    .Y(_03417_),
    .B1(net5847));
 sg13g2_a221oi_1 _20209_ (.B2(net5530),
    .C1(_03413_),
    .B1(_03416_),
    .A1(net5487),
    .Y(_03418_),
    .A2(_03415_));
 sg13g2_nand2_1 _20210_ (.Y(_03419_),
    .A(_03417_),
    .B(_03418_));
 sg13g2_mux4_1 _20211_ (.S0(net5954),
    .A0(\scanline[52][5] ),
    .A1(\scanline[53][5] ),
    .A2(\scanline[54][5] ),
    .A3(\scanline[55][5] ),
    .S1(net5898),
    .X(_03420_));
 sg13g2_nand2_1 _20212_ (.Y(_03421_),
    .A(net5503),
    .B(_03420_));
 sg13g2_mux4_1 _20213_ (.S0(net5927),
    .A0(\scanline[48][5] ),
    .A1(\scanline[49][5] ),
    .A2(\scanline[50][5] ),
    .A3(\scanline[51][5] ),
    .S1(net5870),
    .X(_03422_));
 sg13g2_mux4_1 _20214_ (.S0(net5936),
    .A0(\scanline[56][5] ),
    .A1(\scanline[57][5] ),
    .A2(\scanline[58][5] ),
    .A3(\scanline[59][5] ),
    .S1(net5880),
    .X(_03423_));
 sg13g2_mux4_1 _20215_ (.S0(net5949),
    .A0(\scanline[60][5] ),
    .A1(\scanline[61][5] ),
    .A2(\scanline[62][5] ),
    .A3(\scanline[63][5] ),
    .S1(net5891),
    .X(_03424_));
 sg13g2_a21oi_1 _20216_ (.A1(net5488),
    .A2(_03423_),
    .Y(_03425_),
    .B1(net5554));
 sg13g2_a22oi_1 _20217_ (.Y(_03426_),
    .B1(_03424_),
    .B2(net5531),
    .A2(_03422_),
    .A1(net5519));
 sg13g2_nand3_1 _20218_ (.B(_03425_),
    .C(_03426_),
    .A(_03421_),
    .Y(_03427_));
 sg13g2_nand3_1 _20219_ (.B(_03419_),
    .C(_03427_),
    .A(net5842),
    .Y(_03428_));
 sg13g2_mux4_1 _20220_ (.S0(net5936),
    .A0(\scanline[12][5] ),
    .A1(\scanline[13][5] ),
    .A2(\scanline[14][5] ),
    .A3(\scanline[15][5] ),
    .S1(net5880),
    .X(_03429_));
 sg13g2_mux4_1 _20221_ (.S0(net5933),
    .A0(\scanline[4][5] ),
    .A1(\scanline[5][5] ),
    .A2(\scanline[6][5] ),
    .A3(\scanline[7][5] ),
    .S1(net5876),
    .X(_03430_));
 sg13g2_mux4_1 _20222_ (.S0(net5931),
    .A0(\scanline[8][5] ),
    .A1(\scanline[9][5] ),
    .A2(\scanline[10][5] ),
    .A3(\scanline[11][5] ),
    .S1(net5875),
    .X(_03431_));
 sg13g2_mux4_1 _20223_ (.S0(net5935),
    .A0(\scanline[0][5] ),
    .A1(\scanline[1][5] ),
    .A2(\scanline[2][5] ),
    .A3(\scanline[3][5] ),
    .S1(net5878),
    .X(_03432_));
 sg13g2_a22oi_1 _20224_ (.Y(_03433_),
    .B1(_03432_),
    .B2(net5521),
    .A2(_03430_),
    .A1(net5504));
 sg13g2_a22oi_1 _20225_ (.Y(_03434_),
    .B1(_03431_),
    .B2(net5490),
    .A2(_03429_),
    .A1(net5532));
 sg13g2_a21oi_1 _20226_ (.A1(_03433_),
    .A2(_03434_),
    .Y(_03435_),
    .B1(net5510));
 sg13g2_mux4_1 _20227_ (.S0(net5941),
    .A0(\scanline[28][5] ),
    .A1(\scanline[29][5] ),
    .A2(\scanline[30][5] ),
    .A3(\scanline[31][5] ),
    .S1(net5885),
    .X(_03436_));
 sg13g2_mux4_1 _20228_ (.S0(net5939),
    .A0(\scanline[20][5] ),
    .A1(\scanline[21][5] ),
    .A2(\scanline[22][5] ),
    .A3(\scanline[23][5] ),
    .S1(net5883),
    .X(_03437_));
 sg13g2_mux4_1 _20229_ (.S0(net5941),
    .A0(\scanline[24][5] ),
    .A1(\scanline[25][5] ),
    .A2(\scanline[26][5] ),
    .A3(\scanline[27][5] ),
    .S1(net5885),
    .X(_03438_));
 sg13g2_mux4_1 _20230_ (.S0(net5939),
    .A0(\scanline[16][5] ),
    .A1(\scanline[17][5] ),
    .A2(\scanline[18][5] ),
    .A3(\scanline[19][5] ),
    .S1(net5883),
    .X(_03439_));
 sg13g2_a22oi_1 _20231_ (.Y(_03440_),
    .B1(_03439_),
    .B2(net5520),
    .A2(_03437_),
    .A1(net5505));
 sg13g2_a22oi_1 _20232_ (.Y(_03441_),
    .B1(_03438_),
    .B2(net5489),
    .A2(_03436_),
    .A1(net5533));
 sg13g2_a21oi_2 _20233_ (.B1(net5455),
    .Y(_03442_),
    .A2(_03441_),
    .A1(_03440_));
 sg13g2_nor3_2 _20234_ (.A(net5841),
    .B(_03435_),
    .C(_03442_),
    .Y(_03443_));
 sg13g2_a221oi_1 _20235_ (.B2(_03443_),
    .C1(\hvsync_gen.hpos[9] ),
    .B1(_03428_),
    .A1(_03391_),
    .Y(_03444_),
    .A2(_03408_));
 sg13g2_a21oi_2 _20236_ (.B1(_03444_),
    .Y(_03445_),
    .A2(_03372_),
    .A1(_03351_));
 sg13g2_inv_1 _20237_ (.Y(_03446_),
    .A(net5299));
 sg13g2_mux4_1 _20238_ (.S0(net5922),
    .A0(\scanline[156][4] ),
    .A1(\scanline[157][4] ),
    .A2(\scanline[158][4] ),
    .A3(\scanline[159][4] ),
    .S1(net5866),
    .X(_03447_));
 sg13g2_o21ai_1 _20239_ (.B1(net5844),
    .Y(_03448_),
    .A1(net5526),
    .A2(_03447_));
 sg13g2_mux4_1 _20240_ (.S0(net5918),
    .A0(\scanline[144][4] ),
    .A1(\scanline[145][4] ),
    .A2(\scanline[146][4] ),
    .A3(\scanline[147][4] ),
    .S1(net5864),
    .X(_03449_));
 sg13g2_nor2_1 _20241_ (.A(net5515),
    .B(_03449_),
    .Y(_03450_));
 sg13g2_mux4_1 _20242_ (.S0(net5922),
    .A0(\scanline[152][4] ),
    .A1(\scanline[153][4] ),
    .A2(\scanline[154][4] ),
    .A3(\scanline[155][4] ),
    .S1(net5866),
    .X(_03451_));
 sg13g2_nor2_1 _20243_ (.A(net5483),
    .B(_03451_),
    .Y(_03452_));
 sg13g2_mux4_1 _20244_ (.S0(net5924),
    .A0(\scanline[148][4] ),
    .A1(\scanline[149][4] ),
    .A2(\scanline[150][4] ),
    .A3(\scanline[151][4] ),
    .S1(net5867),
    .X(_03453_));
 sg13g2_nor2_1 _20245_ (.A(net5498),
    .B(_03453_),
    .Y(_03454_));
 sg13g2_nor4_1 _20246_ (.A(_03448_),
    .B(_03450_),
    .C(_03452_),
    .D(_03454_),
    .Y(_03455_));
 sg13g2_mux4_1 _20247_ (.S0(net5918),
    .A0(\scanline[128][4] ),
    .A1(\scanline[129][4] ),
    .A2(\scanline[130][4] ),
    .A3(\scanline[131][4] ),
    .S1(net5864),
    .X(_03456_));
 sg13g2_nor2_1 _20248_ (.A(net5514),
    .B(_03456_),
    .Y(_03457_));
 sg13g2_mux4_1 _20249_ (.S0(net5909),
    .A0(\scanline[136][4] ),
    .A1(\scanline[137][4] ),
    .A2(\scanline[138][4] ),
    .A3(\scanline[139][4] ),
    .S1(net5853),
    .X(_03458_));
 sg13g2_nor2_1 _20250_ (.A(net5483),
    .B(_03458_),
    .Y(_03459_));
 sg13g2_mux4_1 _20251_ (.S0(net5923),
    .A0(\scanline[140][4] ),
    .A1(\scanline[141][4] ),
    .A2(\scanline[142][4] ),
    .A3(\scanline[143][4] ),
    .S1(net5868),
    .X(_03460_));
 sg13g2_nor2_1 _20252_ (.A(net5525),
    .B(_03460_),
    .Y(_03461_));
 sg13g2_mux4_1 _20253_ (.S0(net5909),
    .A0(\scanline[132][4] ),
    .A1(\scanline[133][4] ),
    .A2(\scanline[134][4] ),
    .A3(\scanline[135][4] ),
    .S1(net5853),
    .X(_03462_));
 sg13g2_o21ai_1 _20254_ (.B1(net5553),
    .Y(_03463_),
    .A1(net5497),
    .A2(_03462_));
 sg13g2_nor4_2 _20255_ (.A(_03457_),
    .B(_03459_),
    .C(_03461_),
    .Y(_03464_),
    .D(_03463_));
 sg13g2_o21ai_1 _20256_ (.B1(_08686_),
    .Y(_03465_),
    .A1(_03455_),
    .A2(_03464_));
 sg13g2_mux4_1 _20257_ (.S0(net5955),
    .A0(\scanline[104][4] ),
    .A1(\scanline[105][4] ),
    .A2(\scanline[106][4] ),
    .A3(\scanline[107][4] ),
    .S1(net5896),
    .X(_03466_));
 sg13g2_a21oi_1 _20258_ (.A1(net5493),
    .A2(_03466_),
    .Y(_03467_),
    .B1(net5848));
 sg13g2_nor2b_1 _20259_ (.A(net5949),
    .B_N(\scanline[110][4] ),
    .Y(_03468_));
 sg13g2_a21oi_1 _20260_ (.A1(net5949),
    .A2(\scanline[111][4] ),
    .Y(_03469_),
    .B1(_03468_));
 sg13g2_nand2b_1 _20261_ (.Y(_03470_),
    .B(\scanline[108][4] ),
    .A_N(net5949));
 sg13g2_a21oi_1 _20262_ (.A1(net5949),
    .A2(\scanline[109][4] ),
    .Y(_03471_),
    .B1(net5890));
 sg13g2_a221oi_1 _20263_ (.B2(_03471_),
    .C1(_08689_),
    .B1(_03470_),
    .A1(net5890),
    .Y(_03472_),
    .A2(_03469_));
 sg13g2_mux4_1 _20264_ (.S0(net5952),
    .A0(\scanline[96][4] ),
    .A1(\scanline[97][4] ),
    .A2(\scanline[98][4] ),
    .A3(\scanline[99][4] ),
    .S1(net5893),
    .X(_03473_));
 sg13g2_mux4_1 _20265_ (.S0(net5957),
    .A0(\scanline[100][4] ),
    .A1(\scanline[101][4] ),
    .A2(\scanline[102][4] ),
    .A3(\scanline[103][4] ),
    .S1(net5897),
    .X(_03474_));
 sg13g2_a22oi_1 _20266_ (.Y(_03475_),
    .B1(_03474_),
    .B2(net5507),
    .A2(_03473_),
    .A1(net5523));
 sg13g2_nand3b_1 _20267_ (.B(_03475_),
    .C(_03467_),
    .Y(_03476_),
    .A_N(_03472_));
 sg13g2_mux4_1 _20268_ (.S0(net5964),
    .A0(\scanline[116][4] ),
    .A1(\scanline[117][4] ),
    .A2(\scanline[118][4] ),
    .A3(\scanline[119][4] ),
    .S1(net5903),
    .X(_03477_));
 sg13g2_mux4_1 _20269_ (.S0(net5959),
    .A0(\scanline[124][4] ),
    .A1(\scanline[125][4] ),
    .A2(\scanline[126][4] ),
    .A3(\scanline[127][4] ),
    .S1(net5902),
    .X(_03478_));
 sg13g2_mux4_1 _20270_ (.S0(net5966),
    .A0(\scanline[120][4] ),
    .A1(\scanline[121][4] ),
    .A2(\scanline[122][4] ),
    .A3(\scanline[123][4] ),
    .S1(net5905),
    .X(_03479_));
 sg13g2_mux4_1 _20271_ (.S0(net5962),
    .A0(\scanline[112][4] ),
    .A1(\scanline[113][4] ),
    .A2(\scanline[114][4] ),
    .A3(\scanline[115][4] ),
    .S1(net5901),
    .X(_03480_));
 sg13g2_nand2_1 _20272_ (.Y(_03481_),
    .A(net5522),
    .B(_03480_));
 sg13g2_a21oi_1 _20273_ (.A1(net5491),
    .A2(_03479_),
    .Y(_03482_),
    .B1(net5555));
 sg13g2_a22oi_1 _20274_ (.Y(_03483_),
    .B1(_03478_),
    .B2(net5536),
    .A2(_03477_),
    .A1(net5506));
 sg13g2_nand3_1 _20275_ (.B(_03482_),
    .C(_03483_),
    .A(_03481_),
    .Y(_03484_));
 sg13g2_nand3_1 _20276_ (.B(_03476_),
    .C(_03484_),
    .A(net5842),
    .Y(_03485_));
 sg13g2_mux4_1 _20277_ (.S0(net5963),
    .A0(\scanline[92][4] ),
    .A1(\scanline[93][4] ),
    .A2(\scanline[94][4] ),
    .A3(\scanline[95][4] ),
    .S1(net5901),
    .X(_03486_));
 sg13g2_mux4_1 _20278_ (.S0(net5951),
    .A0(\scanline[84][4] ),
    .A1(\scanline[85][4] ),
    .A2(\scanline[86][4] ),
    .A3(\scanline[87][4] ),
    .S1(net5892),
    .X(_03487_));
 sg13g2_mux4_1 _20279_ (.S0(net5945),
    .A0(\scanline[80][4] ),
    .A1(\scanline[81][4] ),
    .A2(\scanline[82][4] ),
    .A3(\scanline[83][4] ),
    .S1(net5888),
    .X(_03488_));
 sg13g2_mux4_1 _20280_ (.S0(net5943),
    .A0(\scanline[88][4] ),
    .A1(\scanline[89][4] ),
    .A2(\scanline[90][4] ),
    .A3(\scanline[91][4] ),
    .S1(net5889),
    .X(_03489_));
 sg13g2_a22oi_1 _20281_ (.Y(_03490_),
    .B1(_03489_),
    .B2(net5492),
    .A2(_03487_),
    .A1(net5507));
 sg13g2_a22oi_1 _20282_ (.Y(_03491_),
    .B1(_03488_),
    .B2(net5522),
    .A2(_03486_),
    .A1(net5534));
 sg13g2_a21oi_2 _20283_ (.B1(_03393_),
    .Y(_03492_),
    .A2(_03491_),
    .A1(_03490_));
 sg13g2_mux4_1 _20284_ (.S0(net5913),
    .A0(\scanline[64][4] ),
    .A1(\scanline[65][4] ),
    .A2(\scanline[66][4] ),
    .A3(\scanline[67][4] ),
    .S1(net5857),
    .X(_03493_));
 sg13g2_mux4_1 _20285_ (.S0(net5907),
    .A0(\scanline[72][4] ),
    .A1(\scanline[73][4] ),
    .A2(\scanline[74][4] ),
    .A3(\scanline[75][4] ),
    .S1(net5851),
    .X(_03494_));
 sg13g2_mux4_1 _20286_ (.S0(net5913),
    .A0(\scanline[68][4] ),
    .A1(\scanline[69][4] ),
    .A2(\scanline[70][4] ),
    .A3(\scanline[71][4] ),
    .S1(net5857),
    .X(_03495_));
 sg13g2_mux4_1 _20287_ (.S0(net5912),
    .A0(\scanline[76][4] ),
    .A1(\scanline[77][4] ),
    .A2(\scanline[78][4] ),
    .A3(\scanline[79][4] ),
    .S1(net5856),
    .X(_03496_));
 sg13g2_a22oi_1 _20288_ (.Y(_03497_),
    .B1(_03496_),
    .B2(net5529),
    .A2(_03494_),
    .A1(net5486));
 sg13g2_a22oi_1 _20289_ (.Y(_03498_),
    .B1(_03495_),
    .B2(net5500),
    .A2(_03493_),
    .A1(net5517));
 sg13g2_a21oi_2 _20290_ (.B1(net5509),
    .Y(_03499_),
    .A2(_03498_),
    .A1(_03497_));
 sg13g2_nor3_1 _20291_ (.A(net5552),
    .B(_03492_),
    .C(_03499_),
    .Y(_03500_));
 sg13g2_mux4_1 _20292_ (.S0(net5950),
    .A0(\scanline[60][4] ),
    .A1(\scanline[61][4] ),
    .A2(\scanline[62][4] ),
    .A3(\scanline[63][4] ),
    .S1(net5890),
    .X(_03501_));
 sg13g2_a21oi_1 _20293_ (.A1(net5530),
    .A2(_03501_),
    .Y(_03502_),
    .B1(net5554));
 sg13g2_mux4_1 _20294_ (.S0(net5926),
    .A0(\scanline[48][4] ),
    .A1(\scanline[49][4] ),
    .A2(\scanline[50][4] ),
    .A3(\scanline[51][4] ),
    .S1(net5870),
    .X(_03503_));
 sg13g2_nor2b_1 _20295_ (.A(net5949),
    .B_N(\scanline[54][4] ),
    .Y(_03504_));
 sg13g2_a21oi_1 _20296_ (.A1(net5948),
    .A2(\scanline[55][4] ),
    .Y(_03505_),
    .B1(_03504_));
 sg13g2_nand2b_1 _20297_ (.Y(_03506_),
    .B(\scanline[52][4] ),
    .A_N(net5948));
 sg13g2_a21oi_1 _20298_ (.A1(net5948),
    .A2(\scanline[53][4] ),
    .Y(_03507_),
    .B1(net5872));
 sg13g2_a221oi_1 _20299_ (.B2(_03507_),
    .C1(net5499),
    .B1(_03506_),
    .A1(net5891),
    .Y(_03508_),
    .A2(_03505_));
 sg13g2_mux4_1 _20300_ (.S0(net5950),
    .A0(\scanline[56][4] ),
    .A1(\scanline[57][4] ),
    .A2(\scanline[58][4] ),
    .A3(\scanline[59][4] ),
    .S1(net5890),
    .X(_03509_));
 sg13g2_a221oi_1 _20301_ (.B2(net5488),
    .C1(_03508_),
    .B1(_03509_),
    .A1(_08692_),
    .Y(_03510_),
    .A2(_03503_));
 sg13g2_mux4_1 _20302_ (.S0(net5920),
    .A0(\scanline[44][4] ),
    .A1(\scanline[45][4] ),
    .A2(\scanline[46][4] ),
    .A3(\scanline[47][4] ),
    .S1(net5863),
    .X(_03511_));
 sg13g2_mux4_1 _20303_ (.S0(net5936),
    .A0(\scanline[32][4] ),
    .A1(\scanline[33][4] ),
    .A2(\scanline[34][4] ),
    .A3(\scanline[35][4] ),
    .S1(net5880),
    .X(_03512_));
 sg13g2_mux4_1 _20304_ (.S0(net5931),
    .A0(\scanline[36][4] ),
    .A1(\scanline[37][4] ),
    .A2(\scanline[38][4] ),
    .A3(\scanline[39][4] ),
    .S1(net5875),
    .X(_03513_));
 sg13g2_a21oi_1 _20305_ (.A1(net5916),
    .A2(\scanline[41][4] ),
    .Y(_03514_),
    .B1(net5860));
 sg13g2_o21ai_1 _20306_ (.B1(_03514_),
    .Y(_03515_),
    .A1(net5916),
    .A2(_08129_));
 sg13g2_nor2b_1 _20307_ (.A(net5919),
    .B_N(\scanline[42][4] ),
    .Y(_03516_));
 sg13g2_a21oi_1 _20308_ (.A1(net5919),
    .A2(\scanline[43][4] ),
    .Y(_03517_),
    .B1(_03516_));
 sg13g2_a21oi_1 _20309_ (.A1(net5862),
    .A2(_03517_),
    .Y(_03518_),
    .B1(net5484));
 sg13g2_a22oi_1 _20310_ (.Y(_03519_),
    .B1(_03513_),
    .B2(net5501),
    .A2(_03512_),
    .A1(net5518));
 sg13g2_a221oi_1 _20311_ (.B2(_03518_),
    .C1(net5845),
    .B1(_03515_),
    .A1(net5530),
    .Y(_03520_),
    .A2(_03511_));
 sg13g2_a221oi_1 _20312_ (.B2(_03520_),
    .C1(_08117_),
    .B1(_03519_),
    .A1(_03502_),
    .Y(_03521_),
    .A2(_03510_));
 sg13g2_mux4_1 _20313_ (.S0(net5933),
    .A0(\scanline[4][4] ),
    .A1(\scanline[5][4] ),
    .A2(\scanline[6][4] ),
    .A3(\scanline[7][4] ),
    .S1(net5876),
    .X(_03522_));
 sg13g2_mux4_1 _20314_ (.S0(net5935),
    .A0(\scanline[12][4] ),
    .A1(\scanline[13][4] ),
    .A2(\scanline[14][4] ),
    .A3(\scanline[15][4] ),
    .S1(net5878),
    .X(_03523_));
 sg13g2_a22oi_1 _20315_ (.Y(_03524_),
    .B1(_03523_),
    .B2(net5532),
    .A2(_03522_),
    .A1(net5504));
 sg13g2_mux4_1 _20316_ (.S0(net5935),
    .A0(\scanline[0][4] ),
    .A1(\scanline[1][4] ),
    .A2(\scanline[2][4] ),
    .A3(\scanline[3][4] ),
    .S1(net5878),
    .X(_03525_));
 sg13g2_mux4_1 _20317_ (.S0(net5934),
    .A0(\scanline[8][4] ),
    .A1(\scanline[9][4] ),
    .A2(\scanline[10][4] ),
    .A3(\scanline[11][4] ),
    .S1(net5877),
    .X(_03526_));
 sg13g2_a22oi_1 _20318_ (.Y(_03527_),
    .B1(_03526_),
    .B2(net5490),
    .A2(_03525_),
    .A1(net5521));
 sg13g2_a21oi_2 _20319_ (.B1(net5510),
    .Y(_03528_),
    .A2(_03527_),
    .A1(_03524_));
 sg13g2_mux4_1 _20320_ (.S0(net5941),
    .A0(\scanline[24][4] ),
    .A1(\scanline[25][4] ),
    .A2(\scanline[26][4] ),
    .A3(\scanline[27][4] ),
    .S1(net5885),
    .X(_03529_));
 sg13g2_mux4_1 _20321_ (.S0(net5942),
    .A0(\scanline[28][4] ),
    .A1(\scanline[29][4] ),
    .A2(\scanline[30][4] ),
    .A3(\scanline[31][4] ),
    .S1(net5886),
    .X(_03530_));
 sg13g2_a22oi_1 _20322_ (.Y(_03531_),
    .B1(_03530_),
    .B2(net5532),
    .A2(_03529_),
    .A1(net5494));
 sg13g2_mux4_1 _20323_ (.S0(net5939),
    .A0(\scanline[16][4] ),
    .A1(\scanline[17][4] ),
    .A2(\scanline[18][4] ),
    .A3(\scanline[19][4] ),
    .S1(net5883),
    .X(_03532_));
 sg13g2_mux4_1 _20324_ (.S0(net5940),
    .A0(\scanline[20][4] ),
    .A1(\scanline[21][4] ),
    .A2(\scanline[22][4] ),
    .A3(\scanline[23][4] ),
    .S1(net5884),
    .X(_03533_));
 sg13g2_a22oi_1 _20325_ (.Y(_03534_),
    .B1(_03533_),
    .B2(net5505),
    .A2(_03532_),
    .A1(net5520));
 sg13g2_a21oi_2 _20326_ (.B1(net5455),
    .Y(_03535_),
    .A2(_03534_),
    .A1(_03531_));
 sg13g2_nor4_2 _20327_ (.A(net5841),
    .B(_03521_),
    .C(_03528_),
    .Y(_03536_),
    .D(_03535_));
 sg13g2_a21o_1 _20328_ (.A2(_03500_),
    .A1(_03485_),
    .B1(net5839),
    .X(_03537_));
 sg13g2_o21ai_1 _20329_ (.B1(_03465_),
    .Y(_03538_),
    .A1(_03536_),
    .A2(_03537_));
 sg13g2_and2_1 _20330_ (.A(net5513),
    .B(_03538_),
    .X(_03539_));
 sg13g2_nand2_1 _20331_ (.Y(_03540_),
    .A(net5513),
    .B(_03538_));
 sg13g2_nand2b_1 _20332_ (.Y(_03541_),
    .B(\scanline[36][3] ),
    .A_N(net5915));
 sg13g2_a21oi_1 _20333_ (.A1(net5932),
    .A2(\scanline[37][3] ),
    .Y(_03542_),
    .B1(net5860));
 sg13g2_nor2b_1 _20334_ (.A(net5932),
    .B_N(\scanline[38][3] ),
    .Y(_03543_));
 sg13g2_a21oi_1 _20335_ (.A1(net5932),
    .A2(\scanline[39][3] ),
    .Y(_03544_),
    .B1(_03543_));
 sg13g2_a221oi_1 _20336_ (.B2(net5859),
    .C1(net5499),
    .B1(_03544_),
    .A1(_03541_),
    .Y(_03545_),
    .A2(_03542_));
 sg13g2_mux4_1 _20337_ (.S0(net5919),
    .A0(\scanline[32][3] ),
    .A1(\scanline[33][3] ),
    .A2(\scanline[34][3] ),
    .A3(\scanline[35][3] ),
    .S1(net5862),
    .X(_03546_));
 sg13g2_mux4_1 _20338_ (.S0(net5920),
    .A0(\scanline[44][3] ),
    .A1(\scanline[45][3] ),
    .A2(\scanline[46][3] ),
    .A3(\scanline[47][3] ),
    .S1(net5863),
    .X(_03547_));
 sg13g2_mux4_1 _20339_ (.S0(net5915),
    .A0(\scanline[40][3] ),
    .A1(\scanline[41][3] ),
    .A2(\scanline[42][3] ),
    .A3(\scanline[43][3] ),
    .S1(net5859),
    .X(_03548_));
 sg13g2_a22oi_1 _20340_ (.Y(_03549_),
    .B1(_03548_),
    .B2(net5487),
    .A2(_03546_),
    .A1(net5518));
 sg13g2_a21oi_1 _20341_ (.A1(net5529),
    .A2(_03547_),
    .Y(_03550_),
    .B1(net5845));
 sg13g2_nand3b_1 _20342_ (.B(_03549_),
    .C(_03550_),
    .Y(_03551_),
    .A_N(_03545_));
 sg13g2_mux4_1 _20343_ (.S0(net5936),
    .A0(\scanline[56][3] ),
    .A1(\scanline[57][3] ),
    .A2(\scanline[58][3] ),
    .A3(\scanline[59][3] ),
    .S1(net5880),
    .X(_03552_));
 sg13g2_a21oi_1 _20344_ (.A1(net5487),
    .A2(_03552_),
    .Y(_03553_),
    .B1(net5554));
 sg13g2_mux4_1 _20345_ (.S0(net5929),
    .A0(\scanline[52][3] ),
    .A1(\scanline[53][3] ),
    .A2(\scanline[54][3] ),
    .A3(\scanline[55][3] ),
    .S1(net5873),
    .X(_03554_));
 sg13g2_and2_1 _20346_ (.A(net5502),
    .B(_03554_),
    .X(_03555_));
 sg13g2_mux4_1 _20347_ (.S0(net5927),
    .A0(\scanline[48][3] ),
    .A1(\scanline[49][3] ),
    .A2(\scanline[50][3] ),
    .A3(\scanline[51][3] ),
    .S1(net5872),
    .X(_03556_));
 sg13g2_mux4_1 _20348_ (.S0(net5948),
    .A0(\scanline[60][3] ),
    .A1(\scanline[61][3] ),
    .A2(\scanline[62][3] ),
    .A3(\scanline[63][3] ),
    .S1(net5891),
    .X(_03557_));
 sg13g2_a221oi_1 _20349_ (.B2(net5531),
    .C1(_03555_),
    .B1(_03557_),
    .A1(net5519),
    .Y(_03558_),
    .A2(_03556_));
 sg13g2_a21oi_1 _20350_ (.A1(_03553_),
    .A2(_03558_),
    .Y(_03559_),
    .B1(_08117_));
 sg13g2_mux4_1 _20351_ (.S0(net5938),
    .A0(\scanline[24][3] ),
    .A1(\scanline[25][3] ),
    .A2(\scanline[26][3] ),
    .A3(\scanline[27][3] ),
    .S1(net5882),
    .X(_03560_));
 sg13g2_mux4_1 _20352_ (.S0(net5940),
    .A0(\scanline[28][3] ),
    .A1(\scanline[29][3] ),
    .A2(\scanline[30][3] ),
    .A3(\scanline[31][3] ),
    .S1(net5884),
    .X(_03561_));
 sg13g2_mux4_1 _20353_ (.S0(net5940),
    .A0(\scanline[16][3] ),
    .A1(\scanline[17][3] ),
    .A2(\scanline[18][3] ),
    .A3(\scanline[19][3] ),
    .S1(net5884),
    .X(_03562_));
 sg13g2_mux4_1 _20354_ (.S0(net5939),
    .A0(\scanline[20][3] ),
    .A1(\scanline[21][3] ),
    .A2(\scanline[22][3] ),
    .A3(\scanline[23][3] ),
    .S1(net5883),
    .X(_03563_));
 sg13g2_a22oi_1 _20355_ (.Y(_03564_),
    .B1(_03563_),
    .B2(net5505),
    .A2(_03561_),
    .A1(net5533));
 sg13g2_a22oi_1 _20356_ (.Y(_03565_),
    .B1(_03562_),
    .B2(net5520),
    .A2(_03560_),
    .A1(net5489));
 sg13g2_a21oi_2 _20357_ (.B1(net5455),
    .Y(_03566_),
    .A2(_03565_),
    .A1(_03564_));
 sg13g2_mux4_1 _20358_ (.S0(net5935),
    .A0(\scanline[12][3] ),
    .A1(\scanline[13][3] ),
    .A2(\scanline[14][3] ),
    .A3(\scanline[15][3] ),
    .S1(net5878),
    .X(_03567_));
 sg13g2_mux4_1 _20359_ (.S0(net5933),
    .A0(\scanline[4][3] ),
    .A1(\scanline[5][3] ),
    .A2(\scanline[6][3] ),
    .A3(\scanline[7][3] ),
    .S1(net5876),
    .X(_03568_));
 sg13g2_mux4_1 _20360_ (.S0(net5935),
    .A0(\scanline[0][3] ),
    .A1(\scanline[1][3] ),
    .A2(\scanline[2][3] ),
    .A3(\scanline[3][3] ),
    .S1(net5878),
    .X(_03569_));
 sg13g2_mux4_1 _20361_ (.S0(net5933),
    .A0(\scanline[8][3] ),
    .A1(\scanline[9][3] ),
    .A2(\scanline[10][3] ),
    .A3(\scanline[11][3] ),
    .S1(net5876),
    .X(_03570_));
 sg13g2_a22oi_1 _20362_ (.Y(_03571_),
    .B1(_03570_),
    .B2(net5490),
    .A2(_03568_),
    .A1(net5504));
 sg13g2_a22oi_1 _20363_ (.Y(_03572_),
    .B1(_03569_),
    .B2(net5521),
    .A2(_03567_),
    .A1(net5532));
 sg13g2_a21oi_1 _20364_ (.A1(_03571_),
    .A2(_03572_),
    .Y(_03573_),
    .B1(net5510));
 sg13g2_or3_2 _20365_ (.A(net5841),
    .B(_03566_),
    .C(_03573_),
    .X(_03574_));
 sg13g2_a21oi_2 _20366_ (.B1(_03574_),
    .Y(_03575_),
    .A2(_03559_),
    .A1(_03551_));
 sg13g2_nand2b_1 _20367_ (.Y(_03576_),
    .B(\scanline[100][3] ),
    .A_N(net5957));
 sg13g2_a21oi_1 _20368_ (.A1(net5957),
    .A2(\scanline[101][3] ),
    .Y(_03577_),
    .B1(net5897));
 sg13g2_nand2_1 _20369_ (.Y(_03578_),
    .A(net5955),
    .B(\scanline[103][3] ));
 sg13g2_nand2b_1 _20370_ (.Y(_03579_),
    .B(\scanline[102][3] ),
    .A_N(net5955));
 sg13g2_nand3_1 _20371_ (.B(_03578_),
    .C(_03579_),
    .A(net5896),
    .Y(_03580_));
 sg13g2_a21oi_1 _20372_ (.A1(_03576_),
    .A2(_03577_),
    .Y(_03581_),
    .B1(net5499));
 sg13g2_mux4_1 _20373_ (.S0(net5952),
    .A0(\scanline[96][3] ),
    .A1(\scanline[97][3] ),
    .A2(\scanline[98][3] ),
    .A3(\scanline[99][3] ),
    .S1(net5893),
    .X(_03582_));
 sg13g2_mux4_1 _20374_ (.S0(net5957),
    .A0(\scanline[108][3] ),
    .A1(\scanline[109][3] ),
    .A2(\scanline[110][3] ),
    .A3(\scanline[111][3] ),
    .S1(net5897),
    .X(_03583_));
 sg13g2_mux4_1 _20375_ (.S0(net5956),
    .A0(\scanline[104][3] ),
    .A1(\scanline[105][3] ),
    .A2(\scanline[106][3] ),
    .A3(\scanline[107][3] ),
    .S1(net5897),
    .X(_03584_));
 sg13g2_a22oi_1 _20376_ (.Y(_03585_),
    .B1(_03584_),
    .B2(net5491),
    .A2(_03582_),
    .A1(net5523));
 sg13g2_a221oi_1 _20377_ (.B2(net5535),
    .C1(net5847),
    .B1(_03583_),
    .A1(_03580_),
    .Y(_03586_),
    .A2(_03581_));
 sg13g2_mux4_1 _20378_ (.S0(net5964),
    .A0(\scanline[116][3] ),
    .A1(\scanline[117][3] ),
    .A2(\scanline[118][3] ),
    .A3(\scanline[119][3] ),
    .S1(net5903),
    .X(_03587_));
 sg13g2_a21oi_1 _20379_ (.A1(net5507),
    .A2(_03587_),
    .Y(_03588_),
    .B1(net5555));
 sg13g2_mux4_1 _20380_ (.S0(net5966),
    .A0(\scanline[120][3] ),
    .A1(\scanline[121][3] ),
    .A2(\scanline[122][3] ),
    .A3(\scanline[123][3] ),
    .S1(net5904),
    .X(_03589_));
 sg13g2_and2_1 _20381_ (.A(net5491),
    .B(_03589_),
    .X(_03590_));
 sg13g2_mux4_1 _20382_ (.S0(net5961),
    .A0(\scanline[112][3] ),
    .A1(\scanline[113][3] ),
    .A2(\scanline[114][3] ),
    .A3(\scanline[115][3] ),
    .S1(net5900),
    .X(_03591_));
 sg13g2_mux4_1 _20383_ (.S0(net5961),
    .A0(\scanline[124][3] ),
    .A1(\scanline[125][3] ),
    .A2(\scanline[126][3] ),
    .A3(\scanline[127][3] ),
    .S1(net5900),
    .X(_03592_));
 sg13g2_a221oi_1 _20384_ (.B2(net5536),
    .C1(_03590_),
    .B1(_03592_),
    .A1(net5522),
    .Y(_03593_),
    .A2(_03591_));
 sg13g2_a221oi_1 _20385_ (.B2(_03593_),
    .C1(_08117_),
    .B1(_03588_),
    .A1(_03585_),
    .Y(_03594_),
    .A2(_03586_));
 sg13g2_mux4_1 _20386_ (.S0(net5943),
    .A0(\scanline[88][3] ),
    .A1(\scanline[89][3] ),
    .A2(\scanline[90][3] ),
    .A3(\scanline[91][3] ),
    .S1(net5889),
    .X(_03595_));
 sg13g2_mux4_1 _20387_ (.S0(net5944),
    .A0(\scanline[92][3] ),
    .A1(\scanline[93][3] ),
    .A2(\scanline[94][3] ),
    .A3(\scanline[95][3] ),
    .S1(net5887),
    .X(_03596_));
 sg13g2_a22oi_1 _20388_ (.Y(_03597_),
    .B1(_03596_),
    .B2(net5534),
    .A2(_03595_),
    .A1(net5492));
 sg13g2_mux4_1 _20389_ (.S0(net5945),
    .A0(\scanline[80][3] ),
    .A1(\scanline[81][3] ),
    .A2(\scanline[82][3] ),
    .A3(\scanline[83][3] ),
    .S1(net5888),
    .X(_03598_));
 sg13g2_mux4_1 _20390_ (.S0(net5943),
    .A0(\scanline[84][3] ),
    .A1(\scanline[85][3] ),
    .A2(\scanline[86][3] ),
    .A3(\scanline[87][3] ),
    .S1(net5886),
    .X(_03599_));
 sg13g2_a22oi_1 _20391_ (.Y(_03600_),
    .B1(_03599_),
    .B2(net5506),
    .A2(_03598_),
    .A1(net5522));
 sg13g2_a21oi_2 _20392_ (.B1(_03393_),
    .Y(_03601_),
    .A2(_03600_),
    .A1(_03597_));
 sg13g2_mux4_1 _20393_ (.S0(net5914),
    .A0(\scanline[64][3] ),
    .A1(\scanline[65][3] ),
    .A2(\scanline[66][3] ),
    .A3(\scanline[67][3] ),
    .S1(net5858),
    .X(_03602_));
 sg13g2_mux4_1 _20394_ (.S0(net5907),
    .A0(\scanline[72][3] ),
    .A1(\scanline[73][3] ),
    .A2(\scanline[74][3] ),
    .A3(\scanline[75][3] ),
    .S1(net5851),
    .X(_03603_));
 sg13g2_mux4_1 _20395_ (.S0(net5908),
    .A0(\scanline[76][3] ),
    .A1(\scanline[77][3] ),
    .A2(\scanline[78][3] ),
    .A3(\scanline[79][3] ),
    .S1(net5852),
    .X(_03604_));
 sg13g2_mux4_1 _20396_ (.S0(net5913),
    .A0(\scanline[68][3] ),
    .A1(\scanline[69][3] ),
    .A2(\scanline[70][3] ),
    .A3(\scanline[71][3] ),
    .S1(net5857),
    .X(_03605_));
 sg13g2_a22oi_1 _20397_ (.Y(_03606_),
    .B1(_03605_),
    .B2(net5500),
    .A2(_03603_),
    .A1(net5486));
 sg13g2_a22oi_1 _20398_ (.Y(_03607_),
    .B1(_03604_),
    .B2(net5529),
    .A2(_03602_),
    .A1(net5517));
 sg13g2_a21oi_2 _20399_ (.B1(net5509),
    .Y(_03608_),
    .A2(_03607_),
    .A1(_03606_));
 sg13g2_or3_1 _20400_ (.A(net5552),
    .B(_03601_),
    .C(_03608_),
    .X(_03609_));
 sg13g2_o21ai_1 _20401_ (.B1(_08120_),
    .Y(_03610_),
    .A1(_03594_),
    .A2(_03609_));
 sg13g2_mux4_1 _20402_ (.S0(net5923),
    .A0(\scanline[156][3] ),
    .A1(\scanline[157][3] ),
    .A2(\scanline[158][3] ),
    .A3(\scanline[159][3] ),
    .S1(net5868),
    .X(_03611_));
 sg13g2_o21ai_1 _20403_ (.B1(net5844),
    .Y(_03612_),
    .A1(net5527),
    .A2(_03611_));
 sg13g2_mux4_1 _20404_ (.S0(net5924),
    .A0(\scanline[148][3] ),
    .A1(\scanline[149][3] ),
    .A2(\scanline[150][3] ),
    .A3(\scanline[151][3] ),
    .S1(net5869),
    .X(_03613_));
 sg13g2_nor2_1 _20405_ (.A(net5497),
    .B(_03613_),
    .Y(_03614_));
 sg13g2_mux4_1 _20406_ (.S0(net5910),
    .A0(\scanline[144][3] ),
    .A1(\scanline[145][3] ),
    .A2(\scanline[146][3] ),
    .A3(\scanline[147][3] ),
    .S1(net5854),
    .X(_03615_));
 sg13g2_nor2_1 _20407_ (.A(net5515),
    .B(_03615_),
    .Y(_03616_));
 sg13g2_mux4_1 _20408_ (.S0(net5922),
    .A0(\scanline[152][3] ),
    .A1(\scanline[153][3] ),
    .A2(\scanline[154][3] ),
    .A3(\scanline[155][3] ),
    .S1(net5867),
    .X(_03617_));
 sg13g2_nor2_1 _20409_ (.A(net5485),
    .B(_03617_),
    .Y(_03618_));
 sg13g2_nor4_1 _20410_ (.A(_03612_),
    .B(_03614_),
    .C(_03616_),
    .D(_03618_),
    .Y(_03619_));
 sg13g2_mux4_1 _20411_ (.S0(net5909),
    .A0(\scanline[136][3] ),
    .A1(\scanline[137][3] ),
    .A2(\scanline[138][3] ),
    .A3(\scanline[139][3] ),
    .S1(net5853),
    .X(_03620_));
 sg13g2_nor2_1 _20412_ (.A(net5483),
    .B(_03620_),
    .Y(_03621_));
 sg13g2_mux4_1 _20413_ (.S0(net5911),
    .A0(\scanline[132][3] ),
    .A1(\scanline[133][3] ),
    .A2(\scanline[134][3] ),
    .A3(\scanline[135][3] ),
    .S1(net5855),
    .X(_03622_));
 sg13g2_nor2_1 _20414_ (.A(net5497),
    .B(_03622_),
    .Y(_03623_));
 sg13g2_mux4_1 _20415_ (.S0(net5909),
    .A0(\scanline[140][3] ),
    .A1(\scanline[141][3] ),
    .A2(\scanline[142][3] ),
    .A3(\scanline[143][3] ),
    .S1(net5853),
    .X(_03624_));
 sg13g2_o21ai_1 _20416_ (.B1(net5553),
    .Y(_03625_),
    .A1(net5525),
    .A2(_03624_));
 sg13g2_nor3_1 _20417_ (.A(_03621_),
    .B(_03623_),
    .C(_03625_),
    .Y(_03626_));
 sg13g2_nor2_1 _20418_ (.A(_03619_),
    .B(_03626_),
    .Y(_03627_));
 sg13g2_nand2b_1 _20419_ (.Y(_03628_),
    .B(net5918),
    .A_N(\scanline[129][3] ));
 sg13g2_o21ai_1 _20420_ (.B1(_03628_),
    .Y(_03629_),
    .A1(net5918),
    .A2(\scanline[128][3] ));
 sg13g2_mux2_1 _20421_ (.A0(\scanline[130][3] ),
    .A1(\scanline[131][3] ),
    .S(net5918),
    .X(_03630_));
 sg13g2_o21ai_1 _20422_ (.B1(_08694_),
    .Y(_03631_),
    .A1(net5864),
    .A2(_03629_));
 sg13g2_a21oi_1 _20423_ (.A1(net5864),
    .A2(_03630_),
    .Y(_03632_),
    .B1(_03631_));
 sg13g2_or3_1 _20424_ (.A(_08687_),
    .B(_03627_),
    .C(_03632_),
    .X(_03633_));
 sg13g2_o21ai_1 _20425_ (.B1(_03633_),
    .Y(_03634_),
    .A1(_03575_),
    .A2(_03610_));
 sg13g2_and2_1 _20426_ (.A(net5513),
    .B(_03634_),
    .X(_03635_));
 sg13g2_nand2_1 _20427_ (.Y(_03636_),
    .A(net5513),
    .B(_03634_));
 sg13g2_mux4_1 _20428_ (.S0(net5925),
    .A0(\scanline[152][2] ),
    .A1(\scanline[153][2] ),
    .A2(\scanline[154][2] ),
    .A3(\scanline[155][2] ),
    .S1(net5871),
    .X(_03637_));
 sg13g2_o21ai_1 _20429_ (.B1(net5844),
    .Y(_03638_),
    .A1(net5484),
    .A2(_03637_));
 sg13g2_mux4_1 _20430_ (.S0(net5924),
    .A0(\scanline[148][2] ),
    .A1(\scanline[149][2] ),
    .A2(\scanline[150][2] ),
    .A3(\scanline[151][2] ),
    .S1(net5869),
    .X(_03639_));
 sg13g2_nor2_1 _20431_ (.A(net5498),
    .B(_03639_),
    .Y(_03640_));
 sg13g2_mux4_1 _20432_ (.S0(net5918),
    .A0(\scanline[144][2] ),
    .A1(\scanline[145][2] ),
    .A2(\scanline[146][2] ),
    .A3(\scanline[147][2] ),
    .S1(net5864),
    .X(_03641_));
 sg13g2_nor2_1 _20433_ (.A(net5515),
    .B(_03641_),
    .Y(_03642_));
 sg13g2_mux4_1 _20434_ (.S0(net5922),
    .A0(\scanline[156][2] ),
    .A1(\scanline[157][2] ),
    .A2(\scanline[158][2] ),
    .A3(\scanline[159][2] ),
    .S1(net5866),
    .X(_03643_));
 sg13g2_nor2_1 _20435_ (.A(net5526),
    .B(_03643_),
    .Y(_03644_));
 sg13g2_nor4_1 _20436_ (.A(_03638_),
    .B(_03640_),
    .C(_03642_),
    .D(_03644_),
    .Y(_03645_));
 sg13g2_mux4_1 _20437_ (.S0(net5909),
    .A0(\scanline[136][2] ),
    .A1(\scanline[137][2] ),
    .A2(\scanline[138][2] ),
    .A3(\scanline[139][2] ),
    .S1(net5853),
    .X(_03646_));
 sg13g2_o21ai_1 _20438_ (.B1(net5553),
    .Y(_03647_),
    .A1(net5483),
    .A2(_03646_));
 sg13g2_mux4_1 _20439_ (.S0(net5910),
    .A0(\scanline[132][2] ),
    .A1(\scanline[133][2] ),
    .A2(\scanline[134][2] ),
    .A3(\scanline[135][2] ),
    .S1(net5854),
    .X(_03648_));
 sg13g2_nor2_1 _20440_ (.A(net5497),
    .B(_03648_),
    .Y(_03649_));
 sg13g2_mux4_1 _20441_ (.S0(net5923),
    .A0(\scanline[140][2] ),
    .A1(\scanline[141][2] ),
    .A2(\scanline[142][2] ),
    .A3(\scanline[143][2] ),
    .S1(net5868),
    .X(_03650_));
 sg13g2_nor2_1 _20442_ (.A(net5525),
    .B(_03650_),
    .Y(_03651_));
 sg13g2_mux4_1 _20443_ (.S0(net5921),
    .A0(\scanline[128][2] ),
    .A1(\scanline[129][2] ),
    .A2(\scanline[130][2] ),
    .A3(\scanline[131][2] ),
    .S1(net5864),
    .X(_03652_));
 sg13g2_nor2_1 _20444_ (.A(net5514),
    .B(_03652_),
    .Y(_03653_));
 sg13g2_nor4_2 _20445_ (.A(_03647_),
    .B(_03649_),
    .C(_03651_),
    .Y(_03654_),
    .D(_03653_));
 sg13g2_o21ai_1 _20446_ (.B1(_08686_),
    .Y(_03655_),
    .A1(_03645_),
    .A2(_03654_));
 sg13g2_mux4_1 _20447_ (.S0(net5966),
    .A0(\scanline[120][2] ),
    .A1(\scanline[121][2] ),
    .A2(\scanline[122][2] ),
    .A3(\scanline[123][2] ),
    .S1(net5904),
    .X(_03656_));
 sg13g2_and2_1 _20448_ (.A(net5491),
    .B(_03656_),
    .X(_03657_));
 sg13g2_mux4_1 _20449_ (.S0(net5966),
    .A0(\scanline[112][2] ),
    .A1(\scanline[113][2] ),
    .A2(\scanline[114][2] ),
    .A3(\scanline[115][2] ),
    .S1(net5904),
    .X(_03658_));
 sg13g2_nand2b_1 _20450_ (.Y(_03659_),
    .B(\scanline[124][2] ),
    .A_N(net5959));
 sg13g2_a21oi_1 _20451_ (.A1(net5959),
    .A2(\scanline[125][2] ),
    .Y(_03660_),
    .B1(net5899));
 sg13g2_nand2_1 _20452_ (.Y(_03661_),
    .A(net5959),
    .B(\scanline[127][2] ));
 sg13g2_nand2b_1 _20453_ (.Y(_03662_),
    .B(\scanline[126][2] ),
    .A_N(net5960));
 sg13g2_nand3_1 _20454_ (.B(_03661_),
    .C(_03662_),
    .A(net5899),
    .Y(_03663_));
 sg13g2_a21oi_1 _20455_ (.A1(_03659_),
    .A2(_03660_),
    .Y(_03664_),
    .B1(net5528));
 sg13g2_mux4_1 _20456_ (.S0(net5965),
    .A0(\scanline[116][2] ),
    .A1(\scanline[117][2] ),
    .A2(\scanline[118][2] ),
    .A3(\scanline[119][2] ),
    .S1(net5903),
    .X(_03665_));
 sg13g2_a21oi_1 _20457_ (.A1(_03663_),
    .A2(_03664_),
    .Y(_03666_),
    .B1(net5555));
 sg13g2_a221oi_1 _20458_ (.B2(net5506),
    .C1(_03657_),
    .B1(_03665_),
    .A1(net5524),
    .Y(_03667_),
    .A2(_03658_));
 sg13g2_nand2b_1 _20459_ (.Y(_03668_),
    .B(\scanline[108][2] ),
    .A_N(net5953));
 sg13g2_a21oi_1 _20460_ (.A1(net5953),
    .A2(\scanline[109][2] ),
    .Y(_03669_),
    .B1(net5895));
 sg13g2_nand2_1 _20461_ (.Y(_03670_),
    .A(net5954),
    .B(\scanline[111][2] ));
 sg13g2_nand2b_1 _20462_ (.Y(_03671_),
    .B(\scanline[110][2] ),
    .A_N(net5953));
 sg13g2_nand3_1 _20463_ (.B(_03670_),
    .C(_03671_),
    .A(net5898),
    .Y(_03672_));
 sg13g2_a21oi_1 _20464_ (.A1(_03668_),
    .A2(_03669_),
    .Y(_03673_),
    .B1(net5528));
 sg13g2_mux4_1 _20465_ (.S0(net5952),
    .A0(\scanline[96][2] ),
    .A1(\scanline[97][2] ),
    .A2(\scanline[98][2] ),
    .A3(\scanline[99][2] ),
    .S1(net5892),
    .X(_03674_));
 sg13g2_mux4_1 _20466_ (.S0(net5953),
    .A0(\scanline[100][2] ),
    .A1(\scanline[101][2] ),
    .A2(\scanline[102][2] ),
    .A3(\scanline[103][2] ),
    .S1(net5895),
    .X(_03675_));
 sg13g2_mux4_1 _20467_ (.S0(net5955),
    .A0(\scanline[104][2] ),
    .A1(\scanline[105][2] ),
    .A2(\scanline[106][2] ),
    .A3(\scanline[107][2] ),
    .S1(net5896),
    .X(_03676_));
 sg13g2_a22oi_1 _20468_ (.Y(_03677_),
    .B1(_03676_),
    .B2(net5491),
    .A2(_03674_),
    .A1(net5523));
 sg13g2_a221oi_1 _20469_ (.B2(net5502),
    .C1(net5847),
    .B1(_03675_),
    .A1(_03672_),
    .Y(_03678_),
    .A2(_03673_));
 sg13g2_a22oi_1 _20470_ (.Y(_03679_),
    .B1(_03677_),
    .B2(_03678_),
    .A2(_03667_),
    .A1(_03666_));
 sg13g2_mux4_1 _20471_ (.S0(net5943),
    .A0(\scanline[88][2] ),
    .A1(\scanline[89][2] ),
    .A2(\scanline[90][2] ),
    .A3(\scanline[91][2] ),
    .S1(net5886),
    .X(_03680_));
 sg13g2_mux4_1 _20472_ (.S0(net5945),
    .A0(\scanline[80][2] ),
    .A1(\scanline[81][2] ),
    .A2(\scanline[82][2] ),
    .A3(\scanline[83][2] ),
    .S1(net5888),
    .X(_03681_));
 sg13g2_a22oi_1 _20473_ (.Y(_03682_),
    .B1(_03681_),
    .B2(net5520),
    .A2(_03680_),
    .A1(net5489));
 sg13g2_mux4_1 _20474_ (.S0(net5960),
    .A0(\scanline[92][2] ),
    .A1(\scanline[93][2] ),
    .A2(\scanline[94][2] ),
    .A3(\scanline[95][2] ),
    .S1(net5899),
    .X(_03683_));
 sg13g2_mux4_1 _20475_ (.S0(net5960),
    .A0(\scanline[84][2] ),
    .A1(\scanline[85][2] ),
    .A2(\scanline[86][2] ),
    .A3(\scanline[87][2] ),
    .S1(net5899),
    .X(_03684_));
 sg13g2_a22oi_1 _20476_ (.Y(_03685_),
    .B1(_03684_),
    .B2(net5506),
    .A2(_03683_),
    .A1(net5534));
 sg13g2_nand2_2 _20477_ (.Y(_03686_),
    .A(_03682_),
    .B(_03685_));
 sg13g2_mux4_1 _20478_ (.S0(net5914),
    .A0(\scanline[64][2] ),
    .A1(\scanline[65][2] ),
    .A2(\scanline[66][2] ),
    .A3(\scanline[67][2] ),
    .S1(net5858),
    .X(_03687_));
 sg13g2_mux4_1 _20479_ (.S0(net5913),
    .A0(\scanline[68][2] ),
    .A1(\scanline[69][2] ),
    .A2(\scanline[70][2] ),
    .A3(\scanline[71][2] ),
    .S1(net5857),
    .X(_03688_));
 sg13g2_mux4_1 _20480_ (.S0(net5907),
    .A0(\scanline[72][2] ),
    .A1(\scanline[73][2] ),
    .A2(\scanline[74][2] ),
    .A3(\scanline[75][2] ),
    .S1(net5851),
    .X(_03689_));
 sg13g2_mux4_1 _20481_ (.S0(net5908),
    .A0(\scanline[76][2] ),
    .A1(\scanline[77][2] ),
    .A2(\scanline[78][2] ),
    .A3(\scanline[79][2] ),
    .S1(net5852),
    .X(_03690_));
 sg13g2_a22oi_1 _20482_ (.Y(_03691_),
    .B1(_03690_),
    .B2(net5529),
    .A2(_03688_),
    .A1(net5500));
 sg13g2_a22oi_1 _20483_ (.Y(_03692_),
    .B1(_03689_),
    .B2(net5486),
    .A2(_03687_),
    .A1(net5517));
 sg13g2_a21oi_2 _20484_ (.B1(net5509),
    .Y(_03693_),
    .A2(_03692_),
    .A1(_03691_));
 sg13g2_nand2b_1 _20485_ (.Y(_03694_),
    .B(net5840),
    .A_N(_03693_));
 sg13g2_a221oi_1 _20486_ (.B2(_03392_),
    .C1(_03694_),
    .B1(_03686_),
    .A1(\hvsync_gen.hpos[7] ),
    .Y(_03695_),
    .A2(_03679_));
 sg13g2_mux4_1 _20487_ (.S0(net5953),
    .A0(\scanline[52][2] ),
    .A1(\scanline[53][2] ),
    .A2(\scanline[54][2] ),
    .A3(\scanline[55][2] ),
    .S1(net5895),
    .X(_03696_));
 sg13g2_mux4_1 _20488_ (.S0(net5920),
    .A0(\scanline[56][2] ),
    .A1(\scanline[57][2] ),
    .A2(\scanline[58][2] ),
    .A3(\scanline[59][2] ),
    .S1(net5862),
    .X(_03697_));
 sg13g2_mux4_1 _20489_ (.S0(net5926),
    .A0(\scanline[48][2] ),
    .A1(\scanline[49][2] ),
    .A2(\scanline[50][2] ),
    .A3(\scanline[51][2] ),
    .S1(net5870),
    .X(_03698_));
 sg13g2_nand2b_1 _20490_ (.Y(_03699_),
    .B(\scanline[60][2] ),
    .A_N(net5948));
 sg13g2_a21oi_1 _20491_ (.A1(net5948),
    .A2(\scanline[61][2] ),
    .Y(_03700_),
    .B1(net5891));
 sg13g2_nand2_1 _20492_ (.Y(_03701_),
    .A(net5948),
    .B(\scanline[63][2] ));
 sg13g2_nand2b_1 _20493_ (.Y(_03702_),
    .B(\scanline[62][2] ),
    .A_N(net5948));
 sg13g2_nand3_1 _20494_ (.B(_03701_),
    .C(_03702_),
    .A(net5890),
    .Y(_03703_));
 sg13g2_a21oi_1 _20495_ (.A1(_03699_),
    .A2(_03700_),
    .Y(_03704_),
    .B1(net5528));
 sg13g2_a22oi_1 _20496_ (.Y(_03705_),
    .B1(_03698_),
    .B2(net5519),
    .A2(_03697_),
    .A1(net5488));
 sg13g2_a221oi_1 _20497_ (.B2(_03704_),
    .C1(net5554),
    .B1(_03703_),
    .A1(net5502),
    .Y(_03706_),
    .A2(_03696_));
 sg13g2_mux4_1 _20498_ (.S0(net5932),
    .A0(\scanline[36][2] ),
    .A1(\scanline[37][2] ),
    .A2(\scanline[38][2] ),
    .A3(\scanline[39][2] ),
    .S1(net5877),
    .X(_03707_));
 sg13g2_a21oi_1 _20499_ (.A1(net5501),
    .A2(_03707_),
    .Y(_03708_),
    .B1(net5847));
 sg13g2_mux4_1 _20500_ (.S0(net5919),
    .A0(\scanline[32][2] ),
    .A1(\scanline[33][2] ),
    .A2(\scanline[34][2] ),
    .A3(\scanline[35][2] ),
    .S1(net5862),
    .X(_03709_));
 sg13g2_mux4_1 _20501_ (.S0(net5919),
    .A0(\scanline[44][2] ),
    .A1(\scanline[45][2] ),
    .A2(\scanline[46][2] ),
    .A3(\scanline[47][2] ),
    .S1(net5862),
    .X(_03710_));
 sg13g2_and2_1 _20502_ (.A(net5530),
    .B(_03710_),
    .X(_03711_));
 sg13g2_mux4_1 _20503_ (.S0(net5916),
    .A0(\scanline[40][2] ),
    .A1(\scanline[41][2] ),
    .A2(\scanline[42][2] ),
    .A3(\scanline[43][2] ),
    .S1(net5859),
    .X(_03712_));
 sg13g2_a221oi_1 _20504_ (.B2(net5487),
    .C1(_03711_),
    .B1(_03712_),
    .A1(net5518),
    .Y(_03713_),
    .A2(_03709_));
 sg13g2_a221oi_1 _20505_ (.B2(_03713_),
    .C1(_08117_),
    .B1(_03708_),
    .A1(_03705_),
    .Y(_03714_),
    .A2(_03706_));
 sg13g2_mux4_1 _20506_ (.S0(net5938),
    .A0(\scanline[24][2] ),
    .A1(\scanline[25][2] ),
    .A2(\scanline[26][2] ),
    .A3(\scanline[27][2] ),
    .S1(net5882),
    .X(_03715_));
 sg13g2_mux4_1 _20507_ (.S0(net5939),
    .A0(\scanline[16][2] ),
    .A1(\scanline[17][2] ),
    .A2(\scanline[18][2] ),
    .A3(\scanline[19][2] ),
    .S1(net5883),
    .X(_03716_));
 sg13g2_mux4_1 _20508_ (.S0(net5938),
    .A0(\scanline[28][2] ),
    .A1(\scanline[29][2] ),
    .A2(\scanline[30][2] ),
    .A3(\scanline[31][2] ),
    .S1(net5882),
    .X(_03717_));
 sg13g2_mux4_1 _20509_ (.S0(net5939),
    .A0(\scanline[20][2] ),
    .A1(\scanline[21][2] ),
    .A2(\scanline[22][2] ),
    .A3(\scanline[23][2] ),
    .S1(net5883),
    .X(_03718_));
 sg13g2_a22oi_1 _20510_ (.Y(_03719_),
    .B1(_03718_),
    .B2(net5505),
    .A2(_03716_),
    .A1(net5520));
 sg13g2_a22oi_1 _20511_ (.Y(_03720_),
    .B1(_03717_),
    .B2(net5532),
    .A2(_03715_),
    .A1(net5489));
 sg13g2_a21oi_2 _20512_ (.B1(net5455),
    .Y(_03721_),
    .A2(_03720_),
    .A1(_03719_));
 sg13g2_mux4_1 _20513_ (.S0(net5933),
    .A0(\scanline[4][2] ),
    .A1(\scanline[5][2] ),
    .A2(\scanline[6][2] ),
    .A3(\scanline[7][2] ),
    .S1(net5876),
    .X(_03722_));
 sg13g2_mux4_1 _20514_ (.S0(net5935),
    .A0(\scanline[12][2] ),
    .A1(\scanline[13][2] ),
    .A2(\scanline[14][2] ),
    .A3(\scanline[15][2] ),
    .S1(net5879),
    .X(_03723_));
 sg13g2_mux4_1 _20515_ (.S0(net5931),
    .A0(\scanline[8][2] ),
    .A1(\scanline[9][2] ),
    .A2(\scanline[10][2] ),
    .A3(\scanline[11][2] ),
    .S1(net5875),
    .X(_03724_));
 sg13g2_mux4_1 _20516_ (.S0(net5935),
    .A0(\scanline[0][2] ),
    .A1(\scanline[1][2] ),
    .A2(\scanline[2][2] ),
    .A3(\scanline[3][2] ),
    .S1(net5879),
    .X(_03725_));
 sg13g2_a22oi_1 _20517_ (.Y(_03726_),
    .B1(_03725_),
    .B2(net5521),
    .A2(_03723_),
    .A1(net5532));
 sg13g2_a22oi_1 _20518_ (.Y(_03727_),
    .B1(_03724_),
    .B2(net5490),
    .A2(_03722_),
    .A1(net5504));
 sg13g2_a21oi_1 _20519_ (.A1(_03726_),
    .A2(_03727_),
    .Y(_03728_),
    .B1(net5510));
 sg13g2_or3_2 _20520_ (.A(net5841),
    .B(_03721_),
    .C(_03728_),
    .X(_03729_));
 sg13g2_o21ai_1 _20521_ (.B1(_08120_),
    .Y(_03730_),
    .A1(_03714_),
    .A2(_03729_));
 sg13g2_o21ai_1 _20522_ (.B1(_03655_),
    .Y(_03731_),
    .A1(_03695_),
    .A2(_03730_));
 sg13g2_and2_2 _20523_ (.A(net5512),
    .B(net5360),
    .X(_03732_));
 sg13g2_nand2_2 _20524_ (.Y(_03733_),
    .A(net5513),
    .B(_03731_));
 sg13g2_mux4_1 _20525_ (.S0(net5924),
    .A0(\scanline[148][1] ),
    .A1(\scanline[149][1] ),
    .A2(\scanline[150][1] ),
    .A3(\scanline[151][1] ),
    .S1(net5869),
    .X(_03734_));
 sg13g2_nor2_1 _20526_ (.A(net5498),
    .B(_03734_),
    .Y(_03735_));
 sg13g2_mux4_1 _20527_ (.S0(net5923),
    .A0(\scanline[156][1] ),
    .A1(\scanline[157][1] ),
    .A2(\scanline[158][1] ),
    .A3(\scanline[159][1] ),
    .S1(net5867),
    .X(_03736_));
 sg13g2_nor2_1 _20528_ (.A(net5527),
    .B(_03736_),
    .Y(_03737_));
 sg13g2_mux4_1 _20529_ (.S0(net5922),
    .A0(\scanline[144][1] ),
    .A1(\scanline[145][1] ),
    .A2(\scanline[146][1] ),
    .A3(\scanline[147][1] ),
    .S1(net5866),
    .X(_03738_));
 sg13g2_nor2_1 _20530_ (.A(net5515),
    .B(_03738_),
    .Y(_03739_));
 sg13g2_mux4_1 _20531_ (.S0(net5922),
    .A0(\scanline[152][1] ),
    .A1(\scanline[153][1] ),
    .A2(\scanline[154][1] ),
    .A3(\scanline[155][1] ),
    .S1(net5866),
    .X(_03740_));
 sg13g2_nor2_1 _20532_ (.A(net5485),
    .B(_03740_),
    .Y(_03741_));
 sg13g2_mux4_1 _20533_ (.S0(net5911),
    .A0(\scanline[132][1] ),
    .A1(\scanline[133][1] ),
    .A2(\scanline[134][1] ),
    .A3(\scanline[135][1] ),
    .S1(net5855),
    .X(_03742_));
 sg13g2_mux4_1 _20534_ (.S0(net5910),
    .A0(\scanline[140][1] ),
    .A1(\scanline[141][1] ),
    .A2(\scanline[142][1] ),
    .A3(\scanline[143][1] ),
    .S1(net5854),
    .X(_03743_));
 sg13g2_nor2_1 _20535_ (.A(net5525),
    .B(_03743_),
    .Y(_03744_));
 sg13g2_mux4_1 _20536_ (.S0(net5908),
    .A0(\scanline[136][1] ),
    .A1(\scanline[137][1] ),
    .A2(\scanline[138][1] ),
    .A3(\scanline[139][1] ),
    .S1(net5852),
    .X(_03745_));
 sg13g2_nor2_1 _20537_ (.A(net5483),
    .B(_03745_),
    .Y(_03746_));
 sg13g2_mux4_1 _20538_ (.S0(net5910),
    .A0(\scanline[128][1] ),
    .A1(\scanline[129][1] ),
    .A2(\scanline[130][1] ),
    .A3(\scanline[131][1] ),
    .S1(net5854),
    .X(_03747_));
 sg13g2_nor2_1 _20539_ (.A(net5514),
    .B(_03747_),
    .Y(_03748_));
 sg13g2_nor3_1 _20540_ (.A(_03744_),
    .B(_03746_),
    .C(_03748_),
    .Y(_03749_));
 sg13g2_o21ai_1 _20541_ (.B1(_03749_),
    .Y(_03750_),
    .A1(net5497),
    .A2(_03742_));
 sg13g2_nor4_1 _20542_ (.A(_03735_),
    .B(_03737_),
    .C(_03739_),
    .D(_03741_),
    .Y(_03751_));
 sg13g2_o21ai_1 _20543_ (.B1(_08686_),
    .Y(_03752_),
    .A1(net5553),
    .A2(_03751_));
 sg13g2_a21oi_2 _20544_ (.B1(_03752_),
    .Y(_03753_),
    .A2(_03750_),
    .A1(net5553));
 sg13g2_mux4_1 _20545_ (.S0(net5927),
    .A0(\scanline[48][1] ),
    .A1(\scanline[49][1] ),
    .A2(\scanline[50][1] ),
    .A3(\scanline[51][1] ),
    .S1(net5872),
    .X(_03754_));
 sg13g2_nand2_1 _20546_ (.Y(_03755_),
    .A(net5950),
    .B(\scanline[63][1] ));
 sg13g2_nand2b_1 _20547_ (.Y(_03756_),
    .B(\scanline[62][1] ),
    .A_N(net5950));
 sg13g2_nand3_1 _20548_ (.B(_03755_),
    .C(_03756_),
    .A(net5890),
    .Y(_03757_));
 sg13g2_nand2b_1 _20549_ (.Y(_03758_),
    .B(\scanline[60][1] ),
    .A_N(net5950));
 sg13g2_a21oi_1 _20550_ (.A1(net5950),
    .A2(\scanline[61][1] ),
    .Y(_03759_),
    .B1(net5890));
 sg13g2_a21oi_1 _20551_ (.A1(_03758_),
    .A2(_03759_),
    .Y(_03760_),
    .B1(net5528));
 sg13g2_mux4_1 _20552_ (.S0(net5926),
    .A0(\scanline[56][1] ),
    .A1(\scanline[57][1] ),
    .A2(\scanline[58][1] ),
    .A3(\scanline[59][1] ),
    .S1(net5870),
    .X(_03761_));
 sg13g2_and2_1 _20553_ (.A(net5488),
    .B(_03761_),
    .X(_03762_));
 sg13g2_mux4_1 _20554_ (.S0(net5929),
    .A0(\scanline[52][1] ),
    .A1(\scanline[53][1] ),
    .A2(\scanline[54][1] ),
    .A3(\scanline[55][1] ),
    .S1(net5873),
    .X(_03763_));
 sg13g2_a221oi_1 _20555_ (.B2(_03760_),
    .C1(_03762_),
    .B1(_03757_),
    .A1(net5519),
    .Y(_03764_),
    .A2(_03754_));
 sg13g2_a21oi_1 _20556_ (.A1(net5502),
    .A2(_03763_),
    .Y(_03765_),
    .B1(net5553));
 sg13g2_mux4_1 _20557_ (.S0(net5920),
    .A0(\scanline[44][1] ),
    .A1(\scanline[45][1] ),
    .A2(\scanline[46][1] ),
    .A3(\scanline[47][1] ),
    .S1(net5863),
    .X(_03766_));
 sg13g2_mux4_1 _20558_ (.S0(net5916),
    .A0(\scanline[40][1] ),
    .A1(\scanline[41][1] ),
    .A2(\scanline[42][1] ),
    .A3(\scanline[43][1] ),
    .S1(net5860),
    .X(_03767_));
 sg13g2_mux4_1 _20559_ (.S0(net5915),
    .A0(\scanline[36][1] ),
    .A1(\scanline[37][1] ),
    .A2(\scanline[38][1] ),
    .A3(\scanline[39][1] ),
    .S1(net5859),
    .X(_03768_));
 sg13g2_nand2_1 _20560_ (.Y(_03769_),
    .A(net5920),
    .B(\scanline[35][1] ));
 sg13g2_nand2b_1 _20561_ (.Y(_03770_),
    .B(\scanline[34][1] ),
    .A_N(net5920));
 sg13g2_nand3_1 _20562_ (.B(_03769_),
    .C(_03770_),
    .A(net5863),
    .Y(_03771_));
 sg13g2_nand2b_1 _20563_ (.Y(_03772_),
    .B(\scanline[32][1] ),
    .A_N(net5919));
 sg13g2_a21oi_1 _20564_ (.A1(net5920),
    .A2(\scanline[33][1] ),
    .Y(_03773_),
    .B1(net5863));
 sg13g2_a21oi_1 _20565_ (.A1(_03772_),
    .A2(_03773_),
    .Y(_03774_),
    .B1(net5516));
 sg13g2_a22oi_1 _20566_ (.Y(_03775_),
    .B1(_03768_),
    .B2(net5500),
    .A2(_03766_),
    .A1(net5530));
 sg13g2_a221oi_1 _20567_ (.B2(_03774_),
    .C1(net5845),
    .B1(_03771_),
    .A1(net5486),
    .Y(_03776_),
    .A2(_03767_));
 sg13g2_a221oi_1 _20568_ (.B2(_03776_),
    .C1(net5840),
    .B1(_03775_),
    .A1(_03764_),
    .Y(_03777_),
    .A2(_03765_));
 sg13g2_mux4_1 _20569_ (.S0(net5955),
    .A0(\scanline[104][1] ),
    .A1(\scanline[105][1] ),
    .A2(\scanline[106][1] ),
    .A3(\scanline[107][1] ),
    .S1(net5897),
    .X(_03778_));
 sg13g2_mux4_1 _20570_ (.S0(net5952),
    .A0(\scanline[96][1] ),
    .A1(\scanline[97][1] ),
    .A2(\scanline[98][1] ),
    .A3(\scanline[99][1] ),
    .S1(net5892),
    .X(_03779_));
 sg13g2_mux4_1 _20571_ (.S0(net5957),
    .A0(\scanline[100][1] ),
    .A1(\scanline[101][1] ),
    .A2(\scanline[102][1] ),
    .A3(\scanline[103][1] ),
    .S1(net5897),
    .X(_03780_));
 sg13g2_mux4_1 _20572_ (.S0(net5953),
    .A0(\scanline[108][1] ),
    .A1(\scanline[109][1] ),
    .A2(\scanline[110][1] ),
    .A3(\scanline[111][1] ),
    .S1(net5895),
    .X(_03781_));
 sg13g2_a22oi_1 _20573_ (.Y(_03782_),
    .B1(_03781_),
    .B2(net5535),
    .A2(_03778_),
    .A1(net5493));
 sg13g2_a221oi_1 _20574_ (.B2(net5507),
    .C1(net5848),
    .B1(_03780_),
    .A1(net5523),
    .Y(_03783_),
    .A2(_03779_));
 sg13g2_mux4_1 _20575_ (.S0(net5964),
    .A0(\scanline[120][1] ),
    .A1(\scanline[121][1] ),
    .A2(\scanline[122][1] ),
    .A3(\scanline[123][1] ),
    .S1(net5903),
    .X(_03784_));
 sg13g2_a21o_1 _20576_ (.A2(_03784_),
    .A1(net5491),
    .B1(net5554),
    .X(_03785_));
 sg13g2_nand2_1 _20577_ (.Y(_03786_),
    .A(net5959),
    .B(\scanline[127][1] ));
 sg13g2_nand2b_1 _20578_ (.Y(_03787_),
    .B(\scanline[126][1] ),
    .A_N(net5959));
 sg13g2_and3_1 _20579_ (.X(_03788_),
    .A(net5902),
    .B(_03786_),
    .C(_03787_));
 sg13g2_mux2_1 _20580_ (.A0(\scanline[124][1] ),
    .A1(\scanline[125][1] ),
    .S(net5959),
    .X(_03789_));
 sg13g2_o21ai_1 _20581_ (.B1(net5535),
    .Y(_03790_),
    .A1(net5899),
    .A2(_03789_));
 sg13g2_mux4_1 _20582_ (.S0(net5961),
    .A0(\scanline[112][1] ),
    .A1(\scanline[113][1] ),
    .A2(\scanline[114][1] ),
    .A3(\scanline[115][1] ),
    .S1(net5901),
    .X(_03791_));
 sg13g2_mux4_1 _20583_ (.S0(net5964),
    .A0(\scanline[116][1] ),
    .A1(\scanline[117][1] ),
    .A2(\scanline[118][1] ),
    .A3(\scanline[119][1] ),
    .S1(net5904),
    .X(_03792_));
 sg13g2_a22oi_1 _20584_ (.Y(_03793_),
    .B1(_03792_),
    .B2(net5506),
    .A2(_03791_),
    .A1(net5524));
 sg13g2_o21ai_1 _20585_ (.B1(_03793_),
    .Y(_03794_),
    .A1(_03788_),
    .A2(_03790_));
 sg13g2_a21oi_1 _20586_ (.A1(_03782_),
    .A2(_03783_),
    .Y(_03795_),
    .B1(_08119_));
 sg13g2_o21ai_1 _20587_ (.B1(_03795_),
    .Y(_03796_),
    .A1(_03785_),
    .A2(_03794_));
 sg13g2_nand3b_1 _20588_ (.B(_03796_),
    .C(net5843),
    .Y(_03797_),
    .A_N(_03777_));
 sg13g2_mux4_1 _20589_ (.S0(net5937),
    .A0(\scanline[0][1] ),
    .A1(\scanline[1][1] ),
    .A2(\scanline[2][1] ),
    .A3(\scanline[3][1] ),
    .S1(net5879),
    .X(_03798_));
 sg13g2_mux4_1 _20590_ (.S0(net5937),
    .A0(\scanline[12][1] ),
    .A1(\scanline[13][1] ),
    .A2(\scanline[14][1] ),
    .A3(\scanline[15][1] ),
    .S1(net5879),
    .X(_03799_));
 sg13g2_a22oi_1 _20591_ (.Y(_03800_),
    .B1(_03799_),
    .B2(net5535),
    .A2(_03798_),
    .A1(net5523));
 sg13g2_mux4_1 _20592_ (.S0(net5933),
    .A0(\scanline[4][1] ),
    .A1(\scanline[5][1] ),
    .A2(\scanline[6][1] ),
    .A3(\scanline[7][1] ),
    .S1(net5876),
    .X(_03801_));
 sg13g2_mux4_1 _20593_ (.S0(net5931),
    .A0(\scanline[8][1] ),
    .A1(\scanline[9][1] ),
    .A2(\scanline[10][1] ),
    .A3(\scanline[11][1] ),
    .S1(net5875),
    .X(_03802_));
 sg13g2_a22oi_1 _20594_ (.Y(_03803_),
    .B1(_03802_),
    .B2(net5490),
    .A2(_03801_),
    .A1(net5504));
 sg13g2_a21oi_1 _20595_ (.A1(_03800_),
    .A2(_03803_),
    .Y(_03804_),
    .B1(net5847));
 sg13g2_mux4_1 _20596_ (.S0(net5944),
    .A0(\scanline[28][1] ),
    .A1(\scanline[29][1] ),
    .A2(\scanline[30][1] ),
    .A3(\scanline[31][1] ),
    .S1(net5887),
    .X(_03805_));
 sg13g2_mux4_1 _20597_ (.S0(net5944),
    .A0(\scanline[16][1] ),
    .A1(\scanline[17][1] ),
    .A2(\scanline[18][1] ),
    .A3(\scanline[19][1] ),
    .S1(net5887),
    .X(_03806_));
 sg13g2_a22oi_1 _20598_ (.Y(_03807_),
    .B1(_03806_),
    .B2(net5521),
    .A2(_03805_),
    .A1(net5533));
 sg13g2_mux4_1 _20599_ (.S0(net5938),
    .A0(\scanline[24][1] ),
    .A1(\scanline[25][1] ),
    .A2(\scanline[26][1] ),
    .A3(\scanline[27][1] ),
    .S1(net5882),
    .X(_03808_));
 sg13g2_mux4_1 _20600_ (.S0(net5938),
    .A0(\scanline[20][1] ),
    .A1(\scanline[21][1] ),
    .A2(\scanline[22][1] ),
    .A3(\scanline[23][1] ),
    .S1(net5882),
    .X(_03809_));
 sg13g2_a22oi_1 _20601_ (.Y(_03810_),
    .B1(_03809_),
    .B2(net5504),
    .A2(_03808_),
    .A1(net5489));
 sg13g2_a21oi_2 _20602_ (.B1(net5555),
    .Y(_03811_),
    .A2(_03810_),
    .A1(_03807_));
 sg13g2_nor4_2 _20603_ (.A(net5842),
    .B(net5841),
    .C(_03804_),
    .Y(_03812_),
    .D(_03811_));
 sg13g2_mux4_1 _20604_ (.S0(net5918),
    .A0(\scanline[64][1] ),
    .A1(\scanline[65][1] ),
    .A2(\scanline[66][1] ),
    .A3(\scanline[67][1] ),
    .S1(net5864),
    .X(_03813_));
 sg13g2_mux4_1 _20605_ (.S0(net5908),
    .A0(\scanline[76][1] ),
    .A1(\scanline[77][1] ),
    .A2(\scanline[78][1] ),
    .A3(\scanline[79][1] ),
    .S1(net5852),
    .X(_03814_));
 sg13g2_mux4_1 _20606_ (.S0(net5907),
    .A0(\scanline[72][1] ),
    .A1(\scanline[73][1] ),
    .A2(\scanline[74][1] ),
    .A3(\scanline[75][1] ),
    .S1(net5851),
    .X(_03815_));
 sg13g2_mux4_1 _20607_ (.S0(net5913),
    .A0(\scanline[68][1] ),
    .A1(\scanline[69][1] ),
    .A2(\scanline[70][1] ),
    .A3(\scanline[71][1] ),
    .S1(net5857),
    .X(_03816_));
 sg13g2_a22oi_1 _20608_ (.Y(_03817_),
    .B1(_03816_),
    .B2(net5500),
    .A2(_03814_),
    .A1(net5529));
 sg13g2_a221oi_1 _20609_ (.B2(net5486),
    .C1(_03226_),
    .B1(_03815_),
    .A1(net5517),
    .Y(_03818_),
    .A2(_03813_));
 sg13g2_and2_1 _20610_ (.A(_03817_),
    .B(_03818_),
    .X(_03819_));
 sg13g2_nor2b_1 _20611_ (.A(net5942),
    .B_N(\scanline[90][1] ),
    .Y(_03820_));
 sg13g2_a21oi_1 _20612_ (.A1(net5942),
    .A2(\scanline[91][1] ),
    .Y(_03821_),
    .B1(_03820_));
 sg13g2_nand2b_1 _20613_ (.Y(_03822_),
    .B(\scanline[88][1] ),
    .A_N(net5942));
 sg13g2_a21oi_1 _20614_ (.A1(net5942),
    .A2(\scanline[89][1] ),
    .Y(_03823_),
    .B1(net5878));
 sg13g2_a221oi_1 _20615_ (.B2(_03823_),
    .C1(net5485),
    .B1(_03822_),
    .A1(net5878),
    .Y(_03824_),
    .A2(_03821_));
 sg13g2_mux4_1 _20616_ (.S0(net5963),
    .A0(\scanline[92][1] ),
    .A1(\scanline[93][1] ),
    .A2(\scanline[94][1] ),
    .A3(\scanline[95][1] ),
    .S1(net5901),
    .X(_03825_));
 sg13g2_mux4_1 _20617_ (.S0(net5944),
    .A0(\scanline[80][1] ),
    .A1(\scanline[81][1] ),
    .A2(\scanline[82][1] ),
    .A3(\scanline[83][1] ),
    .S1(net5887),
    .X(_03826_));
 sg13g2_mux4_1 _20618_ (.S0(net5951),
    .A0(\scanline[84][1] ),
    .A1(\scanline[85][1] ),
    .A2(\scanline[86][1] ),
    .A3(\scanline[87][1] ),
    .S1(net5892),
    .X(_03827_));
 sg13g2_nand2_1 _20619_ (.Y(_03828_),
    .A(net5507),
    .B(_03827_));
 sg13g2_a22oi_1 _20620_ (.Y(_03829_),
    .B1(_03826_),
    .B2(net5522),
    .A2(_03825_),
    .A1(net5534));
 sg13g2_nand2_1 _20621_ (.Y(_03830_),
    .A(_03828_),
    .B(_03829_));
 sg13g2_nor4_2 _20622_ (.A(net5552),
    .B(net5455),
    .C(_03824_),
    .Y(_03831_),
    .D(_03830_));
 sg13g2_nor4_2 _20623_ (.A(net5839),
    .B(_03812_),
    .C(_03819_),
    .Y(_03832_),
    .D(_03831_));
 sg13g2_a21oi_2 _20624_ (.B1(_03753_),
    .Y(_03833_),
    .A2(_03832_),
    .A1(_03797_));
 sg13g2_a21o_2 _20625_ (.A2(_03832_),
    .A1(_03797_),
    .B1(_03753_),
    .X(_03834_));
 sg13g2_nor2_2 _20626_ (.A(_08697_),
    .B(_03833_),
    .Y(_03835_));
 sg13g2_nand2_2 _20627_ (.Y(_03836_),
    .A(net5512),
    .B(_03834_));
 sg13g2_mux4_1 _20628_ (.S0(net5909),
    .A0(\scanline[140][0] ),
    .A1(\scanline[141][0] ),
    .A2(\scanline[142][0] ),
    .A3(\scanline[143][0] ),
    .S1(net5853),
    .X(_03837_));
 sg13g2_nor2_1 _20629_ (.A(net5525),
    .B(_03837_),
    .Y(_03838_));
 sg13g2_mux4_1 _20630_ (.S0(net5908),
    .A0(\scanline[136][0] ),
    .A1(\scanline[137][0] ),
    .A2(\scanline[138][0] ),
    .A3(\scanline[139][0] ),
    .S1(net5852),
    .X(_03839_));
 sg13g2_nor2_1 _20631_ (.A(net5483),
    .B(_03839_),
    .Y(_03840_));
 sg13g2_mux4_1 _20632_ (.S0(net5911),
    .A0(\scanline[128][0] ),
    .A1(\scanline[129][0] ),
    .A2(\scanline[130][0] ),
    .A3(\scanline[131][0] ),
    .S1(net5855),
    .X(_03841_));
 sg13g2_nor2_1 _20633_ (.A(net5514),
    .B(_03841_),
    .Y(_03842_));
 sg13g2_mux4_1 _20634_ (.S0(net5911),
    .A0(\scanline[132][0] ),
    .A1(\scanline[133][0] ),
    .A2(\scanline[134][0] ),
    .A3(\scanline[135][0] ),
    .S1(net5855),
    .X(_03843_));
 sg13g2_nor2_1 _20635_ (.A(net5497),
    .B(_03843_),
    .Y(_03844_));
 sg13g2_mux4_1 _20636_ (.S0(net5928),
    .A0(\scanline[152][0] ),
    .A1(\scanline[153][0] ),
    .A2(\scanline[154][0] ),
    .A3(\scanline[155][0] ),
    .S1(net5871),
    .X(_03845_));
 sg13g2_nor2_1 _20637_ (.A(net5484),
    .B(_03845_),
    .Y(_03846_));
 sg13g2_mux4_1 _20638_ (.S0(net5925),
    .A0(\scanline[144][0] ),
    .A1(\scanline[145][0] ),
    .A2(\scanline[146][0] ),
    .A3(\scanline[147][0] ),
    .S1(net5871),
    .X(_03847_));
 sg13g2_nor2_1 _20639_ (.A(net5514),
    .B(_03847_),
    .Y(_03848_));
 sg13g2_mux4_1 _20640_ (.S0(net5923),
    .A0(\scanline[156][0] ),
    .A1(\scanline[157][0] ),
    .A2(\scanline[158][0] ),
    .A3(\scanline[159][0] ),
    .S1(net5868),
    .X(_03849_));
 sg13g2_mux4_1 _20641_ (.S0(net5929),
    .A0(\scanline[148][0] ),
    .A1(\scanline[149][0] ),
    .A2(\scanline[150][0] ),
    .A3(\scanline[151][0] ),
    .S1(net5873),
    .X(_03850_));
 sg13g2_nor2_1 _20642_ (.A(net5498),
    .B(_03850_),
    .Y(_03851_));
 sg13g2_nor3_1 _20643_ (.A(_03846_),
    .B(_03848_),
    .C(_03851_),
    .Y(_03852_));
 sg13g2_o21ai_1 _20644_ (.B1(_03852_),
    .Y(_03853_),
    .A1(net5525),
    .A2(_03849_));
 sg13g2_nor4_2 _20645_ (.A(_03838_),
    .B(_03840_),
    .C(_03842_),
    .Y(_03854_),
    .D(_03844_));
 sg13g2_o21ai_1 _20646_ (.B1(_08686_),
    .Y(_03855_),
    .A1(net5844),
    .A2(_03854_));
 sg13g2_a21oi_2 _20647_ (.B1(_03855_),
    .Y(_03856_),
    .A2(_03853_),
    .A1(net5844));
 sg13g2_mux4_1 _20648_ (.S0(net5932),
    .A0(\scanline[32][0] ),
    .A1(\scanline[33][0] ),
    .A2(\scanline[34][0] ),
    .A3(\scanline[35][0] ),
    .S1(net5877),
    .X(_03857_));
 sg13g2_mux4_1 _20649_ (.S0(net5915),
    .A0(\scanline[40][0] ),
    .A1(\scanline[41][0] ),
    .A2(\scanline[42][0] ),
    .A3(\scanline[43][0] ),
    .S1(net5859),
    .X(_03858_));
 sg13g2_mux4_1 _20650_ (.S0(net5926),
    .A0(\scanline[44][0] ),
    .A1(\scanline[45][0] ),
    .A2(\scanline[46][0] ),
    .A3(\scanline[47][0] ),
    .S1(net5870),
    .X(_03859_));
 sg13g2_mux4_1 _20651_ (.S0(net5931),
    .A0(\scanline[36][0] ),
    .A1(\scanline[37][0] ),
    .A2(\scanline[38][0] ),
    .A3(\scanline[39][0] ),
    .S1(net5875),
    .X(_03860_));
 sg13g2_and2_1 _20652_ (.A(net5501),
    .B(_03860_),
    .X(_03861_));
 sg13g2_a21oi_1 _20653_ (.A1(net5531),
    .A2(_03859_),
    .Y(_03862_),
    .B1(net5845));
 sg13g2_a221oi_1 _20654_ (.B2(net5487),
    .C1(_03861_),
    .B1(_03858_),
    .A1(net5518),
    .Y(_03863_),
    .A2(_03857_));
 sg13g2_mux4_1 _20655_ (.S0(net5929),
    .A0(\scanline[52][0] ),
    .A1(\scanline[53][0] ),
    .A2(\scanline[54][0] ),
    .A3(\scanline[55][0] ),
    .S1(net5873),
    .X(_03864_));
 sg13g2_mux4_1 _20656_ (.S0(net5951),
    .A0(\scanline[60][0] ),
    .A1(\scanline[61][0] ),
    .A2(\scanline[62][0] ),
    .A3(\scanline[63][0] ),
    .S1(net5892),
    .X(_03865_));
 sg13g2_mux4_1 _20657_ (.S0(net5950),
    .A0(\scanline[56][0] ),
    .A1(\scanline[57][0] ),
    .A2(\scanline[58][0] ),
    .A3(\scanline[59][0] ),
    .S1(net5890),
    .X(_03866_));
 sg13g2_nand2b_1 _20658_ (.Y(_03867_),
    .B(\scanline[48][0] ),
    .A_N(net5926));
 sg13g2_a21oi_1 _20659_ (.A1(net5926),
    .A2(\scanline[49][0] ),
    .Y(_03868_),
    .B1(net5870));
 sg13g2_nand2_1 _20660_ (.Y(_03869_),
    .A(net5926),
    .B(\scanline[51][0] ));
 sg13g2_nand2b_1 _20661_ (.Y(_03870_),
    .B(\scanline[50][0] ),
    .A_N(net5926));
 sg13g2_nand3_1 _20662_ (.B(_03869_),
    .C(_03870_),
    .A(net5870),
    .Y(_03871_));
 sg13g2_a21oi_1 _20663_ (.A1(_03867_),
    .A2(_03868_),
    .Y(_03872_),
    .B1(net5516));
 sg13g2_a22oi_1 _20664_ (.Y(_03873_),
    .B1(_03866_),
    .B2(net5493),
    .A2(_03865_),
    .A1(net5531));
 sg13g2_a221oi_1 _20665_ (.B2(_03872_),
    .C1(net5556),
    .B1(_03871_),
    .A1(net5502),
    .Y(_03874_),
    .A2(_03864_));
 sg13g2_a22oi_1 _20666_ (.Y(_03875_),
    .B1(_03873_),
    .B2(_03874_),
    .A2(_03863_),
    .A1(_03862_));
 sg13g2_mux4_1 _20667_ (.S0(net5935),
    .A0(\scanline[0][0] ),
    .A1(\scanline[1][0] ),
    .A2(\scanline[2][0] ),
    .A3(\scanline[3][0] ),
    .S1(net5878),
    .X(_03876_));
 sg13g2_mux4_1 _20668_ (.S0(net5933),
    .A0(\scanline[4][0] ),
    .A1(\scanline[5][0] ),
    .A2(\scanline[6][0] ),
    .A3(\scanline[7][0] ),
    .S1(net5876),
    .X(_03877_));
 sg13g2_a22oi_1 _20669_ (.Y(_03878_),
    .B1(_03877_),
    .B2(net5504),
    .A2(_03876_),
    .A1(net5521));
 sg13g2_mux4_1 _20670_ (.S0(net5936),
    .A0(\scanline[12][0] ),
    .A1(\scanline[13][0] ),
    .A2(\scanline[14][0] ),
    .A3(\scanline[15][0] ),
    .S1(net5880),
    .X(_03879_));
 sg13g2_mux4_1 _20671_ (.S0(net5931),
    .A0(\scanline[8][0] ),
    .A1(\scanline[9][0] ),
    .A2(\scanline[10][0] ),
    .A3(\scanline[11][0] ),
    .S1(net5875),
    .X(_03880_));
 sg13g2_a22oi_1 _20672_ (.Y(_03881_),
    .B1(_03880_),
    .B2(net5490),
    .A2(_03879_),
    .A1(net5530));
 sg13g2_a21o_2 _20673_ (.A2(_03881_),
    .A1(_03878_),
    .B1(net5510),
    .X(_03882_));
 sg13g2_mux4_1 _20674_ (.S0(net5938),
    .A0(\scanline[24][0] ),
    .A1(\scanline[25][0] ),
    .A2(\scanline[26][0] ),
    .A3(\scanline[27][0] ),
    .S1(net5882),
    .X(_03883_));
 sg13g2_mux4_1 _20675_ (.S0(net5944),
    .A0(\scanline[16][0] ),
    .A1(\scanline[17][0] ),
    .A2(\scanline[18][0] ),
    .A3(\scanline[19][0] ),
    .S1(net5887),
    .X(_03884_));
 sg13g2_mux4_1 _20676_ (.S0(net5938),
    .A0(\scanline[20][0] ),
    .A1(\scanline[21][0] ),
    .A2(\scanline[22][0] ),
    .A3(\scanline[23][0] ),
    .S1(net5882),
    .X(_03885_));
 sg13g2_mux4_1 _20677_ (.S0(net5939),
    .A0(\scanline[28][0] ),
    .A1(\scanline[29][0] ),
    .A2(\scanline[30][0] ),
    .A3(\scanline[31][0] ),
    .S1(net5883),
    .X(_03886_));
 sg13g2_a22oi_1 _20678_ (.Y(_03887_),
    .B1(_03886_),
    .B2(net5533),
    .A2(_03884_),
    .A1(net5520));
 sg13g2_a22oi_1 _20679_ (.Y(_03888_),
    .B1(_03885_),
    .B2(net5505),
    .A2(_03883_),
    .A1(net5489));
 sg13g2_nand2_2 _20680_ (.Y(_03889_),
    .A(_03887_),
    .B(_03888_));
 sg13g2_a221oi_1 _20681_ (.B2(_03392_),
    .C1(net5841),
    .B1(_03889_),
    .A1(net5842),
    .Y(_03890_),
    .A2(_03875_));
 sg13g2_mux4_1 _20682_ (.S0(net5957),
    .A0(\scanline[104][0] ),
    .A1(\scanline[105][0] ),
    .A2(\scanline[106][0] ),
    .A3(\scanline[107][0] ),
    .S1(net5897),
    .X(_03891_));
 sg13g2_mux4_1 _20683_ (.S0(net5954),
    .A0(\scanline[100][0] ),
    .A1(\scanline[101][0] ),
    .A2(\scanline[102][0] ),
    .A3(\scanline[103][0] ),
    .S1(net5895),
    .X(_03892_));
 sg13g2_mux4_1 _20684_ (.S0(net5953),
    .A0(\scanline[108][0] ),
    .A1(\scanline[109][0] ),
    .A2(\scanline[110][0] ),
    .A3(\scanline[111][0] ),
    .S1(net5895),
    .X(_03893_));
 sg13g2_mux4_1 _20685_ (.S0(net5952),
    .A0(\scanline[96][0] ),
    .A1(\scanline[97][0] ),
    .A2(\scanline[98][0] ),
    .A3(\scanline[99][0] ),
    .S1(net5893),
    .X(_03894_));
 sg13g2_a22oi_1 _20686_ (.Y(_03895_),
    .B1(_03894_),
    .B2(net5523),
    .A2(_03891_),
    .A1(net5493));
 sg13g2_a221oi_1 _20687_ (.B2(net5531),
    .C1(net5847),
    .B1(_03893_),
    .A1(net5502),
    .Y(_03896_),
    .A2(_03892_));
 sg13g2_nand2_1 _20688_ (.Y(_03897_),
    .A(_03895_),
    .B(_03896_));
 sg13g2_mux4_1 _20689_ (.S0(net5966),
    .A0(\scanline[120][0] ),
    .A1(\scanline[121][0] ),
    .A2(\scanline[122][0] ),
    .A3(\scanline[123][0] ),
    .S1(net5904),
    .X(_03898_));
 sg13g2_nand2_1 _20690_ (.Y(_03899_),
    .A(net5491),
    .B(_03898_));
 sg13g2_mux4_1 _20691_ (.S0(net5965),
    .A0(\scanline[116][0] ),
    .A1(\scanline[117][0] ),
    .A2(\scanline[118][0] ),
    .A3(\scanline[119][0] ),
    .S1(net5904),
    .X(_03900_));
 sg13g2_mux4_1 _20692_ (.S0(net5961),
    .A0(\scanline[124][0] ),
    .A1(\scanline[125][0] ),
    .A2(\scanline[126][0] ),
    .A3(\scanline[127][0] ),
    .S1(net5900),
    .X(_03901_));
 sg13g2_nand2_1 _20693_ (.Y(_03902_),
    .A(net5534),
    .B(_03901_));
 sg13g2_a21oi_1 _20694_ (.A1(net5962),
    .A2(\scanline[113][0] ),
    .Y(_03903_),
    .B1(net5900));
 sg13g2_o21ai_1 _20695_ (.B1(_03903_),
    .Y(_03904_),
    .A1(net5962),
    .A2(_08128_));
 sg13g2_nand2_1 _20696_ (.Y(_03905_),
    .A(net5963),
    .B(\scanline[115][0] ));
 sg13g2_nand2b_1 _20697_ (.Y(_03906_),
    .B(\scanline[114][0] ),
    .A_N(net5963));
 sg13g2_nand3_1 _20698_ (.B(_03905_),
    .C(_03906_),
    .A(net5900),
    .Y(_03907_));
 sg13g2_nand3_1 _20699_ (.B(_03904_),
    .C(_03907_),
    .A(net5522),
    .Y(_03908_));
 sg13g2_a21oi_1 _20700_ (.A1(net5508),
    .A2(_03900_),
    .Y(_03909_),
    .B1(net5554));
 sg13g2_nand4_1 _20701_ (.B(_03902_),
    .C(_03908_),
    .A(_03899_),
    .Y(_03910_),
    .D(_03909_));
 sg13g2_nand3_1 _20702_ (.B(_03897_),
    .C(_03910_),
    .A(net5842),
    .Y(_03911_));
 sg13g2_mux4_1 _20703_ (.S0(net5963),
    .A0(\scanline[92][0] ),
    .A1(\scanline[93][0] ),
    .A2(\scanline[94][0] ),
    .A3(\scanline[95][0] ),
    .S1(net5901),
    .X(_03912_));
 sg13g2_mux4_1 _20704_ (.S0(net5960),
    .A0(\scanline[84][0] ),
    .A1(\scanline[85][0] ),
    .A2(\scanline[86][0] ),
    .A3(\scanline[87][0] ),
    .S1(net5899),
    .X(_03913_));
 sg13g2_a22oi_1 _20705_ (.Y(_03914_),
    .B1(_03913_),
    .B2(net5506),
    .A2(_03912_),
    .A1(net5534));
 sg13g2_mux4_1 _20706_ (.S0(net5944),
    .A0(\scanline[80][0] ),
    .A1(\scanline[81][0] ),
    .A2(\scanline[82][0] ),
    .A3(\scanline[83][0] ),
    .S1(net5887),
    .X(_03915_));
 sg13g2_mux4_1 _20707_ (.S0(net5942),
    .A0(\scanline[88][0] ),
    .A1(\scanline[89][0] ),
    .A2(\scanline[90][0] ),
    .A3(\scanline[91][0] ),
    .S1(net5886),
    .X(_03916_));
 sg13g2_a22oi_1 _20708_ (.Y(_03917_),
    .B1(_03916_),
    .B2(net5489),
    .A2(_03915_),
    .A1(net5521));
 sg13g2_a21oi_2 _20709_ (.B1(net5455),
    .Y(_03918_),
    .A2(_03917_),
    .A1(_03914_));
 sg13g2_mux4_1 _20710_ (.S0(net5908),
    .A0(\scanline[76][0] ),
    .A1(\scanline[77][0] ),
    .A2(\scanline[78][0] ),
    .A3(\scanline[79][0] ),
    .S1(net5852),
    .X(_03919_));
 sg13g2_mux4_1 _20711_ (.S0(net5907),
    .A0(\scanline[72][0] ),
    .A1(\scanline[73][0] ),
    .A2(\scanline[74][0] ),
    .A3(\scanline[75][0] ),
    .S1(net5851),
    .X(_03920_));
 sg13g2_mux4_1 _20712_ (.S0(net5913),
    .A0(\scanline[68][0] ),
    .A1(\scanline[69][0] ),
    .A2(\scanline[70][0] ),
    .A3(\scanline[71][0] ),
    .S1(net5857),
    .X(_03921_));
 sg13g2_mux4_1 _20713_ (.S0(net5914),
    .A0(\scanline[64][0] ),
    .A1(\scanline[65][0] ),
    .A2(\scanline[66][0] ),
    .A3(\scanline[67][0] ),
    .S1(net5858),
    .X(_03922_));
 sg13g2_a22oi_1 _20714_ (.Y(_03923_),
    .B1(_03922_),
    .B2(net5517),
    .A2(_03920_),
    .A1(net5486));
 sg13g2_a22oi_1 _20715_ (.Y(_03924_),
    .B1(_03921_),
    .B2(net5500),
    .A2(_03919_),
    .A1(net5529));
 sg13g2_a21oi_2 _20716_ (.B1(net5509),
    .Y(_03925_),
    .A2(_03924_),
    .A1(_03923_));
 sg13g2_nor3_1 _20717_ (.A(net5552),
    .B(_03918_),
    .C(_03925_),
    .Y(_03926_));
 sg13g2_a221oi_1 _20718_ (.B2(_03926_),
    .C1(\hvsync_gen.hpos[9] ),
    .B1(_03911_),
    .A1(_03882_),
    .Y(_03927_),
    .A2(_03890_));
 sg13g2_nor2_1 _20719_ (.A(_03856_),
    .B(_03927_),
    .Y(_03928_));
 sg13g2_or2_2 _20720_ (.X(_03929_),
    .B(_03927_),
    .A(_03856_));
 sg13g2_o21ai_1 _20721_ (.B1(net5512),
    .Y(_03930_),
    .A1(_03856_),
    .A2(_03927_));
 sg13g2_nor2_2 _20722_ (.A(_03833_),
    .B(net5328),
    .Y(_03931_));
 sg13g2_inv_1 _20723_ (.Y(_03932_),
    .A(_03931_));
 sg13g2_a21oi_2 _20724_ (.B1(_03732_),
    .Y(_03933_),
    .A2(_03929_),
    .A1(_03835_));
 sg13g2_and3_1 _20725_ (.X(_03934_),
    .A(net5512),
    .B(net5360),
    .C(_03834_));
 sg13g2_and2_1 _20726_ (.A(_03929_),
    .B(net5326),
    .X(_03935_));
 sg13g2_nand2_2 _20727_ (.Y(_03936_),
    .A(_03929_),
    .B(net5326));
 sg13g2_nand2b_1 _20728_ (.Y(_03937_),
    .B(_03936_),
    .A_N(_03933_));
 sg13g2_o21ai_1 _20729_ (.B1(net5337),
    .Y(_03938_),
    .A1(_03933_),
    .A2(_03935_));
 sg13g2_nand2_1 _20730_ (.Y(_03939_),
    .A(_03835_),
    .B(net5330));
 sg13g2_nor3_2 _20731_ (.A(_08697_),
    .B(net5360),
    .C(_03833_),
    .Y(_03940_));
 sg13g2_nand2_1 _20732_ (.Y(_03941_),
    .A(net5330),
    .B(_03940_));
 sg13g2_nand3_1 _20733_ (.B(_03936_),
    .C(net5285),
    .A(net5333),
    .Y(_03942_));
 sg13g2_nand2_1 _20734_ (.Y(_03943_),
    .A(_03938_),
    .B(_03942_));
 sg13g2_a21oi_1 _20735_ (.A1(net5334),
    .A2(_03937_),
    .Y(_03944_),
    .B1(net5294));
 sg13g2_a21o_1 _20736_ (.A2(net5285),
    .A1(_03936_),
    .B1(net5334),
    .X(_03945_));
 sg13g2_a22oi_1 _20737_ (.Y(_03946_),
    .B1(_03944_),
    .B2(_03945_),
    .A2(_03943_),
    .A1(net5294));
 sg13g2_mux4_1 _20738_ (.S0(net5925),
    .A0(\scanline[152][6] ),
    .A1(\scanline[153][6] ),
    .A2(\scanline[154][6] ),
    .A3(\scanline[155][6] ),
    .S1(net5871),
    .X(_03947_));
 sg13g2_nor2_1 _20739_ (.A(net5484),
    .B(_03947_),
    .Y(_03948_));
 sg13g2_mux4_1 _20740_ (.S0(net5928),
    .A0(\scanline[148][6] ),
    .A1(\scanline[149][6] ),
    .A2(\scanline[150][6] ),
    .A3(\scanline[151][6] ),
    .S1(net5871),
    .X(_03949_));
 sg13g2_mux4_1 _20741_ (.S0(net5922),
    .A0(\scanline[156][6] ),
    .A1(\scanline[157][6] ),
    .A2(\scanline[158][6] ),
    .A3(\scanline[159][6] ),
    .S1(net5866),
    .X(_03950_));
 sg13g2_nor2_1 _20742_ (.A(net5526),
    .B(_03950_),
    .Y(_03951_));
 sg13g2_mux4_1 _20743_ (.S0(net5925),
    .A0(\scanline[144][6] ),
    .A1(\scanline[145][6] ),
    .A2(\scanline[146][6] ),
    .A3(\scanline[147][6] ),
    .S1(net5871),
    .X(_03952_));
 sg13g2_nor2_1 _20744_ (.A(net5514),
    .B(_03952_),
    .Y(_03953_));
 sg13g2_mux4_1 _20745_ (.S0(net5918),
    .A0(\scanline[128][6] ),
    .A1(\scanline[129][6] ),
    .A2(\scanline[130][6] ),
    .A3(\scanline[131][6] ),
    .S1(net5864),
    .X(_03954_));
 sg13g2_nor2_1 _20746_ (.A(net5514),
    .B(_03954_),
    .Y(_03955_));
 sg13g2_mux4_1 _20747_ (.S0(net5909),
    .A0(\scanline[140][6] ),
    .A1(\scanline[141][6] ),
    .A2(\scanline[142][6] ),
    .A3(\scanline[143][6] ),
    .S1(net5853),
    .X(_03956_));
 sg13g2_mux4_1 _20748_ (.S0(net5912),
    .A0(\scanline[136][6] ),
    .A1(\scanline[137][6] ),
    .A2(\scanline[138][6] ),
    .A3(\scanline[139][6] ),
    .S1(net5856),
    .X(_03957_));
 sg13g2_nor2_1 _20749_ (.A(net5483),
    .B(_03957_),
    .Y(_03958_));
 sg13g2_mux4_1 _20750_ (.S0(net5910),
    .A0(\scanline[132][6] ),
    .A1(\scanline[133][6] ),
    .A2(\scanline[134][6] ),
    .A3(\scanline[135][6] ),
    .S1(net5854),
    .X(_03959_));
 sg13g2_nor2_1 _20751_ (.A(net5497),
    .B(_03959_),
    .Y(_03960_));
 sg13g2_nor2_1 _20752_ (.A(_03955_),
    .B(_03960_),
    .Y(_03961_));
 sg13g2_o21ai_1 _20753_ (.B1(_03961_),
    .Y(_03962_),
    .A1(net5525),
    .A2(_03956_));
 sg13g2_o21ai_1 _20754_ (.B1(net5553),
    .Y(_03963_),
    .A1(_03958_),
    .A2(_03962_));
 sg13g2_nor2_1 _20755_ (.A(_03948_),
    .B(_03953_),
    .Y(_03964_));
 sg13g2_o21ai_1 _20756_ (.B1(_03964_),
    .Y(_03965_),
    .A1(net5498),
    .A2(_03949_));
 sg13g2_o21ai_1 _20757_ (.B1(net5844),
    .Y(_03966_),
    .A1(_03951_),
    .A2(_03965_));
 sg13g2_and2_1 _20758_ (.A(_03351_),
    .B(_03966_),
    .X(_03967_));
 sg13g2_mux4_1 _20759_ (.S0(net5953),
    .A0(\scanline[52][6] ),
    .A1(\scanline[53][6] ),
    .A2(\scanline[54][6] ),
    .A3(\scanline[55][6] ),
    .S1(net5895),
    .X(_03968_));
 sg13g2_a21oi_2 _20760_ (.B1(net5554),
    .Y(_03969_),
    .A2(_03968_),
    .A1(net5502));
 sg13g2_mux4_1 _20761_ (.S0(net5936),
    .A0(\scanline[56][6] ),
    .A1(\scanline[57][6] ),
    .A2(\scanline[58][6] ),
    .A3(\scanline[59][6] ),
    .S1(net5880),
    .X(_03970_));
 sg13g2_nand2b_1 _20762_ (.Y(_03971_),
    .B(\scanline[60][6] ),
    .A_N(net5951));
 sg13g2_a21oi_1 _20763_ (.A1(net5951),
    .A2(\scanline[61][6] ),
    .Y(_03972_),
    .B1(net5892));
 sg13g2_nor2b_1 _20764_ (.A(net5951),
    .B_N(\scanline[62][6] ),
    .Y(_03973_));
 sg13g2_a21oi_1 _20765_ (.A1(net5951),
    .A2(\scanline[63][6] ),
    .Y(_03974_),
    .B1(_03973_));
 sg13g2_a221oi_1 _20766_ (.B2(net5892),
    .C1(net5528),
    .B1(_03974_),
    .A1(_03971_),
    .Y(_03975_),
    .A2(_03972_));
 sg13g2_mux4_1 _20767_ (.S0(net5927),
    .A0(\scanline[48][6] ),
    .A1(\scanline[49][6] ),
    .A2(\scanline[50][6] ),
    .A3(\scanline[51][6] ),
    .S1(net5870),
    .X(_03976_));
 sg13g2_a221oi_1 _20768_ (.B2(net5519),
    .C1(_03975_),
    .B1(_03976_),
    .A1(net5488),
    .Y(_03977_),
    .A2(_03970_));
 sg13g2_mux4_1 _20769_ (.S0(net5920),
    .A0(\scanline[44][6] ),
    .A1(\scanline[45][6] ),
    .A2(\scanline[46][6] ),
    .A3(\scanline[47][6] ),
    .S1(net5862),
    .X(_03978_));
 sg13g2_mux4_1 _20770_ (.S0(net5936),
    .A0(\scanline[32][6] ),
    .A1(\scanline[33][6] ),
    .A2(\scanline[34][6] ),
    .A3(\scanline[35][6] ),
    .S1(net5880),
    .X(_03979_));
 sg13g2_mux4_1 _20771_ (.S0(net5931),
    .A0(\scanline[36][6] ),
    .A1(\scanline[37][6] ),
    .A2(\scanline[38][6] ),
    .A3(\scanline[39][6] ),
    .S1(net5875),
    .X(_03980_));
 sg13g2_mux4_1 _20772_ (.S0(net5915),
    .A0(\scanline[40][6] ),
    .A1(\scanline[41][6] ),
    .A2(\scanline[42][6] ),
    .A3(\scanline[43][6] ),
    .S1(net5859),
    .X(_03981_));
 sg13g2_a22oi_1 _20773_ (.Y(_03982_),
    .B1(_03980_),
    .B2(net5501),
    .A2(_03979_),
    .A1(net5518));
 sg13g2_a221oi_1 _20774_ (.B2(net5488),
    .C1(net5845),
    .B1(_03981_),
    .A1(net5531),
    .Y(_03983_),
    .A2(_03978_));
 sg13g2_a221oi_1 _20775_ (.B2(_03983_),
    .C1(_08117_),
    .B1(_03982_),
    .A1(_03969_),
    .Y(_03984_),
    .A2(_03977_));
 sg13g2_mux4_1 _20776_ (.S0(net5939),
    .A0(\scanline[20][6] ),
    .A1(\scanline[21][6] ),
    .A2(\scanline[22][6] ),
    .A3(\scanline[23][6] ),
    .S1(net5883),
    .X(_03985_));
 sg13g2_mux4_1 _20777_ (.S0(net5940),
    .A0(\scanline[16][6] ),
    .A1(\scanline[17][6] ),
    .A2(\scanline[18][6] ),
    .A3(\scanline[19][6] ),
    .S1(net5884),
    .X(_03986_));
 sg13g2_a22oi_1 _20778_ (.Y(_03987_),
    .B1(_03986_),
    .B2(net5520),
    .A2(_03985_),
    .A1(net5505));
 sg13g2_mux4_1 _20779_ (.S0(net5938),
    .A0(\scanline[24][6] ),
    .A1(\scanline[25][6] ),
    .A2(\scanline[26][6] ),
    .A3(\scanline[27][6] ),
    .S1(net5882),
    .X(_03988_));
 sg13g2_mux4_1 _20780_ (.S0(net5942),
    .A0(\scanline[28][6] ),
    .A1(\scanline[29][6] ),
    .A2(\scanline[30][6] ),
    .A3(\scanline[31][6] ),
    .S1(net5886),
    .X(_03989_));
 sg13g2_a22oi_1 _20781_ (.Y(_03990_),
    .B1(_03989_),
    .B2(net5532),
    .A2(_03988_),
    .A1(net5489));
 sg13g2_a21o_2 _20782_ (.A2(_03990_),
    .A1(_03987_),
    .B1(net5455),
    .X(_03991_));
 sg13g2_mux4_1 _20783_ (.S0(net5933),
    .A0(\scanline[4][6] ),
    .A1(\scanline[5][6] ),
    .A2(\scanline[6][6] ),
    .A3(\scanline[7][6] ),
    .S1(net5876),
    .X(_03992_));
 sg13g2_mux4_1 _20784_ (.S0(net5936),
    .A0(\scanline[12][6] ),
    .A1(\scanline[13][6] ),
    .A2(\scanline[14][6] ),
    .A3(\scanline[15][6] ),
    .S1(net5880),
    .X(_03993_));
 sg13g2_mux4_1 _20785_ (.S0(net5931),
    .A0(\scanline[8][6] ),
    .A1(\scanline[9][6] ),
    .A2(\scanline[10][6] ),
    .A3(\scanline[11][6] ),
    .S1(net5875),
    .X(_03994_));
 sg13g2_mux4_1 _20786_ (.S0(net5937),
    .A0(\scanline[0][6] ),
    .A1(\scanline[1][6] ),
    .A2(\scanline[2][6] ),
    .A3(\scanline[3][6] ),
    .S1(net5879),
    .X(_03995_));
 sg13g2_a22oi_1 _20787_ (.Y(_03996_),
    .B1(_03995_),
    .B2(net5517),
    .A2(_03993_),
    .A1(net5532));
 sg13g2_a22oi_1 _20788_ (.Y(_03997_),
    .B1(_03994_),
    .B2(net5490),
    .A2(_03992_),
    .A1(net5504));
 sg13g2_a21oi_2 _20789_ (.B1(net5509),
    .Y(_03998_),
    .A2(_03997_),
    .A1(_03996_));
 sg13g2_nor3_1 _20790_ (.A(net5840),
    .B(_03984_),
    .C(_03998_),
    .Y(_03999_));
 sg13g2_mux4_1 _20791_ (.S0(net5959),
    .A0(\scanline[124][6] ),
    .A1(\scanline[125][6] ),
    .A2(\scanline[126][6] ),
    .A3(\scanline[127][6] ),
    .S1(net5899),
    .X(_04000_));
 sg13g2_mux4_1 _20792_ (.S0(net5964),
    .A0(\scanline[120][6] ),
    .A1(\scanline[121][6] ),
    .A2(\scanline[122][6] ),
    .A3(\scanline[123][6] ),
    .S1(net5903),
    .X(_04001_));
 sg13g2_nand2b_1 _20793_ (.Y(_04002_),
    .B(\scanline[116][6] ),
    .A_N(net5964));
 sg13g2_a21oi_1 _20794_ (.A1(net5964),
    .A2(\scanline[117][6] ),
    .Y(_04003_),
    .B1(net5903));
 sg13g2_nor2b_1 _20795_ (.A(net5965),
    .B_N(\scanline[118][6] ),
    .Y(_04004_));
 sg13g2_a21oi_1 _20796_ (.A1(net5965),
    .A2(\scanline[119][6] ),
    .Y(_04005_),
    .B1(_04004_));
 sg13g2_a221oi_1 _20797_ (.B2(net5903),
    .C1(net5499),
    .B1(_04005_),
    .A1(_04002_),
    .Y(_04006_),
    .A2(_04003_));
 sg13g2_mux4_1 _20798_ (.S0(net5963),
    .A0(\scanline[112][6] ),
    .A1(\scanline[113][6] ),
    .A2(\scanline[114][6] ),
    .A3(\scanline[115][6] ),
    .S1(net5901),
    .X(_04007_));
 sg13g2_nand2_2 _20799_ (.Y(_04008_),
    .A(net5522),
    .B(_04007_));
 sg13g2_nand2b_1 _20800_ (.Y(_04009_),
    .B(net5848),
    .A_N(_04006_));
 sg13g2_a221oi_1 _20801_ (.B2(net5491),
    .C1(_04009_),
    .B1(_04001_),
    .A1(net5535),
    .Y(_04010_),
    .A2(_04000_));
 sg13g2_mux4_1 _20802_ (.S0(net5955),
    .A0(\scanline[100][6] ),
    .A1(\scanline[101][6] ),
    .A2(\scanline[102][6] ),
    .A3(\scanline[103][6] ),
    .S1(net5896),
    .X(_04011_));
 sg13g2_nor2b_1 _20803_ (.A(net5956),
    .B_N(\scanline[106][6] ),
    .Y(_04012_));
 sg13g2_a21oi_1 _20804_ (.A1(net5956),
    .A2(\scanline[107][6] ),
    .Y(_04013_),
    .B1(_04012_));
 sg13g2_nand2b_1 _20805_ (.Y(_04014_),
    .B(\scanline[104][6] ),
    .A_N(net5956));
 sg13g2_a21oi_1 _20806_ (.A1(net5956),
    .A2(\scanline[105][6] ),
    .Y(_04015_),
    .B1(net5896));
 sg13g2_a221oi_1 _20807_ (.B2(_04015_),
    .C1(net5485),
    .B1(_04014_),
    .A1(net5896),
    .Y(_04016_),
    .A2(_04013_));
 sg13g2_mux4_1 _20808_ (.S0(net5951),
    .A0(\scanline[96][6] ),
    .A1(\scanline[97][6] ),
    .A2(\scanline[98][6] ),
    .A3(\scanline[99][6] ),
    .S1(net5892),
    .X(_04017_));
 sg13g2_mux4_1 _20809_ (.S0(net5955),
    .A0(\scanline[108][6] ),
    .A1(\scanline[109][6] ),
    .A2(\scanline[110][6] ),
    .A3(\scanline[111][6] ),
    .S1(net5896),
    .X(_04018_));
 sg13g2_a21oi_1 _20810_ (.A1(net5523),
    .A2(_04017_),
    .Y(_04019_),
    .B1(net5848));
 sg13g2_a221oi_1 _20811_ (.B2(net5535),
    .C1(_04016_),
    .B1(_04018_),
    .A1(net5507),
    .Y(_04020_),
    .A2(_04011_));
 sg13g2_a22oi_1 _20812_ (.Y(_04021_),
    .B1(_04019_),
    .B2(_04020_),
    .A2(_04010_),
    .A1(_04008_));
 sg13g2_nand2_1 _20813_ (.Y(_04022_),
    .A(net5842),
    .B(_04021_));
 sg13g2_mux4_1 _20814_ (.S0(net5945),
    .A0(\scanline[80][6] ),
    .A1(\scanline[81][6] ),
    .A2(\scanline[82][6] ),
    .A3(\scanline[83][6] ),
    .S1(net5888),
    .X(_04023_));
 sg13g2_mux4_1 _20815_ (.S0(net5943),
    .A0(\scanline[88][6] ),
    .A1(\scanline[89][6] ),
    .A2(\scanline[90][6] ),
    .A3(\scanline[91][6] ),
    .S1(net5886),
    .X(_04024_));
 sg13g2_mux4_1 _20816_ (.S0(net5944),
    .A0(\scanline[92][6] ),
    .A1(\scanline[93][6] ),
    .A2(\scanline[94][6] ),
    .A3(\scanline[95][6] ),
    .S1(net5887),
    .X(_04025_));
 sg13g2_mux4_1 _20817_ (.S0(net5943),
    .A0(\scanline[84][6] ),
    .A1(\scanline[85][6] ),
    .A2(\scanline[86][6] ),
    .A3(\scanline[87][6] ),
    .S1(net5886),
    .X(_04026_));
 sg13g2_a22oi_1 _20818_ (.Y(_04027_),
    .B1(_04026_),
    .B2(net5506),
    .A2(_04024_),
    .A1(net5492));
 sg13g2_a22oi_1 _20819_ (.Y(_04028_),
    .B1(_04025_),
    .B2(net5534),
    .A2(_04023_),
    .A1(net5522));
 sg13g2_a21oi_2 _20820_ (.B1(net5455),
    .Y(_04029_),
    .A2(_04028_),
    .A1(_04027_));
 sg13g2_mux4_1 _20821_ (.S0(net5913),
    .A0(\scanline[68][6] ),
    .A1(\scanline[69][6] ),
    .A2(\scanline[70][6] ),
    .A3(\scanline[71][6] ),
    .S1(net5857),
    .X(_04030_));
 sg13g2_mux4_1 _20822_ (.S0(net5914),
    .A0(\scanline[64][6] ),
    .A1(\scanline[65][6] ),
    .A2(\scanline[66][6] ),
    .A3(\scanline[67][6] ),
    .S1(net5858),
    .X(_04031_));
 sg13g2_a22oi_1 _20823_ (.Y(_04032_),
    .B1(_04031_),
    .B2(net5517),
    .A2(_04030_),
    .A1(net5500));
 sg13g2_mux4_1 _20824_ (.S0(net5907),
    .A0(\scanline[72][6] ),
    .A1(\scanline[73][6] ),
    .A2(\scanline[74][6] ),
    .A3(\scanline[75][6] ),
    .S1(net5851),
    .X(_04033_));
 sg13g2_mux4_1 _20825_ (.S0(net5907),
    .A0(\scanline[76][6] ),
    .A1(\scanline[77][6] ),
    .A2(\scanline[78][6] ),
    .A3(\scanline[79][6] ),
    .S1(net5851),
    .X(_04034_));
 sg13g2_a22oi_1 _20826_ (.Y(_04035_),
    .B1(_04034_),
    .B2(net5529),
    .A2(_04033_),
    .A1(net5486));
 sg13g2_a21oi_2 _20827_ (.B1(net5509),
    .Y(_04036_),
    .A2(_04035_),
    .A1(_04032_));
 sg13g2_nor3_1 _20828_ (.A(net5552),
    .B(_04029_),
    .C(_04036_),
    .Y(_04037_));
 sg13g2_a221oi_1 _20829_ (.B2(_04037_),
    .C1(net5839),
    .B1(_04022_),
    .A1(_03991_),
    .Y(_04038_),
    .A2(_03999_));
 sg13g2_a21oi_2 _20830_ (.B1(_04038_),
    .Y(_04039_),
    .A2(_03967_),
    .A1(_03963_));
 sg13g2_a21o_2 _20831_ (.A2(_03967_),
    .A1(_03963_),
    .B1(_04038_),
    .X(_04040_));
 sg13g2_nor2_2 _20832_ (.A(net5331),
    .B(net5330),
    .Y(_04041_));
 sg13g2_inv_1 _20833_ (.Y(_04042_),
    .A(_04041_));
 sg13g2_nor2_1 _20834_ (.A(_03834_),
    .B(net5328),
    .Y(_04043_));
 sg13g2_o21ai_1 _20835_ (.B1(net5301),
    .Y(_04044_),
    .A1(_04041_),
    .A2(net5284));
 sg13g2_and2_1 _20836_ (.A(_04040_),
    .B(_04044_),
    .X(_04045_));
 sg13g2_o21ai_1 _20837_ (.B1(_04045_),
    .Y(_04046_),
    .A1(net5301),
    .A2(_03946_));
 sg13g2_nor3_2 _20838_ (.A(net5360),
    .B(_03834_),
    .C(net5329),
    .Y(_04047_));
 sg13g2_nor3_1 _20839_ (.A(net5292),
    .B(net5327),
    .C(_04047_),
    .Y(_04048_));
 sg13g2_nand2_1 _20840_ (.Y(_04049_),
    .A(_03732_),
    .B(net5330));
 sg13g2_nand2_1 _20841_ (.Y(_04050_),
    .A(net5330),
    .B(net5327));
 sg13g2_nand2b_2 _20842_ (.Y(_04051_),
    .B(_03733_),
    .A_N(net5329));
 sg13g2_nand3_1 _20843_ (.B(_04050_),
    .C(_04051_),
    .A(net5340),
    .Y(_04052_));
 sg13g2_a21oi_1 _20844_ (.A1(net5295),
    .A2(_04052_),
    .Y(_04053_),
    .B1(_04048_));
 sg13g2_nand2_1 _20845_ (.Y(_04054_),
    .A(net5292),
    .B(net5332));
 sg13g2_inv_1 _20846_ (.Y(_04055_),
    .A(net5212));
 sg13g2_o21ai_1 _20847_ (.B1(net5512),
    .Y(_04056_),
    .A1(net5360),
    .A2(_03834_));
 sg13g2_nand2_2 _20848_ (.Y(_04057_),
    .A(net5331),
    .B(_03836_));
 sg13g2_or2_2 _20849_ (.X(_04058_),
    .B(_04056_),
    .A(net5330));
 sg13g2_inv_1 _20850_ (.Y(_04059_),
    .A(_04058_));
 sg13g2_o21ai_1 _20851_ (.B1(_04055_),
    .Y(_04060_),
    .A1(net5327),
    .A2(_04059_));
 sg13g2_nor2_1 _20852_ (.A(net5299),
    .B(net5213),
    .Y(_04061_));
 sg13g2_nor2b_1 _20853_ (.A(_04053_),
    .B_N(net5145),
    .Y(_04062_));
 sg13g2_nor2_1 _20854_ (.A(net5215),
    .B(net5213),
    .Y(_04063_));
 sg13g2_nand2_2 _20855_ (.Y(_04064_),
    .A(net5299),
    .B(_04039_));
 sg13g2_nor2_2 _20856_ (.A(net5337),
    .B(net5327),
    .Y(_04065_));
 sg13g2_and3_1 _20857_ (.X(_04066_),
    .A(net5289),
    .B(_03939_),
    .C(_04065_));
 sg13g2_nand2b_1 _20858_ (.Y(_04067_),
    .B(net5337),
    .A_N(_03538_));
 sg13g2_nor2_1 _20859_ (.A(_03937_),
    .B(net5282),
    .Y(_04068_));
 sg13g2_nor2_1 _20860_ (.A(_04066_),
    .B(_04068_),
    .Y(_04069_));
 sg13g2_nor2_2 _20861_ (.A(net5332),
    .B(net5327),
    .Y(_04070_));
 sg13g2_and2_1 _20862_ (.A(net5331),
    .B(net5328),
    .X(_04071_));
 sg13g2_nand2_2 _20863_ (.Y(_04072_),
    .A(net5331),
    .B(net5329));
 sg13g2_nand3_1 _20864_ (.B(_04070_),
    .C(_04072_),
    .A(net5295),
    .Y(_04073_));
 sg13g2_nor2_1 _20865_ (.A(net5339),
    .B(_03732_),
    .Y(_04074_));
 sg13g2_nand2_1 _20866_ (.Y(_04075_),
    .A(net5334),
    .B(_04071_));
 sg13g2_nand3_1 _20867_ (.B(net5333),
    .C(_04071_),
    .A(net5294),
    .Y(_04076_));
 sg13g2_nand3_1 _20868_ (.B(_04073_),
    .C(_04076_),
    .A(_04069_),
    .Y(_04077_));
 sg13g2_a22oi_1 _20869_ (.Y(_04078_),
    .B1(net5142),
    .B2(_04077_),
    .A2(_04062_),
    .A1(_04060_));
 sg13g2_and2_2 _20870_ (.A(_04046_),
    .B(_04078_),
    .X(_04079_));
 sg13g2_a21oi_2 _20871_ (.B1(net7295),
    .Y(_04080_),
    .A2(_03346_),
    .A1(_03345_));
 sg13g2_nor2_1 _20872_ (.A(_04079_),
    .B(_04080_),
    .Y(_04081_));
 sg13g2_nand2_2 _20873_ (.Y(_04082_),
    .A(_04079_),
    .B(_04080_));
 sg13g2_inv_1 _20874_ (.Y(_04083_),
    .A(_04082_));
 sg13g2_nor3_1 _20875_ (.A(net5408),
    .B(_04081_),
    .C(_04083_),
    .Y(_01157_));
 sg13g2_nand2_2 _20876_ (.Y(_04084_),
    .A(\r_pwm_odd[4] ),
    .B(net5457));
 sg13g2_and3_1 _20877_ (.X(_04085_),
    .A(net5512),
    .B(_03731_),
    .C(_03833_));
 sg13g2_nand2_2 _20878_ (.Y(_04086_),
    .A(_03929_),
    .B(_03940_));
 sg13g2_nand2_1 _20879_ (.Y(_04087_),
    .A(_03836_),
    .B(net5329));
 sg13g2_nand2_1 _20880_ (.Y(_04088_),
    .A(net5328),
    .B(_04056_));
 sg13g2_nand3b_1 _20881_ (.B(_04086_),
    .C(net5281),
    .Y(_04089_),
    .A_N(net5325));
 sg13g2_nand2_1 _20882_ (.Y(_04090_),
    .A(net5291),
    .B(net5338));
 sg13g2_and2_1 _20883_ (.A(net5338),
    .B(_04089_),
    .X(_04091_));
 sg13g2_nor2b_1 _20884_ (.A(_04090_),
    .B_N(_04089_),
    .Y(_04092_));
 sg13g2_nand2_1 _20885_ (.Y(_04093_),
    .A(net5283),
    .B(_04070_));
 sg13g2_and2_1 _20886_ (.A(_04051_),
    .B(_04087_),
    .X(_04094_));
 sg13g2_or2_1 _20887_ (.X(_04095_),
    .B(_04094_),
    .A(net5338));
 sg13g2_a21oi_1 _20888_ (.A1(_04093_),
    .A2(_04095_),
    .Y(_04096_),
    .B1(net5293));
 sg13g2_nand2_1 _20889_ (.Y(_04097_),
    .A(net5333),
    .B(_03836_));
 sg13g2_nand2_1 _20890_ (.Y(_04098_),
    .A(net5336),
    .B(_04056_));
 sg13g2_nor2_1 _20891_ (.A(net5288),
    .B(_04098_),
    .Y(_04099_));
 sg13g2_or3_1 _20892_ (.A(_04092_),
    .B(_04096_),
    .C(_04099_),
    .X(_04100_));
 sg13g2_mux2_2 _20893_ (.A0(_03833_),
    .A1(_03835_),
    .S(net5328),
    .X(_04101_));
 sg13g2_mux2_2 _20894_ (.A0(_03929_),
    .A1(net5328),
    .S(_03836_),
    .X(_04102_));
 sg13g2_nand2_2 _20895_ (.Y(_04103_),
    .A(_03733_),
    .B(_04101_));
 sg13g2_nand2b_1 _20896_ (.Y(_04104_),
    .B(net5300),
    .A_N(net5325));
 sg13g2_nor2b_1 _20897_ (.A(_04104_),
    .B_N(_04103_),
    .Y(_04105_));
 sg13g2_nand2b_2 _20898_ (.Y(_04106_),
    .B(net5332),
    .A_N(_04058_));
 sg13g2_a21oi_1 _20899_ (.A1(net5283),
    .A2(_04070_),
    .Y(_04107_),
    .B1(net5287));
 sg13g2_a221oi_1 _20900_ (.B2(_04107_),
    .C1(net5299),
    .B1(_04106_),
    .A1(net5287),
    .Y(_04108_),
    .A2(_04059_));
 sg13g2_o21ai_1 _20901_ (.B1(net5213),
    .Y(_04109_),
    .A1(_04105_),
    .A2(_04108_));
 sg13g2_o21ai_1 _20902_ (.B1(net5339),
    .Y(_04110_),
    .A1(net5284),
    .A2(_04056_));
 sg13g2_o21ai_1 _20903_ (.B1(net5332),
    .Y(_04111_),
    .A1(_03732_),
    .A2(_04043_));
 sg13g2_a21oi_1 _20904_ (.A1(_04110_),
    .A2(_04111_),
    .Y(_04112_),
    .B1(net5288));
 sg13g2_nor3_1 _20905_ (.A(net5291),
    .B(net5326),
    .C(_04056_),
    .Y(_04113_));
 sg13g2_o21ai_1 _20906_ (.B1(net5144),
    .Y(_04114_),
    .A1(_04112_),
    .A2(_04113_));
 sg13g2_nand2_1 _20907_ (.Y(_04115_),
    .A(_04109_),
    .B(_04114_));
 sg13g2_a21oi_2 _20908_ (.B1(_04115_),
    .Y(_04116_),
    .A2(_04100_),
    .A1(net5143));
 sg13g2_nor2b_1 _20909_ (.A(_04079_),
    .B_N(_04116_),
    .Y(_04117_));
 sg13g2_xnor2_1 _20910_ (.Y(_04118_),
    .A(_04079_),
    .B(_04116_));
 sg13g2_nor2_1 _20911_ (.A(_04084_),
    .B(_04118_),
    .Y(_04119_));
 sg13g2_xor2_1 _20912_ (.B(_04118_),
    .A(_04084_),
    .X(_04120_));
 sg13g2_xnor2_1 _20913_ (.Y(_04121_),
    .A(_04082_),
    .B(_04120_));
 sg13g2_and2_1 _20914_ (.A(net5405),
    .B(_04121_),
    .X(_01158_));
 sg13g2_nand2_2 _20915_ (.Y(_04122_),
    .A(\r_pwm_odd[5] ),
    .B(net5457));
 sg13g2_nand2_2 _20916_ (.Y(_04123_),
    .A(_03732_),
    .B(_04102_));
 sg13g2_and2_1 _20917_ (.A(_04103_),
    .B(_04123_),
    .X(_04124_));
 sg13g2_or2_1 _20918_ (.X(_04125_),
    .B(_04124_),
    .A(net5341));
 sg13g2_a21oi_1 _20919_ (.A1(net5341),
    .A2(_04124_),
    .Y(_04126_),
    .B1(net5297));
 sg13g2_nand2_1 _20920_ (.Y(_04127_),
    .A(_04125_),
    .B(_04126_));
 sg13g2_a21oi_1 _20921_ (.A1(net5286),
    .A2(_04042_),
    .Y(_04128_),
    .B1(net5341));
 sg13g2_a21oi_1 _20922_ (.A1(_03835_),
    .A2(net5330),
    .Y(_04129_),
    .B1(_03940_));
 sg13g2_a21oi_2 _20923_ (.B1(_03836_),
    .Y(_04130_),
    .A2(_03929_),
    .A1(net5360));
 sg13g2_o21ai_1 _20924_ (.B1(net5297),
    .Y(_04131_),
    .A1(net5335),
    .A2(_04130_));
 sg13g2_o21ai_1 _20925_ (.B1(_04127_),
    .Y(_04132_),
    .A1(_04128_),
    .A2(_04131_));
 sg13g2_a21oi_1 _20926_ (.A1(_04057_),
    .A2(_04102_),
    .Y(_04133_),
    .B1(net5342));
 sg13g2_nand2_2 _20927_ (.Y(_04134_),
    .A(net5339),
    .B(net5360));
 sg13g2_nand2b_1 _20928_ (.Y(_04135_),
    .B(_04102_),
    .A_N(_04134_));
 sg13g2_nor2b_1 _20929_ (.A(_04133_),
    .B_N(_04135_),
    .Y(_04136_));
 sg13g2_nor2_1 _20930_ (.A(net5297),
    .B(_04136_),
    .Y(_04137_));
 sg13g2_nand2b_1 _20931_ (.Y(_04138_),
    .B(net5295),
    .A_N(net5325));
 sg13g2_nor2_2 _20932_ (.A(net5339),
    .B(_04085_),
    .Y(_04139_));
 sg13g2_a21oi_1 _20933_ (.A1(net5340),
    .A2(_04041_),
    .Y(_04140_),
    .B1(_04138_));
 sg13g2_o21ai_1 _20934_ (.B1(net5215),
    .Y(_04141_),
    .A1(_04067_),
    .A2(_04086_));
 sg13g2_or3_1 _20935_ (.A(_04137_),
    .B(_04140_),
    .C(_04141_),
    .X(_04142_));
 sg13g2_nand3_1 _20936_ (.B(_04088_),
    .C(_04123_),
    .A(net5302),
    .Y(_04143_));
 sg13g2_and2_1 _20937_ (.A(_04142_),
    .B(_04143_),
    .X(_04144_));
 sg13g2_o21ai_1 _20938_ (.B1(net5342),
    .Y(_04145_),
    .A1(net5331),
    .A2(_04101_));
 sg13g2_nor2_2 _20939_ (.A(_04047_),
    .B(_04145_),
    .Y(_04146_));
 sg13g2_or2_1 _20940_ (.X(_04147_),
    .B(net5328),
    .A(_03634_));
 sg13g2_nand2_1 _20941_ (.Y(_04148_),
    .A(net5296),
    .B(_04147_));
 sg13g2_nand2_1 _20942_ (.Y(_04149_),
    .A(_04049_),
    .B(_04086_));
 sg13g2_nor2_1 _20943_ (.A(net5341),
    .B(_04149_),
    .Y(_04150_));
 sg13g2_nor3_1 _20944_ (.A(net5335),
    .B(_04041_),
    .C(net5325),
    .Y(_04151_));
 sg13g2_nor3_1 _20945_ (.A(net5297),
    .B(_04150_),
    .C(_04151_),
    .Y(_04152_));
 sg13g2_o21ai_1 _20946_ (.B1(net5142),
    .Y(_04153_),
    .A1(_04146_),
    .A2(_04148_));
 sg13g2_nor2_1 _20947_ (.A(_04152_),
    .B(_04153_),
    .Y(_04154_));
 sg13g2_a221oi_1 _20948_ (.B2(_04040_),
    .C1(_04154_),
    .B1(_04144_),
    .A1(net5145),
    .Y(_04155_),
    .A2(_04132_));
 sg13g2_xnor2_1 _20949_ (.Y(_04156_),
    .A(_04117_),
    .B(_04155_));
 sg13g2_nor2_1 _20950_ (.A(_04122_),
    .B(_04156_),
    .Y(_04157_));
 sg13g2_xor2_1 _20951_ (.B(_04156_),
    .A(_04122_),
    .X(_04158_));
 sg13g2_a21oi_2 _20952_ (.B1(_04119_),
    .Y(_04159_),
    .A2(_04120_),
    .A1(_04083_));
 sg13g2_nor2b_1 _20953_ (.A(_04159_),
    .B_N(_04158_),
    .Y(_04160_));
 sg13g2_xor2_1 _20954_ (.B(_04159_),
    .A(_04158_),
    .X(_04161_));
 sg13g2_nor2_1 _20955_ (.A(net5408),
    .B(_04161_),
    .Y(_01159_));
 sg13g2_nand2_2 _20956_ (.Y(_04162_),
    .A(\r_pwm_odd[6] ),
    .B(net5456));
 sg13g2_nor2b_1 _20957_ (.A(_04047_),
    .B_N(_04065_),
    .Y(_04163_));
 sg13g2_a21oi_1 _20958_ (.A1(net5283),
    .A2(_04163_),
    .Y(_04164_),
    .B1(net5296));
 sg13g2_and2_1 _20959_ (.A(_04052_),
    .B(_04164_),
    .X(_04165_));
 sg13g2_nand3_1 _20960_ (.B(_04051_),
    .C(_04070_),
    .A(net5283),
    .Y(_04166_));
 sg13g2_nand2_1 _20961_ (.Y(_04167_),
    .A(net5296),
    .B(_04166_));
 sg13g2_nand2_1 _20962_ (.Y(_04168_),
    .A(net5336),
    .B(_04072_));
 sg13g2_nor2_1 _20963_ (.A(_04041_),
    .B(_04168_),
    .Y(_04169_));
 sg13g2_nor2_1 _20964_ (.A(_04167_),
    .B(_04169_),
    .Y(_04170_));
 sg13g2_o21ai_1 _20965_ (.B1(_03446_),
    .Y(_04171_),
    .A1(_04165_),
    .A2(_04170_));
 sg13g2_nand2_2 _20966_ (.Y(_04172_),
    .A(net5331),
    .B(_03939_));
 sg13g2_and2_1 _20967_ (.A(net5302),
    .B(_04050_),
    .X(_04173_));
 sg13g2_a21oi_1 _20968_ (.A1(_04172_),
    .A2(_04173_),
    .Y(_04174_),
    .B1(_04039_));
 sg13g2_nand2_1 _20969_ (.Y(_04175_),
    .A(_04171_),
    .B(_04174_));
 sg13g2_a21o_1 _20970_ (.A2(_04094_),
    .A1(net5293),
    .B1(_04055_),
    .X(_04176_));
 sg13g2_o21ai_1 _20971_ (.B1(_04176_),
    .Y(_04177_),
    .A1(net5338),
    .A2(_04102_));
 sg13g2_a21oi_2 _20972_ (.B1(net5340),
    .Y(_04178_),
    .A2(_04102_),
    .A1(_03732_));
 sg13g2_nand2_1 _20973_ (.Y(_04179_),
    .A(net5286),
    .B(_04178_));
 sg13g2_nand3_1 _20974_ (.B(_04166_),
    .C(_04179_),
    .A(net5290),
    .Y(_04180_));
 sg13g2_nand3_1 _20975_ (.B(_04177_),
    .C(_04180_),
    .A(net5143),
    .Y(_04181_));
 sg13g2_a21o_1 _20976_ (.A2(_04139_),
    .A1(_04103_),
    .B1(_04167_),
    .X(_04182_));
 sg13g2_nor2_1 _20977_ (.A(net5284),
    .B(net5282),
    .Y(_04183_));
 sg13g2_nand2_1 _20978_ (.Y(_04184_),
    .A(net5283),
    .B(_04183_));
 sg13g2_nor2_2 _20979_ (.A(net5292),
    .B(net5338),
    .Y(_04185_));
 sg13g2_nand2_1 _20980_ (.Y(_04186_),
    .A(_04094_),
    .B(_04185_));
 sg13g2_nand4_1 _20981_ (.B(_04182_),
    .C(_04184_),
    .A(net5144),
    .Y(_04187_),
    .D(_04186_));
 sg13g2_nand3_1 _20982_ (.B(_04181_),
    .C(_04187_),
    .A(_04175_),
    .Y(_04188_));
 sg13g2_a21oi_1 _20983_ (.A1(_04079_),
    .A2(_04116_),
    .Y(_04189_),
    .B1(_04155_));
 sg13g2_nand2_1 _20984_ (.Y(_04190_),
    .A(_04116_),
    .B(_04155_));
 sg13g2_nor2b_1 _20985_ (.A(_04189_),
    .B_N(_04190_),
    .Y(_04191_));
 sg13g2_xnor2_1 _20986_ (.Y(_04192_),
    .A(_04188_),
    .B(_04191_));
 sg13g2_nor2b_1 _20987_ (.A(_04162_),
    .B_N(_04192_),
    .Y(_04193_));
 sg13g2_xnor2_1 _20988_ (.Y(_04194_),
    .A(_04162_),
    .B(_04192_));
 sg13g2_nor2_2 _20989_ (.A(_04157_),
    .B(_04160_),
    .Y(_04195_));
 sg13g2_nor2b_1 _20990_ (.A(_04195_),
    .B_N(_04194_),
    .Y(_04196_));
 sg13g2_xnor2_1 _20991_ (.Y(_04197_),
    .A(_04194_),
    .B(_04195_));
 sg13g2_and2_1 _20992_ (.A(net5405),
    .B(_04197_),
    .X(_01160_));
 sg13g2_nand2_2 _20993_ (.Y(_04198_),
    .A(\r_pwm_odd[7] ),
    .B(net5456));
 sg13g2_nor2_1 _20994_ (.A(net5332),
    .B(_03935_),
    .Y(_04199_));
 sg13g2_nand2b_1 _20995_ (.Y(_04200_),
    .B(_04199_),
    .A_N(_03940_));
 sg13g2_nand2_2 _20996_ (.Y(_04201_),
    .A(net5330),
    .B(net5325));
 sg13g2_a21oi_1 _20997_ (.A1(_03928_),
    .A2(net5325),
    .Y(_04202_),
    .B1(_03940_));
 sg13g2_nand2_1 _20998_ (.Y(_04203_),
    .A(net5332),
    .B(_04202_));
 sg13g2_nand2_1 _20999_ (.Y(_04204_),
    .A(_04200_),
    .B(_04203_));
 sg13g2_nand2_1 _21000_ (.Y(_04205_),
    .A(net5332),
    .B(_04089_));
 sg13g2_nor2_2 _21001_ (.A(net5336),
    .B(_04202_),
    .Y(_04206_));
 sg13g2_nand3b_1 _21002_ (.B(net5291),
    .C(_04205_),
    .Y(_04207_),
    .A_N(_04206_));
 sg13g2_o21ai_1 _21003_ (.B1(_04207_),
    .Y(_04208_),
    .A1(net5291),
    .A2(_04204_));
 sg13g2_nor2_1 _21004_ (.A(_03933_),
    .B(net5326),
    .Y(_04209_));
 sg13g2_and2_1 _21005_ (.A(net5300),
    .B(_04209_),
    .X(_04210_));
 sg13g2_a21oi_1 _21006_ (.A1(net5215),
    .A2(_04208_),
    .Y(_04211_),
    .B1(_04210_));
 sg13g2_nor2_2 _21007_ (.A(net5326),
    .B(_04101_),
    .Y(_04212_));
 sg13g2_a21oi_1 _21008_ (.A1(net5336),
    .A2(_04212_),
    .Y(_04213_),
    .B1(_04206_));
 sg13g2_nor2_1 _21009_ (.A(net5291),
    .B(_04213_),
    .Y(_04214_));
 sg13g2_nor2_1 _21010_ (.A(net5287),
    .B(net5360),
    .Y(_04215_));
 sg13g2_nand3_1 _21011_ (.B(_03932_),
    .C(_04215_),
    .A(net5337),
    .Y(_04216_));
 sg13g2_o21ai_1 _21012_ (.B1(_04216_),
    .Y(_04217_),
    .A1(net5291),
    .A2(_04213_));
 sg13g2_nor2_2 _21013_ (.A(net5327),
    .B(_04041_),
    .Y(_04218_));
 sg13g2_inv_1 _21014_ (.Y(_04219_),
    .A(_04218_));
 sg13g2_nor2b_1 _21015_ (.A(net5212),
    .B_N(net5281),
    .Y(_04220_));
 sg13g2_a21oi_1 _21016_ (.A1(_04218_),
    .A2(_04220_),
    .Y(_04221_),
    .B1(_04217_));
 sg13g2_nor2_1 _21017_ (.A(_04064_),
    .B(_04221_),
    .Y(_04222_));
 sg13g2_nand2_2 _21018_ (.Y(_04223_),
    .A(_03733_),
    .B(_04087_));
 sg13g2_nor2_1 _21019_ (.A(net5282),
    .B(_04223_),
    .Y(_04224_));
 sg13g2_a21oi_1 _21020_ (.A1(_03933_),
    .A2(_04185_),
    .Y(_04225_),
    .B1(_04224_));
 sg13g2_o21ai_1 _21021_ (.B1(net5292),
    .Y(_04226_),
    .A1(_03634_),
    .A2(_04209_));
 sg13g2_o21ai_1 _21022_ (.B1(_04225_),
    .Y(_04227_),
    .A1(_04206_),
    .A2(_04226_));
 sg13g2_a221oi_1 _21023_ (.B2(net5144),
    .C1(_04222_),
    .B1(_04227_),
    .A1(net5213),
    .Y(_04228_),
    .A2(_04211_));
 sg13g2_nor2b_1 _21024_ (.A(_04188_),
    .B_N(_04228_),
    .Y(_04229_));
 sg13g2_xnor2_1 _21025_ (.Y(_04230_),
    .A(_04188_),
    .B(_04228_));
 sg13g2_o21ai_1 _21026_ (.B1(_04190_),
    .Y(_04231_),
    .A1(_04188_),
    .A2(_04189_));
 sg13g2_and2_1 _21027_ (.A(_04230_),
    .B(_04231_),
    .X(_04232_));
 sg13g2_xnor2_1 _21028_ (.Y(_04233_),
    .A(_04230_),
    .B(_04231_));
 sg13g2_xor2_1 _21029_ (.B(_04233_),
    .A(_04198_),
    .X(_04234_));
 sg13g2_nor2_2 _21030_ (.A(_04193_),
    .B(_04196_),
    .Y(_04235_));
 sg13g2_nand2b_1 _21031_ (.Y(_04236_),
    .B(_04234_),
    .A_N(_04235_));
 sg13g2_xor2_1 _21032_ (.B(_04235_),
    .A(_04234_),
    .X(_04237_));
 sg13g2_nor2_1 _21033_ (.A(net5407),
    .B(_04237_),
    .Y(_01161_));
 sg13g2_o21ai_1 _21034_ (.B1(_04236_),
    .Y(_04238_),
    .A1(_04198_),
    .A2(_04233_));
 sg13g2_nand2_1 _21035_ (.Y(_04239_),
    .A(_04134_),
    .B(_04218_));
 sg13g2_o21ai_1 _21036_ (.B1(_04058_),
    .Y(_04240_),
    .A1(_04056_),
    .A2(_04074_));
 sg13g2_a21o_1 _21037_ (.A2(_04240_),
    .A1(net5292),
    .B1(net5300),
    .X(_04241_));
 sg13g2_a21oi_1 _21038_ (.A1(net5287),
    .A2(_04239_),
    .Y(_04242_),
    .B1(_04241_));
 sg13g2_nor2_1 _21039_ (.A(net5215),
    .B(net5326),
    .Y(_04243_));
 sg13g2_o21ai_1 _21040_ (.B1(net5214),
    .Y(_04244_),
    .A1(_04242_),
    .A2(_04243_));
 sg13g2_nor2_1 _21041_ (.A(net5282),
    .B(net5281),
    .Y(_04245_));
 sg13g2_nor2_1 _21042_ (.A(net5337),
    .B(_03933_),
    .Y(_04246_));
 sg13g2_nor3_1 _21043_ (.A(net5287),
    .B(_04219_),
    .C(_04246_),
    .Y(_04247_));
 sg13g2_o21ai_1 _21044_ (.B1(net5144),
    .Y(_04248_),
    .A1(_04245_),
    .A2(_04247_));
 sg13g2_nor2_1 _21045_ (.A(net5292),
    .B(_04240_),
    .Y(_04249_));
 sg13g2_nor2_1 _21046_ (.A(net5212),
    .B(net5281),
    .Y(_04250_));
 sg13g2_o21ai_1 _21047_ (.B1(net5143),
    .Y(_04251_),
    .A1(_04249_),
    .A2(_04250_));
 sg13g2_nand3_1 _21048_ (.B(_04248_),
    .C(_04251_),
    .A(_04244_),
    .Y(_04252_));
 sg13g2_inv_1 _21049_ (.Y(_04253_),
    .A(_04252_));
 sg13g2_xnor2_1 _21050_ (.Y(_04254_),
    .A(_04228_),
    .B(_04252_));
 sg13g2_o21ai_1 _21051_ (.B1(_04254_),
    .Y(_04255_),
    .A1(_04229_),
    .A2(_04232_));
 sg13g2_or3_1 _21052_ (.A(_04229_),
    .B(_04232_),
    .C(_04254_),
    .X(_04256_));
 sg13g2_and2_1 _21053_ (.A(_04255_),
    .B(_04256_),
    .X(_04257_));
 sg13g2_nand2_1 _21054_ (.Y(_04258_),
    .A(_04238_),
    .B(_04257_));
 sg13g2_o21ai_1 _21055_ (.B1(net5403),
    .Y(_04259_),
    .A1(_04238_),
    .A2(_04257_));
 sg13g2_nor2b_1 _21056_ (.A(_04259_),
    .B_N(_04258_),
    .Y(_01162_));
 sg13g2_o21ai_1 _21057_ (.B1(_04253_),
    .Y(_04260_),
    .A1(_04228_),
    .A2(_04232_));
 sg13g2_nand2_1 _21058_ (.Y(_04261_),
    .A(_04252_),
    .B(_04255_));
 sg13g2_and2_1 _21059_ (.A(_04260_),
    .B(_04261_),
    .X(_04262_));
 sg13g2_inv_1 _21060_ (.Y(_04263_),
    .A(_04262_));
 sg13g2_nand3_1 _21061_ (.B(_04257_),
    .C(_04262_),
    .A(_04238_),
    .Y(_04264_));
 sg13g2_nand2_1 _21062_ (.Y(_04265_),
    .A(net5403),
    .B(_04264_));
 sg13g2_a21oi_2 _21063_ (.B1(_04265_),
    .Y(_01163_),
    .A2(_04263_),
    .A1(_04258_));
 sg13g2_a21oi_2 _21064_ (.B1(net5407),
    .Y(_01164_),
    .A2(_04264_),
    .A1(_04260_));
 sg13g2_and3_1 _21065_ (.X(_01165_),
    .A(net2910),
    .B(net5460),
    .C(net5406));
 sg13g2_a21o_1 _21066_ (.A2(_04172_),
    .A1(_04123_),
    .B1(net5333),
    .X(_04266_));
 sg13g2_and2_2 _21067_ (.A(net5302),
    .B(net5290),
    .X(_04267_));
 sg13g2_nand2_2 _21068_ (.Y(_04268_),
    .A(net5299),
    .B(net5288));
 sg13g2_nand2b_2 _21069_ (.Y(_04269_),
    .B(net5325),
    .A_N(net5328));
 sg13g2_nand2_1 _21070_ (.Y(_04270_),
    .A(net5342),
    .B(_04269_));
 sg13g2_nand3_1 _21071_ (.B(_03942_),
    .C(_04270_),
    .A(net5301),
    .Y(_04271_));
 sg13g2_a22oi_1 _21072_ (.Y(_04272_),
    .B1(_04268_),
    .B2(_04271_),
    .A2(_04266_),
    .A1(_03944_));
 sg13g2_nand3_1 _21073_ (.B(_04088_),
    .C(_04269_),
    .A(_04086_),
    .Y(_04273_));
 sg13g2_nor2b_1 _21074_ (.A(_04074_),
    .B_N(_04134_),
    .Y(_04274_));
 sg13g2_a21oi_1 _21075_ (.A1(_04273_),
    .A2(_04274_),
    .Y(_04275_),
    .B1(net5294));
 sg13g2_and4_1 _21076_ (.A(net5294),
    .B(_03938_),
    .C(_04075_),
    .D(_04097_),
    .X(_04276_));
 sg13g2_nor3_1 _21077_ (.A(net5301),
    .B(_04275_),
    .C(_04276_),
    .Y(_04277_));
 sg13g2_o21ai_1 _21078_ (.B1(_04040_),
    .Y(_04278_),
    .A1(_04272_),
    .A2(_04277_));
 sg13g2_nand2_2 _21079_ (.Y(_04279_),
    .A(net5212),
    .B(net5282));
 sg13g2_nand3_1 _21080_ (.B(_04172_),
    .C(_04279_),
    .A(_04123_),
    .Y(_04280_));
 sg13g2_a21o_1 _21081_ (.A2(net5285),
    .A1(_03936_),
    .B1(_04279_),
    .X(_04281_));
 sg13g2_nand3_1 _21082_ (.B(_04280_),
    .C(_04281_),
    .A(net5144),
    .Y(_04282_));
 sg13g2_nor3_1 _21083_ (.A(net5333),
    .B(_04041_),
    .C(net5284),
    .Y(_04283_));
 sg13g2_a21oi_1 _21084_ (.A1(_04058_),
    .A2(net5281),
    .Y(_04284_),
    .B1(net5342));
 sg13g2_o21ai_1 _21085_ (.B1(net5294),
    .Y(_04285_),
    .A1(_04283_),
    .A2(_04284_));
 sg13g2_a21o_1 _21086_ (.A2(_04285_),
    .A1(_04069_),
    .B1(_04064_),
    .X(_04286_));
 sg13g2_nand3_1 _21087_ (.B(_04282_),
    .C(_04286_),
    .A(_04278_),
    .Y(_04287_));
 sg13g2_nand2b_1 _21088_ (.Y(_04288_),
    .B(net5460),
    .A_N(net7269));
 sg13g2_nand2_1 _21089_ (.Y(_04289_),
    .A(_04287_),
    .B(_04288_));
 sg13g2_nor2_2 _21090_ (.A(_04287_),
    .B(_04288_),
    .Y(_04290_));
 sg13g2_inv_1 _21091_ (.Y(_04291_),
    .A(_04290_));
 sg13g2_and3_1 _21092_ (.X(_01166_),
    .A(_03350_),
    .B(_04289_),
    .C(_04291_));
 sg13g2_nand2_1 _21093_ (.Y(_04292_),
    .A(\g_pwm_odd[4] ),
    .B(net5459));
 sg13g2_nor3_1 _21094_ (.A(net5333),
    .B(_03732_),
    .C(_04102_),
    .Y(_04293_));
 sg13g2_a21oi_1 _21095_ (.A1(_03634_),
    .A2(_04085_),
    .Y(_04294_),
    .B1(_04293_));
 sg13g2_nand3_1 _21096_ (.B(_04072_),
    .C(_04101_),
    .A(net5333),
    .Y(_04295_));
 sg13g2_a21oi_1 _21097_ (.A1(_04294_),
    .A2(_04295_),
    .Y(_04296_),
    .B1(net5289));
 sg13g2_o21ai_1 _21098_ (.B1(net5142),
    .Y(_04297_),
    .A1(_04096_),
    .A2(_04296_));
 sg13g2_nor2b_1 _21099_ (.A(_03940_),
    .B_N(_04269_),
    .Y(_04298_));
 sg13g2_or2_1 _21100_ (.X(_04299_),
    .B(_04298_),
    .A(_04279_));
 sg13g2_nand2_1 _21101_ (.Y(_04300_),
    .A(_04130_),
    .B(_04279_));
 sg13g2_a21oi_1 _21102_ (.A1(net5342),
    .A2(_04129_),
    .Y(_04301_),
    .B1(net5295));
 sg13g2_o21ai_1 _21103_ (.B1(net5297),
    .Y(_04302_),
    .A1(net5341),
    .A2(_04130_));
 sg13g2_nand3_1 _21104_ (.B(_04299_),
    .C(_04300_),
    .A(net5145),
    .Y(_04303_));
 sg13g2_nand2_1 _21105_ (.Y(_04304_),
    .A(_04106_),
    .B(_04301_));
 sg13g2_o21ai_1 _21106_ (.B1(net5301),
    .Y(_04305_),
    .A1(_03931_),
    .A2(_04134_));
 sg13g2_nor2b_1 _21107_ (.A(_04305_),
    .B_N(_04106_),
    .Y(_04306_));
 sg13g2_o21ai_1 _21108_ (.B1(_04304_),
    .Y(_04307_),
    .A1(_04267_),
    .A2(_04306_));
 sg13g2_a21oi_1 _21109_ (.A1(net5342),
    .A2(_04059_),
    .Y(_04308_),
    .B1(_04133_));
 sg13g2_nand2_1 _21110_ (.Y(_04309_),
    .A(_03929_),
    .B(_04097_));
 sg13g2_nor2_1 _21111_ (.A(_03538_),
    .B(net5331),
    .Y(_04310_));
 sg13g2_a21oi_1 _21112_ (.A1(_04309_),
    .A2(_04310_),
    .Y(_04311_),
    .B1(net5301));
 sg13g2_o21ai_1 _21113_ (.B1(_04311_),
    .Y(_04312_),
    .A1(net5289),
    .A2(_04308_));
 sg13g2_nand3_1 _21114_ (.B(_04307_),
    .C(_04312_),
    .A(net5214),
    .Y(_04313_));
 sg13g2_and3_2 _21115_ (.X(_04314_),
    .A(_04297_),
    .B(_04303_),
    .C(_04313_));
 sg13g2_nand2_1 _21116_ (.Y(_04315_),
    .A(_04287_),
    .B(_04314_));
 sg13g2_nor2b_1 _21117_ (.A(_04287_),
    .B_N(_04314_),
    .Y(_04316_));
 sg13g2_xnor2_1 _21118_ (.Y(_04317_),
    .A(_04287_),
    .B(_04314_));
 sg13g2_nand2b_1 _21119_ (.Y(_04318_),
    .B(_04317_),
    .A_N(_04292_));
 sg13g2_xor2_1 _21120_ (.B(_04317_),
    .A(_04292_),
    .X(_04319_));
 sg13g2_xnor2_1 _21121_ (.Y(_04320_),
    .A(_04290_),
    .B(_04319_));
 sg13g2_and2_1 _21122_ (.A(net5406),
    .B(_04320_),
    .X(_01167_));
 sg13g2_nand2_2 _21123_ (.Y(_04321_),
    .A(\g_pwm_odd[5] ),
    .B(net5459));
 sg13g2_nand2b_1 _21124_ (.Y(_04322_),
    .B(_04173_),
    .A_N(_04139_));
 sg13g2_a21oi_1 _21125_ (.A1(_04268_),
    .A2(_04322_),
    .Y(_04323_),
    .B1(_04137_));
 sg13g2_nor3_1 _21126_ (.A(net5295),
    .B(_03931_),
    .C(_04218_),
    .Y(_04324_));
 sg13g2_a22oi_1 _21127_ (.Y(_04325_),
    .B1(_04139_),
    .B2(_03932_),
    .A2(_04138_),
    .A1(net5212));
 sg13g2_or2_1 _21128_ (.X(_04326_),
    .B(_04325_),
    .A(net5301));
 sg13g2_a21oi_1 _21129_ (.A1(_04097_),
    .A2(_04324_),
    .Y(_04327_),
    .B1(_04326_));
 sg13g2_o21ai_1 _21130_ (.B1(net5214),
    .Y(_04328_),
    .A1(_04323_),
    .A2(_04327_));
 sg13g2_o21ai_1 _21131_ (.B1(_04057_),
    .Y(_04329_),
    .A1(_03931_),
    .A2(_04218_));
 sg13g2_nand2b_1 _21132_ (.Y(_04330_),
    .B(_04329_),
    .A_N(_04279_));
 sg13g2_o21ai_1 _21133_ (.B1(_04279_),
    .Y(_04331_),
    .A1(net5284),
    .A2(_04056_));
 sg13g2_nand3_1 _21134_ (.B(_04330_),
    .C(_04331_),
    .A(net5145),
    .Y(_04332_));
 sg13g2_a21oi_1 _21135_ (.A1(net5340),
    .A2(_04149_),
    .Y(_04333_),
    .B1(_04302_));
 sg13g2_o21ai_1 _21136_ (.B1(net5142),
    .Y(_04334_),
    .A1(_04152_),
    .A2(_04333_));
 sg13g2_nand3_1 _21137_ (.B(_04332_),
    .C(_04334_),
    .A(_04328_),
    .Y(_04335_));
 sg13g2_xor2_1 _21138_ (.B(_04335_),
    .A(_04315_),
    .X(_04336_));
 sg13g2_xnor2_1 _21139_ (.Y(_04337_),
    .A(_04321_),
    .B(_04336_));
 sg13g2_o21ai_1 _21140_ (.B1(_04318_),
    .Y(_04338_),
    .A1(_04291_),
    .A2(_04319_));
 sg13g2_nand2b_1 _21141_ (.Y(_04339_),
    .B(_04338_),
    .A_N(_04337_));
 sg13g2_xor2_1 _21142_ (.B(_04338_),
    .A(_04337_),
    .X(_04340_));
 sg13g2_nor2_1 _21143_ (.A(net5410),
    .B(_04340_),
    .Y(_01168_));
 sg13g2_nand2_2 _21144_ (.Y(_04341_),
    .A(\g_pwm_odd[6] ),
    .B(net5461));
 sg13g2_nor2b_1 _21145_ (.A(net5284),
    .B_N(_04051_),
    .Y(_04342_));
 sg13g2_nor2_1 _21146_ (.A(net5335),
    .B(_04342_),
    .Y(_04343_));
 sg13g2_nor3_1 _21147_ (.A(net5290),
    .B(_04169_),
    .C(_04343_),
    .Y(_04344_));
 sg13g2_a21o_1 _21148_ (.A2(_04042_),
    .A1(net5340),
    .B1(_04178_),
    .X(_04345_));
 sg13g2_nand3_1 _21149_ (.B(_04072_),
    .C(_04345_),
    .A(net5297),
    .Y(_04346_));
 sg13g2_o21ai_1 _21150_ (.B1(_04346_),
    .Y(_04347_),
    .A1(net5296),
    .A2(_04342_));
 sg13g2_nor3_1 _21151_ (.A(_03446_),
    .B(_04165_),
    .C(_04344_),
    .Y(_04348_));
 sg13g2_a21oi_1 _21152_ (.A1(net5215),
    .A2(_04347_),
    .Y(_04349_),
    .B1(_04348_));
 sg13g2_nor2_1 _21153_ (.A(_04039_),
    .B(_04349_),
    .Y(_04350_));
 sg13g2_nor2b_1 _21154_ (.A(_04124_),
    .B_N(_04279_),
    .Y(_04351_));
 sg13g2_o21ai_1 _21155_ (.B1(net5145),
    .Y(_04352_),
    .A1(_04273_),
    .A2(_04279_));
 sg13g2_a21oi_1 _21156_ (.A1(_04051_),
    .A2(_04070_),
    .Y(_04353_),
    .B1(net5290));
 sg13g2_nand2_1 _21157_ (.Y(_04354_),
    .A(_04125_),
    .B(_04353_));
 sg13g2_nand3_1 _21158_ (.B(_04180_),
    .C(_04354_),
    .A(net5142),
    .Y(_04355_));
 sg13g2_o21ai_1 _21159_ (.B1(_04355_),
    .Y(_04356_),
    .A1(_04351_),
    .A2(_04352_));
 sg13g2_or2_2 _21160_ (.X(_04357_),
    .B(_04356_),
    .A(_04350_));
 sg13g2_nand2_1 _21161_ (.Y(_04358_),
    .A(_04314_),
    .B(_04335_));
 sg13g2_nor2_1 _21162_ (.A(_04316_),
    .B(_04335_),
    .Y(_04359_));
 sg13g2_a21oi_1 _21163_ (.A1(_04314_),
    .A2(_04335_),
    .Y(_04360_),
    .B1(_04359_));
 sg13g2_xnor2_1 _21164_ (.Y(_04361_),
    .A(_04357_),
    .B(_04360_));
 sg13g2_inv_1 _21165_ (.Y(_04362_),
    .A(_04361_));
 sg13g2_nor2_1 _21166_ (.A(_04341_),
    .B(_04362_),
    .Y(_04363_));
 sg13g2_xnor2_1 _21167_ (.Y(_04364_),
    .A(_04341_),
    .B(_04361_));
 sg13g2_o21ai_1 _21168_ (.B1(_04339_),
    .Y(_04365_),
    .A1(_04321_),
    .A2(_04336_));
 sg13g2_xnor2_1 _21169_ (.Y(_04366_),
    .A(_04364_),
    .B(_04365_));
 sg13g2_nor2_1 _21170_ (.A(net5409),
    .B(_04366_),
    .Y(_01169_));
 sg13g2_a221oi_1 _21171_ (.B2(_04090_),
    .C1(net5299),
    .B1(_04212_),
    .A1(net5291),
    .Y(_04367_),
    .A2(_04091_));
 sg13g2_nand2_1 _21172_ (.Y(_04368_),
    .A(net5338),
    .B(_04212_));
 sg13g2_and2_2 _21173_ (.A(net5299),
    .B(net5291),
    .X(_04369_));
 sg13g2_nand3_1 _21174_ (.B(_04368_),
    .C(_04369_),
    .A(_04205_),
    .Y(_04370_));
 sg13g2_o21ai_1 _21175_ (.B1(net5213),
    .Y(_04371_),
    .A1(_04204_),
    .A2(_04268_));
 sg13g2_nor2_1 _21176_ (.A(_04367_),
    .B(_04371_),
    .Y(_04372_));
 sg13g2_nand2b_1 _21177_ (.Y(_04373_),
    .B(_04147_),
    .A_N(_03940_));
 sg13g2_nand2b_1 _21178_ (.Y(_04374_),
    .B(_04373_),
    .A_N(_04104_));
 sg13g2_a21oi_1 _21179_ (.A1(_04268_),
    .A2(_04374_),
    .Y(_04375_),
    .B1(_04214_));
 sg13g2_a21oi_1 _21180_ (.A1(_04086_),
    .A2(_04201_),
    .Y(_04376_),
    .B1(net5299));
 sg13g2_nor3_1 _21181_ (.A(net5213),
    .B(_04375_),
    .C(_04376_),
    .Y(_04377_));
 sg13g2_a21o_2 _21182_ (.A2(_04372_),
    .A1(_04370_),
    .B1(_04377_),
    .X(_04378_));
 sg13g2_nor2_1 _21183_ (.A(_04357_),
    .B(_04378_),
    .Y(_04379_));
 sg13g2_xor2_1 _21184_ (.B(_04378_),
    .A(_04357_),
    .X(_04380_));
 sg13g2_o21ai_1 _21185_ (.B1(_04358_),
    .Y(_04381_),
    .A1(_04357_),
    .A2(_04359_));
 sg13g2_nand2_1 _21186_ (.Y(_04382_),
    .A(_04380_),
    .B(_04381_));
 sg13g2_xnor2_1 _21187_ (.Y(_04383_),
    .A(_04380_),
    .B(_04381_));
 sg13g2_nand2_1 _21188_ (.Y(_04384_),
    .A(\g_pwm_odd[7] ),
    .B(net5462));
 sg13g2_or2_1 _21189_ (.X(_04385_),
    .B(_04384_),
    .A(_04383_));
 sg13g2_xnor2_1 _21190_ (.Y(_04386_),
    .A(_04383_),
    .B(_04384_));
 sg13g2_a21oi_2 _21191_ (.B1(_04363_),
    .Y(_04387_),
    .A2(_04365_),
    .A1(_04364_));
 sg13g2_xnor2_1 _21192_ (.Y(_04388_),
    .A(_04386_),
    .B(_04387_));
 sg13g2_nor2_1 _21193_ (.A(net5410),
    .B(_04388_),
    .Y(_01170_));
 sg13g2_o21ai_1 _21194_ (.B1(_04385_),
    .Y(_04389_),
    .A1(_04386_),
    .A2(_04387_));
 sg13g2_a21oi_1 _21195_ (.A1(_04380_),
    .A2(_04381_),
    .Y(_04390_),
    .B1(_04379_));
 sg13g2_nor3_1 _21196_ (.A(_04064_),
    .B(_04215_),
    .C(_04249_),
    .Y(_04391_));
 sg13g2_nand2_1 _21197_ (.Y(_04392_),
    .A(_03933_),
    .B(_04268_));
 sg13g2_o21ai_1 _21198_ (.B1(_04392_),
    .Y(_04393_),
    .A1(_04239_),
    .A2(_04268_));
 sg13g2_a21oi_1 _21199_ (.A1(net5144),
    .A2(_04219_),
    .Y(_04394_),
    .B1(_04391_));
 sg13g2_o21ai_1 _21200_ (.B1(_04394_),
    .Y(_04395_),
    .A1(_04039_),
    .A2(_04393_));
 sg13g2_xor2_1 _21201_ (.B(_04395_),
    .A(_04378_),
    .X(_04396_));
 sg13g2_nor2_1 _21202_ (.A(_04390_),
    .B(_04396_),
    .Y(_04397_));
 sg13g2_xor2_1 _21203_ (.B(_04396_),
    .A(_04390_),
    .X(_04398_));
 sg13g2_nand2_1 _21204_ (.Y(_04399_),
    .A(_04389_),
    .B(_04398_));
 sg13g2_o21ai_1 _21205_ (.B1(net5404),
    .Y(_04400_),
    .A1(_04389_),
    .A2(_04398_));
 sg13g2_nor2b_1 _21206_ (.A(_04400_),
    .B_N(_04399_),
    .Y(_01171_));
 sg13g2_nand2_1 _21207_ (.Y(_04401_),
    .A(_04378_),
    .B(_04382_));
 sg13g2_nand2_2 _21208_ (.Y(_04402_),
    .A(_04395_),
    .B(_04401_));
 sg13g2_o21ai_1 _21209_ (.B1(_04402_),
    .Y(_04403_),
    .A1(_04395_),
    .A2(_04397_));
 sg13g2_or2_1 _21210_ (.X(_04404_),
    .B(_04403_),
    .A(_04399_));
 sg13g2_nand2_1 _21211_ (.Y(_04405_),
    .A(net5405),
    .B(_04404_));
 sg13g2_a21oi_2 _21212_ (.B1(_04405_),
    .Y(_01172_),
    .A2(_04403_),
    .A1(_04399_));
 sg13g2_a21oi_2 _21213_ (.B1(net5408),
    .Y(_01173_),
    .A2(_04404_),
    .A1(_04402_));
 sg13g2_nand2_1 _21214_ (.Y(_04406_),
    .A(net7314),
    .B(net5459));
 sg13g2_nor3_2 _21215_ (.A(_04054_),
    .B(_04064_),
    .C(_04201_),
    .Y(_04407_));
 sg13g2_nand2_1 _21216_ (.Y(_04408_),
    .A(\b_pwm_odd[1] ),
    .B(net5459));
 sg13g2_nand2_1 _21217_ (.Y(_04409_),
    .A(_04407_),
    .B(_04408_));
 sg13g2_xnor2_1 _21218_ (.Y(_04410_),
    .A(_04406_),
    .B(_04409_));
 sg13g2_nor2_1 _21219_ (.A(net5409),
    .B(net7315),
    .Y(_01174_));
 sg13g2_a221oi_1 _21220_ (.B2(_03937_),
    .C1(_04283_),
    .B1(net5333),
    .A1(net5512),
    .Y(_04411_),
    .A2(_03538_));
 sg13g2_a221oi_1 _21221_ (.B2(_04223_),
    .C1(net5289),
    .B1(_04178_),
    .A1(_04058_),
    .Y(_04412_),
    .A2(_04070_));
 sg13g2_nor3_1 _21222_ (.A(net5301),
    .B(_04411_),
    .C(_04412_),
    .Y(_04413_));
 sg13g2_o21ai_1 _21223_ (.B1(_04267_),
    .Y(_04414_),
    .A1(_04163_),
    .A2(_04293_));
 sg13g2_nand2_1 _21224_ (.Y(_04415_),
    .A(_04052_),
    .B(_04369_));
 sg13g2_o21ai_1 _21225_ (.B1(_04414_),
    .Y(_04416_),
    .A1(_04284_),
    .A2(_04415_));
 sg13g2_o21ai_1 _21226_ (.B1(net5214),
    .Y(_04417_),
    .A1(_04413_),
    .A2(_04416_));
 sg13g2_a21oi_1 _21227_ (.A1(_04051_),
    .A2(_04139_),
    .Y(_04418_),
    .B1(net5289));
 sg13g2_a21oi_1 _21228_ (.A1(_04145_),
    .A2(_04418_),
    .Y(_04419_),
    .B1(_04301_));
 sg13g2_or2_1 _21229_ (.X(_04420_),
    .B(_04419_),
    .A(_04066_));
 sg13g2_nor2_1 _21230_ (.A(net5294),
    .B(_03942_),
    .Y(_04421_));
 sg13g2_a21oi_1 _21231_ (.A1(net5331),
    .A2(_03939_),
    .Y(_04422_),
    .B1(net5282));
 sg13g2_o21ai_1 _21232_ (.B1(_04073_),
    .Y(_04423_),
    .A1(net5212),
    .A2(_04172_));
 sg13g2_or3_1 _21233_ (.A(_04421_),
    .B(_04422_),
    .C(_04423_),
    .X(_04424_));
 sg13g2_a22oi_1 _21234_ (.Y(_04425_),
    .B1(_04424_),
    .B2(net5145),
    .A2(_04420_),
    .A1(net5142));
 sg13g2_nand2_2 _21235_ (.Y(_04426_),
    .A(_04417_),
    .B(_04425_));
 sg13g2_nand2_1 _21236_ (.Y(_04427_),
    .A(\b_pwm_odd[3] ),
    .B(net5461));
 sg13g2_nand2_1 _21237_ (.Y(_04428_),
    .A(_04426_),
    .B(_04427_));
 sg13g2_xor2_1 _21238_ (.B(_04427_),
    .A(_04426_),
    .X(_04429_));
 sg13g2_o21ai_1 _21239_ (.B1(net5459),
    .Y(_04430_),
    .A1(\b_pwm_odd[2] ),
    .A2(net7375));
 sg13g2_nor2b_1 _21240_ (.A(_04430_),
    .B_N(_04407_),
    .Y(_04431_));
 sg13g2_nand2_1 _21241_ (.Y(_04432_),
    .A(_04429_),
    .B(_04431_));
 sg13g2_xnor2_1 _21242_ (.Y(_04433_),
    .A(_04429_),
    .B(_04431_));
 sg13g2_nor2_1 _21243_ (.A(net5409),
    .B(_04433_),
    .Y(_01175_));
 sg13g2_nand2_1 _21244_ (.Y(_04434_),
    .A(\b_pwm_odd[4] ),
    .B(net5461));
 sg13g2_o21ai_1 _21245_ (.B1(net5293),
    .Y(_04435_),
    .A1(net5339),
    .A2(_04103_));
 sg13g2_o21ai_1 _21246_ (.B1(net5340),
    .Y(_04436_),
    .A1(_03732_),
    .A2(net5284));
 sg13g2_nand2_1 _21247_ (.Y(_04437_),
    .A(net5290),
    .B(_04436_));
 sg13g2_a21oi_1 _21248_ (.A1(net5335),
    .A2(_04298_),
    .Y(_04438_),
    .B1(_04437_));
 sg13g2_nor2_1 _21249_ (.A(net5302),
    .B(_04438_),
    .Y(_04439_));
 sg13g2_o21ai_1 _21250_ (.B1(_04439_),
    .Y(_04440_),
    .A1(_04091_),
    .A2(_04435_));
 sg13g2_nand2b_1 _21251_ (.Y(_04441_),
    .B(_04095_),
    .A_N(_04070_));
 sg13g2_nand3_1 _21252_ (.B(_04051_),
    .C(_04201_),
    .A(net5338),
    .Y(_04442_));
 sg13g2_nand2_1 _21253_ (.Y(_04443_),
    .A(_04098_),
    .B(_04442_));
 sg13g2_a221oi_1 _21254_ (.B2(_04369_),
    .C1(net5214),
    .B1(_04443_),
    .A1(_04267_),
    .Y(_04444_),
    .A2(_04441_));
 sg13g2_nand3_1 _21255_ (.B(_04106_),
    .C(_04294_),
    .A(net5289),
    .Y(_04445_));
 sg13g2_nand3_1 _21256_ (.B(_04072_),
    .C(_04201_),
    .A(net5335),
    .Y(_04446_));
 sg13g2_nand3_1 _21257_ (.B(_04436_),
    .C(_04446_),
    .A(net5296),
    .Y(_04447_));
 sg13g2_a21oi_1 _21258_ (.A1(_04445_),
    .A2(_04447_),
    .Y(_04448_),
    .B1(net5302));
 sg13g2_nand2_1 _21259_ (.Y(_04449_),
    .A(_04110_),
    .B(_04369_));
 sg13g2_a21oi_1 _21260_ (.A1(net5286),
    .A2(_04139_),
    .Y(_04450_),
    .B1(_04449_));
 sg13g2_a22oi_1 _21261_ (.Y(_04451_),
    .B1(_04057_),
    .B2(_04065_),
    .A2(_04047_),
    .A1(net5337));
 sg13g2_o21ai_1 _21262_ (.B1(net5213),
    .Y(_04452_),
    .A1(_04268_),
    .A2(_04451_));
 sg13g2_nor3_1 _21263_ (.A(_04448_),
    .B(_04450_),
    .C(_04452_),
    .Y(_04453_));
 sg13g2_a21oi_2 _21264_ (.B1(_04453_),
    .Y(_04454_),
    .A2(_04444_),
    .A1(_04440_));
 sg13g2_a21o_1 _21265_ (.A2(_04425_),
    .A1(_04417_),
    .B1(_04454_),
    .X(_04455_));
 sg13g2_xnor2_1 _21266_ (.Y(_04456_),
    .A(_04426_),
    .B(_04454_));
 sg13g2_nor2_1 _21267_ (.A(_04434_),
    .B(_04456_),
    .Y(_04457_));
 sg13g2_nand2_1 _21268_ (.Y(_04458_),
    .A(_04434_),
    .B(_04456_));
 sg13g2_nand2b_1 _21269_ (.Y(_04459_),
    .B(_04458_),
    .A_N(_04457_));
 sg13g2_o21ai_1 _21270_ (.B1(_04432_),
    .Y(_04460_),
    .A1(_04426_),
    .A2(_04427_));
 sg13g2_xor2_1 _21271_ (.B(_04460_),
    .A(_04459_),
    .X(_04461_));
 sg13g2_nor2_1 _21272_ (.A(net5409),
    .B(_04461_),
    .Y(_01176_));
 sg13g2_nand2_2 _21273_ (.Y(_04462_),
    .A(\b_pwm_odd[5] ),
    .B(net5458));
 sg13g2_nand3b_1 _21274_ (.B(net5296),
    .C(_04135_),
    .Y(_04463_),
    .A_N(_04150_));
 sg13g2_nand3_1 _21275_ (.B(net5285),
    .C(net5283),
    .A(net5340),
    .Y(_04464_));
 sg13g2_nand3_1 _21276_ (.B(_04125_),
    .C(_04464_),
    .A(net5289),
    .Y(_04465_));
 sg13g2_nand3_1 _21277_ (.B(_04463_),
    .C(_04465_),
    .A(net5302),
    .Y(_04466_));
 sg13g2_o21ai_1 _21278_ (.B1(net5281),
    .Y(_04467_),
    .A1(net5334),
    .A2(_04058_));
 sg13g2_a21oi_1 _21279_ (.A1(net5283),
    .A2(_04086_),
    .Y(_04468_),
    .B1(net5341));
 sg13g2_o21ai_1 _21280_ (.B1(net5294),
    .Y(_04469_),
    .A1(_04467_),
    .A2(_04468_));
 sg13g2_a21oi_1 _21281_ (.A1(net5281),
    .A2(_04123_),
    .Y(_04470_),
    .B1(net5282));
 sg13g2_a21oi_1 _21282_ (.A1(net5289),
    .A2(_04133_),
    .Y(_04471_),
    .B1(_04470_));
 sg13g2_nand3_1 _21283_ (.B(_04469_),
    .C(_04471_),
    .A(net5215),
    .Y(_04472_));
 sg13g2_a21oi_1 _21284_ (.A1(_04466_),
    .A2(_04472_),
    .Y(_04473_),
    .B1(_04039_));
 sg13g2_a21oi_1 _21285_ (.A1(net5286),
    .A2(net5283),
    .Y(_04474_),
    .B1(net5212));
 sg13g2_a21oi_1 _21286_ (.A1(net5285),
    .A2(_04042_),
    .Y(_04475_),
    .B1(net5282));
 sg13g2_a221oi_1 _21287_ (.B2(_04329_),
    .C1(_04475_),
    .B1(_04185_),
    .A1(net5297),
    .Y(_04476_),
    .A2(_04146_));
 sg13g2_nand2b_1 _21288_ (.Y(_04477_),
    .B(_04476_),
    .A_N(_04474_));
 sg13g2_nor2_1 _21289_ (.A(_04071_),
    .B(_04145_),
    .Y(_04478_));
 sg13g2_nor2_1 _21290_ (.A(_04468_),
    .B(_04478_),
    .Y(_04479_));
 sg13g2_a221oi_1 _21291_ (.B2(_04267_),
    .C1(net5214),
    .B1(_04479_),
    .A1(net5215),
    .Y(_04480_),
    .A2(_04477_));
 sg13g2_nand4_1 _21292_ (.B(_04050_),
    .C(_04086_),
    .A(net5340),
    .Y(_04481_),
    .D(net5281));
 sg13g2_nand4_1 _21293_ (.B(net5142),
    .C(_04147_),
    .A(net5296),
    .Y(_04482_),
    .D(_04481_));
 sg13g2_o21ai_1 _21294_ (.B1(_04482_),
    .Y(_04483_),
    .A1(_04473_),
    .A2(_04480_));
 sg13g2_inv_1 _21295_ (.Y(_04484_),
    .A(_04483_));
 sg13g2_xnor2_1 _21296_ (.Y(_04485_),
    .A(_04455_),
    .B(_04483_));
 sg13g2_xor2_1 _21297_ (.B(_04485_),
    .A(_04462_),
    .X(_04486_));
 sg13g2_a21oi_2 _21298_ (.B1(_04457_),
    .Y(_04487_),
    .A2(_04460_),
    .A1(_04458_));
 sg13g2_nand2b_1 _21299_ (.Y(_04488_),
    .B(_04486_),
    .A_N(_04487_));
 sg13g2_xor2_1 _21300_ (.B(_04487_),
    .A(_04486_),
    .X(_04489_));
 sg13g2_nor2_1 _21301_ (.A(net5410),
    .B(_04489_),
    .Y(_01177_));
 sg13g2_nand2_2 _21302_ (.Y(_04490_),
    .A(\b_pwm_odd[6] ),
    .B(net5458));
 sg13g2_a21oi_2 _21303_ (.B1(_04454_),
    .Y(_04491_),
    .A2(_04483_),
    .A1(_04426_));
 sg13g2_a21oi_1 _21304_ (.A1(net5285),
    .A2(_04139_),
    .Y(_04492_),
    .B1(net5290));
 sg13g2_nand2_1 _21305_ (.Y(_04493_),
    .A(net5285),
    .B(_04151_));
 sg13g2_a221oi_1 _21306_ (.B2(_04164_),
    .C1(net5302),
    .B1(_04493_),
    .A1(_04266_),
    .Y(_04494_),
    .A2(_04492_));
 sg13g2_o21ai_1 _21307_ (.B1(net5338),
    .Y(_04495_),
    .A1(net5284),
    .A2(net5325));
 sg13g2_a21oi_1 _21308_ (.A1(_04095_),
    .A2(_04495_),
    .Y(_04496_),
    .B1(_04268_));
 sg13g2_nand2_1 _21309_ (.Y(_04497_),
    .A(_04072_),
    .B(_04139_));
 sg13g2_nand3_1 _21310_ (.B(_04369_),
    .C(_04497_),
    .A(_04166_),
    .Y(_04498_));
 sg13g2_nand2b_1 _21311_ (.Y(_04499_),
    .B(_04498_),
    .A_N(_04496_));
 sg13g2_o21ai_1 _21312_ (.B1(net5214),
    .Y(_04500_),
    .A1(_04494_),
    .A2(_04499_));
 sg13g2_nand3_1 _21313_ (.B(_04179_),
    .C(_04200_),
    .A(net5290),
    .Y(_04501_));
 sg13g2_nand3_1 _21314_ (.B(net5285),
    .C(_04269_),
    .A(net5342),
    .Y(_04502_));
 sg13g2_nand3_1 _21315_ (.B(_04097_),
    .C(_04502_),
    .A(net5295),
    .Y(_04503_));
 sg13g2_nand3_1 _21316_ (.B(_04501_),
    .C(_04503_),
    .A(net5142),
    .Y(_04504_));
 sg13g2_a21o_1 _21317_ (.A2(_04273_),
    .A1(net5335),
    .B1(_04146_),
    .X(_04505_));
 sg13g2_o21ai_1 _21318_ (.B1(_04176_),
    .Y(_04506_),
    .A1(_03834_),
    .A2(_04168_));
 sg13g2_and2_1 _21319_ (.A(net5145),
    .B(_04506_),
    .X(_04507_));
 sg13g2_o21ai_1 _21320_ (.B1(_04507_),
    .Y(_04508_),
    .A1(net5296),
    .A2(_04505_));
 sg13g2_and3_2 _21321_ (.X(_04509_),
    .A(_04500_),
    .B(_04504_),
    .C(_04508_));
 sg13g2_nor2_1 _21322_ (.A(_04484_),
    .B(_04509_),
    .Y(_04510_));
 sg13g2_xnor2_1 _21323_ (.Y(_04511_),
    .A(_04483_),
    .B(_04509_));
 sg13g2_xnor2_1 _21324_ (.Y(_04512_),
    .A(_04491_),
    .B(_04511_));
 sg13g2_nor2_1 _21325_ (.A(_04490_),
    .B(_04512_),
    .Y(_04513_));
 sg13g2_xor2_1 _21326_ (.B(_04512_),
    .A(_04490_),
    .X(_04514_));
 sg13g2_o21ai_1 _21327_ (.B1(_04488_),
    .Y(_04515_),
    .A1(_04462_),
    .A2(_04485_));
 sg13g2_xnor2_1 _21328_ (.Y(_04516_),
    .A(_04514_),
    .B(_04515_));
 sg13g2_nor2_1 _21329_ (.A(net5410),
    .B(_04516_),
    .Y(_01178_));
 sg13g2_nand2_1 _21330_ (.Y(_04517_),
    .A(\b_pwm_odd[7] ),
    .B(net5458));
 sg13g2_o21ai_1 _21331_ (.B1(net5337),
    .Y(_04518_),
    .A1(_03933_),
    .A2(net5326));
 sg13g2_nand3_1 _21332_ (.B(_04203_),
    .C(_04518_),
    .A(net5287),
    .Y(_04519_));
 sg13g2_nand2b_1 _21333_ (.Y(_04520_),
    .B(_03938_),
    .A_N(_04226_));
 sg13g2_a21oi_1 _21334_ (.A1(_04519_),
    .A2(_04520_),
    .Y(_04521_),
    .B1(net5300));
 sg13g2_a21oi_1 _21335_ (.A1(_03940_),
    .A2(_04055_),
    .Y(_04522_),
    .B1(net5215));
 sg13g2_nand2_1 _21336_ (.Y(_04523_),
    .A(_04225_),
    .B(_04522_));
 sg13g2_o21ai_1 _21337_ (.B1(net5213),
    .Y(_04524_),
    .A1(_04092_),
    .A2(_04523_));
 sg13g2_o21ai_1 _21338_ (.B1(_04134_),
    .Y(_04525_),
    .A1(net5337),
    .A2(_04212_));
 sg13g2_nor2_1 _21339_ (.A(net5287),
    .B(_04074_),
    .Y(_04526_));
 sg13g2_a22oi_1 _21340_ (.Y(_04527_),
    .B1(_04526_),
    .B2(_04518_),
    .A2(_04525_),
    .A1(net5287));
 sg13g2_and3_1 _21341_ (.X(_04528_),
    .A(net5332),
    .B(_04086_),
    .C(_04201_));
 sg13g2_o21ai_1 _21342_ (.B1(net5288),
    .Y(_04529_),
    .A1(_04206_),
    .A2(_04528_));
 sg13g2_or2_1 _21343_ (.X(_04530_),
    .B(_04223_),
    .A(net5212));
 sg13g2_nand3_1 _21344_ (.B(_04529_),
    .C(_04530_),
    .A(_04216_),
    .Y(_04531_));
 sg13g2_a22oi_1 _21345_ (.Y(_04532_),
    .B1(_04531_),
    .B2(net5144),
    .A2(_04527_),
    .A1(net5143));
 sg13g2_o21ai_1 _21346_ (.B1(_04532_),
    .Y(_04533_),
    .A1(_04521_),
    .A2(_04524_));
 sg13g2_inv_1 _21347_ (.Y(_04534_),
    .A(_04533_));
 sg13g2_xor2_1 _21348_ (.B(_04533_),
    .A(_04509_),
    .X(_04535_));
 sg13g2_a21oi_1 _21349_ (.A1(_04484_),
    .A2(_04509_),
    .Y(_04536_),
    .B1(_04491_));
 sg13g2_nor2_1 _21350_ (.A(_04510_),
    .B(_04536_),
    .Y(_04537_));
 sg13g2_nor3_1 _21351_ (.A(_04510_),
    .B(_04535_),
    .C(_04536_),
    .Y(_04538_));
 sg13g2_xnor2_1 _21352_ (.Y(_04539_),
    .A(_04535_),
    .B(_04537_));
 sg13g2_nand2b_1 _21353_ (.Y(_04540_),
    .B(_04539_),
    .A_N(_04517_));
 sg13g2_xnor2_1 _21354_ (.Y(_04541_),
    .A(_04517_),
    .B(_04539_));
 sg13g2_a21oi_2 _21355_ (.B1(_04513_),
    .Y(_04542_),
    .A2(_04515_),
    .A1(_04514_));
 sg13g2_nand2b_1 _21356_ (.Y(_04543_),
    .B(_04541_),
    .A_N(_04542_));
 sg13g2_nand2b_1 _21357_ (.Y(_04544_),
    .B(_04542_),
    .A_N(_04541_));
 sg13g2_and3_1 _21358_ (.X(_01179_),
    .A(net5404),
    .B(_04543_),
    .C(_04544_));
 sg13g2_nand2_2 _21359_ (.Y(_04545_),
    .A(_04540_),
    .B(_04543_));
 sg13g2_nor3_1 _21360_ (.A(net5292),
    .B(_04070_),
    .C(_04218_),
    .Y(_04546_));
 sg13g2_nor3_1 _21361_ (.A(net5288),
    .B(_04065_),
    .C(_04199_),
    .Y(_04547_));
 sg13g2_nor3_1 _21362_ (.A(net5300),
    .B(_04546_),
    .C(_04547_),
    .Y(_04548_));
 sg13g2_nand2b_1 _21363_ (.Y(_04549_),
    .B(_04216_),
    .A_N(_04099_));
 sg13g2_o21ai_1 _21364_ (.B1(net5300),
    .Y(_04550_),
    .A1(_04245_),
    .A2(_04549_));
 sg13g2_nor2b_1 _21365_ (.A(_04548_),
    .B_N(_04550_),
    .Y(_04551_));
 sg13g2_a21oi_1 _21366_ (.A1(_03538_),
    .A2(net5326),
    .Y(_04552_),
    .B1(_04246_));
 sg13g2_or2_1 _21367_ (.X(_04553_),
    .B(_04552_),
    .A(_04055_));
 sg13g2_a21oi_1 _21368_ (.A1(_04185_),
    .A2(_04218_),
    .Y(_04554_),
    .B1(_04250_));
 sg13g2_o21ai_1 _21369_ (.B1(_04554_),
    .Y(_04555_),
    .A1(net5292),
    .A2(_04057_));
 sg13g2_a22oi_1 _21370_ (.Y(_04556_),
    .B1(_04555_),
    .B2(net5144),
    .A2(_04553_),
    .A1(net5143));
 sg13g2_o21ai_1 _21371_ (.B1(_04556_),
    .Y(_04557_),
    .A1(_04039_),
    .A2(_04551_));
 sg13g2_xor2_1 _21372_ (.B(_04557_),
    .A(_04533_),
    .X(_04558_));
 sg13g2_a21oi_2 _21373_ (.B1(_04538_),
    .Y(_04559_),
    .A2(_04534_),
    .A1(_04509_));
 sg13g2_xnor2_1 _21374_ (.Y(_04560_),
    .A(_04558_),
    .B(_04559_));
 sg13g2_nand2_1 _21375_ (.Y(_04561_),
    .A(_04545_),
    .B(_04560_));
 sg13g2_o21ai_1 _21376_ (.B1(net5404),
    .Y(_04562_),
    .A1(_04545_),
    .A2(_04560_));
 sg13g2_nor2b_1 _21377_ (.A(_04562_),
    .B_N(_04561_),
    .Y(_01180_));
 sg13g2_a21oi_2 _21378_ (.B1(_04557_),
    .Y(_04563_),
    .A2(_04559_),
    .A1(_04533_));
 sg13g2_o21ai_1 _21379_ (.B1(_04557_),
    .Y(_04564_),
    .A1(_04533_),
    .A2(_04559_));
 sg13g2_nand2b_1 _21380_ (.Y(_04565_),
    .B(_04564_),
    .A_N(_04563_));
 sg13g2_and2_1 _21381_ (.A(_04561_),
    .B(_04565_),
    .X(_04566_));
 sg13g2_nor2_1 _21382_ (.A(_04561_),
    .B(_04565_),
    .Y(_04567_));
 sg13g2_nor3_2 _21383_ (.A(net5407),
    .B(_04566_),
    .C(_04567_),
    .Y(_01181_));
 sg13g2_nor2_1 _21384_ (.A(_04563_),
    .B(_04567_),
    .Y(_04568_));
 sg13g2_nor2_2 _21385_ (.A(net5407),
    .B(_04568_),
    .Y(_01182_));
 sg13g2_nand3_1 _21386_ (.B(\r_pwm_even[2] ),
    .C(net5457),
    .A(net2901),
    .Y(_04569_));
 sg13g2_or2_1 _21387_ (.X(_04570_),
    .B(\r_pwm_even[2] ),
    .A(net2901));
 sg13g2_nand3_1 _21388_ (.B(_04569_),
    .C(_04570_),
    .A(net5457),
    .Y(_04571_));
 sg13g2_nand3_1 _21389_ (.B(\r_pwm_odd[1] ),
    .C(net5456),
    .A(net3733),
    .Y(_04572_));
 sg13g2_or2_1 _21390_ (.X(_04573_),
    .B(net3734),
    .A(_04571_));
 sg13g2_nand2_1 _21391_ (.Y(_04574_),
    .A(net5403),
    .B(_04573_));
 sg13g2_a21oi_1 _21392_ (.A1(_04571_),
    .A2(net3734),
    .Y(_01183_),
    .B1(_04574_));
 sg13g2_nand2_1 _21393_ (.Y(_04575_),
    .A(_04569_),
    .B(_04573_));
 sg13g2_nor2b_1 _21394_ (.A(net7338),
    .B_N(_04080_),
    .Y(_04576_));
 sg13g2_nand3_1 _21395_ (.B(net7338),
    .C(net5456),
    .A(net7295),
    .Y(_04577_));
 sg13g2_nand2b_1 _21396_ (.Y(_04578_),
    .B(_04577_),
    .A_N(_04576_));
 sg13g2_and2_1 _21397_ (.A(_04575_),
    .B(_04578_),
    .X(_04579_));
 sg13g2_o21ai_1 _21398_ (.B1(net5403),
    .Y(_04580_),
    .A1(_04575_),
    .A2(_04578_));
 sg13g2_nor2_1 _21399_ (.A(_04579_),
    .B(net7339),
    .Y(_01184_));
 sg13g2_nand2_1 _21400_ (.Y(_04581_),
    .A(\r_pwm_even[4] ),
    .B(net5457));
 sg13g2_nand2b_1 _21401_ (.Y(_04582_),
    .B(_04121_),
    .A_N(_04118_));
 sg13g2_xor2_1 _21402_ (.B(_04084_),
    .A(_04082_),
    .X(_04583_));
 sg13g2_nand2b_1 _21403_ (.Y(_04584_),
    .B(_04583_),
    .A_N(_04581_));
 sg13g2_xnor2_1 _21404_ (.Y(_04585_),
    .A(_04581_),
    .B(_04583_));
 sg13g2_nor2_1 _21405_ (.A(_04081_),
    .B(_04576_),
    .Y(_04586_));
 sg13g2_nand2_1 _21406_ (.Y(_04587_),
    .A(_04585_),
    .B(_04586_));
 sg13g2_xor2_1 _21407_ (.B(_04586_),
    .A(_04585_),
    .X(_04588_));
 sg13g2_nand2_1 _21408_ (.Y(_04589_),
    .A(_04579_),
    .B(_04588_));
 sg13g2_o21ai_1 _21409_ (.B1(net5403),
    .Y(_04590_),
    .A1(_04579_),
    .A2(_04588_));
 sg13g2_nor2b_1 _21410_ (.A(_04590_),
    .B_N(_04589_),
    .Y(_01185_));
 sg13g2_nand2_1 _21411_ (.Y(_04591_),
    .A(_04587_),
    .B(_04589_));
 sg13g2_nand2_1 _21412_ (.Y(_04592_),
    .A(\r_pwm_even[5] ),
    .B(net5456));
 sg13g2_nor2_1 _21413_ (.A(_04156_),
    .B(_04161_),
    .Y(_04593_));
 sg13g2_xnor2_1 _21414_ (.Y(_04594_),
    .A(_04122_),
    .B(_04159_));
 sg13g2_nor2_1 _21415_ (.A(_04592_),
    .B(_04594_),
    .Y(_04595_));
 sg13g2_xor2_1 _21416_ (.B(_04594_),
    .A(_04592_),
    .X(_04596_));
 sg13g2_nand2_1 _21417_ (.Y(_04597_),
    .A(_04582_),
    .B(_04584_));
 sg13g2_nand2_1 _21418_ (.Y(_04598_),
    .A(_04596_),
    .B(_04597_));
 sg13g2_xor2_1 _21419_ (.B(_04597_),
    .A(_04596_),
    .X(_04599_));
 sg13g2_or2_1 _21420_ (.X(_04600_),
    .B(_04599_),
    .A(_04591_));
 sg13g2_nand2_1 _21421_ (.Y(_04601_),
    .A(_04591_),
    .B(_04599_));
 sg13g2_and3_1 _21422_ (.X(_01186_),
    .A(net5405),
    .B(_04600_),
    .C(_04601_));
 sg13g2_nand2_1 _21423_ (.Y(_04602_),
    .A(_04598_),
    .B(_04601_));
 sg13g2_nand2_1 _21424_ (.Y(_04603_),
    .A(\r_pwm_even[6] ),
    .B(net5456));
 sg13g2_xnor2_1 _21425_ (.Y(_04604_),
    .A(_04162_),
    .B(_04195_));
 sg13g2_nor2_1 _21426_ (.A(_04603_),
    .B(_04604_),
    .Y(_04605_));
 sg13g2_xor2_1 _21427_ (.B(_04604_),
    .A(_04603_),
    .X(_04606_));
 sg13g2_nor2_1 _21428_ (.A(_04593_),
    .B(_04595_),
    .Y(_04607_));
 sg13g2_nor2b_1 _21429_ (.A(_04607_),
    .B_N(_04606_),
    .Y(_04608_));
 sg13g2_xnor2_1 _21430_ (.Y(_04609_),
    .A(_04606_),
    .B(_04607_));
 sg13g2_and2_1 _21431_ (.A(_04602_),
    .B(_04609_),
    .X(_04610_));
 sg13g2_o21ai_1 _21432_ (.B1(net5403),
    .Y(_04611_),
    .A1(_04602_),
    .A2(_04609_));
 sg13g2_nor2_1 _21433_ (.A(_04610_),
    .B(_04611_),
    .Y(_01187_));
 sg13g2_or2_1 _21434_ (.X(_04612_),
    .B(_04610_),
    .A(_04608_));
 sg13g2_nand2_1 _21435_ (.Y(_04613_),
    .A(\r_pwm_even[7] ),
    .B(net5456));
 sg13g2_nor2_1 _21436_ (.A(_04233_),
    .B(_04237_),
    .Y(_04614_));
 sg13g2_xnor2_1 _21437_ (.Y(_04615_),
    .A(_04198_),
    .B(_04235_));
 sg13g2_nor2_1 _21438_ (.A(_04613_),
    .B(_04615_),
    .Y(_04616_));
 sg13g2_xor2_1 _21439_ (.B(_04615_),
    .A(_04613_),
    .X(_04617_));
 sg13g2_a21oi_1 _21440_ (.A1(_04192_),
    .A2(_04197_),
    .Y(_04618_),
    .B1(_04605_));
 sg13g2_nor2b_1 _21441_ (.A(_04618_),
    .B_N(_04617_),
    .Y(_04619_));
 sg13g2_xnor2_1 _21442_ (.Y(_04620_),
    .A(_04617_),
    .B(_04618_));
 sg13g2_nor2_1 _21443_ (.A(_04612_),
    .B(_04620_),
    .Y(_04621_));
 sg13g2_a21oi_1 _21444_ (.A1(_04612_),
    .A2(_04620_),
    .Y(_04622_),
    .B1(net5407));
 sg13g2_nor2b_1 _21445_ (.A(_04621_),
    .B_N(_04622_),
    .Y(_01188_));
 sg13g2_a21o_1 _21446_ (.A2(_04620_),
    .A1(_04612_),
    .B1(_04619_),
    .X(_04623_));
 sg13g2_o21ai_1 _21447_ (.B1(_04238_),
    .Y(_04624_),
    .A1(_04614_),
    .A2(_04616_));
 sg13g2_or3_1 _21448_ (.A(_04238_),
    .B(_04614_),
    .C(_04616_),
    .X(_04625_));
 sg13g2_and2_1 _21449_ (.A(_04624_),
    .B(_04625_),
    .X(_04626_));
 sg13g2_nand2_1 _21450_ (.Y(_04627_),
    .A(_04623_),
    .B(_04626_));
 sg13g2_o21ai_1 _21451_ (.B1(net5403),
    .Y(_04628_),
    .A1(_04623_),
    .A2(_04626_));
 sg13g2_nor2b_1 _21452_ (.A(_04628_),
    .B_N(_04627_),
    .Y(_01189_));
 sg13g2_nor2b_1 _21453_ (.A(_04238_),
    .B_N(_04257_),
    .Y(_04629_));
 sg13g2_nand2_1 _21454_ (.Y(_04630_),
    .A(_04262_),
    .B(_04629_));
 sg13g2_xnor2_1 _21455_ (.Y(_04631_),
    .A(_04262_),
    .B(_04629_));
 sg13g2_and2_1 _21456_ (.A(_04624_),
    .B(_04627_),
    .X(_04632_));
 sg13g2_and2_1 _21457_ (.A(_04631_),
    .B(_04632_),
    .X(_04633_));
 sg13g2_nor2_1 _21458_ (.A(_04631_),
    .B(_04632_),
    .Y(_04634_));
 sg13g2_nor3_2 _21459_ (.A(net5407),
    .B(_04633_),
    .C(_04634_),
    .Y(_01190_));
 sg13g2_nand2_1 _21460_ (.Y(_04635_),
    .A(_04260_),
    .B(_04630_));
 sg13g2_nor2_1 _21461_ (.A(_04634_),
    .B(_04635_),
    .Y(_04636_));
 sg13g2_nor3_1 _21462_ (.A(_04260_),
    .B(_04631_),
    .C(_04632_),
    .Y(_04637_));
 sg13g2_nor3_2 _21463_ (.A(net5407),
    .B(_04636_),
    .C(_04637_),
    .Y(_01191_));
 sg13g2_nand3_1 _21464_ (.B(\g_pwm_even[2] ),
    .C(net5460),
    .A(net2910),
    .Y(_04638_));
 sg13g2_or2_1 _21465_ (.X(_04639_),
    .B(\g_pwm_even[2] ),
    .A(net2910));
 sg13g2_nand3_1 _21466_ (.B(_04638_),
    .C(_04639_),
    .A(net5460),
    .Y(_04640_));
 sg13g2_nand3_1 _21467_ (.B(\g_pwm_odd[1] ),
    .C(net5460),
    .A(net3761),
    .Y(_04641_));
 sg13g2_or2_1 _21468_ (.X(_04642_),
    .B(net3762),
    .A(_04640_));
 sg13g2_nand2_1 _21469_ (.Y(_04643_),
    .A(net5406),
    .B(_04642_));
 sg13g2_a21oi_1 _21470_ (.A1(_04640_),
    .A2(net3762),
    .Y(_01192_),
    .B1(_04643_));
 sg13g2_nand2_1 _21471_ (.Y(_04644_),
    .A(_04638_),
    .B(_04642_));
 sg13g2_or2_1 _21472_ (.X(_04645_),
    .B(_04288_),
    .A(\g_pwm_even[3] ));
 sg13g2_nand3_1 _21473_ (.B(\g_pwm_even[3] ),
    .C(net5460),
    .A(net7269),
    .Y(_04646_));
 sg13g2_nand2_1 _21474_ (.Y(_04647_),
    .A(_04645_),
    .B(net7270));
 sg13g2_and2_1 _21475_ (.A(_04644_),
    .B(_04647_),
    .X(_04648_));
 sg13g2_o21ai_1 _21476_ (.B1(net5406),
    .Y(_04649_),
    .A1(_04644_),
    .A2(_04647_));
 sg13g2_nor2_1 _21477_ (.A(_04648_),
    .B(net7271),
    .Y(_01193_));
 sg13g2_nand2_1 _21478_ (.Y(_04650_),
    .A(\g_pwm_even[4] ),
    .B(net5460));
 sg13g2_nand2_1 _21479_ (.Y(_04651_),
    .A(_04317_),
    .B(_04320_));
 sg13g2_xnor2_1 _21480_ (.Y(_04652_),
    .A(_04290_),
    .B(_04292_));
 sg13g2_nand2b_1 _21481_ (.Y(_04653_),
    .B(_04652_),
    .A_N(_04650_));
 sg13g2_xnor2_1 _21482_ (.Y(_04654_),
    .A(_04650_),
    .B(_04652_));
 sg13g2_and2_1 _21483_ (.A(_04289_),
    .B(_04645_),
    .X(_04655_));
 sg13g2_nand2_1 _21484_ (.Y(_04656_),
    .A(_04654_),
    .B(_04655_));
 sg13g2_xor2_1 _21485_ (.B(_04655_),
    .A(_04654_),
    .X(_04657_));
 sg13g2_nand2_1 _21486_ (.Y(_04658_),
    .A(_04648_),
    .B(_04657_));
 sg13g2_o21ai_1 _21487_ (.B1(net5406),
    .Y(_04659_),
    .A1(_04648_),
    .A2(_04657_));
 sg13g2_nor2b_1 _21488_ (.A(_04659_),
    .B_N(_04658_),
    .Y(_01194_));
 sg13g2_nand2_1 _21489_ (.Y(_04660_),
    .A(_04656_),
    .B(_04658_));
 sg13g2_nand2_1 _21490_ (.Y(_04661_),
    .A(\g_pwm_even[5] ),
    .B(net5459));
 sg13g2_nor2_1 _21491_ (.A(_04336_),
    .B(_04340_),
    .Y(_04662_));
 sg13g2_xor2_1 _21492_ (.B(_04338_),
    .A(_04321_),
    .X(_04663_));
 sg13g2_nor2_1 _21493_ (.A(_04661_),
    .B(_04663_),
    .Y(_04664_));
 sg13g2_xor2_1 _21494_ (.B(_04663_),
    .A(_04661_),
    .X(_04665_));
 sg13g2_nand2_1 _21495_ (.Y(_04666_),
    .A(_04651_),
    .B(_04653_));
 sg13g2_and2_1 _21496_ (.A(_04665_),
    .B(_04666_),
    .X(_04667_));
 sg13g2_xor2_1 _21497_ (.B(_04666_),
    .A(_04665_),
    .X(_04668_));
 sg13g2_a21oi_1 _21498_ (.A1(_04660_),
    .A2(_04668_),
    .Y(_04669_),
    .B1(net5409));
 sg13g2_o21ai_1 _21499_ (.B1(_04669_),
    .Y(_04670_),
    .A1(_04660_),
    .A2(_04668_));
 sg13g2_inv_1 _21500_ (.Y(_01195_),
    .A(_04670_));
 sg13g2_a21oi_1 _21501_ (.A1(_04660_),
    .A2(_04668_),
    .Y(_04671_),
    .B1(_04667_));
 sg13g2_nand2_1 _21502_ (.Y(_04672_),
    .A(\g_pwm_even[6] ),
    .B(net5461));
 sg13g2_nor2_1 _21503_ (.A(_04362_),
    .B(_04366_),
    .Y(_04673_));
 sg13g2_xor2_1 _21504_ (.B(_04365_),
    .A(_04341_),
    .X(_04674_));
 sg13g2_nor2_1 _21505_ (.A(_04672_),
    .B(_04674_),
    .Y(_04675_));
 sg13g2_xor2_1 _21506_ (.B(_04674_),
    .A(_04672_),
    .X(_04676_));
 sg13g2_nor2_1 _21507_ (.A(_04662_),
    .B(_04664_),
    .Y(_04677_));
 sg13g2_nor2b_1 _21508_ (.A(_04677_),
    .B_N(_04676_),
    .Y(_04678_));
 sg13g2_xor2_1 _21509_ (.B(_04677_),
    .A(_04676_),
    .X(_04679_));
 sg13g2_nor2_1 _21510_ (.A(_04671_),
    .B(_04679_),
    .Y(_04680_));
 sg13g2_a21oi_1 _21511_ (.A1(_04671_),
    .A2(_04679_),
    .Y(_04681_),
    .B1(net5410));
 sg13g2_nor2b_1 _21512_ (.A(_04680_),
    .B_N(_04681_),
    .Y(_01196_));
 sg13g2_nor2_1 _21513_ (.A(_04678_),
    .B(_04680_),
    .Y(_04682_));
 sg13g2_nand2_1 _21514_ (.Y(_04683_),
    .A(\g_pwm_even[7] ),
    .B(net5461));
 sg13g2_nor2_1 _21515_ (.A(_04383_),
    .B(_04388_),
    .Y(_04684_));
 sg13g2_xnor2_1 _21516_ (.Y(_04685_),
    .A(_04384_),
    .B(_04387_));
 sg13g2_nor2_1 _21517_ (.A(_04683_),
    .B(_04685_),
    .Y(_04686_));
 sg13g2_xor2_1 _21518_ (.B(_04685_),
    .A(_04683_),
    .X(_04687_));
 sg13g2_nor2_1 _21519_ (.A(_04673_),
    .B(_04675_),
    .Y(_04688_));
 sg13g2_nor2b_1 _21520_ (.A(_04688_),
    .B_N(_04687_),
    .Y(_04689_));
 sg13g2_xnor2_1 _21521_ (.Y(_04690_),
    .A(_04687_),
    .B(_04688_));
 sg13g2_nor2b_1 _21522_ (.A(_04690_),
    .B_N(_04682_),
    .Y(_04691_));
 sg13g2_nor2b_1 _21523_ (.A(_04682_),
    .B_N(_04690_),
    .Y(_04692_));
 sg13g2_nor3_1 _21524_ (.A(net5409),
    .B(_04691_),
    .C(_04692_),
    .Y(_01197_));
 sg13g2_or2_1 _21525_ (.X(_04693_),
    .B(_04692_),
    .A(_04689_));
 sg13g2_o21ai_1 _21526_ (.B1(_04389_),
    .Y(_04694_),
    .A1(_04684_),
    .A2(_04686_));
 sg13g2_or3_1 _21527_ (.A(_04389_),
    .B(_04684_),
    .C(_04686_),
    .X(_04695_));
 sg13g2_and2_1 _21528_ (.A(_04694_),
    .B(_04695_),
    .X(_04696_));
 sg13g2_nand2_1 _21529_ (.Y(_04697_),
    .A(_04693_),
    .B(_04696_));
 sg13g2_o21ai_1 _21530_ (.B1(net5406),
    .Y(_04698_),
    .A1(_04693_),
    .A2(_04696_));
 sg13g2_nor2b_1 _21531_ (.A(_04698_),
    .B_N(_04697_),
    .Y(_01198_));
 sg13g2_nand2_1 _21532_ (.Y(_04699_),
    .A(_04694_),
    .B(_04697_));
 sg13g2_nor2b_1 _21533_ (.A(_04389_),
    .B_N(_04398_),
    .Y(_04700_));
 sg13g2_nand2b_1 _21534_ (.Y(_04701_),
    .B(_04700_),
    .A_N(_04403_));
 sg13g2_xnor2_1 _21535_ (.Y(_04702_),
    .A(_04403_),
    .B(_04700_));
 sg13g2_or2_1 _21536_ (.X(_04703_),
    .B(_04702_),
    .A(_04699_));
 sg13g2_nand2_1 _21537_ (.Y(_04704_),
    .A(_04699_),
    .B(_04702_));
 sg13g2_and3_2 _21538_ (.X(_01199_),
    .A(net5404),
    .B(_04703_),
    .C(_04704_));
 sg13g2_nand3_1 _21539_ (.B(_04701_),
    .C(_04704_),
    .A(_04402_),
    .Y(_04705_));
 sg13g2_o21ai_1 _21540_ (.B1(net5404),
    .Y(_04706_),
    .A1(_04402_),
    .A2(_04704_));
 sg13g2_nor2b_2 _21541_ (.A(_04706_),
    .B_N(_04705_),
    .Y(_01200_));
 sg13g2_nor2b_2 _21542_ (.A(tia_vsync_last),
    .B_N(\atari2600.tia.vid_vsync ),
    .Y(_04707_));
 sg13g2_o21ai_1 _21543_ (.B1(net6025),
    .Y(_04708_),
    .A1(\frame_counter[0] ),
    .A2(_04707_));
 sg13g2_a21oi_1 _21544_ (.A1(_08042_),
    .A2(_04707_),
    .Y(_01201_),
    .B1(_04708_));
 sg13g2_o21ai_1 _21545_ (.B1(net6037),
    .Y(_04709_),
    .A1(\frame_counter[1] ),
    .A2(_04707_));
 sg13g2_a21oi_1 _21546_ (.A1(net3528),
    .A2(_04707_),
    .Y(_01202_),
    .B1(_04709_));
 sg13g2_o21ai_1 _21547_ (.B1(net6036),
    .Y(_04710_),
    .A1(net3528),
    .A2(_04707_));
 sg13g2_a21oi_1 _21548_ (.A1(_08041_),
    .A2(_04707_),
    .Y(_01203_),
    .B1(_04710_));
 sg13g2_nand2_2 _21549_ (.Y(_04711_),
    .A(_10480_),
    .B(_03113_));
 sg13g2_mux2_1 _21550_ (.A0(net5791),
    .A1(net4328),
    .S(_04711_),
    .X(_01204_));
 sg13g2_mux2_1 _21551_ (.A0(net5756),
    .A1(net6311),
    .S(_04711_),
    .X(_01205_));
 sg13g2_mux2_1 _21552_ (.A0(net5722),
    .A1(net4394),
    .S(_04711_),
    .X(_01206_));
 sg13g2_mux2_1 _21553_ (.A0(net5693),
    .A1(net6921),
    .S(_04711_),
    .X(_01207_));
 sg13g2_mux2_1 _21554_ (.A0(net5666),
    .A1(net6790),
    .S(_04711_),
    .X(_01208_));
 sg13g2_mux2_1 _21555_ (.A0(net5641),
    .A1(net6865),
    .S(_04711_),
    .X(_01209_));
 sg13g2_mux2_1 _21556_ (.A0(net5607),
    .A1(net7029),
    .S(_04711_),
    .X(_01210_));
 sg13g2_o21ai_1 _21557_ (.B1(net6000),
    .Y(_04712_),
    .A1(net5996),
    .A2(net7091));
 sg13g2_a21oi_1 _21558_ (.A1(net5996),
    .A2(net7),
    .Y(_01211_),
    .B1(_04712_));
 sg13g2_nand2b_1 _21559_ (.Y(_04713_),
    .B(net5996),
    .A_N(net5));
 sg13g2_nand2b_1 _21560_ (.Y(_04714_),
    .B(\atari2600.input_joystick_0[1] ),
    .A_N(net5996));
 sg13g2_nand3_1 _21561_ (.B(_04713_),
    .C(_04714_),
    .A(net6000),
    .Y(_01212_));
 sg13g2_a21oi_1 _21562_ (.A1(\joypmod[2] ),
    .A2(net5995),
    .Y(_04715_),
    .B1(net5978));
 sg13g2_o21ai_1 _21563_ (.B1(_04715_),
    .Y(_01213_),
    .A1(net5995),
    .A2(_08040_));
 sg13g2_nand2b_1 _21564_ (.Y(_04716_),
    .B(net5995),
    .A_N(net1));
 sg13g2_nand2b_1 _21565_ (.Y(_04717_),
    .B(net7020),
    .A_N(net5995));
 sg13g2_nand3_1 _21566_ (.B(_04716_),
    .C(_04717_),
    .A(net5999),
    .Y(_01214_));
 sg13g2_nand2b_1 _21567_ (.Y(_04718_),
    .B(net5996),
    .A_N(net2));
 sg13g2_nand2b_1 _21568_ (.Y(_04719_),
    .B(net7023),
    .A_N(net5996));
 sg13g2_nand3_1 _21569_ (.B(_04718_),
    .C(_04719_),
    .A(net6000),
    .Y(_01215_));
 sg13g2_nand2b_1 _21570_ (.Y(_04720_),
    .B(net5995),
    .A_N(net3));
 sg13g2_nand2b_1 _21571_ (.Y(_04721_),
    .B(net7102),
    .A_N(net5995));
 sg13g2_nand3_1 _21572_ (.B(_04720_),
    .C(_04721_),
    .A(net5999),
    .Y(_01216_));
 sg13g2_nand2b_1 _21573_ (.Y(_04722_),
    .B(net5995),
    .A_N(net4));
 sg13g2_nand2b_1 _21574_ (.Y(_04723_),
    .B(net6986),
    .A_N(net5995));
 sg13g2_nand3_1 _21575_ (.B(_04722_),
    .C(_04723_),
    .A(net5999),
    .Y(_01217_));
 sg13g2_a21oi_1 _21576_ (.A1(net5994),
    .A2(net6969),
    .Y(_04724_),
    .B1(net5978));
 sg13g2_o21ai_1 _21577_ (.B1(_04724_),
    .Y(_01218_),
    .A1(net5994),
    .A2(net1));
 sg13g2_a21oi_1 _21578_ (.A1(net5994),
    .A2(net6997),
    .Y(_04725_),
    .B1(net5976));
 sg13g2_o21ai_1 _21579_ (.B1(_04725_),
    .Y(_01219_),
    .A1(net5994),
    .A2(net2));
 sg13g2_a21oi_1 _21580_ (.A1(net5994),
    .A2(net7094),
    .Y(_04726_),
    .B1(net5976));
 sg13g2_o21ai_1 _21581_ (.B1(_04726_),
    .Y(_01220_),
    .A1(net5994),
    .A2(net3));
 sg13g2_a21oi_1 _21582_ (.A1(net5994),
    .A2(net7044),
    .Y(_04727_),
    .B1(net5976));
 sg13g2_o21ai_1 _21583_ (.B1(_04727_),
    .Y(_01221_),
    .A1(net5994),
    .A2(net4));
 sg13g2_a21oi_1 _21584_ (.A1(net6323),
    .A2(net6),
    .Y(_04728_),
    .B1(net5977));
 sg13g2_o21ai_1 _21585_ (.B1(_04728_),
    .Y(_01222_),
    .A1(net6),
    .A2(net5));
 sg13g2_o21ai_1 _21586_ (.B1(_04409_),
    .Y(_04729_),
    .A1(_08130_),
    .A2(_04408_));
 sg13g2_nand2_1 _21587_ (.Y(_04730_),
    .A(\b_pwm_even[2] ),
    .B(net5459));
 sg13g2_a21oi_1 _21588_ (.A1(\b_pwm_odd[2] ),
    .A2(net5459),
    .Y(_04731_),
    .B1(_04407_));
 sg13g2_nand2b_1 _21589_ (.Y(_04732_),
    .B(_04407_),
    .A_N(_04410_));
 sg13g2_nand2b_1 _21590_ (.Y(_04733_),
    .B(_04732_),
    .A_N(_04731_));
 sg13g2_xor2_1 _21591_ (.B(_04733_),
    .A(_04730_),
    .X(_04734_));
 sg13g2_or2_1 _21592_ (.X(_04735_),
    .B(_04734_),
    .A(_04729_));
 sg13g2_nand2_1 _21593_ (.Y(_04736_),
    .A(_04729_),
    .B(_04734_));
 sg13g2_and3_1 _21594_ (.X(_01223_),
    .A(net5406),
    .B(_04735_),
    .C(_04736_));
 sg13g2_and2_1 _21595_ (.A(\b_pwm_even[3] ),
    .B(net5461),
    .X(_04737_));
 sg13g2_nor2_1 _21596_ (.A(_04426_),
    .B(_04433_),
    .Y(_04738_));
 sg13g2_o21ai_1 _21597_ (.B1(_04428_),
    .Y(_04739_),
    .A1(_04426_),
    .A2(_04433_));
 sg13g2_xnor2_1 _21598_ (.Y(_04740_),
    .A(_04737_),
    .B(_04739_));
 sg13g2_o21ai_1 _21599_ (.B1(_04732_),
    .Y(_04741_),
    .A1(_04730_),
    .A2(_04731_));
 sg13g2_nand2_1 _21600_ (.Y(_04742_),
    .A(_04740_),
    .B(_04741_));
 sg13g2_xnor2_1 _21601_ (.Y(_04743_),
    .A(_04740_),
    .B(_04741_));
 sg13g2_nor2_1 _21602_ (.A(_04736_),
    .B(_04743_),
    .Y(_04744_));
 sg13g2_a21oi_1 _21603_ (.A1(_04736_),
    .A2(_04743_),
    .Y(_04745_),
    .B1(net5409));
 sg13g2_nor2b_1 _21604_ (.A(_04744_),
    .B_N(_04745_),
    .Y(_01224_));
 sg13g2_o21ai_1 _21605_ (.B1(_04742_),
    .Y(_04746_),
    .A1(_04736_),
    .A2(_04743_));
 sg13g2_nand2_1 _21606_ (.Y(_04747_),
    .A(\b_pwm_even[4] ),
    .B(net5461));
 sg13g2_nor2_1 _21607_ (.A(_04456_),
    .B(_04461_),
    .Y(_04748_));
 sg13g2_xor2_1 _21608_ (.B(_04460_),
    .A(_04434_),
    .X(_04749_));
 sg13g2_nor2_1 _21609_ (.A(_04747_),
    .B(_04749_),
    .Y(_04750_));
 sg13g2_xor2_1 _21610_ (.B(_04749_),
    .A(_04747_),
    .X(_04751_));
 sg13g2_a21o_1 _21611_ (.A2(_04737_),
    .A1(_04428_),
    .B1(_04738_),
    .X(_04752_));
 sg13g2_xor2_1 _21612_ (.B(_04752_),
    .A(_04751_),
    .X(_04753_));
 sg13g2_nor2_1 _21613_ (.A(_04746_),
    .B(_04753_),
    .Y(_04754_));
 sg13g2_and2_1 _21614_ (.A(_04746_),
    .B(_04753_),
    .X(_04755_));
 sg13g2_nor3_1 _21615_ (.A(net5409),
    .B(_04754_),
    .C(_04755_),
    .Y(_01225_));
 sg13g2_a21oi_2 _21616_ (.B1(_04755_),
    .Y(_04756_),
    .A2(_04752_),
    .A1(_04751_));
 sg13g2_nand2_1 _21617_ (.Y(_04757_),
    .A(\b_pwm_even[5] ),
    .B(net5458));
 sg13g2_nor2_1 _21618_ (.A(_04485_),
    .B(_04489_),
    .Y(_04758_));
 sg13g2_xnor2_1 _21619_ (.Y(_04759_),
    .A(_04462_),
    .B(_04487_));
 sg13g2_nor2_1 _21620_ (.A(_04757_),
    .B(_04759_),
    .Y(_04760_));
 sg13g2_xor2_1 _21621_ (.B(_04759_),
    .A(_04757_),
    .X(_04761_));
 sg13g2_nor2_1 _21622_ (.A(_04748_),
    .B(_04750_),
    .Y(_04762_));
 sg13g2_o21ai_1 _21623_ (.B1(_04761_),
    .Y(_04763_),
    .A1(_04748_),
    .A2(_04750_));
 sg13g2_xor2_1 _21624_ (.B(_04762_),
    .A(_04761_),
    .X(_04764_));
 sg13g2_o21ai_1 _21625_ (.B1(net5406),
    .Y(_04765_),
    .A1(_04756_),
    .A2(_04764_));
 sg13g2_a21oi_1 _21626_ (.A1(_04756_),
    .A2(_04764_),
    .Y(_01226_),
    .B1(_04765_));
 sg13g2_o21ai_1 _21627_ (.B1(_04763_),
    .Y(_04766_),
    .A1(_04756_),
    .A2(_04764_));
 sg13g2_nand2_1 _21628_ (.Y(_04767_),
    .A(\b_pwm_even[6] ),
    .B(net5458));
 sg13g2_nor2_1 _21629_ (.A(_04512_),
    .B(_04516_),
    .Y(_04768_));
 sg13g2_xor2_1 _21630_ (.B(_04515_),
    .A(_04490_),
    .X(_04769_));
 sg13g2_nor2_1 _21631_ (.A(_04767_),
    .B(_04769_),
    .Y(_04770_));
 sg13g2_xor2_1 _21632_ (.B(_04769_),
    .A(_04767_),
    .X(_04771_));
 sg13g2_nor2_1 _21633_ (.A(_04758_),
    .B(_04760_),
    .Y(_04772_));
 sg13g2_nand2b_1 _21634_ (.Y(_04773_),
    .B(_04771_),
    .A_N(_04772_));
 sg13g2_xnor2_1 _21635_ (.Y(_04774_),
    .A(_04771_),
    .B(_04772_));
 sg13g2_nand2_1 _21636_ (.Y(_04775_),
    .A(_04766_),
    .B(_04774_));
 sg13g2_o21ai_1 _21637_ (.B1(net5404),
    .Y(_04776_),
    .A1(_04766_),
    .A2(_04774_));
 sg13g2_nor2b_1 _21638_ (.A(_04776_),
    .B_N(_04775_),
    .Y(_01227_));
 sg13g2_nand2_1 _21639_ (.Y(_04777_),
    .A(\b_pwm_even[7] ),
    .B(net5458));
 sg13g2_nand3_1 _21640_ (.B(_04543_),
    .C(_04544_),
    .A(_04539_),
    .Y(_04778_));
 sg13g2_xor2_1 _21641_ (.B(_04542_),
    .A(_04517_),
    .X(_04779_));
 sg13g2_nand2b_1 _21642_ (.Y(_04780_),
    .B(_04779_),
    .A_N(_04777_));
 sg13g2_xnor2_1 _21643_ (.Y(_04781_),
    .A(_04777_),
    .B(_04779_));
 sg13g2_nor2_1 _21644_ (.A(_04768_),
    .B(_04770_),
    .Y(_04782_));
 sg13g2_nand2b_1 _21645_ (.Y(_04783_),
    .B(_04781_),
    .A_N(_04782_));
 sg13g2_xor2_1 _21646_ (.B(_04782_),
    .A(_04781_),
    .X(_04784_));
 sg13g2_nand3_1 _21647_ (.B(_04775_),
    .C(_04784_),
    .A(_04773_),
    .Y(_04785_));
 sg13g2_a21o_1 _21648_ (.A2(_04775_),
    .A1(_04773_),
    .B1(_04784_),
    .X(_04786_));
 sg13g2_and3_1 _21649_ (.X(_01228_),
    .A(net5404),
    .B(_04785_),
    .C(_04786_));
 sg13g2_nand2_1 _21650_ (.Y(_04787_),
    .A(_04783_),
    .B(_04786_));
 sg13g2_nand2_1 _21651_ (.Y(_04788_),
    .A(_04778_),
    .B(_04780_));
 sg13g2_xor2_1 _21652_ (.B(_04788_),
    .A(_04545_),
    .X(_04789_));
 sg13g2_and2_1 _21653_ (.A(_04787_),
    .B(_04789_),
    .X(_04790_));
 sg13g2_o21ai_1 _21654_ (.B1(net5404),
    .Y(_04791_),
    .A1(_04787_),
    .A2(_04789_));
 sg13g2_nor2_1 _21655_ (.A(_04790_),
    .B(_04791_),
    .Y(_01229_));
 sg13g2_nor2b_1 _21656_ (.A(_04545_),
    .B_N(_04560_),
    .Y(_04792_));
 sg13g2_xnor2_1 _21657_ (.Y(_04793_),
    .A(_04565_),
    .B(_04792_));
 sg13g2_a21oi_1 _21658_ (.A1(_04545_),
    .A2(_04788_),
    .Y(_04794_),
    .B1(_04790_));
 sg13g2_nor2b_1 _21659_ (.A(_04793_),
    .B_N(_04794_),
    .Y(_04795_));
 sg13g2_nor2b_1 _21660_ (.A(_04794_),
    .B_N(_04793_),
    .Y(_04796_));
 sg13g2_nor3_2 _21661_ (.A(net5408),
    .B(_04795_),
    .C(_04796_),
    .Y(_01230_));
 sg13g2_a21oi_1 _21662_ (.A1(_04564_),
    .A2(_04792_),
    .Y(_04797_),
    .B1(_04563_));
 sg13g2_mux2_1 _21663_ (.A0(_04797_),
    .A1(_04563_),
    .S(_04796_),
    .X(_04798_));
 sg13g2_nor2_2 _21664_ (.A(net5407),
    .B(_04798_),
    .Y(_01231_));
 sg13g2_nand2_2 _21665_ (.Y(_04799_),
    .A(net5424),
    .B(net5417));
 sg13g2_mux2_1 _21666_ (.A0(net5775),
    .A1(net4486),
    .S(_04799_),
    .X(_01232_));
 sg13g2_mux2_1 _21667_ (.A0(net5746),
    .A1(net6690),
    .S(_04799_),
    .X(_01233_));
 sg13g2_mux2_1 _21668_ (.A0(net5715),
    .A1(net6363),
    .S(_04799_),
    .X(_01234_));
 sg13g2_mux2_1 _21669_ (.A0(net5688),
    .A1(net6926),
    .S(_04799_),
    .X(_01235_));
 sg13g2_mux2_1 _21670_ (.A0(net5658),
    .A1(net6155),
    .S(_04799_),
    .X(_01236_));
 sg13g2_mux2_1 _21671_ (.A0(net5631),
    .A1(net6447),
    .S(_04799_),
    .X(_01237_));
 sg13g2_mux2_1 _21672_ (.A0(net5600),
    .A1(net6537),
    .S(_04799_),
    .X(_01238_));
 sg13g2_nor2_2 _21673_ (.A(net5473),
    .B(net5415),
    .Y(_04800_));
 sg13g2_mux2_1 _21674_ (.A0(net3688),
    .A1(net5794),
    .S(_04800_),
    .X(_01239_));
 sg13g2_mux2_1 _21675_ (.A0(net3573),
    .A1(net5766),
    .S(_04800_),
    .X(_01240_));
 sg13g2_mux2_1 _21676_ (.A0(net3294),
    .A1(net5737),
    .S(_04800_),
    .X(_01241_));
 sg13g2_mux2_1 _21677_ (.A0(net3630),
    .A1(net5708),
    .S(_04800_),
    .X(_01242_));
 sg13g2_mux2_1 _21678_ (.A0(net3448),
    .A1(net5680),
    .S(_04800_),
    .X(_01243_));
 sg13g2_mux2_1 _21679_ (.A0(net3332),
    .A1(net5651),
    .S(_04800_),
    .X(_01244_));
 sg13g2_mux2_1 _21680_ (.A0(net3539),
    .A1(net5622),
    .S(_04800_),
    .X(_01245_));
 sg13g2_nand2_2 _21681_ (.Y(_04801_),
    .A(_10497_),
    .B(_03104_));
 sg13g2_mux2_1 _21682_ (.A0(net5786),
    .A1(net6250),
    .S(_04801_),
    .X(_01246_));
 sg13g2_mux2_1 _21683_ (.A0(net5764),
    .A1(net6193),
    .S(_04801_),
    .X(_01247_));
 sg13g2_mux2_1 _21684_ (.A0(net5733),
    .A1(net6916),
    .S(_04801_),
    .X(_01248_));
 sg13g2_mux2_1 _21685_ (.A0(net5704),
    .A1(net6282),
    .S(_04801_),
    .X(_01249_));
 sg13g2_mux2_1 _21686_ (.A0(net5678),
    .A1(net4222),
    .S(_04801_),
    .X(_01250_));
 sg13g2_mux2_1 _21687_ (.A0(net5644),
    .A1(net6252),
    .S(_04801_),
    .X(_01251_));
 sg13g2_mux2_1 _21688_ (.A0(net5619),
    .A1(net6341),
    .S(_04801_),
    .X(_01252_));
 sg13g2_and2_1 _21689_ (.A(net4746),
    .B(_03087_),
    .X(_04802_));
 sg13g2_nor2_1 _21690_ (.A(net3092),
    .B(net4716),
    .Y(_04803_));
 sg13g2_a21oi_1 _21691_ (.A1(net5266),
    .A2(net4716),
    .Y(_01253_),
    .B1(_04803_));
 sg13g2_nor2_1 _21692_ (.A(net3623),
    .B(net4716),
    .Y(_04804_));
 sg13g2_a21oi_1 _21693_ (.A1(net5240),
    .A2(net4716),
    .Y(_01254_),
    .B1(_04804_));
 sg13g2_nor2_1 _21694_ (.A(net3738),
    .B(net4716),
    .Y(_04805_));
 sg13g2_a21oi_1 _21695_ (.A1(net5138),
    .A2(net4716),
    .Y(_01255_),
    .B1(_04805_));
 sg13g2_nor2_1 _21696_ (.A(net3868),
    .B(net4715),
    .Y(_04806_));
 sg13g2_a21oi_1 _21697_ (.A1(net5108),
    .A2(net4715),
    .Y(_01256_),
    .B1(_04806_));
 sg13g2_nor2_1 _21698_ (.A(net3706),
    .B(net4715),
    .Y(_04807_));
 sg13g2_a21oi_1 _21699_ (.A1(net5181),
    .A2(net4715),
    .Y(_01257_),
    .B1(_04807_));
 sg13g2_nor2_1 _21700_ (.A(net3879),
    .B(net4715),
    .Y(_04808_));
 sg13g2_a21oi_1 _21701_ (.A1(net5153),
    .A2(net4715),
    .Y(_01258_),
    .B1(_04808_));
 sg13g2_nor2_1 _21702_ (.A(net3091),
    .B(net4716),
    .Y(_04809_));
 sg13g2_a21oi_1 _21703_ (.A1(net5084),
    .A2(net4716),
    .Y(_01259_),
    .B1(_04809_));
 sg13g2_nor2_1 _21704_ (.A(net3730),
    .B(net4715),
    .Y(_04810_));
 sg13g2_a21oi_1 _21705_ (.A1(net5061),
    .A2(net4715),
    .Y(_01260_),
    .B1(_04810_));
 sg13g2_nor2_2 _21706_ (.A(net4776),
    .B(_03047_),
    .Y(_04811_));
 sg13g2_nand2_2 _21707_ (.Y(_04812_),
    .A(net4747),
    .B(_04811_));
 sg13g2_mux2_1 _21708_ (.A0(net5252),
    .A1(net4504),
    .S(_04812_),
    .X(_01261_));
 sg13g2_mux2_1 _21709_ (.A0(net5231),
    .A1(net4411),
    .S(_04812_),
    .X(_01262_));
 sg13g2_mux2_1 _21710_ (.A0(net5122),
    .A1(net4227),
    .S(_04812_),
    .X(_01263_));
 sg13g2_mux2_1 _21711_ (.A0(net5094),
    .A1(net6658),
    .S(_04812_),
    .X(_01264_));
 sg13g2_mux2_1 _21712_ (.A0(net5190),
    .A1(net6553),
    .S(_04812_),
    .X(_01265_));
 sg13g2_mux2_1 _21713_ (.A0(net5170),
    .A1(net6158),
    .S(_04812_),
    .X(_01266_));
 sg13g2_mux2_1 _21714_ (.A0(net5071),
    .A1(net6816),
    .S(_04812_),
    .X(_01267_));
 sg13g2_mux2_1 _21715_ (.A0(net5053),
    .A1(net6110),
    .S(_04812_),
    .X(_01268_));
 sg13g2_nor2_2 _21716_ (.A(net5036),
    .B(_03164_),
    .Y(_04813_));
 sg13g2_nand2_2 _21717_ (.Y(_04814_),
    .A(net5038),
    .B(_03163_));
 sg13g2_nand2_2 _21718_ (.Y(_04815_),
    .A(net4748),
    .B(_04813_));
 sg13g2_mux2_1 _21719_ (.A0(net5254),
    .A1(net6355),
    .S(_04815_),
    .X(_01269_));
 sg13g2_mux2_1 _21720_ (.A0(net5222),
    .A1(net4255),
    .S(_04815_),
    .X(_01270_));
 sg13g2_mux2_1 _21721_ (.A0(net5119),
    .A1(net4427),
    .S(_04815_),
    .X(_01271_));
 sg13g2_mux2_1 _21722_ (.A0(net5093),
    .A1(net6569),
    .S(_04815_),
    .X(_01272_));
 sg13g2_mux2_1 _21723_ (.A0(net5188),
    .A1(net4449),
    .S(_04815_),
    .X(_01273_));
 sg13g2_mux2_1 _21724_ (.A0(net5162),
    .A1(net6657),
    .S(_04815_),
    .X(_01274_));
 sg13g2_mux2_1 _21725_ (.A0(net5069),
    .A1(net6484),
    .S(_04815_),
    .X(_01275_));
 sg13g2_mux2_1 _21726_ (.A0(net5047),
    .A1(net4175),
    .S(_04815_),
    .X(_01276_));
 sg13g2_nor2_1 _21727_ (.A(_08677_),
    .B(_03008_),
    .Y(_04816_));
 sg13g2_nand2_2 _21728_ (.Y(_04817_),
    .A(_03003_),
    .B(net4734));
 sg13g2_mux2_1 _21729_ (.A0(net5251),
    .A1(net4384),
    .S(_04817_),
    .X(_01277_));
 sg13g2_mux2_1 _21730_ (.A0(net5224),
    .A1(net6085),
    .S(_04817_),
    .X(_01278_));
 sg13g2_mux2_1 _21731_ (.A0(net5123),
    .A1(net6649),
    .S(_04817_),
    .X(_01279_));
 sg13g2_mux2_1 _21732_ (.A0(net5094),
    .A1(net4099),
    .S(_04817_),
    .X(_01280_));
 sg13g2_mux2_1 _21733_ (.A0(net5190),
    .A1(net4040),
    .S(_04817_),
    .X(_01281_));
 sg13g2_mux2_1 _21734_ (.A0(net5163),
    .A1(net4264),
    .S(_04817_),
    .X(_01282_));
 sg13g2_mux2_1 _21735_ (.A0(net5071),
    .A1(net4202),
    .S(_04817_),
    .X(_01283_));
 sg13g2_mux2_1 _21736_ (.A0(net5045),
    .A1(net4259),
    .S(_04817_),
    .X(_01284_));
 sg13g2_nor2_2 _21737_ (.A(_08677_),
    .B(_03089_),
    .Y(_04818_));
 sg13g2_nor2_1 _21738_ (.A(net3786),
    .B(net4714),
    .Y(_04819_));
 sg13g2_a21oi_1 _21739_ (.A1(net5267),
    .A2(_04818_),
    .Y(_01285_),
    .B1(_04819_));
 sg13g2_nor2_1 _21740_ (.A(net3217),
    .B(net4714),
    .Y(_04820_));
 sg13g2_a21oi_1 _21741_ (.A1(net5241),
    .A2(net4714),
    .Y(_01286_),
    .B1(_04820_));
 sg13g2_nor2_1 _21742_ (.A(net3383),
    .B(net4713),
    .Y(_04821_));
 sg13g2_a21oi_1 _21743_ (.A1(net5138),
    .A2(net4713),
    .Y(_01287_),
    .B1(_04821_));
 sg13g2_nor2_1 _21744_ (.A(net3247),
    .B(net4714),
    .Y(_04822_));
 sg13g2_a21oi_1 _21745_ (.A1(net5109),
    .A2(net4714),
    .Y(_01288_),
    .B1(_04822_));
 sg13g2_nor2_1 _21746_ (.A(net3861),
    .B(net4713),
    .Y(_04823_));
 sg13g2_a21oi_1 _21747_ (.A1(net5182),
    .A2(net4713),
    .Y(_01289_),
    .B1(_04823_));
 sg13g2_nor2_1 _21748_ (.A(net3158),
    .B(net4714),
    .Y(_04824_));
 sg13g2_a21oi_1 _21749_ (.A1(net5153),
    .A2(net4714),
    .Y(_01290_),
    .B1(_04824_));
 sg13g2_nor2_1 _21750_ (.A(net3165),
    .B(net4713),
    .Y(_04825_));
 sg13g2_a21oi_1 _21751_ (.A1(net5085),
    .A2(net4713),
    .Y(_01291_),
    .B1(_04825_));
 sg13g2_nor2_1 _21752_ (.A(net2968),
    .B(net4713),
    .Y(_04826_));
 sg13g2_a21oi_1 _21753_ (.A1(net5062),
    .A2(net4713),
    .Y(_01292_),
    .B1(_04826_));
 sg13g2_nand2_2 _21754_ (.Y(_04827_),
    .A(_03003_),
    .B(net4736));
 sg13g2_mux2_1 _21755_ (.A0(net5253),
    .A1(net4541),
    .S(_04827_),
    .X(_01293_));
 sg13g2_mux2_1 _21756_ (.A0(net5225),
    .A1(net6737),
    .S(_04827_),
    .X(_01294_));
 sg13g2_mux2_1 _21757_ (.A0(net5123),
    .A1(net6153),
    .S(_04827_),
    .X(_01295_));
 sg13g2_mux2_1 _21758_ (.A0(net5101),
    .A1(net4155),
    .S(_04827_),
    .X(_01296_));
 sg13g2_mux2_1 _21759_ (.A0(net5195),
    .A1(net6072),
    .S(_04827_),
    .X(_01297_));
 sg13g2_mux2_1 _21760_ (.A0(net5171),
    .A1(net6523),
    .S(_04827_),
    .X(_01298_));
 sg13g2_mux2_1 _21761_ (.A0(net5075),
    .A1(net4437),
    .S(_04827_),
    .X(_01299_));
 sg13g2_mux2_1 _21762_ (.A0(net5054),
    .A1(net4055),
    .S(_04827_),
    .X(_01300_));
 sg13g2_nor2_2 _21763_ (.A(_08580_),
    .B(_03089_),
    .Y(_04828_));
 sg13g2_nor2_1 _21764_ (.A(net3048),
    .B(net4712),
    .Y(_04829_));
 sg13g2_a21oi_1 _21765_ (.A1(net5268),
    .A2(net4712),
    .Y(_01301_),
    .B1(_04829_));
 sg13g2_nor2_1 _21766_ (.A(net3912),
    .B(net4711),
    .Y(_04830_));
 sg13g2_a21oi_1 _21767_ (.A1(net5241),
    .A2(net4711),
    .Y(_01302_),
    .B1(_04830_));
 sg13g2_nor2_1 _21768_ (.A(net3588),
    .B(net4712),
    .Y(_04831_));
 sg13g2_a21oi_1 _21769_ (.A1(net5137),
    .A2(net4712),
    .Y(_01303_),
    .B1(_04831_));
 sg13g2_nor2_1 _21770_ (.A(net3080),
    .B(net4711),
    .Y(_04832_));
 sg13g2_a21oi_1 _21771_ (.A1(net5108),
    .A2(net4711),
    .Y(_01304_),
    .B1(_04832_));
 sg13g2_nor2_1 _21772_ (.A(net3060),
    .B(net4711),
    .Y(_04833_));
 sg13g2_a21oi_1 _21773_ (.A1(net5182),
    .A2(net4711),
    .Y(_01305_),
    .B1(_04833_));
 sg13g2_nor2_1 _21774_ (.A(net3103),
    .B(net4711),
    .Y(_04834_));
 sg13g2_a21oi_1 _21775_ (.A1(net5153),
    .A2(net4711),
    .Y(_01306_),
    .B1(_04834_));
 sg13g2_nor2_1 _21776_ (.A(net3035),
    .B(net4712),
    .Y(_04835_));
 sg13g2_a21oi_1 _21777_ (.A1(net5084),
    .A2(net4712),
    .Y(_01307_),
    .B1(_04835_));
 sg13g2_nor2_1 _21778_ (.A(net3139),
    .B(net4712),
    .Y(_04836_));
 sg13g2_a21oi_1 _21779_ (.A1(net5062),
    .A2(net4712),
    .Y(_01308_),
    .B1(_04836_));
 sg13g2_nor2_1 _21780_ (.A(_03004_),
    .B(net4744),
    .Y(_04837_));
 sg13g2_nor2_1 _21781_ (.A(net3878),
    .B(net4710),
    .Y(_04838_));
 sg13g2_a21oi_1 _21782_ (.A1(net5261),
    .A2(net4710),
    .Y(_01309_),
    .B1(_04838_));
 sg13g2_nor2_1 _21783_ (.A(net3729),
    .B(net4710),
    .Y(_04839_));
 sg13g2_a21oi_1 _21784_ (.A1(net5240),
    .A2(net4710),
    .Y(_01310_),
    .B1(_04839_));
 sg13g2_nor2_1 _21785_ (.A(net3336),
    .B(_04837_),
    .Y(_04840_));
 sg13g2_a21oi_1 _21786_ (.A1(net5137),
    .A2(net4709),
    .Y(_01311_),
    .B1(_04840_));
 sg13g2_nor2_1 _21787_ (.A(net3844),
    .B(net4710),
    .Y(_04841_));
 sg13g2_a21oi_1 _21788_ (.A1(net5109),
    .A2(net4709),
    .Y(_01312_),
    .B1(_04841_));
 sg13g2_nor2_1 _21789_ (.A(net3353),
    .B(net4709),
    .Y(_04842_));
 sg13g2_a21oi_1 _21790_ (.A1(net5181),
    .A2(net4709),
    .Y(_01313_),
    .B1(_04842_));
 sg13g2_nor2_1 _21791_ (.A(net3811),
    .B(net4710),
    .Y(_04843_));
 sg13g2_a21oi_1 _21792_ (.A1(net5152),
    .A2(net4710),
    .Y(_01314_),
    .B1(_04843_));
 sg13g2_nor2_1 _21793_ (.A(net3112),
    .B(net4709),
    .Y(_04844_));
 sg13g2_a21oi_1 _21794_ (.A1(net5083),
    .A2(net4709),
    .Y(_01315_),
    .B1(_04844_));
 sg13g2_nor2_1 _21795_ (.A(net3817),
    .B(net4709),
    .Y(_04845_));
 sg13g2_a21oi_1 _21796_ (.A1(net5060),
    .A2(net4709),
    .Y(_01316_),
    .B1(_04845_));
 sg13g2_nand2_2 _21797_ (.Y(_04846_),
    .A(_03003_),
    .B(net4740));
 sg13g2_mux2_1 _21798_ (.A0(net5252),
    .A1(net6651),
    .S(_04846_),
    .X(_01317_));
 sg13g2_mux2_1 _21799_ (.A0(net5224),
    .A1(net4403),
    .S(_04846_),
    .X(_01318_));
 sg13g2_mux2_1 _21800_ (.A0(net5122),
    .A1(net6745),
    .S(_04846_),
    .X(_01319_));
 sg13g2_mux2_1 _21801_ (.A0(net5094),
    .A1(net6836),
    .S(_04846_),
    .X(_01320_));
 sg13g2_mux2_1 _21802_ (.A0(net5195),
    .A1(net6167),
    .S(_04846_),
    .X(_01321_));
 sg13g2_mux2_1 _21803_ (.A0(net5170),
    .A1(net4217),
    .S(_04846_),
    .X(_01322_));
 sg13g2_mux2_1 _21804_ (.A0(net5075),
    .A1(net4265),
    .S(_04846_),
    .X(_01323_));
 sg13g2_mux2_1 _21805_ (.A0(net5053),
    .A1(net4201),
    .S(_04846_),
    .X(_01324_));
 sg13g2_nand2_2 _21806_ (.Y(_04847_),
    .A(_03003_),
    .B(net4746));
 sg13g2_mux2_1 _21807_ (.A0(net5252),
    .A1(net6141),
    .S(_04847_),
    .X(_01325_));
 sg13g2_mux2_1 _21808_ (.A0(net5224),
    .A1(net6125),
    .S(_04847_),
    .X(_01326_));
 sg13g2_mux2_1 _21809_ (.A0(net5123),
    .A1(net6835),
    .S(_04847_),
    .X(_01327_));
 sg13g2_mux2_1 _21810_ (.A0(net5101),
    .A1(net6333),
    .S(_04847_),
    .X(_01328_));
 sg13g2_mux2_1 _21811_ (.A0(net5195),
    .A1(net6060),
    .S(_04847_),
    .X(_01329_));
 sg13g2_mux2_1 _21812_ (.A0(net5170),
    .A1(net6769),
    .S(_04847_),
    .X(_01330_));
 sg13g2_mux2_1 _21813_ (.A0(net5075),
    .A1(net6526),
    .S(_04847_),
    .X(_01331_));
 sg13g2_mux2_1 _21814_ (.A0(net5053),
    .A1(net6771),
    .S(_04847_),
    .X(_01332_));
 sg13g2_nor2_2 _21815_ (.A(net4742),
    .B(_03088_),
    .Y(_04848_));
 sg13g2_nor2_1 _21816_ (.A(net3088),
    .B(net4708),
    .Y(_04849_));
 sg13g2_a21oi_1 _21817_ (.A1(net5268),
    .A2(net4708),
    .Y(_01333_),
    .B1(_04849_));
 sg13g2_nor2_1 _21818_ (.A(net3833),
    .B(net4707),
    .Y(_04850_));
 sg13g2_a21oi_1 _21819_ (.A1(net5241),
    .A2(net4707),
    .Y(_01334_),
    .B1(_04850_));
 sg13g2_nor2_1 _21820_ (.A(net3079),
    .B(net4708),
    .Y(_04851_));
 sg13g2_a21oi_1 _21821_ (.A1(net5137),
    .A2(net4708),
    .Y(_01335_),
    .B1(_04851_));
 sg13g2_nor2_1 _21822_ (.A(net3666),
    .B(net4707),
    .Y(_04852_));
 sg13g2_a21oi_1 _21823_ (.A1(net5108),
    .A2(net4707),
    .Y(_01336_),
    .B1(_04852_));
 sg13g2_nor2_1 _21824_ (.A(net3008),
    .B(net4707),
    .Y(_04853_));
 sg13g2_a21oi_1 _21825_ (.A1(net5182),
    .A2(net4707),
    .Y(_01337_),
    .B1(_04853_));
 sg13g2_nor2_1 _21826_ (.A(net3039),
    .B(net4707),
    .Y(_04854_));
 sg13g2_a21oi_1 _21827_ (.A1(net5152),
    .A2(net4707),
    .Y(_01338_),
    .B1(_04854_));
 sg13g2_nor2_1 _21828_ (.A(net2997),
    .B(net4708),
    .Y(_04855_));
 sg13g2_a21oi_1 _21829_ (.A1(net5084),
    .A2(net4708),
    .Y(_01339_),
    .B1(_04855_));
 sg13g2_nor2_1 _21830_ (.A(net3210),
    .B(net4708),
    .Y(_04856_));
 sg13g2_a21oi_1 _21831_ (.A1(net5062),
    .A2(net4708),
    .Y(_01340_),
    .B1(_04856_));
 sg13g2_nand2_2 _21832_ (.Y(_04857_),
    .A(_03165_),
    .B(net4733));
 sg13g2_mux2_1 _21833_ (.A0(net5244),
    .A1(net6044),
    .S(_04857_),
    .X(_01341_));
 sg13g2_mux2_1 _21834_ (.A0(net5219),
    .A1(net4234),
    .S(_04857_),
    .X(_01342_));
 sg13g2_mux2_1 _21835_ (.A0(net5116),
    .A1(net4031),
    .S(_04857_),
    .X(_01343_));
 sg13g2_mux2_1 _21836_ (.A0(net5090),
    .A1(net4335),
    .S(_04857_),
    .X(_01344_));
 sg13g2_mux2_1 _21837_ (.A0(net5187),
    .A1(net4324),
    .S(_04857_),
    .X(_01345_));
 sg13g2_mux2_1 _21838_ (.A0(net5157),
    .A1(net4440),
    .S(_04857_),
    .X(_01346_));
 sg13g2_mux2_1 _21839_ (.A0(net5065),
    .A1(net6409),
    .S(_04857_),
    .X(_01347_));
 sg13g2_mux2_1 _21840_ (.A0(net5042),
    .A1(net4321),
    .S(_04857_),
    .X(_01348_));
 sg13g2_o21ai_1 _21841_ (.B1(net6037),
    .Y(_04858_),
    .A1(net5925),
    .A2(_03223_));
 sg13g2_a21oi_1 _21842_ (.A1(net5925),
    .A2(net7180),
    .Y(_01349_),
    .B1(_04858_));
 sg13g2_a21oi_1 _21843_ (.A1(net5925),
    .A2(net7180),
    .Y(_04859_),
    .B1(net5866));
 sg13g2_nand2_1 _21844_ (.Y(_04860_),
    .A(net6037),
    .B(_03224_));
 sg13g2_nor2_1 _21845_ (.A(_04859_),
    .B(_04860_),
    .Y(_01350_));
 sg13g2_xor2_1 _21846_ (.B(_03224_),
    .A(net5850),
    .X(_04861_));
 sg13g2_nor2_1 _21847_ (.A(net5991),
    .B(_04861_),
    .Y(_01351_));
 sg13g2_nor2_1 _21848_ (.A(net3887),
    .B(_03224_),
    .Y(_04862_));
 sg13g2_xnor2_1 _21849_ (.Y(_04863_),
    .A(\hvsync_gen.hpos[5] ),
    .B(_04862_));
 sg13g2_nor2_1 _21850_ (.A(_03231_),
    .B(net3888),
    .Y(_01352_));
 sg13g2_nor2_1 _21851_ (.A(net5527),
    .B(_03224_),
    .Y(_04864_));
 sg13g2_o21ai_1 _21852_ (.B1(_03230_),
    .Y(_04865_),
    .A1(net5846),
    .A2(_04864_));
 sg13g2_a21oi_1 _21853_ (.A1(net5844),
    .A2(_04864_),
    .Y(_01353_),
    .B1(_04865_));
 sg13g2_nor3_1 _21854_ (.A(net3479),
    .B(net5528),
    .C(_03224_),
    .Y(_04866_));
 sg13g2_xnor2_1 _21855_ (.Y(_04867_),
    .A(net5843),
    .B(_04866_));
 sg13g2_nor2_1 _21856_ (.A(_03231_),
    .B(net3480),
    .Y(_01354_));
 sg13g2_nor2_1 _21857_ (.A(_08690_),
    .B(_03224_),
    .Y(_04868_));
 sg13g2_xnor2_1 _21858_ (.Y(_04869_),
    .A(net5840),
    .B(_04868_));
 sg13g2_nor2_1 _21859_ (.A(_03231_),
    .B(_04869_),
    .Y(_01355_));
 sg13g2_nor3_1 _21860_ (.A(net3822),
    .B(_08690_),
    .C(_03224_),
    .Y(_04870_));
 sg13g2_xnor2_1 _21861_ (.Y(_04871_),
    .A(net5839),
    .B(_04870_));
 sg13g2_nor2_1 _21862_ (.A(_03231_),
    .B(net3823),
    .Y(_01356_));
 sg13g2_nand2_2 _21863_ (.Y(_04872_),
    .A(net4739),
    .B(_03165_));
 sg13g2_mux2_1 _21864_ (.A0(net5244),
    .A1(net4396),
    .S(_04872_),
    .X(_01357_));
 sg13g2_mux2_1 _21865_ (.A0(net5219),
    .A1(net4171),
    .S(_04872_),
    .X(_01358_));
 sg13g2_mux2_1 _21866_ (.A0(net5116),
    .A1(net6065),
    .S(_04872_),
    .X(_01359_));
 sg13g2_mux2_1 _21867_ (.A0(net5090),
    .A1(net6948),
    .S(_04872_),
    .X(_01360_));
 sg13g2_mux2_1 _21868_ (.A0(net5187),
    .A1(net4127),
    .S(_04872_),
    .X(_01361_));
 sg13g2_mux2_1 _21869_ (.A0(net5157),
    .A1(net4195),
    .S(_04872_),
    .X(_01362_));
 sg13g2_mux2_1 _21870_ (.A0(net5065),
    .A1(net4017),
    .S(_04872_),
    .X(_01363_));
 sg13g2_mux2_1 _21871_ (.A0(net5042),
    .A1(net6253),
    .S(_04872_),
    .X(_01364_));
 sg13g2_nand4_1 _21872_ (.B(_08289_),
    .C(_08349_),
    .A(_08286_),
    .Y(_04873_),
    .D(_08357_));
 sg13g2_nand2_1 _21873_ (.Y(_04874_),
    .A(_08288_),
    .B(_08524_));
 sg13g2_a21oi_1 _21874_ (.A1(net5971),
    .A2(net5969),
    .Y(_04875_),
    .B1(net5974));
 sg13g2_nor2b_1 _21875_ (.A(_04875_),
    .B_N(\atari2600.cpu.state[2] ),
    .Y(_04876_));
 sg13g2_a21oi_1 _21876_ (.A1(\atari2600.cpu.state[1] ),
    .A2(net5970),
    .Y(_04877_),
    .B1(\atari2600.cpu.state[0] ));
 sg13g2_nor2_1 _21877_ (.A(\atari2600.cpu.state[1] ),
    .B(net5969),
    .Y(_04878_));
 sg13g2_nand2_1 _21878_ (.Y(_04879_),
    .A(net5973),
    .B(net5972));
 sg13g2_o21ai_1 _21879_ (.B1(_04877_),
    .Y(_04880_),
    .A1(_04878_),
    .A2(_04879_));
 sg13g2_o21ai_1 _21880_ (.B1(_08230_),
    .Y(_04881_),
    .A1(net5545),
    .A2(_08294_));
 sg13g2_nand4_1 _21881_ (.B(_08281_),
    .C(_08311_),
    .A(_08172_),
    .Y(_04882_),
    .D(_08414_));
 sg13g2_nand3_1 _21882_ (.B(net5477),
    .C(net5440),
    .A(_08251_),
    .Y(_04883_));
 sg13g2_nor2_2 _21883_ (.A(_08521_),
    .B(_04883_),
    .Y(_04884_));
 sg13g2_o21ai_1 _21884_ (.B1(_04884_),
    .Y(_04885_),
    .A1(_04876_),
    .A2(_04880_));
 sg13g2_or4_1 _21885_ (.A(_08276_),
    .B(_04873_),
    .C(_04882_),
    .D(_04885_),
    .X(_04886_));
 sg13g2_nor2_1 _21886_ (.A(net5479),
    .B(net5402),
    .Y(_04887_));
 sg13g2_nand4_1 _21887_ (.B(_08295_),
    .C(_08424_),
    .A(_08235_),
    .Y(_04888_),
    .D(_04887_));
 sg13g2_nor4_1 _21888_ (.A(_08520_),
    .B(net5388),
    .C(_04886_),
    .D(_04888_),
    .Y(_04889_));
 sg13g2_nand2_2 _21889_ (.Y(_04890_),
    .A(_08172_),
    .B(_08387_));
 sg13g2_nor4_2 _21890_ (.A(net5311),
    .B(_08466_),
    .C(_04889_),
    .Y(_04891_),
    .D(_04890_));
 sg13g2_mux2_1 _21891_ (.A0(net7078),
    .A1(_10396_),
    .S(net5211),
    .X(_01365_));
 sg13g2_mux2_1 _21892_ (.A0(net7107),
    .A1(_10401_),
    .S(net5211),
    .X(_01366_));
 sg13g2_mux2_1 _21893_ (.A0(net7100),
    .A1(_10389_),
    .S(net5211),
    .X(_01367_));
 sg13g2_mux2_1 _21894_ (.A0(net7085),
    .A1(_10411_),
    .S(net5211),
    .X(_01368_));
 sg13g2_nor2_1 _21895_ (.A(net7011),
    .B(_04891_),
    .Y(_04892_));
 sg13g2_a21oi_1 _21896_ (.A1(_08595_),
    .A2(net5210),
    .Y(_01369_),
    .B1(_04892_));
 sg13g2_nand2_2 _21897_ (.Y(_04893_),
    .A(_03007_),
    .B(_03048_));
 sg13g2_nor2_1 _21898_ (.A(_08677_),
    .B(_04893_),
    .Y(_04894_));
 sg13g2_nor2_1 _21899_ (.A(net3292),
    .B(net4705),
    .Y(_04895_));
 sg13g2_a21oi_1 _21900_ (.A1(net5266),
    .A2(net4705),
    .Y(_01370_),
    .B1(_04895_));
 sg13g2_nor2_1 _21901_ (.A(net3747),
    .B(net4705),
    .Y(_04896_));
 sg13g2_a21oi_1 _21902_ (.A1(net5240),
    .A2(net4705),
    .Y(_01371_),
    .B1(_04896_));
 sg13g2_nor2_1 _21903_ (.A(net3019),
    .B(net4705),
    .Y(_04897_));
 sg13g2_a21oi_1 _21904_ (.A1(net5137),
    .A2(net4705),
    .Y(_01372_),
    .B1(_04897_));
 sg13g2_nor2_1 _21905_ (.A(net3026),
    .B(_04894_),
    .Y(_04898_));
 sg13g2_a21oi_1 _21906_ (.A1(net5109),
    .A2(net4706),
    .Y(_01373_),
    .B1(_04898_));
 sg13g2_nor2_1 _21907_ (.A(net3098),
    .B(net4705),
    .Y(_04899_));
 sg13g2_a21oi_1 _21908_ (.A1(net5181),
    .A2(net4705),
    .Y(_01374_),
    .B1(_04899_));
 sg13g2_nor2_1 _21909_ (.A(net3489),
    .B(net4706),
    .Y(_04900_));
 sg13g2_a21oi_1 _21910_ (.A1(net5152),
    .A2(net4706),
    .Y(_01375_),
    .B1(_04900_));
 sg13g2_nor2_1 _21911_ (.A(net3018),
    .B(net4706),
    .Y(_04901_));
 sg13g2_a21oi_1 _21912_ (.A1(net5087),
    .A2(net4706),
    .Y(_01376_),
    .B1(_04901_));
 sg13g2_nor2_1 _21913_ (.A(net2982),
    .B(net4706),
    .Y(_04902_));
 sg13g2_a21oi_1 _21914_ (.A1(net5060),
    .A2(net4706),
    .Y(_01377_),
    .B1(_04902_));
 sg13g2_nand2_2 _21915_ (.Y(_04903_),
    .A(net4737),
    .B(_03165_));
 sg13g2_mux2_1 _21916_ (.A0(net5244),
    .A1(net6169),
    .S(_04903_),
    .X(_01378_));
 sg13g2_mux2_1 _21917_ (.A0(net5222),
    .A1(net6631),
    .S(_04903_),
    .X(_01379_));
 sg13g2_mux2_1 _21918_ (.A0(net5119),
    .A1(net6144),
    .S(_04903_),
    .X(_01380_));
 sg13g2_mux2_1 _21919_ (.A0(net5090),
    .A1(net6566),
    .S(_04903_),
    .X(_01381_));
 sg13g2_mux2_1 _21920_ (.A0(net5188),
    .A1(net6439),
    .S(_04903_),
    .X(_01382_));
 sg13g2_mux2_1 _21921_ (.A0(net5157),
    .A1(net6344),
    .S(_04903_),
    .X(_01383_));
 sg13g2_mux2_1 _21922_ (.A0(net5069),
    .A1(net6429),
    .S(_04903_),
    .X(_01384_));
 sg13g2_mux2_1 _21923_ (.A0(net5042),
    .A1(net4258),
    .S(_04903_),
    .X(_01385_));
 sg13g2_nor2_1 _21924_ (.A(_08580_),
    .B(_04893_),
    .Y(_04904_));
 sg13g2_nor2_1 _21925_ (.A(net3009),
    .B(net4703),
    .Y(_04905_));
 sg13g2_a21oi_1 _21926_ (.A1(net5266),
    .A2(net4703),
    .Y(_01386_),
    .B1(_04905_));
 sg13g2_nor2_1 _21927_ (.A(net3326),
    .B(net4703),
    .Y(_04906_));
 sg13g2_a21oi_1 _21928_ (.A1(net5240),
    .A2(net4703),
    .Y(_01387_),
    .B1(_04906_));
 sg13g2_nor2_1 _21929_ (.A(net3191),
    .B(_04904_),
    .Y(_04907_));
 sg13g2_a21oi_1 _21930_ (.A1(net5137),
    .A2(net4703),
    .Y(_01388_),
    .B1(_04907_));
 sg13g2_nor2_1 _21931_ (.A(net3012),
    .B(net4703),
    .Y(_04908_));
 sg13g2_a21oi_1 _21932_ (.A1(net5109),
    .A2(net4704),
    .Y(_01389_),
    .B1(_04908_));
 sg13g2_nor2_1 _21933_ (.A(net2984),
    .B(net4703),
    .Y(_04909_));
 sg13g2_a21oi_1 _21934_ (.A1(net5181),
    .A2(net4703),
    .Y(_01390_),
    .B1(_04909_));
 sg13g2_nor2_1 _21935_ (.A(net3058),
    .B(net4704),
    .Y(_04910_));
 sg13g2_a21oi_1 _21936_ (.A1(net5152),
    .A2(net4704),
    .Y(_01391_),
    .B1(_04910_));
 sg13g2_nor2_1 _21937_ (.A(net3042),
    .B(net4704),
    .Y(_04911_));
 sg13g2_a21oi_1 _21938_ (.A1(net5087),
    .A2(net4704),
    .Y(_01392_),
    .B1(_04911_));
 sg13g2_nor2_1 _21939_ (.A(net3171),
    .B(net4704),
    .Y(_04912_));
 sg13g2_a21oi_1 _21940_ (.A1(net5060),
    .A2(net4704),
    .Y(_01393_),
    .B1(_04912_));
 sg13g2_nor3_2 _21941_ (.A(net5032),
    .B(_08735_),
    .C(_04893_),
    .Y(_04913_));
 sg13g2_nor2_1 _21942_ (.A(net3162),
    .B(net4701),
    .Y(_04914_));
 sg13g2_a21oi_1 _21943_ (.A1(net5266),
    .A2(net4701),
    .Y(_01394_),
    .B1(_04914_));
 sg13g2_nor2_1 _21944_ (.A(net3004),
    .B(net4702),
    .Y(_04915_));
 sg13g2_a21oi_1 _21945_ (.A1(net5240),
    .A2(_04913_),
    .Y(_01395_),
    .B1(_04915_));
 sg13g2_nor2_1 _21946_ (.A(net3455),
    .B(net4701),
    .Y(_04916_));
 sg13g2_a21oi_1 _21947_ (.A1(net5137),
    .A2(net4701),
    .Y(_01396_),
    .B1(_04916_));
 sg13g2_nor2_1 _21948_ (.A(net3968),
    .B(net4701),
    .Y(_04917_));
 sg13g2_a21oi_1 _21949_ (.A1(net5108),
    .A2(net4701),
    .Y(_01397_),
    .B1(_04917_));
 sg13g2_nor2_1 _21950_ (.A(net3764),
    .B(net4701),
    .Y(_04918_));
 sg13g2_a21oi_1 _21951_ (.A1(net5181),
    .A2(net4701),
    .Y(_01398_),
    .B1(_04918_));
 sg13g2_nor2_1 _21952_ (.A(net3610),
    .B(net4702),
    .Y(_04919_));
 sg13g2_a21oi_1 _21953_ (.A1(net5152),
    .A2(net4702),
    .Y(_01399_),
    .B1(_04919_));
 sg13g2_nor2_1 _21954_ (.A(net3815),
    .B(net4702),
    .Y(_04920_));
 sg13g2_a21oi_1 _21955_ (.A1(net5083),
    .A2(net4702),
    .Y(_01400_),
    .B1(_04920_));
 sg13g2_nor2_1 _21956_ (.A(net3059),
    .B(net4702),
    .Y(_04921_));
 sg13g2_a21oi_1 _21957_ (.A1(net5060),
    .A2(net4702),
    .Y(_01401_),
    .B1(_04921_));
 sg13g2_and2_1 _21958_ (.A(net4747),
    .B(_03048_),
    .X(_04922_));
 sg13g2_nor2_1 _21959_ (.A(net4046),
    .B(net4700),
    .Y(_04923_));
 sg13g2_a21oi_1 _21960_ (.A1(net5266),
    .A2(net4700),
    .Y(_01402_),
    .B1(_04923_));
 sg13g2_nor2_1 _21961_ (.A(net3153),
    .B(net4700),
    .Y(_04924_));
 sg13g2_a21oi_1 _21962_ (.A1(net5240),
    .A2(net4700),
    .Y(_01403_),
    .B1(_04924_));
 sg13g2_nor2_1 _21963_ (.A(net3113),
    .B(net4700),
    .Y(_04925_));
 sg13g2_a21oi_1 _21964_ (.A1(net5137),
    .A2(net4700),
    .Y(_01404_),
    .B1(_04925_));
 sg13g2_nor2_1 _21965_ (.A(net3109),
    .B(net4700),
    .Y(_04926_));
 sg13g2_a21oi_1 _21966_ (.A1(net5109),
    .A2(net4700),
    .Y(_01405_),
    .B1(_04926_));
 sg13g2_nor2_1 _21967_ (.A(net3104),
    .B(net4699),
    .Y(_04927_));
 sg13g2_a21oi_1 _21968_ (.A1(net5181),
    .A2(net4699),
    .Y(_01406_),
    .B1(_04927_));
 sg13g2_nor2_1 _21969_ (.A(net3967),
    .B(net4699),
    .Y(_04928_));
 sg13g2_a21oi_1 _21970_ (.A1(net5152),
    .A2(net4699),
    .Y(_01407_),
    .B1(_04928_));
 sg13g2_nor2_1 _21971_ (.A(net3650),
    .B(net4699),
    .Y(_04929_));
 sg13g2_a21oi_1 _21972_ (.A1(net5083),
    .A2(net4699),
    .Y(_01408_),
    .B1(_04929_));
 sg13g2_nor2_1 _21973_ (.A(net3085),
    .B(net4699),
    .Y(_04930_));
 sg13g2_a21oi_1 _21974_ (.A1(net5060),
    .A2(net4699),
    .Y(_01409_),
    .B1(_04930_));
 sg13g2_nor3_2 _21975_ (.A(net4878),
    .B(net5024),
    .C(_10253_),
    .Y(_04931_));
 sg13g2_nand2_2 _21976_ (.Y(_04932_),
    .A(net4739),
    .B(_04931_));
 sg13g2_mux2_1 _21977_ (.A0(net5255),
    .A1(net6478),
    .S(_04932_),
    .X(_01410_));
 sg13g2_mux2_1 _21978_ (.A0(net5228),
    .A1(net4273),
    .S(_04932_),
    .X(_01411_));
 sg13g2_mux2_1 _21979_ (.A0(net5126),
    .A1(net6145),
    .S(_04932_),
    .X(_01412_));
 sg13g2_mux2_1 _21980_ (.A0(net5098),
    .A1(net4479),
    .S(_04932_),
    .X(_01413_));
 sg13g2_mux2_1 _21981_ (.A0(net5193),
    .A1(net4087),
    .S(_04932_),
    .X(_01414_));
 sg13g2_mux2_1 _21982_ (.A0(net5165),
    .A1(net6281),
    .S(_04932_),
    .X(_01415_));
 sg13g2_mux2_1 _21983_ (.A0(net5072),
    .A1(net6275),
    .S(_04932_),
    .X(_01416_));
 sg13g2_mux2_1 _21984_ (.A0(net5051),
    .A1(net4117),
    .S(_04932_),
    .X(_01417_));
 sg13g2_nand2_2 _21985_ (.Y(_04933_),
    .A(net4736),
    .B(_04931_));
 sg13g2_mux2_1 _21986_ (.A0(net5255),
    .A1(net6703),
    .S(_04933_),
    .X(_01418_));
 sg13g2_mux2_1 _21987_ (.A0(net5228),
    .A1(net6563),
    .S(_04933_),
    .X(_01419_));
 sg13g2_mux2_1 _21988_ (.A0(net5126),
    .A1(net6094),
    .S(_04933_),
    .X(_01420_));
 sg13g2_mux2_1 _21989_ (.A0(net5098),
    .A1(net4205),
    .S(_04933_),
    .X(_01421_));
 sg13g2_mux2_1 _21990_ (.A0(net5193),
    .A1(net6778),
    .S(_04933_),
    .X(_01422_));
 sg13g2_mux2_1 _21991_ (.A0(net5165),
    .A1(net4376),
    .S(_04933_),
    .X(_01423_));
 sg13g2_mux2_1 _21992_ (.A0(net5072),
    .A1(net4475),
    .S(_04933_),
    .X(_01424_));
 sg13g2_mux2_1 _21993_ (.A0(net5050),
    .A1(net4041),
    .S(_04933_),
    .X(_01425_));
 sg13g2_nor2b_1 _21994_ (.A(net4744),
    .B_N(_04931_),
    .Y(_04934_));
 sg13g2_nor2_1 _21995_ (.A(net3128),
    .B(net4698),
    .Y(_04935_));
 sg13g2_a21oi_1 _21996_ (.A1(net5264),
    .A2(net4698),
    .Y(_01426_),
    .B1(_04935_));
 sg13g2_nor2_1 _21997_ (.A(net3049),
    .B(net4698),
    .Y(_04936_));
 sg13g2_a21oi_1 _21998_ (.A1(net5239),
    .A2(net4698),
    .Y(_01427_),
    .B1(_04936_));
 sg13g2_nor2_1 _21999_ (.A(net3036),
    .B(net4697),
    .Y(_04937_));
 sg13g2_a21oi_1 _22000_ (.A1(net5135),
    .A2(net4697),
    .Y(_01428_),
    .B1(_04937_));
 sg13g2_nor2_1 _22001_ (.A(net3976),
    .B(net4697),
    .Y(_04938_));
 sg13g2_a21oi_1 _22002_ (.A1(net5112),
    .A2(net4697),
    .Y(_01429_),
    .B1(_04938_));
 sg13g2_nor2_1 _22003_ (.A(net6408),
    .B(_04934_),
    .Y(_04939_));
 sg13g2_a21oi_1 _22004_ (.A1(net5180),
    .A2(net4698),
    .Y(_01430_),
    .B1(_04939_));
 sg13g2_nor2_1 _22005_ (.A(net4141),
    .B(net4698),
    .Y(_04940_));
 sg13g2_a21oi_1 _22006_ (.A1(net5150),
    .A2(net4698),
    .Y(_01431_),
    .B1(_04940_));
 sg13g2_nor2_1 _22007_ (.A(net3876),
    .B(net4697),
    .Y(_04941_));
 sg13g2_a21oi_1 _22008_ (.A1(net5086),
    .A2(net4697),
    .Y(_01432_),
    .B1(_04941_));
 sg13g2_nor2_1 _22009_ (.A(net3377),
    .B(net4697),
    .Y(_04942_));
 sg13g2_a21oi_1 _22010_ (.A1(net5059),
    .A2(net4697),
    .Y(_01433_),
    .B1(_04942_));
 sg13g2_nand2_2 _22011_ (.Y(_04943_),
    .A(net4740),
    .B(_04813_));
 sg13g2_mux2_1 _22012_ (.A0(net5254),
    .A1(net4370),
    .S(_04943_),
    .X(_01434_));
 sg13g2_mux2_1 _22013_ (.A0(net5222),
    .A1(net4183),
    .S(_04943_),
    .X(_01435_));
 sg13g2_mux2_1 _22014_ (.A0(net5118),
    .A1(net4091),
    .S(_04943_),
    .X(_01436_));
 sg13g2_mux2_1 _22015_ (.A0(net5093),
    .A1(net4144),
    .S(_04943_),
    .X(_01437_));
 sg13g2_mux2_1 _22016_ (.A0(net5188),
    .A1(net6269),
    .S(_04943_),
    .X(_01438_));
 sg13g2_mux2_1 _22017_ (.A0(net5162),
    .A1(net4039),
    .S(_04943_),
    .X(_01439_));
 sg13g2_mux2_1 _22018_ (.A0(net5070),
    .A1(net4170),
    .S(_04943_),
    .X(_01440_));
 sg13g2_mux2_1 _22019_ (.A0(net5047),
    .A1(net6464),
    .S(_04943_),
    .X(_01441_));
 sg13g2_nand2_2 _22020_ (.Y(_04944_),
    .A(net4734),
    .B(_04931_));
 sg13g2_mux2_1 _22021_ (.A0(net5255),
    .A1(net6714),
    .S(_04944_),
    .X(_01442_));
 sg13g2_mux2_1 _22022_ (.A0(net5228),
    .A1(net6575),
    .S(_04944_),
    .X(_01443_));
 sg13g2_mux2_1 _22023_ (.A0(net5126),
    .A1(net6089),
    .S(_04944_),
    .X(_01444_));
 sg13g2_mux2_1 _22024_ (.A0(net5099),
    .A1(net4111),
    .S(_04944_),
    .X(_01445_));
 sg13g2_mux2_1 _22025_ (.A0(net5194),
    .A1(net4103),
    .S(_04944_),
    .X(_01446_));
 sg13g2_mux2_1 _22026_ (.A0(net5167),
    .A1(net4513),
    .S(_04944_),
    .X(_01447_));
 sg13g2_mux2_1 _22027_ (.A0(net5073),
    .A1(net4062),
    .S(_04944_),
    .X(_01448_));
 sg13g2_mux2_1 _22028_ (.A0(net5050),
    .A1(net6638),
    .S(_04944_),
    .X(_01449_));
 sg13g2_nand2_2 _22029_ (.Y(_04945_),
    .A(net4738),
    .B(_04931_));
 sg13g2_mux2_1 _22030_ (.A0(net5255),
    .A1(net4006),
    .S(_04945_),
    .X(_01450_));
 sg13g2_mux2_1 _22031_ (.A0(net5228),
    .A1(net4393),
    .S(_04945_),
    .X(_01451_));
 sg13g2_mux2_1 _22032_ (.A0(net5126),
    .A1(net4422),
    .S(_04945_),
    .X(_01452_));
 sg13g2_mux2_1 _22033_ (.A0(net5099),
    .A1(net4340),
    .S(_04945_),
    .X(_01453_));
 sg13g2_mux2_1 _22034_ (.A0(net5194),
    .A1(net6114),
    .S(_04945_),
    .X(_01454_));
 sg13g2_mux2_1 _22035_ (.A0(net5167),
    .A1(net4225),
    .S(_04945_),
    .X(_01455_));
 sg13g2_mux2_1 _22036_ (.A0(net5073),
    .A1(net4327),
    .S(_04945_),
    .X(_01456_));
 sg13g2_mux2_1 _22037_ (.A0(net5050),
    .A1(net4477),
    .S(_04945_),
    .X(_01457_));
 sg13g2_nor2b_1 _22038_ (.A(net4742),
    .B_N(_04931_),
    .Y(_04946_));
 sg13g2_nor2_1 _22039_ (.A(net3017),
    .B(net4696),
    .Y(_04947_));
 sg13g2_a21oi_1 _22040_ (.A1(net5264),
    .A2(net4696),
    .Y(_01458_),
    .B1(_04947_));
 sg13g2_nor2_1 _22041_ (.A(net3114),
    .B(net4696),
    .Y(_04948_));
 sg13g2_a21oi_1 _22042_ (.A1(net5239),
    .A2(net4696),
    .Y(_01459_),
    .B1(_04948_));
 sg13g2_nor2_1 _22043_ (.A(net3344),
    .B(net4695),
    .Y(_04949_));
 sg13g2_a21oi_1 _22044_ (.A1(net5135),
    .A2(net4695),
    .Y(_01460_),
    .B1(_04949_));
 sg13g2_nor2_1 _22045_ (.A(net3951),
    .B(net4695),
    .Y(_04950_));
 sg13g2_a21oi_1 _22046_ (.A1(net5107),
    .A2(net4695),
    .Y(_01461_),
    .B1(_04950_));
 sg13g2_nor2_1 _22047_ (.A(net4331),
    .B(_04946_),
    .Y(_04951_));
 sg13g2_a21oi_1 _22048_ (.A1(net5180),
    .A2(net4695),
    .Y(_01462_),
    .B1(_04951_));
 sg13g2_nor2_1 _22049_ (.A(net3635),
    .B(net4696),
    .Y(_04952_));
 sg13g2_a21oi_1 _22050_ (.A1(net5150),
    .A2(net4696),
    .Y(_01463_),
    .B1(_04952_));
 sg13g2_nor2_1 _22051_ (.A(net4333),
    .B(net4696),
    .Y(_04953_));
 sg13g2_a21oi_1 _22052_ (.A1(net5083),
    .A2(net4695),
    .Y(_01464_),
    .B1(_04953_));
 sg13g2_nor2_1 _22053_ (.A(net6593),
    .B(net4695),
    .Y(_04954_));
 sg13g2_a21oi_1 _22054_ (.A1(net5059),
    .A2(net4695),
    .Y(_01465_),
    .B1(_04954_));
 sg13g2_nand2_2 _22055_ (.Y(_04955_),
    .A(net4747),
    .B(_04931_));
 sg13g2_mux2_1 _22056_ (.A0(net5255),
    .A1(net4480),
    .S(_04955_),
    .X(_01466_));
 sg13g2_mux2_1 _22057_ (.A0(net5228),
    .A1(net4472),
    .S(_04955_),
    .X(_01467_));
 sg13g2_mux2_1 _22058_ (.A0(net5126),
    .A1(net6922),
    .S(_04955_),
    .X(_01468_));
 sg13g2_mux2_1 _22059_ (.A0(net5099),
    .A1(net4364),
    .S(_04955_),
    .X(_01469_));
 sg13g2_mux2_1 _22060_ (.A0(net5192),
    .A1(net6903),
    .S(_04955_),
    .X(_01470_));
 sg13g2_mux2_1 _22061_ (.A0(net5166),
    .A1(net4160),
    .S(_04955_),
    .X(_01471_));
 sg13g2_mux2_1 _22062_ (.A0(net5073),
    .A1(net6127),
    .S(_04955_),
    .X(_01472_));
 sg13g2_mux2_1 _22063_ (.A0(net5050),
    .A1(net6424),
    .S(_04955_),
    .X(_01473_));
 sg13g2_nor2_2 _22064_ (.A(net4771),
    .B(_03047_),
    .Y(_04956_));
 sg13g2_nand2_2 _22065_ (.Y(_04957_),
    .A(net4739),
    .B(_04956_));
 sg13g2_mux2_1 _22066_ (.A0(net5255),
    .A1(net4294),
    .S(_04957_),
    .X(_01474_));
 sg13g2_mux2_1 _22067_ (.A0(net5229),
    .A1(net4296),
    .S(_04957_),
    .X(_01475_));
 sg13g2_mux2_1 _22068_ (.A0(net5127),
    .A1(net4092),
    .S(_04957_),
    .X(_01476_));
 sg13g2_mux2_1 _22069_ (.A0(net5098),
    .A1(net6135),
    .S(_04957_),
    .X(_01477_));
 sg13g2_mux2_1 _22070_ (.A0(net5193),
    .A1(net4300),
    .S(_04957_),
    .X(_01478_));
 sg13g2_mux2_1 _22071_ (.A0(net5168),
    .A1(net6335),
    .S(_04957_),
    .X(_01479_));
 sg13g2_mux2_1 _22072_ (.A0(net5072),
    .A1(net4110),
    .S(_04957_),
    .X(_01480_));
 sg13g2_mux2_1 _22073_ (.A0(net5050),
    .A1(net4531),
    .S(_04957_),
    .X(_01481_));
 sg13g2_nand2_2 _22074_ (.Y(_04958_),
    .A(net4736),
    .B(_04956_));
 sg13g2_mux2_1 _22075_ (.A0(net5256),
    .A1(net6556),
    .S(_04958_),
    .X(_01482_));
 sg13g2_mux2_1 _22076_ (.A0(net5229),
    .A1(net4497),
    .S(_04958_),
    .X(_01483_));
 sg13g2_mux2_1 _22077_ (.A0(net5127),
    .A1(net6220),
    .S(_04958_),
    .X(_01484_));
 sg13g2_mux2_1 _22078_ (.A0(net5098),
    .A1(net4138),
    .S(_04958_),
    .X(_01485_));
 sg13g2_mux2_1 _22079_ (.A0(net5194),
    .A1(net6346),
    .S(_04958_),
    .X(_01486_));
 sg13g2_mux2_1 _22080_ (.A0(net5165),
    .A1(net4456),
    .S(_04958_),
    .X(_01487_));
 sg13g2_mux2_1 _22081_ (.A0(net5072),
    .A1(net6827),
    .S(_04958_),
    .X(_01488_));
 sg13g2_mux2_1 _22082_ (.A0(net5050),
    .A1(net4063),
    .S(_04958_),
    .X(_01489_));
 sg13g2_nor2b_1 _22083_ (.A(net4744),
    .B_N(_04956_),
    .Y(_04959_));
 sg13g2_nor2_1 _22084_ (.A(net3050),
    .B(net4693),
    .Y(_04960_));
 sg13g2_a21oi_1 _22085_ (.A1(net5264),
    .A2(net4693),
    .Y(_01490_),
    .B1(_04960_));
 sg13g2_nor2_1 _22086_ (.A(net3998),
    .B(net4693),
    .Y(_04961_));
 sg13g2_a21oi_1 _22087_ (.A1(net5238),
    .A2(net4693),
    .Y(_01491_),
    .B1(_04961_));
 sg13g2_nor2_1 _22088_ (.A(net3439),
    .B(net4693),
    .Y(_04962_));
 sg13g2_a21oi_1 _22089_ (.A1(net5136),
    .A2(net4693),
    .Y(_01492_),
    .B1(_04962_));
 sg13g2_nor2_1 _22090_ (.A(net3016),
    .B(net4694),
    .Y(_04963_));
 sg13g2_a21oi_1 _22091_ (.A1(net5112),
    .A2(net4694),
    .Y(_01493_),
    .B1(_04963_));
 sg13g2_nor2_1 _22092_ (.A(net3889),
    .B(net4694),
    .Y(_04964_));
 sg13g2_a21oi_1 _22093_ (.A1(net5180),
    .A2(net4694),
    .Y(_01494_),
    .B1(_04964_));
 sg13g2_nor2_1 _22094_ (.A(net3185),
    .B(net4693),
    .Y(_04965_));
 sg13g2_a21oi_1 _22095_ (.A1(net5150),
    .A2(net4693),
    .Y(_01495_),
    .B1(_04965_));
 sg13g2_nor2_1 _22096_ (.A(net3084),
    .B(net4694),
    .Y(_04966_));
 sg13g2_a21oi_1 _22097_ (.A1(net5086),
    .A2(net4694),
    .Y(_01496_),
    .B1(_04966_));
 sg13g2_nor2_1 _22098_ (.A(net3698),
    .B(net4694),
    .Y(_04967_));
 sg13g2_a21oi_1 _22099_ (.A1(net5063),
    .A2(net4694),
    .Y(_01497_),
    .B1(_04967_));
 sg13g2_nand2_2 _22100_ (.Y(_04968_),
    .A(net4745),
    .B(_04956_));
 sg13g2_mux2_1 _22101_ (.A0(net5255),
    .A1(net6512),
    .S(_04968_),
    .X(_01498_));
 sg13g2_mux2_1 _22102_ (.A0(net5229),
    .A1(net6495),
    .S(_04968_),
    .X(_01499_));
 sg13g2_mux2_1 _22103_ (.A0(net5127),
    .A1(net6628),
    .S(_04968_),
    .X(_01500_));
 sg13g2_mux2_1 _22104_ (.A0(net5098),
    .A1(net4249),
    .S(_04968_),
    .X(_01501_));
 sg13g2_mux2_1 _22105_ (.A0(net5193),
    .A1(net6508),
    .S(_04968_),
    .X(_01502_));
 sg13g2_mux2_1 _22106_ (.A0(net5165),
    .A1(net6633),
    .S(_04968_),
    .X(_01503_));
 sg13g2_mux2_1 _22107_ (.A0(net5072),
    .A1(net6059),
    .S(_04968_),
    .X(_01504_));
 sg13g2_mux2_1 _22108_ (.A0(net5050),
    .A1(net6527),
    .S(_04968_),
    .X(_01505_));
 sg13g2_nand2_2 _22109_ (.Y(_04969_),
    .A(net4734),
    .B(_04956_));
 sg13g2_mux2_1 _22110_ (.A0(net5256),
    .A1(net4074),
    .S(_04969_),
    .X(_01506_));
 sg13g2_mux2_1 _22111_ (.A0(net5229),
    .A1(net4153),
    .S(_04969_),
    .X(_01507_));
 sg13g2_mux2_1 _22112_ (.A0(net5126),
    .A1(net4185),
    .S(_04969_),
    .X(_01508_));
 sg13g2_mux2_1 _22113_ (.A0(net5098),
    .A1(net4203),
    .S(_04969_),
    .X(_01509_));
 sg13g2_mux2_1 _22114_ (.A0(net5192),
    .A1(net4186),
    .S(_04969_),
    .X(_01510_));
 sg13g2_mux2_1 _22115_ (.A0(net5167),
    .A1(net4401),
    .S(_04969_),
    .X(_01511_));
 sg13g2_mux2_1 _22116_ (.A0(net5073),
    .A1(net4451),
    .S(_04969_),
    .X(_01512_));
 sg13g2_mux2_1 _22117_ (.A0(net5051),
    .A1(net4071),
    .S(_04969_),
    .X(_01513_));
 sg13g2_nor3_1 _22118_ (.A(net5037),
    .B(net4743),
    .C(_03164_),
    .Y(_04970_));
 sg13g2_nor2_1 _22119_ (.A(net3807),
    .B(net4692),
    .Y(_04971_));
 sg13g2_a21oi_1 _22120_ (.A1(net5262),
    .A2(net4692),
    .Y(_01514_),
    .B1(_04971_));
 sg13g2_nor2_1 _22121_ (.A(net3096),
    .B(net4691),
    .Y(_04972_));
 sg13g2_a21oi_1 _22122_ (.A1(net5234),
    .A2(net4691),
    .Y(_01515_),
    .B1(_04972_));
 sg13g2_nor2_1 _22123_ (.A(net3901),
    .B(net4691),
    .Y(_04973_));
 sg13g2_a21oi_1 _22124_ (.A1(net5132),
    .A2(net4691),
    .Y(_01516_),
    .B1(_04973_));
 sg13g2_nor2_1 _22125_ (.A(net3029),
    .B(net4691),
    .Y(_04974_));
 sg13g2_a21oi_1 _22126_ (.A1(net5103),
    .A2(net4691),
    .Y(_01517_),
    .B1(_04974_));
 sg13g2_nor2_1 _22127_ (.A(net3295),
    .B(net4692),
    .Y(_04975_));
 sg13g2_a21oi_1 _22128_ (.A1(net5176),
    .A2(net4692),
    .Y(_01518_),
    .B1(_04975_));
 sg13g2_nor2_1 _22129_ (.A(net4001),
    .B(net4691),
    .Y(_04976_));
 sg13g2_a21oi_1 _22130_ (.A1(net5147),
    .A2(net4691),
    .Y(_01519_),
    .B1(_04976_));
 sg13g2_nor2_1 _22131_ (.A(net3231),
    .B(net4692),
    .Y(_04977_));
 sg13g2_a21oi_1 _22132_ (.A1(net5079),
    .A2(net4692),
    .Y(_01520_),
    .B1(_04977_));
 sg13g2_nor2_1 _22133_ (.A(net3325),
    .B(net4692),
    .Y(_04978_));
 sg13g2_a21oi_1 _22134_ (.A1(net5056),
    .A2(net4692),
    .Y(_01521_),
    .B1(_04978_));
 sg13g2_nor2b_1 _22135_ (.A(net4742),
    .B_N(_04956_),
    .Y(_04979_));
 sg13g2_nor2_1 _22136_ (.A(net3669),
    .B(net4689),
    .Y(_04980_));
 sg13g2_a21oi_1 _22137_ (.A1(net5264),
    .A2(net4689),
    .Y(_01522_),
    .B1(_04980_));
 sg13g2_nor2_1 _22138_ (.A(net3143),
    .B(net4689),
    .Y(_04981_));
 sg13g2_a21oi_1 _22139_ (.A1(net5239),
    .A2(net4689),
    .Y(_01523_),
    .B1(_04981_));
 sg13g2_nor2_1 _22140_ (.A(net3339),
    .B(net4689),
    .Y(_04982_));
 sg13g2_a21oi_1 _22141_ (.A1(net5135),
    .A2(net4689),
    .Y(_01524_),
    .B1(_04982_));
 sg13g2_nor2_1 _22142_ (.A(net3662),
    .B(net4690),
    .Y(_04983_));
 sg13g2_a21oi_1 _22143_ (.A1(net5112),
    .A2(net4690),
    .Y(_01525_),
    .B1(_04983_));
 sg13g2_nor2_1 _22144_ (.A(net3129),
    .B(net4690),
    .Y(_04984_));
 sg13g2_a21oi_1 _22145_ (.A1(net5180),
    .A2(net4690),
    .Y(_01526_),
    .B1(_04984_));
 sg13g2_nor2_1 _22146_ (.A(net3166),
    .B(net4689),
    .Y(_04985_));
 sg13g2_a21oi_1 _22147_ (.A1(net5150),
    .A2(net4689),
    .Y(_01527_),
    .B1(_04985_));
 sg13g2_nor2_1 _22148_ (.A(net3281),
    .B(net4690),
    .Y(_04986_));
 sg13g2_a21oi_1 _22149_ (.A1(net5083),
    .A2(net4690),
    .Y(_01528_),
    .B1(_04986_));
 sg13g2_nor2_1 _22150_ (.A(net4003),
    .B(net4690),
    .Y(_04987_));
 sg13g2_a21oi_1 _22151_ (.A1(net5063),
    .A2(net4690),
    .Y(_01529_),
    .B1(_04987_));
 sg13g2_nand2_2 _22152_ (.Y(_04988_),
    .A(net4747),
    .B(_04956_));
 sg13g2_mux2_1 _22153_ (.A0(net5256),
    .A1(net6061),
    .S(_04988_),
    .X(_01530_));
 sg13g2_mux2_1 _22154_ (.A0(net5229),
    .A1(net6966),
    .S(_04988_),
    .X(_01531_));
 sg13g2_mux2_1 _22155_ (.A0(net5126),
    .A1(net4349),
    .S(_04988_),
    .X(_01532_));
 sg13g2_mux2_1 _22156_ (.A0(net5098),
    .A1(net4345),
    .S(_04988_),
    .X(_01533_));
 sg13g2_mux2_1 _22157_ (.A0(net5192),
    .A1(net6814),
    .S(_04988_),
    .X(_01534_));
 sg13g2_mux2_1 _22158_ (.A0(net5167),
    .A1(net4423),
    .S(_04988_),
    .X(_01535_));
 sg13g2_mux2_1 _22159_ (.A0(net5073),
    .A1(net6142),
    .S(_04988_),
    .X(_01536_));
 sg13g2_mux2_1 _22160_ (.A0(net5051),
    .A1(net6276),
    .S(_04988_),
    .X(_01537_));
 sg13g2_nor3_2 _22161_ (.A(net4878),
    .B(net5024),
    .C(_03002_),
    .Y(_04989_));
 sg13g2_nand2_2 _22162_ (.Y(_04990_),
    .A(net4739),
    .B(_04989_));
 sg13g2_mux2_1 _22163_ (.A0(net5246),
    .A1(net6198),
    .S(_04990_),
    .X(_01538_));
 sg13g2_mux2_1 _22164_ (.A0(net5220),
    .A1(net4247),
    .S(_04990_),
    .X(_01539_));
 sg13g2_mux2_1 _22165_ (.A0(net5121),
    .A1(net6560),
    .S(_04990_),
    .X(_01540_));
 sg13g2_mux2_1 _22166_ (.A0(net5092),
    .A1(net4173),
    .S(_04990_),
    .X(_01541_));
 sg13g2_mux2_1 _22167_ (.A0(net5192),
    .A1(net4310),
    .S(_04990_),
    .X(_01542_));
 sg13g2_mux2_1 _22168_ (.A0(net5165),
    .A1(net4371),
    .S(_04990_),
    .X(_01543_));
 sg13g2_mux2_1 _22169_ (.A0(net5074),
    .A1(net4209),
    .S(_04990_),
    .X(_01544_));
 sg13g2_mux2_1 _22170_ (.A0(net5049),
    .A1(net6051),
    .S(_04990_),
    .X(_01545_));
 sg13g2_nand2_2 _22171_ (.Y(_04991_),
    .A(net4736),
    .B(_04989_));
 sg13g2_mux2_1 _22172_ (.A0(net5246),
    .A1(net6516),
    .S(_04991_),
    .X(_01546_));
 sg13g2_mux2_1 _22173_ (.A0(net5220),
    .A1(net4000),
    .S(_04991_),
    .X(_01547_));
 sg13g2_mux2_1 _22174_ (.A0(net5121),
    .A1(net4176),
    .S(_04991_),
    .X(_01548_));
 sg13g2_mux2_1 _22175_ (.A0(net5092),
    .A1(net6124),
    .S(_04991_),
    .X(_01549_));
 sg13g2_mux2_1 _22176_ (.A0(net5192),
    .A1(net4077),
    .S(_04991_),
    .X(_01550_));
 sg13g2_mux2_1 _22177_ (.A0(net5165),
    .A1(net4534),
    .S(_04991_),
    .X(_01551_));
 sg13g2_mux2_1 _22178_ (.A0(net5074),
    .A1(net4120),
    .S(_04991_),
    .X(_01552_));
 sg13g2_mux2_1 _22179_ (.A0(net5049),
    .A1(net6702),
    .S(_04991_),
    .X(_01553_));
 sg13g2_nor2b_1 _22180_ (.A(net4744),
    .B_N(_04989_),
    .Y(_04992_));
 sg13g2_nor2_1 _22181_ (.A(net3703),
    .B(net4688),
    .Y(_04993_));
 sg13g2_a21oi_1 _22182_ (.A1(net5264),
    .A2(net4688),
    .Y(_01554_),
    .B1(_04993_));
 sg13g2_nor2_1 _22183_ (.A(net3500),
    .B(net4688),
    .Y(_04994_));
 sg13g2_a21oi_1 _22184_ (.A1(net5239),
    .A2(net4688),
    .Y(_01555_),
    .B1(_04994_));
 sg13g2_nor2_1 _22185_ (.A(net3426),
    .B(net4687),
    .Y(_04995_));
 sg13g2_a21oi_1 _22186_ (.A1(net5135),
    .A2(net4687),
    .Y(_01556_),
    .B1(_04995_));
 sg13g2_nor2_1 _22187_ (.A(net3604),
    .B(net4687),
    .Y(_04996_));
 sg13g2_a21oi_1 _22188_ (.A1(net5107),
    .A2(net4687),
    .Y(_01557_),
    .B1(_04996_));
 sg13g2_nor2_1 _22189_ (.A(net3778),
    .B(net4687),
    .Y(_04997_));
 sg13g2_a21oi_1 _22190_ (.A1(net5180),
    .A2(net4687),
    .Y(_01558_),
    .B1(_04997_));
 sg13g2_nor2_1 _22191_ (.A(net3724),
    .B(net4688),
    .Y(_04998_));
 sg13g2_a21oi_1 _22192_ (.A1(net5150),
    .A2(net4688),
    .Y(_01559_),
    .B1(_04998_));
 sg13g2_nor2_1 _22193_ (.A(net3245),
    .B(net4688),
    .Y(_04999_));
 sg13g2_a21oi_1 _22194_ (.A1(net5083),
    .A2(net4688),
    .Y(_01560_),
    .B1(_04999_));
 sg13g2_nor2_1 _22195_ (.A(net4057),
    .B(net4687),
    .Y(_05000_));
 sg13g2_a21oi_1 _22196_ (.A1(net5059),
    .A2(net4687),
    .Y(_01561_),
    .B1(_05000_));
 sg13g2_nand2_2 _22197_ (.Y(_05001_),
    .A(net4745),
    .B(_04989_));
 sg13g2_mux2_1 _22198_ (.A0(net5246),
    .A1(net6901),
    .S(_05001_),
    .X(_01562_));
 sg13g2_mux2_1 _22199_ (.A0(net5228),
    .A1(net6640),
    .S(_05001_),
    .X(_01563_));
 sg13g2_mux2_1 _22200_ (.A0(net5121),
    .A1(net6218),
    .S(_05001_),
    .X(_01564_));
 sg13g2_mux2_1 _22201_ (.A0(net5091),
    .A1(net6365),
    .S(_05001_),
    .X(_01565_));
 sg13g2_mux2_1 _22202_ (.A0(net5192),
    .A1(net6422),
    .S(_05001_),
    .X(_01566_));
 sg13g2_mux2_1 _22203_ (.A0(net5165),
    .A1(net4299),
    .S(_05001_),
    .X(_01567_));
 sg13g2_mux2_1 _22204_ (.A0(net5074),
    .A1(net6513),
    .S(_05001_),
    .X(_01568_));
 sg13g2_mux2_1 _22205_ (.A0(net5049),
    .A1(net6221),
    .S(_05001_),
    .X(_01569_));
 sg13g2_nand2_2 _22206_ (.Y(_05002_),
    .A(net4734),
    .B(_04989_));
 sg13g2_mux2_1 _22207_ (.A0(net5249),
    .A1(net6479),
    .S(_05002_),
    .X(_01570_));
 sg13g2_mux2_1 _22208_ (.A0(net5221),
    .A1(net4132),
    .S(_05002_),
    .X(_01571_));
 sg13g2_mux2_1 _22209_ (.A0(net5121),
    .A1(net4488),
    .S(_05002_),
    .X(_01572_));
 sg13g2_mux2_1 _22210_ (.A0(net5092),
    .A1(net4521),
    .S(_05002_),
    .X(_01573_));
 sg13g2_mux2_1 _22211_ (.A0(net5186),
    .A1(net4351),
    .S(_05002_),
    .X(_01574_));
 sg13g2_mux2_1 _22212_ (.A0(net5166),
    .A1(net6859),
    .S(_05002_),
    .X(_01575_));
 sg13g2_mux2_1 _22213_ (.A0(net5074),
    .A1(net6180),
    .S(_05002_),
    .X(_01576_));
 sg13g2_mux2_1 _22214_ (.A0(net5052),
    .A1(net4461),
    .S(_05002_),
    .X(_01577_));
 sg13g2_nand2_2 _22215_ (.Y(_05003_),
    .A(net4738),
    .B(_04989_));
 sg13g2_mux2_1 _22216_ (.A0(net5248),
    .A1(net4084),
    .S(_05003_),
    .X(_01578_));
 sg13g2_mux2_1 _22217_ (.A0(net5221),
    .A1(net4448),
    .S(_05003_),
    .X(_01579_));
 sg13g2_mux2_1 _22218_ (.A0(net5122),
    .A1(net4420),
    .S(_05003_),
    .X(_01580_));
 sg13g2_mux2_1 _22219_ (.A0(net5092),
    .A1(net4168),
    .S(_05003_),
    .X(_01581_));
 sg13g2_mux2_1 _22220_ (.A0(net5186),
    .A1(net4365),
    .S(_05003_),
    .X(_01582_));
 sg13g2_mux2_1 _22221_ (.A0(net5166),
    .A1(net6487),
    .S(_05003_),
    .X(_01583_));
 sg13g2_mux2_1 _22222_ (.A0(net5068),
    .A1(net6104),
    .S(_05003_),
    .X(_01584_));
 sg13g2_mux2_1 _22223_ (.A0(net5052),
    .A1(net6176),
    .S(_05003_),
    .X(_01585_));
 sg13g2_nor2b_1 _22224_ (.A(net4742),
    .B_N(_04989_),
    .Y(_05004_));
 sg13g2_nor2_1 _22225_ (.A(net3123),
    .B(net4686),
    .Y(_05005_));
 sg13g2_a21oi_1 _22226_ (.A1(net5263),
    .A2(net4686),
    .Y(_01586_),
    .B1(_05005_));
 sg13g2_nor2_1 _22227_ (.A(net3621),
    .B(net4685),
    .Y(_05006_));
 sg13g2_a21oi_1 _22228_ (.A1(net5239),
    .A2(net4685),
    .Y(_01587_),
    .B1(_05006_));
 sg13g2_nor2_1 _22229_ (.A(net3840),
    .B(net4686),
    .Y(_05007_));
 sg13g2_a21oi_1 _22230_ (.A1(net5131),
    .A2(net4686),
    .Y(_01588_),
    .B1(_05007_));
 sg13g2_nor2_1 _22231_ (.A(net3298),
    .B(net4686),
    .Y(_05008_));
 sg13g2_a21oi_1 _22232_ (.A1(net5103),
    .A2(net4686),
    .Y(_01589_),
    .B1(_05008_));
 sg13g2_nor2_1 _22233_ (.A(net3909),
    .B(net4685),
    .Y(_05009_));
 sg13g2_a21oi_1 _22234_ (.A1(net5175),
    .A2(net4685),
    .Y(_01590_),
    .B1(_05009_));
 sg13g2_nor2_1 _22235_ (.A(net3136),
    .B(net4685),
    .Y(_05010_));
 sg13g2_a21oi_1 _22236_ (.A1(net5150),
    .A2(net4685),
    .Y(_01591_),
    .B1(_05010_));
 sg13g2_nor2_1 _22237_ (.A(net6391),
    .B(net4686),
    .Y(_05011_));
 sg13g2_a21oi_1 _22238_ (.A1(net5080),
    .A2(_05004_),
    .Y(_01592_),
    .B1(_05011_));
 sg13g2_nor2_1 _22239_ (.A(net3812),
    .B(net4685),
    .Y(_05012_));
 sg13g2_a21oi_1 _22240_ (.A1(net5059),
    .A2(net4685),
    .Y(_01593_),
    .B1(_05012_));
 sg13g2_nand2_2 _22241_ (.Y(_05013_),
    .A(net4745),
    .B(_03165_));
 sg13g2_mux2_1 _22242_ (.A0(net5244),
    .A1(net4398),
    .S(_05013_),
    .X(_01594_));
 sg13g2_mux2_1 _22243_ (.A0(net5219),
    .A1(net6820),
    .S(_05013_),
    .X(_01595_));
 sg13g2_mux2_1 _22244_ (.A0(net5116),
    .A1(net6468),
    .S(_05013_),
    .X(_01596_));
 sg13g2_mux2_1 _22245_ (.A0(net5090),
    .A1(net6296),
    .S(_05013_),
    .X(_01597_));
 sg13g2_mux2_1 _22246_ (.A0(net5185),
    .A1(net6721),
    .S(_05013_),
    .X(_01598_));
 sg13g2_mux2_1 _22247_ (.A0(net5157),
    .A1(net6736),
    .S(_05013_),
    .X(_01599_));
 sg13g2_mux2_1 _22248_ (.A0(net5065),
    .A1(net6251),
    .S(_05013_),
    .X(_01600_));
 sg13g2_mux2_1 _22249_ (.A0(net5042),
    .A1(net4182),
    .S(_05013_),
    .X(_01601_));
 sg13g2_nand2_2 _22250_ (.Y(_05014_),
    .A(net4740),
    .B(_04811_));
 sg13g2_mux2_1 _22251_ (.A0(net5248),
    .A1(net4178),
    .S(_05014_),
    .X(_01602_));
 sg13g2_mux2_1 _22252_ (.A0(net5221),
    .A1(net4248),
    .S(_05014_),
    .X(_01603_));
 sg13g2_mux2_1 _22253_ (.A0(net5122),
    .A1(net4256),
    .S(_05014_),
    .X(_01604_));
 sg13g2_mux2_1 _22254_ (.A0(net5095),
    .A1(net4514),
    .S(_05014_),
    .X(_01605_));
 sg13g2_mux2_1 _22255_ (.A0(net5192),
    .A1(net4316),
    .S(_05014_),
    .X(_01606_));
 sg13g2_mux2_1 _22256_ (.A0(net5166),
    .A1(net4542),
    .S(_05014_),
    .X(_01607_));
 sg13g2_mux2_1 _22257_ (.A0(net5074),
    .A1(net4133),
    .S(_05014_),
    .X(_01608_));
 sg13g2_mux2_1 _22258_ (.A0(net5049),
    .A1(net4261),
    .S(_05014_),
    .X(_01609_));
 sg13g2_nand2_2 _22259_ (.Y(_05015_),
    .A(net4746),
    .B(_04811_));
 sg13g2_mux2_1 _22260_ (.A0(net5248),
    .A1(net6279),
    .S(_05015_),
    .X(_01610_));
 sg13g2_mux2_1 _22261_ (.A0(net5221),
    .A1(net4252),
    .S(_05015_),
    .X(_01611_));
 sg13g2_mux2_1 _22262_ (.A0(net5122),
    .A1(net6655),
    .S(_05015_),
    .X(_01612_));
 sg13g2_mux2_1 _22263_ (.A0(net5095),
    .A1(net6121),
    .S(_05015_),
    .X(_01613_));
 sg13g2_mux2_1 _22264_ (.A0(net5192),
    .A1(net6676),
    .S(_05015_),
    .X(_01614_));
 sg13g2_mux2_1 _22265_ (.A0(net5166),
    .A1(net6607),
    .S(_05015_),
    .X(_01615_));
 sg13g2_mux2_1 _22266_ (.A0(net5074),
    .A1(net6521),
    .S(_05015_),
    .X(_01616_));
 sg13g2_mux2_1 _22267_ (.A0(net5049),
    .A1(net6437),
    .S(_05015_),
    .X(_01617_));
 sg13g2_nand2_2 _22268_ (.Y(_05016_),
    .A(net4736),
    .B(_04811_));
 sg13g2_mux2_1 _22269_ (.A0(net5256),
    .A1(net4529),
    .S(_05016_),
    .X(_01618_));
 sg13g2_mux2_1 _22270_ (.A0(net5230),
    .A1(net6102),
    .S(_05016_),
    .X(_01619_));
 sg13g2_mux2_1 _22271_ (.A0(net5127),
    .A1(net6578),
    .S(_05016_),
    .X(_01620_));
 sg13g2_mux2_1 _22272_ (.A0(net5100),
    .A1(net4226),
    .S(_05016_),
    .X(_01621_));
 sg13g2_mux2_1 _22273_ (.A0(net5195),
    .A1(net6467),
    .S(_05016_),
    .X(_01622_));
 sg13g2_mux2_1 _22274_ (.A0(net5166),
    .A1(net4044),
    .S(_05016_),
    .X(_01623_));
 sg13g2_mux2_1 _22275_ (.A0(net5074),
    .A1(net4078),
    .S(_05016_),
    .X(_01624_));
 sg13g2_mux2_1 _22276_ (.A0(net5049),
    .A1(net4050),
    .S(_05016_),
    .X(_01625_));
 sg13g2_nor2b_1 _22277_ (.A(net4744),
    .B_N(_04811_),
    .Y(_05017_));
 sg13g2_nor2_1 _22278_ (.A(net3720),
    .B(net4684),
    .Y(_05018_));
 sg13g2_a21oi_1 _22279_ (.A1(net5264),
    .A2(net4684),
    .Y(_01626_),
    .B1(_05018_));
 sg13g2_nor2_1 _22280_ (.A(net3854),
    .B(net4683),
    .Y(_05019_));
 sg13g2_a21oi_1 _22281_ (.A1(net5239),
    .A2(net4683),
    .Y(_01627_),
    .B1(_05019_));
 sg13g2_nor2_1 _22282_ (.A(net3126),
    .B(net4684),
    .Y(_05020_));
 sg13g2_a21oi_1 _22283_ (.A1(net5135),
    .A2(net4684),
    .Y(_01628_),
    .B1(_05020_));
 sg13g2_nor2_1 _22284_ (.A(net3032),
    .B(net4684),
    .Y(_05021_));
 sg13g2_a21oi_1 _22285_ (.A1(net5107),
    .A2(net4684),
    .Y(_01629_),
    .B1(_05021_));
 sg13g2_nor2_1 _22286_ (.A(net4210),
    .B(net4684),
    .Y(_05022_));
 sg13g2_a21oi_1 _22287_ (.A1(net5180),
    .A2(net4684),
    .Y(_01630_),
    .B1(_05022_));
 sg13g2_nor2_1 _22288_ (.A(net3895),
    .B(net4683),
    .Y(_05023_));
 sg13g2_a21oi_1 _22289_ (.A1(net5150),
    .A2(net4683),
    .Y(_01631_),
    .B1(_05023_));
 sg13g2_nor2_1 _22290_ (.A(net3566),
    .B(net4683),
    .Y(_05024_));
 sg13g2_a21oi_1 _22291_ (.A1(net5083),
    .A2(net4683),
    .Y(_01632_),
    .B1(_05024_));
 sg13g2_nor2_1 _22292_ (.A(net3041),
    .B(net4683),
    .Y(_05025_));
 sg13g2_a21oi_1 _22293_ (.A1(net5059),
    .A2(net4683),
    .Y(_01633_),
    .B1(_05025_));
 sg13g2_nor2_1 _22294_ (.A(net5577),
    .B(_08212_),
    .Y(_05026_));
 sg13g2_nand2_1 _22295_ (.Y(_05027_),
    .A(\atari2600.cpu.load_reg ),
    .B(_05026_));
 sg13g2_a21oi_2 _22296_ (.B1(net5312),
    .Y(_05028_),
    .A2(_05027_),
    .A1(_08503_));
 sg13g2_nand2_2 _22297_ (.Y(_05029_),
    .A(_08512_),
    .B(_05028_));
 sg13g2_nor2_1 _22298_ (.A(net5572),
    .B(net5478),
    .Y(_05030_));
 sg13g2_a21oi_2 _22299_ (.B1(_05030_),
    .Y(_05031_),
    .A2(net5478),
    .A1(_08191_));
 sg13g2_mux2_1 _22300_ (.A0(_05031_),
    .A1(net3777),
    .S(_05029_),
    .X(_01634_));
 sg13g2_nor2_1 _22301_ (.A(\atari2600.cpu.adc_bcd ),
    .B(_00054_),
    .Y(_05032_));
 sg13g2_nand2b_1 _22302_ (.Y(_05033_),
    .B(_05032_),
    .A_N(\atari2600.cpu.ALU.HC ));
 sg13g2_nand2_1 _22303_ (.Y(_05034_),
    .A(\atari2600.cpu.adc_bcd ),
    .B(\atari2600.cpu.ALU.HC ));
 sg13g2_o21ai_1 _22304_ (.B1(_05033_),
    .Y(_05035_),
    .A1(_00054_),
    .A2(_05034_));
 sg13g2_xnor2_1 _22305_ (.Y(_05036_),
    .A(_00097_),
    .B(_05035_));
 sg13g2_nor2_1 _22306_ (.A(net5478),
    .B(_05036_),
    .Y(_05037_));
 sg13g2_a21oi_2 _22307_ (.B1(_05037_),
    .Y(_05038_),
    .A2(net5478),
    .A1(_08187_));
 sg13g2_mux2_1 _22308_ (.A0(_05038_),
    .A1(net3492),
    .S(_05029_),
    .X(_01635_));
 sg13g2_nand3_1 _22309_ (.B(\atari2600.cpu.adj_bcd ),
    .C(\atari2600.cpu.ALU.HC ),
    .A(\atari2600.cpu.adc_bcd ),
    .Y(_05039_));
 sg13g2_xnor2_1 _22310_ (.Y(_05040_),
    .A(net5571),
    .B(_05039_));
 sg13g2_nand3_1 _22311_ (.B(_05035_),
    .C(_05040_),
    .A(\atari2600.cpu.ADD[1] ),
    .Y(_05041_));
 sg13g2_a21o_1 _22312_ (.A2(_05035_),
    .A1(\atari2600.cpu.ADD[1] ),
    .B1(_05040_),
    .X(_05042_));
 sg13g2_nand3_1 _22313_ (.B(_05041_),
    .C(_05042_),
    .A(net5476),
    .Y(_05043_));
 sg13g2_o21ai_1 _22314_ (.B1(_05043_),
    .Y(_05044_),
    .A1(_08201_),
    .A2(net5476));
 sg13g2_mux2_1 _22315_ (.A0(_05044_),
    .A1(net4392),
    .S(_05029_),
    .X(_01636_));
 sg13g2_o21ai_1 _22316_ (.B1(_05041_),
    .Y(_05045_),
    .A1(_08057_),
    .A2(_05039_));
 sg13g2_xnor2_1 _22317_ (.Y(_05046_),
    .A(_00101_),
    .B(_05033_));
 sg13g2_xnor2_1 _22318_ (.Y(_05047_),
    .A(_05045_),
    .B(_05046_));
 sg13g2_nand2_1 _22319_ (.Y(_05048_),
    .A(net5476),
    .B(_05047_));
 sg13g2_o21ai_1 _22320_ (.B1(_05048_),
    .Y(_05049_),
    .A1(_08196_),
    .A2(net5476));
 sg13g2_mux2_1 _22321_ (.A0(_05049_),
    .A1(net6849),
    .S(_05029_),
    .X(_01637_));
 sg13g2_nor2_1 _22322_ (.A(net5570),
    .B(net5478),
    .Y(_05050_));
 sg13g2_a21oi_2 _22323_ (.B1(_05050_),
    .Y(_05051_),
    .A2(net5478),
    .A1(_08181_));
 sg13g2_mux2_1 _22324_ (.A0(_05051_),
    .A1(net4313),
    .S(_05029_),
    .X(_01638_));
 sg13g2_nand2_1 _22325_ (.Y(_05052_),
    .A(net5351),
    .B(net5478));
 sg13g2_nand2_1 _22326_ (.Y(_05053_),
    .A(\atari2600.cpu.ALU.CO ),
    .B(\atari2600.cpu.adc_bcd ));
 sg13g2_nand2_1 _22327_ (.Y(_05054_),
    .A(_08070_),
    .B(_05032_));
 sg13g2_o21ai_1 _22328_ (.B1(_05054_),
    .Y(_05055_),
    .A1(_00054_),
    .A2(_05053_));
 sg13g2_xnor2_1 _22329_ (.Y(_05056_),
    .A(_08076_),
    .B(_05055_));
 sg13g2_o21ai_1 _22330_ (.B1(_05052_),
    .Y(_05057_),
    .A1(net5478),
    .A2(_05056_));
 sg13g2_mux2_1 _22331_ (.A0(_05057_),
    .A1(net4109),
    .S(_05029_),
    .X(_01639_));
 sg13g2_nand3_1 _22332_ (.B(\atari2600.cpu.adc_bcd ),
    .C(\atari2600.cpu.adj_bcd ),
    .A(\atari2600.cpu.ALU.CO ),
    .Y(_05058_));
 sg13g2_xnor2_1 _22333_ (.Y(_05059_),
    .A(net5568),
    .B(_05058_));
 sg13g2_a21o_1 _22334_ (.A2(_05055_),
    .A1(net5569),
    .B1(_05059_),
    .X(_05060_));
 sg13g2_nand3_1 _22335_ (.B(_05055_),
    .C(_05059_),
    .A(net5569),
    .Y(_05061_));
 sg13g2_nand3_1 _22336_ (.B(_05060_),
    .C(_05061_),
    .A(net5476),
    .Y(_05062_));
 sg13g2_o21ai_1 _22337_ (.B1(_05062_),
    .Y(_05063_),
    .A1(_08244_),
    .A2(net5476));
 sg13g2_mux2_1 _22338_ (.A0(_05063_),
    .A1(net6455),
    .S(_05029_),
    .X(_01640_));
 sg13g2_nor2_1 _22339_ (.A(net5273),
    .B(net5476),
    .Y(_05064_));
 sg13g2_o21ai_1 _22340_ (.B1(_05061_),
    .Y(_05065_),
    .A1(_08072_),
    .A2(_05058_));
 sg13g2_xor2_1 _22341_ (.B(_05054_),
    .A(_00104_),
    .X(_05066_));
 sg13g2_xnor2_1 _22342_ (.Y(_05067_),
    .A(_05065_),
    .B(_05066_));
 sg13g2_a21oi_2 _22343_ (.B1(_05064_),
    .Y(_05068_),
    .A2(_05067_),
    .A1(net5476));
 sg13g2_mux2_1 _22344_ (.A0(_05068_),
    .A1(net6240),
    .S(_05029_),
    .X(_01641_));
 sg13g2_nand2_2 _22345_ (.Y(_05069_),
    .A(net4746),
    .B(net4763));
 sg13g2_mux2_1 _22346_ (.A0(net5253),
    .A1(net4468),
    .S(_05069_),
    .X(_01642_));
 sg13g2_mux2_1 _22347_ (.A0(net5223),
    .A1(net6098),
    .S(_05069_),
    .X(_01643_));
 sg13g2_mux2_1 _22348_ (.A0(net5118),
    .A1(net6501),
    .S(_05069_),
    .X(_01644_));
 sg13g2_mux2_1 _22349_ (.A0(net5095),
    .A1(net4446),
    .S(_05069_),
    .X(_01645_));
 sg13g2_mux2_1 _22350_ (.A0(net5189),
    .A1(net4445),
    .S(_05069_),
    .X(_01646_));
 sg13g2_mux2_1 _22351_ (.A0(net5162),
    .A1(net6166),
    .S(_05069_),
    .X(_01647_));
 sg13g2_mux2_1 _22352_ (.A0(net5070),
    .A1(net6431),
    .S(_05069_),
    .X(_01648_));
 sg13g2_mux2_1 _22353_ (.A0(net5046),
    .A1(net6555),
    .S(_05069_),
    .X(_01649_));
 sg13g2_nand2_2 _22354_ (.Y(_05070_),
    .A(_03041_),
    .B(net4737));
 sg13g2_mux2_1 _22355_ (.A0(net5251),
    .A1(net6118),
    .S(_05070_),
    .X(_01650_));
 sg13g2_mux2_1 _22356_ (.A0(net5225),
    .A1(net4381),
    .S(_05070_),
    .X(_01651_));
 sg13g2_mux2_1 _22357_ (.A0(net5124),
    .A1(net4154),
    .S(_05070_),
    .X(_01652_));
 sg13g2_mux2_1 _22358_ (.A0(net5096),
    .A1(net3996),
    .S(_05070_),
    .X(_01653_));
 sg13g2_mux2_1 _22359_ (.A0(net5191),
    .A1(net4236),
    .S(_05070_),
    .X(_01654_));
 sg13g2_mux2_1 _22360_ (.A0(net5163),
    .A1(net4038),
    .S(_05070_),
    .X(_01655_));
 sg13g2_mux2_1 _22361_ (.A0(net5071),
    .A1(net6082),
    .S(_05070_),
    .X(_01656_));
 sg13g2_mux2_1 _22362_ (.A0(net5045),
    .A1(net4453),
    .S(_05070_),
    .X(_01657_));
 sg13g2_nor3_2 _22363_ (.A(net4876),
    .B(net5021),
    .C(_10253_),
    .Y(_05071_));
 sg13g2_nand2_2 _22364_ (.Y(_05072_),
    .A(net4748),
    .B(_05071_));
 sg13g2_mux2_1 _22365_ (.A0(net5245),
    .A1(net4361),
    .S(_05072_),
    .X(_01658_));
 sg13g2_mux2_1 _22366_ (.A0(net5218),
    .A1(net4269),
    .S(_05072_),
    .X(_01659_));
 sg13g2_mux2_1 _22367_ (.A0(net5115),
    .A1(net4388),
    .S(_05072_),
    .X(_01660_));
 sg13g2_mux2_1 _22368_ (.A0(net5088),
    .A1(net4228),
    .S(_05072_),
    .X(_01661_));
 sg13g2_mux2_1 _22369_ (.A0(net5185),
    .A1(net4238),
    .S(_05072_),
    .X(_01662_));
 sg13g2_mux2_1 _22370_ (.A0(net5158),
    .A1(net6807),
    .S(_05072_),
    .X(_01663_));
 sg13g2_mux2_1 _22371_ (.A0(net5064),
    .A1(net4470),
    .S(_05072_),
    .X(_01664_));
 sg13g2_mux2_1 _22372_ (.A0(net5040),
    .A1(net4263),
    .S(_05072_),
    .X(_01665_));
 sg13g2_nor3_2 _22373_ (.A(net4878),
    .B(net5020),
    .C(_03002_),
    .Y(_05073_));
 sg13g2_nand2_2 _22374_ (.Y(_05074_),
    .A(net4735),
    .B(_05073_));
 sg13g2_mux2_1 _22375_ (.A0(net5248),
    .A1(net4083),
    .S(_05074_),
    .X(_01666_));
 sg13g2_mux2_1 _22376_ (.A0(net5221),
    .A1(net4315),
    .S(_05074_),
    .X(_01667_));
 sg13g2_mux2_1 _22377_ (.A0(net5120),
    .A1(net4130),
    .S(_05074_),
    .X(_01668_));
 sg13g2_mux2_1 _22378_ (.A0(net5097),
    .A1(net4035),
    .S(_05074_),
    .X(_01669_));
 sg13g2_mux2_1 _22379_ (.A0(net5187),
    .A1(net4030),
    .S(_05074_),
    .X(_01670_));
 sg13g2_mux2_1 _22380_ (.A0(net5159),
    .A1(net4408),
    .S(_05074_),
    .X(_01671_));
 sg13g2_mux2_1 _22381_ (.A0(net5066),
    .A1(net6310),
    .S(_05074_),
    .X(_01672_));
 sg13g2_mux2_1 _22382_ (.A0(net5044),
    .A1(net4042),
    .S(_05074_),
    .X(_01673_));
 sg13g2_nor4_2 _22383_ (.A(net5037),
    .B(net4876),
    .C(net5025),
    .Y(_05075_),
    .D(net5021));
 sg13g2_nand2_2 _22384_ (.Y(_05076_),
    .A(net4745),
    .B(_05075_));
 sg13g2_mux2_1 _22385_ (.A0(net5247),
    .A1(net6283),
    .S(_05076_),
    .X(_01674_));
 sg13g2_mux2_1 _22386_ (.A0(net5220),
    .A1(net6761),
    .S(_05076_),
    .X(_01675_));
 sg13g2_mux2_1 _22387_ (.A0(net5120),
    .A1(net4412),
    .S(_05076_),
    .X(_01676_));
 sg13g2_mux2_1 _22388_ (.A0(net5091),
    .A1(net4508),
    .S(_05076_),
    .X(_01677_));
 sg13g2_mux2_1 _22389_ (.A0(net5186),
    .A1(net4334),
    .S(_05076_),
    .X(_01678_));
 sg13g2_mux2_1 _22390_ (.A0(net5160),
    .A1(net6679),
    .S(_05076_),
    .X(_01679_));
 sg13g2_mux2_1 _22391_ (.A0(net5067),
    .A1(net4204),
    .S(_05076_),
    .X(_01680_));
 sg13g2_mux2_1 _22392_ (.A0(net5043),
    .A1(net4356),
    .S(_05076_),
    .X(_01681_));
 sg13g2_nand2_2 _22393_ (.Y(_05077_),
    .A(_03059_),
    .B(net4738));
 sg13g2_mux2_1 _22394_ (.A0(net5258),
    .A1(net4116),
    .S(_05077_),
    .X(_01682_));
 sg13g2_mux2_1 _22395_ (.A0(net5231),
    .A1(net4274),
    .S(_05077_),
    .X(_01683_));
 sg13g2_mux2_1 _22396_ (.A0(net5128),
    .A1(net4052),
    .S(_05077_),
    .X(_01684_));
 sg13g2_mux2_1 _22397_ (.A0(net5100),
    .A1(net6423),
    .S(_05077_),
    .X(_01685_));
 sg13g2_mux2_1 _22398_ (.A0(net5195),
    .A1(net4438),
    .S(_05077_),
    .X(_01686_));
 sg13g2_mux2_1 _22399_ (.A0(net5171),
    .A1(net6492),
    .S(_05077_),
    .X(_01687_));
 sg13g2_mux2_1 _22400_ (.A0(net5076),
    .A1(net4494),
    .S(_05077_),
    .X(_01688_));
 sg13g2_mux2_1 _22401_ (.A0(net5054),
    .A1(net4054),
    .S(_05077_),
    .X(_01689_));
 sg13g2_and2_1 _22402_ (.A(net4747),
    .B(_03087_),
    .X(_05078_));
 sg13g2_nor2_1 _22403_ (.A(net3024),
    .B(net4681),
    .Y(_05079_));
 sg13g2_a21oi_1 _22404_ (.A1(net5267),
    .A2(net4681),
    .Y(_01690_),
    .B1(_05079_));
 sg13g2_nor2_1 _22405_ (.A(net3199),
    .B(net4682),
    .Y(_05080_));
 sg13g2_a21oi_1 _22406_ (.A1(net5241),
    .A2(net4682),
    .Y(_01691_),
    .B1(_05080_));
 sg13g2_nor2_1 _22407_ (.A(net3288),
    .B(net4681),
    .Y(_05081_));
 sg13g2_a21oi_1 _22408_ (.A1(net5137),
    .A2(net4681),
    .Y(_01692_),
    .B1(_05081_));
 sg13g2_nor2_1 _22409_ (.A(net3286),
    .B(net4682),
    .Y(_05082_));
 sg13g2_a21oi_1 _22410_ (.A1(net5108),
    .A2(net4682),
    .Y(_01693_),
    .B1(_05082_));
 sg13g2_nor2_1 _22411_ (.A(net3268),
    .B(_05078_),
    .Y(_05083_));
 sg13g2_a21oi_1 _22412_ (.A1(net5182),
    .A2(net4682),
    .Y(_01694_),
    .B1(_05083_));
 sg13g2_nor2_1 _22413_ (.A(net3918),
    .B(net4682),
    .Y(_05084_));
 sg13g2_a21oi_1 _22414_ (.A1(net5153),
    .A2(net4682),
    .Y(_01695_),
    .B1(_05084_));
 sg13g2_nor2_1 _22415_ (.A(net3853),
    .B(net4681),
    .Y(_05085_));
 sg13g2_a21oi_1 _22416_ (.A1(net5084),
    .A2(net4681),
    .Y(_01696_),
    .B1(_05085_));
 sg13g2_nor2_1 _22417_ (.A(net3100),
    .B(net4681),
    .Y(_05086_));
 sg13g2_a21oi_1 _22418_ (.A1(net5062),
    .A2(net4681),
    .Y(_01697_),
    .B1(_05086_));
 sg13g2_nor2_1 _22419_ (.A(_03166_),
    .B(_04893_),
    .Y(_05087_));
 sg13g2_nor2_1 _22420_ (.A(net3639),
    .B(net4680),
    .Y(_05088_));
 sg13g2_a21oi_1 _22421_ (.A1(net5261),
    .A2(net4680),
    .Y(_01698_),
    .B1(_05088_));
 sg13g2_nor2_1 _22422_ (.A(net3766),
    .B(net4680),
    .Y(_05089_));
 sg13g2_a21oi_1 _22423_ (.A1(net5236),
    .A2(net4680),
    .Y(_01699_),
    .B1(_05089_));
 sg13g2_nor2_1 _22424_ (.A(net2998),
    .B(net4680),
    .Y(_05090_));
 sg13g2_a21oi_1 _22425_ (.A1(net5133),
    .A2(net4680),
    .Y(_01700_),
    .B1(_05090_));
 sg13g2_nor2_1 _22426_ (.A(net3380),
    .B(net4680),
    .Y(_05091_));
 sg13g2_a21oi_1 _22427_ (.A1(net5109),
    .A2(net4680),
    .Y(_01701_),
    .B1(_05091_));
 sg13g2_nor2_1 _22428_ (.A(net2980),
    .B(net4679),
    .Y(_05092_));
 sg13g2_a21oi_1 _22429_ (.A1(net5177),
    .A2(net4679),
    .Y(_01702_),
    .B1(_05092_));
 sg13g2_nor2_1 _22430_ (.A(net3013),
    .B(net4679),
    .Y(_05093_));
 sg13g2_a21oi_1 _22431_ (.A1(net5148),
    .A2(net4679),
    .Y(_01703_),
    .B1(_05093_));
 sg13g2_nor2_1 _22432_ (.A(net3320),
    .B(net4679),
    .Y(_05094_));
 sg13g2_a21oi_1 _22433_ (.A1(net5081),
    .A2(net4679),
    .Y(_01704_),
    .B1(_05094_));
 sg13g2_nor2_1 _22434_ (.A(net3897),
    .B(net4679),
    .Y(_05095_));
 sg13g2_a21oi_1 _22435_ (.A1(net5057),
    .A2(net4679),
    .Y(_01705_),
    .B1(_05095_));
 sg13g2_nand2_2 _22436_ (.Y(_05096_),
    .A(net4745),
    .B(_04931_));
 sg13g2_mux2_1 _22437_ (.A0(net5255),
    .A1(net6318),
    .S(_05096_),
    .X(_01706_));
 sg13g2_mux2_1 _22438_ (.A0(net5228),
    .A1(net4473),
    .S(_05096_),
    .X(_01707_));
 sg13g2_mux2_1 _22439_ (.A0(net5127),
    .A1(net6175),
    .S(_05096_),
    .X(_01708_));
 sg13g2_mux2_1 _22440_ (.A0(net5098),
    .A1(net6146),
    .S(_05096_),
    .X(_01709_));
 sg13g2_mux2_1 _22441_ (.A0(net5193),
    .A1(net4429),
    .S(_05096_),
    .X(_01710_));
 sg13g2_mux2_1 _22442_ (.A0(net5165),
    .A1(net6395),
    .S(_05096_),
    .X(_01711_));
 sg13g2_mux2_1 _22443_ (.A0(net5072),
    .A1(net4509),
    .S(_05096_),
    .X(_01712_));
 sg13g2_mux2_1 _22444_ (.A0(net5051),
    .A1(net6885),
    .S(_05096_),
    .X(_01713_));
 sg13g2_nand2_2 _22445_ (.Y(_05097_),
    .A(net4738),
    .B(_04956_));
 sg13g2_mux2_1 _22446_ (.A0(net5256),
    .A1(net6210),
    .S(_05097_),
    .X(_01714_));
 sg13g2_mux2_1 _22447_ (.A0(net5229),
    .A1(net4212),
    .S(_05097_),
    .X(_01715_));
 sg13g2_mux2_1 _22448_ (.A0(net5126),
    .A1(net4093),
    .S(_05097_),
    .X(_01716_));
 sg13g2_mux2_1 _22449_ (.A0(net5099),
    .A1(net4213),
    .S(_05097_),
    .X(_01717_));
 sg13g2_mux2_1 _22450_ (.A0(net5194),
    .A1(net6073),
    .S(_05097_),
    .X(_01718_));
 sg13g2_mux2_1 _22451_ (.A0(net5166),
    .A1(net4137),
    .S(_05097_),
    .X(_01719_));
 sg13g2_mux2_1 _22452_ (.A0(net5073),
    .A1(net6057),
    .S(_05097_),
    .X(_01720_));
 sg13g2_mux2_1 _22453_ (.A0(net5051),
    .A1(net4047),
    .S(_05097_),
    .X(_01721_));
 sg13g2_nand2_2 _22454_ (.Y(_05098_),
    .A(net4747),
    .B(_04989_));
 sg13g2_mux2_1 _22455_ (.A0(net5249),
    .A1(net6504),
    .S(_05098_),
    .X(_01722_));
 sg13g2_mux2_1 _22456_ (.A0(net5221),
    .A1(net4060),
    .S(_05098_),
    .X(_01723_));
 sg13g2_mux2_1 _22457_ (.A0(net5121),
    .A1(net4459),
    .S(_05098_),
    .X(_01724_));
 sg13g2_mux2_1 _22458_ (.A0(net5092),
    .A1(net6494),
    .S(_05098_),
    .X(_01725_));
 sg13g2_mux2_1 _22459_ (.A0(net5186),
    .A1(net6434),
    .S(_05098_),
    .X(_01726_));
 sg13g2_mux2_1 _22460_ (.A0(net5166),
    .A1(net4245),
    .S(_05098_),
    .X(_01727_));
 sg13g2_mux2_1 _22461_ (.A0(net5074),
    .A1(net6117),
    .S(_05098_),
    .X(_01728_));
 sg13g2_mux2_1 _22462_ (.A0(net5052),
    .A1(net6260),
    .S(_05098_),
    .X(_01729_));
 sg13g2_nor2_1 _22463_ (.A(net4744),
    .B(_03088_),
    .Y(_05099_));
 sg13g2_nor2_1 _22464_ (.A(net3003),
    .B(_05099_),
    .Y(_05100_));
 sg13g2_a21oi_1 _22465_ (.A1(net5266),
    .A2(net4678),
    .Y(_01730_),
    .B1(_05100_));
 sg13g2_nor2_1 _22466_ (.A(net3267),
    .B(net4678),
    .Y(_05101_));
 sg13g2_a21oi_1 _22467_ (.A1(net5240),
    .A2(net4678),
    .Y(_01731_),
    .B1(_05101_));
 sg13g2_nor2_1 _22468_ (.A(net3837),
    .B(net4678),
    .Y(_05102_));
 sg13g2_a21oi_1 _22469_ (.A1(net5139),
    .A2(net4678),
    .Y(_01732_),
    .B1(_05102_));
 sg13g2_nor2_1 _22470_ (.A(net3095),
    .B(net4677),
    .Y(_05103_));
 sg13g2_a21oi_1 _22471_ (.A1(net5108),
    .A2(net4677),
    .Y(_01733_),
    .B1(_05103_));
 sg13g2_nor2_1 _22472_ (.A(net3078),
    .B(net4677),
    .Y(_05104_));
 sg13g2_a21oi_1 _22473_ (.A1(net5182),
    .A2(net4677),
    .Y(_01734_),
    .B1(_05104_));
 sg13g2_nor2_1 _22474_ (.A(net3855),
    .B(net4677),
    .Y(_05105_));
 sg13g2_a21oi_1 _22475_ (.A1(net5152),
    .A2(net4677),
    .Y(_01735_),
    .B1(_05105_));
 sg13g2_nor2_1 _22476_ (.A(net3318),
    .B(net4678),
    .Y(_05106_));
 sg13g2_a21oi_1 _22477_ (.A1(net5084),
    .A2(net4678),
    .Y(_01736_),
    .B1(_05106_));
 sg13g2_nor2_1 _22478_ (.A(net3508),
    .B(net4677),
    .Y(_05107_));
 sg13g2_a21oi_1 _22479_ (.A1(net5060),
    .A2(net4677),
    .Y(_01737_),
    .B1(_05107_));
 sg13g2_nand2_2 _22480_ (.Y(_05108_),
    .A(_03003_),
    .B(net4738));
 sg13g2_mux2_1 _22481_ (.A0(net5253),
    .A1(net4142),
    .S(_05108_),
    .X(_01738_));
 sg13g2_mux2_1 _22482_ (.A0(net5224),
    .A1(net4539),
    .S(_05108_),
    .X(_01739_));
 sg13g2_mux2_1 _22483_ (.A0(net5122),
    .A1(net4114),
    .S(_05108_),
    .X(_01740_));
 sg13g2_mux2_1 _22484_ (.A0(net5095),
    .A1(net4220),
    .S(_05108_),
    .X(_01741_));
 sg13g2_mux2_1 _22485_ (.A0(net5190),
    .A1(net6049),
    .S(_05108_),
    .X(_01742_));
 sg13g2_mux2_1 _22486_ (.A0(net5163),
    .A1(net4523),
    .S(_05108_),
    .X(_01743_));
 sg13g2_mux2_1 _22487_ (.A0(net5071),
    .A1(net6568),
    .S(_05108_),
    .X(_01744_));
 sg13g2_mux2_1 _22488_ (.A0(net5045),
    .A1(net4492),
    .S(_05108_),
    .X(_01745_));
 sg13g2_nor2b_1 _22489_ (.A(net4743),
    .B_N(_05071_),
    .Y(_05109_));
 sg13g2_nor2_1 _22490_ (.A(net4048),
    .B(net4675),
    .Y(_05110_));
 sg13g2_a21oi_1 _22491_ (.A1(net5260),
    .A2(net4675),
    .Y(_01746_),
    .B1(_05110_));
 sg13g2_nor2_1 _22492_ (.A(net3208),
    .B(net4676),
    .Y(_05111_));
 sg13g2_a21oi_1 _22493_ (.A1(net5237),
    .A2(net4676),
    .Y(_01747_),
    .B1(_05111_));
 sg13g2_nor2_1 _22494_ (.A(net3257),
    .B(net4675),
    .Y(_05112_));
 sg13g2_a21oi_1 _22495_ (.A1(net5131),
    .A2(net4675),
    .Y(_01748_),
    .B1(_05112_));
 sg13g2_nor2_1 _22496_ (.A(net3137),
    .B(net4675),
    .Y(_05113_));
 sg13g2_a21oi_1 _22497_ (.A1(net5103),
    .A2(net4675),
    .Y(_01749_),
    .B1(_05113_));
 sg13g2_nor2_1 _22498_ (.A(net3043),
    .B(net4676),
    .Y(_05114_));
 sg13g2_a21oi_1 _22499_ (.A1(net5173),
    .A2(net4676),
    .Y(_01750_),
    .B1(_05114_));
 sg13g2_nor2_1 _22500_ (.A(net3102),
    .B(net4675),
    .Y(_05115_));
 sg13g2_a21oi_1 _22501_ (.A1(net5146),
    .A2(net4675),
    .Y(_01751_),
    .B1(_05115_));
 sg13g2_nor2_1 _22502_ (.A(net3700),
    .B(net4676),
    .Y(_05116_));
 sg13g2_a21oi_1 _22503_ (.A1(net5078),
    .A2(net4676),
    .Y(_01752_),
    .B1(_05116_));
 sg13g2_nor2_1 _22504_ (.A(net4287),
    .B(net4676),
    .Y(_05117_));
 sg13g2_a21oi_1 _22505_ (.A1(net5055),
    .A2(net4676),
    .Y(_01753_),
    .B1(_05117_));
 sg13g2_nand2_1 _22506_ (.Y(_05118_),
    .A(net3117),
    .B(net5312));
 sg13g2_nand3_1 _22507_ (.B(_08331_),
    .C(_08483_),
    .A(_08273_),
    .Y(_05119_));
 sg13g2_nand3_1 _22508_ (.B(_08358_),
    .C(_08518_),
    .A(_08172_),
    .Y(_05120_));
 sg13g2_nor2_1 _22509_ (.A(_05119_),
    .B(_05120_),
    .Y(_05121_));
 sg13g2_nand2_1 _22510_ (.Y(_05122_),
    .A(_08357_),
    .B(_08387_));
 sg13g2_nor4_1 _22511_ (.A(_08316_),
    .B(net5397),
    .C(net5402),
    .D(_05122_),
    .Y(_05123_));
 sg13g2_and3_1 _22512_ (.X(_05124_),
    .A(_04884_),
    .B(_05121_),
    .C(_05123_));
 sg13g2_nand3_1 _22513_ (.B(_05121_),
    .C(_05123_),
    .A(_04884_),
    .Y(_05125_));
 sg13g2_and2_1 _22514_ (.A(net5273),
    .B(_05124_),
    .X(_05126_));
 sg13g2_a21o_1 _22515_ (.A2(net5438),
    .A1(\atari2600.cpu.PC[7] ),
    .B1(_05126_),
    .X(_05127_));
 sg13g2_or2_2 _22516_ (.X(_05128_),
    .B(_08530_),
    .A(_08276_));
 sg13g2_a22oi_1 _22517_ (.Y(_05129_),
    .B1(_05128_),
    .B2(\atari2600.cpu.op[2] ),
    .A2(net5444),
    .A1(\atari2600.cpu.backwards ));
 sg13g2_nand2_1 _22518_ (.Y(_05130_),
    .A(_08585_),
    .B(_05129_));
 sg13g2_nand2_1 _22519_ (.Y(_05131_),
    .A(\atari2600.cpu.op[3] ),
    .B(_05128_));
 sg13g2_xor2_1 _22520_ (.B(net5323),
    .A(_05127_),
    .X(_05132_));
 sg13g2_and2_1 _22521_ (.A(\atari2600.cpu.shift_right ),
    .B(_05128_),
    .X(_05133_));
 sg13g2_o21ai_1 _22522_ (.B1(\atari2600.cpu.ALU.CO ),
    .Y(_05134_),
    .A1(net5444),
    .A2(_08525_));
 sg13g2_nor4_1 _22523_ (.A(_08316_),
    .B(_08381_),
    .C(_08498_),
    .D(_05120_),
    .Y(_05135_));
 sg13g2_a21oi_1 _22524_ (.A1(_08069_),
    .A2(\atari2600.cpu.inc ),
    .Y(_05136_),
    .B1(\atari2600.cpu.rotate ));
 sg13g2_a21oi_1 _22525_ (.A1(_08068_),
    .A2(\atari2600.cpu.rotate ),
    .Y(_05137_),
    .B1(_05136_));
 sg13g2_a21oi_1 _22526_ (.A1(_08056_),
    .A2(_08069_),
    .Y(_05138_),
    .B1(\atari2600.cpu.rotate ));
 sg13g2_nand2b_1 _22527_ (.Y(_05139_),
    .B(\atari2600.cpu.compare ),
    .A_N(\atari2600.cpu.rotate ));
 sg13g2_o21ai_1 _22528_ (.B1(_05139_),
    .Y(_05140_),
    .A1(_00095_),
    .A2(_05138_));
 sg13g2_a22oi_1 _22529_ (.Y(_05141_),
    .B1(_05140_),
    .B2(_08276_),
    .A2(_05137_),
    .A1(_08530_));
 sg13g2_nand3_1 _22530_ (.B(_05135_),
    .C(_05141_),
    .A(_05134_),
    .Y(_05142_));
 sg13g2_and2_1 _22531_ (.A(net5355),
    .B(_05142_),
    .X(_05143_));
 sg13g2_nor3_2 _22532_ (.A(net5480),
    .B(_08283_),
    .C(_05128_),
    .Y(_05144_));
 sg13g2_a21oi_2 _22533_ (.B1(_05144_),
    .Y(_05145_),
    .A2(_05128_),
    .A1(\atari2600.cpu.op[0] ));
 sg13g2_nand2_1 _22534_ (.Y(_05146_),
    .A(_05127_),
    .B(_05145_));
 sg13g2_a21oi_2 _22535_ (.B1(_05144_),
    .Y(_05147_),
    .A2(_05128_),
    .A1(\atari2600.cpu.op[1] ));
 sg13g2_a21o_2 _22536_ (.A2(_05128_),
    .A1(\atari2600.cpu.op[1] ),
    .B1(_05144_),
    .X(_05148_));
 sg13g2_nand3_1 _22537_ (.B(_08059_),
    .C(_05128_),
    .A(\atari2600.cpu.op[0] ),
    .Y(_05149_));
 sg13g2_nand2_1 _22538_ (.Y(_05150_),
    .A(_05146_),
    .B(_05149_));
 sg13g2_nor2_1 _22539_ (.A(_08505_),
    .B(_05119_),
    .Y(_05151_));
 sg13g2_nand2_1 _22540_ (.Y(_05152_),
    .A(_08056_),
    .B(_08276_));
 sg13g2_nor3_1 _22541_ (.A(_08256_),
    .B(_08498_),
    .C(_04890_),
    .Y(_05153_));
 sg13g2_nand3_1 _22542_ (.B(_05152_),
    .C(_05153_),
    .A(_05151_),
    .Y(_05154_));
 sg13g2_a22oi_1 _22543_ (.Y(_05155_),
    .B1(net5361),
    .B2(\atari2600.cpu.ADD[7] ),
    .A2(net5443),
    .A1(\atari2600.cpu.ABH[7] ));
 sg13g2_a22oi_1 _22544_ (.Y(_05156_),
    .B1(_05154_),
    .B2(_08599_),
    .A2(_04881_),
    .A1(net5273));
 sg13g2_and2_1 _22545_ (.A(_05155_),
    .B(_05156_),
    .X(_05157_));
 sg13g2_inv_1 _22546_ (.Y(_05158_),
    .A(_05157_));
 sg13g2_o21ai_1 _22547_ (.B1(_05127_),
    .Y(_05159_),
    .A1(_05147_),
    .A2(_05157_));
 sg13g2_a221oi_1 _22548_ (.B2(_05150_),
    .C1(net5355),
    .B1(_05159_),
    .A1(_05146_),
    .Y(_05160_),
    .A2(_05157_));
 sg13g2_a221oi_1 _22549_ (.B2(_05142_),
    .C1(_05160_),
    .B1(net5355),
    .A1(net5358),
    .Y(_05161_),
    .A2(_05132_));
 sg13g2_nor2_1 _22550_ (.A(net5323),
    .B(net5358),
    .Y(_05162_));
 sg13g2_or2_1 _22551_ (.X(_05163_),
    .B(net5358),
    .A(net5323));
 sg13g2_a21o_1 _22552_ (.A2(_05132_),
    .A1(net5358),
    .B1(_05162_),
    .X(_05164_));
 sg13g2_nand2_1 _22553_ (.Y(_05165_),
    .A(net5363),
    .B(_05164_));
 sg13g2_o21ai_1 _22554_ (.B1(_05118_),
    .Y(_01754_),
    .A1(_05161_),
    .A2(_05165_));
 sg13g2_nor3_2 _22555_ (.A(net7122),
    .B(_08133_),
    .C(net5386),
    .Y(_05166_));
 sg13g2_and2_2 _22556_ (.A(\atari2600.clk_counter[1] ),
    .B(_05166_),
    .X(_05167_));
 sg13g2_nand2_2 _22557_ (.Y(_05168_),
    .A(\atari2600.clk_counter[1] ),
    .B(_05166_));
 sg13g2_nor4_1 _22558_ (.A(\atari2600.pia.reset_timer[4] ),
    .B(\atari2600.pia.reset_timer[3] ),
    .C(\atari2600.pia.reset_timer[2] ),
    .D(\atari2600.pia.reset_timer[1] ),
    .Y(_05169_));
 sg13g2_nor4_2 _22559_ (.A(\atari2600.pia.reset_timer[0] ),
    .B(\atari2600.pia.reset_timer[7] ),
    .C(\atari2600.pia.reset_timer[6] ),
    .Y(_05170_),
    .D(\atari2600.pia.reset_timer[5] ));
 sg13g2_and2_1 _22560_ (.A(_05169_),
    .B(_05170_),
    .X(_05171_));
 sg13g2_nand2_1 _22561_ (.Y(_05172_),
    .A(_05169_),
    .B(_05170_));
 sg13g2_nor2_2 _22562_ (.A(\atari2600.pia.underflow ),
    .B(\atari2600.pia.interval[0] ),
    .Y(_05173_));
 sg13g2_nor3_2 _22563_ (.A(\atari2600.pia.interval[3] ),
    .B(\atari2600.pia.underflow ),
    .C(\atari2600.pia.interval[0] ),
    .Y(_05174_));
 sg13g2_nand2b_2 _22564_ (.Y(_05175_),
    .B(_05173_),
    .A_N(\atari2600.pia.interval[3] ));
 sg13g2_nor2_2 _22565_ (.A(\atari2600.pia.interval[6] ),
    .B(_05175_),
    .Y(_05176_));
 sg13g2_nand2b_1 _22566_ (.Y(_05177_),
    .B(\atari2600.pia.interval[6] ),
    .A_N(\atari2600.pia.underflow ));
 sg13g2_nor2_1 _22567_ (.A(_05174_),
    .B(_05177_),
    .Y(_05178_));
 sg13g2_nor2_1 _22568_ (.A(_05176_),
    .B(_05178_),
    .Y(_05179_));
 sg13g2_o21ai_1 _22569_ (.B1(_00078_),
    .Y(_05180_),
    .A1(_05176_),
    .A2(_05178_));
 sg13g2_nor2b_1 _22570_ (.A(\atari2600.pia.underflow ),
    .B_N(\atari2600.pia.interval[10] ),
    .Y(_05181_));
 sg13g2_and2_1 _22571_ (.A(_00079_),
    .B(_05181_),
    .X(_05182_));
 sg13g2_o21ai_1 _22572_ (.B1(_05175_),
    .Y(_05183_),
    .A1(\atari2600.pia.time_counter[5] ),
    .A2(\atari2600.pia.time_counter[4] ));
 sg13g2_nand3b_1 _22573_ (.B(\atari2600.pia.interval[0] ),
    .C(\atari2600.pia.interval[3] ),
    .Y(_05184_),
    .A_N(\atari2600.pia.underflow ));
 sg13g2_nand3_1 _22574_ (.B(_05175_),
    .C(_05184_),
    .A(\atari2600.pia.time_counter[3] ),
    .Y(_05185_));
 sg13g2_and2_1 _22575_ (.A(\atari2600.pia.time_counter[9] ),
    .B(\atari2600.pia.time_counter[8] ),
    .X(_05186_));
 sg13g2_nand2_1 _22576_ (.Y(_05187_),
    .A(\atari2600.pia.time_counter[5] ),
    .B(\atari2600.pia.time_counter[4] ));
 sg13g2_a21oi_1 _22577_ (.A1(_05175_),
    .A2(_05184_),
    .Y(_05188_),
    .B1(\atari2600.pia.time_counter[3] ));
 sg13g2_and4_1 _22578_ (.A(\atari2600.pia.time_counter[2] ),
    .B(\atari2600.pia.time_counter[1] ),
    .C(\atari2600.pia.time_counter[0] ),
    .D(_05173_),
    .X(_05189_));
 sg13g2_nor4_1 _22579_ (.A(\atari2600.pia.time_counter[2] ),
    .B(\atari2600.pia.time_counter[1] ),
    .C(\atari2600.pia.time_counter[0] ),
    .D(_05173_),
    .Y(_05190_));
 sg13g2_nand4_1 _22580_ (.B(_05174_),
    .C(_05177_),
    .A(\atari2600.pia.time_counter[7] ),
    .Y(_05191_),
    .D(_05182_));
 sg13g2_or3_1 _22581_ (.A(\atari2600.pia.time_counter[7] ),
    .B(_05176_),
    .C(_05182_),
    .X(_05192_));
 sg13g2_a22oi_1 _22582_ (.Y(_05193_),
    .B1(_05191_),
    .B2(_05192_),
    .A2(_05179_),
    .A1(_08050_));
 sg13g2_nor3_1 _22583_ (.A(\atari2600.pia.time_counter[9] ),
    .B(\atari2600.pia.time_counter[8] ),
    .C(_05176_),
    .Y(_05194_));
 sg13g2_a22oi_1 _22584_ (.Y(_05195_),
    .B1(_05194_),
    .B2(_05183_),
    .A2(_05186_),
    .A1(_05176_));
 sg13g2_o21ai_1 _22585_ (.B1(_05185_),
    .Y(_05196_),
    .A1(_05189_),
    .A2(_05190_));
 sg13g2_or4_1 _22586_ (.A(\atari2600.pia.time_counter[23] ),
    .B(\atari2600.pia.time_counter[22] ),
    .C(\atari2600.pia.time_counter[21] ),
    .D(\atari2600.pia.time_counter[20] ),
    .X(_05197_));
 sg13g2_nor3_1 _22587_ (.A(\atari2600.pia.time_counter[14] ),
    .B(\atari2600.pia.time_counter[13] ),
    .C(_05197_),
    .Y(_05198_));
 sg13g2_or4_1 _22588_ (.A(\atari2600.pia.time_counter[19] ),
    .B(\atari2600.pia.time_counter[18] ),
    .C(\atari2600.pia.time_counter[17] ),
    .D(\atari2600.pia.time_counter[16] ),
    .X(_05199_));
 sg13g2_nor4_1 _22589_ (.A(\atari2600.pia.time_counter[15] ),
    .B(\atari2600.pia.time_counter[12] ),
    .C(\atari2600.pia.time_counter[11] ),
    .D(_05199_),
    .Y(_05200_));
 sg13g2_o21ai_1 _22590_ (.B1(_05200_),
    .Y(_05201_),
    .A1(_00079_),
    .A2(_05181_));
 sg13g2_a21oi_1 _22591_ (.A1(_05174_),
    .A2(_05187_),
    .Y(_05202_),
    .B1(_05201_));
 sg13g2_nand4_1 _22592_ (.B(_05193_),
    .C(_05198_),
    .A(_05180_),
    .Y(_05203_),
    .D(_05202_));
 sg13g2_nor4_2 _22593_ (.A(_05188_),
    .B(_05195_),
    .C(_05196_),
    .Y(_05204_),
    .D(_05203_));
 sg13g2_nand2b_1 _22594_ (.Y(_05205_),
    .B(_05171_),
    .A_N(_05204_));
 sg13g2_and2_1 _22595_ (.A(_05167_),
    .B(_05205_),
    .X(_05206_));
 sg13g2_nor2_1 _22596_ (.A(net5980),
    .B(_05206_),
    .Y(_05207_));
 sg13g2_nand2b_2 _22597_ (.Y(_05208_),
    .B(net6001),
    .A_N(_05206_));
 sg13g2_nand2_1 _22598_ (.Y(_05209_),
    .A(net7026),
    .B(net5141));
 sg13g2_mux2_1 _22599_ (.A0(net6538),
    .A1(net7026),
    .S(net5322),
    .X(_05210_));
 sg13g2_nand2_2 _22600_ (.Y(_05211_),
    .A(net6000),
    .B(_05206_));
 sg13g2_o21ai_1 _22601_ (.B1(_05209_),
    .Y(_01755_),
    .A1(_05210_),
    .A2(_05211_));
 sg13g2_nand2_1 _22602_ (.Y(_05212_),
    .A(net7087),
    .B(net5141));
 sg13g2_mux2_1 _22603_ (.A0(\atari2600.pia.reset_timer[1] ),
    .A1(\atari2600.pia.diag[1] ),
    .S(net5322),
    .X(_05213_));
 sg13g2_or2_1 _22604_ (.X(_05214_),
    .B(_05213_),
    .A(_05210_));
 sg13g2_xor2_1 _22605_ (.B(_05213_),
    .A(_05210_),
    .X(_05215_));
 sg13g2_o21ai_1 _22606_ (.B1(_05212_),
    .Y(_01756_),
    .A1(_05211_),
    .A2(_05215_));
 sg13g2_nand2_1 _22607_ (.Y(_05216_),
    .A(net7115),
    .B(net5141));
 sg13g2_mux2_1 _22608_ (.A0(\atari2600.pia.reset_timer[2] ),
    .A1(\atari2600.pia.diag[2] ),
    .S(net5322),
    .X(_05217_));
 sg13g2_xor2_1 _22609_ (.B(_05217_),
    .A(_05214_),
    .X(_05218_));
 sg13g2_o21ai_1 _22610_ (.B1(_05216_),
    .Y(_01757_),
    .A1(_05211_),
    .A2(_05218_));
 sg13g2_nand2_1 _22611_ (.Y(_05219_),
    .A(net7074),
    .B(net5141));
 sg13g2_mux2_1 _22612_ (.A0(\atari2600.pia.reset_timer[3] ),
    .A1(\atari2600.pia.diag[3] ),
    .S(net5322),
    .X(_05220_));
 sg13g2_nor3_2 _22613_ (.A(_05214_),
    .B(_05217_),
    .C(_05220_),
    .Y(_05221_));
 sg13g2_o21ai_1 _22614_ (.B1(_05220_),
    .Y(_05222_),
    .A1(_05214_),
    .A2(_05217_));
 sg13g2_nor2b_1 _22615_ (.A(_05221_),
    .B_N(_05222_),
    .Y(_05223_));
 sg13g2_o21ai_1 _22616_ (.B1(_05219_),
    .Y(_01758_),
    .A1(_05211_),
    .A2(_05223_));
 sg13g2_nand2_1 _22617_ (.Y(_05224_),
    .A(net3829),
    .B(net5141));
 sg13g2_nor2_1 _22618_ (.A(\atari2600.pia.reset_timer[4] ),
    .B(net5322),
    .Y(_05225_));
 sg13g2_nand2b_1 _22619_ (.Y(_05226_),
    .B(_05204_),
    .A_N(\atari2600.pia.diag[4] ));
 sg13g2_nor2b_1 _22620_ (.A(_05225_),
    .B_N(_05226_),
    .Y(_05227_));
 sg13g2_nand2b_1 _22621_ (.Y(_05228_),
    .B(_05221_),
    .A_N(_05227_));
 sg13g2_xnor2_1 _22622_ (.Y(_05229_),
    .A(_05221_),
    .B(_05227_));
 sg13g2_o21ai_1 _22623_ (.B1(_05224_),
    .Y(_01759_),
    .A1(_05211_),
    .A2(_05229_));
 sg13g2_nand2_1 _22624_ (.Y(_05230_),
    .A(net7075),
    .B(_05207_));
 sg13g2_mux2_1 _22625_ (.A0(\atari2600.pia.reset_timer[5] ),
    .A1(\atari2600.pia.diag[5] ),
    .S(net5322),
    .X(_05231_));
 sg13g2_nor2_1 _22626_ (.A(_05228_),
    .B(_05231_),
    .Y(_05232_));
 sg13g2_xor2_1 _22627_ (.B(_05231_),
    .A(_05228_),
    .X(_05233_));
 sg13g2_o21ai_1 _22628_ (.B1(_05230_),
    .Y(_01760_),
    .A1(_05211_),
    .A2(_05233_));
 sg13g2_nand2_1 _22629_ (.Y(_05234_),
    .A(net7060),
    .B(net5141));
 sg13g2_mux2_1 _22630_ (.A0(\atari2600.pia.reset_timer[6] ),
    .A1(\atari2600.pia.diag[6] ),
    .S(net5322),
    .X(_05235_));
 sg13g2_nor3_1 _22631_ (.A(_05228_),
    .B(_05231_),
    .C(_05235_),
    .Y(_05236_));
 sg13g2_xnor2_1 _22632_ (.Y(_05237_),
    .A(_05232_),
    .B(_05235_));
 sg13g2_o21ai_1 _22633_ (.B1(_05234_),
    .Y(_01761_),
    .A1(_05211_),
    .A2(_05237_));
 sg13g2_nand2_1 _22634_ (.Y(_05238_),
    .A(net6951),
    .B(net5141));
 sg13g2_mux2_1 _22635_ (.A0(\atari2600.pia.reset_timer[7] ),
    .A1(\atari2600.pia.diag[7] ),
    .S(net5322),
    .X(_05239_));
 sg13g2_xnor2_1 _22636_ (.Y(_05240_),
    .A(_05236_),
    .B(_05239_));
 sg13g2_o21ai_1 _22637_ (.B1(_05238_),
    .Y(_01762_),
    .A1(_05211_),
    .A2(_05240_));
 sg13g2_nand2_1 _22638_ (.Y(_05241_),
    .A(_05167_),
    .B(_05172_));
 sg13g2_a21oi_1 _22639_ (.A1(_05167_),
    .A2(_05172_),
    .Y(_05242_),
    .B1(net5980));
 sg13g2_nand2_2 _22640_ (.Y(_05243_),
    .A(net6001),
    .B(_05241_));
 sg13g2_nor3_1 _22641_ (.A(\atari2600.pia.diag[2] ),
    .B(\atari2600.pia.diag[1] ),
    .C(net7377),
    .Y(_05244_));
 sg13g2_nor4_1 _22642_ (.A(\atari2600.pia.diag[7] ),
    .B(\atari2600.pia.diag[6] ),
    .C(\atari2600.pia.diag[5] ),
    .D(\atari2600.pia.diag[3] ),
    .Y(_05245_));
 sg13g2_nand3_1 _22643_ (.B(_05244_),
    .C(_05245_),
    .A(net6000),
    .Y(_05246_));
 sg13g2_nor3_1 _22644_ (.A(_05168_),
    .B(_05226_),
    .C(net7378),
    .Y(_05247_));
 sg13g2_a21o_1 _22645_ (.A2(net5209),
    .A1(net3644),
    .B1(_05247_),
    .X(_01763_));
 sg13g2_and2_1 _22646_ (.A(_10403_),
    .B(_03006_),
    .X(_05248_));
 sg13g2_nand2_2 _22647_ (.Y(_05249_),
    .A(net5344),
    .B(net4762));
 sg13g2_nor2_2 _22648_ (.A(_08589_),
    .B(net4732),
    .Y(_05250_));
 sg13g2_and3_2 _22649_ (.X(_05251_),
    .A(_03005_),
    .B(_04813_),
    .C(_05250_));
 sg13g2_nand3_1 _22650_ (.B(_04813_),
    .C(_05250_),
    .A(_03005_),
    .Y(_05252_));
 sg13g2_nand3_1 _22651_ (.B(net5352),
    .C(net4762),
    .A(net6002),
    .Y(_05253_));
 sg13g2_inv_1 _22652_ (.Y(_05254_),
    .A(_05253_));
 sg13g2_nor2_1 _22653_ (.A(net4019),
    .B(_05251_),
    .Y(_05255_));
 sg13g2_nor2_1 _22654_ (.A(_08677_),
    .B(_04814_),
    .Y(_05256_));
 sg13g2_nor2_2 _22655_ (.A(_08565_),
    .B(net4935),
    .Y(_05257_));
 sg13g2_nand2_2 _22656_ (.Y(_05258_),
    .A(net4911),
    .B(_08746_));
 sg13g2_nor2_2 _22657_ (.A(_03166_),
    .B(_04814_),
    .Y(_05259_));
 sg13g2_nor2_2 _22658_ (.A(_08735_),
    .B(net4928),
    .Y(_05260_));
 sg13g2_nand2_2 _22659_ (.Y(_05261_),
    .A(net4826),
    .B(_08746_));
 sg13g2_nor2_2 _22660_ (.A(_03164_),
    .B(_05261_),
    .Y(_05262_));
 sg13g2_nand2_2 _22661_ (.Y(_05263_),
    .A(_03163_),
    .B(_05260_));
 sg13g2_and2_1 _22662_ (.A(\atari2600.input_joystick_0[0] ),
    .B(_05262_),
    .X(_05264_));
 sg13g2_a221oi_1 _22663_ (.B2(net3941),
    .C1(_05264_),
    .B1(_05259_),
    .A1(\atari2600.pia.diag[0] ),
    .Y(_05265_),
    .A2(net4674));
 sg13g2_a21oi_1 _22664_ (.A1(net7101),
    .A2(_10251_),
    .Y(_05266_),
    .B1(_05252_));
 sg13g2_a21oi_1 _22665_ (.A1(_05265_),
    .A2(_05266_),
    .Y(_01764_),
    .B1(_05255_));
 sg13g2_nor2_1 _22666_ (.A(net3987),
    .B(_05251_),
    .Y(_05267_));
 sg13g2_and2_1 _22667_ (.A(net2995),
    .B(_05262_),
    .X(_05268_));
 sg13g2_a221oi_1 _22668_ (.B2(net3920),
    .C1(_05268_),
    .B1(_05259_),
    .A1(\atari2600.pia.diag[1] ),
    .Y(_05269_),
    .A2(net4674));
 sg13g2_a21oi_1 _22669_ (.A1(net7023),
    .A2(_10251_),
    .Y(_05270_),
    .B1(_05252_));
 sg13g2_a21oi_1 _22670_ (.A1(_05269_),
    .A2(_05270_),
    .Y(_01765_),
    .B1(_05267_));
 sg13g2_nor2_1 _22671_ (.A(net3313),
    .B(_05251_),
    .Y(_05271_));
 sg13g2_nor3_2 _22672_ (.A(net5029),
    .B(net4948),
    .C(_04814_),
    .Y(_05272_));
 sg13g2_a21o_1 _22673_ (.A2(_05272_),
    .A1(net3244),
    .B1(_05262_),
    .X(_05273_));
 sg13g2_a221oi_1 _22674_ (.B2(\atari2600.pia.swa_dir[2] ),
    .C1(_05273_),
    .B1(_05259_),
    .A1(\atari2600.pia.diag[2] ),
    .Y(_05274_),
    .A2(net4674));
 sg13g2_a21oi_1 _22675_ (.A1(\atari2600.input_joystick_0[5] ),
    .A2(_10251_),
    .Y(_05275_),
    .B1(_05252_));
 sg13g2_a21oi_1 _22676_ (.A1(_05274_),
    .A2(_05275_),
    .Y(_01766_),
    .B1(_05271_));
 sg13g2_nor2_1 _22677_ (.A(net6223),
    .B(_05251_),
    .Y(_05276_));
 sg13g2_and2_1 _22678_ (.A(\atari2600.input_switches[2] ),
    .B(_05262_),
    .X(_05277_));
 sg13g2_a221oi_1 _22679_ (.B2(net3351),
    .C1(_05277_),
    .B1(_05259_),
    .A1(\atari2600.pia.diag[3] ),
    .Y(_05278_),
    .A2(net4674));
 sg13g2_a21oi_1 _22680_ (.A1(\atari2600.input_joystick_0[6] ),
    .A2(_10251_),
    .Y(_05279_),
    .B1(_05252_));
 sg13g2_a21oi_1 _22681_ (.A1(_05278_),
    .A2(_05279_),
    .Y(_01767_),
    .B1(_05276_));
 sg13g2_nand2_1 _22682_ (.Y(_05280_),
    .A(net3086),
    .B(_05272_));
 sg13g2_a22oi_1 _22683_ (.Y(_05281_),
    .B1(_05259_),
    .B2(net3916),
    .A2(_05256_),
    .A1(\atari2600.pia.diag[4] ));
 sg13g2_nand4_1 _22684_ (.B(_05266_),
    .C(_05280_),
    .A(_05263_),
    .Y(_05282_),
    .D(_05281_));
 sg13g2_o21ai_1 _22685_ (.B1(_05282_),
    .Y(_05283_),
    .A1(net6599),
    .A2(_05251_));
 sg13g2_inv_1 _22686_ (.Y(_01768_),
    .A(_05283_));
 sg13g2_a21oi_1 _22687_ (.A1(net3044),
    .A2(_05259_),
    .Y(_05284_),
    .B1(_05262_));
 sg13g2_a22oi_1 _22688_ (.Y(_05285_),
    .B1(_05272_),
    .B2(net3845),
    .A2(net4674),
    .A1(\atari2600.pia.diag[5] ));
 sg13g2_nand3_1 _22689_ (.B(_05284_),
    .C(_05285_),
    .A(_05270_),
    .Y(_05286_));
 sg13g2_o21ai_1 _22690_ (.B1(_05286_),
    .Y(_05287_),
    .A1(net4532),
    .A2(_05251_));
 sg13g2_inv_1 _22691_ (.Y(_01769_),
    .A(_05287_));
 sg13g2_nor2_1 _22692_ (.A(net3065),
    .B(_05251_),
    .Y(_05288_));
 sg13g2_nand3_1 _22693_ (.B(_08583_),
    .C(_03163_),
    .A(\atari2600.pia.instat[0] ),
    .Y(_05289_));
 sg13g2_o21ai_1 _22694_ (.B1(_05289_),
    .Y(_05290_),
    .A1(\atari2600.input_switches[1] ),
    .A2(_05263_));
 sg13g2_a221oi_1 _22695_ (.B2(\atari2600.pia.swa_dir[6] ),
    .C1(_05290_),
    .B1(_05259_),
    .A1(\atari2600.pia.diag[6] ),
    .Y(_05291_),
    .A2(net4674));
 sg13g2_a21oi_1 _22696_ (.A1(_05275_),
    .A2(_05291_),
    .Y(_01770_),
    .B1(_05288_));
 sg13g2_nor2_1 _22697_ (.A(net3409),
    .B(_05251_),
    .Y(_05292_));
 sg13g2_nand3_1 _22698_ (.B(_08583_),
    .C(_03163_),
    .A(\atari2600.pia.instat[1] ),
    .Y(_05293_));
 sg13g2_o21ai_1 _22699_ (.B1(_05293_),
    .Y(_05294_),
    .A1(\atari2600.input_switches[0] ),
    .A2(_05263_));
 sg13g2_a221oi_1 _22700_ (.B2(\atari2600.pia.swa_dir[7] ),
    .C1(_05294_),
    .B1(_05259_),
    .A1(\atari2600.pia.diag[7] ),
    .Y(_05295_),
    .A2(net4674));
 sg13g2_a21oi_1 _22701_ (.A1(_05279_),
    .A2(_05295_),
    .Y(_01771_),
    .B1(_05292_));
 sg13g2_nor2_2 _22702_ (.A(_05168_),
    .B(_05205_),
    .Y(_05296_));
 sg13g2_nor2_1 _22703_ (.A(net7117),
    .B(_05296_),
    .Y(_05297_));
 sg13g2_and2_1 _22704_ (.A(net7117),
    .B(_05167_),
    .X(_05298_));
 sg13g2_nor3_1 _22705_ (.A(net5980),
    .B(_05297_),
    .C(_05298_),
    .Y(_01772_));
 sg13g2_xnor2_1 _22706_ (.Y(_05299_),
    .A(net7208),
    .B(_05298_));
 sg13g2_nor2_1 _22707_ (.A(_05243_),
    .B(_05299_),
    .Y(_01773_));
 sg13g2_a21oi_1 _22708_ (.A1(\atari2600.pia.time_counter[1] ),
    .A2(_05298_),
    .Y(_05300_),
    .B1(net6989));
 sg13g2_and4_1 _22709_ (.A(net6989),
    .B(\atari2600.pia.time_counter[1] ),
    .C(\atari2600.pia.time_counter[0] ),
    .D(_05167_),
    .X(_05301_));
 sg13g2_nor3_1 _22710_ (.A(_05243_),
    .B(net6990),
    .C(_05301_),
    .Y(_01774_));
 sg13g2_nor2_1 _22711_ (.A(net7071),
    .B(_05301_),
    .Y(_05302_));
 sg13g2_nand4_1 _22712_ (.B(\atari2600.pia.time_counter[2] ),
    .C(\atari2600.pia.time_counter[1] ),
    .A(net7071),
    .Y(_05303_),
    .D(\atari2600.pia.time_counter[0] ));
 sg13g2_nor2_2 _22713_ (.A(_05168_),
    .B(_05303_),
    .Y(_05304_));
 sg13g2_nor3_1 _22714_ (.A(_05208_),
    .B(net7072),
    .C(_05304_),
    .Y(_01775_));
 sg13g2_a21oi_1 _22715_ (.A1(net7172),
    .A2(_05304_),
    .Y(_05305_),
    .B1(_05243_));
 sg13g2_o21ai_1 _22716_ (.B1(_05305_),
    .Y(_05306_),
    .A1(net7172),
    .A2(_05304_));
 sg13g2_inv_1 _22717_ (.Y(_01776_),
    .A(net7173));
 sg13g2_a21oi_1 _22718_ (.A1(\atari2600.pia.time_counter[4] ),
    .A2(_05304_),
    .Y(_05307_),
    .B1(net3168));
 sg13g2_nor2_2 _22719_ (.A(_05187_),
    .B(_05303_),
    .Y(_05308_));
 sg13g2_and2_1 _22720_ (.A(_05167_),
    .B(_05308_),
    .X(_05309_));
 sg13g2_nor3_1 _22721_ (.A(_05243_),
    .B(net3169),
    .C(_05309_),
    .Y(_01777_));
 sg13g2_xnor2_1 _22722_ (.Y(_05310_),
    .A(_00078_),
    .B(_05308_));
 sg13g2_a22oi_1 _22723_ (.Y(_05311_),
    .B1(_05296_),
    .B2(_05310_),
    .A2(_05168_),
    .A1(net3883));
 sg13g2_nor2_1 _22724_ (.A(net5980),
    .B(net3884),
    .Y(_01778_));
 sg13g2_and3_1 _22725_ (.X(_05312_),
    .A(net3883),
    .B(_05167_),
    .C(_05308_));
 sg13g2_nor2_1 _22726_ (.A(net7159),
    .B(_05312_),
    .Y(_05313_));
 sg13g2_and2_1 _22727_ (.A(net7159),
    .B(_05312_),
    .X(_05314_));
 sg13g2_nor3_1 _22728_ (.A(_05208_),
    .B(_05313_),
    .C(_05314_),
    .Y(_01779_));
 sg13g2_o21ai_1 _22729_ (.B1(net5141),
    .Y(_05315_),
    .A1(net6150),
    .A2(_05314_));
 sg13g2_a21oi_1 _22730_ (.A1(net6150),
    .A2(_05314_),
    .Y(_01780_),
    .B1(_05315_));
 sg13g2_a21oi_1 _22731_ (.A1(\atari2600.pia.time_counter[8] ),
    .A2(_05314_),
    .Y(_05316_),
    .B1(net3870));
 sg13g2_nand4_1 _22732_ (.B(net3883),
    .C(_05186_),
    .A(\atari2600.pia.time_counter[7] ),
    .Y(_05317_),
    .D(_05308_));
 sg13g2_nor2_1 _22733_ (.A(_05168_),
    .B(_05317_),
    .Y(_05318_));
 sg13g2_and2_1 _22734_ (.A(\atari2600.pia.time_counter[7] ),
    .B(_05186_),
    .X(_05319_));
 sg13g2_nor3_1 _22735_ (.A(_05208_),
    .B(net3871),
    .C(_05318_),
    .Y(_01781_));
 sg13g2_xor2_1 _22736_ (.B(_05317_),
    .A(_00079_),
    .X(_05320_));
 sg13g2_a22oi_1 _22737_ (.Y(_05321_),
    .B1(_05296_),
    .B2(_05320_),
    .A2(_05168_),
    .A1(net6960));
 sg13g2_nor2_1 _22738_ (.A(net5980),
    .B(net6961),
    .Y(_01782_));
 sg13g2_a21oi_1 _22739_ (.A1(\atari2600.pia.time_counter[10] ),
    .A2(_05318_),
    .Y(_05322_),
    .B1(net4022));
 sg13g2_and4_1 _22740_ (.A(net4022),
    .B(net6960),
    .C(_05312_),
    .D(_05319_),
    .X(_05323_));
 sg13g2_nor3_1 _22741_ (.A(_05208_),
    .B(net4023),
    .C(_05323_),
    .Y(_01783_));
 sg13g2_nor2_1 _22742_ (.A(net6970),
    .B(_05323_),
    .Y(_05324_));
 sg13g2_and4_1 _22743_ (.A(net6970),
    .B(net4022),
    .C(net6960),
    .D(_05318_),
    .X(_05325_));
 sg13g2_nand2b_1 _22744_ (.Y(_05326_),
    .B(net5208),
    .A_N(_05325_));
 sg13g2_nor2_1 _22745_ (.A(_05324_),
    .B(_05326_),
    .Y(_01784_));
 sg13g2_nand2b_1 _22746_ (.Y(_05327_),
    .B(net6001),
    .A_N(net6993));
 sg13g2_a21oi_1 _22747_ (.A1(_05171_),
    .A2(_05325_),
    .Y(_05328_),
    .B1(net6993));
 sg13g2_a21oi_1 _22748_ (.A1(_05326_),
    .A2(_05327_),
    .Y(_01785_),
    .B1(net6994));
 sg13g2_a21oi_1 _22749_ (.A1(\atari2600.pia.time_counter[13] ),
    .A2(_05325_),
    .Y(_05329_),
    .B1(net3794));
 sg13g2_and4_1 _22750_ (.A(net3794),
    .B(net6993),
    .C(net6970),
    .D(_05323_),
    .X(_05330_));
 sg13g2_and2_1 _22751_ (.A(\atari2600.pia.time_counter[14] ),
    .B(\atari2600.pia.time_counter[13] ),
    .X(_05331_));
 sg13g2_nor3_1 _22752_ (.A(_05243_),
    .B(net3795),
    .C(_05330_),
    .Y(_01786_));
 sg13g2_and2_1 _22753_ (.A(net7109),
    .B(_05330_),
    .X(_05332_));
 sg13g2_o21ai_1 _22754_ (.B1(net5208),
    .Y(_05333_),
    .A1(net7109),
    .A2(_05330_));
 sg13g2_nor2_1 _22755_ (.A(_05332_),
    .B(_05333_),
    .Y(_01787_));
 sg13g2_nor2_1 _22756_ (.A(net7062),
    .B(_05332_),
    .Y(_05334_));
 sg13g2_and4_1 _22757_ (.A(\atari2600.pia.time_counter[16] ),
    .B(\atari2600.pia.time_counter[15] ),
    .C(_05325_),
    .D(_05331_),
    .X(_05335_));
 sg13g2_nand2b_1 _22758_ (.Y(_05336_),
    .B(net5208),
    .A_N(_05335_));
 sg13g2_nor2_1 _22759_ (.A(net7063),
    .B(_05336_),
    .Y(_01788_));
 sg13g2_nand2b_1 _22760_ (.Y(_05337_),
    .B(net6000),
    .A_N(net4180));
 sg13g2_a21oi_1 _22761_ (.A1(_05171_),
    .A2(_05335_),
    .Y(_05338_),
    .B1(net4180));
 sg13g2_a21oi_1 _22762_ (.A1(_05336_),
    .A2(_05337_),
    .Y(_01789_),
    .B1(net4181));
 sg13g2_a21oi_1 _22763_ (.A1(\atari2600.pia.time_counter[17] ),
    .A2(_05335_),
    .Y(_05339_),
    .B1(net3414));
 sg13g2_and4_2 _22764_ (.A(net3414),
    .B(net4180),
    .C(\atari2600.pia.time_counter[16] ),
    .D(_05332_),
    .X(_05340_));
 sg13g2_nor3_1 _22765_ (.A(_05243_),
    .B(net3415),
    .C(_05340_),
    .Y(_01790_));
 sg13g2_o21ai_1 _22766_ (.B1(net5208),
    .Y(_05341_),
    .A1(net6534),
    .A2(_05340_));
 sg13g2_a21oi_1 _22767_ (.A1(net6534),
    .A2(_05340_),
    .Y(_01791_),
    .B1(_05341_));
 sg13g2_a21oi_1 _22768_ (.A1(\atari2600.pia.time_counter[19] ),
    .A2(_05340_),
    .Y(_05342_),
    .B1(net3580));
 sg13g2_and3_1 _22769_ (.X(_05343_),
    .A(net3580),
    .B(net6534),
    .C(_05340_));
 sg13g2_nor3_1 _22770_ (.A(_05243_),
    .B(net3581),
    .C(_05343_),
    .Y(_01792_));
 sg13g2_and2_1 _22771_ (.A(net7095),
    .B(_05343_),
    .X(_05344_));
 sg13g2_o21ai_1 _22772_ (.B1(net5208),
    .Y(_05345_),
    .A1(net7095),
    .A2(_05343_));
 sg13g2_nor2_1 _22773_ (.A(_05344_),
    .B(_05345_),
    .Y(_01793_));
 sg13g2_nand2_1 _22774_ (.Y(_05346_),
    .A(net7121),
    .B(_05344_));
 sg13g2_o21ai_1 _22775_ (.B1(net5208),
    .Y(_05347_),
    .A1(net7121),
    .A2(_05344_));
 sg13g2_nor2b_1 _22776_ (.A(_05347_),
    .B_N(_05346_),
    .Y(_01794_));
 sg13g2_and3_1 _22777_ (.X(_05348_),
    .A(net7237),
    .B(_05241_),
    .C(_05346_));
 sg13g2_nor3_1 _22778_ (.A(net7237),
    .B(_05172_),
    .C(_05346_),
    .Y(_05349_));
 sg13g2_o21ai_1 _22779_ (.B1(net6000),
    .Y(_05350_),
    .A1(_05348_),
    .A2(_05349_));
 sg13g2_inv_1 _22780_ (.Y(_01795_),
    .A(_05350_));
 sg13g2_nand3_1 _22781_ (.B(net5344),
    .C(net4762),
    .A(_08589_),
    .Y(_05351_));
 sg13g2_and4_1 _22782_ (.A(net5030),
    .B(_08589_),
    .C(net4763),
    .D(_05254_),
    .X(_05352_));
 sg13g2_nand4_1 _22783_ (.B(_08589_),
    .C(net4763),
    .A(net5030),
    .Y(_05353_),
    .D(_05254_));
 sg13g2_nand3_1 _22784_ (.B(net6001),
    .C(net4578),
    .A(net7331),
    .Y(_05354_));
 sg13g2_a21oi_1 _22785_ (.A1(_05250_),
    .A2(net4674),
    .Y(_05355_),
    .B1(_05354_));
 sg13g2_or2_1 _22786_ (.X(_01796_),
    .B(_05355_),
    .A(_05247_));
 sg13g2_nand2_1 _22787_ (.Y(_05356_),
    .A(net6538),
    .B(net5976));
 sg13g2_a21oi_1 _22788_ (.A1(net6538),
    .A2(_05249_),
    .Y(_05357_),
    .B1(net4581));
 sg13g2_o21ai_1 _22789_ (.B1(net5207),
    .Y(_05358_),
    .A1(net5254),
    .A2(net4579));
 sg13g2_o21ai_1 _22790_ (.B1(_05356_),
    .Y(_01797_),
    .A1(_05357_),
    .A2(_05358_));
 sg13g2_nand2_1 _22791_ (.Y(_05359_),
    .A(net5976),
    .B(net4179));
 sg13g2_nand2_2 _22792_ (.Y(_05360_),
    .A(net6008),
    .B(net5230));
 sg13g2_a21oi_1 _22793_ (.A1(net4179),
    .A2(net4732),
    .Y(_05361_),
    .B1(net4581));
 sg13g2_o21ai_1 _22794_ (.B1(net5207),
    .Y(_05362_),
    .A1(net5223),
    .A2(net4578));
 sg13g2_o21ai_1 _22795_ (.B1(_05359_),
    .Y(_01798_),
    .A1(_05361_),
    .A2(_05362_));
 sg13g2_nand2_1 _22796_ (.Y(_05363_),
    .A(net5977),
    .B(net7096));
 sg13g2_a21oi_1 _22797_ (.A1(net7096),
    .A2(net4732),
    .Y(_05364_),
    .B1(net4581));
 sg13g2_o21ai_1 _22798_ (.B1(net5207),
    .Y(_05365_),
    .A1(net5119),
    .A2(net4578));
 sg13g2_o21ai_1 _22799_ (.B1(_05363_),
    .Y(_01799_),
    .A1(_05364_),
    .A2(_05365_));
 sg13g2_nand2_1 _22800_ (.Y(_05366_),
    .A(net5976),
    .B(net6209));
 sg13g2_a21oi_1 _22801_ (.A1(net6209),
    .A2(net4732),
    .Y(_05367_),
    .B1(net4581));
 sg13g2_o21ai_1 _22802_ (.B1(net5207),
    .Y(_05368_),
    .A1(net5093),
    .A2(net4578));
 sg13g2_o21ai_1 _22803_ (.B1(_05366_),
    .Y(_01800_),
    .A1(_05367_),
    .A2(_05368_));
 sg13g2_nand2_1 _22804_ (.Y(_05369_),
    .A(net5976),
    .B(net6345));
 sg13g2_a21oi_1 _22805_ (.A1(net6345),
    .A2(net4732),
    .Y(_05370_),
    .B1(net4580));
 sg13g2_o21ai_1 _22806_ (.B1(net5207),
    .Y(_05371_),
    .A1(net5189),
    .A2(net4579));
 sg13g2_o21ai_1 _22807_ (.B1(_05369_),
    .Y(_01801_),
    .A1(_05370_),
    .A2(_05371_));
 sg13g2_nand2_1 _22808_ (.Y(_05372_),
    .A(net5981),
    .B(net6700));
 sg13g2_a21oi_1 _22809_ (.A1(net6700),
    .A2(net4732),
    .Y(_05373_),
    .B1(net4580));
 sg13g2_o21ai_1 _22810_ (.B1(net5207),
    .Y(_05374_),
    .A1(net5164),
    .A2(net4579));
 sg13g2_o21ai_1 _22811_ (.B1(_05372_),
    .Y(_01802_),
    .A1(_05373_),
    .A2(_05374_));
 sg13g2_nand2_1 _22812_ (.Y(_05375_),
    .A(net5976),
    .B(net6418));
 sg13g2_a21oi_1 _22813_ (.A1(net6418),
    .A2(net4732),
    .Y(_05376_),
    .B1(net4580));
 sg13g2_o21ai_1 _22814_ (.B1(net5207),
    .Y(_05377_),
    .A1(net5070),
    .A2(net4579));
 sg13g2_o21ai_1 _22815_ (.B1(_05375_),
    .Y(_01803_),
    .A1(_05376_),
    .A2(_05377_));
 sg13g2_nand2_1 _22816_ (.Y(_05378_),
    .A(net5980),
    .B(net7034));
 sg13g2_a21oi_1 _22817_ (.A1(net7034),
    .A2(net4732),
    .Y(_05379_),
    .B1(net4580));
 sg13g2_o21ai_1 _22818_ (.B1(net5207),
    .Y(_05380_),
    .A1(net5047),
    .A2(net4579));
 sg13g2_o21ai_1 _22819_ (.B1(_05378_),
    .Y(_01804_),
    .A1(_05379_),
    .A2(_05380_));
 sg13g2_nor3_1 _22820_ (.A(_03166_),
    .B(_04814_),
    .C(_05351_),
    .Y(_05381_));
 sg13g2_nor2_1 _22821_ (.A(net3941),
    .B(net4672),
    .Y(_05382_));
 sg13g2_a21oi_1 _22822_ (.A1(net5262),
    .A2(net4672),
    .Y(_01805_),
    .B1(_05382_));
 sg13g2_nor2_1 _22823_ (.A(net3920),
    .B(net4672),
    .Y(_05383_));
 sg13g2_a21oi_1 _22824_ (.A1(net5235),
    .A2(net4672),
    .Y(_01806_),
    .B1(_05383_));
 sg13g2_nor2_1 _22825_ (.A(net3602),
    .B(net4673),
    .Y(_05384_));
 sg13g2_a21oi_1 _22826_ (.A1(net5133),
    .A2(net4673),
    .Y(_01807_),
    .B1(_05384_));
 sg13g2_nor2_1 _22827_ (.A(net3351),
    .B(net4672),
    .Y(_05385_));
 sg13g2_a21oi_1 _22828_ (.A1(net5104),
    .A2(net4672),
    .Y(_01808_),
    .B1(_05385_));
 sg13g2_nor2_1 _22829_ (.A(net3916),
    .B(net4673),
    .Y(_05386_));
 sg13g2_a21oi_1 _22830_ (.A1(net5178),
    .A2(net4673),
    .Y(_01809_),
    .B1(_05386_));
 sg13g2_nor2_1 _22831_ (.A(net3044),
    .B(net4672),
    .Y(_05387_));
 sg13g2_a21oi_1 _22832_ (.A1(net5147),
    .A2(net4672),
    .Y(_01810_),
    .B1(_05387_));
 sg13g2_nor2_1 _22833_ (.A(net3701),
    .B(net4673),
    .Y(_05388_));
 sg13g2_a21oi_1 _22834_ (.A1(net5079),
    .A2(net4673),
    .Y(_01811_),
    .B1(_05388_));
 sg13g2_nor2_1 _22835_ (.A(net3990),
    .B(net4673),
    .Y(_05389_));
 sg13g2_a21oi_1 _22836_ (.A1(net5056),
    .A2(net4673),
    .Y(_01812_),
    .B1(_05389_));
 sg13g2_nor2_2 _22837_ (.A(net5425),
    .B(_03077_),
    .Y(_05390_));
 sg13g2_mux2_1 _22838_ (.A0(net3649),
    .A1(net5792),
    .S(_05390_),
    .X(_01813_));
 sg13g2_mux2_1 _22839_ (.A0(net3615),
    .A1(net5757),
    .S(_05390_),
    .X(_01814_));
 sg13g2_mux2_1 _22840_ (.A0(net3228),
    .A1(net5728),
    .S(_05390_),
    .X(_01815_));
 sg13g2_mux2_1 _22841_ (.A0(net3317),
    .A1(net5698),
    .S(_05390_),
    .X(_01816_));
 sg13g2_mux2_1 _22842_ (.A0(net3324),
    .A1(net5673),
    .S(_05390_),
    .X(_01817_));
 sg13g2_mux2_1 _22843_ (.A0(net3715),
    .A1(net5648),
    .S(_05390_),
    .X(_01818_));
 sg13g2_mux2_1 _22844_ (.A0(net3385),
    .A1(net5614),
    .S(_05390_),
    .X(_01819_));
 sg13g2_nor2_1 _22845_ (.A(net4948),
    .B(net4944),
    .Y(_05391_));
 sg13g2_nand2_2 _22846_ (.Y(_05392_),
    .A(net4862),
    .B(_08741_));
 sg13g2_nor2_1 _22847_ (.A(_08606_),
    .B(net4775),
    .Y(_05393_));
 sg13g2_nand2_2 _22848_ (.Y(_05394_),
    .A(_08605_),
    .B(_08753_));
 sg13g2_nor2_1 _22849_ (.A(_05392_),
    .B(_05394_),
    .Y(_05395_));
 sg13g2_nor2_2 _22850_ (.A(_08635_),
    .B(net4775),
    .Y(_05396_));
 sg13g2_nand2b_2 _22851_ (.Y(_05397_),
    .B(_08753_),
    .A_N(_08635_));
 sg13g2_nor2_2 _22852_ (.A(_05392_),
    .B(_05397_),
    .Y(_05398_));
 sg13g2_nand2_2 _22853_ (.Y(_05399_),
    .A(_05391_),
    .B(_05396_));
 sg13g2_nand2_1 _22854_ (.Y(_05400_),
    .A(net6004),
    .B(net4731));
 sg13g2_nand2_1 _22855_ (.Y(_05401_),
    .A(net2947),
    .B(net4670));
 sg13g2_o21ai_1 _22856_ (.B1(_05401_),
    .Y(_01820_),
    .A1(_08005_),
    .A2(net4671));
 sg13g2_nand2_1 _22857_ (.Y(_05402_),
    .A(net2989),
    .B(net4670));
 sg13g2_o21ai_1 _22858_ (.B1(_05402_),
    .Y(_01821_),
    .A1(_08004_),
    .A2(net4670));
 sg13g2_nand2_1 _22859_ (.Y(_05403_),
    .A(net2940),
    .B(net4670));
 sg13g2_o21ai_1 _22860_ (.B1(_05403_),
    .Y(_01822_),
    .A1(_08003_),
    .A2(net4671));
 sg13g2_nand2_1 _22861_ (.Y(_05404_),
    .A(net3054),
    .B(net4670));
 sg13g2_o21ai_1 _22862_ (.B1(_05404_),
    .Y(_01823_),
    .A1(_08002_),
    .A2(net4670));
 sg13g2_mux2_1 _22863_ (.A0(net4317),
    .A1(\atari2600.tia.old_grp1[4] ),
    .S(net4671),
    .X(_01824_));
 sg13g2_mux2_1 _22864_ (.A0(\atari2600.tia.diag[101] ),
    .A1(net6659),
    .S(net4671),
    .X(_01825_));
 sg13g2_nand2_1 _22865_ (.Y(_05405_),
    .A(net2964),
    .B(net4671));
 sg13g2_o21ai_1 _22866_ (.B1(_05405_),
    .Y(_01826_),
    .A1(_08001_),
    .A2(net4671));
 sg13g2_nand2_1 _22867_ (.Y(_05406_),
    .A(net2934),
    .B(net4670));
 sg13g2_o21ai_1 _22868_ (.B1(_05406_),
    .Y(_01827_),
    .A1(_08000_),
    .A2(net4670));
 sg13g2_nor2_2 _22869_ (.A(net5425),
    .B(_03119_),
    .Y(_05407_));
 sg13g2_mux2_1 _22870_ (.A0(net3343),
    .A1(net5792),
    .S(_05407_),
    .X(_01828_));
 sg13g2_mux2_1 _22871_ (.A0(net3361),
    .A1(net5757),
    .S(_05407_),
    .X(_01829_));
 sg13g2_mux2_1 _22872_ (.A0(net4004),
    .A1(net5728),
    .S(_05407_),
    .X(_01830_));
 sg13g2_mux2_1 _22873_ (.A0(net3787),
    .A1(net5698),
    .S(_05407_),
    .X(_01831_));
 sg13g2_mux2_1 _22874_ (.A0(net3251),
    .A1(net5673),
    .S(_05407_),
    .X(_01832_));
 sg13g2_mux2_1 _22875_ (.A0(net3892),
    .A1(net5648),
    .S(_05407_),
    .X(_01833_));
 sg13g2_mux2_1 _22876_ (.A0(net3164),
    .A1(net5614),
    .S(_05407_),
    .X(_01834_));
 sg13g2_a21oi_1 _22877_ (.A1(_08659_),
    .A2(_08666_),
    .Y(_05408_),
    .B1(_08163_));
 sg13g2_o21ai_1 _22878_ (.B1(net5265),
    .Y(_05409_),
    .A1(net5129),
    .A2(net5230));
 sg13g2_and2_1 _22879_ (.A(_08681_),
    .B(_05408_),
    .X(_05410_));
 sg13g2_inv_1 _22880_ (.Y(_05411_),
    .A(_05410_));
 sg13g2_o21ai_1 _22881_ (.B1(net6013),
    .Y(_05412_),
    .A1(_05409_),
    .A2(_05411_));
 sg13g2_a21oi_1 _22882_ (.A1(_08038_),
    .A2(_05411_),
    .Y(_01835_),
    .B1(_05412_));
 sg13g2_o21ai_1 _22883_ (.B1(net6013),
    .Y(_05413_),
    .A1(net7255),
    .A2(_05410_));
 sg13g2_a21oi_1 _22884_ (.A1(_08666_),
    .A2(_05410_),
    .Y(_01836_),
    .B1(_05413_));
 sg13g2_nand3_1 _22885_ (.B(net5129),
    .C(net5238),
    .A(net5265),
    .Y(_05414_));
 sg13g2_o21ai_1 _22886_ (.B1(net6012),
    .Y(_05415_),
    .A1(net7256),
    .A2(_05410_));
 sg13g2_a21oi_1 _22887_ (.A1(_05410_),
    .A2(_05414_),
    .Y(_01837_),
    .B1(_05415_));
 sg13g2_or2_1 _22888_ (.X(_05416_),
    .B(net4723),
    .A(net7324));
 sg13g2_nand2_2 _22889_ (.Y(_05417_),
    .A(net4723),
    .B(_08657_));
 sg13g2_and3_1 _22890_ (.X(_01838_),
    .A(net6029),
    .B(_05416_),
    .C(_05417_));
 sg13g2_nand2_1 _22891_ (.Y(_05418_),
    .A(net7198),
    .B(_08638_));
 sg13g2_nand2_2 _22892_ (.Y(_05419_),
    .A(net6008),
    .B(net5238));
 sg13g2_o21ai_1 _22893_ (.B1(_05418_),
    .Y(_01839_),
    .A1(_05417_),
    .A2(_05419_));
 sg13g2_nand2_1 _22894_ (.Y(_05420_),
    .A(net7184),
    .B(_08638_));
 sg13g2_o21ai_1 _22895_ (.B1(_05420_),
    .Y(_01840_),
    .A1(_05360_),
    .A2(_05417_));
 sg13g2_nand2_1 _22896_ (.Y(_05421_),
    .A(net5837),
    .B(_08638_));
 sg13g2_o21ai_1 _22897_ (.B1(_05421_),
    .Y(_01841_),
    .A1(_05417_),
    .A2(_05419_));
 sg13g2_nand2_1 _22898_ (.Y(_05422_),
    .A(net2924),
    .B(_08638_));
 sg13g2_o21ai_1 _22899_ (.B1(_05422_),
    .Y(_01842_),
    .A1(_05360_),
    .A2(_05417_));
 sg13g2_nand2_1 _22900_ (.Y(_05423_),
    .A(net5835),
    .B(_08682_));
 sg13g2_nand2_2 _22901_ (.Y(_05424_),
    .A(_08657_),
    .B(_08680_));
 sg13g2_o21ai_1 _22902_ (.B1(_05423_),
    .Y(_01843_),
    .A1(_05419_),
    .A2(_05424_));
 sg13g2_nand2_1 _22903_ (.Y(_05425_),
    .A(net5834),
    .B(_08682_));
 sg13g2_o21ai_1 _22904_ (.B1(_05425_),
    .Y(_01844_),
    .A1(_05360_),
    .A2(_05424_));
 sg13g2_o21ai_1 _22905_ (.B1(_05424_),
    .Y(_05426_),
    .A1(net7319),
    .A2(_08681_));
 sg13g2_nor2_1 _22906_ (.A(net5983),
    .B(_05426_),
    .Y(_01845_));
 sg13g2_nand2_1 _22907_ (.Y(_05427_),
    .A(net7154),
    .B(_08682_));
 sg13g2_o21ai_1 _22908_ (.B1(_05427_),
    .Y(_01846_),
    .A1(_05419_),
    .A2(_05424_));
 sg13g2_nand2_1 _22909_ (.Y(_05428_),
    .A(net7145),
    .B(_08682_));
 sg13g2_o21ai_1 _22910_ (.B1(_05428_),
    .Y(_01847_),
    .A1(_05360_),
    .A2(_05424_));
 sg13g2_nand3_1 _22911_ (.B(net6000),
    .C(net4578),
    .A(net7009),
    .Y(_05429_));
 sg13g2_o21ai_1 _22912_ (.B1(_05429_),
    .Y(_01848_),
    .A1(_08565_),
    .A2(net4578));
 sg13g2_nor2_1 _22913_ (.A(net7082),
    .B(net4580),
    .Y(_05430_));
 sg13g2_nor2_1 _22914_ (.A(net4807),
    .B(net4578),
    .Y(_05431_));
 sg13g2_nor3_1 _22915_ (.A(net5980),
    .B(_05430_),
    .C(_05431_),
    .Y(_01849_));
 sg13g2_nor2_1 _22916_ (.A(net6876),
    .B(net4580),
    .Y(_05432_));
 sg13g2_nor2_1 _22917_ (.A(net4845),
    .B(net4578),
    .Y(_05433_));
 sg13g2_nor3_1 _22918_ (.A(net5980),
    .B(_05432_),
    .C(_05433_),
    .Y(_01850_));
 sg13g2_nand2_2 _22919_ (.Y(_05434_),
    .A(net5179),
    .B(net5151));
 sg13g2_o21ai_1 _22920_ (.B1(net6030),
    .Y(_05435_),
    .A1(net7129),
    .A2(net4724));
 sg13g2_a21oi_1 _22921_ (.A1(net4723),
    .A2(_05434_),
    .Y(_01851_),
    .B1(_05435_));
 sg13g2_nand2_2 _22922_ (.Y(_05436_),
    .A(net5193),
    .B(net5151));
 sg13g2_o21ai_1 _22923_ (.B1(net6028),
    .Y(_05437_),
    .A1(net7127),
    .A2(net4723));
 sg13g2_a21oi_1 _22924_ (.A1(net4723),
    .A2(_05436_),
    .Y(_01852_),
    .B1(_05437_));
 sg13g2_nand2_2 _22925_ (.Y(_05438_),
    .A(net5179),
    .B(net5169));
 sg13g2_o21ai_1 _22926_ (.B1(net6030),
    .Y(_05439_),
    .A1(net7177),
    .A2(net4723));
 sg13g2_a21oi_1 _22927_ (.A1(net4723),
    .A2(_05438_),
    .Y(_01853_),
    .B1(_05439_));
 sg13g2_nand2_2 _22928_ (.Y(_05440_),
    .A(net5193),
    .B(net5169));
 sg13g2_o21ai_1 _22929_ (.B1(net6030),
    .Y(_05441_),
    .A1(net7170),
    .A2(net4723));
 sg13g2_a21oi_1 _22930_ (.A1(net4724),
    .A2(_05440_),
    .Y(_01854_),
    .B1(_05441_));
 sg13g2_o21ai_1 _22931_ (.B1(net6007),
    .Y(_05442_),
    .A1(net7152),
    .A2(_08681_));
 sg13g2_a21oi_1 _22932_ (.A1(_08680_),
    .A2(_05434_),
    .Y(_01855_),
    .B1(_05442_));
 sg13g2_o21ai_1 _22933_ (.B1(net6007),
    .Y(_05443_),
    .A1(net7149),
    .A2(_08681_));
 sg13g2_a21oi_1 _22934_ (.A1(_08680_),
    .A2(_05436_),
    .Y(_01856_),
    .B1(_05443_));
 sg13g2_o21ai_1 _22935_ (.B1(net6007),
    .Y(_05444_),
    .A1(net7130),
    .A2(_08681_));
 sg13g2_a21oi_1 _22936_ (.A1(_08680_),
    .A2(_05438_),
    .Y(_01857_),
    .B1(_05444_));
 sg13g2_o21ai_1 _22937_ (.B1(net6007),
    .Y(_05445_),
    .A1(net7207),
    .A2(_08681_));
 sg13g2_a21oi_1 _22938_ (.A1(_08680_),
    .A2(_05440_),
    .Y(_01858_),
    .B1(_05445_));
 sg13g2_nor2_2 _22939_ (.A(_08735_),
    .B(net4944),
    .Y(_05446_));
 sg13g2_nand2_1 _22940_ (.Y(_05447_),
    .A(net4817),
    .B(_08741_));
 sg13g2_nor2_2 _22941_ (.A(_08637_),
    .B(_05447_),
    .Y(_05448_));
 sg13g2_nand2_2 _22942_ (.Y(_05449_),
    .A(_08636_),
    .B(_05446_));
 sg13g2_nand2b_1 _22943_ (.Y(_05450_),
    .B(_05449_),
    .A_N(net7238));
 sg13g2_a21oi_1 _22944_ (.A1(_05434_),
    .A2(_05448_),
    .Y(_05451_),
    .B1(net5992));
 sg13g2_and2_1 _22945_ (.A(_05450_),
    .B(_05451_),
    .X(_01859_));
 sg13g2_nand2b_1 _22946_ (.Y(_05452_),
    .B(_05449_),
    .A_N(net7227));
 sg13g2_a21oi_1 _22947_ (.A1(_05436_),
    .A2(_05448_),
    .Y(_05453_),
    .B1(net5992));
 sg13g2_and2_1 _22948_ (.A(_05452_),
    .B(_05453_),
    .X(_01860_));
 sg13g2_a21o_1 _22949_ (.A2(_05448_),
    .A1(_05438_),
    .B1(net5992),
    .X(_05454_));
 sg13g2_a21oi_1 _22950_ (.A1(_08035_),
    .A2(net4730),
    .Y(_01861_),
    .B1(_05454_));
 sg13g2_nand2b_1 _22951_ (.Y(_05455_),
    .B(net4730),
    .A_N(net7253));
 sg13g2_a21oi_1 _22952_ (.A1(_05440_),
    .A2(_05448_),
    .Y(_05456_),
    .B1(net5992));
 sg13g2_and2_1 _22953_ (.A(_05455_),
    .B(_05456_),
    .X(_01862_));
 sg13g2_nor2_2 _22954_ (.A(_10373_),
    .B(net5425),
    .Y(_05457_));
 sg13g2_mux2_1 _22955_ (.A0(net3167),
    .A1(net5792),
    .S(_05457_),
    .X(_01863_));
 sg13g2_mux2_1 _22956_ (.A0(net3513),
    .A1(net5757),
    .S(_05457_),
    .X(_01864_));
 sg13g2_mux2_1 _22957_ (.A0(net3282),
    .A1(net5728),
    .S(_05457_),
    .X(_01865_));
 sg13g2_mux2_1 _22958_ (.A0(net3428),
    .A1(net5698),
    .S(_05457_),
    .X(_01866_));
 sg13g2_mux2_1 _22959_ (.A0(net3765),
    .A1(net5673),
    .S(_05457_),
    .X(_01867_));
 sg13g2_mux2_1 _22960_ (.A0(net3752),
    .A1(net5648),
    .S(_05457_),
    .X(_01868_));
 sg13g2_mux2_1 _22961_ (.A0(net3142),
    .A1(net5614),
    .S(_05457_),
    .X(_01869_));
 sg13g2_nand2_2 _22962_ (.Y(_05458_),
    .A(net5432),
    .B(net5411));
 sg13g2_mux2_1 _22963_ (.A0(net5773),
    .A1(net6113),
    .S(_05458_),
    .X(_01870_));
 sg13g2_mux2_1 _22964_ (.A0(net5745),
    .A1(net6554),
    .S(_05458_),
    .X(_01871_));
 sg13g2_mux2_1 _22965_ (.A0(net5717),
    .A1(net6597),
    .S(_05458_),
    .X(_01872_));
 sg13g2_mux2_1 _22966_ (.A0(net5689),
    .A1(net6342),
    .S(_05458_),
    .X(_01873_));
 sg13g2_mux2_1 _22967_ (.A0(net5658),
    .A1(net6321),
    .S(_05458_),
    .X(_01874_));
 sg13g2_mux2_1 _22968_ (.A0(net5628),
    .A1(net6517),
    .S(_05458_),
    .X(_01875_));
 sg13g2_mux2_1 _22969_ (.A0(net5601),
    .A1(net4169),
    .S(_05458_),
    .X(_01876_));
 sg13g2_nand2_2 _22970_ (.Y(_05459_),
    .A(_10480_),
    .B(_03124_));
 sg13g2_mux2_1 _22971_ (.A0(net5792),
    .A1(net6858),
    .S(_05459_),
    .X(_01877_));
 sg13g2_mux2_1 _22972_ (.A0(net5757),
    .A1(net6536),
    .S(_05459_),
    .X(_01878_));
 sg13g2_mux2_1 _22973_ (.A0(net5727),
    .A1(net6295),
    .S(_05459_),
    .X(_01879_));
 sg13g2_mux2_1 _22974_ (.A0(net5698),
    .A1(net6466),
    .S(_05459_),
    .X(_01880_));
 sg13g2_mux2_1 _22975_ (.A0(net5673),
    .A1(net6441),
    .S(_05459_),
    .X(_01881_));
 sg13g2_mux2_1 _22976_ (.A0(net5648),
    .A1(net6914),
    .S(_05459_),
    .X(_01882_));
 sg13g2_mux2_1 _22977_ (.A0(net5614),
    .A1(net6241),
    .S(_05459_),
    .X(_01883_));
 sg13g2_nor2_2 _22978_ (.A(net5425),
    .B(_03101_),
    .Y(_05460_));
 sg13g2_mux2_1 _22979_ (.A0(net3551),
    .A1(net5791),
    .S(_05460_),
    .X(_01884_));
 sg13g2_mux2_1 _22980_ (.A0(net4230),
    .A1(net5751),
    .S(_05460_),
    .X(_01885_));
 sg13g2_mux2_1 _22981_ (.A0(net3820),
    .A1(net5727),
    .S(_05460_),
    .X(_01886_));
 sg13g2_mux2_1 _22982_ (.A0(net3891),
    .A1(net5699),
    .S(_05460_),
    .X(_01887_));
 sg13g2_mux2_1 _22983_ (.A0(net4075),
    .A1(net5663),
    .S(_05460_),
    .X(_01888_));
 sg13g2_mux2_1 _22984_ (.A0(net3593),
    .A1(net5636),
    .S(_05460_),
    .X(_01889_));
 sg13g2_mux2_1 _22985_ (.A0(net3238),
    .A1(net5614),
    .S(_05460_),
    .X(_01890_));
 sg13g2_nand2_2 _22986_ (.Y(_05461_),
    .A(_10480_),
    .B(net5419));
 sg13g2_mux2_1 _22987_ (.A0(net5791),
    .A1(net6503),
    .S(_05461_),
    .X(_01891_));
 sg13g2_mux2_1 _22988_ (.A0(net5751),
    .A1(net6544),
    .S(_05461_),
    .X(_01892_));
 sg13g2_mux2_1 _22989_ (.A0(net5727),
    .A1(net6356),
    .S(_05461_),
    .X(_01893_));
 sg13g2_mux2_1 _22990_ (.A0(net5699),
    .A1(net6490),
    .S(_05461_),
    .X(_01894_));
 sg13g2_mux2_1 _22991_ (.A0(net5663),
    .A1(net6929),
    .S(_05461_),
    .X(_01895_));
 sg13g2_mux2_1 _22992_ (.A0(net5636),
    .A1(net6635),
    .S(_05461_),
    .X(_01896_));
 sg13g2_mux2_1 _22993_ (.A0(net5614),
    .A1(net4369),
    .S(_05461_),
    .X(_01897_));
 sg13g2_nand2_2 _22994_ (.Y(_05462_),
    .A(net5469),
    .B(net5411));
 sg13g2_mux2_1 _22995_ (.A0(net5785),
    .A1(net6747),
    .S(_05462_),
    .X(_01898_));
 sg13g2_mux2_1 _22996_ (.A0(net5753),
    .A1(net6735),
    .S(_05462_),
    .X(_01899_));
 sg13g2_mux2_1 _22997_ (.A0(net5724),
    .A1(net4206),
    .S(_05462_),
    .X(_01900_));
 sg13g2_mux2_1 _22998_ (.A0(net5695),
    .A1(net6842),
    .S(_05462_),
    .X(_01901_));
 sg13g2_mux2_1 _22999_ (.A0(net5667),
    .A1(net6913),
    .S(_05462_),
    .X(_01902_));
 sg13g2_mux2_1 _23000_ (.A0(net5639),
    .A1(net6438),
    .S(_05462_),
    .X(_01903_));
 sg13g2_mux2_1 _23001_ (.A0(net5609),
    .A1(net6329),
    .S(_05462_),
    .X(_01904_));
 sg13g2_nand2_2 _23002_ (.Y(_05463_),
    .A(_10480_),
    .B(net5424));
 sg13g2_mux2_1 _23003_ (.A0(net5777),
    .A1(net6899),
    .S(_05463_),
    .X(_01905_));
 sg13g2_mux2_1 _23004_ (.A0(net5751),
    .A1(net6477),
    .S(_05463_),
    .X(_01906_));
 sg13g2_mux2_1 _23005_ (.A0(net5720),
    .A1(net4503),
    .S(_05463_),
    .X(_01907_));
 sg13g2_mux2_1 _23006_ (.A0(net5699),
    .A1(net6430),
    .S(_05463_),
    .X(_01908_));
 sg13g2_mux2_1 _23007_ (.A0(net5663),
    .A1(net6459),
    .S(_05463_),
    .X(_01909_));
 sg13g2_mux2_1 _23008_ (.A0(net5636),
    .A1(net6667),
    .S(_05463_),
    .X(_01910_));
 sg13g2_mux2_1 _23009_ (.A0(net5605),
    .A1(net6893),
    .S(_05463_),
    .X(_01911_));
 sg13g2_nand2_2 _23010_ (.Y(_05464_),
    .A(net4747),
    .B(_03059_));
 sg13g2_mux2_1 _23011_ (.A0(net5256),
    .A1(net4436),
    .S(_05464_),
    .X(_01912_));
 sg13g2_mux2_1 _23012_ (.A0(net5231),
    .A1(net6456),
    .S(_05464_),
    .X(_01913_));
 sg13g2_mux2_1 _23013_ (.A0(net5128),
    .A1(net6289),
    .S(_05464_),
    .X(_01914_));
 sg13g2_mux2_1 _23014_ (.A0(net5100),
    .A1(net6670),
    .S(_05464_),
    .X(_01915_));
 sg13g2_mux2_1 _23015_ (.A0(net5195),
    .A1(net6314),
    .S(_05464_),
    .X(_01916_));
 sg13g2_mux2_1 _23016_ (.A0(net5171),
    .A1(net4266),
    .S(_05464_),
    .X(_01917_));
 sg13g2_mux2_1 _23017_ (.A0(net5076),
    .A1(net4522),
    .S(_05464_),
    .X(_01918_));
 sg13g2_mux2_1 _23018_ (.A0(net5054),
    .A1(net6696),
    .S(_05464_),
    .X(_01919_));
 sg13g2_nor2_1 _23019_ (.A(\flash_rom.addr[8] ),
    .B(net5395),
    .Y(_05465_));
 sg13g2_nor2_1 _23020_ (.A(net4165),
    .B(net5427),
    .Y(_05466_));
 sg13g2_nor3_1 _23021_ (.A(net4570),
    .B(_05465_),
    .C(_05466_),
    .Y(_01920_));
 sg13g2_nor2_1 _23022_ (.A(net3021),
    .B(net5394),
    .Y(_05467_));
 sg13g2_nor2_1 _23023_ (.A(\flash_rom.addr[13] ),
    .B(net5428),
    .Y(_05468_));
 sg13g2_nor3_1 _23024_ (.A(net4570),
    .B(_05467_),
    .C(_05468_),
    .Y(_01921_));
 sg13g2_nor2_1 _23025_ (.A(net4066),
    .B(net5395),
    .Y(_05469_));
 sg13g2_nor2_1 _23026_ (.A(net3646),
    .B(net5427),
    .Y(_05470_));
 sg13g2_nor3_1 _23027_ (.A(net4570),
    .B(_05469_),
    .C(_05470_),
    .Y(_01922_));
 sg13g2_nor2_1 _23028_ (.A(net3846),
    .B(net5395),
    .Y(_05471_));
 sg13g2_nor2_1 _23029_ (.A(\flash_rom.addr[15] ),
    .B(net5427),
    .Y(_05472_));
 sg13g2_nor3_1 _23030_ (.A(net4570),
    .B(_05471_),
    .C(_05472_),
    .Y(_01923_));
 sg13g2_nand2_1 _23031_ (.Y(_05473_),
    .A(_08034_),
    .B(net5394));
 sg13g2_o21ai_1 _23032_ (.B1(_05473_),
    .Y(_05474_),
    .A1(net4221),
    .A2(net5394));
 sg13g2_nand2b_1 _23033_ (.Y(_01924_),
    .B(_05474_),
    .A_N(net4571));
 sg13g2_nor2_2 _23034_ (.A(net5472),
    .B(_10499_),
    .Y(_05475_));
 sg13g2_mux2_1 _23035_ (.A0(net3995),
    .A1(net5775),
    .S(_05475_),
    .X(_01925_));
 sg13g2_mux2_1 _23036_ (.A0(net3742),
    .A1(net5747),
    .S(_05475_),
    .X(_01926_));
 sg13g2_mux2_1 _23037_ (.A0(net3907),
    .A1(net5721),
    .S(_05475_),
    .X(_01927_));
 sg13g2_mux2_1 _23038_ (.A0(net3756),
    .A1(net5690),
    .S(_05475_),
    .X(_01928_));
 sg13g2_mux2_1 _23039_ (.A0(net3782),
    .A1(net5660),
    .S(_05475_),
    .X(_01929_));
 sg13g2_mux2_1 _23040_ (.A0(net3626),
    .A1(net5632),
    .S(_05475_),
    .X(_01930_));
 sg13g2_mux2_1 _23041_ (.A0(net3848),
    .A1(net5603),
    .S(_05475_),
    .X(_01931_));
 sg13g2_nor2_2 _23042_ (.A(_10499_),
    .B(net5471),
    .Y(_05476_));
 sg13g2_mux2_1 _23043_ (.A0(net3655),
    .A1(net5777),
    .S(_05476_),
    .X(_01932_));
 sg13g2_mux2_1 _23044_ (.A0(net3264),
    .A1(net5747),
    .S(_05476_),
    .X(_01933_));
 sg13g2_mux2_1 _23045_ (.A0(net3423),
    .A1(net5718),
    .S(_05476_),
    .X(_01934_));
 sg13g2_mux2_1 _23046_ (.A0(net3259),
    .A1(net5688),
    .S(_05476_),
    .X(_01935_));
 sg13g2_mux2_1 _23047_ (.A0(net3886),
    .A1(net5660),
    .S(_05476_),
    .X(_01936_));
 sg13g2_mux2_1 _23048_ (.A0(net3819),
    .A1(net5632),
    .S(_05476_),
    .X(_01937_));
 sg13g2_mux2_1 _23049_ (.A0(net3640),
    .A1(net5603),
    .S(_05476_),
    .X(_01938_));
 sg13g2_nor2_2 _23050_ (.A(_10499_),
    .B(net5467),
    .Y(_05477_));
 sg13g2_mux2_1 _23051_ (.A0(net3605),
    .A1(net5777),
    .S(_05477_),
    .X(_01939_));
 sg13g2_mux2_1 _23052_ (.A0(net3182),
    .A1(net5747),
    .S(_05477_),
    .X(_01940_));
 sg13g2_mux2_1 _23053_ (.A0(net3107),
    .A1(net5718),
    .S(_05477_),
    .X(_01941_));
 sg13g2_mux2_1 _23054_ (.A0(net3785),
    .A1(net5688),
    .S(_05477_),
    .X(_01942_));
 sg13g2_mux2_1 _23055_ (.A0(net3291),
    .A1(net5660),
    .S(_05477_),
    .X(_01943_));
 sg13g2_mux2_1 _23056_ (.A0(net3152),
    .A1(net5632),
    .S(_05477_),
    .X(_01944_));
 sg13g2_mux2_1 _23057_ (.A0(net3654),
    .A1(net5603),
    .S(_05477_),
    .X(_01945_));
 sg13g2_nand2_2 _23058_ (.Y(_05478_),
    .A(net5423),
    .B(net5468));
 sg13g2_mux2_1 _23059_ (.A0(net5777),
    .A1(net6149),
    .S(_05478_),
    .X(_01946_));
 sg13g2_mux2_1 _23060_ (.A0(net5747),
    .A1(net6947),
    .S(_05478_),
    .X(_01947_));
 sg13g2_mux2_1 _23061_ (.A0(net5718),
    .A1(net6614),
    .S(_05478_),
    .X(_01948_));
 sg13g2_mux2_1 _23062_ (.A0(net5688),
    .A1(net6884),
    .S(_05478_),
    .X(_01949_));
 sg13g2_mux2_1 _23063_ (.A0(net5660),
    .A1(net6715),
    .S(_05478_),
    .X(_01950_));
 sg13g2_mux2_1 _23064_ (.A0(net5632),
    .A1(net6097),
    .S(_05478_),
    .X(_01951_));
 sg13g2_mux2_1 _23065_ (.A0(net5603),
    .A1(net6502),
    .S(_05478_),
    .X(_01952_));
 sg13g2_nand2_2 _23066_ (.Y(_05479_),
    .A(net4739),
    .B(_05073_));
 sg13g2_mux2_1 _23067_ (.A0(net5248),
    .A1(net4251),
    .S(_05479_),
    .X(_01953_));
 sg13g2_mux2_1 _23068_ (.A0(net5221),
    .A1(net4386),
    .S(_05479_),
    .X(_01954_));
 sg13g2_mux2_1 _23069_ (.A0(net5116),
    .A1(net4140),
    .S(_05479_),
    .X(_01955_));
 sg13g2_mux2_1 _23070_ (.A0(net5092),
    .A1(net4462),
    .S(_05479_),
    .X(_01956_));
 sg13g2_mux2_1 _23071_ (.A0(net5187),
    .A1(net4101),
    .S(_05479_),
    .X(_01957_));
 sg13g2_mux2_1 _23072_ (.A0(net5159),
    .A1(net6078),
    .S(_05479_),
    .X(_01958_));
 sg13g2_mux2_1 _23073_ (.A0(net5066),
    .A1(net4149),
    .S(_05479_),
    .X(_01959_));
 sg13g2_mux2_1 _23074_ (.A0(net5044),
    .A1(net4082),
    .S(_05479_),
    .X(_01960_));
 sg13g2_nor2_1 _23075_ (.A(net4743),
    .B(_04814_),
    .Y(_05480_));
 sg13g2_nor2_1 _23076_ (.A(net3899),
    .B(net4668),
    .Y(_05481_));
 sg13g2_a21oi_1 _23077_ (.A1(net5262),
    .A2(net4668),
    .Y(_01961_),
    .B1(_05481_));
 sg13g2_nor2_1 _23078_ (.A(net3269),
    .B(net4668),
    .Y(_05482_));
 sg13g2_a21oi_1 _23079_ (.A1(net5235),
    .A2(net4668),
    .Y(_01962_),
    .B1(_05482_));
 sg13g2_nor2_1 _23080_ (.A(net3969),
    .B(net4668),
    .Y(_05483_));
 sg13g2_a21oi_1 _23081_ (.A1(net5132),
    .A2(net4668),
    .Y(_01963_),
    .B1(_05483_));
 sg13g2_nor2_1 _23082_ (.A(net3304),
    .B(net4668),
    .Y(_05484_));
 sg13g2_a21oi_1 _23083_ (.A1(net5104),
    .A2(net4668),
    .Y(_01964_),
    .B1(_05484_));
 sg13g2_nor2_1 _23084_ (.A(net3797),
    .B(net4669),
    .Y(_05485_));
 sg13g2_a21oi_1 _23085_ (.A1(net5178),
    .A2(net4669),
    .Y(_01965_),
    .B1(_05485_));
 sg13g2_nor2_1 _23086_ (.A(net3660),
    .B(net4669),
    .Y(_05486_));
 sg13g2_a21oi_1 _23087_ (.A1(net5147),
    .A2(net4669),
    .Y(_01966_),
    .B1(_05486_));
 sg13g2_nor2_1 _23088_ (.A(net3485),
    .B(net4669),
    .Y(_05487_));
 sg13g2_a21oi_1 _23089_ (.A1(net5079),
    .A2(net4669),
    .Y(_01967_),
    .B1(_05487_));
 sg13g2_nor2_1 _23090_ (.A(net3147),
    .B(net4669),
    .Y(_05488_));
 sg13g2_a21oi_1 _23091_ (.A1(net5056),
    .A2(net4669),
    .Y(_01968_),
    .B1(_05488_));
 sg13g2_nand2_2 _23092_ (.Y(_05489_),
    .A(_03041_),
    .B(net4733));
 sg13g2_mux2_1 _23093_ (.A0(net5251),
    .A1(net4095),
    .S(_05489_),
    .X(_01969_));
 sg13g2_mux2_1 _23094_ (.A0(net5225),
    .A1(net4390),
    .S(_05489_),
    .X(_01970_));
 sg13g2_mux2_1 _23095_ (.A0(net5124),
    .A1(net6716),
    .S(_05489_),
    .X(_01971_));
 sg13g2_mux2_1 _23096_ (.A0(net5096),
    .A1(net4079),
    .S(_05489_),
    .X(_01972_));
 sg13g2_mux2_1 _23097_ (.A0(net5191),
    .A1(net4405),
    .S(_05489_),
    .X(_01973_));
 sg13g2_mux2_1 _23098_ (.A0(net5163),
    .A1(net6257),
    .S(_05489_),
    .X(_01974_));
 sg13g2_mux2_1 _23099_ (.A0(net5071),
    .A1(net4121),
    .S(_05489_),
    .X(_01975_));
 sg13g2_mux2_1 _23100_ (.A0(net5045),
    .A1(net4524),
    .S(_05489_),
    .X(_01976_));
 sg13g2_nand2_2 _23101_ (.Y(_05490_),
    .A(_10478_),
    .B(net5422));
 sg13g2_mux2_1 _23102_ (.A0(net5781),
    .A1(net6558),
    .S(_05490_),
    .X(_01977_));
 sg13g2_mux2_1 _23103_ (.A0(net5752),
    .A1(net6812),
    .S(_05490_),
    .X(_01978_));
 sg13g2_mux2_1 _23104_ (.A0(net5722),
    .A1(net6112),
    .S(_05490_),
    .X(_01979_));
 sg13g2_mux2_1 _23105_ (.A0(net5693),
    .A1(net6576),
    .S(_05490_),
    .X(_01980_));
 sg13g2_mux2_1 _23106_ (.A0(net5659),
    .A1(net6669),
    .S(_05490_),
    .X(_01981_));
 sg13g2_mux2_1 _23107_ (.A0(net5630),
    .A1(net6622),
    .S(_05490_),
    .X(_01982_));
 sg13g2_mux2_1 _23108_ (.A0(net5602),
    .A1(net4483),
    .S(_05490_),
    .X(_01983_));
 sg13g2_nand2_2 _23109_ (.Y(_05491_),
    .A(_10381_),
    .B(net5422));
 sg13g2_mux2_1 _23110_ (.A0(net5781),
    .A1(net6823),
    .S(_05491_),
    .X(_01984_));
 sg13g2_mux2_1 _23111_ (.A0(net5752),
    .A1(net6672),
    .S(_05491_),
    .X(_01985_));
 sg13g2_mux2_1 _23112_ (.A0(net5722),
    .A1(net6574),
    .S(_05491_),
    .X(_01986_));
 sg13g2_mux2_1 _23113_ (.A0(net5693),
    .A1(net6433),
    .S(_05491_),
    .X(_01987_));
 sg13g2_mux2_1 _23114_ (.A0(net5659),
    .A1(net6096),
    .S(_05491_),
    .X(_01988_));
 sg13g2_mux2_1 _23115_ (.A0(net5630),
    .A1(net6389),
    .S(_05491_),
    .X(_01989_));
 sg13g2_mux2_1 _23116_ (.A0(net5602),
    .A1(net6322),
    .S(_05491_),
    .X(_01990_));
 sg13g2_nand2_2 _23117_ (.Y(_05492_),
    .A(net5422),
    .B(_02995_));
 sg13g2_mux2_1 _23118_ (.A0(net5781),
    .A1(net4447),
    .S(_05492_),
    .X(_01991_));
 sg13g2_mux2_1 _23119_ (.A0(net5752),
    .A1(net6709),
    .S(_05492_),
    .X(_01992_));
 sg13g2_mux2_1 _23120_ (.A0(net5718),
    .A1(net6522),
    .S(_05492_),
    .X(_01993_));
 sg13g2_mux2_1 _23121_ (.A0(net5693),
    .A1(net6381),
    .S(_05492_),
    .X(_01994_));
 sg13g2_mux2_1 _23122_ (.A0(net5659),
    .A1(net6793),
    .S(_05492_),
    .X(_01995_));
 sg13g2_mux2_1 _23123_ (.A0(net5630),
    .A1(net6682),
    .S(_05492_),
    .X(_01996_));
 sg13g2_mux2_1 _23124_ (.A0(net5602),
    .A1(net6851),
    .S(_05492_),
    .X(_01997_));
 sg13g2_nand2_2 _23125_ (.Y(_05493_),
    .A(net5422),
    .B(net5412));
 sg13g2_mux2_1 _23126_ (.A0(net5781),
    .A1(net6374),
    .S(_05493_),
    .X(_01998_));
 sg13g2_mux2_1 _23127_ (.A0(net5747),
    .A1(net6133),
    .S(_05493_),
    .X(_01999_));
 sg13g2_mux2_1 _23128_ (.A0(net5717),
    .A1(net4426),
    .S(_05493_),
    .X(_02000_));
 sg13g2_mux2_1 _23129_ (.A0(net5689),
    .A1(net6809),
    .S(_05493_),
    .X(_02001_));
 sg13g2_mux2_1 _23130_ (.A0(net5659),
    .A1(net6385),
    .S(_05493_),
    .X(_02002_));
 sg13g2_mux2_1 _23131_ (.A0(net5630),
    .A1(net6319),
    .S(_05493_),
    .X(_02003_));
 sg13g2_mux2_1 _23132_ (.A0(net5602),
    .A1(net4455),
    .S(_05493_),
    .X(_02004_));
 sg13g2_nand2_2 _23133_ (.Y(_05494_),
    .A(net5469),
    .B(_03100_));
 sg13g2_mux2_1 _23134_ (.A0(net5787),
    .A1(net6681),
    .S(_05494_),
    .X(_02005_));
 sg13g2_mux2_1 _23135_ (.A0(net5754),
    .A1(net6904),
    .S(_05494_),
    .X(_02006_));
 sg13g2_mux2_1 _23136_ (.A0(net5731),
    .A1(net6888),
    .S(_05494_),
    .X(_02007_));
 sg13g2_mux2_1 _23137_ (.A0(net5705),
    .A1(net6320),
    .S(_05494_),
    .X(_02008_));
 sg13g2_mux2_1 _23138_ (.A0(net5668),
    .A1(net6643),
    .S(_05494_),
    .X(_02009_));
 sg13g2_mux2_1 _23139_ (.A0(net5638),
    .A1(net6243),
    .S(_05494_),
    .X(_02010_));
 sg13g2_mux2_1 _23140_ (.A0(net5609),
    .A1(net6924),
    .S(_05494_),
    .X(_02011_));
 sg13g2_nor2_1 _23141_ (.A(net5989),
    .B(net5354),
    .Y(_05495_));
 sg13g2_nand2_1 _23142_ (.Y(_05496_),
    .A(\atari2600.tia.audio_left_counter[0] ),
    .B(net5280));
 sg13g2_nor2_2 _23143_ (.A(\atari2600.tia.audc0[3] ),
    .B(\atari2600.tia.audc0[2] ),
    .Y(_05497_));
 sg13g2_nor2_1 _23144_ (.A(\atari2600.tia.audc0[1] ),
    .B(\atari2600.tia.audc0[0] ),
    .Y(_05498_));
 sg13g2_nand2_1 _23145_ (.Y(_05499_),
    .A(_05497_),
    .B(_05498_));
 sg13g2_nor2b_1 _23146_ (.A(\atari2600.tia.audc0[2] ),
    .B_N(\atari2600.tia.audc0[3] ),
    .Y(_05500_));
 sg13g2_nand3_1 _23147_ (.B(\atari2600.tia.audc0[0] ),
    .C(_05500_),
    .A(\atari2600.tia.audc0[1] ),
    .Y(_05501_));
 sg13g2_nand2_2 _23148_ (.Y(_05502_),
    .A(_05499_),
    .B(_05501_));
 sg13g2_and4_2 _23149_ (.A(\atari2600.tia.audf0[3] ),
    .B(\atari2600.tia.audf0[2] ),
    .C(\atari2600.tia.audf0[1] ),
    .D(net5582),
    .X(_05503_));
 sg13g2_nand4_1 _23150_ (.B(\atari2600.tia.audf0[2] ),
    .C(\atari2600.tia.audf0[1] ),
    .A(\atari2600.tia.audf0[3] ),
    .Y(_05504_),
    .D(net5582));
 sg13g2_and3_1 _23151_ (.X(_05505_),
    .A(\atari2600.tia.audf0[2] ),
    .B(\atari2600.tia.audf0[1] ),
    .C(net5582));
 sg13g2_o21ai_1 _23152_ (.B1(_05504_),
    .Y(_05506_),
    .A1(\atari2600.tia.audf0[3] ),
    .A2(_05505_));
 sg13g2_inv_1 _23153_ (.Y(_05507_),
    .A(_05506_));
 sg13g2_a21oi_1 _23154_ (.A1(\atari2600.tia.audf0[1] ),
    .A2(net5582),
    .Y(_05508_),
    .B1(\atari2600.tia.audf0[2] ));
 sg13g2_nor2_1 _23155_ (.A(_05505_),
    .B(_05508_),
    .Y(_05509_));
 sg13g2_nor2_1 _23156_ (.A(_00112_),
    .B(_05506_),
    .Y(_05510_));
 sg13g2_a21oi_1 _23157_ (.A1(\atari2600.tia.audf0[4] ),
    .A2(_05503_),
    .Y(_05511_),
    .B1(_05510_));
 sg13g2_nor2b_1 _23158_ (.A(_05511_),
    .B_N(_05509_),
    .Y(_05512_));
 sg13g2_nand2b_1 _23159_ (.Y(_05513_),
    .B(_05507_),
    .A_N(_05512_));
 sg13g2_xor2_1 _23160_ (.B(net5582),
    .A(\atari2600.tia.audf0[1] ),
    .X(_05514_));
 sg13g2_nand2_1 _23161_ (.Y(_05515_),
    .A(\atari2600.tia.audf0[3] ),
    .B(_05509_));
 sg13g2_nor4_1 _23162_ (.A(_07951_),
    .B(_08100_),
    .C(_05505_),
    .D(_05508_),
    .Y(_05516_));
 sg13g2_nand2_1 _23163_ (.Y(_05517_),
    .A(_00112_),
    .B(_05504_));
 sg13g2_a21o_1 _23164_ (.A2(_05517_),
    .A1(_05506_),
    .B1(_05516_),
    .X(_05518_));
 sg13g2_nand2_2 _23165_ (.Y(_05519_),
    .A(_05514_),
    .B(_05518_));
 sg13g2_xor2_1 _23166_ (.B(_05511_),
    .A(_05509_),
    .X(_05520_));
 sg13g2_nor2_1 _23167_ (.A(_05519_),
    .B(_05520_),
    .Y(_05521_));
 sg13g2_or2_1 _23168_ (.X(_05522_),
    .B(_05520_),
    .A(_05519_));
 sg13g2_nor4_2 _23169_ (.A(_07951_),
    .B(\atari2600.tia.audf0[2] ),
    .C(_07953_),
    .Y(_05523_),
    .D(net5582));
 sg13g2_nand2_1 _23170_ (.Y(_05524_),
    .A(\atari2600.tia.audf0[2] ),
    .B(_05514_));
 sg13g2_inv_1 _23171_ (.Y(_05525_),
    .A(_05524_));
 sg13g2_xnor2_1 _23172_ (.Y(_05526_),
    .A(_00112_),
    .B(_05503_));
 sg13g2_xnor2_1 _23173_ (.Y(_05527_),
    .A(_08100_),
    .B(_05503_));
 sg13g2_mux2_1 _23174_ (.A0(_00112_),
    .A1(_05526_),
    .S(_05506_),
    .X(_05528_));
 sg13g2_mux2_1 _23175_ (.A0(_08100_),
    .A1(_05527_),
    .S(_05506_),
    .X(_05529_));
 sg13g2_nand3_1 _23176_ (.B(_05525_),
    .C(_05528_),
    .A(_07951_),
    .Y(_05530_));
 sg13g2_a221oi_1 _23177_ (.B2(_05515_),
    .C1(_05516_),
    .B1(_05529_),
    .A1(_07951_),
    .Y(_05531_),
    .A2(_05525_));
 sg13g2_nor3_1 _23178_ (.A(\atari2600.tia.audf0[3] ),
    .B(_05524_),
    .C(_05528_),
    .Y(_05532_));
 sg13g2_o21ai_1 _23179_ (.B1(_00107_),
    .Y(_05533_),
    .A1(_05531_),
    .A2(_05532_));
 sg13g2_or3_1 _23180_ (.A(_00107_),
    .B(_05531_),
    .C(_05532_),
    .X(_05534_));
 sg13g2_and3_1 _23181_ (.X(_05535_),
    .A(_05523_),
    .B(_05533_),
    .C(_05534_));
 sg13g2_nand3_1 _23182_ (.B(_05533_),
    .C(_05534_),
    .A(_05523_),
    .Y(_05536_));
 sg13g2_xnor2_1 _23183_ (.Y(_05537_),
    .A(_05514_),
    .B(_05518_));
 sg13g2_a21oi_2 _23184_ (.B1(_05537_),
    .Y(_05538_),
    .A2(_05533_),
    .A1(_05530_));
 sg13g2_a21o_1 _23185_ (.A2(_05533_),
    .A1(_05530_),
    .B1(_05537_),
    .X(_05539_));
 sg13g2_xor2_1 _23186_ (.B(_05520_),
    .A(_05519_),
    .X(_05540_));
 sg13g2_xnor2_1 _23187_ (.Y(_05541_),
    .A(_05519_),
    .B(_05520_));
 sg13g2_a21oi_2 _23188_ (.B1(_05541_),
    .Y(_05542_),
    .A2(_05539_),
    .A1(_05536_));
 sg13g2_o21ai_1 _23189_ (.B1(_05540_),
    .Y(_05543_),
    .A1(_05535_),
    .A2(_05538_));
 sg13g2_a21oi_2 _23190_ (.B1(_05513_),
    .Y(_05544_),
    .A2(_05543_),
    .A1(_05522_));
 sg13g2_and3_1 _23191_ (.X(_05545_),
    .A(_05513_),
    .B(_05522_),
    .C(_05543_));
 sg13g2_nor2_2 _23192_ (.A(_05544_),
    .B(_05545_),
    .Y(_05546_));
 sg13g2_o21ai_1 _23193_ (.B1(_05510_),
    .Y(_05547_),
    .A1(_05535_),
    .A2(_05538_));
 sg13g2_a21oi_1 _23194_ (.A1(_05507_),
    .A2(_05521_),
    .Y(_05548_),
    .B1(_05512_));
 sg13g2_a21oi_2 _23195_ (.B1(_05527_),
    .Y(_05549_),
    .A2(_05548_),
    .A1(_05547_));
 sg13g2_and3_1 _23196_ (.X(_05550_),
    .A(_05527_),
    .B(_05547_),
    .C(_05548_));
 sg13g2_nor2_2 _23197_ (.A(_05549_),
    .B(_05550_),
    .Y(_05551_));
 sg13g2_nor2_2 _23198_ (.A(_07967_),
    .B(\atari2600.tia.audc0[0] ),
    .Y(_05552_));
 sg13g2_nand2_2 _23199_ (.Y(_05553_),
    .A(\atari2600.tia.audc0[1] ),
    .B(_07968_));
 sg13g2_nor2_2 _23200_ (.A(_05497_),
    .B(_05553_),
    .Y(_05554_));
 sg13g2_nand2b_2 _23201_ (.Y(_05555_),
    .B(net5454),
    .A_N(_05497_));
 sg13g2_nand2_1 _23202_ (.Y(_05556_),
    .A(_05551_),
    .B(_05552_));
 sg13g2_nand2_1 _23203_ (.Y(_05557_),
    .A(_05546_),
    .B(net5454));
 sg13g2_nand2_1 _23204_ (.Y(_05558_),
    .A(_05546_),
    .B(_05554_));
 sg13g2_nor3_1 _23205_ (.A(_05549_),
    .B(_05550_),
    .C(_05558_),
    .Y(_05559_));
 sg13g2_a21o_2 _23206_ (.A2(_05503_),
    .A1(_08100_),
    .B1(_05549_),
    .X(_05560_));
 sg13g2_a22oi_1 _23207_ (.Y(_05561_),
    .B1(_05560_),
    .B2(net5454),
    .A2(_05554_),
    .A1(_05551_));
 sg13g2_nor2_1 _23208_ (.A(_05559_),
    .B(_05561_),
    .Y(_05562_));
 sg13g2_and2_2 _23209_ (.A(\atari2600.tia.audc0[3] ),
    .B(\atari2600.tia.audc0[2] ),
    .X(_05563_));
 sg13g2_nand2_1 _23210_ (.Y(_05564_),
    .A(\atari2600.tia.audc0[3] ),
    .B(\atari2600.tia.audc0[2] ));
 sg13g2_nor2_2 _23211_ (.A(net5454),
    .B(_05563_),
    .Y(_05565_));
 sg13g2_nand2_2 _23212_ (.Y(_05566_),
    .A(_05553_),
    .B(net5482));
 sg13g2_a21oi_1 _23213_ (.A1(_05556_),
    .A2(_05558_),
    .Y(_05567_),
    .B1(_05559_));
 sg13g2_a21oi_2 _23214_ (.B1(_05567_),
    .Y(_05568_),
    .A2(_05566_),
    .A1(_05560_));
 sg13g2_nand2_1 _23215_ (.Y(_05569_),
    .A(\atari2600.tia.audc0[2] ),
    .B(_07967_));
 sg13g2_o21ai_1 _23216_ (.B1(_05569_),
    .Y(_05570_),
    .A1(_07968_),
    .A2(net5482));
 sg13g2_a22oi_1 _23217_ (.Y(_05571_),
    .B1(\atari2600.tia.audc0[0] ),
    .B2(_05563_),
    .A2(_07967_),
    .A1(\atari2600.tia.audc0[2] ));
 sg13g2_a21oi_2 _23218_ (.B1(_05570_),
    .Y(_05572_),
    .A2(net5482),
    .A1(_05552_));
 sg13g2_o21ai_1 _23219_ (.B1(_05571_),
    .Y(_05573_),
    .A1(net5453),
    .A2(_05563_));
 sg13g2_a22oi_1 _23220_ (.Y(_05574_),
    .B1(_05573_),
    .B2(_05551_),
    .A2(_05571_),
    .A1(_05560_));
 sg13g2_nand2_1 _23221_ (.Y(_05575_),
    .A(_05546_),
    .B(_05566_));
 sg13g2_nor2_1 _23222_ (.A(_05574_),
    .B(_05575_),
    .Y(_05576_));
 sg13g2_a22oi_1 _23223_ (.Y(_05577_),
    .B1(_05573_),
    .B2(_05560_),
    .A2(_05566_),
    .A1(_05551_));
 sg13g2_nor2_1 _23224_ (.A(_05576_),
    .B(_05577_),
    .Y(_05578_));
 sg13g2_nor3_2 _23225_ (.A(_05535_),
    .B(_05538_),
    .C(_05540_),
    .Y(_05579_));
 sg13g2_nor2_2 _23226_ (.A(_05542_),
    .B(_05579_),
    .Y(_05580_));
 sg13g2_nand2_1 _23227_ (.Y(_05581_),
    .A(net5454),
    .B(_05580_));
 sg13g2_nand3_1 _23228_ (.B(_05554_),
    .C(_05580_),
    .A(_05546_),
    .Y(_05582_));
 sg13g2_o21ai_1 _23229_ (.B1(_05557_),
    .Y(_05583_),
    .A1(_05497_),
    .A2(_05581_));
 sg13g2_and2_1 _23230_ (.A(_05582_),
    .B(_05583_),
    .X(_05584_));
 sg13g2_a21o_1 _23231_ (.A2(_05584_),
    .A1(_05578_),
    .B1(_05576_),
    .X(_05585_));
 sg13g2_nand2b_1 _23232_ (.Y(_05586_),
    .B(_05585_),
    .A_N(_05568_));
 sg13g2_xor2_1 _23233_ (.B(_05585_),
    .A(_05568_),
    .X(_05587_));
 sg13g2_o21ai_1 _23234_ (.B1(_05586_),
    .Y(_05588_),
    .A1(_05582_),
    .A2(_05587_));
 sg13g2_and2_1 _23235_ (.A(_05562_),
    .B(_05588_),
    .X(_05589_));
 sg13g2_nor2_1 _23236_ (.A(net5482),
    .B(_05581_),
    .Y(_05590_));
 sg13g2_xor2_1 _23237_ (.B(_05588_),
    .A(_05562_),
    .X(_05591_));
 sg13g2_a21oi_1 _23238_ (.A1(_05590_),
    .A2(_05591_),
    .Y(_05592_),
    .B1(_05589_));
 sg13g2_a21oi_1 _23239_ (.A1(_05554_),
    .A2(_05560_),
    .Y(_05593_),
    .B1(_05559_));
 sg13g2_nor2_1 _23240_ (.A(_05557_),
    .B(net5481),
    .Y(_05594_));
 sg13g2_nor2b_1 _23241_ (.A(_05593_),
    .B_N(_05594_),
    .Y(_05595_));
 sg13g2_xnor2_1 _23242_ (.Y(_05596_),
    .A(_05593_),
    .B(_05594_));
 sg13g2_nand2b_1 _23243_ (.Y(_05597_),
    .B(_05596_),
    .A_N(_05592_));
 sg13g2_xnor2_1 _23244_ (.Y(_05598_),
    .A(_05592_),
    .B(_05596_));
 sg13g2_xor2_1 _23245_ (.B(_05575_),
    .A(_05574_),
    .X(_05599_));
 sg13g2_nor3_1 _23246_ (.A(_05544_),
    .B(_05545_),
    .C(_05570_),
    .Y(_05600_));
 sg13g2_nor3_1 _23247_ (.A(_05549_),
    .B(_05550_),
    .C(_05570_),
    .Y(_05601_));
 sg13g2_nor3_2 _23248_ (.A(_05544_),
    .B(_05545_),
    .C(_05572_),
    .Y(_05602_));
 sg13g2_nand2_1 _23249_ (.Y(_05603_),
    .A(_05601_),
    .B(_05602_));
 sg13g2_nand2_1 _23250_ (.Y(_05604_),
    .A(_05566_),
    .B(_05580_));
 sg13g2_xnor2_1 _23251_ (.Y(_05605_),
    .A(_05601_),
    .B(_05602_));
 sg13g2_o21ai_1 _23252_ (.B1(_05603_),
    .Y(_05606_),
    .A1(_05604_),
    .A2(_05605_));
 sg13g2_nand2_1 _23253_ (.Y(_05607_),
    .A(_05599_),
    .B(_05606_));
 sg13g2_nand3_1 _23254_ (.B(_05533_),
    .C(_05537_),
    .A(_05530_),
    .Y(_05608_));
 sg13g2_nand3_1 _23255_ (.B(_05539_),
    .C(_05608_),
    .A(_05536_),
    .Y(_05609_));
 sg13g2_nor2_1 _23256_ (.A(net5453),
    .B(_05609_),
    .Y(_05610_));
 sg13g2_or2_1 _23257_ (.X(_05611_),
    .B(_05609_),
    .A(_05555_));
 sg13g2_nor3_2 _23258_ (.A(_05542_),
    .B(_05579_),
    .C(_05611_),
    .Y(_05612_));
 sg13g2_a21o_1 _23259_ (.A2(_05611_),
    .A1(_05581_),
    .B1(_05612_),
    .X(_05613_));
 sg13g2_xnor2_1 _23260_ (.Y(_05614_),
    .A(_05599_),
    .B(_05606_));
 sg13g2_o21ai_1 _23261_ (.B1(_05607_),
    .Y(_05615_),
    .A1(_05613_),
    .A2(_05614_));
 sg13g2_xnor2_1 _23262_ (.Y(_05616_),
    .A(_05578_),
    .B(_05584_));
 sg13g2_nor2b_1 _23263_ (.A(_05616_),
    .B_N(_05615_),
    .Y(_05617_));
 sg13g2_xor2_1 _23264_ (.B(_05616_),
    .A(_05615_),
    .X(_05618_));
 sg13g2_inv_1 _23265_ (.Y(_05619_),
    .A(_05618_));
 sg13g2_a21oi_1 _23266_ (.A1(_05612_),
    .A2(_05619_),
    .Y(_05620_),
    .B1(_05617_));
 sg13g2_xor2_1 _23267_ (.B(_05587_),
    .A(_05582_),
    .X(_05621_));
 sg13g2_nor2b_1 _23268_ (.A(_05620_),
    .B_N(_05621_),
    .Y(_05622_));
 sg13g2_nor3_2 _23269_ (.A(_05553_),
    .B(net5481),
    .C(_05609_),
    .Y(_05623_));
 sg13g2_xnor2_1 _23270_ (.Y(_05624_),
    .A(_05620_),
    .B(_05621_));
 sg13g2_a21oi_1 _23271_ (.A1(_05623_),
    .A2(_05624_),
    .Y(_05625_),
    .B1(_05622_));
 sg13g2_xnor2_1 _23272_ (.Y(_05626_),
    .A(_05590_),
    .B(_05591_));
 sg13g2_nor2_1 _23273_ (.A(_05625_),
    .B(_05626_),
    .Y(_05627_));
 sg13g2_a21oi_1 _23274_ (.A1(_07952_),
    .A2(_07953_),
    .Y(_05628_),
    .B1(_05525_));
 sg13g2_xnor2_1 _23275_ (.Y(_05629_),
    .A(\atari2600.tia.audf0[3] ),
    .B(_05628_));
 sg13g2_xnor2_1 _23276_ (.Y(_05630_),
    .A(_07951_),
    .B(_05628_));
 sg13g2_nand2_1 _23277_ (.Y(_05631_),
    .A(_05573_),
    .B(_05630_));
 sg13g2_xnor2_1 _23278_ (.Y(_05632_),
    .A(\atari2600.tia.audf0[2] ),
    .B(net5582));
 sg13g2_nor2_1 _23279_ (.A(net5401),
    .B(_05632_),
    .Y(_05633_));
 sg13g2_nor2_1 _23280_ (.A(net5401),
    .B(_05629_),
    .Y(_05634_));
 sg13g2_nor2_1 _23281_ (.A(_05572_),
    .B(_05632_),
    .Y(_05635_));
 sg13g2_xnor2_1 _23282_ (.Y(_05636_),
    .A(_00107_),
    .B(_05514_));
 sg13g2_xnor2_1 _23283_ (.Y(_05637_),
    .A(_05634_),
    .B(_05635_));
 sg13g2_nor3_1 _23284_ (.A(_05565_),
    .B(_05636_),
    .C(_05637_),
    .Y(_05638_));
 sg13g2_a21oi_1 _23285_ (.A1(_05634_),
    .A2(_05635_),
    .Y(_05639_),
    .B1(_05638_));
 sg13g2_nor2_1 _23286_ (.A(_05565_),
    .B(_05632_),
    .Y(_05640_));
 sg13g2_a21oi_1 _23287_ (.A1(_05533_),
    .A2(_05534_),
    .Y(_05641_),
    .B1(_05523_));
 sg13g2_or2_1 _23288_ (.X(_05642_),
    .B(_05641_),
    .A(_05535_));
 sg13g2_nor2_1 _23289_ (.A(_05572_),
    .B(_05642_),
    .Y(_05643_));
 sg13g2_nor2_1 _23290_ (.A(net5401),
    .B(net5321),
    .Y(_05644_));
 sg13g2_nor3_1 _23291_ (.A(net5401),
    .B(_05631_),
    .C(net5321),
    .Y(_05645_));
 sg13g2_o21ai_1 _23292_ (.B1(_05631_),
    .Y(_05646_),
    .A1(net5401),
    .A2(net5321));
 sg13g2_nor2b_1 _23293_ (.A(_05645_),
    .B_N(_05646_),
    .Y(_05647_));
 sg13g2_xnor2_1 _23294_ (.Y(_05648_),
    .A(_05640_),
    .B(_05647_));
 sg13g2_nor2_1 _23295_ (.A(_05639_),
    .B(_05648_),
    .Y(_05649_));
 sg13g2_nand2b_1 _23296_ (.Y(_05650_),
    .B(net5454),
    .A_N(_05636_));
 sg13g2_nor2_1 _23297_ (.A(_05555_),
    .B(_05636_),
    .Y(_05651_));
 sg13g2_nand2_1 _23298_ (.Y(_05652_),
    .A(_07954_),
    .B(_05651_));
 sg13g2_inv_1 _23299_ (.Y(_05653_),
    .A(_05652_));
 sg13g2_o21ai_1 _23300_ (.B1(_05650_),
    .Y(_05654_),
    .A1(net5582),
    .A2(_05555_));
 sg13g2_and2_1 _23301_ (.A(_05652_),
    .B(_05654_),
    .X(_05655_));
 sg13g2_xor2_1 _23302_ (.B(_05648_),
    .A(_05639_),
    .X(_05656_));
 sg13g2_a21oi_1 _23303_ (.A1(_05655_),
    .A2(_05656_),
    .Y(_05657_),
    .B1(_05649_));
 sg13g2_nor2_1 _23304_ (.A(net5453),
    .B(_05632_),
    .Y(_05658_));
 sg13g2_nor2_1 _23305_ (.A(_05555_),
    .B(_05632_),
    .Y(_05659_));
 sg13g2_nand2b_1 _23306_ (.Y(_05660_),
    .B(_05651_),
    .A_N(_05632_));
 sg13g2_o21ai_1 _23307_ (.B1(_05660_),
    .Y(_05661_),
    .A1(_05651_),
    .A2(_05658_));
 sg13g2_a21o_1 _23308_ (.A2(_05646_),
    .A1(_05640_),
    .B1(_05645_),
    .X(_05662_));
 sg13g2_nor2_1 _23309_ (.A(_05565_),
    .B(_05629_),
    .Y(_05663_));
 sg13g2_nor2_1 _23310_ (.A(_05572_),
    .B(_05609_),
    .Y(_05664_));
 sg13g2_nor2_1 _23311_ (.A(net5401),
    .B(_05609_),
    .Y(_05665_));
 sg13g2_xor2_1 _23312_ (.B(_05665_),
    .A(_05643_),
    .X(_05666_));
 sg13g2_xnor2_1 _23313_ (.Y(_05667_),
    .A(_05663_),
    .B(_05666_));
 sg13g2_nand2b_1 _23314_ (.Y(_05668_),
    .B(_05662_),
    .A_N(_05667_));
 sg13g2_xor2_1 _23315_ (.B(_05667_),
    .A(_05662_),
    .X(_05669_));
 sg13g2_xor2_1 _23316_ (.B(_05669_),
    .A(_05661_),
    .X(_05670_));
 sg13g2_nor2b_1 _23317_ (.A(_05657_),
    .B_N(_05670_),
    .Y(_05671_));
 sg13g2_xnor2_1 _23318_ (.Y(_05672_),
    .A(_05657_),
    .B(_05670_));
 sg13g2_a21oi_1 _23319_ (.A1(_05653_),
    .A2(_05672_),
    .Y(_05673_),
    .B1(_05671_));
 sg13g2_o21ai_1 _23320_ (.B1(_05668_),
    .Y(_05674_),
    .A1(_05661_),
    .A2(_05669_));
 sg13g2_nand2_1 _23321_ (.Y(_05675_),
    .A(_05554_),
    .B(_05630_));
 sg13g2_nor2_1 _23322_ (.A(_05632_),
    .B(_05675_),
    .Y(_05676_));
 sg13g2_a21oi_1 _23323_ (.A1(net5454),
    .A2(_05630_),
    .Y(_05677_),
    .B1(_05659_));
 sg13g2_or2_1 _23324_ (.X(_05678_),
    .B(_05677_),
    .A(_05676_));
 sg13g2_inv_1 _23325_ (.Y(_05679_),
    .A(_05678_));
 sg13g2_a22oi_1 _23326_ (.Y(_05680_),
    .B1(_05666_),
    .B2(_05663_),
    .A2(_05664_),
    .A1(_05644_));
 sg13g2_nor2_1 _23327_ (.A(_05565_),
    .B(net5321),
    .Y(_05681_));
 sg13g2_nand2_1 _23328_ (.Y(_05682_),
    .A(_05573_),
    .B(_05580_));
 sg13g2_nor3_2 _23329_ (.A(_05542_),
    .B(net5401),
    .C(_05579_),
    .Y(_05683_));
 sg13g2_xor2_1 _23330_ (.B(_05683_),
    .A(_05664_),
    .X(_05684_));
 sg13g2_and2_1 _23331_ (.A(_05681_),
    .B(_05684_),
    .X(_05685_));
 sg13g2_xnor2_1 _23332_ (.Y(_05686_),
    .A(_05681_),
    .B(_05684_));
 sg13g2_nor2_1 _23333_ (.A(_05680_),
    .B(_05686_),
    .Y(_05687_));
 sg13g2_xor2_1 _23334_ (.B(_05686_),
    .A(_05680_),
    .X(_05688_));
 sg13g2_xnor2_1 _23335_ (.Y(_05689_),
    .A(_05678_),
    .B(_05688_));
 sg13g2_xnor2_1 _23336_ (.Y(_05690_),
    .A(_05674_),
    .B(_05689_));
 sg13g2_nor2_1 _23337_ (.A(_05660_),
    .B(_05690_),
    .Y(_05691_));
 sg13g2_xnor2_1 _23338_ (.Y(_05692_),
    .A(_05660_),
    .B(_05690_));
 sg13g2_nor2_1 _23339_ (.A(_05673_),
    .B(_05692_),
    .Y(_05693_));
 sg13g2_nor2_1 _23340_ (.A(_08098_),
    .B(net5453),
    .Y(_05694_));
 sg13g2_nand2_1 _23341_ (.Y(_05695_),
    .A(_00107_),
    .B(net5454));
 sg13g2_nor2_1 _23342_ (.A(net5481),
    .B(_05695_),
    .Y(_05696_));
 sg13g2_xor2_1 _23343_ (.B(_05692_),
    .A(_05673_),
    .X(_05697_));
 sg13g2_a21oi_1 _23344_ (.A1(_05696_),
    .A2(_05697_),
    .Y(_05698_),
    .B1(_05693_));
 sg13g2_nor2_1 _23345_ (.A(net5481),
    .B(_05650_),
    .Y(_05699_));
 sg13g2_a21oi_1 _23346_ (.A1(_05674_),
    .A2(_05689_),
    .Y(_05700_),
    .B1(_05691_));
 sg13g2_a21oi_1 _23347_ (.A1(_05679_),
    .A2(_05688_),
    .Y(_05701_),
    .B1(_05687_));
 sg13g2_or2_1 _23348_ (.X(_05702_),
    .B(net5321),
    .A(net5453));
 sg13g2_nor2_1 _23349_ (.A(_05555_),
    .B(net5321),
    .Y(_05703_));
 sg13g2_nor2_1 _23350_ (.A(net5321),
    .B(_05675_),
    .Y(_05704_));
 sg13g2_a21oi_1 _23351_ (.A1(_05675_),
    .A2(_05702_),
    .Y(_05705_),
    .B1(_05704_));
 sg13g2_a21oi_1 _23352_ (.A1(_05664_),
    .A2(_05683_),
    .Y(_05706_),
    .B1(_05685_));
 sg13g2_nand2b_1 _23353_ (.Y(_05707_),
    .B(_05566_),
    .A_N(_05609_));
 sg13g2_nand2_1 _23354_ (.Y(_05708_),
    .A(_05602_),
    .B(_05683_));
 sg13g2_xor2_1 _23355_ (.B(_05682_),
    .A(_05600_),
    .X(_05709_));
 sg13g2_xor2_1 _23356_ (.B(_05709_),
    .A(_05707_),
    .X(_05710_));
 sg13g2_nor2b_1 _23357_ (.A(_05706_),
    .B_N(_05710_),
    .Y(_05711_));
 sg13g2_xnor2_1 _23358_ (.Y(_05712_),
    .A(_05706_),
    .B(_05710_));
 sg13g2_xnor2_1 _23359_ (.Y(_05713_),
    .A(_05705_),
    .B(_05712_));
 sg13g2_nor2_1 _23360_ (.A(_05701_),
    .B(_05713_),
    .Y(_05714_));
 sg13g2_xor2_1 _23361_ (.B(_05713_),
    .A(_05701_),
    .X(_05715_));
 sg13g2_xnor2_1 _23362_ (.Y(_05716_),
    .A(_05676_),
    .B(_05715_));
 sg13g2_nor2_1 _23363_ (.A(_05700_),
    .B(_05716_),
    .Y(_05717_));
 sg13g2_xor2_1 _23364_ (.B(_05716_),
    .A(_05700_),
    .X(_05718_));
 sg13g2_xnor2_1 _23365_ (.Y(_05719_),
    .A(_05699_),
    .B(_05718_));
 sg13g2_nor2_1 _23366_ (.A(_05698_),
    .B(_05719_),
    .Y(_05720_));
 sg13g2_xnor2_1 _23367_ (.Y(_05721_),
    .A(_05655_),
    .B(_05656_));
 sg13g2_nor2_1 _23368_ (.A(net5401),
    .B(_05636_),
    .Y(_05722_));
 sg13g2_nor2_1 _23369_ (.A(_05572_),
    .B(_05636_),
    .Y(_05723_));
 sg13g2_nor2_1 _23370_ (.A(_08098_),
    .B(_05565_),
    .Y(_05724_));
 sg13g2_xor2_1 _23371_ (.B(_05723_),
    .A(_05633_),
    .X(_05725_));
 sg13g2_a22oi_1 _23372_ (.Y(_05726_),
    .B1(_05724_),
    .B2(_05725_),
    .A2(_05722_),
    .A1(_05635_));
 sg13g2_o21ai_1 _23373_ (.B1(_05637_),
    .Y(_05727_),
    .A1(_05565_),
    .A2(_05636_));
 sg13g2_nand2b_1 _23374_ (.Y(_05728_),
    .B(_05727_),
    .A_N(_05638_));
 sg13g2_nor2_1 _23375_ (.A(_05726_),
    .B(_05728_),
    .Y(_05729_));
 sg13g2_xor2_1 _23376_ (.B(_05728_),
    .A(_05726_),
    .X(_05730_));
 sg13g2_a21oi_1 _23377_ (.A1(_05694_),
    .A2(_05730_),
    .Y(_05731_),
    .B1(_05729_));
 sg13g2_nor2_1 _23378_ (.A(_05721_),
    .B(_05731_),
    .Y(_05732_));
 sg13g2_xnor2_1 _23379_ (.Y(_05733_),
    .A(_05652_),
    .B(_05672_));
 sg13g2_nand2_1 _23380_ (.Y(_05734_),
    .A(_05732_),
    .B(_05733_));
 sg13g2_xnor2_1 _23381_ (.Y(_05735_),
    .A(_05696_),
    .B(_05697_));
 sg13g2_nor2_1 _23382_ (.A(_05734_),
    .B(_05735_),
    .Y(_05736_));
 sg13g2_nor4_2 _23383_ (.A(_08098_),
    .B(_05514_),
    .C(net5453),
    .Y(_05737_),
    .D(_05563_));
 sg13g2_xor2_1 _23384_ (.B(_05725_),
    .A(_05724_),
    .X(_05738_));
 sg13g2_nand2_1 _23385_ (.Y(_05739_),
    .A(_05737_),
    .B(_05738_));
 sg13g2_xnor2_1 _23386_ (.Y(_05740_),
    .A(_05695_),
    .B(_05730_));
 sg13g2_nand2b_1 _23387_ (.Y(_05741_),
    .B(_05740_),
    .A_N(_05739_));
 sg13g2_xnor2_1 _23388_ (.Y(_05742_),
    .A(_05721_),
    .B(_05731_));
 sg13g2_nor2_1 _23389_ (.A(_05741_),
    .B(_05742_),
    .Y(_05743_));
 sg13g2_nand2_1 _23390_ (.Y(_05744_),
    .A(_05733_),
    .B(_05743_));
 sg13g2_inv_1 _23391_ (.Y(_05745_),
    .A(_05744_));
 sg13g2_xor2_1 _23392_ (.B(_05735_),
    .A(_05734_),
    .X(_05746_));
 sg13g2_a21o_1 _23393_ (.A2(_05746_),
    .A1(_05745_),
    .B1(_05736_),
    .X(_05747_));
 sg13g2_xor2_1 _23394_ (.B(_05719_),
    .A(_05698_),
    .X(_05748_));
 sg13g2_a21oi_2 _23395_ (.B1(_05720_),
    .Y(_05749_),
    .A2(_05748_),
    .A1(_05747_));
 sg13g2_nor3_1 _23396_ (.A(net5453),
    .B(net5481),
    .C(_05632_),
    .Y(_05750_));
 sg13g2_a21oi_1 _23397_ (.A1(_05676_),
    .A2(_05715_),
    .Y(_05751_),
    .B1(_05714_));
 sg13g2_a21oi_1 _23398_ (.A1(_05705_),
    .A2(_05712_),
    .Y(_05752_),
    .B1(_05711_));
 sg13g2_or2_1 _23399_ (.X(_05753_),
    .B(net5321),
    .A(_05611_));
 sg13g2_o21ai_1 _23400_ (.B1(_05753_),
    .Y(_05754_),
    .A1(_05610_),
    .A2(_05703_));
 sg13g2_o21ai_1 _23401_ (.B1(_05708_),
    .Y(_05755_),
    .A1(_05707_),
    .A2(_05709_));
 sg13g2_xnor2_1 _23402_ (.Y(_05756_),
    .A(_05604_),
    .B(_05605_));
 sg13g2_nand2b_1 _23403_ (.Y(_05757_),
    .B(_05755_),
    .A_N(_05756_));
 sg13g2_xor2_1 _23404_ (.B(_05756_),
    .A(_05755_),
    .X(_05758_));
 sg13g2_xor2_1 _23405_ (.B(_05758_),
    .A(_05754_),
    .X(_05759_));
 sg13g2_nor2b_1 _23406_ (.A(_05752_),
    .B_N(_05759_),
    .Y(_05760_));
 sg13g2_xnor2_1 _23407_ (.Y(_05761_),
    .A(_05752_),
    .B(_05759_));
 sg13g2_xnor2_1 _23408_ (.Y(_05762_),
    .A(_05704_),
    .B(_05761_));
 sg13g2_nor2_1 _23409_ (.A(_05751_),
    .B(_05762_),
    .Y(_05763_));
 sg13g2_xor2_1 _23410_ (.B(_05762_),
    .A(_05751_),
    .X(_05764_));
 sg13g2_xnor2_1 _23411_ (.Y(_05765_),
    .A(_05750_),
    .B(_05764_));
 sg13g2_a21oi_1 _23412_ (.A1(_05699_),
    .A2(_05718_),
    .Y(_05766_),
    .B1(_05717_));
 sg13g2_or2_1 _23413_ (.X(_05767_),
    .B(_05766_),
    .A(_05765_));
 sg13g2_xnor2_1 _23414_ (.Y(_05768_),
    .A(_05765_),
    .B(_05766_));
 sg13g2_a21oi_1 _23415_ (.A1(_05750_),
    .A2(_05764_),
    .Y(_05769_),
    .B1(_05763_));
 sg13g2_nor3_2 _23416_ (.A(net5453),
    .B(net5481),
    .C(_05629_),
    .Y(_05770_));
 sg13g2_a21oi_1 _23417_ (.A1(_05704_),
    .A2(_05761_),
    .Y(_05771_),
    .B1(_05760_));
 sg13g2_o21ai_1 _23418_ (.B1(_05757_),
    .Y(_05772_),
    .A1(_05754_),
    .A2(_05758_));
 sg13g2_xnor2_1 _23419_ (.Y(_05773_),
    .A(_05613_),
    .B(_05614_));
 sg13g2_nand2b_1 _23420_ (.Y(_05774_),
    .B(_05772_),
    .A_N(_05773_));
 sg13g2_xor2_1 _23421_ (.B(_05773_),
    .A(_05772_),
    .X(_05775_));
 sg13g2_xnor2_1 _23422_ (.Y(_05776_),
    .A(_05753_),
    .B(_05775_));
 sg13g2_nor2_1 _23423_ (.A(_05771_),
    .B(_05776_),
    .Y(_05777_));
 sg13g2_xor2_1 _23424_ (.B(_05776_),
    .A(_05771_),
    .X(_05778_));
 sg13g2_xnor2_1 _23425_ (.Y(_05779_),
    .A(_05770_),
    .B(_05778_));
 sg13g2_nand2_1 _23426_ (.Y(_05780_),
    .A(_05769_),
    .B(_05779_));
 sg13g2_or2_1 _23427_ (.X(_05781_),
    .B(_05779_),
    .A(_05769_));
 sg13g2_nand2_1 _23428_ (.Y(_05782_),
    .A(_05780_),
    .B(_05781_));
 sg13g2_nor3_2 _23429_ (.A(_05749_),
    .B(_05768_),
    .C(_05782_),
    .Y(_05783_));
 sg13g2_nand2b_1 _23430_ (.Y(_05784_),
    .B(_05780_),
    .A_N(_05767_));
 sg13g2_nand2_1 _23431_ (.Y(_05785_),
    .A(_05781_),
    .B(_05784_));
 sg13g2_nor2_1 _23432_ (.A(_05783_),
    .B(_05785_),
    .Y(_05786_));
 sg13g2_nor2_1 _23433_ (.A(net5481),
    .B(_05702_),
    .Y(_05787_));
 sg13g2_o21ai_1 _23434_ (.B1(_05774_),
    .Y(_05788_),
    .A1(_05753_),
    .A2(_05775_));
 sg13g2_xor2_1 _23435_ (.B(_05618_),
    .A(_05612_),
    .X(_05789_));
 sg13g2_nor2b_1 _23436_ (.A(_05789_),
    .B_N(_05788_),
    .Y(_05790_));
 sg13g2_xor2_1 _23437_ (.B(_05789_),
    .A(_05788_),
    .X(_05791_));
 sg13g2_nor3_1 _23438_ (.A(net5481),
    .B(_05702_),
    .C(_05791_),
    .Y(_05792_));
 sg13g2_xor2_1 _23439_ (.B(_05791_),
    .A(_05787_),
    .X(_05793_));
 sg13g2_a21oi_1 _23440_ (.A1(_05770_),
    .A2(_05778_),
    .Y(_05794_),
    .B1(_05777_));
 sg13g2_nor2_1 _23441_ (.A(_05793_),
    .B(_05794_),
    .Y(_05795_));
 sg13g2_inv_1 _23442_ (.Y(_05796_),
    .A(_05795_));
 sg13g2_xnor2_1 _23443_ (.Y(_05797_),
    .A(_05793_),
    .B(_05794_));
 sg13g2_inv_1 _23444_ (.Y(_05798_),
    .A(_05797_));
 sg13g2_nor2_1 _23445_ (.A(_05790_),
    .B(_05792_),
    .Y(_05799_));
 sg13g2_xnor2_1 _23446_ (.Y(_05800_),
    .A(_05623_),
    .B(_05624_));
 sg13g2_or2_1 _23447_ (.X(_05801_),
    .B(_05800_),
    .A(_05799_));
 sg13g2_inv_1 _23448_ (.Y(_05802_),
    .A(_05801_));
 sg13g2_nand2_1 _23449_ (.Y(_05803_),
    .A(_05799_),
    .B(_05800_));
 sg13g2_xor2_1 _23450_ (.B(_05800_),
    .A(_05799_),
    .X(_05804_));
 sg13g2_and2_1 _23451_ (.A(_05798_),
    .B(_05804_),
    .X(_05805_));
 sg13g2_o21ai_1 _23452_ (.B1(_05805_),
    .Y(_05806_),
    .A1(_05783_),
    .A2(_05785_));
 sg13g2_a21oi_1 _23453_ (.A1(_05795_),
    .A2(_05803_),
    .Y(_05807_),
    .B1(_05802_));
 sg13g2_xor2_1 _23454_ (.B(_05626_),
    .A(_05625_),
    .X(_05808_));
 sg13g2_inv_1 _23455_ (.Y(_05809_),
    .A(_05808_));
 sg13g2_a21oi_1 _23456_ (.A1(_05806_),
    .A2(_05807_),
    .Y(_05810_),
    .B1(_05809_));
 sg13g2_o21ai_1 _23457_ (.B1(_05598_),
    .Y(_05811_),
    .A1(_05627_),
    .A2(_05810_));
 sg13g2_nand2_2 _23458_ (.Y(_05812_),
    .A(_05597_),
    .B(_05811_));
 sg13g2_a21oi_1 _23459_ (.A1(_05554_),
    .A2(_05560_),
    .Y(_05813_),
    .B1(_05563_));
 sg13g2_nor3_2 _23460_ (.A(_05556_),
    .B(_05595_),
    .C(_05813_),
    .Y(_05814_));
 sg13g2_xor2_1 _23461_ (.B(_05814_),
    .A(_05812_),
    .X(_05815_));
 sg13g2_xnor2_1 _23462_ (.Y(_05816_),
    .A(_05812_),
    .B(_05814_));
 sg13g2_nand2_1 _23463_ (.Y(_05817_),
    .A(_00122_),
    .B(_05815_));
 sg13g2_or3_1 _23464_ (.A(_05598_),
    .B(_05627_),
    .C(_05810_),
    .X(_05818_));
 sg13g2_and2_2 _23465_ (.A(_05811_),
    .B(_05818_),
    .X(_05819_));
 sg13g2_xor2_1 _23466_ (.B(_05819_),
    .A(_00121_),
    .X(_05820_));
 sg13g2_nand3_1 _23467_ (.B(_05807_),
    .C(_05809_),
    .A(_05806_),
    .Y(_05821_));
 sg13g2_nand2b_2 _23468_ (.Y(_05822_),
    .B(_05821_),
    .A_N(_05810_));
 sg13g2_nor2b_1 _23469_ (.A(_00120_),
    .B_N(_05822_),
    .Y(_05823_));
 sg13g2_xnor2_1 _23470_ (.Y(_05824_),
    .A(_00120_),
    .B(_05822_));
 sg13g2_nand2_1 _23471_ (.Y(_05825_),
    .A(_05820_),
    .B(_05824_));
 sg13g2_o21ai_1 _23472_ (.B1(_05798_),
    .Y(_05826_),
    .A1(_05783_),
    .A2(_05785_));
 sg13g2_a21o_1 _23473_ (.A2(_05826_),
    .A1(_05796_),
    .B1(_05804_),
    .X(_05827_));
 sg13g2_nand3_1 _23474_ (.B(_05804_),
    .C(_05826_),
    .A(_05796_),
    .Y(_05828_));
 sg13g2_nand2_1 _23475_ (.Y(_05829_),
    .A(_05827_),
    .B(_05828_));
 sg13g2_a21o_1 _23476_ (.A2(_05828_),
    .A1(_05827_),
    .B1(_08102_),
    .X(_05830_));
 sg13g2_nand3_1 _23477_ (.B(_05827_),
    .C(_05828_),
    .A(_08102_),
    .Y(_05831_));
 sg13g2_xnor2_1 _23478_ (.Y(_05832_),
    .A(_05786_),
    .B(_05797_));
 sg13g2_xnor2_1 _23479_ (.Y(_05833_),
    .A(_00118_),
    .B(_05832_));
 sg13g2_and3_1 _23480_ (.X(_05834_),
    .A(_05830_),
    .B(_05831_),
    .C(_05833_));
 sg13g2_o21ai_1 _23481_ (.B1(_05767_),
    .Y(_05835_),
    .A1(_05749_),
    .A2(_05768_));
 sg13g2_xnor2_1 _23482_ (.Y(_05836_),
    .A(_05782_),
    .B(_05835_));
 sg13g2_nand2b_1 _23483_ (.Y(_05837_),
    .B(\atari2600.tia.audio_left_counter[10] ),
    .A_N(_05836_));
 sg13g2_xnor2_1 _23484_ (.Y(_05838_),
    .A(_00117_),
    .B(_05836_));
 sg13g2_inv_1 _23485_ (.Y(_05839_),
    .A(_05838_));
 sg13g2_xor2_1 _23486_ (.B(_05768_),
    .A(_05749_),
    .X(_05840_));
 sg13g2_and2_1 _23487_ (.A(_00116_),
    .B(_05840_),
    .X(_05841_));
 sg13g2_nand2_1 _23488_ (.Y(_05842_),
    .A(_00116_),
    .B(_05840_));
 sg13g2_xnor2_1 _23489_ (.Y(_05843_),
    .A(_05744_),
    .B(_05746_));
 sg13g2_and2_1 _23490_ (.A(_00114_),
    .B(_05843_),
    .X(_05844_));
 sg13g2_xor2_1 _23491_ (.B(_05748_),
    .A(_05747_),
    .X(_05845_));
 sg13g2_xnor2_1 _23492_ (.Y(_05846_),
    .A(_00115_),
    .B(_05845_));
 sg13g2_or2_1 _23493_ (.X(_05847_),
    .B(_05846_),
    .A(_05844_));
 sg13g2_nor2_1 _23494_ (.A(_00114_),
    .B(_05843_),
    .Y(_05848_));
 sg13g2_nor2_1 _23495_ (.A(_05732_),
    .B(_05743_),
    .Y(_05849_));
 sg13g2_xnor2_1 _23496_ (.Y(_05850_),
    .A(_05733_),
    .B(_05849_));
 sg13g2_nor2b_1 _23497_ (.A(_05850_),
    .B_N(\atari2600.tia.audio_left_counter[6] ),
    .Y(_05851_));
 sg13g2_xnor2_1 _23498_ (.Y(_05852_),
    .A(_00113_),
    .B(_05850_));
 sg13g2_xor2_1 _23499_ (.B(_05742_),
    .A(_05741_),
    .X(_05853_));
 sg13g2_or2_1 _23500_ (.X(_05854_),
    .B(_05853_),
    .A(_00111_));
 sg13g2_nand2_1 _23501_ (.Y(_05855_),
    .A(_00111_),
    .B(_05853_));
 sg13g2_xor2_1 _23502_ (.B(_05740_),
    .A(_05739_),
    .X(_05856_));
 sg13g2_nand2_1 _23503_ (.Y(_05857_),
    .A(\atari2600.tia.audio_left_counter[4] ),
    .B(_05856_));
 sg13g2_xor2_1 _23504_ (.B(_05856_),
    .A(_00110_),
    .X(_05858_));
 sg13g2_xor2_1 _23505_ (.B(_05738_),
    .A(_05737_),
    .X(_05859_));
 sg13g2_or2_1 _23506_ (.X(_05860_),
    .B(_05859_),
    .A(_00109_));
 sg13g2_nand2_1 _23507_ (.Y(_05861_),
    .A(_00109_),
    .B(_05859_));
 sg13g2_nand2_2 _23508_ (.Y(_05862_),
    .A(_00107_),
    .B(_05571_));
 sg13g2_nor2_1 _23509_ (.A(\atari2600.tia.audio_left_counter[1] ),
    .B(_05862_),
    .Y(_05863_));
 sg13g2_a21oi_1 _23510_ (.A1(_00107_),
    .A2(_05573_),
    .Y(_05864_),
    .B1(_05722_));
 sg13g2_nor2_2 _23511_ (.A(_05737_),
    .B(_05864_),
    .Y(_05865_));
 sg13g2_xnor2_1 _23512_ (.Y(_05866_),
    .A(_00108_),
    .B(_05865_));
 sg13g2_nor2_1 _23513_ (.A(_05863_),
    .B(_05866_),
    .Y(_05867_));
 sg13g2_o21ai_1 _23514_ (.B1(_05860_),
    .Y(_05868_),
    .A1(_08033_),
    .A2(_05865_));
 sg13g2_o21ai_1 _23515_ (.B1(_05861_),
    .Y(_05869_),
    .A1(_05867_),
    .A2(_05868_));
 sg13g2_o21ai_1 _23516_ (.B1(_05857_),
    .Y(_05870_),
    .A1(_05858_),
    .A2(_05869_));
 sg13g2_nand2_1 _23517_ (.Y(_05871_),
    .A(_05855_),
    .B(_05870_));
 sg13g2_a21oi_1 _23518_ (.A1(_05854_),
    .A2(_05871_),
    .Y(_05872_),
    .B1(_05852_));
 sg13g2_nor3_1 _23519_ (.A(_05848_),
    .B(_05851_),
    .C(_05872_),
    .Y(_05873_));
 sg13g2_nor3_1 _23520_ (.A(_05844_),
    .B(_05846_),
    .C(_05873_),
    .Y(_05874_));
 sg13g2_nor2_1 _23521_ (.A(_00116_),
    .B(_05840_),
    .Y(_05875_));
 sg13g2_nand2b_1 _23522_ (.Y(_05876_),
    .B(\atari2600.tia.audio_left_counter[8] ),
    .A_N(_05845_));
 sg13g2_o21ai_1 _23523_ (.B1(_05876_),
    .Y(_05877_),
    .A1(_00116_),
    .A2(_05840_));
 sg13g2_o21ai_1 _23524_ (.B1(_05842_),
    .Y(_05878_),
    .A1(_05874_),
    .A2(_05877_));
 sg13g2_o21ai_1 _23525_ (.B1(_05837_),
    .Y(_05879_),
    .A1(_05838_),
    .A2(_05878_));
 sg13g2_nand4_1 _23526_ (.B(_05831_),
    .C(_05833_),
    .A(_05830_),
    .Y(_05880_),
    .D(_05879_));
 sg13g2_nand4_1 _23527_ (.B(_05830_),
    .C(_05831_),
    .A(_08101_),
    .Y(_05881_),
    .D(_05832_));
 sg13g2_nand3_1 _23528_ (.B(_05827_),
    .C(_05828_),
    .A(\atari2600.tia.audio_left_counter[12] ),
    .Y(_05882_));
 sg13g2_nand3_1 _23529_ (.B(_05881_),
    .C(_05882_),
    .A(_05880_),
    .Y(_05883_));
 sg13g2_nand3_1 _23530_ (.B(_05824_),
    .C(_05883_),
    .A(_05820_),
    .Y(_05884_));
 sg13g2_nor2_1 _23531_ (.A(_00122_),
    .B(_05815_),
    .Y(_05885_));
 sg13g2_nor2b_1 _23532_ (.A(_05819_),
    .B_N(\atari2600.tia.audio_left_counter[14] ),
    .Y(_05886_));
 sg13g2_a221oi_1 _23533_ (.B2(_05823_),
    .C1(_05886_),
    .B1(_05820_),
    .A1(_08103_),
    .Y(_05887_),
    .A2(_05816_));
 sg13g2_a22oi_1 _23534_ (.Y(_05888_),
    .B1(_05884_),
    .B2(_05887_),
    .A2(_05815_),
    .A1(_00122_));
 sg13g2_nor3_1 _23535_ (.A(\atari2600.tia.audio_left_counter[0] ),
    .B(_05502_),
    .C(_05888_),
    .Y(_05889_));
 sg13g2_a21oi_1 _23536_ (.A1(net3464),
    .A2(_05502_),
    .Y(_05890_),
    .B1(_05889_));
 sg13g2_o21ai_1 _23537_ (.B1(_05496_),
    .Y(_02012_),
    .A1(net5306),
    .A2(net3465));
 sg13g2_nand2_1 _23538_ (.Y(_05891_),
    .A(net7021),
    .B(net5280));
 sg13g2_nand2b_1 _23539_ (.Y(_05892_),
    .B(_05888_),
    .A_N(_05502_));
 sg13g2_nand2_1 _23540_ (.Y(_05893_),
    .A(\atari2600.tia.audio_left_counter[1] ),
    .B(\atari2600.tia.audio_left_counter[0] ));
 sg13g2_or2_1 _23541_ (.X(_05894_),
    .B(\atari2600.tia.audio_left_counter[0] ),
    .A(net7021));
 sg13g2_nand3_1 _23542_ (.B(_05893_),
    .C(_05894_),
    .A(net4552),
    .Y(_05895_));
 sg13g2_o21ai_1 _23543_ (.B1(_05891_),
    .Y(_02013_),
    .A1(net5306),
    .A2(_05895_));
 sg13g2_nand2_1 _23544_ (.Y(_05896_),
    .A(net3933),
    .B(net5279));
 sg13g2_nor2_1 _23545_ (.A(_00108_),
    .B(_05893_),
    .Y(_05897_));
 sg13g2_xor2_1 _23546_ (.B(_05893_),
    .A(_00108_),
    .X(_05898_));
 sg13g2_nand3_1 _23547_ (.B(net4552),
    .C(_05898_),
    .A(net5344),
    .Y(_05899_));
 sg13g2_nand2_1 _23548_ (.Y(_02014_),
    .A(_05896_),
    .B(_05899_));
 sg13g2_xor2_1 _23549_ (.B(_05897_),
    .A(_00109_),
    .X(_05900_));
 sg13g2_nor2_1 _23550_ (.A(net5306),
    .B(_05900_),
    .Y(_05901_));
 sg13g2_a22oi_1 _23551_ (.Y(_05902_),
    .B1(net4552),
    .B2(_05901_),
    .A2(net5278),
    .A1(net3411));
 sg13g2_inv_1 _23552_ (.Y(_02015_),
    .A(net3412));
 sg13g2_nand2_1 _23553_ (.Y(_05903_),
    .A(net3133),
    .B(net5278));
 sg13g2_nand4_1 _23554_ (.B(\atari2600.tia.audio_left_counter[2] ),
    .C(\atari2600.tia.audio_left_counter[1] ),
    .A(\atari2600.tia.audio_left_counter[3] ),
    .Y(_05904_),
    .D(\atari2600.tia.audio_left_counter[0] ));
 sg13g2_nor2_1 _23555_ (.A(_00110_),
    .B(_05904_),
    .Y(_05905_));
 sg13g2_xor2_1 _23556_ (.B(_05904_),
    .A(_00110_),
    .X(_05906_));
 sg13g2_nand3_1 _23557_ (.B(net4552),
    .C(_05906_),
    .A(net5343),
    .Y(_05907_));
 sg13g2_nand2_1 _23558_ (.Y(_02016_),
    .A(_05903_),
    .B(_05907_));
 sg13g2_xor2_1 _23559_ (.B(_05905_),
    .A(_00111_),
    .X(_05908_));
 sg13g2_nor2_1 _23560_ (.A(net5306),
    .B(_05908_),
    .Y(_05909_));
 sg13g2_a22oi_1 _23561_ (.Y(_05910_),
    .B1(net4552),
    .B2(_05909_),
    .A2(net5278),
    .A1(net3473));
 sg13g2_inv_1 _23562_ (.Y(_02017_),
    .A(net3474));
 sg13g2_nand2_1 _23563_ (.Y(_05911_),
    .A(net3992),
    .B(net5278));
 sg13g2_nand2_1 _23564_ (.Y(_05912_),
    .A(\atari2600.tia.audio_left_counter[5] ),
    .B(\atari2600.tia.audio_left_counter[4] ));
 sg13g2_nor2_2 _23565_ (.A(_05904_),
    .B(_05912_),
    .Y(_05913_));
 sg13g2_nor3_1 _23566_ (.A(_00113_),
    .B(_05904_),
    .C(_05912_),
    .Y(_05914_));
 sg13g2_xnor2_1 _23567_ (.Y(_05915_),
    .A(_00113_),
    .B(_05913_));
 sg13g2_nand3_1 _23568_ (.B(net4552),
    .C(_05915_),
    .A(net5343),
    .Y(_05916_));
 sg13g2_nand2_1 _23569_ (.Y(_02018_),
    .A(_05911_),
    .B(_05916_));
 sg13g2_xor2_1 _23570_ (.B(_05914_),
    .A(_00114_),
    .X(_05917_));
 sg13g2_nor2_1 _23571_ (.A(net5303),
    .B(_05917_),
    .Y(_05918_));
 sg13g2_a22oi_1 _23572_ (.Y(_05919_),
    .B1(net4552),
    .B2(_05918_),
    .A2(net5278),
    .A1(net3069));
 sg13g2_inv_1 _23573_ (.Y(_02019_),
    .A(net3070));
 sg13g2_nand2_1 _23574_ (.Y(_05920_),
    .A(net3145),
    .B(net5277));
 sg13g2_and2_1 _23575_ (.A(\atari2600.tia.audio_left_counter[7] ),
    .B(\atari2600.tia.audio_left_counter[6] ),
    .X(_05921_));
 sg13g2_nand2_1 _23576_ (.Y(_05922_),
    .A(_05913_),
    .B(_05921_));
 sg13g2_nor2_1 _23577_ (.A(_00115_),
    .B(_05922_),
    .Y(_05923_));
 sg13g2_xor2_1 _23578_ (.B(_05922_),
    .A(_00115_),
    .X(_05924_));
 sg13g2_nand3_1 _23579_ (.B(net4552),
    .C(_05924_),
    .A(net5343),
    .Y(_05925_));
 sg13g2_nand2_1 _23580_ (.Y(_02020_),
    .A(_05920_),
    .B(_05925_));
 sg13g2_xor2_1 _23581_ (.B(_05923_),
    .A(_00116_),
    .X(_05926_));
 sg13g2_nor2_1 _23582_ (.A(net5303),
    .B(_05926_),
    .Y(_05927_));
 sg13g2_a22oi_1 _23583_ (.Y(_05928_),
    .B1(net4553),
    .B2(_05927_),
    .A2(net5276),
    .A1(net3905));
 sg13g2_inv_1 _23584_ (.Y(_02021_),
    .A(net3906));
 sg13g2_nand2_1 _23585_ (.Y(_05929_),
    .A(net3805),
    .B(net5276));
 sg13g2_nand4_1 _23586_ (.B(net3145),
    .C(_05913_),
    .A(\atari2600.tia.audio_left_counter[9] ),
    .Y(_05930_),
    .D(_05921_));
 sg13g2_inv_1 _23587_ (.Y(_05931_),
    .A(_05930_));
 sg13g2_nor2_1 _23588_ (.A(_00117_),
    .B(_05930_),
    .Y(_05932_));
 sg13g2_xor2_1 _23589_ (.B(_05930_),
    .A(_00117_),
    .X(_05933_));
 sg13g2_nand3_1 _23590_ (.B(net4553),
    .C(_05933_),
    .A(net5343),
    .Y(_05934_));
 sg13g2_nand2_1 _23591_ (.Y(_02022_),
    .A(_05929_),
    .B(_05934_));
 sg13g2_xnor2_1 _23592_ (.Y(_05935_),
    .A(_08101_),
    .B(_05932_));
 sg13g2_nor2_1 _23593_ (.A(net5303),
    .B(_05935_),
    .Y(_05936_));
 sg13g2_a22oi_1 _23594_ (.Y(_05937_),
    .B1(net4553),
    .B2(_05936_),
    .A2(net5276),
    .A1(net3328));
 sg13g2_inv_1 _23595_ (.Y(_02023_),
    .A(net3329));
 sg13g2_nand2_1 _23596_ (.Y(_05938_),
    .A(net3118),
    .B(net5276));
 sg13g2_nand3_1 _23597_ (.B(\atari2600.tia.audio_left_counter[10] ),
    .C(_05931_),
    .A(\atari2600.tia.audio_left_counter[11] ),
    .Y(_05939_));
 sg13g2_inv_1 _23598_ (.Y(_05940_),
    .A(_05939_));
 sg13g2_nor2_1 _23599_ (.A(_00119_),
    .B(_05939_),
    .Y(_05941_));
 sg13g2_xnor2_1 _23600_ (.Y(_05942_),
    .A(_08102_),
    .B(_05939_));
 sg13g2_nand3_1 _23601_ (.B(net4553),
    .C(_05942_),
    .A(net5343),
    .Y(_05943_));
 sg13g2_nand2_1 _23602_ (.Y(_02024_),
    .A(_05938_),
    .B(_05943_));
 sg13g2_xor2_1 _23603_ (.B(_05941_),
    .A(_00120_),
    .X(_05944_));
 sg13g2_nor2_1 _23604_ (.A(net5304),
    .B(_05944_),
    .Y(_05945_));
 sg13g2_a22oi_1 _23605_ (.Y(_05946_),
    .B1(net4553),
    .B2(_05945_),
    .A2(net5276),
    .A1(net3676));
 sg13g2_inv_1 _23606_ (.Y(_02025_),
    .A(net3677));
 sg13g2_nand2_1 _23607_ (.Y(_05947_),
    .A(net2974),
    .B(net5276));
 sg13g2_nand3_1 _23608_ (.B(\atari2600.tia.audio_left_counter[12] ),
    .C(_05940_),
    .A(\atari2600.tia.audio_left_counter[13] ),
    .Y(_05948_));
 sg13g2_nor2_1 _23609_ (.A(_00121_),
    .B(_05948_),
    .Y(_05949_));
 sg13g2_xor2_1 _23610_ (.B(_05948_),
    .A(_00121_),
    .X(_05950_));
 sg13g2_nand3_1 _23611_ (.B(net4553),
    .C(_05950_),
    .A(net5343),
    .Y(_05951_));
 sg13g2_nand2_1 _23612_ (.Y(_02026_),
    .A(_05947_),
    .B(_05951_));
 sg13g2_xnor2_1 _23613_ (.Y(_05952_),
    .A(_08103_),
    .B(_05949_));
 sg13g2_nor2_1 _23614_ (.A(net5303),
    .B(_05952_),
    .Y(_05953_));
 sg13g2_a22oi_1 _23615_ (.Y(_05954_),
    .B1(net4553),
    .B2(_05953_),
    .A2(net5278),
    .A1(net2970));
 sg13g2_inv_1 _23616_ (.Y(_02027_),
    .A(net2971));
 sg13g2_nand2_1 _23617_ (.Y(_05955_),
    .A(\atari2600.tia.audio_right_counter[0] ),
    .B(net5279));
 sg13g2_nor2_1 _23618_ (.A(_07965_),
    .B(\atari2600.tia.audc1[0] ),
    .Y(_05956_));
 sg13g2_nand2_1 _23619_ (.Y(_05957_),
    .A(\atari2600.tia.audc1[1] ),
    .B(_07966_));
 sg13g2_nor2_1 _23620_ (.A(_07963_),
    .B(net5583),
    .Y(_05958_));
 sg13g2_nor2_2 _23621_ (.A(\atari2600.tia.audc1[3] ),
    .B(net5583),
    .Y(_05959_));
 sg13g2_a22oi_1 _23622_ (.Y(_05960_),
    .B1(_05959_),
    .B2(_07966_),
    .A2(_05958_),
    .A1(\atari2600.tia.audc1[1] ));
 sg13g2_nor3_1 _23623_ (.A(\atari2600.tia.audc1[3] ),
    .B(net5583),
    .C(\atari2600.tia.audc1[1] ),
    .Y(_05961_));
 sg13g2_nor2_2 _23624_ (.A(_05956_),
    .B(_05960_),
    .Y(_05962_));
 sg13g2_and2_1 _23625_ (.A(net5578),
    .B(net5580),
    .X(_05963_));
 sg13g2_nand3_1 _23626_ (.B(\atari2600.tia.audf1[1] ),
    .C(net5580),
    .A(net5578),
    .Y(_05964_));
 sg13g2_nand4_1 _23627_ (.B(net5578),
    .C(net5579),
    .A(\atari2600.tia.audf1[3] ),
    .Y(_05965_),
    .D(net5580));
 sg13g2_inv_1 _23628_ (.Y(_05966_),
    .A(_05965_));
 sg13g2_nor2_1 _23629_ (.A(_00140_),
    .B(_05965_),
    .Y(_05967_));
 sg13g2_nand2_1 _23630_ (.Y(_05968_),
    .A(_00140_),
    .B(_05965_));
 sg13g2_nor2b_1 _23631_ (.A(_05967_),
    .B_N(_05968_),
    .Y(_05969_));
 sg13g2_nor2_1 _23632_ (.A(net5578),
    .B(net5580),
    .Y(_05970_));
 sg13g2_nor2_1 _23633_ (.A(\atari2600.tia.audf1[2] ),
    .B(net5579),
    .Y(_05971_));
 sg13g2_a21oi_1 _23634_ (.A1(net5579),
    .A2(net5580),
    .Y(_05972_),
    .B1(net5578));
 sg13g2_nor2b_1 _23635_ (.A(_05972_),
    .B_N(_05964_),
    .Y(_05973_));
 sg13g2_a22oi_1 _23636_ (.Y(_05974_),
    .B1(_05972_),
    .B2(\atari2600.tia.audf1[3] ),
    .A2(_05963_),
    .A1(net5579));
 sg13g2_xor2_1 _23637_ (.B(_05974_),
    .A(_00140_),
    .X(_05975_));
 sg13g2_xor2_1 _23638_ (.B(_05975_),
    .A(_00139_),
    .X(_05976_));
 sg13g2_xor2_1 _23639_ (.B(net5580),
    .A(net5579),
    .X(_05977_));
 sg13g2_xnor2_1 _23640_ (.Y(_05978_),
    .A(net5579),
    .B(net5580));
 sg13g2_nor3_1 _23641_ (.A(\atari2600.tia.audf1[3] ),
    .B(_07947_),
    .C(_05978_),
    .Y(_05979_));
 sg13g2_nand2_1 _23642_ (.Y(_05980_),
    .A(_05976_),
    .B(_05979_));
 sg13g2_xnor2_1 _23643_ (.Y(_05981_),
    .A(_05976_),
    .B(_05979_));
 sg13g2_nor4_2 _23644_ (.A(_07946_),
    .B(net5578),
    .C(_07948_),
    .Y(_05982_),
    .D(net5580));
 sg13g2_nand4_1 _23645_ (.B(net5579),
    .C(_05970_),
    .A(\atari2600.tia.audf1[3] ),
    .Y(_05983_),
    .D(_05976_));
 sg13g2_and2_1 _23646_ (.A(\atari2600.tia.audf1[3] ),
    .B(_05973_),
    .X(_05984_));
 sg13g2_a22oi_1 _23647_ (.Y(_05985_),
    .B1(_05984_),
    .B2(_00140_),
    .A2(_05975_),
    .A1(_00139_));
 sg13g2_xnor2_1 _23648_ (.Y(_05986_),
    .A(_07946_),
    .B(_05964_));
 sg13g2_nand2_1 _23649_ (.Y(_05987_),
    .A(_05968_),
    .B(_05986_));
 sg13g2_xnor2_1 _23650_ (.Y(_05988_),
    .A(_05978_),
    .B(_05987_));
 sg13g2_xnor2_1 _23651_ (.Y(_05989_),
    .A(_05985_),
    .B(_05988_));
 sg13g2_o21ai_1 _23652_ (.B1(_05983_),
    .Y(_05990_),
    .A1(_05980_),
    .A2(_05989_));
 sg13g2_nand2b_1 _23653_ (.Y(_05991_),
    .B(_05990_),
    .A_N(_00140_));
 sg13g2_a21oi_1 _23654_ (.A1(\atari2600.tia.audf1[4] ),
    .A2(_05966_),
    .Y(_05992_),
    .B1(_05973_));
 sg13g2_a22oi_1 _23655_ (.Y(_05993_),
    .B1(_05978_),
    .B2(_05986_),
    .A2(_05965_),
    .A1(_00140_));
 sg13g2_nor2b_1 _23656_ (.A(_05992_),
    .B_N(_05993_),
    .Y(_05994_));
 sg13g2_xor2_1 _23657_ (.B(_05993_),
    .A(_05992_),
    .X(_05995_));
 sg13g2_nor3_1 _23658_ (.A(_05985_),
    .B(_05988_),
    .C(_05995_),
    .Y(_05996_));
 sg13g2_nor2_1 _23659_ (.A(_05994_),
    .B(_05996_),
    .Y(_05997_));
 sg13g2_o21ai_1 _23660_ (.B1(_05991_),
    .Y(_05998_),
    .A1(_05986_),
    .A2(_05997_));
 sg13g2_a21oi_2 _23661_ (.B1(_05967_),
    .Y(_05999_),
    .A2(_05998_),
    .A1(_05968_));
 sg13g2_inv_1 _23662_ (.Y(_06000_),
    .A(_05999_));
 sg13g2_nor2_1 _23663_ (.A(net5450),
    .B(_05999_),
    .Y(_06001_));
 sg13g2_and2_1 _23664_ (.A(_05980_),
    .B(_05989_),
    .X(_06002_));
 sg13g2_nor2_2 _23665_ (.A(_05990_),
    .B(_06002_),
    .Y(_06003_));
 sg13g2_or2_2 _23666_ (.X(_06004_),
    .B(_06002_),
    .A(_05990_));
 sg13g2_nor2_1 _23667_ (.A(_07963_),
    .B(_07964_),
    .Y(_06005_));
 sg13g2_o21ai_1 _23668_ (.B1(_05995_),
    .Y(_06006_),
    .A1(_05985_),
    .A2(_05988_));
 sg13g2_nand2b_1 _23669_ (.Y(_06007_),
    .B(_06006_),
    .A_N(_05996_));
 sg13g2_a21oi_1 _23670_ (.A1(_05990_),
    .A2(_06006_),
    .Y(_06008_),
    .B1(_05996_));
 sg13g2_xnor2_1 _23671_ (.Y(_06009_),
    .A(_05986_),
    .B(_05994_));
 sg13g2_xnor2_1 _23672_ (.Y(_06010_),
    .A(_06008_),
    .B(_06009_));
 sg13g2_and2_1 _23673_ (.A(net5452),
    .B(_06010_),
    .X(_06011_));
 sg13g2_nand2_1 _23674_ (.Y(_06012_),
    .A(net5451),
    .B(_06010_));
 sg13g2_nor2_1 _23675_ (.A(net5450),
    .B(_06004_),
    .Y(_06013_));
 sg13g2_nor4_2 _23676_ (.A(_07963_),
    .B(_07964_),
    .C(_06004_),
    .Y(_06014_),
    .D(_06012_));
 sg13g2_xnor2_1 _23677_ (.Y(_06015_),
    .A(_05969_),
    .B(_05998_));
 sg13g2_xnor2_1 _23678_ (.Y(_06016_),
    .A(_05990_),
    .B(_06007_));
 sg13g2_nand3_1 _23679_ (.B(net5447),
    .C(net5320),
    .A(net5451),
    .Y(_06017_));
 sg13g2_nor2_1 _23680_ (.A(net5450),
    .B(_06015_),
    .Y(_06018_));
 sg13g2_or2_1 _23681_ (.X(_06019_),
    .B(_06017_),
    .A(_06015_));
 sg13g2_nor2_2 _23682_ (.A(net5449),
    .B(_05959_),
    .Y(_06020_));
 sg13g2_nand2b_1 _23683_ (.Y(_06021_),
    .B(net5452),
    .A_N(_05959_));
 sg13g2_o21ai_1 _23684_ (.B1(_06017_),
    .Y(_06022_),
    .A1(_06015_),
    .A2(_06021_));
 sg13g2_and2_1 _23685_ (.A(_06019_),
    .B(_06022_),
    .X(_06023_));
 sg13g2_and2_1 _23686_ (.A(_06014_),
    .B(_06023_),
    .X(_06024_));
 sg13g2_xor2_1 _23687_ (.B(_06023_),
    .A(_06014_),
    .X(_06025_));
 sg13g2_xnor2_1 _23688_ (.Y(_06026_),
    .A(_06001_),
    .B(_06025_));
 sg13g2_xnor2_1 _23689_ (.Y(_06027_),
    .A(_05981_),
    .B(_05982_));
 sg13g2_xor2_1 _23690_ (.B(_05982_),
    .A(_05981_),
    .X(_06028_));
 sg13g2_nand2_1 _23691_ (.Y(_06029_),
    .A(net5451),
    .B(_06027_));
 sg13g2_nor4_2 _23692_ (.A(_07963_),
    .B(_07964_),
    .C(net5449),
    .Y(_06030_),
    .D(_06028_));
 sg13g2_nand2_1 _23693_ (.Y(_06031_),
    .A(net5320),
    .B(_06030_));
 sg13g2_a22oi_1 _23694_ (.Y(_06032_),
    .B1(_06020_),
    .B2(_06010_),
    .A2(_06013_),
    .A1(net5448));
 sg13g2_or2_1 _23695_ (.X(_06033_),
    .B(_06032_),
    .A(_06014_));
 sg13g2_or2_1 _23696_ (.X(_06034_),
    .B(_06033_),
    .A(_06031_));
 sg13g2_xnor2_1 _23697_ (.Y(_06035_),
    .A(_06031_),
    .B(_06033_));
 sg13g2_nor2_2 _23698_ (.A(net5451),
    .B(net5448),
    .Y(_06036_));
 sg13g2_or2_2 _23699_ (.X(_06037_),
    .B(net5448),
    .A(net5451));
 sg13g2_a21oi_1 _23700_ (.A1(_06000_),
    .A2(_06037_),
    .Y(_06038_),
    .B1(_06018_));
 sg13g2_o21ai_1 _23701_ (.B1(_06034_),
    .Y(_06039_),
    .A1(_06035_),
    .A2(_06038_));
 sg13g2_nand2b_1 _23702_ (.Y(_06040_),
    .B(_06039_),
    .A_N(_06026_));
 sg13g2_xor2_1 _23703_ (.B(_06039_),
    .A(_06026_),
    .X(_06041_));
 sg13g2_a21oi_1 _23704_ (.A1(net5578),
    .A2(_05977_),
    .Y(_06042_),
    .B1(_05971_));
 sg13g2_xnor2_1 _23705_ (.Y(_06043_),
    .A(\atari2600.tia.audf1[3] ),
    .B(_06042_));
 sg13g2_xnor2_1 _23706_ (.Y(_06044_),
    .A(_07946_),
    .B(_06042_));
 sg13g2_nor2_2 _23707_ (.A(net5449),
    .B(_06043_),
    .Y(_06045_));
 sg13g2_and2_1 _23708_ (.A(net5447),
    .B(_06045_),
    .X(_06046_));
 sg13g2_nand2_1 _23709_ (.Y(_06047_),
    .A(_06003_),
    .B(_06046_));
 sg13g2_and2_1 _23710_ (.A(net5320),
    .B(_06020_),
    .X(_06048_));
 sg13g2_o21ai_1 _23711_ (.B1(_06031_),
    .Y(_06049_),
    .A1(_06030_),
    .A2(_06048_));
 sg13g2_nor2_1 _23712_ (.A(_06047_),
    .B(_06049_),
    .Y(_06050_));
 sg13g2_nor2_1 _23713_ (.A(net5449),
    .B(net5447),
    .Y(_06051_));
 sg13g2_nand2_1 _23714_ (.Y(_06052_),
    .A(_07963_),
    .B(\atari2600.tia.audc1[1] ));
 sg13g2_and3_2 _23715_ (.X(_06053_),
    .A(\atari2600.tia.audc1[2] ),
    .B(net5449),
    .C(_06052_));
 sg13g2_nand3_1 _23716_ (.B(net5449),
    .C(_06052_),
    .A(net5583),
    .Y(_06054_));
 sg13g2_nor2_2 _23717_ (.A(_06051_),
    .B(_06053_),
    .Y(_06055_));
 sg13g2_nand2b_2 _23718_ (.Y(_06056_),
    .B(_06054_),
    .A_N(_06051_));
 sg13g2_nor2_1 _23719_ (.A(_06012_),
    .B(_06015_),
    .Y(_06057_));
 sg13g2_o21ai_1 _23720_ (.B1(_06012_),
    .Y(_06058_),
    .A1(_06015_),
    .A2(_06036_));
 sg13g2_nand2b_1 _23721_ (.Y(_06059_),
    .B(_06058_),
    .A_N(_06057_));
 sg13g2_o21ai_1 _23722_ (.B1(_06059_),
    .Y(_06060_),
    .A1(_05999_),
    .A2(_06055_));
 sg13g2_xor2_1 _23723_ (.B(_06049_),
    .A(_06047_),
    .X(_06061_));
 sg13g2_a21oi_1 _23724_ (.A1(_06060_),
    .A2(_06061_),
    .Y(_06062_),
    .B1(_06050_));
 sg13g2_xor2_1 _23725_ (.B(_06038_),
    .A(_06035_),
    .X(_06063_));
 sg13g2_nor2b_1 _23726_ (.A(_06062_),
    .B_N(_06063_),
    .Y(_06064_));
 sg13g2_xnor2_1 _23727_ (.Y(_06065_),
    .A(_06062_),
    .B(_06063_));
 sg13g2_a21oi_1 _23728_ (.A1(_06057_),
    .A2(_06065_),
    .Y(_06066_),
    .B1(_06064_));
 sg13g2_nor2_1 _23729_ (.A(_06041_),
    .B(_06066_),
    .Y(_06067_));
 sg13g2_a21oi_1 _23730_ (.A1(_06001_),
    .A2(_06025_),
    .Y(_06068_),
    .B1(_06024_));
 sg13g2_a22oi_1 _23731_ (.Y(_06069_),
    .B1(_06020_),
    .B2(_06000_),
    .A2(_06011_),
    .A1(net5447));
 sg13g2_or2_1 _23732_ (.X(_06070_),
    .B(_06069_),
    .A(_06019_));
 sg13g2_xor2_1 _23733_ (.B(_06069_),
    .A(_06019_),
    .X(_06071_));
 sg13g2_inv_1 _23734_ (.Y(_06072_),
    .A(_06071_));
 sg13g2_nand2_1 _23735_ (.Y(_06073_),
    .A(_06068_),
    .B(_06071_));
 sg13g2_xor2_1 _23736_ (.B(_06073_),
    .A(_06040_),
    .X(_06074_));
 sg13g2_xnor2_1 _23737_ (.Y(_06075_),
    .A(_06057_),
    .B(_06065_));
 sg13g2_nor2_2 _23738_ (.A(_05963_),
    .B(_05970_),
    .Y(_06076_));
 sg13g2_nand2_1 _23739_ (.Y(_06077_),
    .A(net5452),
    .B(net5446));
 sg13g2_nand3_1 _23740_ (.B(net5448),
    .C(_06076_),
    .A(net5451),
    .Y(_06078_));
 sg13g2_nand2_1 _23741_ (.Y(_06079_),
    .A(_06030_),
    .B(_06076_));
 sg13g2_nor2_1 _23742_ (.A(_06004_),
    .B(_06021_),
    .Y(_06080_));
 sg13g2_o21ai_1 _23743_ (.B1(_06047_),
    .Y(_06081_),
    .A1(_06046_),
    .A2(_06080_));
 sg13g2_nor2_1 _23744_ (.A(_06015_),
    .B(_06055_),
    .Y(_06082_));
 sg13g2_a22oi_1 _23745_ (.Y(_06083_),
    .B1(_06037_),
    .B2(_06010_),
    .A2(net5320),
    .A1(net5451));
 sg13g2_a21oi_1 _23746_ (.A1(_06011_),
    .A2(_06016_),
    .Y(_06084_),
    .B1(_06083_));
 sg13g2_and2_1 _23747_ (.A(_06082_),
    .B(_06084_),
    .X(_06085_));
 sg13g2_xnor2_1 _23748_ (.Y(_06086_),
    .A(_06082_),
    .B(_06084_));
 sg13g2_xor2_1 _23749_ (.B(_06081_),
    .A(_06079_),
    .X(_06087_));
 sg13g2_nand2b_1 _23750_ (.Y(_06088_),
    .B(_06087_),
    .A_N(_06086_));
 sg13g2_o21ai_1 _23751_ (.B1(_06088_),
    .Y(_06089_),
    .A1(_06079_),
    .A2(_06081_));
 sg13g2_xnor2_1 _23752_ (.Y(_06090_),
    .A(_06060_),
    .B(_06061_));
 sg13g2_nand2b_1 _23753_ (.Y(_06091_),
    .B(_06089_),
    .A_N(_06090_));
 sg13g2_a21o_1 _23754_ (.A2(_06016_),
    .A1(_06011_),
    .B1(_06085_),
    .X(_06092_));
 sg13g2_xor2_1 _23755_ (.B(_06090_),
    .A(_06089_),
    .X(_06093_));
 sg13g2_nand2b_1 _23756_ (.Y(_06094_),
    .B(_06092_),
    .A_N(_06093_));
 sg13g2_a21oi_1 _23757_ (.A1(_06091_),
    .A2(_06094_),
    .Y(_06095_),
    .B1(_06075_));
 sg13g2_inv_1 _23758_ (.Y(_06096_),
    .A(_06095_));
 sg13g2_xnor2_1 _23759_ (.Y(_06097_),
    .A(_06041_),
    .B(_06066_));
 sg13g2_nor2_1 _23760_ (.A(_06096_),
    .B(_06097_),
    .Y(_06098_));
 sg13g2_xnor2_1 _23761_ (.Y(_06099_),
    .A(_06092_),
    .B(_06093_));
 sg13g2_xnor2_1 _23762_ (.Y(_06100_),
    .A(_00139_),
    .B(_05977_));
 sg13g2_nor2_2 _23763_ (.A(net5449),
    .B(_06100_),
    .Y(_06101_));
 sg13g2_nor2b_1 _23764_ (.A(_06100_),
    .B_N(_06046_),
    .Y(_06102_));
 sg13g2_nand2_1 _23765_ (.Y(_06103_),
    .A(_06020_),
    .B(_06027_));
 sg13g2_a22oi_1 _23766_ (.Y(_06104_),
    .B1(_06078_),
    .B2(_06103_),
    .A2(net5446),
    .A1(_06030_));
 sg13g2_and2_1 _23767_ (.A(_06102_),
    .B(_06104_),
    .X(_06105_));
 sg13g2_nand2_1 _23768_ (.Y(_06106_),
    .A(_06010_),
    .B(_06056_));
 sg13g2_a21oi_1 _23769_ (.A1(net5451),
    .A2(_06003_),
    .Y(_06107_),
    .B1(net5320));
 sg13g2_nor3_1 _23770_ (.A(net5450),
    .B(_06004_),
    .C(_06007_),
    .Y(_06108_));
 sg13g2_nor3_1 _23771_ (.A(_06036_),
    .B(_06107_),
    .C(_06108_),
    .Y(_06109_));
 sg13g2_nor2b_1 _23772_ (.A(_06106_),
    .B_N(_06109_),
    .Y(_06110_));
 sg13g2_xnor2_1 _23773_ (.Y(_06111_),
    .A(_06106_),
    .B(_06109_));
 sg13g2_or2_1 _23774_ (.X(_06112_),
    .B(_06104_),
    .A(_06102_));
 sg13g2_nand2b_1 _23775_ (.Y(_06113_),
    .B(_06112_),
    .A_N(_06105_));
 sg13g2_a21oi_1 _23776_ (.A1(_06111_),
    .A2(_06112_),
    .Y(_06114_),
    .B1(_06105_));
 sg13g2_xnor2_1 _23777_ (.Y(_06115_),
    .A(_06086_),
    .B(_06087_));
 sg13g2_nor2b_1 _23778_ (.A(_06114_),
    .B_N(_06115_),
    .Y(_06116_));
 sg13g2_nor2_1 _23779_ (.A(_06108_),
    .B(_06110_),
    .Y(_06117_));
 sg13g2_xor2_1 _23780_ (.B(_06115_),
    .A(_06114_),
    .X(_06118_));
 sg13g2_nor2_1 _23781_ (.A(_06117_),
    .B(_06118_),
    .Y(_06119_));
 sg13g2_nor2_2 _23782_ (.A(_06116_),
    .B(_06119_),
    .Y(_06120_));
 sg13g2_nand2b_1 _23783_ (.Y(_06121_),
    .B(_06099_),
    .A_N(_06120_));
 sg13g2_nand3_1 _23784_ (.B(_06091_),
    .C(_06094_),
    .A(_06075_),
    .Y(_06122_));
 sg13g2_nand2_1 _23785_ (.Y(_06123_),
    .A(_06096_),
    .B(_06122_));
 sg13g2_or2_1 _23786_ (.X(_06124_),
    .B(_06123_),
    .A(_06121_));
 sg13g2_xnor2_1 _23787_ (.Y(_06125_),
    .A(_06099_),
    .B(_06120_));
 sg13g2_nor2_1 _23788_ (.A(net5581),
    .B(net5449),
    .Y(_06126_));
 sg13g2_and3_1 _23789_ (.X(_06127_),
    .A(\atari2600.tia.audf1[2] ),
    .B(net5447),
    .C(_06126_));
 sg13g2_a22oi_1 _23790_ (.Y(_06128_),
    .B1(_06101_),
    .B2(net5447),
    .A2(_06044_),
    .A1(_06020_));
 sg13g2_or2_1 _23791_ (.X(_06129_),
    .B(_06128_),
    .A(_06102_));
 sg13g2_inv_1 _23792_ (.Y(_06130_),
    .A(_06129_));
 sg13g2_xor2_1 _23793_ (.B(_06129_),
    .A(_06127_),
    .X(_06131_));
 sg13g2_nand2_1 _23794_ (.Y(_06132_),
    .A(net5320),
    .B(_06056_));
 sg13g2_nor3_1 _23795_ (.A(_05990_),
    .B(_06002_),
    .C(_06036_),
    .Y(_06133_));
 sg13g2_mux2_1 _23796_ (.A0(_06004_),
    .A1(_06133_),
    .S(_06029_),
    .X(_06134_));
 sg13g2_nor2b_1 _23797_ (.A(_06132_),
    .B_N(_06134_),
    .Y(_06135_));
 sg13g2_xnor2_1 _23798_ (.Y(_06136_),
    .A(_06132_),
    .B(_06134_));
 sg13g2_nor2b_1 _23799_ (.A(_06131_),
    .B_N(_06136_),
    .Y(_06137_));
 sg13g2_a21oi_1 _23800_ (.A1(_06127_),
    .A2(_06130_),
    .Y(_06138_),
    .B1(_06137_));
 sg13g2_xor2_1 _23801_ (.B(_06113_),
    .A(_06111_),
    .X(_06139_));
 sg13g2_a21oi_1 _23802_ (.A1(_06013_),
    .A2(_06027_),
    .Y(_06140_),
    .B1(_06135_));
 sg13g2_xor2_1 _23803_ (.B(_06139_),
    .A(_06138_),
    .X(_06141_));
 sg13g2_nand2b_1 _23804_ (.Y(_06142_),
    .B(_06141_),
    .A_N(_06140_));
 sg13g2_o21ai_1 _23805_ (.B1(_06142_),
    .Y(_06143_),
    .A1(_06138_),
    .A2(_06139_));
 sg13g2_xor2_1 _23806_ (.B(_06118_),
    .A(_06117_),
    .X(_06144_));
 sg13g2_nor2_1 _23807_ (.A(_05999_),
    .B(_06053_),
    .Y(_06145_));
 sg13g2_xnor2_1 _23808_ (.Y(_06146_),
    .A(_06143_),
    .B(_06144_));
 sg13g2_nor3_1 _23809_ (.A(_05999_),
    .B(_06053_),
    .C(_06146_),
    .Y(_06147_));
 sg13g2_a21o_1 _23810_ (.A2(_06144_),
    .A1(_06143_),
    .B1(_06147_),
    .X(_06148_));
 sg13g2_and2_1 _23811_ (.A(_06125_),
    .B(_06148_),
    .X(_06149_));
 sg13g2_xnor2_1 _23812_ (.Y(_06150_),
    .A(_06028_),
    .B(_06045_));
 sg13g2_and4_1 _23813_ (.A(_06003_),
    .B(_06037_),
    .C(_06056_),
    .D(_06150_),
    .X(_06151_));
 sg13g2_a22oi_1 _23814_ (.Y(_06152_),
    .B1(_06150_),
    .B2(_06037_),
    .A2(_06056_),
    .A1(_06003_));
 sg13g2_a22oi_1 _23815_ (.Y(_06153_),
    .B1(_06126_),
    .B2(net5447),
    .A2(net5446),
    .A1(_06020_));
 sg13g2_or2_1 _23816_ (.X(_06154_),
    .B(_06153_),
    .A(_06127_));
 sg13g2_or3_1 _23817_ (.A(_06151_),
    .B(_06152_),
    .C(_06154_),
    .X(_06155_));
 sg13g2_xor2_1 _23818_ (.B(_06136_),
    .A(_06131_),
    .X(_06156_));
 sg13g2_nor2_1 _23819_ (.A(_06155_),
    .B(_06156_),
    .Y(_06157_));
 sg13g2_a21o_1 _23820_ (.A2(_06045_),
    .A1(_06027_),
    .B1(_06151_),
    .X(_06158_));
 sg13g2_xor2_1 _23821_ (.B(_06156_),
    .A(_06155_),
    .X(_06159_));
 sg13g2_a21oi_1 _23822_ (.A1(_06158_),
    .A2(_06159_),
    .Y(_06160_),
    .B1(_06157_));
 sg13g2_xor2_1 _23823_ (.B(_06141_),
    .A(_06140_),
    .X(_06161_));
 sg13g2_nor2_1 _23824_ (.A(_06160_),
    .B(_06161_),
    .Y(_06162_));
 sg13g2_nor2_2 _23825_ (.A(_06015_),
    .B(_06053_),
    .Y(_06163_));
 sg13g2_xor2_1 _23826_ (.B(_06161_),
    .A(_06160_),
    .X(_06164_));
 sg13g2_a21oi_2 _23827_ (.B1(_06162_),
    .Y(_06165_),
    .A2(_06164_),
    .A1(_06163_));
 sg13g2_xor2_1 _23828_ (.B(_06146_),
    .A(_06145_),
    .X(_06166_));
 sg13g2_nor2_1 _23829_ (.A(_06165_),
    .B(_06166_),
    .Y(_06167_));
 sg13g2_o21ai_1 _23830_ (.B1(_06154_),
    .Y(_06168_),
    .A1(_06151_),
    .A2(_06152_));
 sg13g2_nand2_1 _23831_ (.Y(_06169_),
    .A(_06045_),
    .B(net5446));
 sg13g2_o21ai_1 _23832_ (.B1(_06077_),
    .Y(_06170_),
    .A1(_06036_),
    .A2(_06043_));
 sg13g2_nand2_1 _23833_ (.Y(_06171_),
    .A(_06169_),
    .B(_06170_));
 sg13g2_nand4_1 _23834_ (.B(_06056_),
    .C(_06169_),
    .A(_06027_),
    .Y(_06172_),
    .D(_06170_));
 sg13g2_o21ai_1 _23835_ (.B1(_06171_),
    .Y(_06173_),
    .A1(_06028_),
    .A2(_06055_));
 sg13g2_nor2_1 _23836_ (.A(_06021_),
    .B(_06100_),
    .Y(_06174_));
 sg13g2_and3_1 _23837_ (.X(_06175_),
    .A(_06172_),
    .B(_06173_),
    .C(_06174_));
 sg13g2_nand3_1 _23838_ (.B(_06168_),
    .C(_06175_),
    .A(_06155_),
    .Y(_06176_));
 sg13g2_nand2_1 _23839_ (.Y(_06177_),
    .A(_06169_),
    .B(_06172_));
 sg13g2_a21o_1 _23840_ (.A2(_06168_),
    .A1(_06155_),
    .B1(_06175_),
    .X(_06178_));
 sg13g2_nand3_1 _23841_ (.B(_06177_),
    .C(_06178_),
    .A(_06176_),
    .Y(_06179_));
 sg13g2_nand2_1 _23842_ (.Y(_06180_),
    .A(_06176_),
    .B(_06179_));
 sg13g2_xnor2_1 _23843_ (.Y(_06181_),
    .A(_06158_),
    .B(_06159_));
 sg13g2_nand2b_1 _23844_ (.Y(_06182_),
    .B(_06180_),
    .A_N(_06181_));
 sg13g2_nand2_1 _23845_ (.Y(_06183_),
    .A(_06010_),
    .B(_06054_));
 sg13g2_xor2_1 _23846_ (.B(_06181_),
    .A(_06180_),
    .X(_06184_));
 sg13g2_o21ai_1 _23847_ (.B1(_06182_),
    .Y(_06185_),
    .A1(_06183_),
    .A2(_06184_));
 sg13g2_xnor2_1 _23848_ (.Y(_06186_),
    .A(_06163_),
    .B(_06164_));
 sg13g2_nand2b_1 _23849_ (.Y(_06187_),
    .B(_06185_),
    .A_N(_06186_));
 sg13g2_nand2_1 _23850_ (.Y(_06188_),
    .A(net5446),
    .B(_06101_));
 sg13g2_or2_1 _23851_ (.X(_06189_),
    .B(_06101_),
    .A(net5446));
 sg13g2_nand3_1 _23852_ (.B(_06188_),
    .C(_06189_),
    .A(_06037_),
    .Y(_06190_));
 sg13g2_nand2_1 _23853_ (.Y(_06191_),
    .A(_06044_),
    .B(_06056_));
 sg13g2_xor2_1 _23854_ (.B(_06191_),
    .A(_06190_),
    .X(_06192_));
 sg13g2_nand3_1 _23855_ (.B(_06020_),
    .C(_06192_),
    .A(_00139_),
    .Y(_06193_));
 sg13g2_a21oi_1 _23856_ (.A1(_06172_),
    .A2(_06173_),
    .Y(_06194_),
    .B1(_06174_));
 sg13g2_or3_1 _23857_ (.A(_06175_),
    .B(_06193_),
    .C(_06194_),
    .X(_06195_));
 sg13g2_o21ai_1 _23858_ (.B1(_06188_),
    .Y(_06196_),
    .A1(_06190_),
    .A2(_06191_));
 sg13g2_o21ai_1 _23859_ (.B1(_06193_),
    .Y(_06197_),
    .A1(_06175_),
    .A2(_06194_));
 sg13g2_and3_1 _23860_ (.X(_06198_),
    .A(_06195_),
    .B(_06196_),
    .C(_06197_));
 sg13g2_nand3_1 _23861_ (.B(_06196_),
    .C(_06197_),
    .A(_06195_),
    .Y(_06199_));
 sg13g2_nand2_1 _23862_ (.Y(_06200_),
    .A(_06195_),
    .B(_06199_));
 sg13g2_a21o_1 _23863_ (.A2(_06178_),
    .A1(_06176_),
    .B1(_06177_),
    .X(_06201_));
 sg13g2_and3_1 _23864_ (.X(_06202_),
    .A(_06179_),
    .B(_06200_),
    .C(_06201_));
 sg13g2_nand3_1 _23865_ (.B(_06200_),
    .C(_06201_),
    .A(_06179_),
    .Y(_06203_));
 sg13g2_and2_1 _23866_ (.A(net5320),
    .B(net5400),
    .X(_06204_));
 sg13g2_nand2_1 _23867_ (.Y(_06205_),
    .A(net5320),
    .B(net5400));
 sg13g2_a21oi_1 _23868_ (.A1(_06179_),
    .A2(_06201_),
    .Y(_06206_),
    .B1(_06200_));
 sg13g2_a21o_1 _23869_ (.A2(_06201_),
    .A1(_06179_),
    .B1(_06200_),
    .X(_06207_));
 sg13g2_nor3_1 _23870_ (.A(_06202_),
    .B(_06205_),
    .C(_06206_),
    .Y(_06208_));
 sg13g2_o21ai_1 _23871_ (.B1(_06203_),
    .Y(_06209_),
    .A1(_06205_),
    .A2(_06206_));
 sg13g2_xor2_1 _23872_ (.B(_06184_),
    .A(_06183_),
    .X(_06210_));
 sg13g2_and2_1 _23873_ (.A(_06209_),
    .B(_06210_),
    .X(_06211_));
 sg13g2_nand2_1 _23874_ (.Y(_06212_),
    .A(_07949_),
    .B(_06101_));
 sg13g2_nand2_1 _23875_ (.Y(_06213_),
    .A(_06056_),
    .B(net5446));
 sg13g2_nor2_1 _23876_ (.A(_06036_),
    .B(_06100_),
    .Y(_06214_));
 sg13g2_o21ai_1 _23877_ (.B1(_06212_),
    .Y(_06215_),
    .A1(_06126_),
    .A2(_06214_));
 sg13g2_o21ai_1 _23878_ (.B1(_06212_),
    .Y(_06216_),
    .A1(_06213_),
    .A2(_06215_));
 sg13g2_a21o_1 _23879_ (.A2(_06020_),
    .A1(_00139_),
    .B1(_06192_),
    .X(_06217_));
 sg13g2_nand2_1 _23880_ (.Y(_06218_),
    .A(_06193_),
    .B(_06217_));
 sg13g2_nand2b_1 _23881_ (.Y(_06219_),
    .B(_06216_),
    .A_N(_06218_));
 sg13g2_a21oi_2 _23882_ (.B1(_06196_),
    .Y(_06220_),
    .A2(_06197_),
    .A1(_06195_));
 sg13g2_nor3_2 _23883_ (.A(_06198_),
    .B(_06219_),
    .C(_06220_),
    .Y(_06221_));
 sg13g2_or3_1 _23884_ (.A(_06198_),
    .B(_06219_),
    .C(_06220_),
    .X(_06222_));
 sg13g2_o21ai_1 _23885_ (.B1(_06219_),
    .Y(_06223_),
    .A1(_06198_),
    .A2(_06220_));
 sg13g2_and4_2 _23886_ (.A(_06003_),
    .B(net5400),
    .C(_06222_),
    .D(_06223_),
    .X(_06224_));
 sg13g2_nor2_1 _23887_ (.A(_06221_),
    .B(_06224_),
    .Y(_06225_));
 sg13g2_a21oi_1 _23888_ (.A1(_06203_),
    .A2(_06207_),
    .Y(_06226_),
    .B1(_06204_));
 sg13g2_nor3_1 _23889_ (.A(_06202_),
    .B(_06204_),
    .C(_06206_),
    .Y(_06227_));
 sg13g2_a21oi_1 _23890_ (.A1(_06203_),
    .A2(_06207_),
    .Y(_06228_),
    .B1(_06205_));
 sg13g2_nor3_1 _23891_ (.A(_06208_),
    .B(_06225_),
    .C(_06226_),
    .Y(_06229_));
 sg13g2_or3_1 _23892_ (.A(_06208_),
    .B(_06225_),
    .C(_06226_),
    .X(_06230_));
 sg13g2_xnor2_1 _23893_ (.Y(_06231_),
    .A(_06216_),
    .B(_06218_));
 sg13g2_nor2_1 _23894_ (.A(_06055_),
    .B(_06100_),
    .Y(_06232_));
 sg13g2_nor2_1 _23895_ (.A(net5581),
    .B(_06036_),
    .Y(_06233_));
 sg13g2_nand2_1 _23896_ (.Y(_06234_),
    .A(_06232_),
    .B(_06233_));
 sg13g2_xnor2_1 _23897_ (.Y(_06235_),
    .A(_06213_),
    .B(_06215_));
 sg13g2_nor2_1 _23898_ (.A(_06234_),
    .B(_06235_),
    .Y(_06236_));
 sg13g2_nand2_1 _23899_ (.Y(_06237_),
    .A(_06027_),
    .B(net5400));
 sg13g2_xnor2_1 _23900_ (.Y(_06238_),
    .A(_06231_),
    .B(_06236_));
 sg13g2_nor2_1 _23901_ (.A(_06237_),
    .B(_06238_),
    .Y(_06239_));
 sg13g2_a21oi_1 _23902_ (.A1(_06231_),
    .A2(_06236_),
    .Y(_06240_),
    .B1(_06239_));
 sg13g2_a22oi_1 _23903_ (.Y(_06241_),
    .B1(_06222_),
    .B2(_06223_),
    .A2(net5400),
    .A1(_06003_));
 sg13g2_nor3_1 _23904_ (.A(_06224_),
    .B(_06240_),
    .C(_06241_),
    .Y(_06242_));
 sg13g2_nand2_1 _23905_ (.Y(_06243_),
    .A(_06044_),
    .B(net5400));
 sg13g2_xor2_1 _23906_ (.B(_06235_),
    .A(_06234_),
    .X(_06244_));
 sg13g2_nand2b_1 _23907_ (.Y(_06245_),
    .B(_06244_),
    .A_N(_06243_));
 sg13g2_xnor2_1 _23908_ (.Y(_06246_),
    .A(_06243_),
    .B(_06244_));
 sg13g2_nand2_1 _23909_ (.Y(_06247_),
    .A(net5400),
    .B(net5446));
 sg13g2_xnor2_1 _23910_ (.Y(_06248_),
    .A(_06232_),
    .B(_06233_));
 sg13g2_nor2_1 _23911_ (.A(_06247_),
    .B(_06248_),
    .Y(_06249_));
 sg13g2_xor2_1 _23912_ (.B(_06248_),
    .A(_06247_),
    .X(_06250_));
 sg13g2_inv_1 _23913_ (.Y(_06251_),
    .A(_06250_));
 sg13g2_nand3_1 _23914_ (.B(_05978_),
    .C(_06051_),
    .A(_00139_),
    .Y(_06252_));
 sg13g2_nor2_1 _23915_ (.A(_06251_),
    .B(_06252_),
    .Y(_06253_));
 sg13g2_o21ai_1 _23916_ (.B1(_06246_),
    .Y(_06254_),
    .A1(_06249_),
    .A2(_06253_));
 sg13g2_and2_1 _23917_ (.A(_06245_),
    .B(_06254_),
    .X(_06255_));
 sg13g2_xnor2_1 _23918_ (.Y(_06256_),
    .A(_06237_),
    .B(_06238_));
 sg13g2_nor2_1 _23919_ (.A(_06255_),
    .B(_06256_),
    .Y(_06257_));
 sg13g2_o21ai_1 _23920_ (.B1(_06240_),
    .Y(_06258_),
    .A1(_06224_),
    .A2(_06241_));
 sg13g2_nor2b_1 _23921_ (.A(_06242_),
    .B_N(_06258_),
    .Y(_06259_));
 sg13g2_a21oi_1 _23922_ (.A1(_06257_),
    .A2(_06258_),
    .Y(_06260_),
    .B1(_06242_));
 sg13g2_nor4_2 _23923_ (.A(_06221_),
    .B(_06224_),
    .C(_06227_),
    .Y(_06261_),
    .D(_06228_));
 sg13g2_nor3_1 _23924_ (.A(_06229_),
    .B(_06260_),
    .C(_06261_),
    .Y(_06262_));
 sg13g2_o21ai_1 _23925_ (.B1(_06230_),
    .Y(_06263_),
    .A1(_06260_),
    .A2(_06261_));
 sg13g2_xor2_1 _23926_ (.B(_06210_),
    .A(_06209_),
    .X(_06264_));
 sg13g2_a21oi_1 _23927_ (.A1(_06263_),
    .A2(_06264_),
    .Y(_06265_),
    .B1(_06211_));
 sg13g2_xor2_1 _23928_ (.B(_06186_),
    .A(_06185_),
    .X(_06266_));
 sg13g2_o21ai_1 _23929_ (.B1(_06187_),
    .Y(_06267_),
    .A1(_06265_),
    .A2(_06266_));
 sg13g2_nand2_1 _23930_ (.Y(_06268_),
    .A(_06165_),
    .B(_06166_));
 sg13g2_xnor2_1 _23931_ (.Y(_06269_),
    .A(_06165_),
    .B(_06166_));
 sg13g2_a21o_1 _23932_ (.A2(_06268_),
    .A1(_06267_),
    .B1(_06167_),
    .X(_06270_));
 sg13g2_xor2_1 _23933_ (.B(_06148_),
    .A(_06125_),
    .X(_06271_));
 sg13g2_a21oi_1 _23934_ (.A1(_06270_),
    .A2(_06271_),
    .Y(_06272_),
    .B1(_06149_));
 sg13g2_and2_1 _23935_ (.A(_06121_),
    .B(_06123_),
    .X(_06273_));
 sg13g2_xor2_1 _23936_ (.B(_06123_),
    .A(_06121_),
    .X(_06274_));
 sg13g2_o21ai_1 _23937_ (.B1(_06124_),
    .Y(_06275_),
    .A1(_06272_),
    .A2(_06273_));
 sg13g2_xnor2_1 _23938_ (.Y(_06276_),
    .A(_06095_),
    .B(_06097_));
 sg13g2_a21oi_1 _23939_ (.A1(_06275_),
    .A2(_06276_),
    .Y(_06277_),
    .B1(_06098_));
 sg13g2_xnor2_1 _23940_ (.Y(_06278_),
    .A(_06067_),
    .B(_06074_));
 sg13g2_nor2_1 _23941_ (.A(_06277_),
    .B(_06278_),
    .Y(_06279_));
 sg13g2_a21oi_1 _23942_ (.A1(_06067_),
    .A2(_06074_),
    .Y(_06280_),
    .B1(_06279_));
 sg13g2_a21oi_1 _23943_ (.A1(_06040_),
    .A2(_06068_),
    .Y(_06281_),
    .B1(_06072_));
 sg13g2_nand3_1 _23944_ (.B(_06018_),
    .C(_06070_),
    .A(net5447),
    .Y(_06282_));
 sg13g2_xnor2_1 _23945_ (.Y(_06283_),
    .A(_06281_),
    .B(_06282_));
 sg13g2_xnor2_1 _23946_ (.Y(_06284_),
    .A(_06280_),
    .B(_06283_));
 sg13g2_xnor2_1 _23947_ (.Y(_06285_),
    .A(_06275_),
    .B(_06276_));
 sg13g2_nor2_1 _23948_ (.A(_08105_),
    .B(_06285_),
    .Y(_06286_));
 sg13g2_xor2_1 _23949_ (.B(_06271_),
    .A(_06270_),
    .X(_06287_));
 sg13g2_nor2_1 _23950_ (.A(_00132_),
    .B(_06287_),
    .Y(_06288_));
 sg13g2_nand2_1 _23951_ (.Y(_06289_),
    .A(_00132_),
    .B(_06287_));
 sg13g2_xor2_1 _23952_ (.B(_06266_),
    .A(_06265_),
    .X(_06290_));
 sg13g2_or2_1 _23953_ (.X(_06291_),
    .B(_06290_),
    .A(_00130_));
 sg13g2_xnor2_1 _23954_ (.Y(_06292_),
    .A(_06263_),
    .B(_06264_));
 sg13g2_and2_1 _23955_ (.A(\atari2600.tia.audio_right_counter[8] ),
    .B(_06292_),
    .X(_06293_));
 sg13g2_xor2_1 _23956_ (.B(_06292_),
    .A(_00129_),
    .X(_06294_));
 sg13g2_o21ai_1 _23957_ (.B1(_06260_),
    .Y(_06295_),
    .A1(_06229_),
    .A2(_06261_));
 sg13g2_nand2b_1 _23958_ (.Y(_06296_),
    .B(_06295_),
    .A_N(_06262_));
 sg13g2_nor2_1 _23959_ (.A(_08104_),
    .B(_06296_),
    .Y(_06297_));
 sg13g2_xnor2_1 _23960_ (.Y(_06298_),
    .A(_06257_),
    .B(_06259_));
 sg13g2_xor2_1 _23961_ (.B(_06256_),
    .A(_06255_),
    .X(_06299_));
 sg13g2_or3_1 _23962_ (.A(_06246_),
    .B(_06249_),
    .C(_06253_),
    .X(_06300_));
 sg13g2_and2_1 _23963_ (.A(_06254_),
    .B(_06300_),
    .X(_06301_));
 sg13g2_nand2_1 _23964_ (.Y(_06302_),
    .A(_00139_),
    .B(_06056_));
 sg13g2_o21ai_1 _23965_ (.B1(_06302_),
    .Y(_06303_),
    .A1(_06053_),
    .A2(_06100_));
 sg13g2_nand2_1 _23966_ (.Y(_06304_),
    .A(_06252_),
    .B(_06303_));
 sg13g2_nand3b_1 _23967_ (.B(_00139_),
    .C(net5400),
    .Y(_06305_),
    .A_N(\atari2600.tia.audio_right_counter[1] ));
 sg13g2_xnor2_1 _23968_ (.Y(_06306_),
    .A(_00123_),
    .B(_06304_));
 sg13g2_xnor2_1 _23969_ (.Y(_06307_),
    .A(_06250_),
    .B(_06252_));
 sg13g2_nor2_1 _23970_ (.A(_00124_),
    .B(_06307_),
    .Y(_06308_));
 sg13g2_a221oi_1 _23971_ (.B2(_06306_),
    .C1(_06308_),
    .B1(_06305_),
    .A1(\atari2600.tia.audio_right_counter[2] ),
    .Y(_06309_),
    .A2(_06304_));
 sg13g2_a21oi_1 _23972_ (.A1(_00124_),
    .A2(_06307_),
    .Y(_06310_),
    .B1(_06309_));
 sg13g2_a21oi_1 _23973_ (.A1(_00125_),
    .A2(_06310_),
    .Y(_06311_),
    .B1(\atari2600.tia.audio_right_counter[4] ));
 sg13g2_nor2b_1 _23974_ (.A(_00125_),
    .B_N(_06310_),
    .Y(_06312_));
 sg13g2_nor2_1 _23975_ (.A(_06301_),
    .B(_06311_),
    .Y(_06313_));
 sg13g2_a21oi_1 _23976_ (.A1(_06301_),
    .A2(_06312_),
    .Y(_06314_),
    .B1(_06313_));
 sg13g2_a21o_1 _23977_ (.A2(_06299_),
    .A1(_00126_),
    .B1(_06314_),
    .X(_06315_));
 sg13g2_o21ai_1 _23978_ (.B1(_06315_),
    .Y(_06316_),
    .A1(_00126_),
    .A2(_06299_));
 sg13g2_and2_1 _23979_ (.A(\atari2600.tia.audio_right_counter[6] ),
    .B(_06298_),
    .X(_06317_));
 sg13g2_xnor2_1 _23980_ (.Y(_06318_),
    .A(_00127_),
    .B(_06298_));
 sg13g2_a221oi_1 _23981_ (.B2(_06318_),
    .C1(_06317_),
    .B1(_06316_),
    .A1(_08104_),
    .Y(_06319_),
    .A2(_06296_));
 sg13g2_nor3_1 _23982_ (.A(_06294_),
    .B(_06297_),
    .C(_06319_),
    .Y(_06320_));
 sg13g2_nand2_1 _23983_ (.Y(_06321_),
    .A(_00130_),
    .B(_06290_));
 sg13g2_o21ai_1 _23984_ (.B1(_06321_),
    .Y(_06322_),
    .A1(_06293_),
    .A2(_06320_));
 sg13g2_xnor2_1 _23985_ (.Y(_06323_),
    .A(_06267_),
    .B(_06269_));
 sg13g2_xnor2_1 _23986_ (.Y(_06324_),
    .A(_00131_),
    .B(_06323_));
 sg13g2_a21oi_1 _23987_ (.A1(_06291_),
    .A2(_06322_),
    .Y(_06325_),
    .B1(_06324_));
 sg13g2_nor2b_1 _23988_ (.A(_06323_),
    .B_N(\atari2600.tia.audio_right_counter[10] ),
    .Y(_06326_));
 sg13g2_or3_1 _23989_ (.A(_06288_),
    .B(_06325_),
    .C(_06326_),
    .X(_06327_));
 sg13g2_xnor2_1 _23990_ (.Y(_06328_),
    .A(_06272_),
    .B(_06274_));
 sg13g2_xor2_1 _23991_ (.B(_06328_),
    .A(_00133_),
    .X(_06329_));
 sg13g2_nand3_1 _23992_ (.B(_06327_),
    .C(_06329_),
    .A(_06289_),
    .Y(_06330_));
 sg13g2_nor2b_1 _23993_ (.A(_06328_),
    .B_N(\atari2600.tia.audio_right_counter[12] ),
    .Y(_06331_));
 sg13g2_a21oi_1 _23994_ (.A1(_08105_),
    .A2(_06285_),
    .Y(_06332_),
    .B1(_06331_));
 sg13g2_a21oi_1 _23995_ (.A1(_06330_),
    .A2(_06332_),
    .Y(_06333_),
    .B1(_06286_));
 sg13g2_xnor2_1 _23996_ (.Y(_06334_),
    .A(_06277_),
    .B(_06278_));
 sg13g2_xnor2_1 _23997_ (.Y(_06335_),
    .A(_00135_),
    .B(_06334_));
 sg13g2_a22oi_1 _23998_ (.Y(_06336_),
    .B1(_06335_),
    .B2(_06333_),
    .A2(_06334_),
    .A1(\atari2600.tia.audio_right_counter[14] ));
 sg13g2_a21o_1 _23999_ (.A2(_06284_),
    .A1(_00136_),
    .B1(_06336_),
    .X(_06337_));
 sg13g2_o21ai_1 _24000_ (.B1(_06337_),
    .Y(_06338_),
    .A1(_00136_),
    .A2(_06284_));
 sg13g2_nor2_2 _24001_ (.A(_05962_),
    .B(_06338_),
    .Y(_06339_));
 sg13g2_a22oi_1 _24002_ (.Y(_06340_),
    .B1(_06339_),
    .B2(_08032_),
    .A2(_05962_),
    .A1(net2903));
 sg13g2_o21ai_1 _24003_ (.B1(_05955_),
    .Y(_02028_),
    .A1(net5306),
    .A2(net2904));
 sg13g2_nor2b_1 _24004_ (.A(_05962_),
    .B_N(_06338_),
    .Y(_06341_));
 sg13g2_nand2_1 _24005_ (.Y(_06342_),
    .A(\atari2600.tia.audio_right_counter[1] ),
    .B(\atari2600.tia.audio_right_counter[0] ));
 sg13g2_xnor2_1 _24006_ (.Y(_06343_),
    .A(net7244),
    .B(\atari2600.tia.audio_right_counter[0] ));
 sg13g2_nor3_1 _24007_ (.A(net5306),
    .B(net4554),
    .C(_06343_),
    .Y(_06344_));
 sg13g2_a21o_1 _24008_ (.A2(net5279),
    .A1(net7244),
    .B1(_06344_),
    .X(_02029_));
 sg13g2_nor2_1 _24009_ (.A(_00123_),
    .B(_06342_),
    .Y(_06345_));
 sg13g2_and2_1 _24010_ (.A(_00123_),
    .B(_06342_),
    .X(_06346_));
 sg13g2_nor4_1 _24011_ (.A(net5306),
    .B(net4554),
    .C(_06345_),
    .D(_06346_),
    .Y(_06347_));
 sg13g2_a21o_1 _24012_ (.A2(net5279),
    .A1(net6889),
    .B1(_06347_),
    .X(_02030_));
 sg13g2_xor2_1 _24013_ (.B(_06345_),
    .A(_00124_),
    .X(_06348_));
 sg13g2_nor3_1 _24014_ (.A(net5306),
    .B(net4554),
    .C(_06348_),
    .Y(_06349_));
 sg13g2_a21o_1 _24015_ (.A2(net5279),
    .A1(net3838),
    .B1(_06349_),
    .X(_02031_));
 sg13g2_nand4_1 _24016_ (.B(\atari2600.tia.audio_right_counter[2] ),
    .C(\atari2600.tia.audio_right_counter[1] ),
    .A(\atari2600.tia.audio_right_counter[3] ),
    .Y(_06350_),
    .D(\atari2600.tia.audio_right_counter[0] ));
 sg13g2_nor2_1 _24017_ (.A(_00125_),
    .B(_06350_),
    .Y(_06351_));
 sg13g2_and2_1 _24018_ (.A(_00125_),
    .B(_06350_),
    .X(_06352_));
 sg13g2_nor4_1 _24019_ (.A(net5305),
    .B(net4554),
    .C(_06351_),
    .D(_06352_),
    .Y(_06353_));
 sg13g2_a21o_1 _24020_ (.A2(net5279),
    .A1(net6284),
    .B1(_06353_),
    .X(_02032_));
 sg13g2_xor2_1 _24021_ (.B(_06351_),
    .A(_00126_),
    .X(_06354_));
 sg13g2_nor3_1 _24022_ (.A(net5305),
    .B(net4554),
    .C(_06354_),
    .Y(_06355_));
 sg13g2_a21o_1 _24023_ (.A2(net5279),
    .A1(net4135),
    .B1(_06355_),
    .X(_02033_));
 sg13g2_nand2_1 _24024_ (.Y(_06356_),
    .A(\atari2600.tia.audio_right_counter[5] ),
    .B(\atari2600.tia.audio_right_counter[4] ));
 sg13g2_nor2_1 _24025_ (.A(_06350_),
    .B(_06356_),
    .Y(_06357_));
 sg13g2_nor2b_1 _24026_ (.A(_06357_),
    .B_N(_00127_),
    .Y(_06358_));
 sg13g2_nor3_1 _24027_ (.A(_00127_),
    .B(_06350_),
    .C(_06356_),
    .Y(_06359_));
 sg13g2_nor4_1 _24028_ (.A(net5305),
    .B(net4554),
    .C(_06358_),
    .D(_06359_),
    .Y(_06360_));
 sg13g2_a21o_1 _24029_ (.A2(net5277),
    .A1(net6832),
    .B1(_06360_),
    .X(_02034_));
 sg13g2_xnor2_1 _24030_ (.Y(_06361_),
    .A(_08104_),
    .B(_06359_));
 sg13g2_nor3_1 _24031_ (.A(net5305),
    .B(net4554),
    .C(_06361_),
    .Y(_06362_));
 sg13g2_a21o_1 _24032_ (.A2(net5277),
    .A1(net3926),
    .B1(_06362_),
    .X(_02035_));
 sg13g2_nand3_1 _24033_ (.B(\atari2600.tia.audio_right_counter[6] ),
    .C(_06357_),
    .A(net3926),
    .Y(_06363_));
 sg13g2_inv_1 _24034_ (.Y(_06364_),
    .A(_06363_));
 sg13g2_and2_1 _24035_ (.A(_00129_),
    .B(_06363_),
    .X(_06365_));
 sg13g2_nor2_1 _24036_ (.A(_00129_),
    .B(_06363_),
    .Y(_06366_));
 sg13g2_nor4_1 _24037_ (.A(net5305),
    .B(net4555),
    .C(_06365_),
    .D(_06366_),
    .Y(_06367_));
 sg13g2_a21o_1 _24038_ (.A2(net5277),
    .A1(net6791),
    .B1(_06367_),
    .X(_02036_));
 sg13g2_xor2_1 _24039_ (.B(_06366_),
    .A(_00130_),
    .X(_06368_));
 sg13g2_nor3_1 _24040_ (.A(net5303),
    .B(net4555),
    .C(_06368_),
    .Y(_06369_));
 sg13g2_a21o_1 _24041_ (.A2(net5277),
    .A1(net3982),
    .B1(_06369_),
    .X(_02037_));
 sg13g2_nand3_1 _24042_ (.B(\atari2600.tia.audio_right_counter[8] ),
    .C(_06364_),
    .A(net3982),
    .Y(_06370_));
 sg13g2_inv_1 _24043_ (.Y(_06371_),
    .A(_06370_));
 sg13g2_and2_1 _24044_ (.A(_00131_),
    .B(_06370_),
    .X(_06372_));
 sg13g2_nor2_1 _24045_ (.A(_00131_),
    .B(_06370_),
    .Y(_06373_));
 sg13g2_nor4_1 _24046_ (.A(net5303),
    .B(net4555),
    .C(_06372_),
    .D(_06373_),
    .Y(_06374_));
 sg13g2_a21o_1 _24047_ (.A2(net5277),
    .A1(net6203),
    .B1(_06374_),
    .X(_02038_));
 sg13g2_xor2_1 _24048_ (.B(_06373_),
    .A(_00132_),
    .X(_06375_));
 sg13g2_nor3_1 _24049_ (.A(net5303),
    .B(net4555),
    .C(_06375_),
    .Y(_06376_));
 sg13g2_a21o_1 _24050_ (.A2(net5277),
    .A1(net3754),
    .B1(_06376_),
    .X(_02039_));
 sg13g2_and3_1 _24051_ (.X(_06377_),
    .A(\atari2600.tia.audio_right_counter[11] ),
    .B(\atari2600.tia.audio_right_counter[10] ),
    .C(_06371_));
 sg13g2_nor2b_1 _24052_ (.A(_06377_),
    .B_N(_00133_),
    .Y(_06378_));
 sg13g2_nor2b_1 _24053_ (.A(_00133_),
    .B_N(_06377_),
    .Y(_06379_));
 sg13g2_nor4_1 _24054_ (.A(net5304),
    .B(net4554),
    .C(_06378_),
    .D(_06379_),
    .Y(_06380_));
 sg13g2_a21o_1 _24055_ (.A2(net5280),
    .A1(net6998),
    .B1(_06380_),
    .X(_02040_));
 sg13g2_xnor2_1 _24056_ (.Y(_06381_),
    .A(_08105_),
    .B(_06379_));
 sg13g2_nor3_1 _24057_ (.A(net5303),
    .B(net4555),
    .C(_06381_),
    .Y(_06382_));
 sg13g2_a21o_1 _24058_ (.A2(net5276),
    .A1(net3856),
    .B1(_06382_),
    .X(_02041_));
 sg13g2_nand3_1 _24059_ (.B(\atari2600.tia.audio_right_counter[12] ),
    .C(_06377_),
    .A(net3856),
    .Y(_06383_));
 sg13g2_and2_1 _24060_ (.A(_00135_),
    .B(_06383_),
    .X(_06384_));
 sg13g2_nor2_1 _24061_ (.A(_00135_),
    .B(_06383_),
    .Y(_06385_));
 sg13g2_nor4_1 _24062_ (.A(net5304),
    .B(net4555),
    .C(_06384_),
    .D(_06385_),
    .Y(_06386_));
 sg13g2_a21o_1 _24063_ (.A2(net5276),
    .A1(net4007),
    .B1(_06386_),
    .X(_02042_));
 sg13g2_xor2_1 _24064_ (.B(_06385_),
    .A(_00136_),
    .X(_06387_));
 sg13g2_nor3_1 _24065_ (.A(net5304),
    .B(net4555),
    .C(_06387_),
    .Y(_06388_));
 sg13g2_a21o_1 _24066_ (.A2(net5278),
    .A1(net3000),
    .B1(_06388_),
    .X(_02043_));
 sg13g2_o21ai_1 _24067_ (.B1(net5354),
    .Y(_06389_),
    .A1(_05502_),
    .A2(_05888_));
 sg13g2_nor2_1 _24068_ (.A(\atari2600.tia.audc0[1] ),
    .B(_07968_),
    .Y(_06390_));
 sg13g2_nor3_1 _24069_ (.A(\atari2600.tia.audc0[3] ),
    .B(_07967_),
    .C(_07968_),
    .Y(_06391_));
 sg13g2_a22oi_1 _24070_ (.Y(_06392_),
    .B1(_06391_),
    .B2(\atari2600.tia.audc0[2] ),
    .A2(_06390_),
    .A1(_05500_));
 sg13g2_nand2_1 _24071_ (.Y(_06393_),
    .A(_05498_),
    .B(_05500_));
 sg13g2_mux2_1 _24072_ (.A0(\atari2600.tia.p5_l ),
    .A1(_00167_),
    .S(_06392_),
    .X(_06394_));
 sg13g2_nand2_1 _24073_ (.Y(_06395_),
    .A(_05497_),
    .B(_06390_));
 sg13g2_mux2_1 _24074_ (.A0(\atari2600.tia.p9_l ),
    .A1(_06394_),
    .S(_06393_),
    .X(_06396_));
 sg13g2_mux2_1 _24075_ (.A0(\atari2600.tia.p4_l ),
    .A1(_06396_),
    .S(_06395_),
    .X(_06397_));
 sg13g2_or2_1 _24076_ (.X(_06398_),
    .B(_06397_),
    .A(_05502_));
 sg13g2_o21ai_1 _24077_ (.B1(net6022),
    .Y(_06399_),
    .A1(_06389_),
    .A2(_06398_));
 sg13g2_a21oi_1 _24078_ (.A1(_08031_),
    .A2(_06389_),
    .Y(_02044_),
    .B1(_06399_));
 sg13g2_nor2_1 _24079_ (.A(_08163_),
    .B(_06339_),
    .Y(_06400_));
 sg13g2_nor3_1 _24080_ (.A(_07963_),
    .B(net5583),
    .C(\atari2600.tia.audc1[1] ),
    .Y(_06401_));
 sg13g2_nor3_1 _24081_ (.A(\atari2600.tia.audc1[3] ),
    .B(_07965_),
    .C(_07966_),
    .Y(_06402_));
 sg13g2_a22oi_1 _24082_ (.Y(_06403_),
    .B1(_06402_),
    .B2(net5583),
    .A2(_06401_),
    .A1(\atari2600.tia.audc1[0] ));
 sg13g2_a221oi_1 _24083_ (.B2(net5583),
    .C1(_00166_),
    .B1(_06402_),
    .A1(_07965_),
    .Y(_06404_),
    .A2(_05958_));
 sg13g2_nor2_1 _24084_ (.A(\atari2600.tia.p9_r ),
    .B(\atari2600.tia.audc1[0] ),
    .Y(_06405_));
 sg13g2_a22oi_1 _24085_ (.Y(_06406_),
    .B1(_06401_),
    .B2(_06405_),
    .A2(_05961_),
    .A1(\atari2600.tia.audc1[0] ));
 sg13g2_o21ai_1 _24086_ (.B1(_06406_),
    .Y(_06407_),
    .A1(\atari2600.tia.p5_r ),
    .A2(_06403_));
 sg13g2_nand3_1 _24087_ (.B(\atari2600.tia.audc1[0] ),
    .C(_05961_),
    .A(\atari2600.tia.p4_r ),
    .Y(_06408_));
 sg13g2_o21ai_1 _24088_ (.B1(_06408_),
    .Y(_06409_),
    .A1(_06404_),
    .A2(_06407_));
 sg13g2_nor2_1 _24089_ (.A(_05962_),
    .B(_06409_),
    .Y(_06410_));
 sg13g2_o21ai_1 _24090_ (.B1(net6035),
    .Y(_06411_),
    .A1(net5833),
    .A2(_06400_));
 sg13g2_a21oi_1 _24091_ (.A1(_06400_),
    .A2(_06410_),
    .Y(_02045_),
    .B1(_06411_));
 sg13g2_o21ai_1 _24092_ (.B1(net6931),
    .Y(_06412_),
    .A1(_10252_),
    .A2(_10254_));
 sg13g2_a21oi_1 _24093_ (.A1(_10256_),
    .A2(_06412_),
    .Y(_02046_),
    .B1(net5993));
 sg13g2_nor3_2 _24094_ (.A(_08632_),
    .B(net5230),
    .C(_05258_),
    .Y(_06413_));
 sg13g2_a21oi_1 _24095_ (.A1(_08636_),
    .A2(_05257_),
    .Y(_06414_),
    .B1(net3083));
 sg13g2_nor3_1 _24096_ (.A(net5989),
    .B(_06413_),
    .C(_06414_),
    .Y(_02047_));
 sg13g2_a21oi_1 _24097_ (.A1(_08636_),
    .A2(_05260_),
    .Y(_06415_),
    .B1(net7364));
 sg13g2_and3_2 _24098_ (.X(_06416_),
    .A(_10184_),
    .B(_10201_),
    .C(net5424));
 sg13g2_nor3_1 _24099_ (.A(net5984),
    .B(_06415_),
    .C(_06416_),
    .Y(_02048_));
 sg13g2_nor4_2 _24100_ (.A(net5029),
    .B(net4948),
    .C(_04814_),
    .Y(_06417_),
    .D(_05351_));
 sg13g2_nor2_1 _24101_ (.A(net3244),
    .B(_06417_),
    .Y(_06418_));
 sg13g2_a21oi_1 _24102_ (.A1(net5132),
    .A2(_06417_),
    .Y(_02049_),
    .B1(_06418_));
 sg13g2_nor2_1 _24103_ (.A(net3086),
    .B(_06417_),
    .Y(_06419_));
 sg13g2_a21oi_1 _24104_ (.A1(net5178),
    .A2(_06417_),
    .Y(_02050_),
    .B1(_06419_));
 sg13g2_nor2_1 _24105_ (.A(net3845),
    .B(_06417_),
    .Y(_06420_));
 sg13g2_a21oi_1 _24106_ (.A1(net5147),
    .A2(_06417_),
    .Y(_02051_),
    .B1(_06420_));
 sg13g2_nand2_2 _24107_ (.Y(_06421_),
    .A(net4911),
    .B(_08741_));
 sg13g2_nor2_1 _24108_ (.A(_08632_),
    .B(_06421_),
    .Y(_06422_));
 sg13g2_o21ai_1 _24109_ (.B1(net6021),
    .Y(_06423_),
    .A1(net7059),
    .A2(net4667));
 sg13g2_a21oi_1 _24110_ (.A1(net5243),
    .A2(net4667),
    .Y(_02052_),
    .B1(_06423_));
 sg13g2_o21ai_1 _24111_ (.B1(net6020),
    .Y(_06424_),
    .A1(net6987),
    .A2(net4666));
 sg13g2_a21oi_1 _24112_ (.A1(net5139),
    .A2(net4667),
    .Y(_02053_),
    .B1(_06424_));
 sg13g2_o21ai_1 _24113_ (.B1(net6018),
    .Y(_06425_),
    .A1(net6978),
    .A2(net4667));
 sg13g2_a21oi_1 _24114_ (.A1(net5111),
    .A2(net4667),
    .Y(_02054_),
    .B1(_06425_));
 sg13g2_o21ai_1 _24115_ (.B1(net6013),
    .Y(_06426_),
    .A1(net6982),
    .A2(net4667));
 sg13g2_a21oi_1 _24116_ (.A1(net5179),
    .A2(net4666),
    .Y(_02055_),
    .B1(_06426_));
 sg13g2_o21ai_1 _24117_ (.B1(net6013),
    .Y(_06427_),
    .A1(net7014),
    .A2(net4666));
 sg13g2_a21oi_1 _24118_ (.A1(net5155),
    .A2(net4666),
    .Y(_02056_),
    .B1(_06427_));
 sg13g2_o21ai_1 _24119_ (.B1(net6019),
    .Y(_06428_),
    .A1(net7076),
    .A2(net4666));
 sg13g2_a21oi_1 _24120_ (.A1(net5085),
    .A2(net4666),
    .Y(_02057_),
    .B1(_06428_));
 sg13g2_o21ai_1 _24121_ (.B1(net6019),
    .Y(_06429_),
    .A1(net7043),
    .A2(net4666));
 sg13g2_a21oi_1 _24122_ (.A1(net5062),
    .A2(net4666),
    .Y(_02058_),
    .B1(_06429_));
 sg13g2_nor2_2 _24123_ (.A(net5015),
    .B(_08735_),
    .Y(_06430_));
 sg13g2_nand2_2 _24124_ (.Y(_06431_),
    .A(_08581_),
    .B(net4816));
 sg13g2_nor2_1 _24125_ (.A(net4751),
    .B(_06431_),
    .Y(_06432_));
 sg13g2_nand3_1 _24126_ (.B(_08631_),
    .C(_06430_),
    .A(_08605_),
    .Y(_06433_));
 sg13g2_nor2_1 _24127_ (.A(_08637_),
    .B(_06431_),
    .Y(_06434_));
 sg13g2_o21ai_1 _24128_ (.B1(net6019),
    .Y(_06435_),
    .A1(net5232),
    .A2(net4729));
 sg13g2_a21oi_1 _24129_ (.A1(_08030_),
    .A2(net4729),
    .Y(_02059_),
    .B1(_06435_));
 sg13g2_o21ai_1 _24130_ (.B1(net6019),
    .Y(_06436_),
    .A1(net5129),
    .A2(_06433_));
 sg13g2_a21oi_1 _24131_ (.A1(_08029_),
    .A2(_06433_),
    .Y(_02060_),
    .B1(_06436_));
 sg13g2_o21ai_1 _24132_ (.B1(net6019),
    .Y(_06437_),
    .A1(net5101),
    .A2(net4729));
 sg13g2_a21oi_1 _24133_ (.A1(_08028_),
    .A2(net4729),
    .Y(_02061_),
    .B1(_06437_));
 sg13g2_o21ai_1 _24134_ (.B1(net6013),
    .Y(_06438_),
    .A1(net7192),
    .A2(_06434_));
 sg13g2_a21oi_1 _24135_ (.A1(net5184),
    .A2(_06434_),
    .Y(_02062_),
    .B1(_06438_));
 sg13g2_o21ai_1 _24136_ (.B1(net6012),
    .Y(_06439_),
    .A1(net7217),
    .A2(_06434_));
 sg13g2_a21oi_1 _24137_ (.A1(net5151),
    .A2(_06432_),
    .Y(_02063_),
    .B1(_06439_));
 sg13g2_o21ai_1 _24138_ (.B1(net6018),
    .Y(_06440_),
    .A1(net5075),
    .A2(net4729));
 sg13g2_a21oi_1 _24139_ (.A1(_08025_),
    .A2(net4729),
    .Y(_02064_),
    .B1(_06440_));
 sg13g2_o21ai_1 _24140_ (.B1(net6018),
    .Y(_06441_),
    .A1(net5054),
    .A2(net4729));
 sg13g2_a21oi_1 _24141_ (.A1(_08024_),
    .A2(net4729),
    .Y(_02065_),
    .B1(_06441_));
 sg13g2_nor2_2 _24142_ (.A(net5016),
    .B(net4948),
    .Y(_06442_));
 sg13g2_nand2_1 _24143_ (.Y(_06443_),
    .A(_08581_),
    .B(net4862));
 sg13g2_nor2_1 _24144_ (.A(net4751),
    .B(_06443_),
    .Y(_06444_));
 sg13g2_nor2_1 _24145_ (.A(_08637_),
    .B(_06443_),
    .Y(_06445_));
 sg13g2_nand2_2 _24146_ (.Y(_06446_),
    .A(_08636_),
    .B(_06442_));
 sg13g2_o21ai_1 _24147_ (.B1(net6021),
    .Y(_06447_),
    .A1(net5232),
    .A2(_06446_));
 sg13g2_a21oi_1 _24148_ (.A1(_08023_),
    .A2(_06446_),
    .Y(_02066_),
    .B1(_06447_));
 sg13g2_o21ai_1 _24149_ (.B1(net6012),
    .Y(_06448_),
    .A1(net7205),
    .A2(_06445_));
 sg13g2_a21oi_1 _24150_ (.A1(net5135),
    .A2(_06444_),
    .Y(_02067_),
    .B1(_06448_));
 sg13g2_o21ai_1 _24151_ (.B1(net6017),
    .Y(_06449_),
    .A1(net5101),
    .A2(_06446_));
 sg13g2_a21oi_1 _24152_ (.A1(_08022_),
    .A2(_06446_),
    .Y(_02068_),
    .B1(_06449_));
 sg13g2_o21ai_1 _24153_ (.B1(net6012),
    .Y(_06450_),
    .A1(net7186),
    .A2(_06445_));
 sg13g2_a21oi_1 _24154_ (.A1(net5179),
    .A2(_06444_),
    .Y(_02069_),
    .B1(_06450_));
 sg13g2_o21ai_1 _24155_ (.B1(net6012),
    .Y(_06451_),
    .A1(net7158),
    .A2(_06445_));
 sg13g2_a21oi_1 _24156_ (.A1(net5155),
    .A2(_06444_),
    .Y(_02070_),
    .B1(_06451_));
 sg13g2_o21ai_1 _24157_ (.B1(net6017),
    .Y(_06452_),
    .A1(net5075),
    .A2(_06446_));
 sg13g2_a21oi_1 _24158_ (.A1(_08019_),
    .A2(_06446_),
    .Y(_02071_),
    .B1(_06452_));
 sg13g2_o21ai_1 _24159_ (.B1(net6017),
    .Y(_06453_),
    .A1(net5054),
    .A2(_06446_));
 sg13g2_a21oi_1 _24160_ (.A1(_08018_),
    .A2(_06446_),
    .Y(_02072_),
    .B1(_06453_));
 sg13g2_nor2_2 _24161_ (.A(_08676_),
    .B(net4945),
    .Y(_06454_));
 sg13g2_nand2_2 _24162_ (.Y(_06455_),
    .A(net4992),
    .B(_08741_));
 sg13g2_nor2_1 _24163_ (.A(net4751),
    .B(_06455_),
    .Y(_06456_));
 sg13g2_o21ai_1 _24164_ (.B1(net6020),
    .Y(_06457_),
    .A1(net7116),
    .A2(net4665));
 sg13g2_a21oi_1 _24165_ (.A1(net5243),
    .A2(net4665),
    .Y(_02073_),
    .B1(_06457_));
 sg13g2_o21ai_1 _24166_ (.B1(net6020),
    .Y(_06458_),
    .A1(net7092),
    .A2(net4665));
 sg13g2_a21oi_1 _24167_ (.A1(net5135),
    .A2(net4665),
    .Y(_02074_),
    .B1(_06458_));
 sg13g2_o21ai_1 _24168_ (.B1(net6019),
    .Y(_06459_),
    .A1(net7164),
    .A2(net4664));
 sg13g2_a21oi_1 _24169_ (.A1(net5111),
    .A2(net4664),
    .Y(_02075_),
    .B1(_06459_));
 sg13g2_o21ai_1 _24170_ (.B1(net6013),
    .Y(_06460_),
    .A1(net7097),
    .A2(net4665));
 sg13g2_a21oi_1 _24171_ (.A1(net5184),
    .A2(net4665),
    .Y(_02076_),
    .B1(_06460_));
 sg13g2_o21ai_1 _24172_ (.B1(net6019),
    .Y(_06461_),
    .A1(net7157),
    .A2(net4664));
 sg13g2_a21oi_1 _24173_ (.A1(net5155),
    .A2(net4664),
    .Y(_02077_),
    .B1(_06461_));
 sg13g2_o21ai_1 _24174_ (.B1(net6020),
    .Y(_06462_),
    .A1(net7233),
    .A2(net4664));
 sg13g2_a21oi_1 _24175_ (.A1(net5085),
    .A2(net4664),
    .Y(_02078_),
    .B1(_06462_));
 sg13g2_o21ai_1 _24176_ (.B1(net6019),
    .Y(_06463_),
    .A1(net7190),
    .A2(net4664));
 sg13g2_a21oi_1 _24177_ (.A1(net5062),
    .A2(net4664),
    .Y(_02079_),
    .B1(_06463_));
 sg13g2_nor3_1 _24178_ (.A(_08565_),
    .B(net4955),
    .C(_05394_),
    .Y(_06464_));
 sg13g2_o21ai_1 _24179_ (.B1(net6010),
    .Y(_06465_),
    .A1(net7169),
    .A2(_06464_));
 sg13g2_a21oi_1 _24180_ (.A1(net5238),
    .A2(_06464_),
    .Y(_02080_),
    .B1(_06465_));
 sg13g2_nor3_1 _24181_ (.A(net4955),
    .B(_08735_),
    .C(_05394_),
    .Y(_06466_));
 sg13g2_o21ai_1 _24182_ (.B1(net6010),
    .Y(_06467_),
    .A1(net7232),
    .A2(_06466_));
 sg13g2_a21oi_1 _24183_ (.A1(net5238),
    .A2(_06466_),
    .Y(_02081_),
    .B1(_06467_));
 sg13g2_nor3_1 _24184_ (.A(net4955),
    .B(net4948),
    .C(_05394_),
    .Y(_06468_));
 sg13g2_o21ai_1 _24185_ (.B1(net6010),
    .Y(_06469_),
    .A1(net7239),
    .A2(_06468_));
 sg13g2_a21oi_1 _24186_ (.A1(net5238),
    .A2(_06468_),
    .Y(_02082_),
    .B1(_06469_));
 sg13g2_nand2_2 _24187_ (.Y(_06470_),
    .A(net5422),
    .B(_03118_));
 sg13g2_mux2_1 _24188_ (.A0(net5781),
    .A1(net6875),
    .S(_06470_),
    .X(_02083_));
 sg13g2_mux2_1 _24189_ (.A0(net5752),
    .A1(net6259),
    .S(_06470_),
    .X(_02084_));
 sg13g2_mux2_1 _24190_ (.A0(net5722),
    .A1(net6465),
    .S(_06470_),
    .X(_02085_));
 sg13g2_mux2_1 _24191_ (.A0(net5693),
    .A1(net6115),
    .S(_06470_),
    .X(_02086_));
 sg13g2_mux2_1 _24192_ (.A0(net5665),
    .A1(net6070),
    .S(_06470_),
    .X(_02087_));
 sg13g2_mux2_1 _24193_ (.A0(net5638),
    .A1(net4350),
    .S(_06470_),
    .X(_02088_));
 sg13g2_mux2_1 _24194_ (.A0(net5607),
    .A1(net6988),
    .S(_06470_),
    .X(_02089_));
 sg13g2_nor2_2 _24195_ (.A(_08606_),
    .B(net4771),
    .Y(_06471_));
 sg13g2_nand2_2 _24196_ (.Y(_06472_),
    .A(_08605_),
    .B(_08782_));
 sg13g2_nor3_1 _24197_ (.A(_08584_),
    .B(net5257),
    .C(_06472_),
    .Y(_06473_));
 sg13g2_a21oi_1 _24198_ (.A1(_08583_),
    .A2(_06471_),
    .Y(_06474_),
    .B1(net7292));
 sg13g2_nor3_1 _24199_ (.A(net5984),
    .B(_06473_),
    .C(_06474_),
    .Y(_02090_));
 sg13g2_nor2_2 _24200_ (.A(_06431_),
    .B(_06472_),
    .Y(_06475_));
 sg13g2_o21ai_1 _24201_ (.B1(net6005),
    .Y(_06476_),
    .A1(net7288),
    .A2(_06475_));
 sg13g2_a21oi_1 _24202_ (.A1(net5264),
    .A2(_06475_),
    .Y(_02091_),
    .B1(_06476_));
 sg13g2_nor2_1 _24203_ (.A(net4751),
    .B(_05392_),
    .Y(_06477_));
 sg13g2_o21ai_1 _24204_ (.B1(net6010),
    .Y(_06478_),
    .A1(net6138),
    .A2(_06477_));
 sg13g2_a21oi_1 _24205_ (.A1(net5107),
    .A2(_06477_),
    .Y(_02092_),
    .B1(_06478_));
 sg13g2_nor2_2 _24206_ (.A(_08676_),
    .B(net4954),
    .Y(_06479_));
 sg13g2_nor2b_1 _24207_ (.A(net4751),
    .B_N(_06479_),
    .Y(_06480_));
 sg13g2_o21ai_1 _24208_ (.B1(net6004),
    .Y(_06481_),
    .A1(net4105),
    .A2(_06480_));
 sg13g2_a21oi_1 _24209_ (.A1(net5107),
    .A2(_06480_),
    .Y(_02093_),
    .B1(_06481_));
 sg13g2_o21ai_1 _24210_ (.B1(net6032),
    .Y(_06482_),
    .A1(net5257),
    .A2(net4730));
 sg13g2_a21oi_1 _24211_ (.A1(_08010_),
    .A2(net4730),
    .Y(_02094_),
    .B1(_06482_));
 sg13g2_o21ai_1 _24212_ (.B1(net6009),
    .Y(_06483_),
    .A1(net5230),
    .A2(net4730));
 sg13g2_a21oi_1 _24213_ (.A1(net5565),
    .A2(net4730),
    .Y(_02095_),
    .B1(_06483_));
 sg13g2_o21ai_1 _24214_ (.B1(net6033),
    .Y(_06484_),
    .A1(net5130),
    .A2(net4730));
 sg13g2_a21oi_1 _24215_ (.A1(_08008_),
    .A2(net4730),
    .Y(_02096_),
    .B1(_06484_));
 sg13g2_o21ai_1 _24216_ (.B1(net6016),
    .Y(_06485_),
    .A1(net7093),
    .A2(net4731));
 sg13g2_a21oi_1 _24217_ (.A1(net5265),
    .A2(net4731),
    .Y(_02097_),
    .B1(_06485_));
 sg13g2_o21ai_1 _24218_ (.B1(net6016),
    .Y(_06486_),
    .A1(net5229),
    .A2(_05399_));
 sg13g2_a21oi_1 _24219_ (.A1(_08007_),
    .A2(_05399_),
    .Y(_02098_),
    .B1(_06486_));
 sg13g2_o21ai_1 _24220_ (.B1(net6004),
    .Y(_06487_),
    .A1(net7171),
    .A2(net4731));
 sg13g2_a21oi_1 _24221_ (.A1(net5136),
    .A2(net4731),
    .Y(_02099_),
    .B1(_06487_));
 sg13g2_o21ai_1 _24222_ (.B1(net6010),
    .Y(_06488_),
    .A1(net7183),
    .A2(net4731));
 sg13g2_a21oi_1 _24223_ (.A1(net5107),
    .A2(net4731),
    .Y(_02100_),
    .B1(_06488_));
 sg13g2_o21ai_1 _24224_ (.B1(net6010),
    .Y(_06489_),
    .A1(net7098),
    .A2(_05398_));
 sg13g2_a21oi_1 _24225_ (.A1(net5179),
    .A2(_05395_),
    .Y(_02101_),
    .B1(_06489_));
 sg13g2_o21ai_1 _24226_ (.B1(net6010),
    .Y(_06490_),
    .A1(net7131),
    .A2(net4731));
 sg13g2_a21oi_1 _24227_ (.A1(net5151),
    .A2(_05395_),
    .Y(_02102_),
    .B1(_06490_));
 sg13g2_o21ai_1 _24228_ (.B1(net6016),
    .Y(_06491_),
    .A1(net5073),
    .A2(_05399_));
 sg13g2_a21oi_1 _24229_ (.A1(_08006_),
    .A2(_05399_),
    .Y(_02103_),
    .B1(_06491_));
 sg13g2_o21ai_1 _24230_ (.B1(net6016),
    .Y(_06492_),
    .A1(net7108),
    .A2(_05398_));
 sg13g2_a21oi_1 _24231_ (.A1(net5059),
    .A2(_05398_),
    .Y(_02104_),
    .B1(_06492_));
 sg13g2_and2_2 _24232_ (.A(_05393_),
    .B(_06479_),
    .X(_06493_));
 sg13g2_and2_1 _24233_ (.A(_05396_),
    .B(_06479_),
    .X(_06494_));
 sg13g2_nand2_1 _24234_ (.Y(_06495_),
    .A(_05396_),
    .B(_06479_));
 sg13g2_o21ai_1 _24235_ (.B1(net6003),
    .Y(_06496_),
    .A1(net5257),
    .A2(net4727));
 sg13g2_a21oi_1 _24236_ (.A1(_08005_),
    .A2(net4727),
    .Y(_02105_),
    .B1(_06496_));
 sg13g2_o21ai_1 _24237_ (.B1(net6003),
    .Y(_06497_),
    .A1(net5228),
    .A2(net4727));
 sg13g2_a21oi_1 _24238_ (.A1(_08004_),
    .A2(net4727),
    .Y(_02106_),
    .B1(_06497_));
 sg13g2_o21ai_1 _24239_ (.B1(net6003),
    .Y(_06498_),
    .A1(net5129),
    .A2(net4727));
 sg13g2_a21oi_1 _24240_ (.A1(_08003_),
    .A2(net4727),
    .Y(_02107_),
    .B1(_06498_));
 sg13g2_o21ai_1 _24241_ (.B1(net6003),
    .Y(_06499_),
    .A1(net5102),
    .A2(net4727));
 sg13g2_a21oi_1 _24242_ (.A1(_08002_),
    .A2(net4727),
    .Y(_02108_),
    .B1(_06499_));
 sg13g2_o21ai_1 _24243_ (.B1(net6004),
    .Y(_06500_),
    .A1(net4317),
    .A2(_06494_));
 sg13g2_a21oi_1 _24244_ (.A1(net5179),
    .A2(_06493_),
    .Y(_02109_),
    .B1(_06500_));
 sg13g2_o21ai_1 _24245_ (.B1(net6004),
    .Y(_06501_),
    .A1(net7106),
    .A2(_06494_));
 sg13g2_a21oi_1 _24246_ (.A1(net5151),
    .A2(_06493_),
    .Y(_02110_),
    .B1(_06501_));
 sg13g2_o21ai_1 _24247_ (.B1(net6004),
    .Y(_06502_),
    .A1(net5072),
    .A2(net4728));
 sg13g2_a21oi_1 _24248_ (.A1(_08001_),
    .A2(net4728),
    .Y(_02111_),
    .B1(_06502_));
 sg13g2_o21ai_1 _24249_ (.B1(net6003),
    .Y(_06503_),
    .A1(net5050),
    .A2(net4728));
 sg13g2_a21oi_1 _24250_ (.A1(_08000_),
    .A2(net4728),
    .Y(_02112_),
    .B1(_06503_));
 sg13g2_nand2_1 _24251_ (.Y(_06504_),
    .A(\atari2600.tia.colup0[0] ),
    .B(_10210_));
 sg13g2_a21oi_1 _24252_ (.A1(\atari2600.tia.colup1[0] ),
    .A2(_10211_),
    .Y(_06505_),
    .B1(net5565));
 sg13g2_a22oi_1 _24253_ (.Y(_06506_),
    .B1(_06504_),
    .B2(_06505_),
    .A2(_08017_),
    .A1(net5566));
 sg13g2_mux2_1 _24254_ (.A0(\atari2600.tia.colubk[0] ),
    .A1(_06506_),
    .S(net5114),
    .X(_06507_));
 sg13g2_a21oi_1 _24255_ (.A1(_09820_),
    .A2(_06507_),
    .Y(_06508_),
    .B1(net4583));
 sg13g2_o21ai_1 _24256_ (.B1(_06508_),
    .Y(_06509_),
    .A1(_08023_),
    .A2(net4769));
 sg13g2_and2_1 _24257_ (.A(\atari2600.tia.pf_priority ),
    .B(net5114),
    .X(_06510_));
 sg13g2_a21oi_1 _24258_ (.A1(_08030_),
    .A2(net4582),
    .Y(_06511_),
    .B1(net5019));
 sg13g2_nand2_1 _24259_ (.Y(_06512_),
    .A(_06509_),
    .B(_06511_));
 sg13g2_a21oi_1 _24260_ (.A1(_06506_),
    .A2(net5019),
    .Y(_06513_),
    .B1(net4767));
 sg13g2_o21ai_1 _24261_ (.B1(net4783),
    .Y(_06514_),
    .A1(\atari2600.tia.colup1[0] ),
    .A2(_10052_));
 sg13g2_a21oi_1 _24262_ (.A1(_06512_),
    .A2(_06513_),
    .Y(_06515_),
    .B1(_06514_));
 sg13g2_a21oi_1 _24263_ (.A1(\atari2600.tia.vid_ypos[2] ),
    .A2(\atari2600.tia.vid_ypos[1] ),
    .Y(_06516_),
    .B1(\atari2600.tia.vid_ypos[3] ));
 sg13g2_nand2b_1 _24264_ (.Y(_06517_),
    .B(\atari2600.tia.vid_ypos[4] ),
    .A_N(_06516_));
 sg13g2_and4_1 _24265_ (.A(_08043_),
    .B(_00143_),
    .C(_08139_),
    .D(_06517_),
    .X(_06518_));
 sg13g2_nor3_2 _24266_ (.A(_09827_),
    .B(net5474),
    .C(_06518_),
    .Y(_06519_));
 sg13g2_nand3b_1 _24267_ (.B(net5511),
    .C(_09826_),
    .Y(_06520_),
    .A_N(_06518_));
 sg13g2_nand2_1 _24268_ (.Y(_06521_),
    .A(net5779),
    .B(_06520_));
 sg13g2_o21ai_1 _24269_ (.B1(net4764),
    .Y(_06522_),
    .A1(_08030_),
    .A2(net4782));
 sg13g2_nor2_1 _24270_ (.A(_06515_),
    .B(_06522_),
    .Y(_06523_));
 sg13g2_o21ai_1 _24271_ (.B1(_06519_),
    .Y(_06524_),
    .A1(net7116),
    .A2(net4764));
 sg13g2_o21ai_1 _24272_ (.B1(_06521_),
    .Y(_02113_),
    .A1(_06523_),
    .A2(_06524_));
 sg13g2_nand2_1 _24273_ (.Y(_06525_),
    .A(\atari2600.tia.colup0[1] ),
    .B(net5511));
 sg13g2_a21oi_1 _24274_ (.A1(\atari2600.tia.colup1[1] ),
    .A2(net5474),
    .Y(_06526_),
    .B1(net5566));
 sg13g2_a22oi_1 _24275_ (.Y(_06527_),
    .B1(_06525_),
    .B2(_06526_),
    .A2(_08016_),
    .A1(net5566));
 sg13g2_mux2_1 _24276_ (.A0(\atari2600.tia.colubk[1] ),
    .A1(_06527_),
    .S(net5114),
    .X(_06528_));
 sg13g2_nand2_1 _24277_ (.Y(_06529_),
    .A(\atari2600.tia.colup1[1] ),
    .B(_09821_));
 sg13g2_a21oi_1 _24278_ (.A1(net4769),
    .A2(_06528_),
    .Y(_06530_),
    .B1(net4582));
 sg13g2_a221oi_1 _24279_ (.B2(_06530_),
    .C1(net5018),
    .B1(_06529_),
    .A1(_08029_),
    .Y(_06531_),
    .A2(net4582));
 sg13g2_a21oi_1 _24280_ (.A1(net5018),
    .A2(_06527_),
    .Y(_06532_),
    .B1(_06531_));
 sg13g2_nand2_1 _24281_ (.Y(_06533_),
    .A(\atari2600.tia.colup1[1] ),
    .B(net4767));
 sg13g2_o21ai_1 _24282_ (.B1(_06533_),
    .Y(_06534_),
    .A1(net4767),
    .A2(_06532_));
 sg13g2_mux2_1 _24283_ (.A0(\atari2600.tia.colup0[1] ),
    .A1(_06534_),
    .S(net4782),
    .X(_06535_));
 sg13g2_inv_1 _24284_ (.Y(_06536_),
    .A(_06535_));
 sg13g2_o21ai_1 _24285_ (.B1(_06519_),
    .Y(_06537_),
    .A1(net7092),
    .A2(net4765));
 sg13g2_a21oi_1 _24286_ (.A1(net4765),
    .A2(_06536_),
    .Y(_06538_),
    .B1(_06537_));
 sg13g2_a21o_1 _24287_ (.A2(_06520_),
    .A1(net5744),
    .B1(_06538_),
    .X(_02114_));
 sg13g2_nand2_1 _24288_ (.Y(_06539_),
    .A(\atari2600.tia.colup0[2] ),
    .B(net5511));
 sg13g2_a21oi_1 _24289_ (.A1(\atari2600.tia.colup1[2] ),
    .A2(net5474),
    .Y(_06540_),
    .B1(net5565));
 sg13g2_a22oi_1 _24290_ (.Y(_06541_),
    .B1(_06539_),
    .B2(_06540_),
    .A2(_08015_),
    .A1(net5565));
 sg13g2_mux2_1 _24291_ (.A0(\atari2600.tia.colubk[2] ),
    .A1(_06541_),
    .S(net5114),
    .X(_06542_));
 sg13g2_a21oi_1 _24292_ (.A1(net4770),
    .A2(_06542_),
    .Y(_06543_),
    .B1(net4583));
 sg13g2_o21ai_1 _24293_ (.B1(_06543_),
    .Y(_06544_),
    .A1(_08022_),
    .A2(net4770));
 sg13g2_a21oi_1 _24294_ (.A1(_08028_),
    .A2(net4583),
    .Y(_06545_),
    .B1(net5019));
 sg13g2_a22oi_1 _24295_ (.Y(_06546_),
    .B1(_06544_),
    .B2(_06545_),
    .A2(_06541_),
    .A1(net5019));
 sg13g2_nor2_1 _24296_ (.A(_10051_),
    .B(_06546_),
    .Y(_06547_));
 sg13g2_a21oi_1 _24297_ (.A1(\atari2600.tia.colup1[2] ),
    .A2(net4767),
    .Y(_06548_),
    .B1(_06547_));
 sg13g2_nand2_1 _24298_ (.Y(_06549_),
    .A(net4783),
    .B(_06548_));
 sg13g2_o21ai_1 _24299_ (.B1(_06549_),
    .Y(_06550_),
    .A1(\atari2600.tia.colup0[2] ),
    .A2(net4783));
 sg13g2_o21ai_1 _24300_ (.B1(_06519_),
    .Y(_06551_),
    .A1(net7164),
    .A2(net4764));
 sg13g2_a21oi_1 _24301_ (.A1(net4764),
    .A2(_06550_),
    .Y(_06552_),
    .B1(_06551_));
 sg13g2_a21o_1 _24302_ (.A2(_06520_),
    .A1(net5714),
    .B1(_06552_),
    .X(_02115_));
 sg13g2_nand2_1 _24303_ (.Y(_06553_),
    .A(\atari2600.tia.colup0[3] ),
    .B(net5511));
 sg13g2_a21oi_1 _24304_ (.A1(\atari2600.tia.colup1[3] ),
    .A2(net5474),
    .Y(_06554_),
    .B1(net5566));
 sg13g2_a22oi_1 _24305_ (.Y(_06555_),
    .B1(_06553_),
    .B2(_06554_),
    .A2(_08014_),
    .A1(net5566));
 sg13g2_mux2_1 _24306_ (.A0(\atari2600.tia.colubk[3] ),
    .A1(_06555_),
    .S(net5114),
    .X(_06556_));
 sg13g2_a21oi_1 _24307_ (.A1(net4769),
    .A2(_06556_),
    .Y(_06557_),
    .B1(net4582));
 sg13g2_o21ai_1 _24308_ (.B1(_06557_),
    .Y(_06558_),
    .A1(_08021_),
    .A2(net4769));
 sg13g2_a21oi_1 _24309_ (.A1(_08027_),
    .A2(net4582),
    .Y(_06559_),
    .B1(net5018));
 sg13g2_a22oi_1 _24310_ (.Y(_06560_),
    .B1(_06558_),
    .B2(_06559_),
    .A2(_06555_),
    .A1(net5018));
 sg13g2_nor2_1 _24311_ (.A(net4767),
    .B(_06560_),
    .Y(_06561_));
 sg13g2_a21oi_1 _24312_ (.A1(\atari2600.tia.colup1[3] ),
    .A2(net4767),
    .Y(_06562_),
    .B1(_06561_));
 sg13g2_nand2_1 _24313_ (.Y(_06563_),
    .A(net4782),
    .B(_06562_));
 sg13g2_o21ai_1 _24314_ (.B1(_06563_),
    .Y(_06564_),
    .A1(\atari2600.tia.colup0[3] ),
    .A2(net4782));
 sg13g2_o21ai_1 _24315_ (.B1(_06519_),
    .Y(_06565_),
    .A1(net7097),
    .A2(net4765));
 sg13g2_a21oi_1 _24316_ (.A1(net4765),
    .A2(_06564_),
    .Y(_06566_),
    .B1(_06565_));
 sg13g2_a21o_1 _24317_ (.A2(_06520_),
    .A1(net5687),
    .B1(_06566_),
    .X(_02116_));
 sg13g2_nand2_1 _24318_ (.Y(_06567_),
    .A(\atari2600.tia.colup0[4] ),
    .B(net5511));
 sg13g2_a21oi_1 _24319_ (.A1(\atari2600.tia.colup1[4] ),
    .A2(net5474),
    .Y(_06568_),
    .B1(net5566));
 sg13g2_a22oi_1 _24320_ (.Y(_06569_),
    .B1(_06567_),
    .B2(_06568_),
    .A2(_08013_),
    .A1(net5566));
 sg13g2_mux2_1 _24321_ (.A0(\atari2600.tia.colubk[4] ),
    .A1(_06569_),
    .S(net5114),
    .X(_06570_));
 sg13g2_a21oi_1 _24322_ (.A1(net4769),
    .A2(_06570_),
    .Y(_06571_),
    .B1(net4582));
 sg13g2_o21ai_1 _24323_ (.B1(_06571_),
    .Y(_06572_),
    .A1(_08020_),
    .A2(net4769));
 sg13g2_a21oi_1 _24324_ (.A1(_08026_),
    .A2(net4582),
    .Y(_06573_),
    .B1(net5018));
 sg13g2_a22oi_1 _24325_ (.Y(_06574_),
    .B1(_06572_),
    .B2(_06573_),
    .A2(_06569_),
    .A1(net5018));
 sg13g2_nor2_1 _24326_ (.A(net4767),
    .B(_06574_),
    .Y(_06575_));
 sg13g2_a21oi_1 _24327_ (.A1(\atari2600.tia.colup1[4] ),
    .A2(net4767),
    .Y(_06576_),
    .B1(_06575_));
 sg13g2_nand2_1 _24328_ (.Y(_06577_),
    .A(net4782),
    .B(_06576_));
 sg13g2_o21ai_1 _24329_ (.B1(_06577_),
    .Y(_06578_),
    .A1(\atari2600.tia.colup0[4] ),
    .A2(net4782));
 sg13g2_o21ai_1 _24330_ (.B1(_06519_),
    .Y(_06579_),
    .A1(net7157),
    .A2(net4764));
 sg13g2_a21oi_1 _24331_ (.A1(net4764),
    .A2(_06578_),
    .Y(_06580_),
    .B1(_06579_));
 sg13g2_a21o_1 _24332_ (.A2(_06520_),
    .A1(net5657),
    .B1(_06580_),
    .X(_02117_));
 sg13g2_nand2_1 _24333_ (.Y(_06581_),
    .A(net5634),
    .B(_06520_));
 sg13g2_nand2_1 _24334_ (.Y(_06582_),
    .A(\atari2600.tia.colup0[5] ),
    .B(net5511));
 sg13g2_a21oi_1 _24335_ (.A1(\atari2600.tia.colup1[5] ),
    .A2(net5474),
    .Y(_06583_),
    .B1(net5565));
 sg13g2_a22oi_1 _24336_ (.Y(_06584_),
    .B1(_06582_),
    .B2(_06583_),
    .A2(_08012_),
    .A1(net5565));
 sg13g2_mux2_1 _24337_ (.A0(\atari2600.tia.colubk[5] ),
    .A1(_06584_),
    .S(net5114),
    .X(_06585_));
 sg13g2_nand2_1 _24338_ (.Y(_06586_),
    .A(net4769),
    .B(_06585_));
 sg13g2_o21ai_1 _24339_ (.B1(_06586_),
    .Y(_06587_),
    .A1(_08019_),
    .A2(net4769));
 sg13g2_a21oi_1 _24340_ (.A1(_08025_),
    .A2(net4583),
    .Y(_06588_),
    .B1(net5018));
 sg13g2_o21ai_1 _24341_ (.B1(_06588_),
    .Y(_06589_),
    .A1(net4582),
    .A2(_06587_));
 sg13g2_a21oi_1 _24342_ (.A1(net5019),
    .A2(_06584_),
    .Y(_06590_),
    .B1(net4768));
 sg13g2_o21ai_1 _24343_ (.B1(net4782),
    .Y(_06591_),
    .A1(\atari2600.tia.colup1[5] ),
    .A2(_10052_));
 sg13g2_a21oi_1 _24344_ (.A1(_06589_),
    .A2(_06590_),
    .Y(_06592_),
    .B1(_06591_));
 sg13g2_o21ai_1 _24345_ (.B1(net4766),
    .Y(_06593_),
    .A1(_08025_),
    .A2(net4783));
 sg13g2_nor2_1 _24346_ (.A(_06592_),
    .B(_06593_),
    .Y(_06594_));
 sg13g2_o21ai_1 _24347_ (.B1(_06519_),
    .Y(_06595_),
    .A1(net7233),
    .A2(net4764));
 sg13g2_o21ai_1 _24348_ (.B1(_06581_),
    .Y(_02118_),
    .A1(_06594_),
    .A2(_06595_));
 sg13g2_nand2_1 _24349_ (.Y(_06596_),
    .A(net5599),
    .B(_06520_));
 sg13g2_nand2_1 _24350_ (.Y(_06597_),
    .A(\atari2600.tia.colup0[6] ),
    .B(net5511));
 sg13g2_a21oi_1 _24351_ (.A1(\atari2600.tia.colup1[6] ),
    .A2(net5474),
    .Y(_06598_),
    .B1(net5565));
 sg13g2_a22oi_1 _24352_ (.Y(_06599_),
    .B1(_06597_),
    .B2(_06598_),
    .A2(_08011_),
    .A1(net5565));
 sg13g2_mux2_1 _24353_ (.A0(\atari2600.tia.colubk[6] ),
    .A1(_06599_),
    .S(net5114),
    .X(_06600_));
 sg13g2_nand2_1 _24354_ (.Y(_06601_),
    .A(net4770),
    .B(_06600_));
 sg13g2_o21ai_1 _24355_ (.B1(_06601_),
    .Y(_06602_),
    .A1(_08018_),
    .A2(net4770));
 sg13g2_a21oi_1 _24356_ (.A1(_08024_),
    .A2(net4583),
    .Y(_06603_),
    .B1(net5019));
 sg13g2_o21ai_1 _24357_ (.B1(_06603_),
    .Y(_06604_),
    .A1(net4583),
    .A2(_06602_));
 sg13g2_a21oi_1 _24358_ (.A1(net5018),
    .A2(_06599_),
    .Y(_06605_),
    .B1(net4768));
 sg13g2_o21ai_1 _24359_ (.B1(net4782),
    .Y(_06606_),
    .A1(\atari2600.tia.colup1[6] ),
    .A2(_10052_));
 sg13g2_a21oi_1 _24360_ (.A1(_06604_),
    .A2(_06605_),
    .Y(_06607_),
    .B1(_06606_));
 sg13g2_o21ai_1 _24361_ (.B1(net4766),
    .Y(_06608_),
    .A1(_08024_),
    .A2(net4783));
 sg13g2_nor2_1 _24362_ (.A(_06607_),
    .B(_06608_),
    .Y(_06609_));
 sg13g2_o21ai_1 _24363_ (.B1(_06519_),
    .Y(_06610_),
    .A1(net7190),
    .A2(net4764));
 sg13g2_o21ai_1 _24364_ (.B1(_06596_),
    .Y(_02119_),
    .A1(_06609_),
    .A2(_06610_));
 sg13g2_and3_1 _24365_ (.X(_06611_),
    .A(net6010),
    .B(net5354),
    .C(_06493_));
 sg13g2_mux2_1 _24366_ (.A0(net3461),
    .A1(\atari2600.tia.diag[104] ),
    .S(net4663),
    .X(_02120_));
 sg13g2_nor2_1 _24367_ (.A(\atari2600.tia.old_grp0[1] ),
    .B(net4663),
    .Y(_06612_));
 sg13g2_a21oi_1 _24368_ (.A1(_08007_),
    .A2(net4663),
    .Y(_02121_),
    .B1(_06612_));
 sg13g2_mux2_1 _24369_ (.A0(net3627),
    .A1(\atari2600.tia.diag[106] ),
    .S(net4663),
    .X(_02122_));
 sg13g2_mux2_1 _24370_ (.A0(net3201),
    .A1(\atari2600.tia.diag[107] ),
    .S(net4663),
    .X(_02123_));
 sg13g2_mux2_1 _24371_ (.A0(net3364),
    .A1(\atari2600.tia.diag[108] ),
    .S(net4663),
    .X(_02124_));
 sg13g2_mux2_1 _24372_ (.A0(net3218),
    .A1(\atari2600.tia.diag[109] ),
    .S(net4663),
    .X(_02125_));
 sg13g2_nor2_1 _24373_ (.A(net3239),
    .B(_06611_),
    .Y(_06613_));
 sg13g2_a21oi_1 _24374_ (.A1(_08006_),
    .A2(_06611_),
    .Y(_02126_),
    .B1(_06613_));
 sg13g2_mux2_1 _24375_ (.A0(net3271),
    .A1(\atari2600.tia.diag[111] ),
    .S(net4663),
    .X(_02127_));
 sg13g2_nor2_1 _24376_ (.A(_08676_),
    .B(net4934),
    .Y(_06614_));
 sg13g2_nand2_2 _24377_ (.Y(_06615_),
    .A(net4992),
    .B(_08746_));
 sg13g2_nor2_2 _24378_ (.A(net4771),
    .B(_05447_),
    .Y(_06616_));
 sg13g2_nand2_2 _24379_ (.Y(_06617_),
    .A(_08782_),
    .B(_05446_));
 sg13g2_nor2_1 _24380_ (.A(_08606_),
    .B(_06617_),
    .Y(_06618_));
 sg13g2_nand2_1 _24381_ (.Y(_06619_),
    .A(_08605_),
    .B(net4755));
 sg13g2_o21ai_1 _24382_ (.B1(_06619_),
    .Y(_06620_),
    .A1(_05394_),
    .A2(_06615_));
 sg13g2_o21ai_1 _24383_ (.B1(_06619_),
    .Y(_06621_),
    .A1(_05397_),
    .A2(_06615_));
 sg13g2_o21ai_1 _24384_ (.B1(net6006),
    .Y(_06622_),
    .A1(net7285),
    .A2(net4662));
 sg13g2_nand2_2 _24385_ (.Y(_06623_),
    .A(net5511),
    .B(_06617_));
 sg13g2_nor2_2 _24386_ (.A(net5829),
    .B(net4726),
    .Y(_06624_));
 sg13g2_nand2b_1 _24387_ (.Y(_06625_),
    .B(\atari2600.tia.hmp0[0] ),
    .A_N(\atari2600.tia.diag[64] ));
 sg13g2_xor2_1 _24388_ (.B(\atari2600.tia.diag[64] ),
    .A(net7162),
    .X(_06626_));
 sg13g2_a21oi_1 _24389_ (.A1(net4754),
    .A2(_06626_),
    .Y(_06627_),
    .B1(_06624_));
 sg13g2_a21oi_1 _24390_ (.A1(_06621_),
    .A2(_06627_),
    .Y(_02128_),
    .B1(_06622_));
 sg13g2_o21ai_1 _24391_ (.B1(net6006),
    .Y(_06628_),
    .A1(net7296),
    .A2(net4662));
 sg13g2_a21oi_2 _24392_ (.B1(net4726),
    .Y(_06629_),
    .A2(_10319_),
    .A1(_10317_));
 sg13g2_nor2_1 _24393_ (.A(\atari2600.tia.hmp0[1] ),
    .B(_07999_),
    .Y(_06630_));
 sg13g2_xnor2_1 _24394_ (.Y(_06631_),
    .A(\atari2600.tia.hmp0[1] ),
    .B(\atari2600.tia.diag[65] ));
 sg13g2_xor2_1 _24395_ (.B(_06631_),
    .A(_06625_),
    .X(_06632_));
 sg13g2_a21oi_1 _24396_ (.A1(net4754),
    .A2(_06632_),
    .Y(_06633_),
    .B1(_06629_));
 sg13g2_a21oi_1 _24397_ (.A1(_06621_),
    .A2(_06633_),
    .Y(_02129_),
    .B1(_06628_));
 sg13g2_o21ai_1 _24398_ (.B1(net6006),
    .Y(_06634_),
    .A1(net5596),
    .A2(net4662));
 sg13g2_nand2_1 _24399_ (.Y(_06635_),
    .A(net5561),
    .B(_10261_));
 sg13g2_a21oi_2 _24400_ (.B1(net4726),
    .Y(_06636_),
    .A2(_06635_),
    .A1(_10332_));
 sg13g2_xnor2_1 _24401_ (.Y(_06637_),
    .A(\atari2600.tia.hmp0[2] ),
    .B(net5596));
 sg13g2_a21oi_1 _24402_ (.A1(_06625_),
    .A2(_06631_),
    .Y(_06638_),
    .B1(_06630_));
 sg13g2_nor2b_1 _24403_ (.A(_06638_),
    .B_N(_06637_),
    .Y(_06639_));
 sg13g2_xor2_1 _24404_ (.B(_06638_),
    .A(_06637_),
    .X(_06640_));
 sg13g2_o21ai_1 _24405_ (.B1(net4662),
    .Y(_06641_),
    .A1(_06617_),
    .A2(_06640_));
 sg13g2_nor2_1 _24406_ (.A(_06636_),
    .B(_06641_),
    .Y(_06642_));
 sg13g2_nor2_1 _24407_ (.A(_06634_),
    .B(_06642_),
    .Y(_02130_));
 sg13g2_o21ai_1 _24408_ (.B1(net6004),
    .Y(_06643_),
    .A1(net5595),
    .A2(net4662));
 sg13g2_xnor2_1 _24409_ (.Y(_06644_),
    .A(net5821),
    .B(_10326_));
 sg13g2_nor2_2 _24410_ (.A(net4726),
    .B(_06644_),
    .Y(_06645_));
 sg13g2_xnor2_1 _24411_ (.Y(_06646_),
    .A(net5588),
    .B(net5595));
 sg13g2_a21oi_2 _24412_ (.B1(_06639_),
    .Y(_06647_),
    .A2(net5596),
    .A1(_07977_));
 sg13g2_nor2b_1 _24413_ (.A(_06647_),
    .B_N(_06646_),
    .Y(_06648_));
 sg13g2_xnor2_1 _24414_ (.Y(_06649_),
    .A(_06646_),
    .B(_06647_));
 sg13g2_a21oi_1 _24415_ (.A1(net4754),
    .A2(_06649_),
    .Y(_06650_),
    .B1(_06645_));
 sg13g2_a21oi_1 _24416_ (.A1(_06621_),
    .A2(_06650_),
    .Y(_02131_),
    .B1(_06643_));
 sg13g2_o21ai_1 _24417_ (.B1(net6004),
    .Y(_06651_),
    .A1(net5594),
    .A2(_06620_));
 sg13g2_and3_1 _24418_ (.X(_06652_),
    .A(net5821),
    .B(net5817),
    .C(_06635_));
 sg13g2_a21oi_1 _24419_ (.A1(net5821),
    .A2(_06635_),
    .Y(_06653_),
    .B1(net5817));
 sg13g2_nor3_2 _24420_ (.A(net4726),
    .B(_06652_),
    .C(_06653_),
    .Y(_06654_));
 sg13g2_xnor2_1 _24421_ (.Y(_06655_),
    .A(net5588),
    .B(net5594));
 sg13g2_a21oi_1 _24422_ (.A1(_07976_),
    .A2(net5595),
    .Y(_06656_),
    .B1(_06648_));
 sg13g2_nor2b_1 _24423_ (.A(_06656_),
    .B_N(_06655_),
    .Y(_06657_));
 sg13g2_xor2_1 _24424_ (.B(_06656_),
    .A(_06655_),
    .X(_06658_));
 sg13g2_o21ai_1 _24425_ (.B1(_06620_),
    .Y(_06659_),
    .A1(_06617_),
    .A2(_06658_));
 sg13g2_nor2_1 _24426_ (.A(_06654_),
    .B(_06659_),
    .Y(_06660_));
 sg13g2_nor2_1 _24427_ (.A(_06651_),
    .B(_06660_),
    .Y(_02132_));
 sg13g2_o21ai_1 _24428_ (.B1(net6014),
    .Y(_06661_),
    .A1(net5593),
    .A2(net4662));
 sg13g2_xor2_1 _24429_ (.B(_06652_),
    .A(net5809),
    .X(_06662_));
 sg13g2_nor2_2 _24430_ (.A(net4726),
    .B(_06662_),
    .Y(_06663_));
 sg13g2_a21oi_1 _24431_ (.A1(_07976_),
    .A2(net5594),
    .Y(_06664_),
    .B1(_06657_));
 sg13g2_nand2_1 _24432_ (.Y(_06665_),
    .A(\atari2600.tia.hmp0[3] ),
    .B(_07996_));
 sg13g2_xnor2_1 _24433_ (.Y(_06666_),
    .A(net5588),
    .B(net5593));
 sg13g2_xnor2_1 _24434_ (.Y(_06667_),
    .A(_06664_),
    .B(_06666_));
 sg13g2_a21oi_1 _24435_ (.A1(net4755),
    .A2(_06667_),
    .Y(_06668_),
    .B1(_06663_));
 sg13g2_a21oi_1 _24436_ (.A1(_06621_),
    .A2(_06668_),
    .Y(_02133_),
    .B1(_06661_));
 sg13g2_o21ai_1 _24437_ (.B1(net6014),
    .Y(_06669_),
    .A1(net7355),
    .A2(_06620_));
 sg13g2_nand2_1 _24438_ (.Y(_06670_),
    .A(net5812),
    .B(_06652_));
 sg13g2_or2_1 _24439_ (.X(_06671_),
    .B(_06670_),
    .A(net5803));
 sg13g2_a21oi_1 _24440_ (.A1(net5803),
    .A2(_06670_),
    .Y(_06672_),
    .B1(net4726));
 sg13g2_and2_2 _24441_ (.A(_06671_),
    .B(_06672_),
    .X(_06673_));
 sg13g2_xnor2_1 _24442_ (.Y(_06674_),
    .A(net5588),
    .B(\atari2600.tia.diag[70] ));
 sg13g2_o21ai_1 _24443_ (.B1(_06664_),
    .Y(_06675_),
    .A1(net5588),
    .A2(_07996_));
 sg13g2_a21oi_1 _24444_ (.A1(_06665_),
    .A2(_06675_),
    .Y(_06676_),
    .B1(_06674_));
 sg13g2_nand3_1 _24445_ (.B(_06674_),
    .C(_06675_),
    .A(_06665_),
    .Y(_06677_));
 sg13g2_nand2_1 _24446_ (.Y(_06678_),
    .A(net4755),
    .B(_06677_));
 sg13g2_o21ai_1 _24447_ (.B1(net4662),
    .Y(_06679_),
    .A1(_06676_),
    .A2(_06678_));
 sg13g2_nor2_1 _24448_ (.A(_06673_),
    .B(_06679_),
    .Y(_06680_));
 sg13g2_nor2_1 _24449_ (.A(_06669_),
    .B(_06680_),
    .Y(_02134_));
 sg13g2_o21ai_1 _24450_ (.B1(net6014),
    .Y(_06681_),
    .A1(net7337),
    .A2(net4662));
 sg13g2_xnor2_1 _24451_ (.Y(_06682_),
    .A(_00150_),
    .B(_06671_));
 sg13g2_nor2_2 _24452_ (.A(_06623_),
    .B(_06682_),
    .Y(_06683_));
 sg13g2_o21ai_1 _24453_ (.B1(_06677_),
    .Y(_06684_),
    .A1(net5588),
    .A2(_07995_));
 sg13g2_xor2_1 _24454_ (.B(\atari2600.tia.diag[71] ),
    .A(\atari2600.tia.hmp0[3] ),
    .X(_06685_));
 sg13g2_xnor2_1 _24455_ (.Y(_06686_),
    .A(_06684_),
    .B(_06685_));
 sg13g2_a21oi_1 _24456_ (.A1(net4755),
    .A2(_06686_),
    .Y(_06687_),
    .B1(_06683_));
 sg13g2_a21oi_1 _24457_ (.A1(_06621_),
    .A2(_06687_),
    .Y(_02135_),
    .B1(_06681_));
 sg13g2_o21ai_1 _24458_ (.B1(_06619_),
    .Y(_06688_),
    .A1(_05258_),
    .A2(_05394_));
 sg13g2_o21ai_1 _24459_ (.B1(net6028),
    .Y(_06689_),
    .A1(net7247),
    .A2(net4661));
 sg13g2_nand2b_1 _24460_ (.Y(_06690_),
    .B(\atari2600.tia.hmp1[0] ),
    .A_N(\atari2600.tia.diag[56] ));
 sg13g2_xor2_1 _24461_ (.B(\atari2600.tia.diag[56] ),
    .A(net7150),
    .X(_06691_));
 sg13g2_a21oi_1 _24462_ (.A1(net4757),
    .A2(_06691_),
    .Y(_06692_),
    .B1(_06624_));
 sg13g2_a21oi_1 _24463_ (.A1(net4661),
    .A2(_06692_),
    .Y(_02136_),
    .B1(_06689_));
 sg13g2_o21ai_1 _24464_ (.B1(net6029),
    .Y(_06693_),
    .A1(net7289),
    .A2(net4661));
 sg13g2_nor2b_1 _24465_ (.A(\atari2600.tia.hmp1[1] ),
    .B_N(\atari2600.tia.diag[57] ),
    .Y(_06694_));
 sg13g2_xnor2_1 _24466_ (.Y(_06695_),
    .A(\atari2600.tia.hmp1[1] ),
    .B(\atari2600.tia.diag[57] ));
 sg13g2_xor2_1 _24467_ (.B(_06695_),
    .A(_06690_),
    .X(_06696_));
 sg13g2_a21oi_1 _24468_ (.A1(net4756),
    .A2(_06696_),
    .Y(_06697_),
    .B1(_06629_));
 sg13g2_a21oi_1 _24469_ (.A1(net4661),
    .A2(_06697_),
    .Y(_02137_),
    .B1(_06693_));
 sg13g2_o21ai_1 _24470_ (.B1(net6027),
    .Y(_06698_),
    .A1(net7330),
    .A2(net4661));
 sg13g2_xnor2_1 _24471_ (.Y(_06699_),
    .A(\atari2600.tia.hmp1[2] ),
    .B(\atari2600.tia.diag[58] ));
 sg13g2_a21oi_1 _24472_ (.A1(_06690_),
    .A2(_06695_),
    .Y(_06700_),
    .B1(_06694_));
 sg13g2_nor2b_1 _24473_ (.A(_06700_),
    .B_N(_06699_),
    .Y(_06701_));
 sg13g2_xnor2_1 _24474_ (.Y(_06702_),
    .A(_06699_),
    .B(_06700_));
 sg13g2_a21oi_1 _24475_ (.A1(net4756),
    .A2(_06702_),
    .Y(_06703_),
    .B1(_06636_));
 sg13g2_a21oi_1 _24476_ (.A1(net4661),
    .A2(_06703_),
    .Y(_02138_),
    .B1(_06698_));
 sg13g2_o21ai_1 _24477_ (.B1(net6029),
    .Y(_06704_),
    .A1(net5592),
    .A2(net4660));
 sg13g2_xnor2_1 _24478_ (.Y(_06705_),
    .A(net5587),
    .B(net5592));
 sg13g2_a21oi_2 _24479_ (.B1(_06701_),
    .Y(_06706_),
    .A2(\atari2600.tia.diag[58] ),
    .A1(_07975_));
 sg13g2_nor2b_1 _24480_ (.A(_06706_),
    .B_N(_06705_),
    .Y(_06707_));
 sg13g2_xnor2_1 _24481_ (.Y(_06708_),
    .A(_06705_),
    .B(_06706_));
 sg13g2_a21oi_1 _24482_ (.A1(net4756),
    .A2(_06708_),
    .Y(_06709_),
    .B1(_06645_));
 sg13g2_a21oi_1 _24483_ (.A1(net4661),
    .A2(_06709_),
    .Y(_02139_),
    .B1(_06704_));
 sg13g2_o21ai_1 _24484_ (.B1(net6032),
    .Y(_06710_),
    .A1(net5590),
    .A2(_06688_));
 sg13g2_xnor2_1 _24485_ (.Y(_06711_),
    .A(net5587),
    .B(net5590));
 sg13g2_a21oi_1 _24486_ (.A1(_07974_),
    .A2(net5592),
    .Y(_06712_),
    .B1(_06707_));
 sg13g2_nor2b_1 _24487_ (.A(_06712_),
    .B_N(_06711_),
    .Y(_06713_));
 sg13g2_xnor2_1 _24488_ (.Y(_06714_),
    .A(_06711_),
    .B(_06712_));
 sg13g2_a21oi_1 _24489_ (.A1(net4759),
    .A2(_06714_),
    .Y(_06715_),
    .B1(_06654_));
 sg13g2_a21oi_1 _24490_ (.A1(net4660),
    .A2(_06715_),
    .Y(_02140_),
    .B1(_06710_));
 sg13g2_o21ai_1 _24491_ (.B1(net6032),
    .Y(_06716_),
    .A1(net7327),
    .A2(net4660));
 sg13g2_a21oi_1 _24492_ (.A1(_07974_),
    .A2(net5590),
    .Y(_06717_),
    .B1(_06713_));
 sg13g2_nand2_1 _24493_ (.Y(_06718_),
    .A(\atari2600.tia.hmp1[3] ),
    .B(_07993_));
 sg13g2_xnor2_1 _24494_ (.Y(_06719_),
    .A(net5587),
    .B(\atari2600.tia.diag[61] ));
 sg13g2_xnor2_1 _24495_ (.Y(_06720_),
    .A(_06717_),
    .B(_06719_));
 sg13g2_a21oi_1 _24496_ (.A1(net4759),
    .A2(_06720_),
    .Y(_06721_),
    .B1(_06663_));
 sg13g2_a21oi_1 _24497_ (.A1(net4660),
    .A2(_06721_),
    .Y(_02141_),
    .B1(_06716_));
 sg13g2_o21ai_1 _24498_ (.B1(net6032),
    .Y(_06722_),
    .A1(net5589),
    .A2(net4660));
 sg13g2_xnor2_1 _24499_ (.Y(_06723_),
    .A(net5587),
    .B(net5589));
 sg13g2_o21ai_1 _24500_ (.B1(_06717_),
    .Y(_06724_),
    .A1(net5587),
    .A2(_07993_));
 sg13g2_a21oi_1 _24501_ (.A1(_06718_),
    .A2(_06724_),
    .Y(_06725_),
    .B1(_06723_));
 sg13g2_nand3_1 _24502_ (.B(_06723_),
    .C(_06724_),
    .A(_06718_),
    .Y(_06726_));
 sg13g2_nor2b_1 _24503_ (.A(_06725_),
    .B_N(_06726_),
    .Y(_06727_));
 sg13g2_a21oi_1 _24504_ (.A1(net4758),
    .A2(_06727_),
    .Y(_06728_),
    .B1(_06673_));
 sg13g2_a21oi_1 _24505_ (.A1(net4660),
    .A2(_06728_),
    .Y(_02142_),
    .B1(_06722_));
 sg13g2_o21ai_1 _24506_ (.B1(net6032),
    .Y(_06729_),
    .A1(net7346),
    .A2(net4660));
 sg13g2_o21ai_1 _24507_ (.B1(_06726_),
    .Y(_06730_),
    .A1(net5587),
    .A2(_07992_));
 sg13g2_xor2_1 _24508_ (.B(\atari2600.tia.diag[63] ),
    .A(net5587),
    .X(_06731_));
 sg13g2_xnor2_1 _24509_ (.Y(_06732_),
    .A(_06730_),
    .B(_06731_));
 sg13g2_a21oi_1 _24510_ (.A1(net4758),
    .A2(_06732_),
    .Y(_06733_),
    .B1(_06683_));
 sg13g2_a21oi_1 _24511_ (.A1(net4660),
    .A2(_06733_),
    .Y(_02143_),
    .B1(_06729_));
 sg13g2_a21oi_1 _24512_ (.A1(_05260_),
    .A2(_05393_),
    .Y(_06734_),
    .B1(_06618_));
 sg13g2_a221oi_1 _24513_ (.B2(_06471_),
    .C1(_06618_),
    .B1(_06454_),
    .A1(_05260_),
    .Y(_06735_),
    .A2(_05393_));
 sg13g2_o21ai_1 _24514_ (.B1(_06734_),
    .Y(_06736_),
    .A1(_06455_),
    .A2(_06472_));
 sg13g2_nor2_2 _24515_ (.A(net4771),
    .B(_06455_),
    .Y(_06737_));
 sg13g2_nand2_1 _24516_ (.Y(_06738_),
    .A(_08782_),
    .B(_06454_));
 sg13g2_o21ai_1 _24517_ (.B1(net6005),
    .Y(_06739_),
    .A1(net7305),
    .A2(_06736_));
 sg13g2_nand2_1 _24518_ (.Y(_06740_),
    .A(_06624_),
    .B(net4753));
 sg13g2_nor2b_1 _24519_ (.A(\atari2600.tia.diag[48] ),
    .B_N(\atari2600.tia.hmm0[0] ),
    .Y(_06741_));
 sg13g2_xor2_1 _24520_ (.B(\atari2600.tia.diag[48] ),
    .A(net7126),
    .X(_06742_));
 sg13g2_a221oi_1 _24521_ (.B2(net4754),
    .C1(net4658),
    .B1(_06742_),
    .A1(net7285),
    .Y(_06743_),
    .A2(_06737_));
 sg13g2_a21oi_1 _24522_ (.A1(_06740_),
    .A2(_06743_),
    .Y(_02144_),
    .B1(_06739_));
 sg13g2_o21ai_1 _24523_ (.B1(net6006),
    .Y(_06744_),
    .A1(net7329),
    .A2(_06736_));
 sg13g2_nand2_1 _24524_ (.Y(_06745_),
    .A(_06629_),
    .B(net4753));
 sg13g2_xor2_1 _24525_ (.B(\atari2600.tia.diag[49] ),
    .A(\atari2600.tia.hmm0[1] ),
    .X(_06746_));
 sg13g2_nor2_1 _24526_ (.A(_06741_),
    .B(_06746_),
    .Y(_06747_));
 sg13g2_xor2_1 _24527_ (.B(_06746_),
    .A(_06741_),
    .X(_06748_));
 sg13g2_a221oi_1 _24528_ (.B2(net4754),
    .C1(net4658),
    .B1(_06748_),
    .A1(net7296),
    .Y(_06749_),
    .A2(_06737_));
 sg13g2_a21oi_1 _24529_ (.A1(_06745_),
    .A2(_06749_),
    .Y(_02145_),
    .B1(_06744_));
 sg13g2_nand2_1 _24530_ (.Y(_06750_),
    .A(_06636_),
    .B(net4753));
 sg13g2_xor2_1 _24531_ (.B(\atari2600.tia.p0_w[3] ),
    .A(net5596),
    .X(_06751_));
 sg13g2_nand2b_1 _24532_ (.Y(_06752_),
    .B(\atari2600.tia.diag[50] ),
    .A_N(\atari2600.tia.hmm0[2] ));
 sg13g2_xor2_1 _24533_ (.B(\atari2600.tia.diag[50] ),
    .A(\atari2600.tia.hmm0[2] ),
    .X(_06753_));
 sg13g2_a21oi_1 _24534_ (.A1(_07973_),
    .A2(\atari2600.tia.diag[49] ),
    .Y(_06754_),
    .B1(_06747_));
 sg13g2_or2_1 _24535_ (.X(_06755_),
    .B(_06754_),
    .A(_06753_));
 sg13g2_a21oi_1 _24536_ (.A1(_06753_),
    .A2(_06754_),
    .Y(_06756_),
    .B1(_06617_));
 sg13g2_a221oi_1 _24537_ (.B2(_06756_),
    .C1(net4658),
    .B1(_06755_),
    .A1(_06737_),
    .Y(_06757_),
    .A2(_06751_));
 sg13g2_o21ai_1 _24538_ (.B1(net6006),
    .Y(_06758_),
    .A1(net7301),
    .A2(_06736_));
 sg13g2_a21oi_1 _24539_ (.A1(_06750_),
    .A2(_06757_),
    .Y(_02146_),
    .B1(_06758_));
 sg13g2_nand2_1 _24540_ (.Y(_06759_),
    .A(_06645_),
    .B(net4753));
 sg13g2_xor2_1 _24541_ (.B(\atari2600.tia.diag[51] ),
    .A(net5586),
    .X(_06760_));
 sg13g2_nand3_1 _24542_ (.B(_06755_),
    .C(_06760_),
    .A(_06752_),
    .Y(_06761_));
 sg13g2_a21oi_1 _24543_ (.A1(_06752_),
    .A2(_06755_),
    .Y(_06762_),
    .B1(_06760_));
 sg13g2_nor2_1 _24544_ (.A(_06617_),
    .B(_06762_),
    .Y(_06763_));
 sg13g2_nand2_1 _24545_ (.Y(_06764_),
    .A(net5595),
    .B(\atari2600.tia.p0_w[4] ));
 sg13g2_xor2_1 _24546_ (.B(\atari2600.tia.p0_w[4] ),
    .A(net5595),
    .X(_06765_));
 sg13g2_nand3_1 _24547_ (.B(\atari2600.tia.p0_w[3] ),
    .C(_06765_),
    .A(\atari2600.tia.diag[66] ),
    .Y(_06766_));
 sg13g2_a21oi_1 _24548_ (.A1(net5596),
    .A2(\atari2600.tia.p0_w[3] ),
    .Y(_06767_),
    .B1(_06765_));
 sg13g2_nor2_1 _24549_ (.A(net4753),
    .B(_06767_),
    .Y(_06768_));
 sg13g2_a221oi_1 _24550_ (.B2(_06768_),
    .C1(net4658),
    .B1(_06766_),
    .A1(_06761_),
    .Y(_06769_),
    .A2(_06763_));
 sg13g2_o21ai_1 _24551_ (.B1(net6008),
    .Y(_06770_),
    .A1(net7309),
    .A2(_06736_));
 sg13g2_a21oi_1 _24552_ (.A1(_06759_),
    .A2(_06769_),
    .Y(_02147_),
    .B1(_06770_));
 sg13g2_nand2_1 _24553_ (.Y(_06771_),
    .A(_06654_),
    .B(net4753));
 sg13g2_xor2_1 _24554_ (.B(\atari2600.tia.diag[52] ),
    .A(net5586),
    .X(_06772_));
 sg13g2_a21o_1 _24555_ (.A2(\atari2600.tia.diag[51] ),
    .A1(_07972_),
    .B1(_06762_),
    .X(_06773_));
 sg13g2_nand2b_1 _24556_ (.Y(_06774_),
    .B(_06773_),
    .A_N(_06772_));
 sg13g2_xnor2_1 _24557_ (.Y(_06775_),
    .A(_06772_),
    .B(_06773_));
 sg13g2_nand2_1 _24558_ (.Y(_06776_),
    .A(net5594),
    .B(\atari2600.tia.p0_w[5] ));
 sg13g2_xnor2_1 _24559_ (.Y(_06777_),
    .A(net5594),
    .B(\atari2600.tia.p0_w[5] ));
 sg13g2_a21oi_2 _24560_ (.B1(_06777_),
    .Y(_06778_),
    .A2(_06766_),
    .A1(_06764_));
 sg13g2_nand3_1 _24561_ (.B(_06766_),
    .C(_06777_),
    .A(_06764_),
    .Y(_06779_));
 sg13g2_nor2b_1 _24562_ (.A(_06778_),
    .B_N(_06779_),
    .Y(_06780_));
 sg13g2_a221oi_1 _24563_ (.B2(_06737_),
    .C1(net4658),
    .B1(_06780_),
    .A1(net4754),
    .Y(_06781_),
    .A2(_06775_));
 sg13g2_a221oi_1 _24564_ (.B2(_06781_),
    .C1(net5983),
    .B1(_06771_),
    .A1(_07990_),
    .Y(_02148_),
    .A2(net4658));
 sg13g2_nand2_1 _24565_ (.Y(_06782_),
    .A(_06663_),
    .B(_06738_));
 sg13g2_o21ai_1 _24566_ (.B1(_06774_),
    .Y(_06783_),
    .A1(net5586),
    .A2(_07990_));
 sg13g2_xor2_1 _24567_ (.B(\atari2600.tia.diag[53] ),
    .A(net5586),
    .X(_06784_));
 sg13g2_xnor2_1 _24568_ (.Y(_06785_),
    .A(_06783_),
    .B(_06784_));
 sg13g2_a21oi_1 _24569_ (.A1(net5594),
    .A2(\atari2600.tia.p0_w[5] ),
    .Y(_06786_),
    .B1(_06778_));
 sg13g2_xnor2_1 _24570_ (.Y(_06787_),
    .A(net5593),
    .B(_06786_));
 sg13g2_a221oi_1 _24571_ (.B2(_06737_),
    .C1(net4659),
    .B1(_06787_),
    .A1(net4755),
    .Y(_06788_),
    .A2(_06785_));
 sg13g2_a221oi_1 _24572_ (.B2(_06788_),
    .C1(net5983),
    .B1(_06782_),
    .A1(_07989_),
    .Y(_02149_),
    .A2(net4659));
 sg13g2_nand2_1 _24573_ (.Y(_06789_),
    .A(_06673_),
    .B(net4753));
 sg13g2_nor2_1 _24574_ (.A(\atari2600.tia.hmm0[3] ),
    .B(_07988_),
    .Y(_06790_));
 sg13g2_nand2_1 _24575_ (.Y(_06791_),
    .A(net5586),
    .B(_07988_));
 sg13g2_nand2b_1 _24576_ (.Y(_06792_),
    .B(_06791_),
    .A_N(_06790_));
 sg13g2_o21ai_1 _24577_ (.B1(_06783_),
    .Y(_06793_),
    .A1(_07972_),
    .A2(\atari2600.tia.diag[53] ));
 sg13g2_o21ai_1 _24578_ (.B1(_06793_),
    .Y(_06794_),
    .A1(net5586),
    .A2(_07989_));
 sg13g2_xnor2_1 _24579_ (.Y(_06795_),
    .A(_06792_),
    .B(_06794_));
 sg13g2_nand2_1 _24580_ (.Y(_06796_),
    .A(net5593),
    .B(_06778_));
 sg13g2_o21ai_1 _24581_ (.B1(_06796_),
    .Y(_06797_),
    .A1(_00161_),
    .A2(_06776_));
 sg13g2_nand2_1 _24582_ (.Y(_06798_),
    .A(\atari2600.tia.diag[70] ),
    .B(_06797_));
 sg13g2_xnor2_1 _24583_ (.Y(_06799_),
    .A(_07995_),
    .B(_06797_));
 sg13g2_a221oi_1 _24584_ (.B2(_06737_),
    .C1(net4659),
    .B1(_06799_),
    .A1(net4754),
    .Y(_06800_),
    .A2(_06795_));
 sg13g2_a221oi_1 _24585_ (.B2(_06800_),
    .C1(net5983),
    .B1(_06789_),
    .A1(_07988_),
    .Y(_02150_),
    .A2(net4659));
 sg13g2_nand2_1 _24586_ (.Y(_06801_),
    .A(_06683_),
    .B(net4753));
 sg13g2_a21oi_1 _24587_ (.A1(_06791_),
    .A2(_06794_),
    .Y(_06802_),
    .B1(_06790_));
 sg13g2_xnor2_1 _24588_ (.Y(_06803_),
    .A(net5586),
    .B(\atari2600.tia.diag[55] ));
 sg13g2_xnor2_1 _24589_ (.Y(_06804_),
    .A(_06802_),
    .B(_06803_));
 sg13g2_xor2_1 _24590_ (.B(_06798_),
    .A(_00162_),
    .X(_06805_));
 sg13g2_a221oi_1 _24591_ (.B2(_06737_),
    .C1(net4658),
    .B1(_06805_),
    .A1(net4754),
    .Y(_06806_),
    .A2(_06804_));
 sg13g2_a221oi_1 _24592_ (.B2(_06806_),
    .C1(net5983),
    .B1(_06801_),
    .A1(_07987_),
    .Y(_02151_),
    .A2(net4658));
 sg13g2_nor2_2 _24593_ (.A(net4948),
    .B(net4932),
    .Y(_06807_));
 sg13g2_nor2_2 _24594_ (.A(net4771),
    .B(_06421_),
    .Y(_06808_));
 sg13g2_or2_2 _24595_ (.X(_06809_),
    .B(_06421_),
    .A(net4771));
 sg13g2_a221oi_1 _24596_ (.B2(_08753_),
    .C1(_06808_),
    .B1(_06807_),
    .A1(_08782_),
    .Y(_06810_),
    .A2(_05446_));
 sg13g2_nor2_2 _24597_ (.A(_08606_),
    .B(_06810_),
    .Y(_06811_));
 sg13g2_nor3_1 _24598_ (.A(net5829),
    .B(net4726),
    .C(_06808_),
    .Y(_06812_));
 sg13g2_nand2b_1 _24599_ (.Y(_06813_),
    .B(\atari2600.tia.hmm1[0] ),
    .A_N(\atari2600.tia.diag[40] ));
 sg13g2_xor2_1 _24600_ (.B(\atari2600.tia.diag[40] ),
    .A(net7161),
    .X(_06814_));
 sg13g2_a221oi_1 _24601_ (.B2(net4756),
    .C1(_06812_),
    .B1(_06814_),
    .A1(net7247),
    .Y(_06815_),
    .A2(_06808_));
 sg13g2_o21ai_1 _24602_ (.B1(net6028),
    .Y(_06816_),
    .A1(net7278),
    .A2(net4656));
 sg13g2_a21oi_1 _24603_ (.A1(net4656),
    .A2(_06815_),
    .Y(_02152_),
    .B1(_06816_));
 sg13g2_nor2b_1 _24604_ (.A(\atari2600.tia.hmm1[1] ),
    .B_N(\atari2600.tia.diag[41] ),
    .Y(_06817_));
 sg13g2_xnor2_1 _24605_ (.Y(_06818_),
    .A(\atari2600.tia.hmm1[1] ),
    .B(\atari2600.tia.diag[41] ));
 sg13g2_xor2_1 _24606_ (.B(_06818_),
    .A(_06813_),
    .X(_06819_));
 sg13g2_and2_1 _24607_ (.A(\atari2600.tia.diag[57] ),
    .B(_06808_),
    .X(_06820_));
 sg13g2_a221oi_1 _24608_ (.B2(net4756),
    .C1(_06820_),
    .B1(_06819_),
    .A1(_06629_),
    .Y(_06821_),
    .A2(net4752));
 sg13g2_o21ai_1 _24609_ (.B1(net6028),
    .Y(_06822_),
    .A1(net7273),
    .A2(net4656));
 sg13g2_a21oi_1 _24610_ (.A1(net4656),
    .A2(_06821_),
    .Y(_02153_),
    .B1(_06822_));
 sg13g2_nand2b_1 _24611_ (.Y(_06823_),
    .B(\atari2600.tia.diag[42] ),
    .A_N(\atari2600.tia.hmm1[2] ));
 sg13g2_xor2_1 _24612_ (.B(\atari2600.tia.diag[42] ),
    .A(\atari2600.tia.hmm1[2] ),
    .X(_06824_));
 sg13g2_a21oi_1 _24613_ (.A1(_06813_),
    .A2(_06818_),
    .Y(_06825_),
    .B1(_06817_));
 sg13g2_xor2_1 _24614_ (.B(_06825_),
    .A(_06824_),
    .X(_06826_));
 sg13g2_nand2_1 _24615_ (.Y(_06827_),
    .A(\atari2600.tia.diag[58] ),
    .B(\atari2600.tia.p1_w[3] ));
 sg13g2_or2_1 _24616_ (.X(_06828_),
    .B(\atari2600.tia.p1_w[3] ),
    .A(\atari2600.tia.diag[58] ));
 sg13g2_and3_1 _24617_ (.X(_06829_),
    .A(_06808_),
    .B(_06827_),
    .C(_06828_));
 sg13g2_a221oi_1 _24618_ (.B2(net4756),
    .C1(_06829_),
    .B1(_06826_),
    .A1(_06636_),
    .Y(_06830_),
    .A2(net4752));
 sg13g2_o21ai_1 _24619_ (.B1(net6028),
    .Y(_06831_),
    .A1(net7312),
    .A2(net4656));
 sg13g2_a21oi_1 _24620_ (.A1(net4656),
    .A2(_06830_),
    .Y(_02154_),
    .B1(_06831_));
 sg13g2_nand2_1 _24621_ (.Y(_06832_),
    .A(_07971_),
    .B(\atari2600.tia.diag[43] ));
 sg13g2_xor2_1 _24622_ (.B(\atari2600.tia.diag[43] ),
    .A(net5585),
    .X(_06833_));
 sg13g2_o21ai_1 _24623_ (.B1(_06823_),
    .Y(_06834_),
    .A1(_06824_),
    .A2(_06825_));
 sg13g2_nand2b_1 _24624_ (.Y(_06835_),
    .B(_06834_),
    .A_N(_06833_));
 sg13g2_xnor2_1 _24625_ (.Y(_06836_),
    .A(_06833_),
    .B(_06834_));
 sg13g2_nand2_1 _24626_ (.Y(_06837_),
    .A(net5592),
    .B(\atari2600.tia.p1_w[4] ));
 sg13g2_xor2_1 _24627_ (.B(\atari2600.tia.p1_w[4] ),
    .A(net5592),
    .X(_06838_));
 sg13g2_nand2b_1 _24628_ (.Y(_06839_),
    .B(_06838_),
    .A_N(_06827_));
 sg13g2_xor2_1 _24629_ (.B(_06838_),
    .A(_06827_),
    .X(_06840_));
 sg13g2_nor2_1 _24630_ (.A(net4752),
    .B(_06840_),
    .Y(_06841_));
 sg13g2_a221oi_1 _24631_ (.B2(net4756),
    .C1(_06841_),
    .B1(_06836_),
    .A1(_06645_),
    .Y(_06842_),
    .A2(net4752));
 sg13g2_o21ai_1 _24632_ (.B1(net6028),
    .Y(_06843_),
    .A1(net7284),
    .A2(net4656));
 sg13g2_a21oi_1 _24633_ (.A1(net4656),
    .A2(_06842_),
    .Y(_02155_),
    .B1(_06843_));
 sg13g2_nand2_1 _24634_ (.Y(_06844_),
    .A(net5591),
    .B(\atari2600.tia.p1_w[5] ));
 sg13g2_xnor2_1 _24635_ (.Y(_06845_),
    .A(net5590),
    .B(\atari2600.tia.p1_w[5] ));
 sg13g2_a21oi_1 _24636_ (.A1(_06837_),
    .A2(_06839_),
    .Y(_06846_),
    .B1(_06845_));
 sg13g2_and3_1 _24637_ (.X(_06847_),
    .A(_06837_),
    .B(_06839_),
    .C(_06845_));
 sg13g2_nor3_1 _24638_ (.A(_06809_),
    .B(_06846_),
    .C(_06847_),
    .Y(_06848_));
 sg13g2_xor2_1 _24639_ (.B(\atari2600.tia.diag[44] ),
    .A(net5585),
    .X(_06849_));
 sg13g2_a21oi_1 _24640_ (.A1(_06832_),
    .A2(_06835_),
    .Y(_06850_),
    .B1(_06849_));
 sg13g2_nand3_1 _24641_ (.B(_06835_),
    .C(_06849_),
    .A(_06832_),
    .Y(_06851_));
 sg13g2_nor2b_1 _24642_ (.A(_06850_),
    .B_N(_06851_),
    .Y(_06852_));
 sg13g2_a221oi_1 _24643_ (.B2(net4757),
    .C1(_06848_),
    .B1(_06852_),
    .A1(_06654_),
    .Y(_06853_),
    .A2(net4752));
 sg13g2_o21ai_1 _24644_ (.B1(net6029),
    .Y(_06854_),
    .A1(net7254),
    .A2(net4657));
 sg13g2_a21oi_1 _24645_ (.A1(net4657),
    .A2(_06853_),
    .Y(_02156_),
    .B1(_06854_));
 sg13g2_a21oi_1 _24646_ (.A1(_07971_),
    .A2(\atari2600.tia.diag[44] ),
    .Y(_06855_),
    .B1(_06850_));
 sg13g2_xnor2_1 _24647_ (.Y(_06856_),
    .A(net5585),
    .B(\atari2600.tia.diag[45] ));
 sg13g2_xnor2_1 _24648_ (.Y(_06857_),
    .A(_06855_),
    .B(_06856_));
 sg13g2_a21oi_1 _24649_ (.A1(net5590),
    .A2(\atari2600.tia.p1_w[5] ),
    .Y(_06858_),
    .B1(_06846_));
 sg13g2_xnor2_1 _24650_ (.Y(_06859_),
    .A(_07993_),
    .B(_06858_));
 sg13g2_nor2_1 _24651_ (.A(_06809_),
    .B(_06859_),
    .Y(_06860_));
 sg13g2_a221oi_1 _24652_ (.B2(net4759),
    .C1(_06860_),
    .B1(_06857_),
    .A1(_06663_),
    .Y(_06861_),
    .A2(net4752));
 sg13g2_o21ai_1 _24653_ (.B1(net6031),
    .Y(_06862_),
    .A1(net7318),
    .A2(net4657));
 sg13g2_a21oi_1 _24654_ (.A1(net4657),
    .A2(_06861_),
    .Y(_02157_),
    .B1(_06862_));
 sg13g2_nor2_1 _24655_ (.A(net5585),
    .B(_07984_),
    .Y(_06863_));
 sg13g2_nand2_1 _24656_ (.Y(_06864_),
    .A(net5585),
    .B(_07984_));
 sg13g2_nand2b_1 _24657_ (.Y(_06865_),
    .B(_06864_),
    .A_N(_06863_));
 sg13g2_a21oi_1 _24658_ (.A1(net5585),
    .A2(_07985_),
    .Y(_06866_),
    .B1(_06855_));
 sg13g2_a21o_1 _24659_ (.A2(\atari2600.tia.diag[45] ),
    .A1(_07971_),
    .B1(_06866_),
    .X(_06867_));
 sg13g2_xnor2_1 _24660_ (.Y(_06868_),
    .A(_06865_),
    .B(_06867_));
 sg13g2_nand2_1 _24661_ (.Y(_06869_),
    .A(\atari2600.tia.diag[61] ),
    .B(_06846_));
 sg13g2_o21ai_1 _24662_ (.B1(_06869_),
    .Y(_06870_),
    .A1(_00157_),
    .A2(_06844_));
 sg13g2_nand2b_1 _24663_ (.Y(_06871_),
    .B(_07992_),
    .A_N(_06870_));
 sg13g2_nand2_1 _24664_ (.Y(_06872_),
    .A(net5589),
    .B(_06870_));
 sg13g2_and3_1 _24665_ (.X(_06873_),
    .A(_06808_),
    .B(_06871_),
    .C(_06872_));
 sg13g2_a221oi_1 _24666_ (.B2(net4758),
    .C1(_06873_),
    .B1(_06868_),
    .A1(_06673_),
    .Y(_06874_),
    .A2(_06809_));
 sg13g2_o21ai_1 _24667_ (.B1(net6029),
    .Y(_06875_),
    .A1(net7235),
    .A2(net4657));
 sg13g2_a21oi_1 _24668_ (.A1(net4657),
    .A2(_06874_),
    .Y(_02158_),
    .B1(_06875_));
 sg13g2_a21oi_1 _24669_ (.A1(_06864_),
    .A2(_06867_),
    .Y(_06876_),
    .B1(_06863_));
 sg13g2_xnor2_1 _24670_ (.Y(_06877_),
    .A(net5585),
    .B(\atari2600.tia.diag[47] ));
 sg13g2_xnor2_1 _24671_ (.Y(_06878_),
    .A(_06876_),
    .B(_06877_));
 sg13g2_xnor2_1 _24672_ (.Y(_06879_),
    .A(_00158_),
    .B(_06872_));
 sg13g2_nor2_1 _24673_ (.A(net4752),
    .B(_06879_),
    .Y(_06880_));
 sg13g2_a221oi_1 _24674_ (.B2(net4758),
    .C1(_06880_),
    .B1(_06878_),
    .A1(_06683_),
    .Y(_06881_),
    .A2(net4752));
 sg13g2_o21ai_1 _24675_ (.B1(net6029),
    .Y(_06882_),
    .A1(net7287),
    .A2(net4657));
 sg13g2_a21oi_1 _24676_ (.A1(net4657),
    .A2(_06881_),
    .Y(_02159_),
    .B1(_06882_));
 sg13g2_o21ai_1 _24677_ (.B1(_06619_),
    .Y(_06883_),
    .A1(_08679_),
    .A2(_05394_));
 sg13g2_o21ai_1 _24678_ (.B1(net6030),
    .Y(_06884_),
    .A1(net7303),
    .A2(net4655));
 sg13g2_nand2b_1 _24679_ (.Y(_06885_),
    .B(\atari2600.tia.hmbl[0] ),
    .A_N(\atari2600.tia.diag[32] ));
 sg13g2_xor2_1 _24680_ (.B(\atari2600.tia.diag[32] ),
    .A(net7201),
    .X(_06886_));
 sg13g2_a21oi_1 _24681_ (.A1(net4757),
    .A2(_06886_),
    .Y(_06887_),
    .B1(_06624_));
 sg13g2_a21oi_1 _24682_ (.A1(net4655),
    .A2(_06887_),
    .Y(_02160_),
    .B1(_06884_));
 sg13g2_o21ai_1 _24683_ (.B1(net6030),
    .Y(_06888_),
    .A1(net7298),
    .A2(net4655));
 sg13g2_nor2b_1 _24684_ (.A(\atari2600.tia.hmbl[1] ),
    .B_N(\atari2600.tia.diag[33] ),
    .Y(_06889_));
 sg13g2_xnor2_1 _24685_ (.Y(_06890_),
    .A(\atari2600.tia.hmbl[1] ),
    .B(\atari2600.tia.diag[33] ));
 sg13g2_xor2_1 _24686_ (.B(_06890_),
    .A(_06885_),
    .X(_06891_));
 sg13g2_a21oi_1 _24687_ (.A1(net4756),
    .A2(_06891_),
    .Y(_06892_),
    .B1(_06629_));
 sg13g2_a21oi_1 _24688_ (.A1(net4655),
    .A2(_06892_),
    .Y(_02161_),
    .B1(_06888_));
 sg13g2_o21ai_1 _24689_ (.B1(net6030),
    .Y(_06893_),
    .A1(net7316),
    .A2(net4655));
 sg13g2_xnor2_1 _24690_ (.Y(_06894_),
    .A(\atari2600.tia.hmbl[2] ),
    .B(\atari2600.tia.diag[34] ));
 sg13g2_a21oi_1 _24691_ (.A1(_06885_),
    .A2(_06890_),
    .Y(_06895_),
    .B1(_06889_));
 sg13g2_nor2b_1 _24692_ (.A(_06895_),
    .B_N(_06894_),
    .Y(_06896_));
 sg13g2_xnor2_1 _24693_ (.Y(_06897_),
    .A(_06894_),
    .B(_06895_));
 sg13g2_a21oi_1 _24694_ (.A1(net4757),
    .A2(_06897_),
    .Y(_06898_),
    .B1(_06636_));
 sg13g2_a21oi_1 _24695_ (.A1(net4655),
    .A2(_06898_),
    .Y(_02162_),
    .B1(_06893_));
 sg13g2_o21ai_1 _24696_ (.B1(net6031),
    .Y(_06899_),
    .A1(net7317),
    .A2(net4654));
 sg13g2_xnor2_1 _24697_ (.Y(_06900_),
    .A(net5584),
    .B(\atari2600.tia.diag[35] ));
 sg13g2_a21oi_2 _24698_ (.B1(_06896_),
    .Y(_06901_),
    .A2(\atari2600.tia.diag[34] ),
    .A1(_07970_));
 sg13g2_nor2b_1 _24699_ (.A(_06901_),
    .B_N(_06900_),
    .Y(_06902_));
 sg13g2_xnor2_1 _24700_ (.Y(_06903_),
    .A(_06900_),
    .B(_06901_));
 sg13g2_a21oi_1 _24701_ (.A1(net4757),
    .A2(_06903_),
    .Y(_06904_),
    .B1(_06645_));
 sg13g2_a21oi_1 _24702_ (.A1(net4655),
    .A2(_06904_),
    .Y(_02163_),
    .B1(_06899_));
 sg13g2_o21ai_1 _24703_ (.B1(net6030),
    .Y(_06905_),
    .A1(net7222),
    .A2(net4654));
 sg13g2_xnor2_1 _24704_ (.Y(_06906_),
    .A(net5584),
    .B(\atari2600.tia.diag[36] ));
 sg13g2_a21oi_1 _24705_ (.A1(_07969_),
    .A2(\atari2600.tia.diag[35] ),
    .Y(_06907_),
    .B1(_06902_));
 sg13g2_nor2b_1 _24706_ (.A(_06907_),
    .B_N(_06906_),
    .Y(_06908_));
 sg13g2_xnor2_1 _24707_ (.Y(_06909_),
    .A(_06906_),
    .B(_06907_));
 sg13g2_a21oi_1 _24708_ (.A1(net4758),
    .A2(_06909_),
    .Y(_06910_),
    .B1(_06654_));
 sg13g2_a21oi_1 _24709_ (.A1(net4654),
    .A2(_06910_),
    .Y(_02164_),
    .B1(_06905_));
 sg13g2_o21ai_1 _24710_ (.B1(net6030),
    .Y(_06911_),
    .A1(net7304),
    .A2(net4654));
 sg13g2_a21oi_1 _24711_ (.A1(_07969_),
    .A2(\atari2600.tia.diag[36] ),
    .Y(_06912_),
    .B1(_06908_));
 sg13g2_nand2_1 _24712_ (.Y(_06913_),
    .A(net5584),
    .B(_07979_));
 sg13g2_xnor2_1 _24713_ (.Y(_06914_),
    .A(net5584),
    .B(\atari2600.tia.diag[37] ));
 sg13g2_xnor2_1 _24714_ (.Y(_06915_),
    .A(_06912_),
    .B(_06914_));
 sg13g2_a21oi_1 _24715_ (.A1(net4758),
    .A2(_06915_),
    .Y(_06916_),
    .B1(_06663_));
 sg13g2_a21oi_1 _24716_ (.A1(_06883_),
    .A2(_06916_),
    .Y(_02165_),
    .B1(_06911_));
 sg13g2_o21ai_1 _24717_ (.B1(net6033),
    .Y(_06917_),
    .A1(net7251),
    .A2(net4654));
 sg13g2_xnor2_1 _24718_ (.Y(_06918_),
    .A(net5584),
    .B(\atari2600.tia.diag[38] ));
 sg13g2_o21ai_1 _24719_ (.B1(_06912_),
    .Y(_06919_),
    .A1(net5584),
    .A2(_07979_));
 sg13g2_a21oi_1 _24720_ (.A1(_06913_),
    .A2(_06919_),
    .Y(_06920_),
    .B1(_06918_));
 sg13g2_nand3_1 _24721_ (.B(_06918_),
    .C(_06919_),
    .A(_06913_),
    .Y(_06921_));
 sg13g2_nor2b_1 _24722_ (.A(_06920_),
    .B_N(_06921_),
    .Y(_06922_));
 sg13g2_a21oi_1 _24723_ (.A1(net4758),
    .A2(_06922_),
    .Y(_06923_),
    .B1(_06673_));
 sg13g2_a21oi_1 _24724_ (.A1(net4654),
    .A2(_06923_),
    .Y(_02166_),
    .B1(_06917_));
 sg13g2_o21ai_1 _24725_ (.B1(net6033),
    .Y(_06924_),
    .A1(net7249),
    .A2(net4654));
 sg13g2_o21ai_1 _24726_ (.B1(_06921_),
    .Y(_06925_),
    .A1(net5584),
    .A2(_07978_));
 sg13g2_xor2_1 _24727_ (.B(\atari2600.tia.diag[39] ),
    .A(\atari2600.tia.hmbl[3] ),
    .X(_06926_));
 sg13g2_xnor2_1 _24728_ (.Y(_06927_),
    .A(_06925_),
    .B(_06926_));
 sg13g2_a21oi_1 _24729_ (.A1(net4758),
    .A2(_06927_),
    .Y(_06928_),
    .B1(_06683_));
 sg13g2_a21oi_1 _24730_ (.A1(net4654),
    .A2(_06928_),
    .Y(_02167_),
    .B1(_06924_));
 sg13g2_nor3_1 _24731_ (.A(net4751),
    .B(net4954),
    .C(net4948),
    .Y(_06929_));
 sg13g2_o21ai_1 _24732_ (.B1(net6012),
    .Y(_06930_),
    .A1(net7046),
    .A2(net4652));
 sg13g2_a21oi_1 _24733_ (.A1(net5264),
    .A2(net4652),
    .Y(_02168_),
    .B1(_06930_));
 sg13g2_o21ai_1 _24734_ (.B1(net6009),
    .Y(_06931_),
    .A1(net6822),
    .A2(net4652));
 sg13g2_a21oi_1 _24735_ (.A1(net5238),
    .A2(net4653),
    .Y(_02169_),
    .B1(_06931_));
 sg13g2_o21ai_1 _24736_ (.B1(net6009),
    .Y(_06932_),
    .A1(net7030),
    .A2(net4653));
 sg13g2_a21oi_1 _24737_ (.A1(net5136),
    .A2(net4653),
    .Y(_02170_),
    .B1(_06932_));
 sg13g2_o21ai_1 _24738_ (.B1(net6009),
    .Y(_06933_),
    .A1(net7025),
    .A2(net4653));
 sg13g2_a21oi_1 _24739_ (.A1(net5107),
    .A2(net4653),
    .Y(_02171_),
    .B1(_06933_));
 sg13g2_o21ai_1 _24740_ (.B1(net6012),
    .Y(_06934_),
    .A1(net7048),
    .A2(net4653));
 sg13g2_a21oi_1 _24741_ (.A1(net5179),
    .A2(net4653),
    .Y(_02172_),
    .B1(_06934_));
 sg13g2_o21ai_1 _24742_ (.B1(net6012),
    .Y(_06935_),
    .A1(net6957),
    .A2(_06929_));
 sg13g2_a21oi_1 _24743_ (.A1(net5151),
    .A2(net4652),
    .Y(_02173_),
    .B1(_06935_));
 sg13g2_nand2_1 _24744_ (.Y(_06936_),
    .A(net5086),
    .B(net4652));
 sg13g2_o21ai_1 _24745_ (.B1(_06936_),
    .Y(_06937_),
    .A1(net7015),
    .A2(net4652));
 sg13g2_nor2_1 _24746_ (.A(net5983),
    .B(_06937_),
    .Y(_02174_));
 sg13g2_nand2_1 _24747_ (.Y(_06938_),
    .A(net5059),
    .B(net4652));
 sg13g2_o21ai_1 _24748_ (.B1(_06938_),
    .Y(_06939_),
    .A1(net7047),
    .A2(net4652));
 sg13g2_nor2_1 _24749_ (.A(net5983),
    .B(_06939_),
    .Y(_02175_));
 sg13g2_a21oi_2 _24750_ (.B1(_06472_),
    .Y(_06940_),
    .A2(_06615_),
    .A1(_05392_));
 sg13g2_nand2_2 _24751_ (.Y(_06941_),
    .A(_08782_),
    .B(_05391_));
 sg13g2_nand2_2 _24752_ (.Y(_06942_),
    .A(net5193),
    .B(_06941_));
 sg13g2_o21ai_1 _24753_ (.B1(net6006),
    .Y(_06943_),
    .A1(net7162),
    .A2(_06940_));
 sg13g2_a21oi_1 _24754_ (.A1(_06940_),
    .A2(_06942_),
    .Y(_02176_),
    .B1(_06943_));
 sg13g2_nand2_2 _24755_ (.Y(_06944_),
    .A(net5169),
    .B(_06941_));
 sg13g2_o21ai_1 _24756_ (.B1(net6006),
    .Y(_06945_),
    .A1(net7191),
    .A2(_06940_));
 sg13g2_a21oi_1 _24757_ (.A1(_06940_),
    .A2(_06944_),
    .Y(_02177_),
    .B1(_06945_));
 sg13g2_nand2_2 _24758_ (.Y(_06946_),
    .A(net5072),
    .B(_06941_));
 sg13g2_o21ai_1 _24759_ (.B1(net6003),
    .Y(_06947_),
    .A1(net7160),
    .A2(_06940_));
 sg13g2_a21oi_1 _24760_ (.A1(_06940_),
    .A2(_06946_),
    .Y(_02178_),
    .B1(_06947_));
 sg13g2_nand2_2 _24761_ (.Y(_06948_),
    .A(net5051),
    .B(_06941_));
 sg13g2_o21ai_1 _24762_ (.B1(net6005),
    .Y(_06949_),
    .A1(net5588),
    .A2(_06940_));
 sg13g2_a21oi_1 _24763_ (.A1(_06940_),
    .A2(_06948_),
    .Y(_02179_),
    .B1(_06949_));
 sg13g2_a21oi_2 _24764_ (.B1(_06472_),
    .Y(_06950_),
    .A2(_05392_),
    .A1(_05258_));
 sg13g2_o21ai_1 _24765_ (.B1(net6027),
    .Y(_06951_),
    .A1(net7150),
    .A2(_06950_));
 sg13g2_a21oi_1 _24766_ (.A1(_06942_),
    .A2(_06950_),
    .Y(_02180_),
    .B1(_06951_));
 sg13g2_o21ai_1 _24767_ (.B1(net6027),
    .Y(_06952_),
    .A1(net7144),
    .A2(_06950_));
 sg13g2_a21oi_1 _24768_ (.A1(_06944_),
    .A2(_06950_),
    .Y(_02181_),
    .B1(_06952_));
 sg13g2_o21ai_1 _24769_ (.B1(net6027),
    .Y(_06953_),
    .A1(net7125),
    .A2(_06950_));
 sg13g2_a21oi_1 _24770_ (.A1(_06946_),
    .A2(_06950_),
    .Y(_02182_),
    .B1(_06953_));
 sg13g2_o21ai_1 _24771_ (.B1(net6008),
    .Y(_06954_),
    .A1(net7212),
    .A2(_06950_));
 sg13g2_a21oi_1 _24772_ (.A1(_06948_),
    .A2(_06950_),
    .Y(_02183_),
    .B1(_06954_));
 sg13g2_a21oi_2 _24773_ (.B1(_06472_),
    .Y(_06955_),
    .A2(_05392_),
    .A1(_05261_));
 sg13g2_o21ai_1 _24774_ (.B1(net6003),
    .Y(_06956_),
    .A1(net7126),
    .A2(_06955_));
 sg13g2_a21oi_1 _24775_ (.A1(_06942_),
    .A2(_06955_),
    .Y(_02184_),
    .B1(_06956_));
 sg13g2_o21ai_1 _24776_ (.B1(net6003),
    .Y(_06957_),
    .A1(net7134),
    .A2(_06955_));
 sg13g2_a21oi_1 _24777_ (.A1(_06944_),
    .A2(_06955_),
    .Y(_02185_),
    .B1(_06957_));
 sg13g2_o21ai_1 _24778_ (.B1(net6005),
    .Y(_06958_),
    .A1(net7114),
    .A2(_06955_));
 sg13g2_a21oi_1 _24779_ (.A1(_06946_),
    .A2(_06955_),
    .Y(_02186_),
    .B1(_06958_));
 sg13g2_nand2_1 _24780_ (.Y(_06959_),
    .A(_06948_),
    .B(_06955_));
 sg13g2_o21ai_1 _24781_ (.B1(_06959_),
    .Y(_06960_),
    .A1(net7118),
    .A2(_06955_));
 sg13g2_nor2_1 _24782_ (.A(net5984),
    .B(_06960_),
    .Y(_02187_));
 sg13g2_and2_2 _24783_ (.A(_03043_),
    .B(_06471_),
    .X(_06961_));
 sg13g2_o21ai_1 _24784_ (.B1(net6007),
    .Y(_06962_),
    .A1(net7161),
    .A2(_06961_));
 sg13g2_a21oi_1 _24785_ (.A1(_06942_),
    .A2(_06961_),
    .Y(_02188_),
    .B1(_06962_));
 sg13g2_o21ai_1 _24786_ (.B1(net6027),
    .Y(_06963_),
    .A1(net7182),
    .A2(_06961_));
 sg13g2_a21oi_1 _24787_ (.A1(_06944_),
    .A2(_06961_),
    .Y(_02189_),
    .B1(_06963_));
 sg13g2_o21ai_1 _24788_ (.B1(net6028),
    .Y(_06964_),
    .A1(net7165),
    .A2(_06961_));
 sg13g2_a21oi_1 _24789_ (.A1(_06946_),
    .A2(_06961_),
    .Y(_02190_),
    .B1(_06964_));
 sg13g2_o21ai_1 _24790_ (.B1(net6007),
    .Y(_06965_),
    .A1(net5585),
    .A2(_06961_));
 sg13g2_a21oi_1 _24791_ (.A1(_06948_),
    .A2(_06961_),
    .Y(_02191_),
    .B1(_06965_));
 sg13g2_a21oi_2 _24792_ (.B1(_06472_),
    .Y(_06966_),
    .A2(_05392_),
    .A1(_08679_));
 sg13g2_o21ai_1 _24793_ (.B1(net6027),
    .Y(_06967_),
    .A1(net7201),
    .A2(_06966_));
 sg13g2_a21oi_1 _24794_ (.A1(_06942_),
    .A2(_06966_),
    .Y(_02192_),
    .B1(_06967_));
 sg13g2_o21ai_1 _24795_ (.B1(net6027),
    .Y(_06968_),
    .A1(net7219),
    .A2(_06966_));
 sg13g2_a21oi_1 _24796_ (.A1(_06944_),
    .A2(_06966_),
    .Y(_02193_),
    .B1(_06968_));
 sg13g2_o21ai_1 _24797_ (.B1(net6027),
    .Y(_06969_),
    .A1(net7252),
    .A2(_06966_));
 sg13g2_a21oi_1 _24798_ (.A1(_06946_),
    .A2(_06966_),
    .Y(_02194_),
    .B1(_06969_));
 sg13g2_o21ai_1 _24799_ (.B1(net6006),
    .Y(_06970_),
    .A1(net7302),
    .A2(_06966_));
 sg13g2_a21oi_1 _24800_ (.A1(_06948_),
    .A2(_06966_),
    .Y(_02195_),
    .B1(_06970_));
 sg13g2_nand2_1 _24801_ (.Y(_06971_),
    .A(net2963),
    .B(net5280));
 sg13g2_nor2_1 _24802_ (.A(net5982),
    .B(net5037),
    .Y(_02856_));
 sg13g2_nand3_1 _24803_ (.B(_06471_),
    .C(_06479_),
    .A(net6018),
    .Y(_06972_));
 sg13g2_nand2_1 _24804_ (.Y(_02196_),
    .A(_06971_),
    .B(_06972_));
 sg13g2_nor2_2 _24805_ (.A(_08584_),
    .B(_05397_),
    .Y(_06973_));
 sg13g2_inv_1 _24806_ (.Y(_06974_),
    .A(_06973_));
 sg13g2_o21ai_1 _24807_ (.B1(net6024),
    .Y(_06975_),
    .A1(net7277),
    .A2(_06973_));
 sg13g2_a21oi_1 _24808_ (.A1(net5268),
    .A2(_06973_),
    .Y(_02197_),
    .B1(_06975_));
 sg13g2_o21ai_1 _24809_ (.B1(net6024),
    .Y(_06976_),
    .A1(net5232),
    .A2(_06974_));
 sg13g2_a21oi_1 _24810_ (.A1(_07967_),
    .A2(_06974_),
    .Y(_02198_),
    .B1(_06976_));
 sg13g2_o21ai_1 _24811_ (.B1(net6024),
    .Y(_06977_),
    .A1(net7293),
    .A2(_06973_));
 sg13g2_a21oi_1 _24812_ (.A1(net5139),
    .A2(_06973_),
    .Y(_02199_),
    .B1(_06977_));
 sg13g2_o21ai_1 _24813_ (.B1(net6024),
    .Y(_06978_),
    .A1(net7283),
    .A2(_06973_));
 sg13g2_a21oi_1 _24814_ (.A1(net5111),
    .A2(_06973_),
    .Y(_02200_),
    .B1(_06978_));
 sg13g2_nand2_2 _24815_ (.Y(_06979_),
    .A(_05396_),
    .B(_06430_));
 sg13g2_o21ai_1 _24816_ (.B1(net6035),
    .Y(_06980_),
    .A1(net5258),
    .A2(_06979_));
 sg13g2_a21oi_1 _24817_ (.A1(_07966_),
    .A2(_06979_),
    .Y(_02201_),
    .B1(_06980_));
 sg13g2_o21ai_1 _24818_ (.B1(net6035),
    .Y(_06981_),
    .A1(net5232),
    .A2(_06979_));
 sg13g2_a21oi_1 _24819_ (.A1(_07965_),
    .A2(_06979_),
    .Y(_02202_),
    .B1(_06981_));
 sg13g2_o21ai_1 _24820_ (.B1(net6035),
    .Y(_06982_),
    .A1(net5129),
    .A2(_06979_));
 sg13g2_a21oi_1 _24821_ (.A1(_07964_),
    .A2(_06979_),
    .Y(_02203_),
    .B1(_06982_));
 sg13g2_o21ai_1 _24822_ (.B1(net6035),
    .Y(_06983_),
    .A1(net5101),
    .A2(_06979_));
 sg13g2_a21oi_1 _24823_ (.A1(_07963_),
    .A2(_06979_),
    .Y(_02204_),
    .B1(_06983_));
 sg13g2_or2_2 _24824_ (.X(_06984_),
    .B(_06421_),
    .A(_05397_));
 sg13g2_o21ai_1 _24825_ (.B1(net6022),
    .Y(_06985_),
    .A1(net5259),
    .A2(_06984_));
 sg13g2_a21oi_1 _24826_ (.A1(_07962_),
    .A2(_06984_),
    .Y(_02205_),
    .B1(_06985_));
 sg13g2_o21ai_1 _24827_ (.B1(net6022),
    .Y(_06986_),
    .A1(net5233),
    .A2(_06984_));
 sg13g2_a21oi_1 _24828_ (.A1(_07961_),
    .A2(_06984_),
    .Y(_02206_),
    .B1(_06986_));
 sg13g2_o21ai_1 _24829_ (.B1(net6022),
    .Y(_06987_),
    .A1(net5130),
    .A2(_06984_));
 sg13g2_a21oi_1 _24830_ (.A1(_07960_),
    .A2(_06984_),
    .Y(_02207_),
    .B1(_06987_));
 sg13g2_o21ai_1 _24831_ (.B1(net6022),
    .Y(_06988_),
    .A1(net5102),
    .A2(_06984_));
 sg13g2_a21oi_1 _24832_ (.A1(_07959_),
    .A2(_06984_),
    .Y(_02208_),
    .B1(_06988_));
 sg13g2_nand2_2 _24833_ (.Y(_06989_),
    .A(_05396_),
    .B(_05446_));
 sg13g2_o21ai_1 _24834_ (.B1(net6017),
    .Y(_06990_),
    .A1(net5258),
    .A2(_06989_));
 sg13g2_a21oi_1 _24835_ (.A1(_07958_),
    .A2(_06989_),
    .Y(_02209_),
    .B1(_06990_));
 sg13g2_o21ai_1 _24836_ (.B1(net6023),
    .Y(_06991_),
    .A1(net5232),
    .A2(_06989_));
 sg13g2_a21oi_1 _24837_ (.A1(_07957_),
    .A2(_06989_),
    .Y(_02210_),
    .B1(_06991_));
 sg13g2_o21ai_1 _24838_ (.B1(net6023),
    .Y(_06992_),
    .A1(net5128),
    .A2(_06989_));
 sg13g2_a21oi_1 _24839_ (.A1(_07956_),
    .A2(_06989_),
    .Y(_02211_),
    .B1(_06992_));
 sg13g2_o21ai_1 _24840_ (.B1(net6023),
    .Y(_06993_),
    .A1(net5100),
    .A2(_06989_));
 sg13g2_a21oi_1 _24841_ (.A1(_07955_),
    .A2(_06989_),
    .Y(_02212_),
    .B1(_06993_));
 sg13g2_nand2_2 _24842_ (.Y(_06994_),
    .A(_05396_),
    .B(_06442_));
 sg13g2_o21ai_1 _24843_ (.B1(net6024),
    .Y(_06995_),
    .A1(net5258),
    .A2(net4725));
 sg13g2_a21oi_1 _24844_ (.A1(_07954_),
    .A2(net4725),
    .Y(_02213_),
    .B1(_06995_));
 sg13g2_o21ai_1 _24845_ (.B1(net6024),
    .Y(_06996_),
    .A1(net5232),
    .A2(net4725));
 sg13g2_a21oi_1 _24846_ (.A1(_07953_),
    .A2(net4725),
    .Y(_02214_),
    .B1(_06996_));
 sg13g2_o21ai_1 _24847_ (.B1(net6024),
    .Y(_06997_),
    .A1(net5129),
    .A2(net4725));
 sg13g2_a21oi_1 _24848_ (.A1(_07952_),
    .A2(net4725),
    .Y(_02215_),
    .B1(_06997_));
 sg13g2_o21ai_1 _24849_ (.B1(net6024),
    .Y(_06998_),
    .A1(net5101),
    .A2(_06994_));
 sg13g2_a21oi_1 _24850_ (.A1(_07951_),
    .A2(net4725),
    .Y(_02216_),
    .B1(_06998_));
 sg13g2_o21ai_1 _24851_ (.B1(net6025),
    .Y(_06999_),
    .A1(net5196),
    .A2(_06994_));
 sg13g2_a21oi_1 _24852_ (.A1(_07950_),
    .A2(net4725),
    .Y(_02217_),
    .B1(_06999_));
 sg13g2_nor2_2 _24853_ (.A(_05397_),
    .B(_06455_),
    .Y(_07000_));
 sg13g2_nand2_2 _24854_ (.Y(_07001_),
    .A(_05396_),
    .B(_06454_));
 sg13g2_o21ai_1 _24855_ (.B1(net6034),
    .Y(_07002_),
    .A1(net5258),
    .A2(_07001_));
 sg13g2_a21oi_1 _24856_ (.A1(_07949_),
    .A2(_07001_),
    .Y(_02218_),
    .B1(_07002_));
 sg13g2_o21ai_1 _24857_ (.B1(net6034),
    .Y(_07003_),
    .A1(net5232),
    .A2(_07001_));
 sg13g2_a21oi_1 _24858_ (.A1(_07948_),
    .A2(_07001_),
    .Y(_02219_),
    .B1(_07003_));
 sg13g2_o21ai_1 _24859_ (.B1(net6034),
    .Y(_07004_),
    .A1(net5129),
    .A2(_07001_));
 sg13g2_a21oi_1 _24860_ (.A1(_07947_),
    .A2(_07001_),
    .Y(_02220_),
    .B1(_07004_));
 sg13g2_o21ai_1 _24861_ (.B1(net6034),
    .Y(_07005_),
    .A1(net5101),
    .A2(_07001_));
 sg13g2_a21oi_1 _24862_ (.A1(_07946_),
    .A2(_07001_),
    .Y(_02221_),
    .B1(_07005_));
 sg13g2_o21ai_1 _24863_ (.B1(net6034),
    .Y(_07006_),
    .A1(net7041),
    .A2(_07000_));
 sg13g2_a21oi_1 _24864_ (.A1(net5184),
    .A2(_07000_),
    .Y(_02222_),
    .B1(_07006_));
 sg13g2_a21oi_1 _24865_ (.A1(\atari2600.tia.audio_left_counter[1] ),
    .A2(_05862_),
    .Y(_07007_),
    .B1(_08099_));
 sg13g2_nand4_1 _24866_ (.B(_05861_),
    .C(_05867_),
    .A(_05860_),
    .Y(_07008_),
    .D(_07007_));
 sg13g2_nor2_1 _24867_ (.A(_05858_),
    .B(_07008_),
    .Y(_07009_));
 sg13g2_nand3_1 _24868_ (.B(_05855_),
    .C(_07009_),
    .A(_05854_),
    .Y(_07010_));
 sg13g2_or3_1 _24869_ (.A(_05848_),
    .B(_05852_),
    .C(_07010_),
    .X(_07011_));
 sg13g2_nor4_1 _24870_ (.A(_05841_),
    .B(_05847_),
    .C(_05875_),
    .D(_07011_),
    .Y(_07012_));
 sg13g2_nand4_1 _24871_ (.B(_05834_),
    .C(_05839_),
    .A(_05817_),
    .Y(_07013_),
    .D(_07012_));
 sg13g2_nor3_2 _24872_ (.A(_05825_),
    .B(_05885_),
    .C(_07013_),
    .Y(_07014_));
 sg13g2_nor4_1 _24873_ (.A(_05841_),
    .B(_05847_),
    .C(_05875_),
    .D(_07011_),
    .Y(_07015_));
 sg13g2_nand3_1 _24874_ (.B(_05834_),
    .C(_07015_),
    .A(_05817_),
    .Y(_07016_));
 sg13g2_or4_2 _24875_ (.A(_05825_),
    .B(_05838_),
    .C(_05885_),
    .D(_07016_),
    .X(_07017_));
 sg13g2_a21oi_1 _24876_ (.A1(net6891),
    .A2(net4549),
    .Y(_07018_),
    .B1(net5987));
 sg13g2_o21ai_1 _24877_ (.B1(_07018_),
    .Y(_02223_),
    .A1(_07945_),
    .A2(net4549));
 sg13g2_a21oi_1 _24878_ (.A1(net3865),
    .A2(net4549),
    .Y(_07019_),
    .B1(net5987));
 sg13g2_o21ai_1 _24879_ (.B1(_07019_),
    .Y(_02224_),
    .A1(_07944_),
    .A2(_07017_));
 sg13g2_a21oi_1 _24880_ (.A1(\atari2600.tia.poly4_l.x[3] ),
    .A2(net4551),
    .Y(_07020_),
    .B1(net5987));
 sg13g2_o21ai_1 _24881_ (.B1(_07020_),
    .Y(_02225_),
    .A1(_07944_),
    .A2(net4551));
 sg13g2_xnor2_1 _24882_ (.Y(_07021_),
    .A(net3865),
    .B(net6891));
 sg13g2_a21oi_1 _24883_ (.A1(net7017),
    .A2(net4549),
    .Y(_07022_),
    .B1(net5987));
 sg13g2_o21ai_1 _24884_ (.B1(_07022_),
    .Y(_02226_),
    .A1(_07017_),
    .A2(_07021_));
 sg13g2_a21oi_1 _24885_ (.A1(\atari2600.tia.p5_l ),
    .A2(net4547),
    .Y(_07023_),
    .B1(net5986));
 sg13g2_o21ai_1 _24886_ (.B1(_07023_),
    .Y(_02227_),
    .A1(_07943_),
    .A2(net4547));
 sg13g2_a21oi_1 _24887_ (.A1(net3930),
    .A2(net4550),
    .Y(_07024_),
    .B1(net5986));
 sg13g2_o21ai_1 _24888_ (.B1(_07024_),
    .Y(_02228_),
    .A1(_07943_),
    .A2(net4550));
 sg13g2_a21oi_1 _24889_ (.A1(net3930),
    .A2(net4547),
    .Y(_07025_),
    .B1(net5986));
 sg13g2_o21ai_1 _24890_ (.B1(_07025_),
    .Y(_02229_),
    .A1(_07942_),
    .A2(net4547));
 sg13g2_a21oi_1 _24891_ (.A1(\atari2600.tia.poly5_l.x[4] ),
    .A2(net4550),
    .Y(_07026_),
    .B1(net5986));
 sg13g2_o21ai_1 _24892_ (.B1(_07026_),
    .Y(_02230_),
    .A1(_07942_),
    .A2(net4550));
 sg13g2_xnor2_1 _24893_ (.Y(_07027_),
    .A(net3930),
    .B(\atari2600.tia.p5_l ));
 sg13g2_a21oi_1 _24894_ (.A1(net6854),
    .A2(net4547),
    .Y(_07028_),
    .B1(net5986));
 sg13g2_o21ai_1 _24895_ (.B1(_07028_),
    .Y(_02231_),
    .A1(net4547),
    .A2(_07027_));
 sg13g2_a21oi_1 _24896_ (.A1(\atari2600.tia.p9_l ),
    .A2(net4549),
    .Y(_07029_),
    .B1(net5985));
 sg13g2_o21ai_1 _24897_ (.B1(_07029_),
    .Y(_02232_),
    .A1(_07941_),
    .A2(net4549));
 sg13g2_a21oi_1 _24898_ (.A1(net3241),
    .A2(net4551),
    .Y(_07030_),
    .B1(net5986));
 sg13g2_o21ai_1 _24899_ (.B1(_07030_),
    .Y(_02233_),
    .A1(_07941_),
    .A2(net4551));
 sg13g2_a21oi_1 _24900_ (.A1(net3241),
    .A2(net4548),
    .Y(_07031_),
    .B1(net5985));
 sg13g2_o21ai_1 _24901_ (.B1(_07031_),
    .Y(_02234_),
    .A1(_07940_),
    .A2(net4548));
 sg13g2_a21oi_1 _24902_ (.A1(net4098),
    .A2(net4550),
    .Y(_07032_),
    .B1(net5985));
 sg13g2_o21ai_1 _24903_ (.B1(_07032_),
    .Y(_02235_),
    .A1(_07940_),
    .A2(net4551));
 sg13g2_a21oi_1 _24904_ (.A1(net4098),
    .A2(net4548),
    .Y(_07033_),
    .B1(net5985));
 sg13g2_o21ai_1 _24905_ (.B1(_07033_),
    .Y(_02236_),
    .A1(_07939_),
    .A2(net4548));
 sg13g2_a21oi_1 _24906_ (.A1(net4187),
    .A2(net4550),
    .Y(_07034_),
    .B1(net5985));
 sg13g2_o21ai_1 _24907_ (.B1(_07034_),
    .Y(_02237_),
    .A1(_07939_),
    .A2(net4550));
 sg13g2_a21oi_1 _24908_ (.A1(net4187),
    .A2(net4547),
    .Y(_07035_),
    .B1(net5985));
 sg13g2_o21ai_1 _24909_ (.B1(_07035_),
    .Y(_02238_),
    .A1(_07938_),
    .A2(net4548));
 sg13g2_a21oi_1 _24910_ (.A1(net3942),
    .A2(net4550),
    .Y(_07036_),
    .B1(net5985));
 sg13g2_o21ai_1 _24911_ (.B1(_07036_),
    .Y(_02239_),
    .A1(_07938_),
    .A2(net4551));
 sg13g2_xnor2_1 _24912_ (.Y(_07037_),
    .A(net4098),
    .B(net7006));
 sg13g2_a21oi_1 _24913_ (.A1(net3942),
    .A2(net4547),
    .Y(_07038_),
    .B1(net5985));
 sg13g2_o21ai_1 _24914_ (.B1(_07038_),
    .Y(_02240_),
    .A1(net4548),
    .A2(_07037_));
 sg13g2_xor2_1 _24915_ (.B(_05819_),
    .A(_00135_),
    .X(_07039_));
 sg13g2_xor2_1 _24916_ (.B(_05832_),
    .A(_00132_),
    .X(_07040_));
 sg13g2_and2_1 _24917_ (.A(_00129_),
    .B(_05845_),
    .X(_07041_));
 sg13g2_nor2_1 _24918_ (.A(_00129_),
    .B(_05845_),
    .Y(_07042_));
 sg13g2_nand2_1 _24919_ (.Y(_07043_),
    .A(_00128_),
    .B(_05843_));
 sg13g2_nor2_1 _24920_ (.A(_00128_),
    .B(_05843_),
    .Y(_07044_));
 sg13g2_or2_1 _24921_ (.X(_07045_),
    .B(_05850_),
    .A(_00127_));
 sg13g2_xnor2_1 _24922_ (.Y(_07046_),
    .A(_00125_),
    .B(_05856_));
 sg13g2_or2_1 _24923_ (.X(_07047_),
    .B(_05865_),
    .A(_00123_));
 sg13g2_o21ai_1 _24924_ (.B1(_08032_),
    .Y(_07048_),
    .A1(\atari2600.tia.audio_right_counter[1] ),
    .A2(_05862_));
 sg13g2_a221oi_1 _24925_ (.B2(_00123_),
    .C1(_07048_),
    .B1(_05865_),
    .A1(\atari2600.tia.audio_right_counter[1] ),
    .Y(_07049_),
    .A2(_05862_));
 sg13g2_xor2_1 _24926_ (.B(_05859_),
    .A(_00124_),
    .X(_07050_));
 sg13g2_nand4_1 _24927_ (.B(_07047_),
    .C(_07049_),
    .A(_07046_),
    .Y(_07051_),
    .D(_07050_));
 sg13g2_a21oi_1 _24928_ (.A1(_00126_),
    .A2(_05853_),
    .Y(_07052_),
    .B1(_07051_));
 sg13g2_nor2_1 _24929_ (.A(_00126_),
    .B(_05853_),
    .Y(_07053_));
 sg13g2_nor2_1 _24930_ (.A(_08105_),
    .B(_05822_),
    .Y(_07054_));
 sg13g2_and2_1 _24931_ (.A(_08105_),
    .B(_05822_),
    .X(_07055_));
 sg13g2_xor2_1 _24932_ (.B(_05829_),
    .A(_00133_),
    .X(_07056_));
 sg13g2_a21oi_1 _24933_ (.A1(_00127_),
    .A2(_05850_),
    .Y(_07057_),
    .B1(_07053_));
 sg13g2_nand4_1 _24934_ (.B(_07045_),
    .C(_07052_),
    .A(_07043_),
    .Y(_07058_),
    .D(_07057_));
 sg13g2_nor4_1 _24935_ (.A(_07041_),
    .B(_07042_),
    .C(_07044_),
    .D(_07058_),
    .Y(_07059_));
 sg13g2_o21ai_1 _24936_ (.B1(_07059_),
    .Y(_07060_),
    .A1(_00130_),
    .A2(_05840_));
 sg13g2_a221oi_1 _24937_ (.B2(_00130_),
    .C1(_07060_),
    .B1(_05840_),
    .A1(_00131_),
    .Y(_07061_),
    .A2(_05836_));
 sg13g2_o21ai_1 _24938_ (.B1(_07061_),
    .Y(_07062_),
    .A1(_00131_),
    .A2(_05836_));
 sg13g2_nor4_1 _24939_ (.A(_07040_),
    .B(_07054_),
    .C(_07055_),
    .D(_07062_),
    .Y(_07063_));
 sg13g2_nand2_1 _24940_ (.Y(_07064_),
    .A(_00136_),
    .B(_05815_));
 sg13g2_and4_1 _24941_ (.A(_07039_),
    .B(_07056_),
    .C(_07063_),
    .D(_07064_),
    .X(_07065_));
 sg13g2_o21ai_1 _24942_ (.B1(_07065_),
    .Y(_07066_),
    .A1(_00136_),
    .A2(_05815_));
 sg13g2_a21oi_1 _24943_ (.A1(\atari2600.tia.p4_r ),
    .A2(net4546),
    .Y(_07067_),
    .B1(net5990));
 sg13g2_o21ai_1 _24944_ (.B1(_07067_),
    .Y(_02241_),
    .A1(_07937_),
    .A2(net4544));
 sg13g2_o21ai_1 _24945_ (.B1(net6036),
    .Y(_07068_),
    .A1(_07936_),
    .A2(net4544));
 sg13g2_a21o_1 _24946_ (.A2(net4544),
    .A1(net6877),
    .B1(_07068_),
    .X(_02242_));
 sg13g2_mux2_1 _24947_ (.A0(net6748),
    .A1(net7001),
    .S(net4544),
    .X(_07069_));
 sg13g2_or2_1 _24948_ (.X(_02243_),
    .B(_07069_),
    .A(net5990));
 sg13g2_nand2_1 _24949_ (.Y(_07070_),
    .A(net6748),
    .B(net4546));
 sg13g2_xor2_1 _24950_ (.B(\atari2600.tia.p4_r ),
    .A(\atari2600.tia.poly4_r.x[1] ),
    .X(_07071_));
 sg13g2_nand2b_1 _24951_ (.Y(_07072_),
    .B(_07071_),
    .A_N(net4546));
 sg13g2_nand3_1 _24952_ (.B(_07070_),
    .C(_07072_),
    .A(net6036),
    .Y(_02244_));
 sg13g2_o21ai_1 _24953_ (.B1(net6038),
    .Y(_07073_),
    .A1(_07935_),
    .A2(net4543));
 sg13g2_a21o_1 _24954_ (.A2(net4543),
    .A1(net7167),
    .B1(_07073_),
    .X(_02245_));
 sg13g2_a21oi_1 _24955_ (.A1(\atari2600.tia.poly5_r.x[1] ),
    .A2(net4543),
    .Y(_07074_),
    .B1(net5990));
 sg13g2_o21ai_1 _24956_ (.B1(_07074_),
    .Y(_02246_),
    .A1(_07934_),
    .A2(net4543));
 sg13g2_o21ai_1 _24957_ (.B1(net6036),
    .Y(_07075_),
    .A1(_07933_),
    .A2(net4543));
 sg13g2_a21o_1 _24958_ (.A2(net4543),
    .A1(net3056),
    .B1(_07075_),
    .X(_02247_));
 sg13g2_mux2_1 _24959_ (.A0(net6872),
    .A1(net7016),
    .S(net4543),
    .X(_07076_));
 sg13g2_or2_1 _24960_ (.X(_02248_),
    .B(_07076_),
    .A(net5990));
 sg13g2_nand2_1 _24961_ (.Y(_07077_),
    .A(net6872),
    .B(net4543));
 sg13g2_xor2_1 _24962_ (.B(\atari2600.tia.p5_r ),
    .A(net3056),
    .X(_07078_));
 sg13g2_nand2b_1 _24963_ (.Y(_07079_),
    .B(_07078_),
    .A_N(net4544));
 sg13g2_nand3_1 _24964_ (.B(_07077_),
    .C(_07079_),
    .A(net6036),
    .Y(_02249_));
 sg13g2_o21ai_1 _24965_ (.B1(net6036),
    .Y(_07080_),
    .A1(_07932_),
    .A2(net4545));
 sg13g2_a21o_1 _24966_ (.A2(net4545),
    .A1(net7240),
    .B1(_07080_),
    .X(_02250_));
 sg13g2_mux2_1 _24967_ (.A0(net7257),
    .A1(\atari2600.tia.poly9_r.x[1] ),
    .S(net4545),
    .X(_07081_));
 sg13g2_or2_1 _24968_ (.X(_02251_),
    .B(net7258),
    .A(net5990));
 sg13g2_mux2_1 _24969_ (.A0(net4414),
    .A1(net7257),
    .S(net4545),
    .X(_07082_));
 sg13g2_or2_1 _24970_ (.X(_02252_),
    .B(_07082_),
    .A(net5990));
 sg13g2_a21oi_1 _24971_ (.A1(net4414),
    .A2(net4545),
    .Y(_07083_),
    .B1(net5990));
 sg13g2_o21ai_1 _24972_ (.B1(_07083_),
    .Y(_02253_),
    .A1(_07931_),
    .A2(net4545));
 sg13g2_o21ai_1 _24973_ (.B1(net6036),
    .Y(_07084_),
    .A1(_07930_),
    .A2(net4546));
 sg13g2_a21o_1 _24974_ (.A2(net4545),
    .A1(net6939),
    .B1(_07084_),
    .X(_02254_));
 sg13g2_mux2_1 _24975_ (.A0(\atari2600.tia.poly9_r.x[6] ),
    .A1(net7264),
    .S(_07066_),
    .X(_07085_));
 sg13g2_or2_1 _24976_ (.X(_02255_),
    .B(net7265),
    .A(net5990));
 sg13g2_mux2_1 _24977_ (.A0(net7259),
    .A1(net7276),
    .S(net4546),
    .X(_07086_));
 sg13g2_or2_1 _24978_ (.X(_02256_),
    .B(_07086_),
    .A(net5991));
 sg13g2_mux2_1 _24979_ (.A0(net4357),
    .A1(net7259),
    .S(net4546),
    .X(_07087_));
 sg13g2_or2_1 _24980_ (.X(_02257_),
    .B(_07087_),
    .A(net5991));
 sg13g2_xor2_1 _24981_ (.B(\atari2600.tia.p9_r ),
    .A(\atari2600.tia.poly9_r.x[4] ),
    .X(_07088_));
 sg13g2_nand2_1 _24982_ (.Y(_07089_),
    .A(net4357),
    .B(net4546));
 sg13g2_nand2b_1 _24983_ (.Y(_07090_),
    .B(_07088_),
    .A_N(net4545));
 sg13g2_nand3_1 _24984_ (.B(_07089_),
    .C(_07090_),
    .A(net6036),
    .Y(_02258_));
 sg13g2_nand2_2 _24985_ (.Y(_07091_),
    .A(net5432),
    .B(_03100_));
 sg13g2_mux2_1 _24986_ (.A0(net5773),
    .A1(net6687),
    .S(_07091_),
    .X(_02259_));
 sg13g2_mux2_1 _24987_ (.A0(net5748),
    .A1(net6547),
    .S(_07091_),
    .X(_02260_));
 sg13g2_mux2_1 _24988_ (.A0(net5717),
    .A1(net6773),
    .S(_07091_),
    .X(_02261_));
 sg13g2_mux2_1 _24989_ (.A0(net5689),
    .A1(net6225),
    .S(_07091_),
    .X(_02262_));
 sg13g2_mux2_1 _24990_ (.A0(net5658),
    .A1(net6837),
    .S(_07091_),
    .X(_02263_));
 sg13g2_mux2_1 _24991_ (.A0(net5629),
    .A1(net6641),
    .S(_07091_),
    .X(_02264_));
 sg13g2_mux2_1 _24992_ (.A0(net5601),
    .A1(net6274),
    .S(_07091_),
    .X(_02265_));
 sg13g2_nand2_2 _24993_ (.Y(_07092_),
    .A(net5469),
    .B(_02995_));
 sg13g2_mux2_1 _24994_ (.A0(net5782),
    .A1(net6821),
    .S(_07092_),
    .X(_02266_));
 sg13g2_mux2_1 _24995_ (.A0(net5753),
    .A1(net4501),
    .S(_07092_),
    .X(_02267_));
 sg13g2_mux2_1 _24996_ (.A0(net5724),
    .A1(net6453),
    .S(_07092_),
    .X(_02268_));
 sg13g2_mux2_1 _24997_ (.A0(net5695),
    .A1(net6270),
    .S(_07092_),
    .X(_02269_));
 sg13g2_mux2_1 _24998_ (.A0(net5667),
    .A1(net6719),
    .S(_07092_),
    .X(_02270_));
 sg13g2_mux2_1 _24999_ (.A0(net5638),
    .A1(net6268),
    .S(_07092_),
    .X(_02271_));
 sg13g2_mux2_1 _25000_ (.A0(net5607),
    .A1(net6846),
    .S(_07092_),
    .X(_02272_));
 sg13g2_nand2_2 _25001_ (.Y(_07093_),
    .A(net5431),
    .B(net5419));
 sg13g2_mux2_1 _25002_ (.A0(net5773),
    .A1(net6863),
    .S(_07093_),
    .X(_02273_));
 sg13g2_mux2_1 _25003_ (.A0(net5747),
    .A1(net6549),
    .S(_07093_),
    .X(_02274_));
 sg13g2_mux2_1 _25004_ (.A0(net5717),
    .A1(net6162),
    .S(_07093_),
    .X(_02275_));
 sg13g2_mux2_1 _25005_ (.A0(net5689),
    .A1(net6256),
    .S(_07093_),
    .X(_02276_));
 sg13g2_mux2_1 _25006_ (.A0(net5658),
    .A1(net6664),
    .S(_07093_),
    .X(_02277_));
 sg13g2_mux2_1 _25007_ (.A0(net5628),
    .A1(net6394),
    .S(_07093_),
    .X(_02278_));
 sg13g2_mux2_1 _25008_ (.A0(net5601),
    .A1(net6583),
    .S(_07093_),
    .X(_02279_));
 sg13g2_nand2_2 _25009_ (.Y(_07094_),
    .A(net5469),
    .B(_03118_));
 sg13g2_mux2_1 _25010_ (.A0(net5785),
    .A1(net6868),
    .S(_07094_),
    .X(_02280_));
 sg13g2_mux2_1 _25011_ (.A0(net5753),
    .A1(net4322),
    .S(_07094_),
    .X(_02281_));
 sg13g2_mux2_1 _25012_ (.A0(net5724),
    .A1(net6306),
    .S(_07094_),
    .X(_02282_));
 sg13g2_mux2_1 _25013_ (.A0(net5695),
    .A1(net6974),
    .S(_07094_),
    .X(_02283_));
 sg13g2_mux2_1 _25014_ (.A0(net5668),
    .A1(net6505),
    .S(_07094_),
    .X(_02284_));
 sg13g2_mux2_1 _25015_ (.A0(net5638),
    .A1(net6586),
    .S(_07094_),
    .X(_02285_));
 sg13g2_mux2_1 _25016_ (.A0(net5609),
    .A1(net6677),
    .S(_07094_),
    .X(_02286_));
 sg13g2_nor2_2 _25017_ (.A(_10481_),
    .B(net5471),
    .Y(_07095_));
 sg13g2_mux2_1 _25018_ (.A0(net3874),
    .A1(net5790),
    .S(_07095_),
    .X(_02287_));
 sg13g2_mux2_1 _25019_ (.A0(net3408),
    .A1(net5756),
    .S(_07095_),
    .X(_02288_));
 sg13g2_mux2_1 _25020_ (.A0(net3565),
    .A1(net5727),
    .S(_07095_),
    .X(_02289_));
 sg13g2_mux2_1 _25021_ (.A0(net3221),
    .A1(net5698),
    .S(_07095_),
    .X(_02290_));
 sg13g2_mux2_1 _25022_ (.A0(net3882),
    .A1(net5670),
    .S(_07095_),
    .X(_02291_));
 sg13g2_mux2_1 _25023_ (.A0(net3939),
    .A1(net5647),
    .S(_07095_),
    .X(_02292_));
 sg13g2_mux2_1 _25024_ (.A0(net3138),
    .A1(net5613),
    .S(_07095_),
    .X(_02293_));
 sg13g2_nor2_2 _25025_ (.A(net5473),
    .B(net5425),
    .Y(_07096_));
 sg13g2_mux2_1 _25026_ (.A0(net3556),
    .A1(net5790),
    .S(_07096_),
    .X(_02294_));
 sg13g2_mux2_1 _25027_ (.A0(net3571),
    .A1(net5756),
    .S(_07096_),
    .X(_02295_));
 sg13g2_mux2_1 _25028_ (.A0(net3597),
    .A1(net5727),
    .S(_07096_),
    .X(_02296_));
 sg13g2_mux2_1 _25029_ (.A0(net3648),
    .A1(net5698),
    .S(_07096_),
    .X(_02297_));
 sg13g2_mux2_1 _25030_ (.A0(net3467),
    .A1(net5670),
    .S(_07096_),
    .X(_02298_));
 sg13g2_mux2_1 _25031_ (.A0(net3732),
    .A1(net5646),
    .S(_07096_),
    .X(_02299_));
 sg13g2_mux2_1 _25032_ (.A0(net3511),
    .A1(net5613),
    .S(_07096_),
    .X(_02300_));
 sg13g2_nor3_1 _25033_ (.A(\atari2600.pia.interval[0] ),
    .B(net5977),
    .C(net4580),
    .Y(_07097_));
 sg13g2_a221oi_1 _25034_ (.B2(net4580),
    .C1(_07097_),
    .B1(_08676_),
    .A1(_08039_),
    .Y(_02301_),
    .A2(net5977));
 sg13g2_nand2_2 _25035_ (.Y(_07098_),
    .A(_10372_),
    .B(net5422));
 sg13g2_mux2_1 _25036_ (.A0(net5781),
    .A1(net6722),
    .S(_07098_),
    .X(_02302_));
 sg13g2_mux2_1 _25037_ (.A0(net5752),
    .A1(net6265),
    .S(_07098_),
    .X(_02303_));
 sg13g2_mux2_1 _25038_ (.A0(net5722),
    .A1(net6540),
    .S(_07098_),
    .X(_02304_));
 sg13g2_mux2_1 _25039_ (.A0(net5693),
    .A1(net4413),
    .S(_07098_),
    .X(_02305_));
 sg13g2_mux2_1 _25040_ (.A0(net5665),
    .A1(net6782),
    .S(_07098_),
    .X(_02306_));
 sg13g2_mux2_1 _25041_ (.A0(net5638),
    .A1(net4493),
    .S(_07098_),
    .X(_02307_));
 sg13g2_mux2_1 _25042_ (.A0(net5607),
    .A1(net6596),
    .S(_07098_),
    .X(_02308_));
 sg13g2_nand3_1 _25043_ (.B(_03163_),
    .C(_05250_),
    .A(_08583_),
    .Y(_07099_));
 sg13g2_nand3_1 _25044_ (.B(net5209),
    .C(_07099_),
    .A(net3155),
    .Y(_07100_));
 sg13g2_nand2b_1 _25045_ (.Y(_02309_),
    .B(_07100_),
    .A_N(_05247_));
 sg13g2_nand2_2 _25046_ (.Y(_07101_),
    .A(net5422),
    .B(_03124_));
 sg13g2_mux2_1 _25047_ (.A0(net5781),
    .A1(net6729),
    .S(_07101_),
    .X(_02310_));
 sg13g2_mux2_1 _25048_ (.A0(net5752),
    .A1(net6708),
    .S(_07101_),
    .X(_02311_));
 sg13g2_mux2_1 _25049_ (.A0(net5722),
    .A1(net4286),
    .S(_07101_),
    .X(_02312_));
 sg13g2_mux2_1 _25050_ (.A0(net5693),
    .A1(net6496),
    .S(_07101_),
    .X(_02313_));
 sg13g2_mux2_1 _25051_ (.A0(net5665),
    .A1(net6143),
    .S(_07101_),
    .X(_02314_));
 sg13g2_mux2_1 _25052_ (.A0(net5638),
    .A1(net4417),
    .S(_07101_),
    .X(_02315_));
 sg13g2_mux2_1 _25053_ (.A0(net5607),
    .A1(net4377),
    .S(_07101_),
    .X(_02316_));
 sg13g2_nand2_2 _25054_ (.Y(_07102_),
    .A(net5431),
    .B(net5416));
 sg13g2_mux2_1 _25055_ (.A0(net5773),
    .A1(net6680),
    .S(_07102_),
    .X(_02317_));
 sg13g2_mux2_1 _25056_ (.A0(net5748),
    .A1(net6377),
    .S(_07102_),
    .X(_02318_));
 sg13g2_mux2_1 _25057_ (.A0(net5717),
    .A1(net6838),
    .S(_07102_),
    .X(_02319_));
 sg13g2_mux2_1 _25058_ (.A0(net5688),
    .A1(net6813),
    .S(_07102_),
    .X(_02320_));
 sg13g2_mux2_1 _25059_ (.A0(net5658),
    .A1(net6967),
    .S(_07102_),
    .X(_02321_));
 sg13g2_mux2_1 _25060_ (.A0(net5628),
    .A1(net6056),
    .S(_07102_),
    .X(_02322_));
 sg13g2_mux2_1 _25061_ (.A0(net5601),
    .A1(net4442),
    .S(_07102_),
    .X(_02323_));
 sg13g2_nand2_2 _25062_ (.Y(_07103_),
    .A(net5431),
    .B(net5424));
 sg13g2_mux2_1 _25063_ (.A0(net5773),
    .A1(net6666),
    .S(_07103_),
    .X(_02324_));
 sg13g2_mux2_1 _25064_ (.A0(net5748),
    .A1(net4515),
    .S(_07103_),
    .X(_02325_));
 sg13g2_mux2_1 _25065_ (.A0(net5716),
    .A1(net6776),
    .S(_07103_),
    .X(_02326_));
 sg13g2_mux2_1 _25066_ (.A0(net5689),
    .A1(net6606),
    .S(_07103_),
    .X(_02327_));
 sg13g2_mux2_1 _25067_ (.A0(net5658),
    .A1(net6475),
    .S(_07103_),
    .X(_02328_));
 sg13g2_mux2_1 _25068_ (.A0(net5629),
    .A1(net6499),
    .S(_07103_),
    .X(_02329_));
 sg13g2_mux2_1 _25069_ (.A0(net5601),
    .A1(net6625),
    .S(_07103_),
    .X(_02330_));
 sg13g2_nor4_2 _25070_ (.A(net5038),
    .B(net4876),
    .C(net5027),
    .Y(_07104_),
    .D(net5021));
 sg13g2_nand2_2 _25071_ (.Y(_07105_),
    .A(net4748),
    .B(_07104_));
 sg13g2_mux2_1 _25072_ (.A0(net5244),
    .A1(net6620),
    .S(_07105_),
    .X(_02331_));
 sg13g2_mux2_1 _25073_ (.A0(net5218),
    .A1(net4391),
    .S(_07105_),
    .X(_02332_));
 sg13g2_mux2_1 _25074_ (.A0(net5115),
    .A1(net6976),
    .S(_07105_),
    .X(_02333_));
 sg13g2_mux2_1 _25075_ (.A0(net5088),
    .A1(net6817),
    .S(_07105_),
    .X(_02334_));
 sg13g2_mux2_1 _25076_ (.A0(net5185),
    .A1(net4457),
    .S(_07105_),
    .X(_02335_));
 sg13g2_mux2_1 _25077_ (.A0(net5157),
    .A1(net6474),
    .S(_07105_),
    .X(_02336_));
 sg13g2_mux2_1 _25078_ (.A0(net5068),
    .A1(net6392),
    .S(_07105_),
    .X(_02337_));
 sg13g2_mux2_1 _25079_ (.A0(net5040),
    .A1(net4421),
    .S(_07105_),
    .X(_02338_));
 sg13g2_nor2b_1 _25080_ (.A(net4741),
    .B_N(_07104_),
    .Y(_07106_));
 sg13g2_nor2_1 _25081_ (.A(net3051),
    .B(net4650),
    .Y(_07107_));
 sg13g2_a21oi_1 _25082_ (.A1(net5260),
    .A2(net4650),
    .Y(_02339_),
    .B1(_07107_));
 sg13g2_nor2_1 _25083_ (.A(net3798),
    .B(net4651),
    .Y(_07108_));
 sg13g2_a21oi_1 _25084_ (.A1(net5234),
    .A2(net4651),
    .Y(_02340_),
    .B1(_07108_));
 sg13g2_nor2_1 _25085_ (.A(net3186),
    .B(net4650),
    .Y(_07109_));
 sg13g2_a21oi_1 _25086_ (.A1(net5131),
    .A2(net4650),
    .Y(_02341_),
    .B1(_07109_));
 sg13g2_nor2_1 _25087_ (.A(net3279),
    .B(net4650),
    .Y(_07110_));
 sg13g2_a21oi_1 _25088_ (.A1(net5103),
    .A2(net4650),
    .Y(_02342_),
    .B1(_07110_));
 sg13g2_nor2_1 _25089_ (.A(net3151),
    .B(net4651),
    .Y(_07111_));
 sg13g2_a21oi_1 _25090_ (.A1(net5173),
    .A2(net4651),
    .Y(_02343_),
    .B1(_07111_));
 sg13g2_nor2_1 _25091_ (.A(net3921),
    .B(net4651),
    .Y(_07112_));
 sg13g2_a21oi_1 _25092_ (.A1(net5146),
    .A2(net4651),
    .Y(_02344_),
    .B1(_07112_));
 sg13g2_nor2_1 _25093_ (.A(net3452),
    .B(net4651),
    .Y(_07113_));
 sg13g2_a21oi_1 _25094_ (.A1(net5078),
    .A2(net4651),
    .Y(_02345_),
    .B1(_07113_));
 sg13g2_nor2_1 _25095_ (.A(net3875),
    .B(net4650),
    .Y(_07114_));
 sg13g2_a21oi_1 _25096_ (.A1(net5055),
    .A2(net4650),
    .Y(_02346_),
    .B1(_07114_));
 sg13g2_nand2_2 _25097_ (.Y(_07115_),
    .A(net4737),
    .B(_07104_));
 sg13g2_mux2_1 _25098_ (.A0(net5244),
    .A1(net4021),
    .S(_07115_),
    .X(_02347_));
 sg13g2_mux2_1 _25099_ (.A0(net5218),
    .A1(net6139),
    .S(_07115_),
    .X(_02348_));
 sg13g2_mux2_1 _25100_ (.A0(net5116),
    .A1(net4188),
    .S(_07115_),
    .X(_02349_));
 sg13g2_mux2_1 _25101_ (.A0(net5088),
    .A1(net4068),
    .S(_07115_),
    .X(_02350_));
 sg13g2_mux2_1 _25102_ (.A0(net5185),
    .A1(net4028),
    .S(_07115_),
    .X(_02351_));
 sg13g2_mux2_1 _25103_ (.A0(net5157),
    .A1(net4069),
    .S(_07115_),
    .X(_02352_));
 sg13g2_mux2_1 _25104_ (.A0(net5065),
    .A1(net4241),
    .S(_07115_),
    .X(_02353_));
 sg13g2_mux2_1 _25105_ (.A0(net5040),
    .A1(net4107),
    .S(_07115_),
    .X(_02354_));
 sg13g2_nand2_2 _25106_ (.Y(_07116_),
    .A(net4733),
    .B(_07104_));
 sg13g2_mux2_1 _25107_ (.A0(net5244),
    .A1(net4463),
    .S(_07116_),
    .X(_02355_));
 sg13g2_mux2_1 _25108_ (.A0(net5218),
    .A1(net4125),
    .S(_07116_),
    .X(_02356_));
 sg13g2_mux2_1 _25109_ (.A0(net5116),
    .A1(net7077),
    .S(_07116_),
    .X(_02357_));
 sg13g2_mux2_1 _25110_ (.A0(net5089),
    .A1(net4033),
    .S(_07116_),
    .X(_02358_));
 sg13g2_mux2_1 _25111_ (.A0(net5185),
    .A1(net4489),
    .S(_07116_),
    .X(_02359_));
 sg13g2_mux2_1 _25112_ (.A0(net5157),
    .A1(net4281),
    .S(_07116_),
    .X(_02360_));
 sg13g2_mux2_1 _25113_ (.A0(net5064),
    .A1(net4250),
    .S(_07116_),
    .X(_02361_));
 sg13g2_mux2_1 _25114_ (.A0(net5040),
    .A1(net4108),
    .S(_07116_),
    .X(_02362_));
 sg13g2_nor2_2 _25115_ (.A(_03042_),
    .B(net4741),
    .Y(_07117_));
 sg13g2_nor2_1 _25116_ (.A(net3230),
    .B(net4648),
    .Y(_07118_));
 sg13g2_a21oi_1 _25117_ (.A1(net5261),
    .A2(net4648),
    .Y(_02363_),
    .B1(_07118_));
 sg13g2_nor2_1 _25118_ (.A(net3075),
    .B(net4649),
    .Y(_07119_));
 sg13g2_a21oi_1 _25119_ (.A1(net5235),
    .A2(net4649),
    .Y(_02364_),
    .B1(_07119_));
 sg13g2_nor2_1 _25120_ (.A(net3076),
    .B(net4649),
    .Y(_07120_));
 sg13g2_a21oi_1 _25121_ (.A1(net5134),
    .A2(net4649),
    .Y(_02365_),
    .B1(_07120_));
 sg13g2_nor2_1 _25122_ (.A(net3772),
    .B(net4649),
    .Y(_07121_));
 sg13g2_a21oi_1 _25123_ (.A1(net5105),
    .A2(net4649),
    .Y(_02366_),
    .B1(_07121_));
 sg13g2_nor2_1 _25124_ (.A(net3971),
    .B(net4649),
    .Y(_07122_));
 sg13g2_a21oi_1 _25125_ (.A1(net5178),
    .A2(net4649),
    .Y(_02367_),
    .B1(_07122_));
 sg13g2_nor2_1 _25126_ (.A(net2994),
    .B(net4648),
    .Y(_07123_));
 sg13g2_a21oi_1 _25127_ (.A1(net5148),
    .A2(net4648),
    .Y(_02368_),
    .B1(_07123_));
 sg13g2_nor2_1 _25128_ (.A(net3237),
    .B(net4648),
    .Y(_07124_));
 sg13g2_a21oi_1 _25129_ (.A1(net5080),
    .A2(net4648),
    .Y(_02369_),
    .B1(_07124_));
 sg13g2_nor2_1 _25130_ (.A(net3407),
    .B(net4648),
    .Y(_07125_));
 sg13g2_a21oi_1 _25131_ (.A1(net5057),
    .A2(net4648),
    .Y(_02370_),
    .B1(_07125_));
 sg13g2_nand2_2 _25132_ (.Y(_07126_),
    .A(_08514_),
    .B(_05028_));
 sg13g2_mux2_1 _25133_ (.A0(_05031_),
    .A1(net3557),
    .S(_07126_),
    .X(_02371_));
 sg13g2_mux2_1 _25134_ (.A0(_05038_),
    .A1(net3491),
    .S(_07126_),
    .X(_02372_));
 sg13g2_mux2_1 _25135_ (.A0(_05044_),
    .A1(net6804),
    .S(_07126_),
    .X(_02373_));
 sg13g2_mux2_1 _25136_ (.A0(_05049_),
    .A1(net4231),
    .S(_07126_),
    .X(_02374_));
 sg13g2_mux2_1 _25137_ (.A0(_05051_),
    .A1(net4387),
    .S(_07126_),
    .X(_02375_));
 sg13g2_mux2_1 _25138_ (.A0(_05057_),
    .A1(net6843),
    .S(_07126_),
    .X(_02376_));
 sg13g2_mux2_1 _25139_ (.A0(_05063_),
    .A1(net4253),
    .S(_07126_),
    .X(_02377_));
 sg13g2_mux2_1 _25140_ (.A0(_05068_),
    .A1(net4276),
    .S(_07126_),
    .X(_02378_));
 sg13g2_nor3_1 _25141_ (.A(_08565_),
    .B(_08637_),
    .C(net4954),
    .Y(_07127_));
 sg13g2_nand3_1 _25142_ (.B(_08579_),
    .C(_08636_),
    .A(net5036),
    .Y(_07128_));
 sg13g2_o21ai_1 _25143_ (.B1(net6009),
    .Y(_07129_),
    .A1(net7049),
    .A2(_07127_));
 sg13g2_a21oi_1 _25144_ (.A1(net5179),
    .A2(_07127_),
    .Y(_02379_),
    .B1(_07129_));
 sg13g2_o21ai_1 _25145_ (.B1(net6016),
    .Y(_07130_),
    .A1(net5172),
    .A2(_07128_));
 sg13g2_a21oi_1 _25146_ (.A1(_07929_),
    .A2(_07128_),
    .Y(_02380_),
    .B1(_07130_));
 sg13g2_o21ai_1 _25147_ (.B1(net6011),
    .Y(_07131_),
    .A1(net5073),
    .A2(_07128_));
 sg13g2_a21oi_1 _25148_ (.A1(_07928_),
    .A2(_07128_),
    .Y(_02381_),
    .B1(_07131_));
 sg13g2_o21ai_1 _25149_ (.B1(net6011),
    .Y(_07132_),
    .A1(net5054),
    .A2(_07128_));
 sg13g2_a21oi_1 _25150_ (.A1(_07927_),
    .A2(_07128_),
    .Y(_02382_),
    .B1(_07132_));
 sg13g2_nor3_1 _25151_ (.A(net4751),
    .B(net4954),
    .C(_08735_),
    .Y(_07133_));
 sg13g2_nand2_1 _25152_ (.Y(_07134_),
    .A(net5059),
    .B(_07133_));
 sg13g2_o21ai_1 _25153_ (.B1(_07134_),
    .Y(_07135_),
    .A1(net7070),
    .A2(net4647));
 sg13g2_nor2_1 _25154_ (.A(net5984),
    .B(_07135_),
    .Y(_02383_));
 sg13g2_nand2_1 _25155_ (.Y(_07136_),
    .A(net5086),
    .B(net4646));
 sg13g2_o21ai_1 _25156_ (.B1(_07136_),
    .Y(_07137_),
    .A1(net7007),
    .A2(net4646));
 sg13g2_nor2_1 _25157_ (.A(net5984),
    .B(_07137_),
    .Y(_02384_));
 sg13g2_o21ai_1 _25158_ (.B1(net6009),
    .Y(_07138_),
    .A1(net6942),
    .A2(net4646));
 sg13g2_a21oi_1 _25159_ (.A1(net5151),
    .A2(net4646),
    .Y(_02385_),
    .B1(_07138_));
 sg13g2_o21ai_1 _25160_ (.B1(net6011),
    .Y(_07139_),
    .A1(net7010),
    .A2(net4646));
 sg13g2_a21oi_1 _25161_ (.A1(net5180),
    .A2(net4646),
    .Y(_02386_),
    .B1(_07139_));
 sg13g2_o21ai_1 _25162_ (.B1(net6016),
    .Y(_07140_),
    .A1(net7099),
    .A2(net4647));
 sg13g2_a21oi_1 _25163_ (.A1(net5107),
    .A2(net4647),
    .Y(_02387_),
    .B1(_07140_));
 sg13g2_o21ai_1 _25164_ (.B1(net6016),
    .Y(_07141_),
    .A1(net6170),
    .A2(net4647));
 sg13g2_a21oi_1 _25165_ (.A1(net5135),
    .A2(net4647),
    .Y(_02388_),
    .B1(_07141_));
 sg13g2_o21ai_1 _25166_ (.B1(net6009),
    .Y(_07142_),
    .A1(net7067),
    .A2(net4647));
 sg13g2_a21oi_1 _25167_ (.A1(net5239),
    .A2(net4647),
    .Y(_02389_),
    .B1(_07142_));
 sg13g2_o21ai_1 _25168_ (.B1(net6009),
    .Y(_07143_),
    .A1(net7050),
    .A2(net4646));
 sg13g2_a21oi_1 _25169_ (.A1(net5265),
    .A2(net4646),
    .Y(_02390_),
    .B1(_07143_));
 sg13g2_nand2_2 _25170_ (.Y(_07144_),
    .A(_08511_),
    .B(_05028_));
 sg13g2_mux2_1 _25171_ (.A0(_05031_),
    .A1(net3501),
    .S(_07144_),
    .X(_02391_));
 sg13g2_mux2_1 _25172_ (.A0(_05038_),
    .A1(net3749),
    .S(_07144_),
    .X(_02392_));
 sg13g2_mux2_1 _25173_ (.A0(_05044_),
    .A1(net4454),
    .S(_07144_),
    .X(_02393_));
 sg13g2_mux2_1 _25174_ (.A0(_05049_),
    .A1(net4112),
    .S(_07144_),
    .X(_02394_));
 sg13g2_mux2_1 _25175_ (.A0(_05051_),
    .A1(net4283),
    .S(_07144_),
    .X(_02395_));
 sg13g2_mux2_1 _25176_ (.A0(_05057_),
    .A1(net6372),
    .S(_07144_),
    .X(_02396_));
 sg13g2_mux2_1 _25177_ (.A0(_05063_),
    .A1(net6550),
    .S(_07144_),
    .X(_02397_));
 sg13g2_mux2_1 _25178_ (.A0(_05068_),
    .A1(net6707),
    .S(_07144_),
    .X(_02398_));
 sg13g2_nand2_2 _25179_ (.Y(_07145_),
    .A(_03041_),
    .B(net4740));
 sg13g2_mux2_1 _25180_ (.A0(net5248),
    .A1(net4184),
    .S(_07145_),
    .X(_02399_));
 sg13g2_mux2_1 _25181_ (.A0(net5222),
    .A1(net6712),
    .S(_07145_),
    .X(_02400_));
 sg13g2_mux2_1 _25182_ (.A0(net5118),
    .A1(net4194),
    .S(_07145_),
    .X(_02401_));
 sg13g2_mux2_1 _25183_ (.A0(net5094),
    .A1(net4325),
    .S(_07145_),
    .X(_02402_));
 sg13g2_mux2_1 _25184_ (.A0(net5188),
    .A1(net4196),
    .S(_07145_),
    .X(_02403_));
 sg13g2_mux2_1 _25185_ (.A0(net5159),
    .A1(net4012),
    .S(_07145_),
    .X(_02404_));
 sg13g2_mux2_1 _25186_ (.A0(net5066),
    .A1(net4161),
    .S(_07145_),
    .X(_02405_));
 sg13g2_mux2_1 _25187_ (.A0(net5044),
    .A1(net4051),
    .S(_07145_),
    .X(_02406_));
 sg13g2_nor2_2 _25188_ (.A(_10417_),
    .B(_10425_),
    .Y(_07146_));
 sg13g2_nor2_2 _25189_ (.A(net4760),
    .B(_07146_),
    .Y(_07147_));
 sg13g2_mux2_1 _25190_ (.A0(\atari2600.rom_data[0] ),
    .A1(net6691),
    .S(net4781),
    .X(_07148_));
 sg13g2_a22oi_1 _25191_ (.Y(_07149_),
    .B1(_07147_),
    .B2(net6692),
    .A2(net4761),
    .A1(net4019));
 sg13g2_inv_1 _25192_ (.Y(_02407_),
    .A(_07149_));
 sg13g2_mux2_1 _25193_ (.A0(net4229),
    .A1(net7065),
    .S(net4781),
    .X(_07150_));
 sg13g2_a22oi_1 _25194_ (.Y(_07151_),
    .B1(_07147_),
    .B2(_07150_),
    .A2(net4760),
    .A1(net3987));
 sg13g2_inv_1 _25195_ (.Y(_02408_),
    .A(_07151_));
 sg13g2_mux2_1 _25196_ (.A0(\atari2600.rom_data[2] ),
    .A1(net6066),
    .S(_10424_),
    .X(_07152_));
 sg13g2_a22oi_1 _25197_ (.Y(_07153_),
    .B1(_07147_),
    .B2(net6067),
    .A2(net4760),
    .A1(net3313));
 sg13g2_inv_1 _25198_ (.Y(_02409_),
    .A(_07153_));
 sg13g2_mux2_1 _25199_ (.A0(net3958),
    .A1(net6946),
    .S(net4781),
    .X(_07154_));
 sg13g2_a22oi_1 _25200_ (.Y(_07155_),
    .B1(_07147_),
    .B2(_07154_),
    .A2(net4760),
    .A1(net6223));
 sg13g2_inv_1 _25201_ (.Y(_02410_),
    .A(_07155_));
 sg13g2_mux2_1 _25202_ (.A0(net3172),
    .A1(\atari2600.ram_data[4] ),
    .S(net4781),
    .X(_07156_));
 sg13g2_a22oi_1 _25203_ (.Y(_07157_),
    .B1(_07147_),
    .B2(_07156_),
    .A2(net4761),
    .A1(net6599));
 sg13g2_inv_1 _25204_ (.Y(_02411_),
    .A(net6600));
 sg13g2_mux2_1 _25205_ (.A0(net3001),
    .A1(\atari2600.ram_data[5] ),
    .S(net4781),
    .X(_07158_));
 sg13g2_a22oi_1 _25206_ (.Y(_07159_),
    .B1(_07147_),
    .B2(_07158_),
    .A2(net4760),
    .A1(net4532));
 sg13g2_inv_1 _25207_ (.Y(_02412_),
    .A(net4533));
 sg13g2_a21oi_1 _25208_ (.A1(net3965),
    .A2(_10425_),
    .Y(_07160_),
    .B1(net4760));
 sg13g2_a22oi_1 _25209_ (.Y(_07161_),
    .B1(_07146_),
    .B2(net2956),
    .A2(_03006_),
    .A1(net7031));
 sg13g2_a22oi_1 _25210_ (.Y(_02413_),
    .B1(_07160_),
    .B2(_07161_),
    .A2(net4761),
    .A1(_08125_));
 sg13g2_a21oi_1 _25211_ (.A1(net3354),
    .A2(_10425_),
    .Y(_07162_),
    .B1(net4760));
 sg13g2_a22oi_1 _25212_ (.Y(_07163_),
    .B1(_07146_),
    .B2(net2972),
    .A2(_03006_),
    .A1(net7224));
 sg13g2_a22oi_1 _25213_ (.Y(_02414_),
    .B1(_07162_),
    .B2(_07163_),
    .A2(net4760),
    .A1(_08126_));
 sg13g2_nor2_1 _25214_ (.A(net7002),
    .B(net5362),
    .Y(_07164_));
 sg13g2_a21oi_1 _25215_ (.A1(net5362),
    .A2(net5274),
    .Y(_02415_),
    .B1(_07164_));
 sg13g2_nor2_1 _25216_ (.A(net7113),
    .B(net5362),
    .Y(_07165_));
 sg13g2_a21oi_1 _25217_ (.A1(net5362),
    .A2(net5199),
    .Y(_02416_),
    .B1(_07165_));
 sg13g2_nor2_1 _25218_ (.A(net6962),
    .B(net5362),
    .Y(_07166_));
 sg13g2_a21oi_1 _25219_ (.A1(net5362),
    .A2(net5204),
    .Y(_02417_),
    .B1(_07166_));
 sg13g2_nand2_1 _25220_ (.Y(_07167_),
    .A(net5577),
    .B(net5346));
 sg13g2_o21ai_1 _25221_ (.B1(_07167_),
    .Y(_02418_),
    .A1(_08219_),
    .A2(_08259_));
 sg13g2_nand3_1 _25222_ (.B(net5199),
    .C(_08405_),
    .A(net5272),
    .Y(_07168_));
 sg13g2_o21ai_1 _25223_ (.B1(_07168_),
    .Y(_02419_),
    .A1(_08075_),
    .A2(net5271));
 sg13g2_nand4_1 _25224_ (.B(net5270),
    .C(_08216_),
    .A(net5204),
    .Y(_07169_),
    .D(net5199));
 sg13g2_nor3_1 _25225_ (.A(_08175_),
    .B(net5203),
    .C(_07169_),
    .Y(_07170_));
 sg13g2_a21o_1 _25226_ (.A2(net5348),
    .A1(net3970),
    .B1(_07170_),
    .X(_02420_));
 sg13g2_nor3_1 _25227_ (.A(net5274),
    .B(net5203),
    .C(_07169_),
    .Y(_07171_));
 sg13g2_a21o_1 _25228_ (.A2(net5346),
    .A1(net4102),
    .B1(_07171_),
    .X(_02421_));
 sg13g2_nand2_1 _25229_ (.Y(_07172_),
    .A(net2923),
    .B(net5346));
 sg13g2_nor2_2 _25230_ (.A(net5204),
    .B(_08247_),
    .Y(_07173_));
 sg13g2_nand2b_2 _25231_ (.Y(_07174_),
    .B(_08246_),
    .A_N(net5206));
 sg13g2_nand2_1 _25232_ (.Y(_07175_),
    .A(_08216_),
    .B(_07173_));
 sg13g2_nand2_1 _25233_ (.Y(_07176_),
    .A(net5274),
    .B(_08382_));
 sg13g2_o21ai_1 _25234_ (.B1(_07172_),
    .Y(_02422_),
    .A1(_07175_),
    .A2(_07176_));
 sg13g2_nand2_1 _25235_ (.Y(_07177_),
    .A(net2966),
    .B(net5346));
 sg13g2_nand2_1 _25236_ (.Y(_07178_),
    .A(_08175_),
    .B(_08382_));
 sg13g2_o21ai_1 _25237_ (.B1(_07177_),
    .Y(_02423_),
    .A1(_07175_),
    .A2(_07178_));
 sg13g2_nand2_1 _25238_ (.Y(_07179_),
    .A(net2983),
    .B(net5347));
 sg13g2_nand3_1 _25239_ (.B(_08216_),
    .C(_08246_),
    .A(net5206),
    .Y(_07180_));
 sg13g2_o21ai_1 _25240_ (.B1(_07179_),
    .Y(_02424_),
    .A1(_07176_),
    .A2(_07180_));
 sg13g2_nand2_1 _25241_ (.Y(_07181_),
    .A(net3028),
    .B(net5348));
 sg13g2_o21ai_1 _25242_ (.B1(_07181_),
    .Y(_02425_),
    .A1(_07178_),
    .A2(_07180_));
 sg13g2_nand2_2 _25243_ (.Y(_07182_),
    .A(net5423),
    .B(_03100_));
 sg13g2_mux2_1 _25244_ (.A0(net5789),
    .A1(net6874),
    .S(_07182_),
    .X(_02426_));
 sg13g2_mux2_1 _25245_ (.A0(net5755),
    .A1(net4491),
    .S(_07182_),
    .X(_02427_));
 sg13g2_mux2_1 _25246_ (.A0(net5723),
    .A1(net6611),
    .S(_07182_),
    .X(_02428_));
 sg13g2_mux2_1 _25247_ (.A0(net5694),
    .A1(net6100),
    .S(_07182_),
    .X(_02429_));
 sg13g2_mux2_1 _25248_ (.A0(net5665),
    .A1(net6717),
    .S(_07182_),
    .X(_02430_));
 sg13g2_mux2_1 _25249_ (.A0(net5640),
    .A1(net6897),
    .S(_07182_),
    .X(_02431_));
 sg13g2_mux2_1 _25250_ (.A0(net5608),
    .A1(net4389),
    .S(_07182_),
    .X(_02432_));
 sg13g2_nand2_1 _25251_ (.Y(_07183_),
    .A(net7004),
    .B(net5348));
 sg13g2_nor2_1 _25252_ (.A(net5206),
    .B(_08246_),
    .Y(_07184_));
 sg13g2_nand2b_1 _25253_ (.Y(_07185_),
    .B(net5199),
    .A_N(net5205));
 sg13g2_nor2_2 _25254_ (.A(net5275),
    .B(_07185_),
    .Y(_07186_));
 sg13g2_nand2_1 _25255_ (.Y(_07187_),
    .A(_08183_),
    .B(_07186_));
 sg13g2_o21ai_1 _25256_ (.B1(_07183_),
    .Y(_02433_),
    .A1(_08219_),
    .A2(_07187_));
 sg13g2_mux2_1 _25257_ (.A0(net6992),
    .A1(_08450_),
    .S(net5270),
    .X(_02434_));
 sg13g2_nand2_1 _25258_ (.Y(_07188_),
    .A(net6841),
    .B(net5348));
 sg13g2_nor2b_1 _25259_ (.A(_08223_),
    .B_N(_08446_),
    .Y(_07189_));
 sg13g2_nand3_1 _25260_ (.B(net5272),
    .C(_07189_),
    .A(net5205),
    .Y(_07190_));
 sg13g2_o21ai_1 _25261_ (.B1(_07188_),
    .Y(_02435_),
    .A1(net5274),
    .A2(_07190_));
 sg13g2_nand3_1 _25262_ (.B(_08246_),
    .C(_08446_),
    .A(net5204),
    .Y(_07191_));
 sg13g2_nand2_1 _25263_ (.Y(_07192_),
    .A(net5270),
    .B(_07191_));
 sg13g2_o21ai_1 _25264_ (.B1(_07192_),
    .Y(_07193_),
    .A1(net7103),
    .A2(net5270));
 sg13g2_inv_1 _25265_ (.Y(_02436_),
    .A(_07193_));
 sg13g2_nand2_1 _25266_ (.Y(_07194_),
    .A(net5203),
    .B(_08199_));
 sg13g2_nor3_1 _25267_ (.A(_08215_),
    .B(_07174_),
    .C(_07194_),
    .Y(_07195_));
 sg13g2_nor2_2 _25268_ (.A(_08183_),
    .B(_07174_),
    .Y(_07196_));
 sg13g2_a21oi_1 _25269_ (.A1(_08242_),
    .A2(_07196_),
    .Y(_07197_),
    .B1(_07195_));
 sg13g2_nand3_1 _25270_ (.B(net5201),
    .C(_07173_),
    .A(net5275),
    .Y(_07198_));
 sg13g2_nand3_1 _25271_ (.B(_07197_),
    .C(_07198_),
    .A(net5270),
    .Y(_07199_));
 sg13g2_o21ai_1 _25272_ (.B1(_07199_),
    .Y(_07200_),
    .A1(net7221),
    .A2(net5271));
 sg13g2_inv_1 _25273_ (.Y(_02437_),
    .A(_07200_));
 sg13g2_nor2_2 _25274_ (.A(net5271),
    .B(_08332_),
    .Y(_07201_));
 sg13g2_nand2_1 _25275_ (.Y(_07202_),
    .A(net7139),
    .B(_07201_));
 sg13g2_nand2_1 _25276_ (.Y(_07203_),
    .A(net6733),
    .B(net5204));
 sg13g2_nand3b_1 _25277_ (.B(_08248_),
    .C(net5201),
    .Y(_07204_),
    .A_N(_07201_));
 sg13g2_o21ai_1 _25278_ (.B1(_07202_),
    .Y(_02438_),
    .A1(_07203_),
    .A2(_07204_));
 sg13g2_o21ai_1 _25279_ (.B1(_07190_),
    .Y(_02439_),
    .A1(_08069_),
    .A2(net5271));
 sg13g2_nand2_1 _25280_ (.Y(_07205_),
    .A(net6996),
    .B(_07201_));
 sg13g2_nand2_1 _25281_ (.Y(_02440_),
    .A(_07204_),
    .B(_07205_));
 sg13g2_nor2_1 _25282_ (.A(net5349),
    .B(_08447_),
    .Y(_07206_));
 sg13g2_nand3_1 _25283_ (.B(_07173_),
    .C(_07206_),
    .A(_08175_),
    .Y(_07207_));
 sg13g2_a22oi_1 _25284_ (.Y(_07208_),
    .B1(_08218_),
    .B2(_07196_),
    .A2(net5347),
    .A1(net6973));
 sg13g2_nand2_1 _25285_ (.Y(_02441_),
    .A(_07207_),
    .B(_07208_));
 sg13g2_nor2_1 _25286_ (.A(net5347),
    .B(_07186_),
    .Y(_07209_));
 sg13g2_a21oi_1 _25287_ (.A1(_08056_),
    .A2(net5347),
    .Y(_02442_),
    .B1(_07209_));
 sg13g2_a22oi_1 _25288_ (.Y(_07210_),
    .B1(_07185_),
    .B2(_07206_),
    .A2(net5348),
    .A1(net4410));
 sg13g2_inv_1 _25289_ (.Y(_02443_),
    .A(_07210_));
 sg13g2_a21oi_1 _25290_ (.A1(_08194_),
    .A2(net5202),
    .Y(_07211_),
    .B1(net5200));
 sg13g2_nand2_2 _25291_ (.Y(_07212_),
    .A(net5275),
    .B(_07184_));
 sg13g2_inv_1 _25292_ (.Y(_07213_),
    .A(_07212_));
 sg13g2_nor3_1 _25293_ (.A(net5350),
    .B(_07211_),
    .C(_07212_),
    .Y(_07214_));
 sg13g2_a21o_1 _25294_ (.A2(net5350),
    .A1(net7225),
    .B1(_07214_),
    .X(_02444_));
 sg13g2_nor2_1 _25295_ (.A(net5203),
    .B(_07185_),
    .Y(_07215_));
 sg13g2_nand4_1 _25296_ (.B(net5272),
    .C(net5200),
    .A(_08204_),
    .Y(_07216_),
    .D(_07194_));
 sg13g2_a22oi_1 _25297_ (.Y(_07217_),
    .B1(_07206_),
    .B2(_07215_),
    .A2(net5347),
    .A1(net6937));
 sg13g2_nand2_1 _25298_ (.Y(_02445_),
    .A(_07216_),
    .B(_07217_));
 sg13g2_nor2_2 _25299_ (.A(net7228),
    .B(net5982),
    .Y(_07218_));
 sg13g2_a21oi_1 _25300_ (.A1(net6039),
    .A2(net5271),
    .Y(_02446_),
    .B1(_07218_));
 sg13g2_and2_1 _25301_ (.A(net4746),
    .B(_03048_),
    .X(_07219_));
 sg13g2_nor2_1 _25302_ (.A(net3023),
    .B(net4645),
    .Y(_07220_));
 sg13g2_a21oi_1 _25303_ (.A1(net5262),
    .A2(net4645),
    .Y(_02447_),
    .B1(_07220_));
 sg13g2_nor2_1 _25304_ (.A(net3757),
    .B(net4645),
    .Y(_07221_));
 sg13g2_a21oi_1 _25305_ (.A1(net5236),
    .A2(net4645),
    .Y(_02448_),
    .B1(_07221_));
 sg13g2_nor2_1 _25306_ (.A(net3425),
    .B(net4644),
    .Y(_07222_));
 sg13g2_a21oi_1 _25307_ (.A1(net5133),
    .A2(net4644),
    .Y(_02449_),
    .B1(_07222_));
 sg13g2_nor2_1 _25308_ (.A(net3132),
    .B(net4644),
    .Y(_07223_));
 sg13g2_a21oi_1 _25309_ (.A1(net5105),
    .A2(net4644),
    .Y(_02450_),
    .B1(_07223_));
 sg13g2_nor2_1 _25310_ (.A(net3372),
    .B(_07219_),
    .Y(_07224_));
 sg13g2_a21oi_1 _25311_ (.A1(net5177),
    .A2(net4645),
    .Y(_02451_),
    .B1(_07224_));
 sg13g2_nor2_1 _25312_ (.A(net3488),
    .B(net4645),
    .Y(_07225_));
 sg13g2_a21oi_1 _25313_ (.A1(net5148),
    .A2(net4645),
    .Y(_02452_),
    .B1(_07225_));
 sg13g2_nor2_1 _25314_ (.A(net3947),
    .B(net4644),
    .Y(_07226_));
 sg13g2_a21oi_1 _25315_ (.A1(net5081),
    .A2(net4644),
    .Y(_02453_),
    .B1(_07226_));
 sg13g2_nor2_1 _25316_ (.A(net3047),
    .B(net4644),
    .Y(_07227_));
 sg13g2_a21oi_1 _25317_ (.A1(net5057),
    .A2(net4644),
    .Y(_02454_),
    .B1(_07227_));
 sg13g2_o21ai_1 _25318_ (.B1(_07186_),
    .Y(_07228_),
    .A1(_08184_),
    .A2(net5202));
 sg13g2_nor2_1 _25319_ (.A(_08193_),
    .B(_07228_),
    .Y(_07229_));
 sg13g2_nand4_1 _25320_ (.B(_08205_),
    .C(_08446_),
    .A(net5275),
    .Y(_07230_),
    .D(_07196_));
 sg13g2_nand2_1 _25321_ (.Y(_07231_),
    .A(net5272),
    .B(_07230_));
 sg13g2_o21ai_1 _25322_ (.B1(net5203),
    .Y(_07232_),
    .A1(net5205),
    .A2(_08190_));
 sg13g2_a21oi_1 _25323_ (.A1(_07212_),
    .A2(_07232_),
    .Y(_07233_),
    .B1(_08206_));
 sg13g2_nor2_1 _25324_ (.A(_08454_),
    .B(_07187_),
    .Y(_07234_));
 sg13g2_o21ai_1 _25325_ (.B1(net5200),
    .Y(_07235_),
    .A1(_08175_),
    .A2(net5205));
 sg13g2_o21ai_1 _25326_ (.B1(_07235_),
    .Y(_07236_),
    .A1(_08454_),
    .A2(_07187_));
 sg13g2_nor2_1 _25327_ (.A(net5349),
    .B(_07234_),
    .Y(_07237_));
 sg13g2_nor4_2 _25328_ (.A(_07229_),
    .B(_07231_),
    .C(_07233_),
    .Y(_07238_),
    .D(_07236_));
 sg13g2_a21oi_1 _25329_ (.A1(_08116_),
    .A2(net5346),
    .Y(_02455_),
    .B1(_07238_));
 sg13g2_and2_1 _25330_ (.A(net5576),
    .B(net5997),
    .X(_07239_));
 sg13g2_and3_1 _25331_ (.X(_07240_),
    .A(net5997),
    .B(net5380),
    .C(_04890_));
 sg13g2_a21o_1 _25332_ (.A2(_07239_),
    .A1(net5349),
    .B1(net5319),
    .X(_02456_));
 sg13g2_nor2_1 _25333_ (.A(net6971),
    .B(net5318),
    .Y(_07241_));
 sg13g2_a21oi_1 _25334_ (.A1(_08191_),
    .A2(net5318),
    .Y(_02457_),
    .B1(_07241_));
 sg13g2_nor2_1 _25335_ (.A(net7032),
    .B(net5318),
    .Y(_07242_));
 sg13g2_a21oi_1 _25336_ (.A1(_08187_),
    .A2(net5318),
    .Y(_02458_),
    .B1(_07242_));
 sg13g2_nor2_1 _25337_ (.A(net6917),
    .B(net5319),
    .Y(_07243_));
 sg13g2_a21oi_1 _25338_ (.A1(_08201_),
    .A2(net5319),
    .Y(_02459_),
    .B1(_07243_));
 sg13g2_nor2_1 _25339_ (.A(net6928),
    .B(net5319),
    .Y(_07244_));
 sg13g2_a21oi_1 _25340_ (.A1(_08196_),
    .A2(net5319),
    .Y(_02460_),
    .B1(_07244_));
 sg13g2_nor2_1 _25341_ (.A(net6975),
    .B(net5318),
    .Y(_07245_));
 sg13g2_a21oi_1 _25342_ (.A1(_08181_),
    .A2(net5318),
    .Y(_02461_),
    .B1(_07245_));
 sg13g2_mux2_1 _25343_ (.A0(net6404),
    .A1(net5351),
    .S(net5318),
    .X(_02462_));
 sg13g2_nor2_1 _25344_ (.A(net6634),
    .B(net5319),
    .Y(_07246_));
 sg13g2_a21oi_1 _25345_ (.A1(_08244_),
    .A2(net5319),
    .Y(_02463_),
    .B1(_07246_));
 sg13g2_mux2_1 _25346_ (.A0(net3071),
    .A1(\atari2600.cpu.DI[7] ),
    .S(net5318),
    .X(_02464_));
 sg13g2_nor2_2 _25347_ (.A(net5480),
    .B(net5445),
    .Y(_07247_));
 sg13g2_inv_1 _25348_ (.Y(_07248_),
    .A(_07247_));
 sg13g2_nor2_1 _25349_ (.A(\atari2600.cpu.cld ),
    .B(\atari2600.cpu.sed ),
    .Y(_07249_));
 sg13g2_a21oi_1 _25350_ (.A1(_05026_),
    .A2(_07249_),
    .Y(_07250_),
    .B1(_07247_));
 sg13g2_mux2_1 _25351_ (.A0(_00055_),
    .A1(\atari2600.cpu.ADD[3] ),
    .S(net5577),
    .X(_07251_));
 sg13g2_nor2_1 _25352_ (.A(net5445),
    .B(_07251_),
    .Y(_07252_));
 sg13g2_a21oi_1 _25353_ (.A1(_08196_),
    .A2(net5445),
    .Y(_07253_),
    .B1(_07252_));
 sg13g2_mux2_1 _25354_ (.A0(net6733),
    .A1(_07253_),
    .S(_07250_),
    .X(_07254_));
 sg13g2_and2_1 _25355_ (.A(_07218_),
    .B(_07254_),
    .X(_02465_));
 sg13g2_nor3_1 _25356_ (.A(\atari2600.cpu.sei ),
    .B(\atari2600.cpu.cli ),
    .C(_08279_),
    .Y(_07255_));
 sg13g2_a221oi_1 _25357_ (.B2(_07247_),
    .C1(_07255_),
    .B1(_08453_),
    .A1(net5973),
    .Y(_07256_),
    .A2(_00145_));
 sg13g2_nand2_1 _25358_ (.Y(_07257_),
    .A(\atari2600.cpu.ADD[2] ),
    .B(_08453_));
 sg13g2_a21oi_1 _25359_ (.A1(_00056_),
    .A2(_08452_),
    .Y(_07258_),
    .B1(_08335_));
 sg13g2_o21ai_1 _25360_ (.B1(_07256_),
    .Y(_07259_),
    .A1(\atari2600.cpu.DIMUX[2] ),
    .A2(_08336_));
 sg13g2_a21o_1 _25361_ (.A2(_07258_),
    .A1(_07257_),
    .B1(_07259_),
    .X(_07260_));
 sg13g2_nand2b_1 _25362_ (.Y(_07261_),
    .B(net4146),
    .A_N(_07256_));
 sg13g2_nand3_1 _25363_ (.B(_07260_),
    .C(net4147),
    .A(_08311_),
    .Y(_02466_));
 sg13g2_a21oi_1 _25364_ (.A1(\atari2600.cpu.bit_ins ),
    .A2(_08276_),
    .Y(_07262_),
    .B1(_07248_));
 sg13g2_nor2_1 _25365_ (.A(\atari2600.cpu.plp ),
    .B(\atari2600.cpu.clv ),
    .Y(_07263_));
 sg13g2_nor3_1 _25366_ (.A(net5577),
    .B(\atari2600.cpu.adc_sbc ),
    .C(\atari2600.cpu.clv ),
    .Y(_07264_));
 sg13g2_a21oi_1 _25367_ (.A1(net5480),
    .A2(_07264_),
    .Y(_07265_),
    .B1(_07262_));
 sg13g2_xor2_1 _25368_ (.B(\atari2600.cpu.ALU.AI7 ),
    .A(\atari2600.cpu.ALU.BI7 ),
    .X(_07266_));
 sg13g2_xor2_1 _25369_ (.B(_00104_),
    .A(\atari2600.cpu.ALU.CO ),
    .X(_07267_));
 sg13g2_xnor2_1 _25370_ (.Y(_07268_),
    .A(_07266_),
    .B(_07267_));
 sg13g2_a221oi_1 _25371_ (.B2(_07268_),
    .C1(_08212_),
    .B1(_07263_),
    .A1(net5568),
    .Y(_07269_),
    .A2(\atari2600.cpu.plp ));
 sg13g2_a21oi_1 _25372_ (.A1(_08212_),
    .A2(_08244_),
    .Y(_07270_),
    .B1(_07269_));
 sg13g2_mux2_1 _25373_ (.A0(net3684),
    .A1(_07270_),
    .S(_07265_),
    .X(_02467_));
 sg13g2_nand2_1 _25374_ (.Y(_07271_),
    .A(_08232_),
    .B(_07262_));
 sg13g2_nor3_1 _25375_ (.A(\atari2600.cpu.compare ),
    .B(net5577),
    .C(_08212_),
    .Y(_07272_));
 sg13g2_o21ai_1 _25376_ (.B1(_07272_),
    .Y(_07273_),
    .A1(_08116_),
    .A2(_08514_));
 sg13g2_nand2_1 _25377_ (.Y(_07274_),
    .A(_07271_),
    .B(_07273_));
 sg13g2_nor3_1 _25378_ (.A(net5273),
    .B(net5480),
    .C(net5479),
    .Y(_07275_));
 sg13g2_a21oi_1 _25379_ (.A1(_08212_),
    .A2(_08232_),
    .Y(_07276_),
    .B1(\atari2600.cpu.ADD[7] ));
 sg13g2_nor3_1 _25380_ (.A(_07274_),
    .B(_07275_),
    .C(_07276_),
    .Y(_07277_));
 sg13g2_a21o_1 _25381_ (.A2(_07274_),
    .A1(net4089),
    .B1(_07277_),
    .X(_02468_));
 sg13g2_nand2_1 _25382_ (.Y(_07278_),
    .A(_08232_),
    .B(_07247_));
 sg13g2_o21ai_1 _25383_ (.B1(_07278_),
    .Y(_07279_),
    .A1(\atari2600.cpu.bit_ins ),
    .A2(_07273_));
 sg13g2_nor4_1 _25384_ (.A(net5568),
    .B(\atari2600.cpu.ADD[7] ),
    .C(net5569),
    .D(net5570),
    .Y(_07280_));
 sg13g2_nor4_1 _25385_ (.A(net5571),
    .B(\atari2600.cpu.ADD[3] ),
    .C(\atari2600.cpu.ADD[1] ),
    .D(net5572),
    .Y(_07281_));
 sg13g2_nand2_1 _25386_ (.Y(_07282_),
    .A(_07280_),
    .B(_07281_));
 sg13g2_nand2b_1 _25387_ (.Y(_07283_),
    .B(_07282_),
    .A_N(net5577));
 sg13g2_a21oi_1 _25388_ (.A1(_08061_),
    .A2(\atari2600.cpu.plp ),
    .Y(_07284_),
    .B1(net5445));
 sg13g2_a22oi_1 _25389_ (.Y(_07285_),
    .B1(_07283_),
    .B2(_07284_),
    .A2(net5445),
    .A1(\atari2600.cpu.DIMUX[1] ));
 sg13g2_nand2_1 _25390_ (.Y(_07286_),
    .A(net5479),
    .B(_07282_));
 sg13g2_a21oi_1 _25391_ (.A1(_08232_),
    .A2(_07285_),
    .Y(_07287_),
    .B1(_07279_));
 sg13g2_a22oi_1 _25392_ (.Y(_07288_),
    .B1(_07286_),
    .B2(_07287_),
    .A2(_07279_),
    .A1(net3931));
 sg13g2_inv_1 _25393_ (.Y(_02469_),
    .A(net3932));
 sg13g2_a22oi_1 _25394_ (.Y(_07289_),
    .B1(net5479),
    .B2(net7146),
    .A2(net5480),
    .A1(net7280));
 sg13g2_nor3_1 _25395_ (.A(\atari2600.cpu.shift ),
    .B(\atari2600.cpu.compare ),
    .C(\atari2600.cpu.adc_sbc ),
    .Y(_07290_));
 sg13g2_nor3_1 _25396_ (.A(\atari2600.cpu.clc ),
    .B(net5577),
    .C(\atari2600.cpu.sec ),
    .Y(_07291_));
 sg13g2_a21oi_1 _25397_ (.A1(_07290_),
    .A2(_07291_),
    .Y(_07292_),
    .B1(_07289_));
 sg13g2_mux2_1 _25398_ (.A0(_00057_),
    .A1(net5572),
    .S(net5577),
    .X(_07293_));
 sg13g2_nand2_1 _25399_ (.Y(_07294_),
    .A(_07290_),
    .B(_07293_));
 sg13g2_o21ai_1 _25400_ (.B1(_07294_),
    .Y(_07295_),
    .A1(_08070_),
    .A2(_07290_));
 sg13g2_o21ai_1 _25401_ (.B1(_08336_),
    .Y(_07296_),
    .A1(_08068_),
    .A2(_07292_));
 sg13g2_a21oi_1 _25402_ (.A1(_07292_),
    .A2(_07295_),
    .Y(_07297_),
    .B1(_07296_));
 sg13g2_a21oi_1 _25403_ (.A1(_08191_),
    .A2(net5445),
    .Y(_02470_),
    .B1(net7281));
 sg13g2_nand2_2 _25404_ (.Y(_07298_),
    .A(net5423),
    .B(net5419));
 sg13g2_mux2_1 _25405_ (.A0(net5783),
    .A1(net4284),
    .S(_07298_),
    .X(_02471_));
 sg13g2_mux2_1 _25406_ (.A0(net5752),
    .A1(net4243),
    .S(_07298_),
    .X(_02472_));
 sg13g2_mux2_1 _25407_ (.A0(net5723),
    .A1(net6288),
    .S(_07298_),
    .X(_02473_));
 sg13g2_mux2_1 _25408_ (.A0(net5694),
    .A1(net6219),
    .S(_07298_),
    .X(_02474_));
 sg13g2_mux2_1 _25409_ (.A0(net5666),
    .A1(net6515),
    .S(_07298_),
    .X(_02475_));
 sg13g2_mux2_1 _25410_ (.A0(net5641),
    .A1(net6764),
    .S(_07298_),
    .X(_02476_));
 sg13g2_mux2_1 _25411_ (.A0(net5608),
    .A1(net6401),
    .S(_07298_),
    .X(_02477_));
 sg13g2_a21o_1 _25412_ (.A2(net5315),
    .A1(\atari2600.cpu.backwards ),
    .B1(_08177_),
    .X(_02478_));
 sg13g2_mux2_1 _25413_ (.A0(net4279),
    .A1(_08561_),
    .S(net5211),
    .X(_02479_));
 sg13g2_mux2_1 _25414_ (.A0(net7008),
    .A1(_08552_),
    .S(net5211),
    .X(_02480_));
 sg13g2_mux2_1 _25415_ (.A0(net4291),
    .A1(_08574_),
    .S(net5210),
    .X(_02481_));
 sg13g2_mux2_1 _25416_ (.A0(net3430),
    .A1(_08541_),
    .S(net5210),
    .X(_02482_));
 sg13g2_mux2_1 _25417_ (.A0(net3487),
    .A1(_08626_),
    .S(net5210),
    .X(_02483_));
 sg13g2_mux2_1 _25418_ (.A0(net3908),
    .A1(_08614_),
    .S(net5210),
    .X(_02484_));
 sg13g2_mux2_1 _25419_ (.A0(net3371),
    .A1(_08724_),
    .S(net5210),
    .X(_02485_));
 sg13g2_mux2_1 _25420_ (.A0(net4126),
    .A1(_08604_),
    .S(net5210),
    .X(_02486_));
 sg13g2_nor2_1 _25421_ (.A(net6091),
    .B(net5363),
    .Y(_07299_));
 sg13g2_a21oi_1 _25422_ (.A1(net5363),
    .A2(_05157_),
    .Y(_02487_),
    .B1(_07299_));
 sg13g2_a21oi_1 _25423_ (.A1(_08585_),
    .A2(_05129_),
    .Y(_07300_),
    .B1(net5358));
 sg13g2_nand2b_1 _25424_ (.Y(_07301_),
    .B(_05142_),
    .A_N(net5355));
 sg13g2_nor2_1 _25425_ (.A(_07300_),
    .B(_07301_),
    .Y(_07302_));
 sg13g2_nand2b_1 _25426_ (.Y(_07303_),
    .B(_05154_),
    .A_N(_08546_));
 sg13g2_a22oi_1 _25427_ (.Y(_07304_),
    .B1(net5361),
    .B2(\atari2600.cpu.ADD[1] ),
    .A2(net5441),
    .A1(\atari2600.cpu.ABH[1] ));
 sg13g2_nand2_1 _25428_ (.Y(_07305_),
    .A(_07303_),
    .B(_07304_));
 sg13g2_a21oi_2 _25429_ (.B1(_07305_),
    .Y(_07306_),
    .A2(net5402),
    .A1(\atari2600.cpu.DIMUX[1] ));
 sg13g2_nor2b_1 _25430_ (.A(_07306_),
    .B_N(net5355),
    .Y(_07307_));
 sg13g2_nand2_1 _25431_ (.Y(_07308_),
    .A(\atari2600.cpu.PC[0] ),
    .B(net5438));
 sg13g2_o21ai_1 _25432_ (.B1(_07308_),
    .Y(_07309_),
    .A1(_08191_),
    .A2(_05125_));
 sg13g2_nand2_1 _25433_ (.Y(_07310_),
    .A(_05145_),
    .B(_07309_));
 sg13g2_nand2_1 _25434_ (.Y(_07311_),
    .A(_05149_),
    .B(_07310_));
 sg13g2_a22oi_1 _25435_ (.Y(_07312_),
    .B1(net5361),
    .B2(net5572),
    .A2(net5444),
    .A1(\atari2600.cpu.ABH[0] ));
 sg13g2_inv_1 _25436_ (.Y(_07313_),
    .A(_07312_));
 sg13g2_a221oi_1 _25437_ (.B2(_08555_),
    .C1(_07313_),
    .B1(_05154_),
    .A1(\atari2600.cpu.DIMUX[0] ),
    .Y(_07314_),
    .A2(net5402));
 sg13g2_o21ai_1 _25438_ (.B1(_07309_),
    .Y(_07315_),
    .A1(_05147_),
    .A2(_07314_));
 sg13g2_a221oi_1 _25439_ (.B2(_07311_),
    .C1(net5355),
    .B1(_07315_),
    .A1(_07310_),
    .Y(_07316_),
    .A2(_07314_));
 sg13g2_nor2_1 _25440_ (.A(_07307_),
    .B(_07316_),
    .Y(_07317_));
 sg13g2_o21ai_1 _25441_ (.B1(net5358),
    .Y(_07318_),
    .A1(net5323),
    .A2(_07309_));
 sg13g2_a21o_1 _25442_ (.A2(_07309_),
    .A1(net5323),
    .B1(_07318_),
    .X(_07319_));
 sg13g2_a21o_1 _25443_ (.A2(_07319_),
    .A1(_05163_),
    .B1(_07317_),
    .X(_07320_));
 sg13g2_inv_1 _25444_ (.Y(_07321_),
    .A(_07320_));
 sg13g2_nand2_1 _25445_ (.Y(_07322_),
    .A(_07317_),
    .B(_07319_));
 sg13g2_and3_1 _25446_ (.X(_07323_),
    .A(_07302_),
    .B(_07320_),
    .C(_07322_));
 sg13g2_a21oi_1 _25447_ (.A1(_07320_),
    .A2(_07322_),
    .Y(_07324_),
    .B1(_07302_));
 sg13g2_nor3_1 _25448_ (.A(net5313),
    .B(_07323_),
    .C(_07324_),
    .Y(_07325_));
 sg13g2_a21o_1 _25449_ (.A2(net5313),
    .A1(net5572),
    .B1(_07325_),
    .X(_02488_));
 sg13g2_nor2_1 _25450_ (.A(net7308),
    .B(net5364),
    .Y(_07326_));
 sg13g2_nor2_1 _25451_ (.A(_07321_),
    .B(_07323_),
    .Y(_07327_));
 sg13g2_a22oi_1 _25452_ (.Y(_07328_),
    .B1(net5361),
    .B2(net5571),
    .A2(net5441),
    .A1(\atari2600.cpu.ABH[2] ));
 sg13g2_a22oi_1 _25453_ (.Y(_07329_),
    .B1(_05154_),
    .B2(_08568_),
    .A2(_04881_),
    .A1(\atari2600.cpu.DIMUX[2] ));
 sg13g2_nand2_1 _25454_ (.Y(_07330_),
    .A(_07328_),
    .B(_07329_));
 sg13g2_nand2_1 _25455_ (.Y(_07331_),
    .A(\atari2600.cpu.PC[1] ),
    .B(net5438));
 sg13g2_o21ai_1 _25456_ (.B1(_07331_),
    .Y(_07332_),
    .A1(_08187_),
    .A2(_05125_));
 sg13g2_nand2_1 _25457_ (.Y(_07333_),
    .A(_05145_),
    .B(_07332_));
 sg13g2_nand2_1 _25458_ (.Y(_07334_),
    .A(_05149_),
    .B(_07333_));
 sg13g2_o21ai_1 _25459_ (.B1(_07332_),
    .Y(_07335_),
    .A1(_05147_),
    .A2(_07306_));
 sg13g2_a221oi_1 _25460_ (.B2(_07335_),
    .C1(net5355),
    .B1(_07334_),
    .A1(_07306_),
    .Y(_07336_),
    .A2(_07333_));
 sg13g2_a21oi_1 _25461_ (.A1(net5357),
    .A2(_07330_),
    .Y(_07337_),
    .B1(_07336_));
 sg13g2_o21ai_1 _25462_ (.B1(net5358),
    .Y(_07338_),
    .A1(net5323),
    .A2(_07332_));
 sg13g2_a21o_1 _25463_ (.A2(_07332_),
    .A1(net5323),
    .B1(_07338_),
    .X(_07339_));
 sg13g2_a21oi_1 _25464_ (.A1(_05163_),
    .A2(_07339_),
    .Y(_07340_),
    .B1(_07337_));
 sg13g2_a21o_1 _25465_ (.A2(_07339_),
    .A1(_07337_),
    .B1(_07340_),
    .X(_07341_));
 sg13g2_nor2_1 _25466_ (.A(_07327_),
    .B(_07341_),
    .Y(_07342_));
 sg13g2_xnor2_1 _25467_ (.Y(_07343_),
    .A(_07327_),
    .B(_07341_));
 sg13g2_a21oi_1 _25468_ (.A1(net5364),
    .A2(_07343_),
    .Y(_02489_),
    .B1(_07326_));
 sg13g2_nor2_1 _25469_ (.A(net5571),
    .B(net5364),
    .Y(_07344_));
 sg13g2_a22oi_1 _25470_ (.Y(_07345_),
    .B1(net5361),
    .B2(\atari2600.cpu.ADD[3] ),
    .A2(net5442),
    .A1(\atari2600.cpu.ABH[3] ));
 sg13g2_a22oi_1 _25471_ (.Y(_07346_),
    .B1(_05154_),
    .B2(_08517_),
    .A2(net5402),
    .A1(\atari2600.cpu.DIMUX[3] ));
 sg13g2_nand2_2 _25472_ (.Y(_07347_),
    .A(_07345_),
    .B(_07346_));
 sg13g2_a22oi_1 _25473_ (.Y(_07348_),
    .B1(_05124_),
    .B2(\atari2600.cpu.DIMUX[2] ),
    .A2(net5438),
    .A1(_08058_));
 sg13g2_nand2b_1 _25474_ (.Y(_07349_),
    .B(_05145_),
    .A_N(_07348_));
 sg13g2_a21oi_1 _25475_ (.A1(_05148_),
    .A2(_07330_),
    .Y(_07350_),
    .B1(_07348_));
 sg13g2_a21oi_1 _25476_ (.A1(_05149_),
    .A2(_07349_),
    .Y(_07351_),
    .B1(_07350_));
 sg13g2_nor2b_1 _25477_ (.A(_07330_),
    .B_N(_07349_),
    .Y(_07352_));
 sg13g2_nor3_1 _25478_ (.A(net5356),
    .B(_07351_),
    .C(_07352_),
    .Y(_07353_));
 sg13g2_a21oi_1 _25479_ (.A1(net5356),
    .A2(_07347_),
    .Y(_07354_),
    .B1(_07353_));
 sg13g2_xnor2_1 _25480_ (.Y(_07355_),
    .A(net5323),
    .B(_07348_));
 sg13g2_nand2_1 _25481_ (.Y(_07356_),
    .A(net5359),
    .B(_07355_));
 sg13g2_a21o_1 _25482_ (.A2(_07356_),
    .A1(_05163_),
    .B1(_07354_),
    .X(_07357_));
 sg13g2_nand2_1 _25483_ (.Y(_07358_),
    .A(_07354_),
    .B(_07356_));
 sg13g2_nand2_1 _25484_ (.Y(_07359_),
    .A(_07357_),
    .B(_07358_));
 sg13g2_nor2_1 _25485_ (.A(_07340_),
    .B(_07342_),
    .Y(_07360_));
 sg13g2_xnor2_1 _25486_ (.Y(_07361_),
    .A(_07359_),
    .B(_07360_));
 sg13g2_a21oi_1 _25487_ (.A1(net5364),
    .A2(_07361_),
    .Y(_02490_),
    .B1(_07344_));
 sg13g2_nor2_1 _25488_ (.A(net7349),
    .B(net5367),
    .Y(_07362_));
 sg13g2_a22oi_1 _25489_ (.Y(_07363_),
    .B1(_08522_),
    .B2(net5570),
    .A2(net5441),
    .A1(\atari2600.cpu.ABH[4] ));
 sg13g2_a22oi_1 _25490_ (.Y(_07364_),
    .B1(_05154_),
    .B2(_08620_),
    .A2(net5402),
    .A1(\atari2600.cpu.DIMUX[4] ));
 sg13g2_and2_1 _25491_ (.A(_07363_),
    .B(_07364_),
    .X(_07365_));
 sg13g2_inv_1 _25492_ (.Y(_07366_),
    .A(_07365_));
 sg13g2_nand2_1 _25493_ (.Y(_07367_),
    .A(\atari2600.cpu.PC[3] ),
    .B(net5438));
 sg13g2_o21ai_1 _25494_ (.B1(_07367_),
    .Y(_07368_),
    .A1(_08196_),
    .A2(_05125_));
 sg13g2_nand2_1 _25495_ (.Y(_07369_),
    .A(_05145_),
    .B(_07368_));
 sg13g2_nand2_1 _25496_ (.Y(_07370_),
    .A(_05148_),
    .B(_07347_));
 sg13g2_a22oi_1 _25497_ (.Y(_07371_),
    .B1(_07370_),
    .B2(_07368_),
    .A2(_07369_),
    .A1(_05149_));
 sg13g2_nor2b_1 _25498_ (.A(_07347_),
    .B_N(_07369_),
    .Y(_07372_));
 sg13g2_nor3_1 _25499_ (.A(net5356),
    .B(_07371_),
    .C(_07372_),
    .Y(_07373_));
 sg13g2_a21oi_1 _25500_ (.A1(net5357),
    .A2(_07366_),
    .Y(_07374_),
    .B1(_07373_));
 sg13g2_o21ai_1 _25501_ (.B1(net5359),
    .Y(_07375_),
    .A1(net5324),
    .A2(_07368_));
 sg13g2_a21oi_1 _25502_ (.A1(net5324),
    .A2(_07368_),
    .Y(_07376_),
    .B1(_07375_));
 sg13g2_inv_1 _25503_ (.Y(_07377_),
    .A(_07376_));
 sg13g2_a21o_1 _25504_ (.A2(_07377_),
    .A1(_05163_),
    .B1(_07374_),
    .X(_07378_));
 sg13g2_nand2_1 _25505_ (.Y(_07379_),
    .A(_07374_),
    .B(_07377_));
 sg13g2_nand2_1 _25506_ (.Y(_07380_),
    .A(_07378_),
    .B(_07379_));
 sg13g2_o21ai_1 _25507_ (.B1(_07357_),
    .Y(_07381_),
    .A1(_07359_),
    .A2(_07360_));
 sg13g2_nand2b_1 _25508_ (.Y(_07382_),
    .B(_07381_),
    .A_N(_07380_));
 sg13g2_xor2_1 _25509_ (.B(_07381_),
    .A(_07380_),
    .X(_07383_));
 sg13g2_a21oi_1 _25510_ (.A1(net5367),
    .A2(_07383_),
    .Y(_02491_),
    .B1(_07362_));
 sg13g2_nand2_1 _25511_ (.Y(_07384_),
    .A(net5570),
    .B(net5313));
 sg13g2_a22oi_1 _25512_ (.Y(_07385_),
    .B1(net5361),
    .B2(net5569),
    .A2(net5443),
    .A1(\atari2600.cpu.ABH[5] ));
 sg13g2_a22oi_1 _25513_ (.Y(_07386_),
    .B1(_05154_),
    .B2(_08609_),
    .A2(net5402),
    .A1(net5351));
 sg13g2_nand2_1 _25514_ (.Y(_07387_),
    .A(_07385_),
    .B(_07386_));
 sg13g2_nand2_1 _25515_ (.Y(_07388_),
    .A(\atari2600.cpu.PC[4] ),
    .B(net5437));
 sg13g2_o21ai_1 _25516_ (.B1(_07388_),
    .Y(_07389_),
    .A1(_08181_),
    .A2(_05125_));
 sg13g2_nand2_1 _25517_ (.Y(_07390_),
    .A(_05145_),
    .B(_07389_));
 sg13g2_nand2_1 _25518_ (.Y(_07391_),
    .A(_05149_),
    .B(_07390_));
 sg13g2_o21ai_1 _25519_ (.B1(_07389_),
    .Y(_07392_),
    .A1(_05147_),
    .A2(_07365_));
 sg13g2_a221oi_1 _25520_ (.B2(_07392_),
    .C1(net5357),
    .B1(_07391_),
    .A1(_07365_),
    .Y(_07393_),
    .A2(_07390_));
 sg13g2_a21oi_1 _25521_ (.A1(net5356),
    .A2(_07387_),
    .Y(_07394_),
    .B1(_07393_));
 sg13g2_o21ai_1 _25522_ (.B1(net5359),
    .Y(_07395_),
    .A1(net5324),
    .A2(_07389_));
 sg13g2_a21oi_1 _25523_ (.A1(net5324),
    .A2(_07389_),
    .Y(_07396_),
    .B1(_07395_));
 sg13g2_nor2_1 _25524_ (.A(_05162_),
    .B(_07396_),
    .Y(_07397_));
 sg13g2_mux2_1 _25525_ (.A0(_07397_),
    .A1(_07396_),
    .S(_07394_),
    .X(_07398_));
 sg13g2_nand2_1 _25526_ (.Y(_07399_),
    .A(\atari2600.cpu.adc_bcd ),
    .B(_08276_));
 sg13g2_a21oi_1 _25527_ (.A1(_07343_),
    .A2(_07361_),
    .Y(_07400_),
    .B1(_07399_));
 sg13g2_nand2b_1 _25528_ (.Y(_07401_),
    .B(_07400_),
    .A_N(_07383_));
 sg13g2_and3_2 _25529_ (.X(_07402_),
    .A(_07378_),
    .B(_07382_),
    .C(_07401_));
 sg13g2_nand2b_1 _25530_ (.Y(_07403_),
    .B(_07398_),
    .A_N(_07402_));
 sg13g2_xor2_1 _25531_ (.B(_07402_),
    .A(_07398_),
    .X(_07404_));
 sg13g2_o21ai_1 _25532_ (.B1(_07384_),
    .Y(_02492_),
    .A1(net5313),
    .A2(_07404_));
 sg13g2_nor2_1 _25533_ (.A(net5569),
    .B(net5364),
    .Y(_07405_));
 sg13g2_o21ai_1 _25534_ (.B1(_07403_),
    .Y(_07406_),
    .A1(_07394_),
    .A2(_07397_));
 sg13g2_a22oi_1 _25535_ (.Y(_07407_),
    .B1(net5361),
    .B2(net5568),
    .A2(net5443),
    .A1(\atari2600.cpu.ABH[6] ));
 sg13g2_a22oi_1 _25536_ (.Y(_07408_),
    .B1(_05154_),
    .B2(_08718_),
    .A2(net5402),
    .A1(\atari2600.cpu.DIMUX[6] ));
 sg13g2_nand2_1 _25537_ (.Y(_07409_),
    .A(_07407_),
    .B(_07408_));
 sg13g2_a22oi_1 _25538_ (.Y(_07410_),
    .B1(_05124_),
    .B2(net5351),
    .A2(net5437),
    .A1(\atari2600.cpu.PC[5] ));
 sg13g2_nand2b_1 _25539_ (.Y(_07411_),
    .B(_05145_),
    .A_N(_07410_));
 sg13g2_a21oi_1 _25540_ (.A1(_05148_),
    .A2(_07387_),
    .Y(_07412_),
    .B1(_07410_));
 sg13g2_a21oi_1 _25541_ (.A1(_05149_),
    .A2(_07411_),
    .Y(_07413_),
    .B1(_07412_));
 sg13g2_nor2b_1 _25542_ (.A(_07387_),
    .B_N(_07411_),
    .Y(_07414_));
 sg13g2_nor3_1 _25543_ (.A(net5356),
    .B(_07413_),
    .C(_07414_),
    .Y(_07415_));
 sg13g2_a21oi_1 _25544_ (.A1(net5356),
    .A2(_07409_),
    .Y(_07416_),
    .B1(_07415_));
 sg13g2_xnor2_1 _25545_ (.Y(_07417_),
    .A(net5324),
    .B(_07410_));
 sg13g2_and2_1 _25546_ (.A(net5358),
    .B(_07417_),
    .X(_07418_));
 sg13g2_nor2_1 _25547_ (.A(_05162_),
    .B(_07418_),
    .Y(_07419_));
 sg13g2_or2_1 _25548_ (.X(_07420_),
    .B(_07419_),
    .A(_07416_));
 sg13g2_mux2_1 _25549_ (.A0(_07419_),
    .A1(_07418_),
    .S(_07416_),
    .X(_07421_));
 sg13g2_nand2_1 _25550_ (.Y(_07422_),
    .A(_07406_),
    .B(_07421_));
 sg13g2_xnor2_1 _25551_ (.Y(_07423_),
    .A(_07406_),
    .B(_07421_));
 sg13g2_a21oi_1 _25552_ (.A1(net5364),
    .A2(_07423_),
    .Y(_02493_),
    .B1(_07405_));
 sg13g2_nor2_1 _25553_ (.A(net5568),
    .B(net5364),
    .Y(_07424_));
 sg13g2_nand2_1 _25554_ (.Y(_07425_),
    .A(\atari2600.cpu.PC[6] ),
    .B(net5437));
 sg13g2_o21ai_1 _25555_ (.B1(_07425_),
    .Y(_07426_),
    .A1(_08244_),
    .A2(_05125_));
 sg13g2_nand2_1 _25556_ (.Y(_07427_),
    .A(_05145_),
    .B(_07426_));
 sg13g2_nand2_1 _25557_ (.Y(_07428_),
    .A(_05148_),
    .B(_07409_));
 sg13g2_a22oi_1 _25558_ (.Y(_07429_),
    .B1(_07428_),
    .B2(_07426_),
    .A2(_07427_),
    .A1(_05149_));
 sg13g2_nor2b_1 _25559_ (.A(_07409_),
    .B_N(_07427_),
    .Y(_07430_));
 sg13g2_nor3_1 _25560_ (.A(net5356),
    .B(_07429_),
    .C(_07430_),
    .Y(_07431_));
 sg13g2_a21oi_1 _25561_ (.A1(net5356),
    .A2(_05158_),
    .Y(_07432_),
    .B1(_07431_));
 sg13g2_o21ai_1 _25562_ (.B1(net5359),
    .Y(_07433_),
    .A1(net5324),
    .A2(_07426_));
 sg13g2_a21o_1 _25563_ (.A2(_07426_),
    .A1(net5324),
    .B1(_07433_),
    .X(_07434_));
 sg13g2_a21oi_1 _25564_ (.A1(_05163_),
    .A2(_07434_),
    .Y(_07435_),
    .B1(_07432_));
 sg13g2_a21o_1 _25565_ (.A2(_07434_),
    .A1(_07432_),
    .B1(_07435_),
    .X(_07436_));
 sg13g2_a21oi_1 _25566_ (.A1(_07420_),
    .A2(_07422_),
    .Y(_07437_),
    .B1(_07436_));
 sg13g2_nand3_1 _25567_ (.B(_07422_),
    .C(_07436_),
    .A(_07420_),
    .Y(_07438_));
 sg13g2_nand2b_1 _25568_ (.Y(_07439_),
    .B(_07438_),
    .A_N(_07437_));
 sg13g2_a21oi_1 _25569_ (.A1(net5367),
    .A2(_07439_),
    .Y(_02494_),
    .B1(_07424_));
 sg13g2_nand2_1 _25570_ (.Y(_07440_),
    .A(net7279),
    .B(net5313));
 sg13g2_o21ai_1 _25571_ (.B1(_05164_),
    .Y(_07441_),
    .A1(_05143_),
    .A2(_05160_));
 sg13g2_nand2b_1 _25572_ (.Y(_07442_),
    .B(_07441_),
    .A_N(_05161_));
 sg13g2_or2_1 _25573_ (.X(_07443_),
    .B(_07437_),
    .A(_07435_));
 sg13g2_inv_1 _25574_ (.Y(_07444_),
    .A(_07443_));
 sg13g2_xor2_1 _25575_ (.B(_07443_),
    .A(_07442_),
    .X(_07445_));
 sg13g2_o21ai_1 _25576_ (.B1(_07440_),
    .Y(_02495_),
    .A1(net5313),
    .A2(_07445_));
 sg13g2_nor2_1 _25577_ (.A(net7042),
    .B(net5362),
    .Y(_07446_));
 sg13g2_a21oi_1 _25578_ (.A1(net5362),
    .A2(_07402_),
    .Y(_02496_),
    .B1(_07446_));
 sg13g2_nor2b_1 _25579_ (.A(_07314_),
    .B_N(net5355),
    .Y(_07447_));
 sg13g2_o21ai_1 _25580_ (.B1(_07441_),
    .Y(_07448_),
    .A1(_05161_),
    .A2(_07444_));
 sg13g2_xnor2_1 _25581_ (.Y(_07449_),
    .A(_07447_),
    .B(_07448_));
 sg13g2_a21oi_1 _25582_ (.A1(_07423_),
    .A2(_07439_),
    .Y(_07450_),
    .B1(_07399_));
 sg13g2_nand2b_1 _25583_ (.Y(_07451_),
    .B(_07450_),
    .A_N(_07445_));
 sg13g2_and2_1 _25584_ (.A(net5364),
    .B(_07451_),
    .X(_07452_));
 sg13g2_a22oi_1 _25585_ (.Y(_02497_),
    .B1(_07449_),
    .B2(_07452_),
    .A2(net5312),
    .A1(_08070_));
 sg13g2_nor2_1 _25586_ (.A(net7123),
    .B(net5363),
    .Y(_07453_));
 sg13g2_nor3_1 _25587_ (.A(net5437),
    .B(_08391_),
    .C(_08440_),
    .Y(_07454_));
 sg13g2_nor2_1 _25588_ (.A(_08211_),
    .B(_08270_),
    .Y(_07455_));
 sg13g2_nand3_1 _25589_ (.B(_07454_),
    .C(_07455_),
    .A(_08482_),
    .Y(_07456_));
 sg13g2_nand3_1 _25590_ (.B(_08414_),
    .C(_08524_),
    .A(_08311_),
    .Y(_07457_));
 sg13g2_nor2_1 _25591_ (.A(_07456_),
    .B(_07457_),
    .Y(_07458_));
 sg13g2_nand3_1 _25592_ (.B(net5440),
    .C(_08524_),
    .A(_08288_),
    .Y(_07459_));
 sg13g2_nand2b_2 _25593_ (.Y(_07460_),
    .B(net5475),
    .A_N(_07459_));
 sg13g2_nor2_1 _25594_ (.A(_08413_),
    .B(_07460_),
    .Y(_07461_));
 sg13g2_nor3_1 _25595_ (.A(_00065_),
    .B(net5435),
    .C(_07460_),
    .Y(_07462_));
 sg13g2_a221oi_1 _25596_ (.B2(net5572),
    .C1(_07462_),
    .B1(_07459_),
    .A1(\atari2600.cpu.PC[0] ),
    .Y(_07463_),
    .A2(net5435));
 sg13g2_nor2_1 _25597_ (.A(_07458_),
    .B(_07463_),
    .Y(_07464_));
 sg13g2_xnor2_1 _25598_ (.Y(_07465_),
    .A(_07458_),
    .B(_07463_));
 sg13g2_a21oi_1 _25599_ (.A1(net5363),
    .A2(_07465_),
    .Y(_02498_),
    .B1(_07453_));
 sg13g2_nor2_1 _25600_ (.A(net7055),
    .B(net5365),
    .Y(_07466_));
 sg13g2_nor2_1 _25601_ (.A(_00064_),
    .B(_07460_),
    .Y(_07467_));
 sg13g2_a21oi_1 _25602_ (.A1(_08288_),
    .A2(_08524_),
    .Y(_07468_),
    .B1(_08061_));
 sg13g2_nor2_1 _25603_ (.A(\atari2600.cpu.res ),
    .B(net5475),
    .Y(_07469_));
 sg13g2_nor4_2 _25604_ (.A(_08548_),
    .B(_07467_),
    .C(_07468_),
    .Y(_07470_),
    .D(_07469_));
 sg13g2_nand2b_1 _25605_ (.Y(_07471_),
    .B(_07464_),
    .A_N(_07470_));
 sg13g2_xor2_1 _25606_ (.B(_07470_),
    .A(_07464_),
    .X(_07472_));
 sg13g2_a21oi_1 _25607_ (.A1(net5365),
    .A2(_07472_),
    .Y(_02499_),
    .B1(_07466_));
 sg13g2_o21ai_1 _25608_ (.B1(net5475),
    .Y(_07473_),
    .A1(_00099_),
    .A2(net5439));
 sg13g2_a21oi_1 _25609_ (.A1(net5571),
    .A2(net5387),
    .Y(_07474_),
    .B1(_07473_));
 sg13g2_o21ai_1 _25610_ (.B1(_07474_),
    .Y(_07475_),
    .A1(_00082_),
    .A2(_07459_));
 sg13g2_nor2b_1 _25611_ (.A(_07475_),
    .B_N(_07471_),
    .Y(_07476_));
 sg13g2_nor2b_2 _25612_ (.A(_07471_),
    .B_N(_07475_),
    .Y(_07477_));
 sg13g2_nor3_1 _25613_ (.A(net5314),
    .B(_07476_),
    .C(_07477_),
    .Y(_07478_));
 sg13g2_a21o_1 _25614_ (.A2(net5314),
    .A1(net6980),
    .B1(_07478_),
    .X(_02500_));
 sg13g2_o21ai_1 _25615_ (.B1(_08314_),
    .Y(_07479_),
    .A1(_00101_),
    .A2(net5439));
 sg13g2_a21oi_1 _25616_ (.A1(\atari2600.cpu.ADD[3] ),
    .A2(net5388),
    .Y(_07480_),
    .B1(_07479_));
 sg13g2_o21ai_1 _25617_ (.B1(_07480_),
    .Y(_07481_),
    .A1(_00066_),
    .A2(_07459_));
 sg13g2_nand2_2 _25618_ (.Y(_07482_),
    .A(_07477_),
    .B(_07481_));
 sg13g2_o21ai_1 _25619_ (.B1(net5365),
    .Y(_07483_),
    .A1(_07477_),
    .A2(_07481_));
 sg13g2_nor2b_1 _25620_ (.A(_07483_),
    .B_N(_07482_),
    .Y(_07484_));
 sg13g2_a21o_1 _25621_ (.A2(net5314),
    .A1(net7155),
    .B1(_07484_),
    .X(_02501_));
 sg13g2_nor2_1 _25622_ (.A(net7189),
    .B(net5382),
    .Y(_07485_));
 sg13g2_o21ai_1 _25623_ (.B1(net5475),
    .Y(_07486_),
    .A1(_00067_),
    .A2(_07459_));
 sg13g2_a21oi_2 _25624_ (.B1(_07486_),
    .Y(_07487_),
    .A2(_07459_),
    .A1(net5570));
 sg13g2_xnor2_1 _25625_ (.Y(_07488_),
    .A(_07482_),
    .B(_07487_));
 sg13g2_a21oi_1 _25626_ (.A1(net5381),
    .A2(_07488_),
    .Y(_02502_),
    .B1(_07485_));
 sg13g2_nand2_1 _25627_ (.Y(_07489_),
    .A(net5569),
    .B(net5387));
 sg13g2_o21ai_1 _25628_ (.B1(_07489_),
    .Y(_07490_),
    .A1(_00068_),
    .A2(_07460_));
 sg13g2_nor3_1 _25629_ (.A(_08313_),
    .B(_08610_),
    .C(_07490_),
    .Y(_07491_));
 sg13g2_o21ai_1 _25630_ (.B1(_07491_),
    .Y(_07492_),
    .A1(_07482_),
    .A2(_07487_));
 sg13g2_or3_1 _25631_ (.A(_07482_),
    .B(_07487_),
    .C(_07491_),
    .X(_07493_));
 sg13g2_a21oi_1 _25632_ (.A1(_07492_),
    .A2(_07493_),
    .Y(_07494_),
    .B1(net5314));
 sg13g2_a21oi_1 _25633_ (.A1(_08073_),
    .A2(net5314),
    .Y(_02503_),
    .B1(_07494_));
 sg13g2_nor2_1 _25634_ (.A(net7079),
    .B(net5365),
    .Y(_07495_));
 sg13g2_o21ai_1 _25635_ (.B1(_08314_),
    .Y(_07496_),
    .A1(_00103_),
    .A2(net5440));
 sg13g2_a21oi_1 _25636_ (.A1(net5568),
    .A2(net5387),
    .Y(_07497_),
    .B1(_07496_));
 sg13g2_o21ai_1 _25637_ (.B1(_07497_),
    .Y(_07498_),
    .A1(_00069_),
    .A2(_07459_));
 sg13g2_nor2b_1 _25638_ (.A(_07493_),
    .B_N(_07498_),
    .Y(_07499_));
 sg13g2_xor2_1 _25639_ (.B(_07498_),
    .A(_07493_),
    .X(_07500_));
 sg13g2_a21oi_1 _25640_ (.A1(net5365),
    .A2(_07500_),
    .Y(_02504_),
    .B1(_07495_));
 sg13g2_nor2_1 _25641_ (.A(net7068),
    .B(net5365),
    .Y(_07501_));
 sg13g2_a21oi_1 _25642_ (.A1(\atari2600.cpu.ADD[7] ),
    .A2(net5387),
    .Y(_07502_),
    .B1(_08313_));
 sg13g2_o21ai_1 _25643_ (.B1(_07502_),
    .Y(_07503_),
    .A1(_00070_),
    .A2(_07460_));
 sg13g2_nor2_1 _25644_ (.A(_08600_),
    .B(_07503_),
    .Y(_07504_));
 sg13g2_nor2b_2 _25645_ (.A(_07504_),
    .B_N(_07499_),
    .Y(_07505_));
 sg13g2_xor2_1 _25646_ (.B(_07504_),
    .A(_07499_),
    .X(_07506_));
 sg13g2_a21oi_1 _25647_ (.A1(net5365),
    .A2(_07506_),
    .Y(_02505_),
    .B1(_07501_));
 sg13g2_nand2_1 _25648_ (.Y(_07507_),
    .A(\atari2600.cpu.DIMUX[0] ),
    .B(net5388));
 sg13g2_nor2_1 _25649_ (.A(_08313_),
    .B(net5317),
    .Y(_07508_));
 sg13g2_o21ai_1 _25650_ (.B1(net5475),
    .Y(_07509_),
    .A1(net5435),
    .A2(_07459_));
 sg13g2_a221oi_1 _25651_ (.B2(net5572),
    .C1(_07509_),
    .B1(net5435),
    .A1(\atari2600.cpu.ABH[0] ),
    .Y(_07510_),
    .A2(net5441));
 sg13g2_a22oi_1 _25652_ (.Y(_07511_),
    .B1(_07507_),
    .B2(_07510_),
    .A2(_07461_),
    .A1(_00071_));
 sg13g2_nand2_1 _25653_ (.Y(_07512_),
    .A(_07505_),
    .B(_07511_));
 sg13g2_o21ai_1 _25654_ (.B1(net5381),
    .Y(_07513_),
    .A1(_07505_),
    .A2(_07511_));
 sg13g2_nor2b_1 _25655_ (.A(_07513_),
    .B_N(_07512_),
    .Y(_07514_));
 sg13g2_a21o_1 _25656_ (.A2(net5314),
    .A1(net7064),
    .B1(_07514_),
    .X(_02506_));
 sg13g2_nand2_1 _25657_ (.Y(_07515_),
    .A(net4058),
    .B(net5314));
 sg13g2_nand2_1 _25658_ (.Y(_07516_),
    .A(\atari2600.cpu.DIMUX[1] ),
    .B(net5388));
 sg13g2_a221oi_1 _25659_ (.B2(_08074_),
    .C1(_07509_),
    .B1(net5435),
    .A1(\atari2600.cpu.ABH[1] ),
    .Y(_07517_),
    .A2(net5441));
 sg13g2_a22oi_1 _25660_ (.Y(_07518_),
    .B1(_07516_),
    .B2(_07517_),
    .A2(net5317),
    .A1(_00072_));
 sg13g2_nor2b_1 _25661_ (.A(_07512_),
    .B_N(_07518_),
    .Y(_07519_));
 sg13g2_xor2_1 _25662_ (.B(_07518_),
    .A(_07512_),
    .X(_07520_));
 sg13g2_o21ai_1 _25663_ (.B1(_07515_),
    .Y(_02507_),
    .A1(net5313),
    .A2(_07520_));
 sg13g2_nor2_1 _25664_ (.A(net6999),
    .B(net5381),
    .Y(_07521_));
 sg13g2_or2_1 _25665_ (.X(_07522_),
    .B(_08414_),
    .A(_00099_));
 sg13g2_a221oi_1 _25666_ (.B2(\atari2600.cpu.DIMUX[2] ),
    .C1(_07509_),
    .B1(net5387),
    .A1(\atari2600.cpu.ABH[2] ),
    .Y(_07523_),
    .A2(net5441));
 sg13g2_a22oi_1 _25667_ (.Y(_07524_),
    .B1(_07522_),
    .B2(_07523_),
    .A2(net5317),
    .A1(_00073_));
 sg13g2_nand2_1 _25668_ (.Y(_07525_),
    .A(_07519_),
    .B(_07524_));
 sg13g2_xnor2_1 _25669_ (.Y(_07526_),
    .A(_07519_),
    .B(_07524_));
 sg13g2_a21oi_1 _25670_ (.A1(net5381),
    .A2(_07526_),
    .Y(_02508_),
    .B1(_07521_));
 sg13g2_nor2_1 _25671_ (.A(net7089),
    .B(net5381),
    .Y(_07527_));
 sg13g2_a21oi_1 _25672_ (.A1(\atari2600.cpu.ABH[3] ),
    .A2(net5442),
    .Y(_07528_),
    .B1(_07509_));
 sg13g2_o21ai_1 _25673_ (.B1(_07528_),
    .Y(_07529_),
    .A1(_00101_),
    .A2(_08414_));
 sg13g2_a21oi_1 _25674_ (.A1(\atari2600.cpu.DIMUX[3] ),
    .A2(net5388),
    .Y(_07530_),
    .B1(_07529_));
 sg13g2_a21oi_1 _25675_ (.A1(_00074_),
    .A2(net5317),
    .Y(_07531_),
    .B1(_07530_));
 sg13g2_nand3_1 _25676_ (.B(_07524_),
    .C(_07531_),
    .A(_07519_),
    .Y(_07532_));
 sg13g2_xor2_1 _25677_ (.B(_07531_),
    .A(_07525_),
    .X(_07533_));
 sg13g2_a21oi_1 _25678_ (.A1(net5381),
    .A2(_07533_),
    .Y(_02509_),
    .B1(_07527_));
 sg13g2_nor2_1 _25679_ (.A(net6919),
    .B(net5381),
    .Y(_07534_));
 sg13g2_nand2_1 _25680_ (.Y(_07535_),
    .A(\atari2600.cpu.DIMUX[4] ),
    .B(net5388));
 sg13g2_a221oi_1 _25681_ (.B2(net5570),
    .C1(_07509_),
    .B1(net5435),
    .A1(\atari2600.cpu.ABH[4] ),
    .Y(_07536_),
    .A2(net5442));
 sg13g2_a22oi_1 _25682_ (.Y(_07537_),
    .B1(_07535_),
    .B2(_07536_),
    .A2(net5317),
    .A1(_00075_));
 sg13g2_nor2b_2 _25683_ (.A(_07532_),
    .B_N(_07537_),
    .Y(_07538_));
 sg13g2_xor2_1 _25684_ (.B(_07537_),
    .A(_07532_),
    .X(_07539_));
 sg13g2_a21oi_1 _25685_ (.A1(net5381),
    .A2(_07539_),
    .Y(_02510_),
    .B1(_07534_));
 sg13g2_nand2_1 _25686_ (.Y(_07540_),
    .A(net5351),
    .B(net5387));
 sg13g2_a221oi_1 _25687_ (.B2(_08076_),
    .C1(_07509_),
    .B1(net5435),
    .A1(\atari2600.cpu.ABH[5] ),
    .Y(_07541_),
    .A2(net5443));
 sg13g2_a22oi_1 _25688_ (.Y(_07542_),
    .B1(_07540_),
    .B2(_07541_),
    .A2(net5317),
    .A1(_00076_));
 sg13g2_nand2_1 _25689_ (.Y(_07543_),
    .A(_07538_),
    .B(_07542_));
 sg13g2_o21ai_1 _25690_ (.B1(net5365),
    .Y(_07544_),
    .A1(_07538_),
    .A2(_07542_));
 sg13g2_nor2b_1 _25691_ (.A(_07544_),
    .B_N(_07543_),
    .Y(_07545_));
 sg13g2_a21o_1 _25692_ (.A2(net5313),
    .A1(net6581),
    .B1(_07545_),
    .X(_02511_));
 sg13g2_nor2_1 _25693_ (.A(net7052),
    .B(net5366),
    .Y(_07546_));
 sg13g2_a21oi_1 _25694_ (.A1(\atari2600.cpu.ABH[6] ),
    .A2(net5443),
    .Y(_07547_),
    .B1(_07509_));
 sg13g2_o21ai_1 _25695_ (.B1(_07547_),
    .Y(_07548_),
    .A1(_00103_),
    .A2(_08414_));
 sg13g2_a21oi_1 _25696_ (.A1(\atari2600.cpu.DIMUX[6] ),
    .A2(net5387),
    .Y(_07549_),
    .B1(_07548_));
 sg13g2_a21oi_1 _25697_ (.A1(_08121_),
    .A2(net5317),
    .Y(_07550_),
    .B1(_07549_));
 sg13g2_nor2b_1 _25698_ (.A(_07543_),
    .B_N(_07550_),
    .Y(_07551_));
 sg13g2_xor2_1 _25699_ (.B(_07550_),
    .A(_07543_),
    .X(_07552_));
 sg13g2_a21oi_1 _25700_ (.A1(net5366),
    .A2(_07552_),
    .Y(_02512_),
    .B1(_07546_));
 sg13g2_nor2_1 _25701_ (.A(net7083),
    .B(net5366),
    .Y(_07553_));
 sg13g2_o21ai_1 _25702_ (.B1(_07508_),
    .Y(_07554_),
    .A1(_00104_),
    .A2(_08414_));
 sg13g2_a221oi_1 _25703_ (.B2(net5273),
    .C1(_07554_),
    .B1(net5387),
    .A1(\atari2600.cpu.ABH[7] ),
    .Y(_07555_),
    .A2(net5443));
 sg13g2_a21oi_1 _25704_ (.A1(_08123_),
    .A2(net5317),
    .Y(_07556_),
    .B1(_07555_));
 sg13g2_xnor2_1 _25705_ (.Y(_07557_),
    .A(_07551_),
    .B(_07556_));
 sg13g2_a21oi_1 _25706_ (.A1(net5366),
    .A2(_07557_),
    .Y(_02513_),
    .B1(_07553_));
 sg13g2_nand2_2 _25707_ (.Y(_07558_),
    .A(net4748),
    .B(_03158_));
 sg13g2_mux2_1 _25708_ (.A0(net5251),
    .A1(net6055),
    .S(_07558_),
    .X(_02514_));
 sg13g2_mux2_1 _25709_ (.A0(net5223),
    .A1(net4464),
    .S(_07558_),
    .X(_02515_));
 sg13g2_mux2_1 _25710_ (.A0(net5119),
    .A1(net6214),
    .S(_07558_),
    .X(_02516_));
 sg13g2_mux2_1 _25711_ (.A0(net5093),
    .A1(net6741),
    .S(_07558_),
    .X(_02517_));
 sg13g2_mux2_1 _25712_ (.A0(net5189),
    .A1(net6308),
    .S(_07558_),
    .X(_02518_));
 sg13g2_mux2_1 _25713_ (.A0(net5163),
    .A1(net6471),
    .S(_07558_),
    .X(_02519_));
 sg13g2_mux2_1 _25714_ (.A0(net5069),
    .A1(net6552),
    .S(_07558_),
    .X(_02520_));
 sg13g2_mux2_1 _25715_ (.A0(net5045),
    .A1(net4336),
    .S(_07558_),
    .X(_02521_));
 sg13g2_nor2_1 _25716_ (.A(_10252_),
    .B(_04893_),
    .Y(_07559_));
 sg13g2_nor2_1 _25717_ (.A(net3203),
    .B(net4642),
    .Y(_07560_));
 sg13g2_a21oi_1 _25718_ (.A1(net5263),
    .A2(net4642),
    .Y(_02522_),
    .B1(_07560_));
 sg13g2_nor2_1 _25719_ (.A(net2999),
    .B(net4643),
    .Y(_07561_));
 sg13g2_a21oi_1 _25720_ (.A1(net5236),
    .A2(net4642),
    .Y(_02523_),
    .B1(_07561_));
 sg13g2_nor2_1 _25721_ (.A(net3256),
    .B(net4642),
    .Y(_07562_));
 sg13g2_a21oi_1 _25722_ (.A1(net5133),
    .A2(net4642),
    .Y(_02524_),
    .B1(_07562_));
 sg13g2_nor2_1 _25723_ (.A(net3144),
    .B(net4642),
    .Y(_07563_));
 sg13g2_a21oi_1 _25724_ (.A1(net5105),
    .A2(net4642),
    .Y(_02525_),
    .B1(_07563_));
 sg13g2_nor2_1 _25725_ (.A(net3249),
    .B(net4642),
    .Y(_07564_));
 sg13g2_a21oi_1 _25726_ (.A1(net5177),
    .A2(_07559_),
    .Y(_02526_),
    .B1(_07564_));
 sg13g2_nor2_1 _25727_ (.A(net3207),
    .B(net4643),
    .Y(_07565_));
 sg13g2_a21oi_1 _25728_ (.A1(net5148),
    .A2(net4643),
    .Y(_02527_),
    .B1(_07565_));
 sg13g2_nor2_1 _25729_ (.A(net3497),
    .B(net4643),
    .Y(_07566_));
 sg13g2_a21oi_1 _25730_ (.A1(net5081),
    .A2(net4643),
    .Y(_02528_),
    .B1(_07566_));
 sg13g2_nor2_1 _25731_ (.A(net3061),
    .B(net4643),
    .Y(_07567_));
 sg13g2_a21oi_1 _25732_ (.A1(net5057),
    .A2(net4643),
    .Y(_02529_),
    .B1(_07567_));
 sg13g2_nand2_2 _25733_ (.Y(_07568_),
    .A(net5423),
    .B(net5416));
 sg13g2_mux2_1 _25734_ (.A0(net5783),
    .A1(net6584),
    .S(_07568_),
    .X(_02530_));
 sg13g2_mux2_1 _25735_ (.A0(net5755),
    .A1(net4428),
    .S(_07568_),
    .X(_02531_));
 sg13g2_mux2_1 _25736_ (.A0(net5723),
    .A1(net6671),
    .S(_07568_),
    .X(_02532_));
 sg13g2_mux2_1 _25737_ (.A0(net5694),
    .A1(net6860),
    .S(_07568_),
    .X(_02533_));
 sg13g2_mux2_1 _25738_ (.A0(net5666),
    .A1(net6815),
    .S(_07568_),
    .X(_02534_));
 sg13g2_mux2_1 _25739_ (.A0(net5640),
    .A1(net6337),
    .S(_07568_),
    .X(_02535_));
 sg13g2_mux2_1 _25740_ (.A0(net5608),
    .A1(net6819),
    .S(_07568_),
    .X(_02536_));
 sg13g2_nand2_2 _25741_ (.Y(_07569_),
    .A(net4745),
    .B(_07104_));
 sg13g2_mux2_1 _25742_ (.A0(net5245),
    .A1(net4346),
    .S(_07569_),
    .X(_02537_));
 sg13g2_mux2_1 _25743_ (.A0(net5218),
    .A1(net4214),
    .S(_07569_),
    .X(_02538_));
 sg13g2_mux2_1 _25744_ (.A0(net5117),
    .A1(net6546),
    .S(_07569_),
    .X(_02539_));
 sg13g2_mux2_1 _25745_ (.A0(net5089),
    .A1(net6172),
    .S(_07569_),
    .X(_02540_));
 sg13g2_mux2_1 _25746_ (.A0(net5185),
    .A1(net6370),
    .S(_07569_),
    .X(_02541_));
 sg13g2_mux2_1 _25747_ (.A0(net5158),
    .A1(net6388),
    .S(_07569_),
    .X(_02542_));
 sg13g2_mux2_1 _25748_ (.A0(net5064),
    .A1(net6302),
    .S(_07569_),
    .X(_02543_));
 sg13g2_mux2_1 _25749_ (.A0(net5041),
    .A1(net6571),
    .S(_07569_),
    .X(_02544_));
 sg13g2_nor2b_1 _25750_ (.A(net4743),
    .B_N(_07104_),
    .Y(_07570_));
 sg13g2_nor2_1 _25751_ (.A(net3554),
    .B(net4640),
    .Y(_07571_));
 sg13g2_a21oi_1 _25752_ (.A1(net5260),
    .A2(net4640),
    .Y(_02545_),
    .B1(_07571_));
 sg13g2_nor2_1 _25753_ (.A(net3687),
    .B(net4641),
    .Y(_07572_));
 sg13g2_a21oi_1 _25754_ (.A1(net5237),
    .A2(net4641),
    .Y(_02546_),
    .B1(_07572_));
 sg13g2_nor2_1 _25755_ (.A(net3226),
    .B(net4641),
    .Y(_07573_));
 sg13g2_a21oi_1 _25756_ (.A1(net5131),
    .A2(net4641),
    .Y(_02547_),
    .B1(_07573_));
 sg13g2_nor2_1 _25757_ (.A(net3780),
    .B(net4641),
    .Y(_07574_));
 sg13g2_a21oi_1 _25758_ (.A1(net5106),
    .A2(net4641),
    .Y(_02548_),
    .B1(_07574_));
 sg13g2_nor2_1 _25759_ (.A(net3175),
    .B(net4640),
    .Y(_07575_));
 sg13g2_a21oi_1 _25760_ (.A1(net5173),
    .A2(net4640),
    .Y(_02549_),
    .B1(_07575_));
 sg13g2_nor2_1 _25761_ (.A(net3348),
    .B(net4640),
    .Y(_07576_));
 sg13g2_a21oi_1 _25762_ (.A1(net5146),
    .A2(net4640),
    .Y(_02550_),
    .B1(_07576_));
 sg13g2_nor2_1 _25763_ (.A(net3775),
    .B(net4641),
    .Y(_07577_));
 sg13g2_a21oi_1 _25764_ (.A1(net5078),
    .A2(net4641),
    .Y(_02551_),
    .B1(_07577_));
 sg13g2_nor2_1 _25765_ (.A(net3810),
    .B(net4640),
    .Y(_07578_));
 sg13g2_a21oi_1 _25766_ (.A1(net5055),
    .A2(net4640),
    .Y(_02552_),
    .B1(_07578_));
 sg13g2_nor2_1 _25767_ (.A(_03089_),
    .B(_03166_),
    .Y(_07579_));
 sg13g2_nor2_1 _25768_ (.A(net2977),
    .B(net4639),
    .Y(_07580_));
 sg13g2_a21oi_1 _25769_ (.A1(net5266),
    .A2(net4639),
    .Y(_02553_),
    .B1(_07580_));
 sg13g2_nor2_1 _25770_ (.A(net2973),
    .B(net4639),
    .Y(_07581_));
 sg13g2_a21oi_1 _25771_ (.A1(net5240),
    .A2(net4639),
    .Y(_02554_),
    .B1(_07581_));
 sg13g2_nor2_1 _25772_ (.A(net3957),
    .B(net4639),
    .Y(_07582_));
 sg13g2_a21oi_1 _25773_ (.A1(net5139),
    .A2(net4639),
    .Y(_02555_),
    .B1(_07582_));
 sg13g2_nor2_1 _25774_ (.A(net3195),
    .B(net4638),
    .Y(_07583_));
 sg13g2_a21oi_1 _25775_ (.A1(net5108),
    .A2(net4638),
    .Y(_02556_),
    .B1(_07583_));
 sg13g2_nor2_1 _25776_ (.A(net3031),
    .B(net4638),
    .Y(_07584_));
 sg13g2_a21oi_1 _25777_ (.A1(net5181),
    .A2(net4638),
    .Y(_02557_),
    .B1(_07584_));
 sg13g2_nor2_1 _25778_ (.A(net3825),
    .B(net4638),
    .Y(_07585_));
 sg13g2_a21oi_1 _25779_ (.A1(net5152),
    .A2(net4638),
    .Y(_02558_),
    .B1(_07585_));
 sg13g2_nor2_1 _25780_ (.A(net3062),
    .B(net4639),
    .Y(_07586_));
 sg13g2_a21oi_1 _25781_ (.A1(net5084),
    .A2(net4639),
    .Y(_02559_),
    .B1(_07586_));
 sg13g2_nor2_1 _25782_ (.A(net3300),
    .B(net4638),
    .Y(_07587_));
 sg13g2_a21oi_1 _25783_ (.A1(net5060),
    .A2(net4638),
    .Y(_02560_),
    .B1(_07587_));
 sg13g2_a21oi_1 _25784_ (.A1(net7122),
    .A2(net5386),
    .Y(_07588_),
    .B1(_05166_));
 sg13g2_nor2_1 _25785_ (.A(net5988),
    .B(_07588_),
    .Y(_02561_));
 sg13g2_a21oi_1 _25786_ (.A1(\atari2600.clk_counter[1] ),
    .A2(net7122),
    .Y(_07589_),
    .B1(_08133_));
 sg13g2_nand2b_1 _25787_ (.Y(_07590_),
    .B(_07589_),
    .A_N(_09655_));
 sg13g2_o21ai_1 _25788_ (.B1(net6017),
    .Y(_07591_),
    .A1(\atari2600.clk_counter[1] ),
    .A2(_08161_));
 sg13g2_a21oi_1 _25789_ (.A1(_08161_),
    .A2(_07590_),
    .Y(_02562_),
    .B1(_07591_));
 sg13g2_and3_1 _25790_ (.X(_02563_),
    .A(net2913),
    .B(net6026),
    .C(net5385));
 sg13g2_and3_1 _25791_ (.X(_02564_),
    .A(net2907),
    .B(net6026),
    .C(net5385));
 sg13g2_and3_1 _25792_ (.X(_02565_),
    .A(net2927),
    .B(net6026),
    .C(net5385));
 sg13g2_and3_1 _25793_ (.X(_02566_),
    .A(net2938),
    .B(net6026),
    .C(net5385));
 sg13g2_and3_1 _25794_ (.X(_02567_),
    .A(net2898),
    .B(net6017),
    .C(net5385));
 sg13g2_and3_1 _25795_ (.X(_02568_),
    .A(net2902),
    .B(net6017),
    .C(net5386));
 sg13g2_and2_1 _25796_ (.A(\atari2600.clk_counter[8] ),
    .B(net5386),
    .X(_07592_));
 sg13g2_nor2b_1 _25797_ (.A(net3159),
    .B_N(_07589_),
    .Y(_07593_));
 sg13g2_a22oi_1 _25798_ (.Y(_07594_),
    .B1(_07593_),
    .B2(_08669_),
    .A2(_07592_),
    .A1(net6017));
 sg13g2_inv_1 _25799_ (.Y(_02569_),
    .A(net3160));
 sg13g2_nor2_1 _25800_ (.A(net4741),
    .B(_04814_),
    .Y(_07595_));
 sg13g2_nor2_1 _25801_ (.A(net3108),
    .B(net4636),
    .Y(_07596_));
 sg13g2_a21oi_1 _25802_ (.A1(net5262),
    .A2(net4636),
    .Y(_02570_),
    .B1(_07596_));
 sg13g2_nor2_1 _25803_ (.A(net3946),
    .B(net4636),
    .Y(_07597_));
 sg13g2_a21oi_1 _25804_ (.A1(net5235),
    .A2(net4636),
    .Y(_02571_),
    .B1(_07597_));
 sg13g2_nor2_1 _25805_ (.A(net3532),
    .B(net4637),
    .Y(_07598_));
 sg13g2_a21oi_1 _25806_ (.A1(net5132),
    .A2(net4637),
    .Y(_02572_),
    .B1(_07598_));
 sg13g2_nor2_1 _25807_ (.A(net3849),
    .B(net4636),
    .Y(_07599_));
 sg13g2_a21oi_1 _25808_ (.A1(net5104),
    .A2(net4636),
    .Y(_02573_),
    .B1(_07599_));
 sg13g2_nor2_1 _25809_ (.A(net3835),
    .B(net4637),
    .Y(_07600_));
 sg13g2_a21oi_1 _25810_ (.A1(net5176),
    .A2(net4637),
    .Y(_02574_),
    .B1(_07600_));
 sg13g2_nor2_1 _25811_ (.A(net3359),
    .B(net4636),
    .Y(_07601_));
 sg13g2_a21oi_1 _25812_ (.A1(net5147),
    .A2(net4636),
    .Y(_02575_),
    .B1(_07601_));
 sg13g2_nor2_1 _25813_ (.A(net3454),
    .B(net4637),
    .Y(_07602_));
 sg13g2_a21oi_1 _25814_ (.A1(net5079),
    .A2(net4637),
    .Y(_02576_),
    .B1(_07602_));
 sg13g2_nor2_1 _25815_ (.A(net3064),
    .B(net4637),
    .Y(_07603_));
 sg13g2_a21oi_1 _25816_ (.A1(net5056),
    .A2(net4637),
    .Y(_02577_),
    .B1(_07603_));
 sg13g2_nor2_1 _25817_ (.A(_03004_),
    .B(net4742),
    .Y(_07604_));
 sg13g2_nor2_1 _25818_ (.A(net3275),
    .B(net4634),
    .Y(_07605_));
 sg13g2_a21oi_1 _25819_ (.A1(net5261),
    .A2(net4634),
    .Y(_02578_),
    .B1(_07605_));
 sg13g2_nor2_1 _25820_ (.A(net3697),
    .B(net4634),
    .Y(_07606_));
 sg13g2_a21oi_1 _25821_ (.A1(net5235),
    .A2(net4634),
    .Y(_02579_),
    .B1(_07606_));
 sg13g2_nor2_1 _25822_ (.A(net3382),
    .B(net4635),
    .Y(_07607_));
 sg13g2_a21oi_1 _25823_ (.A1(net5133),
    .A2(net4635),
    .Y(_02580_),
    .B1(_07607_));
 sg13g2_nor2_1 _25824_ (.A(net3953),
    .B(net4635),
    .Y(_07608_));
 sg13g2_a21oi_1 _25825_ (.A1(net5104),
    .A2(net4635),
    .Y(_02581_),
    .B1(_07608_));
 sg13g2_nor2_1 _25826_ (.A(net3125),
    .B(net4635),
    .Y(_07609_));
 sg13g2_a21oi_1 _25827_ (.A1(net5177),
    .A2(_07604_),
    .Y(_02582_),
    .B1(_07609_));
 sg13g2_nor2_1 _25828_ (.A(net4211),
    .B(net4634),
    .Y(_07610_));
 sg13g2_a21oi_1 _25829_ (.A1(net5148),
    .A2(net4634),
    .Y(_02583_),
    .B1(_07610_));
 sg13g2_nor2_1 _25830_ (.A(net3880),
    .B(net4635),
    .Y(_07611_));
 sg13g2_a21oi_1 _25831_ (.A1(net5080),
    .A2(net4635),
    .Y(_02584_),
    .B1(_07611_));
 sg13g2_nor2_1 _25832_ (.A(net3176),
    .B(net4634),
    .Y(_07612_));
 sg13g2_a21oi_1 _25833_ (.A1(net5056),
    .A2(net4634),
    .Y(_02585_),
    .B1(_07612_));
 sg13g2_nor2_1 _25834_ (.A(net7138),
    .B(\hvsync_gen.vga.vpos[0] ),
    .Y(_07613_));
 sg13g2_nand3_1 _25835_ (.B(\hvsync_gen.vga.vpos[2] ),
    .C(_07613_),
    .A(\hvsync_gen.vga.vpos[3] ),
    .Y(_07614_));
 sg13g2_nor4_1 _25836_ (.A(_08047_),
    .B(\hvsync_gen.vga.vpos[5] ),
    .C(\hvsync_gen.vga.vpos[4] ),
    .D(_07614_),
    .Y(_07615_));
 sg13g2_a21o_1 _25837_ (.A2(_07615_),
    .A1(_08493_),
    .B1(net5989),
    .X(_07616_));
 sg13g2_or2_1 _25838_ (.X(_07617_),
    .B(_07616_),
    .A(_03229_));
 sg13g2_inv_1 _25839_ (.Y(_07618_),
    .A(_07617_));
 sg13g2_a22oi_1 _25840_ (.Y(_07619_),
    .B1(_07618_),
    .B2(net2893),
    .A2(_03230_),
    .A1(\hvsync_gen.vga.vpos[0] ));
 sg13g2_inv_1 _25841_ (.Y(_02586_),
    .A(net2894));
 sg13g2_and2_1 _25842_ (.A(net7138),
    .B(\hvsync_gen.vga.vpos[0] ),
    .X(_07620_));
 sg13g2_nor3_1 _25843_ (.A(_07613_),
    .B(_07617_),
    .C(_07620_),
    .Y(_07621_));
 sg13g2_a21o_1 _25844_ (.A2(_03230_),
    .A1(net7138),
    .B1(_07621_),
    .X(_02587_));
 sg13g2_and3_1 _25845_ (.X(_07622_),
    .A(net7163),
    .B(_03231_),
    .C(_07620_));
 sg13g2_and2_2 _25846_ (.A(_03231_),
    .B(_07616_),
    .X(_07623_));
 sg13g2_a21oi_1 _25847_ (.A1(_03231_),
    .A2(_07620_),
    .Y(_07624_),
    .B1(net7163));
 sg13g2_nor3_1 _25848_ (.A(_07622_),
    .B(_07623_),
    .C(_07624_),
    .Y(_02588_));
 sg13g2_nor2_1 _25849_ (.A(net7236),
    .B(_07622_),
    .Y(_07625_));
 sg13g2_and2_1 _25850_ (.A(net7236),
    .B(_07622_),
    .X(_07626_));
 sg13g2_nor3_1 _25851_ (.A(_07623_),
    .B(_07625_),
    .C(_07626_),
    .Y(_02589_));
 sg13g2_nor2_1 _25852_ (.A(net7147),
    .B(_07626_),
    .Y(_07627_));
 sg13g2_nand4_1 _25853_ (.B(\hvsync_gen.vga.vpos[3] ),
    .C(\hvsync_gen.vga.vpos[2] ),
    .A(net7147),
    .Y(_07628_),
    .D(_07620_));
 sg13g2_nor2_1 _25854_ (.A(_03230_),
    .B(_07628_),
    .Y(_07629_));
 sg13g2_nor3_1 _25855_ (.A(_07623_),
    .B(net7148),
    .C(_07629_),
    .Y(_02590_));
 sg13g2_and2_1 _25856_ (.A(net7187),
    .B(_07629_),
    .X(_07630_));
 sg13g2_nor2_1 _25857_ (.A(net7187),
    .B(_07629_),
    .Y(_07631_));
 sg13g2_nor3_1 _25858_ (.A(_07623_),
    .B(_07630_),
    .C(net7188),
    .Y(_02591_));
 sg13g2_xnor2_1 _25859_ (.Y(_07632_),
    .A(net7218),
    .B(_07630_));
 sg13g2_nor2_1 _25860_ (.A(_07623_),
    .B(_07632_),
    .Y(_02592_));
 sg13g2_and3_1 _25861_ (.X(_07633_),
    .A(net7039),
    .B(net7376),
    .C(_07630_));
 sg13g2_a21oi_1 _25862_ (.A1(\hvsync_gen.vga.vpos[6] ),
    .A2(_07630_),
    .Y(_07634_),
    .B1(net7039));
 sg13g2_nor3_1 _25863_ (.A(_07623_),
    .B(_07633_),
    .C(net7040),
    .Y(_02593_));
 sg13g2_a21oi_1 _25864_ (.A1(net7176),
    .A2(_07633_),
    .Y(_07635_),
    .B1(_07623_));
 sg13g2_o21ai_1 _25865_ (.B1(_07635_),
    .Y(_07636_),
    .A1(net7176),
    .A2(_07633_));
 sg13g2_inv_1 _25866_ (.Y(_02594_),
    .A(_07636_));
 sg13g2_nor4_1 _25867_ (.A(net7142),
    .B(_08699_),
    .C(_07617_),
    .D(_07628_),
    .Y(_07637_));
 sg13g2_a21o_1 _25868_ (.A2(_07635_),
    .A1(net7142),
    .B1(_07637_),
    .X(_02595_));
 sg13g2_o21ai_1 _25869_ (.B1(net5999),
    .Y(_07638_),
    .A1(net5537),
    .A2(_10444_));
 sg13g2_and2_1 _25870_ (.A(_08077_),
    .B(_10349_),
    .X(_07639_));
 sg13g2_nand2_1 _25871_ (.Y(_07640_),
    .A(_08077_),
    .B(_10349_));
 sg13g2_nand2_1 _25872_ (.Y(_07641_),
    .A(net5567),
    .B(_10352_));
 sg13g2_nor3_2 _25873_ (.A(net7199),
    .B(\flash_rom.nibbles_remaining[1] ),
    .C(net7174),
    .Y(_07642_));
 sg13g2_nand4_1 _25874_ (.B(net5567),
    .C(_10352_),
    .A(net7229),
    .Y(_07643_),
    .D(_07642_));
 sg13g2_a21oi_1 _25875_ (.A1(_07640_),
    .A2(net7230),
    .Y(_02596_),
    .B1(net4572));
 sg13g2_nand2_2 _25876_ (.Y(_07644_),
    .A(net4748),
    .B(_03041_));
 sg13g2_mux2_1 _25877_ (.A0(net5251),
    .A1(net6378),
    .S(_07644_),
    .X(_02597_));
 sg13g2_mux2_1 _25878_ (.A0(net5225),
    .A1(net4500),
    .S(_07644_),
    .X(_02598_));
 sg13g2_mux2_1 _25879_ (.A0(net5124),
    .A1(net4474),
    .S(_07644_),
    .X(_02599_));
 sg13g2_mux2_1 _25880_ (.A0(net5095),
    .A1(net6743),
    .S(_07644_),
    .X(_02600_));
 sg13g2_mux2_1 _25881_ (.A0(net5190),
    .A1(net4525),
    .S(_07644_),
    .X(_02601_));
 sg13g2_mux2_1 _25882_ (.A0(net5163),
    .A1(net4338),
    .S(_07644_),
    .X(_02602_));
 sg13g2_mux2_1 _25883_ (.A0(net5071),
    .A1(net4341),
    .S(_07644_),
    .X(_02603_));
 sg13g2_mux2_1 _25884_ (.A0(net5045),
    .A1(net6237),
    .S(_07644_),
    .X(_02604_));
 sg13g2_nand2_2 _25885_ (.Y(_07645_),
    .A(net4739),
    .B(_05071_));
 sg13g2_mux2_1 _25886_ (.A0(net5245),
    .A1(net6358),
    .S(_07645_),
    .X(_02605_));
 sg13g2_mux2_1 _25887_ (.A0(net5217),
    .A1(net6206),
    .S(_07645_),
    .X(_02606_));
 sg13g2_mux2_1 _25888_ (.A0(net5115),
    .A1(net4239),
    .S(_07645_),
    .X(_02607_));
 sg13g2_mux2_1 _25889_ (.A0(net5088),
    .A1(net4277),
    .S(_07645_),
    .X(_02608_));
 sg13g2_mux2_1 _25890_ (.A0(net5185),
    .A1(net4065),
    .S(_07645_),
    .X(_02609_));
 sg13g2_mux2_1 _25891_ (.A0(net5158),
    .A1(net6626),
    .S(_07645_),
    .X(_02610_));
 sg13g2_mux2_1 _25892_ (.A0(net5065),
    .A1(net6040),
    .S(_07645_),
    .X(_02611_));
 sg13g2_mux2_1 _25893_ (.A0(net5041),
    .A1(net4157),
    .S(_07645_),
    .X(_02612_));
 sg13g2_nor2b_1 _25894_ (.A(net4741),
    .B_N(net4763),
    .Y(_07646_));
 sg13g2_nor2_1 _25895_ (.A(net3800),
    .B(net4633),
    .Y(_07647_));
 sg13g2_a21oi_1 _25896_ (.A1(net5261),
    .A2(net4633),
    .Y(_02613_),
    .B1(_07647_));
 sg13g2_nor2_1 _25897_ (.A(net3692),
    .B(net4633),
    .Y(_07648_));
 sg13g2_a21oi_1 _25898_ (.A1(net5236),
    .A2(net4633),
    .Y(_02614_),
    .B1(_07648_));
 sg13g2_nor2_1 _25899_ (.A(net3174),
    .B(net4633),
    .Y(_07649_));
 sg13g2_a21oi_1 _25900_ (.A1(net5132),
    .A2(net4633),
    .Y(_02615_),
    .B1(_07649_));
 sg13g2_nor2_1 _25901_ (.A(net3773),
    .B(_07646_),
    .Y(_07650_));
 sg13g2_a21oi_1 _25902_ (.A1(net5104),
    .A2(net4633),
    .Y(_02616_),
    .B1(_07650_));
 sg13g2_nor2_1 _25903_ (.A(net3252),
    .B(net4632),
    .Y(_07651_));
 sg13g2_a21oi_1 _25904_ (.A1(net5176),
    .A2(net4632),
    .Y(_02617_),
    .B1(_07651_));
 sg13g2_nor2_1 _25905_ (.A(net3253),
    .B(net4632),
    .Y(_07652_));
 sg13g2_a21oi_1 _25906_ (.A1(net5148),
    .A2(net4632),
    .Y(_02618_),
    .B1(_07652_));
 sg13g2_nor2_1 _25907_ (.A(net4499),
    .B(net4632),
    .Y(_07653_));
 sg13g2_a21oi_1 _25908_ (.A1(net5078),
    .A2(net4632),
    .Y(_02619_),
    .B1(_07653_));
 sg13g2_nor2_1 _25909_ (.A(net3472),
    .B(net4632),
    .Y(_07654_));
 sg13g2_a21oi_1 _25910_ (.A1(net5057),
    .A2(net4632),
    .Y(_02620_),
    .B1(_07654_));
 sg13g2_nor2_1 _25911_ (.A(_03042_),
    .B(net4743),
    .Y(_07655_));
 sg13g2_nor2_1 _25912_ (.A(net3576),
    .B(_07655_),
    .Y(_07656_));
 sg13g2_a21oi_1 _25913_ (.A1(net5263),
    .A2(net4631),
    .Y(_02621_),
    .B1(_07656_));
 sg13g2_nor2_1 _25914_ (.A(net3898),
    .B(net4630),
    .Y(_07657_));
 sg13g2_a21oi_1 _25915_ (.A1(net5234),
    .A2(net4630),
    .Y(_02622_),
    .B1(_07657_));
 sg13g2_nor2_1 _25916_ (.A(net3082),
    .B(net4631),
    .Y(_07658_));
 sg13g2_a21oi_1 _25917_ (.A1(net5131),
    .A2(net4631),
    .Y(_02623_),
    .B1(_07658_));
 sg13g2_nor2_1 _25918_ (.A(net3890),
    .B(net4630),
    .Y(_07659_));
 sg13g2_a21oi_1 _25919_ (.A1(net5105),
    .A2(net4630),
    .Y(_02624_),
    .B1(_07659_));
 sg13g2_nor2_1 _25920_ (.A(net3863),
    .B(net4631),
    .Y(_07660_));
 sg13g2_a21oi_1 _25921_ (.A1(net5177),
    .A2(net4631),
    .Y(_02625_),
    .B1(_07660_));
 sg13g2_nor2_1 _25922_ (.A(net4053),
    .B(net4631),
    .Y(_07661_));
 sg13g2_a21oi_1 _25923_ (.A1(net5146),
    .A2(net4631),
    .Y(_02626_),
    .B1(_07661_));
 sg13g2_nor2_1 _25924_ (.A(net3366),
    .B(net4630),
    .Y(_07662_));
 sg13g2_a21oi_1 _25925_ (.A1(net5080),
    .A2(net4630),
    .Y(_02627_),
    .B1(_07662_));
 sg13g2_nor2_1 _25926_ (.A(net3188),
    .B(net4630),
    .Y(_07663_));
 sg13g2_a21oi_1 _25927_ (.A1(net5058),
    .A2(net4630),
    .Y(_02628_),
    .B1(_07663_));
 sg13g2_nand2_1 _25928_ (.Y(_07664_),
    .A(net4735),
    .B(_05071_));
 sg13g2_mux2_1 _25929_ (.A0(net5245),
    .A1(net6420),
    .S(net4629),
    .X(_02629_));
 sg13g2_mux2_1 _25930_ (.A0(net5217),
    .A1(net6325),
    .S(net4629),
    .X(_02630_));
 sg13g2_mux2_1 _25931_ (.A0(net5115),
    .A1(net6048),
    .S(net4629),
    .X(_02631_));
 sg13g2_mux2_1 _25932_ (.A0(net5088),
    .A1(net6458),
    .S(net4629),
    .X(_02632_));
 sg13g2_nand2_1 _25933_ (.Y(_07665_),
    .A(net2951),
    .B(net4629));
 sg13g2_o21ai_1 _25934_ (.B1(_07665_),
    .Y(_02633_),
    .A1(net5175),
    .A2(net4629));
 sg13g2_mux2_1 _25935_ (.A0(net5158),
    .A1(net6580),
    .S(net4629),
    .X(_02634_));
 sg13g2_mux2_1 _25936_ (.A0(net5064),
    .A1(net6185),
    .S(_07664_),
    .X(_02635_));
 sg13g2_mux2_1 _25937_ (.A0(net5041),
    .A1(net6228),
    .S(net4629),
    .X(_02636_));
 sg13g2_nand2_1 _25938_ (.Y(_07666_),
    .A(_03041_),
    .B(net4735));
 sg13g2_mux2_1 _25939_ (.A0(net5251),
    .A1(net6881),
    .S(net4628),
    .X(_02637_));
 sg13g2_mux2_1 _25940_ (.A0(net5224),
    .A1(net4235),
    .S(_07666_),
    .X(_02638_));
 sg13g2_mux2_1 _25941_ (.A0(net5124),
    .A1(net4100),
    .S(net4628),
    .X(_02639_));
 sg13g2_mux2_1 _25942_ (.A0(net5094),
    .A1(net6393),
    .S(net4628),
    .X(_02640_));
 sg13g2_nand2_1 _25943_ (.Y(_07667_),
    .A(net2942),
    .B(net4628));
 sg13g2_o21ai_1 _25944_ (.B1(_07667_),
    .Y(_02641_),
    .A1(net5177),
    .A2(net4628));
 sg13g2_mux2_1 _25945_ (.A0(net5159),
    .A1(net4027),
    .S(net4628),
    .X(_02642_));
 sg13g2_mux2_1 _25946_ (.A0(net5066),
    .A1(net6862),
    .S(net4628),
    .X(_02643_));
 sg13g2_mux2_1 _25947_ (.A0(net5043),
    .A1(net6103),
    .S(net4628),
    .X(_02644_));
 sg13g2_nand2_1 _25948_ (.Y(_07668_),
    .A(net4745),
    .B(_05071_));
 sg13g2_mux2_1 _25949_ (.A0(net5245),
    .A1(net4314),
    .S(net4627),
    .X(_02645_));
 sg13g2_mux2_1 _25950_ (.A0(net5217),
    .A1(net4295),
    .S(net4627),
    .X(_02646_));
 sg13g2_mux2_1 _25951_ (.A0(net5115),
    .A1(net4285),
    .S(net4627),
    .X(_02647_));
 sg13g2_mux2_1 _25952_ (.A0(net5088),
    .A1(net6273),
    .S(net4627),
    .X(_02648_));
 sg13g2_nand2_1 _25953_ (.Y(_07669_),
    .A(net2928),
    .B(net4627));
 sg13g2_o21ai_1 _25954_ (.B1(_07669_),
    .Y(_02649_),
    .A1(net5173),
    .A2(net4627));
 sg13g2_mux2_1 _25955_ (.A0(net5158),
    .A1(net6132),
    .S(net4627),
    .X(_02650_));
 sg13g2_mux2_1 _25956_ (.A0(net5064),
    .A1(net6825),
    .S(_07668_),
    .X(_02651_));
 sg13g2_mux2_1 _25957_ (.A0(net5041),
    .A1(net6419),
    .S(net4627),
    .X(_02652_));
 sg13g2_nand2_2 _25958_ (.Y(_07670_),
    .A(_08515_),
    .B(_05028_));
 sg13g2_mux2_1 _25959_ (.A0(_05031_),
    .A1(net3804),
    .S(_07670_),
    .X(_02653_));
 sg13g2_mux2_1 _25960_ (.A0(_05038_),
    .A1(net3923),
    .S(_07670_),
    .X(_02654_));
 sg13g2_mux2_1 _25961_ (.A0(_05044_),
    .A1(net6045),
    .S(_07670_),
    .X(_02655_));
 sg13g2_mux2_1 _25962_ (.A0(_05049_),
    .A1(net6673),
    .S(_07670_),
    .X(_02656_));
 sg13g2_mux2_1 _25963_ (.A0(_05051_),
    .A1(net4425),
    .S(_07670_),
    .X(_02657_));
 sg13g2_mux2_1 _25964_ (.A0(_05057_),
    .A1(net6122),
    .S(_07670_),
    .X(_02658_));
 sg13g2_mux2_1 _25965_ (.A0(_05063_),
    .A1(net6785),
    .S(_07670_),
    .X(_02659_));
 sg13g2_mux2_1 _25966_ (.A0(_05068_),
    .A1(net6482),
    .S(_07670_),
    .X(_02660_));
 sg13g2_nand2_1 _25967_ (.Y(_07671_),
    .A(_04813_),
    .B(net4733));
 sg13g2_mux2_1 _25968_ (.A0(net5254),
    .A1(net4378),
    .S(net4577),
    .X(_02661_));
 sg13g2_mux2_1 _25969_ (.A0(net5222),
    .A1(net4496),
    .S(net4577),
    .X(_02662_));
 sg13g2_mux2_1 _25970_ (.A0(net5119),
    .A1(net6685),
    .S(_07671_),
    .X(_02663_));
 sg13g2_mux2_1 _25971_ (.A0(net5093),
    .A1(net4354),
    .S(net4577),
    .X(_02664_));
 sg13g2_nand2_1 _25972_ (.Y(_07672_),
    .A(net2914),
    .B(net4577));
 sg13g2_o21ai_1 _25973_ (.B1(_07672_),
    .Y(_02665_),
    .A1(net5176),
    .A2(net4577));
 sg13g2_mux2_1 _25974_ (.A0(net5162),
    .A1(net4177),
    .S(net4577),
    .X(_02666_));
 sg13g2_mux2_1 _25975_ (.A0(net5069),
    .A1(net4537),
    .S(net4577),
    .X(_02667_));
 sg13g2_mux2_1 _25976_ (.A0(net5047),
    .A1(net6130),
    .S(net4577),
    .X(_02668_));
 sg13g2_nor2b_1 _25977_ (.A(net4743),
    .B_N(_05073_),
    .Y(_07673_));
 sg13g2_nor2_1 _25978_ (.A(net4096),
    .B(net4626),
    .Y(_07674_));
 sg13g2_a21oi_1 _25979_ (.A1(net5260),
    .A2(net4626),
    .Y(_02669_),
    .B1(_07674_));
 sg13g2_nor2_1 _25980_ (.A(net3652),
    .B(net4625),
    .Y(_07675_));
 sg13g2_a21oi_1 _25981_ (.A1(net5234),
    .A2(net4625),
    .Y(_02670_),
    .B1(_07675_));
 sg13g2_nor2_1 _25982_ (.A(net4064),
    .B(net4625),
    .Y(_07676_));
 sg13g2_a21oi_1 _25983_ (.A1(net5134),
    .A2(net4625),
    .Y(_02671_),
    .B1(_07676_));
 sg13g2_nor2_1 _25984_ (.A(net3530),
    .B(net4625),
    .Y(_07677_));
 sg13g2_a21oi_1 _25985_ (.A1(net5103),
    .A2(net4625),
    .Y(_02672_),
    .B1(_07677_));
 sg13g2_mux2_1 _25986_ (.A0(net3533),
    .A1(net5186),
    .S(net4625),
    .X(_02673_));
 sg13g2_nor2_1 _25987_ (.A(net3663),
    .B(net4626),
    .Y(_07678_));
 sg13g2_a21oi_1 _25988_ (.A1(net5146),
    .A2(net4626),
    .Y(_02674_),
    .B1(_07678_));
 sg13g2_nor2_1 _25989_ (.A(net3124),
    .B(net4626),
    .Y(_07679_));
 sg13g2_a21oi_1 _25990_ (.A1(net5080),
    .A2(net4625),
    .Y(_02675_),
    .B1(_07679_));
 sg13g2_nor2_1 _25991_ (.A(net3596),
    .B(net4626),
    .Y(_07680_));
 sg13g2_a21oi_1 _25992_ (.A1(net5055),
    .A2(net4626),
    .Y(_02676_),
    .B1(_07680_));
 sg13g2_nand2_1 _25993_ (.Y(_07681_),
    .A(net4745),
    .B(_05073_));
 sg13g2_mux2_1 _25994_ (.A0(net5248),
    .A1(net6336),
    .S(_07681_),
    .X(_02677_));
 sg13g2_mux2_1 _25995_ (.A0(net5221),
    .A1(net6348),
    .S(net4624),
    .X(_02678_));
 sg13g2_mux2_1 _25996_ (.A0(net5120),
    .A1(net6171),
    .S(net4624),
    .X(_02679_));
 sg13g2_mux2_1 _25997_ (.A0(net5092),
    .A1(net6601),
    .S(net4624),
    .X(_02680_));
 sg13g2_nand2_1 _25998_ (.Y(_07682_),
    .A(net2912),
    .B(net4624));
 sg13g2_o21ai_1 _25999_ (.B1(_07682_),
    .Y(_02681_),
    .A1(net5175),
    .A2(net4624));
 sg13g2_mux2_1 _26000_ (.A0(net5159),
    .A1(net4517),
    .S(net4624),
    .X(_02682_));
 sg13g2_mux2_1 _26001_ (.A0(net5066),
    .A1(net4379),
    .S(net4624),
    .X(_02683_));
 sg13g2_mux2_1 _26002_ (.A0(net5044),
    .A1(net6403),
    .S(net4624),
    .X(_02684_));
 sg13g2_nand2_1 _26003_ (.Y(_07683_),
    .A(net4734),
    .B(_05073_));
 sg13g2_mux2_1 _26004_ (.A0(net5247),
    .A1(net4113),
    .S(_07683_),
    .X(_02685_));
 sg13g2_mux2_1 _26005_ (.A0(net5220),
    .A1(net6509),
    .S(net4623),
    .X(_02686_));
 sg13g2_mux2_1 _26006_ (.A0(net5121),
    .A1(net4270),
    .S(net4623),
    .X(_02687_));
 sg13g2_mux2_1 _26007_ (.A0(net5091),
    .A1(net4320),
    .S(net4623),
    .X(_02688_));
 sg13g2_nand2_1 _26008_ (.Y(_07684_),
    .A(net2921),
    .B(net4623));
 sg13g2_o21ai_1 _26009_ (.B1(_07684_),
    .Y(_02689_),
    .A1(net5174),
    .A2(net4623));
 sg13g2_mux2_1 _26010_ (.A0(net5160),
    .A1(net4498),
    .S(net4623),
    .X(_02690_));
 sg13g2_mux2_1 _26011_ (.A0(net5066),
    .A1(net6400),
    .S(net4623),
    .X(_02691_));
 sg13g2_mux2_1 _26012_ (.A0(net5043),
    .A1(net6795),
    .S(net4623),
    .X(_02692_));
 sg13g2_nand2_1 _26013_ (.Y(_07685_),
    .A(net4738),
    .B(_05073_));
 sg13g2_mux2_1 _26014_ (.A0(net5247),
    .A1(net6244),
    .S(net4622),
    .X(_02693_));
 sg13g2_mux2_1 _26015_ (.A0(net5220),
    .A1(net3985),
    .S(net4622),
    .X(_02694_));
 sg13g2_mux2_1 _26016_ (.A0(net5120),
    .A1(net6368),
    .S(net4622),
    .X(_02695_));
 sg13g2_mux2_1 _26017_ (.A0(net5091),
    .A1(net4056),
    .S(_07685_),
    .X(_02696_));
 sg13g2_nand2_1 _26018_ (.Y(_07686_),
    .A(net2909),
    .B(net4622));
 sg13g2_o21ai_1 _26019_ (.B1(_07686_),
    .Y(_02697_),
    .A1(net5174),
    .A2(net4622));
 sg13g2_mux2_1 _26020_ (.A0(net5159),
    .A1(net4208),
    .S(net4622),
    .X(_02698_));
 sg13g2_mux2_1 _26021_ (.A0(net5067),
    .A1(net6178),
    .S(net4622),
    .X(_02699_));
 sg13g2_mux2_1 _26022_ (.A0(net5049),
    .A1(net6054),
    .S(net4622),
    .X(_02700_));
 sg13g2_nor2b_1 _26023_ (.A(net4742),
    .B_N(_05073_),
    .Y(_07687_));
 sg13g2_nor2_1 _26024_ (.A(net4159),
    .B(net4621),
    .Y(_07688_));
 sg13g2_a21oi_1 _26025_ (.A1(net5260),
    .A2(net4621),
    .Y(_02701_),
    .B1(_07688_));
 sg13g2_nor2_1 _26026_ (.A(net3668),
    .B(net4620),
    .Y(_07689_));
 sg13g2_a21oi_1 _26027_ (.A1(net5234),
    .A2(net4620),
    .Y(_02702_),
    .B1(_07689_));
 sg13g2_nor2_1 _26028_ (.A(net3011),
    .B(net4620),
    .Y(_07690_));
 sg13g2_a21oi_1 _26029_ (.A1(net5131),
    .A2(net4620),
    .Y(_02703_),
    .B1(_07690_));
 sg13g2_nor2_1 _26030_ (.A(net3106),
    .B(net4621),
    .Y(_07691_));
 sg13g2_a21oi_1 _26031_ (.A1(net5106),
    .A2(net4620),
    .Y(_02704_),
    .B1(_07691_));
 sg13g2_mux2_1 _26032_ (.A0(net3197),
    .A1(net5186),
    .S(net4620),
    .X(_02705_));
 sg13g2_nor2_1 _26033_ (.A(net3262),
    .B(net4621),
    .Y(_07692_));
 sg13g2_a21oi_1 _26034_ (.A1(net5150),
    .A2(net4621),
    .Y(_02706_),
    .B1(_07692_));
 sg13g2_nor2_1 _26035_ (.A(net3149),
    .B(net4621),
    .Y(_07693_));
 sg13g2_a21oi_1 _26036_ (.A1(net5080),
    .A2(net4621),
    .Y(_02707_),
    .B1(_07693_));
 sg13g2_nor2_1 _26037_ (.A(net3632),
    .B(net4620),
    .Y(_07694_));
 sg13g2_a21oi_1 _26038_ (.A1(net5055),
    .A2(net4620),
    .Y(_02708_),
    .B1(_07694_));
 sg13g2_nand2_1 _26039_ (.Y(_07695_),
    .A(net4747),
    .B(_05073_));
 sg13g2_mux2_1 _26040_ (.A0(net5247),
    .A1(net6207),
    .S(_07695_),
    .X(_02709_));
 sg13g2_mux2_1 _26041_ (.A0(net5220),
    .A1(net4016),
    .S(net4619),
    .X(_02710_));
 sg13g2_mux2_1 _26042_ (.A0(net5120),
    .A1(net4375),
    .S(net4619),
    .X(_02711_));
 sg13g2_mux2_1 _26043_ (.A0(net5091),
    .A1(net4025),
    .S(net4619),
    .X(_02712_));
 sg13g2_nand2_1 _26044_ (.Y(_07696_),
    .A(net2955),
    .B(net4619));
 sg13g2_o21ai_1 _26045_ (.B1(_07696_),
    .Y(_02713_),
    .A1(net5174),
    .A2(net4619));
 sg13g2_mux2_1 _26046_ (.A0(net5159),
    .A1(net4237),
    .S(net4619),
    .X(_02714_));
 sg13g2_mux2_1 _26047_ (.A0(net5066),
    .A1(net6457),
    .S(net4619),
    .X(_02715_));
 sg13g2_mux2_1 _26048_ (.A0(net5049),
    .A1(net4306),
    .S(net4619),
    .X(_02716_));
 sg13g2_nand2_1 _26049_ (.Y(_07697_),
    .A(net4739),
    .B(_05075_));
 sg13g2_mux2_1 _26050_ (.A0(net5246),
    .A1(net4326),
    .S(_07697_),
    .X(_02717_));
 sg13g2_mux2_1 _26051_ (.A0(net5220),
    .A1(net4465),
    .S(net4618),
    .X(_02718_));
 sg13g2_mux2_1 _26052_ (.A0(net5117),
    .A1(net4304),
    .S(net4618),
    .X(_02719_));
 sg13g2_mux2_1 _26053_ (.A0(net5091),
    .A1(net6076),
    .S(net4618),
    .X(_02720_));
 sg13g2_nand2_1 _26054_ (.Y(_07698_),
    .A(net2961),
    .B(net4618));
 sg13g2_o21ai_1 _26055_ (.B1(_07698_),
    .Y(_02721_),
    .A1(net5174),
    .A2(net4618));
 sg13g2_mux2_1 _26056_ (.A0(net5160),
    .A1(net4309),
    .S(net4618),
    .X(_02722_));
 sg13g2_mux2_1 _26057_ (.A0(net5067),
    .A1(net4193),
    .S(net4618),
    .X(_02723_));
 sg13g2_mux2_1 _26058_ (.A0(net5043),
    .A1(net4122),
    .S(net4618),
    .X(_02724_));
 sg13g2_nand2_1 _26059_ (.Y(_07699_),
    .A(net4735),
    .B(_05075_));
 sg13g2_mux2_1 _26060_ (.A0(net5246),
    .A1(net4424),
    .S(_07699_),
    .X(_02725_));
 sg13g2_mux2_1 _26061_ (.A0(net5220),
    .A1(net4312),
    .S(net4617),
    .X(_02726_));
 sg13g2_mux2_1 _26062_ (.A0(net5120),
    .A1(net6309),
    .S(net4617),
    .X(_02727_));
 sg13g2_mux2_1 _26063_ (.A0(net5091),
    .A1(net4128),
    .S(net4617),
    .X(_02728_));
 sg13g2_nand2_1 _26064_ (.Y(_07700_),
    .A(net2919),
    .B(net4617));
 sg13g2_o21ai_1 _26065_ (.B1(_07700_),
    .Y(_02729_),
    .A1(net5174),
    .A2(net4617));
 sg13g2_mux2_1 _26066_ (.A0(net5160),
    .A1(net4347),
    .S(net4617),
    .X(_02730_));
 sg13g2_mux2_1 _26067_ (.A0(net5067),
    .A1(net6445),
    .S(net4617),
    .X(_02731_));
 sg13g2_mux2_1 _26068_ (.A0(net5043),
    .A1(net6213),
    .S(net4617),
    .X(_02732_));
 sg13g2_nor2b_1 _26069_ (.A(net4743),
    .B_N(_05075_),
    .Y(_07701_));
 sg13g2_nor2_1 _26070_ (.A(net3052),
    .B(net4616),
    .Y(_07702_));
 sg13g2_a21oi_1 _26071_ (.A1(net5260),
    .A2(net4616),
    .Y(_02733_),
    .B1(_07702_));
 sg13g2_nor2_1 _26072_ (.A(net3053),
    .B(net4615),
    .Y(_07703_));
 sg13g2_a21oi_1 _26073_ (.A1(net5234),
    .A2(net4615),
    .Y(_02734_),
    .B1(_07703_));
 sg13g2_nor2_1 _26074_ (.A(net3040),
    .B(net4615),
    .Y(_07704_));
 sg13g2_a21oi_1 _26075_ (.A1(net5134),
    .A2(net4615),
    .Y(_02735_),
    .B1(_07704_));
 sg13g2_nor2_1 _26076_ (.A(net3759),
    .B(net4615),
    .Y(_07705_));
 sg13g2_a21oi_1 _26077_ (.A1(net5103),
    .A2(net4615),
    .Y(_02736_),
    .B1(_07705_));
 sg13g2_mux2_1 _26078_ (.A0(net3179),
    .A1(net5186),
    .S(net4615),
    .X(_02737_));
 sg13g2_nor2_1 _26079_ (.A(net3960),
    .B(net4616),
    .Y(_07706_));
 sg13g2_a21oi_1 _26080_ (.A1(net5146),
    .A2(net4616),
    .Y(_02738_),
    .B1(_07706_));
 sg13g2_nor2_1 _26081_ (.A(net3193),
    .B(net4616),
    .Y(_07707_));
 sg13g2_a21oi_1 _26082_ (.A1(net5080),
    .A2(net4615),
    .Y(_02739_),
    .B1(_07707_));
 sg13g2_nor2_1 _26083_ (.A(net3030),
    .B(net4616),
    .Y(_07708_));
 sg13g2_a21oi_1 _26084_ (.A1(net5055),
    .A2(net4616),
    .Y(_02740_),
    .B1(_07708_));
 sg13g2_nand2_1 _26085_ (.Y(_07709_),
    .A(net4737),
    .B(_04813_));
 sg13g2_mux2_1 _26086_ (.A0(net5254),
    .A1(net4034),
    .S(net4576),
    .X(_02741_));
 sg13g2_mux2_1 _26087_ (.A0(net5222),
    .A1(net4174),
    .S(net4576),
    .X(_02742_));
 sg13g2_mux2_1 _26088_ (.A0(net5119),
    .A1(net4152),
    .S(net4576),
    .X(_02743_));
 sg13g2_mux2_1 _26089_ (.A0(net5093),
    .A1(net6421),
    .S(net4576),
    .X(_02744_));
 sg13g2_nand2_1 _26090_ (.Y(_07710_),
    .A(net2939),
    .B(net4576));
 sg13g2_o21ai_1 _26091_ (.B1(_07710_),
    .Y(_02745_),
    .A1(net5176),
    .A2(_07709_));
 sg13g2_mux2_1 _26092_ (.A0(net5162),
    .A1(net6119),
    .S(net4576),
    .X(_02746_));
 sg13g2_mux2_1 _26093_ (.A0(net5069),
    .A1(net4432),
    .S(net4576),
    .X(_02747_));
 sg13g2_mux2_1 _26094_ (.A0(net5047),
    .A1(net4233),
    .S(net4576),
    .X(_02748_));
 sg13g2_nand2_1 _26095_ (.Y(_07711_),
    .A(net4733),
    .B(_05075_));
 sg13g2_mux2_1 _26096_ (.A0(net5246),
    .A1(net4043),
    .S(_07711_),
    .X(_02749_));
 sg13g2_mux2_1 _26097_ (.A0(net5217),
    .A1(net6339),
    .S(net4614),
    .X(_02750_));
 sg13g2_mux2_1 _26098_ (.A0(net5117),
    .A1(net4443),
    .S(net4614),
    .X(_02751_));
 sg13g2_mux2_1 _26099_ (.A0(net5089),
    .A1(net6360),
    .S(net4614),
    .X(_02752_));
 sg13g2_nand2_1 _26100_ (.Y(_07712_),
    .A(net2915),
    .B(net4614));
 sg13g2_o21ai_1 _26101_ (.B1(_07712_),
    .Y(_02753_),
    .A1(net5174),
    .A2(net4614));
 sg13g2_mux2_1 _26102_ (.A0(net5160),
    .A1(net4431),
    .S(net4614),
    .X(_02754_));
 sg13g2_mux2_1 _26103_ (.A0(net5067),
    .A1(net6109),
    .S(net4614),
    .X(_02755_));
 sg13g2_mux2_1 _26104_ (.A0(net5043),
    .A1(net4450),
    .S(net4614),
    .X(_02756_));
 sg13g2_nand2_1 _26105_ (.Y(_07713_),
    .A(net4737),
    .B(_05075_));
 sg13g2_mux2_1 _26106_ (.A0(net5246),
    .A1(net4495),
    .S(_07713_),
    .X(_02757_));
 sg13g2_mux2_1 _26107_ (.A0(net5217),
    .A1(net4045),
    .S(net4613),
    .X(_02758_));
 sg13g2_mux2_1 _26108_ (.A0(net5120),
    .A1(net4151),
    .S(net4613),
    .X(_02759_));
 sg13g2_mux2_1 _26109_ (.A0(net5091),
    .A1(net4297),
    .S(net4613),
    .X(_02760_));
 sg13g2_nand2_1 _26110_ (.Y(_07714_),
    .A(net2944),
    .B(net4613));
 sg13g2_o21ai_1 _26111_ (.B1(_07714_),
    .Y(_02761_),
    .A1(net5174),
    .A2(net4613));
 sg13g2_mux2_1 _26112_ (.A0(net5160),
    .A1(net4011),
    .S(net4613),
    .X(_02762_));
 sg13g2_mux2_1 _26113_ (.A0(net5067),
    .A1(net4482),
    .S(net4613),
    .X(_02763_));
 sg13g2_mux2_1 _26114_ (.A0(net5043),
    .A1(net4106),
    .S(net4613),
    .X(_02764_));
 sg13g2_nor2b_1 _26115_ (.A(net4741),
    .B_N(_05075_),
    .Y(_07715_));
 sg13g2_nor2_1 _26116_ (.A(net3115),
    .B(net4612),
    .Y(_07716_));
 sg13g2_a21oi_1 _26117_ (.A1(net5263),
    .A2(net4612),
    .Y(_02765_),
    .B1(_07716_));
 sg13g2_nor2_1 _26118_ (.A(net3033),
    .B(net4611),
    .Y(_07717_));
 sg13g2_a21oi_1 _26119_ (.A1(net5237),
    .A2(net4611),
    .Y(_02766_),
    .B1(_07717_));
 sg13g2_nor2_1 _26120_ (.A(net3572),
    .B(net4611),
    .Y(_07718_));
 sg13g2_a21oi_1 _26121_ (.A1(net5134),
    .A2(net4611),
    .Y(_02767_),
    .B1(_07718_));
 sg13g2_nor2_1 _26122_ (.A(net3963),
    .B(net4611),
    .Y(_07719_));
 sg13g2_a21oi_1 _26123_ (.A1(net5106),
    .A2(net4611),
    .Y(_02768_),
    .B1(_07719_));
 sg13g2_mux2_1 _26124_ (.A0(net3330),
    .A1(net5186),
    .S(net4611),
    .X(_02769_));
 sg13g2_nor2_1 _26125_ (.A(net3447),
    .B(net4612),
    .Y(_07720_));
 sg13g2_a21oi_1 _26126_ (.A1(net5149),
    .A2(net4612),
    .Y(_02770_),
    .B1(_07720_));
 sg13g2_nor2_1 _26127_ (.A(net3063),
    .B(net4612),
    .Y(_07721_));
 sg13g2_a21oi_1 _26128_ (.A1(net5080),
    .A2(net4612),
    .Y(_02771_),
    .B1(_07721_));
 sg13g2_nor2_1 _26129_ (.A(net3994),
    .B(net4612),
    .Y(_07722_));
 sg13g2_a21oi_1 _26130_ (.A1(net5058),
    .A2(net4611),
    .Y(_02772_),
    .B1(_07722_));
 sg13g2_nand2_1 _26131_ (.Y(_07723_),
    .A(net4748),
    .B(_05075_));
 sg13g2_mux2_1 _26132_ (.A0(net5246),
    .A1(net6069),
    .S(_07723_),
    .X(_02773_));
 sg13g2_mux2_1 _26133_ (.A0(net5217),
    .A1(net4254),
    .S(net4610),
    .X(_02774_));
 sg13g2_mux2_1 _26134_ (.A0(net5120),
    .A1(net4343),
    .S(net4610),
    .X(_02775_));
 sg13g2_mux2_1 _26135_ (.A0(net5089),
    .A1(net6426),
    .S(net4610),
    .X(_02776_));
 sg13g2_nand2_1 _26136_ (.Y(_07724_),
    .A(net2960),
    .B(net4610));
 sg13g2_o21ai_1 _26137_ (.B1(_07724_),
    .Y(_02777_),
    .A1(net5174),
    .A2(net4610));
 sg13g2_mux2_1 _26138_ (.A0(net5160),
    .A1(net6235),
    .S(net4610),
    .X(_02778_));
 sg13g2_mux2_1 _26139_ (.A0(net5067),
    .A1(net4536),
    .S(net4610),
    .X(_02779_));
 sg13g2_mux2_1 _26140_ (.A0(net5043),
    .A1(net6128),
    .S(net4610),
    .X(_02780_));
 sg13g2_nand2_1 _26141_ (.Y(_07725_),
    .A(_03059_),
    .B(net4740));
 sg13g2_mux2_1 _26142_ (.A0(net5258),
    .A1(net4086),
    .S(net4609),
    .X(_02781_));
 sg13g2_mux2_1 _26143_ (.A0(net5231),
    .A1(net4097),
    .S(net4609),
    .X(_02782_));
 sg13g2_mux2_1 _26144_ (.A0(net5128),
    .A1(net4409),
    .S(net4609),
    .X(_02783_));
 sg13g2_mux2_1 _26145_ (.A0(net5100),
    .A1(net6222),
    .S(net4609),
    .X(_02784_));
 sg13g2_nand2_1 _26146_ (.Y(_07726_),
    .A(net2922),
    .B(net4609));
 sg13g2_o21ai_1 _26147_ (.B1(_07726_),
    .Y(_02785_),
    .A1(net5183),
    .A2(net4609));
 sg13g2_mux2_1 _26148_ (.A0(net5170),
    .A1(net6148),
    .S(net4609),
    .X(_02786_));
 sg13g2_mux2_1 _26149_ (.A0(net5076),
    .A1(net4240),
    .S(_07725_),
    .X(_02787_));
 sg13g2_mux2_1 _26150_ (.A0(net5053),
    .A1(net6572),
    .S(net4609),
    .X(_02788_));
 sg13g2_nand2_1 _26151_ (.Y(_07727_),
    .A(_03059_),
    .B(net4735));
 sg13g2_mux2_1 _26152_ (.A0(net5258),
    .A1(net4118),
    .S(net4608),
    .X(_02789_));
 sg13g2_mux2_1 _26153_ (.A0(net5231),
    .A1(net6205),
    .S(net4608),
    .X(_02790_));
 sg13g2_mux2_1 _26154_ (.A0(net5128),
    .A1(net4190),
    .S(net4608),
    .X(_02791_));
 sg13g2_mux2_1 _26155_ (.A0(net5100),
    .A1(net6086),
    .S(net4608),
    .X(_02792_));
 sg13g2_nand2_1 _26156_ (.Y(_07728_),
    .A(net2943),
    .B(net4608));
 sg13g2_o21ai_1 _26157_ (.B1(_07728_),
    .Y(_02793_),
    .A1(net5183),
    .A2(net4608));
 sg13g2_mux2_1 _26158_ (.A0(net5170),
    .A1(net6427),
    .S(net4608),
    .X(_02794_));
 sg13g2_mux2_1 _26159_ (.A0(net5076),
    .A1(net6665),
    .S(net4608),
    .X(_02795_));
 sg13g2_mux2_1 _26160_ (.A0(net5053),
    .A1(net4260),
    .S(_07727_),
    .X(_02796_));
 sg13g2_nor2_1 _26161_ (.A(net4744),
    .B(_03060_),
    .Y(_07729_));
 sg13g2_nor2_1 _26162_ (.A(net6179),
    .B(net4607),
    .Y(_07730_));
 sg13g2_a21oi_1 _26163_ (.A1(net5267),
    .A2(net4607),
    .Y(_02797_),
    .B1(_07730_));
 sg13g2_nor2_1 _26164_ (.A(net3111),
    .B(net4606),
    .Y(_07731_));
 sg13g2_a21oi_1 _26165_ (.A1(net5242),
    .A2(net4606),
    .Y(_02798_),
    .B1(_07731_));
 sg13g2_nor2_1 _26166_ (.A(net6154),
    .B(net4607),
    .Y(_07732_));
 sg13g2_a21oi_1 _26167_ (.A1(net5138),
    .A2(net4606),
    .Y(_02799_),
    .B1(_07732_));
 sg13g2_nor2_1 _26168_ (.A(net3046),
    .B(net4606),
    .Y(_07733_));
 sg13g2_a21oi_1 _26169_ (.A1(net5110),
    .A2(net4606),
    .Y(_02800_),
    .B1(_07733_));
 sg13g2_mux2_1 _26170_ (.A0(net3496),
    .A1(net5195),
    .S(net4607),
    .X(_02801_));
 sg13g2_nor2_1 _26171_ (.A(net3397),
    .B(net4606),
    .Y(_07734_));
 sg13g2_a21oi_1 _26172_ (.A1(net5154),
    .A2(net4606),
    .Y(_02802_),
    .B1(_07734_));
 sg13g2_nor2_1 _26173_ (.A(net3744),
    .B(net4607),
    .Y(_07735_));
 sg13g2_a21oi_1 _26174_ (.A1(net5083),
    .A2(net4607),
    .Y(_02803_),
    .B1(_07735_));
 sg13g2_nor2_1 _26175_ (.A(net3027),
    .B(net4607),
    .Y(_07736_));
 sg13g2_a21oi_1 _26176_ (.A1(net5061),
    .A2(net4606),
    .Y(_02804_),
    .B1(_07736_));
 sg13g2_nand2_1 _26177_ (.Y(_07737_),
    .A(net4746),
    .B(_03059_));
 sg13g2_mux2_1 _26178_ (.A0(net5258),
    .A1(net6120),
    .S(net4605),
    .X(_02805_));
 sg13g2_mux2_1 _26179_ (.A0(net5231),
    .A1(net6343),
    .S(net4605),
    .X(_02806_));
 sg13g2_mux2_1 _26180_ (.A0(net5128),
    .A1(net6160),
    .S(net4605),
    .X(_02807_));
 sg13g2_mux2_1 _26181_ (.A0(net5100),
    .A1(net6470),
    .S(net4605),
    .X(_02808_));
 sg13g2_nand2_1 _26182_ (.Y(_07738_),
    .A(net2952),
    .B(net4605));
 sg13g2_o21ai_1 _26183_ (.B1(_07738_),
    .Y(_02809_),
    .A1(net5183),
    .A2(net4605));
 sg13g2_mux2_1 _26184_ (.A0(net5170),
    .A1(net4540),
    .S(net4605),
    .X(_02810_));
 sg13g2_mux2_1 _26185_ (.A0(net5076),
    .A1(net6266),
    .S(_07737_),
    .X(_02811_));
 sg13g2_mux2_1 _26186_ (.A0(net5053),
    .A1(net6519),
    .S(net4605),
    .X(_02812_));
 sg13g2_nand2_1 _26187_ (.Y(_07739_),
    .A(_03059_),
    .B(net4734));
 sg13g2_mux2_1 _26188_ (.A0(net5256),
    .A1(net6095),
    .S(net4604),
    .X(_02813_));
 sg13g2_mux2_1 _26189_ (.A0(net5231),
    .A1(net6063),
    .S(net4604),
    .X(_02814_));
 sg13g2_mux2_1 _26190_ (.A0(net5128),
    .A1(net4272),
    .S(net4604),
    .X(_02815_));
 sg13g2_mux2_1 _26191_ (.A0(net5100),
    .A1(net4139),
    .S(net4604),
    .X(_02816_));
 sg13g2_nand2_1 _26192_ (.Y(_07740_),
    .A(net2926),
    .B(net4604));
 sg13g2_o21ai_1 _26193_ (.B1(_07740_),
    .Y(_02817_),
    .A1(net5183),
    .A2(_07739_));
 sg13g2_mux2_1 _26194_ (.A0(net5171),
    .A1(net4067),
    .S(net4604),
    .X(_02818_));
 sg13g2_mux2_1 _26195_ (.A0(net5075),
    .A1(net6332),
    .S(net4604),
    .X(_02819_));
 sg13g2_mux2_1 _26196_ (.A0(net5054),
    .A1(net4452),
    .S(net4604),
    .X(_02820_));
 sg13g2_nand2_1 _26197_ (.Y(_07741_),
    .A(_03158_),
    .B(net4733));
 sg13g2_mux2_1 _26198_ (.A0(net5251),
    .A1(net4145),
    .S(net4603),
    .X(_02821_));
 sg13g2_mux2_1 _26199_ (.A0(net5223),
    .A1(net4076),
    .S(net4603),
    .X(_02822_));
 sg13g2_mux2_1 _26200_ (.A0(net5118),
    .A1(net4129),
    .S(net4603),
    .X(_02823_));
 sg13g2_mux2_1 _26201_ (.A0(net5093),
    .A1(net6351),
    .S(net4603),
    .X(_02824_));
 sg13g2_nand2_1 _26202_ (.Y(_07742_),
    .A(net2949),
    .B(_07741_));
 sg13g2_o21ai_1 _26203_ (.B1(_07742_),
    .Y(_02825_),
    .A1(net5176),
    .A2(net4603));
 sg13g2_mux2_1 _26204_ (.A0(net5163),
    .A1(net4362),
    .S(net4603),
    .X(_02826_));
 sg13g2_mux2_1 _26205_ (.A0(net5069),
    .A1(net4124),
    .S(net4603),
    .X(_02827_));
 sg13g2_mux2_1 _26206_ (.A0(net5045),
    .A1(net4385),
    .S(net4603),
    .X(_02828_));
 sg13g2_nor3_1 _26207_ (.A(_03008_),
    .B(_03166_),
    .C(_04814_),
    .Y(_07743_));
 sg13g2_nor2_1 _26208_ (.A(net3713),
    .B(net4602),
    .Y(_07744_));
 sg13g2_a21oi_1 _26209_ (.A1(net5262),
    .A2(net4602),
    .Y(_02829_),
    .B1(_07744_));
 sg13g2_nor2_1 _26210_ (.A(net2987),
    .B(net4602),
    .Y(_07745_));
 sg13g2_a21oi_1 _26211_ (.A1(net5235),
    .A2(net4602),
    .Y(_02830_),
    .B1(_07745_));
 sg13g2_nor2_1 _26212_ (.A(net3421),
    .B(net4601),
    .Y(_07746_));
 sg13g2_a21oi_1 _26213_ (.A1(net5132),
    .A2(net4601),
    .Y(_02831_),
    .B1(_07746_));
 sg13g2_nor2_1 _26214_ (.A(net4026),
    .B(net4602),
    .Y(_07747_));
 sg13g2_a21oi_1 _26215_ (.A1(net5104),
    .A2(net4602),
    .Y(_02832_),
    .B1(_07747_));
 sg13g2_mux2_1 _26216_ (.A0(net3322),
    .A1(net5189),
    .S(net4602),
    .X(_02833_));
 sg13g2_nor2_1 _26217_ (.A(net3081),
    .B(net4601),
    .Y(_07748_));
 sg13g2_a21oi_1 _26218_ (.A1(net5147),
    .A2(net4601),
    .Y(_02834_),
    .B1(_07748_));
 sg13g2_nor2_1 _26219_ (.A(net3101),
    .B(net4601),
    .Y(_07749_));
 sg13g2_a21oi_1 _26220_ (.A1(net5079),
    .A2(net4601),
    .Y(_02835_),
    .B1(_07749_));
 sg13g2_nor2_1 _26221_ (.A(net3015),
    .B(net4601),
    .Y(_07750_));
 sg13g2_a21oi_1 _26222_ (.A1(net5056),
    .A2(net4601),
    .Y(_02836_),
    .B1(_07750_));
 sg13g2_nor2b_1 _26223_ (.A(net4743),
    .B_N(net4763),
    .Y(_07751_));
 sg13g2_nor2_1 _26224_ (.A(net3824),
    .B(net4600),
    .Y(_07752_));
 sg13g2_a21oi_1 _26225_ (.A1(net5261),
    .A2(net4600),
    .Y(_02837_),
    .B1(_07752_));
 sg13g2_nor2_1 _26226_ (.A(net3068),
    .B(net4599),
    .Y(_07753_));
 sg13g2_a21oi_1 _26227_ (.A1(net5235),
    .A2(net4599),
    .Y(_02838_),
    .B1(_07753_));
 sg13g2_nor2_1 _26228_ (.A(net3340),
    .B(net4599),
    .Y(_07754_));
 sg13g2_a21oi_1 _26229_ (.A1(net5132),
    .A2(net4599),
    .Y(_02839_),
    .B1(_07754_));
 sg13g2_nor2_1 _26230_ (.A(net3928),
    .B(net4600),
    .Y(_07755_));
 sg13g2_a21oi_1 _26231_ (.A1(net5104),
    .A2(net4600),
    .Y(_02840_),
    .B1(_07755_));
 sg13g2_mux2_1 _26232_ (.A0(net3243),
    .A1(net5188),
    .S(net4600),
    .X(_02841_));
 sg13g2_nor2_1 _26233_ (.A(net4218),
    .B(net4599),
    .Y(_07756_));
 sg13g2_a21oi_1 _26234_ (.A1(net5147),
    .A2(net4599),
    .Y(_02842_),
    .B1(_07756_));
 sg13g2_nor2_1 _26235_ (.A(net3456),
    .B(net4599),
    .Y(_07757_));
 sg13g2_a21oi_1 _26236_ (.A1(net5078),
    .A2(net4599),
    .Y(_02843_),
    .B1(_07757_));
 sg13g2_nor2_1 _26237_ (.A(net4005),
    .B(net4600),
    .Y(_07758_));
 sg13g2_a21oi_1 _26238_ (.A1(net5056),
    .A2(net4600),
    .Y(_02844_),
    .B1(_07758_));
 sg13g2_nand2_1 _26239_ (.Y(_07759_),
    .A(net4763),
    .B(net4735));
 sg13g2_mux2_1 _26240_ (.A0(net5254),
    .A1(net4518),
    .S(net4598),
    .X(_02845_));
 sg13g2_mux2_1 _26241_ (.A0(net5223),
    .A1(net4207),
    .S(net4598),
    .X(_02846_));
 sg13g2_mux2_1 _26242_ (.A0(net5118),
    .A1(net4081),
    .S(net4598),
    .X(_02847_));
 sg13g2_mux2_1 _26243_ (.A0(net5093),
    .A1(net4526),
    .S(net4598),
    .X(_02848_));
 sg13g2_nand2_1 _26244_ (.Y(_07760_),
    .A(net2959),
    .B(_07759_));
 sg13g2_o21ai_1 _26245_ (.B1(_07760_),
    .Y(_02849_),
    .A1(net5176),
    .A2(net4598));
 sg13g2_mux2_1 _26246_ (.A0(net5162),
    .A1(net6347),
    .S(net4598),
    .X(_02850_));
 sg13g2_mux2_1 _26247_ (.A0(net5070),
    .A1(net6105),
    .S(net4598),
    .X(_02851_));
 sg13g2_mux2_1 _26248_ (.A0(net5046),
    .A1(net6945),
    .S(net4598),
    .X(_02852_));
 sg13g2_nor2_1 _26249_ (.A(net5979),
    .B(_08563_),
    .Y(_02853_));
 sg13g2_nor2_1 _26250_ (.A(net5979),
    .B(_08554_),
    .Y(_02854_));
 sg13g2_nor2_1 _26251_ (.A(net5982),
    .B(net5032),
    .Y(_02855_));
 sg13g2_nor2_1 _26252_ (.A(net5982),
    .B(net5026),
    .Y(_02857_));
 sg13g2_nor2_1 _26253_ (.A(net5981),
    .B(net4877),
    .Y(_02858_));
 sg13g2_nor2_1 _26254_ (.A(net5982),
    .B(net5024),
    .Y(_02859_));
 sg13g2_and2_1 _26255_ (.A(net5998),
    .B(_10417_),
    .X(_02860_));
 sg13g2_nor2_1 _26256_ (.A(net5979),
    .B(_10398_),
    .Y(_02861_));
 sg13g2_nor2_1 _26257_ (.A(net5979),
    .B(_10404_),
    .Y(_02862_));
 sg13g2_and2_1 _26258_ (.A(net5998),
    .B(_10390_),
    .X(_02863_));
 sg13g2_and2_1 _26259_ (.A(net5998),
    .B(_10412_),
    .X(_02864_));
 sg13g2_nor2_1 _26260_ (.A(net5979),
    .B(net4781),
    .Y(_02865_));
 sg13g2_nand2_1 _26261_ (.Y(_07761_),
    .A(net4740),
    .B(net4763));
 sg13g2_mux2_1 _26262_ (.A0(net5253),
    .A1(net4200),
    .S(net4597),
    .X(_02866_));
 sg13g2_mux2_1 _26263_ (.A0(net5223),
    .A1(net4268),
    .S(net4597),
    .X(_02867_));
 sg13g2_mux2_1 _26264_ (.A0(net5118),
    .A1(net6083),
    .S(net4597),
    .X(_02868_));
 sg13g2_mux2_1 _26265_ (.A0(net5095),
    .A1(net6588),
    .S(net4597),
    .X(_02869_));
 sg13g2_nand2_1 _26266_ (.Y(_07762_),
    .A(net2937),
    .B(_07761_));
 sg13g2_o21ai_1 _26267_ (.B1(_07762_),
    .Y(_02870_),
    .A1(net5176),
    .A2(net4597));
 sg13g2_mux2_1 _26268_ (.A0(net5162),
    .A1(net6694),
    .S(net4597),
    .X(_02871_));
 sg13g2_mux2_1 _26269_ (.A0(net5070),
    .A1(net6075),
    .S(net4597),
    .X(_02872_));
 sg13g2_mux2_1 _26270_ (.A0(net5046),
    .A1(net4162),
    .S(net4597),
    .X(_02873_));
 sg13g2_nand2_1 _26271_ (.Y(_07763_),
    .A(net4748),
    .B(_03165_));
 sg13g2_mux2_1 _26272_ (.A0(net5244),
    .A1(net6227),
    .S(net4575),
    .X(_02874_));
 sg13g2_mux2_1 _26273_ (.A0(net5219),
    .A1(net6636),
    .S(net4575),
    .X(_02875_));
 sg13g2_mux2_1 _26274_ (.A0(net5115),
    .A1(net6354),
    .S(net4575),
    .X(_02876_));
 sg13g2_mux2_1 _26275_ (.A0(net5090),
    .A1(net4395),
    .S(net4575),
    .X(_02877_));
 sg13g2_nand2_1 _26276_ (.Y(_07764_),
    .A(net2979),
    .B(_07763_));
 sg13g2_o21ai_1 _26277_ (.B1(_07764_),
    .Y(_02878_),
    .A1(net5175),
    .A2(net4575));
 sg13g2_mux2_1 _26278_ (.A0(net5157),
    .A1(net6446),
    .S(net4575),
    .X(_02879_));
 sg13g2_mux2_1 _26279_ (.A0(net5065),
    .A1(net4418),
    .S(net4575),
    .X(_02880_));
 sg13g2_mux2_1 _26280_ (.A0(net5042),
    .A1(net6108),
    .S(net4575),
    .X(_02881_));
 sg13g2_nor2b_1 _26281_ (.A(net4741),
    .B_N(_04811_),
    .Y(_07765_));
 sg13g2_nor2_1 _26282_ (.A(net3979),
    .B(net4595),
    .Y(_07766_));
 sg13g2_a21oi_1 _26283_ (.A1(net5261),
    .A2(net4595),
    .Y(_02882_),
    .B1(_07766_));
 sg13g2_nor2_1 _26284_ (.A(net3653),
    .B(net4596),
    .Y(_07767_));
 sg13g2_a21oi_1 _26285_ (.A1(net5242),
    .A2(net4596),
    .Y(_02883_),
    .B1(_07767_));
 sg13g2_nor2_1 _26286_ (.A(net3633),
    .B(net4595),
    .Y(_07768_));
 sg13g2_a21oi_1 _26287_ (.A1(net5133),
    .A2(net4595),
    .Y(_02884_),
    .B1(_07768_));
 sg13g2_nor2_1 _26288_ (.A(net4049),
    .B(net4595),
    .Y(_07769_));
 sg13g2_a21oi_1 _26289_ (.A1(net5110),
    .A2(net4595),
    .Y(_02885_),
    .B1(_07769_));
 sg13g2_mux2_1 _26290_ (.A0(net3568),
    .A1(net5195),
    .S(net4596),
    .X(_02886_));
 sg13g2_nor2_1 _26291_ (.A(net3090),
    .B(net4596),
    .Y(_07770_));
 sg13g2_a21oi_1 _26292_ (.A1(net5154),
    .A2(net4596),
    .Y(_02887_),
    .B1(_07770_));
 sg13g2_nor2_1 _26293_ (.A(net3781),
    .B(net4595),
    .Y(_07771_));
 sg13g2_a21oi_1 _26294_ (.A1(net5087),
    .A2(net4595),
    .Y(_02888_),
    .B1(_07771_));
 sg13g2_nor2_1 _26295_ (.A(net3859),
    .B(net4596),
    .Y(_07772_));
 sg13g2_a21oi_1 _26296_ (.A1(net5061),
    .A2(net4596),
    .Y(_02889_),
    .B1(_07772_));
 sg13g2_nor3_1 _26297_ (.A(net5038),
    .B(net4741),
    .C(_03164_),
    .Y(_07773_));
 sg13g2_nor2_1 _26298_ (.A(net3094),
    .B(net4593),
    .Y(_07774_));
 sg13g2_a21oi_1 _26299_ (.A1(net5260),
    .A2(net4593),
    .Y(_02890_),
    .B1(_07774_));
 sg13g2_nor2_1 _26300_ (.A(net3406),
    .B(net4593),
    .Y(_07775_));
 sg13g2_a21oi_1 _26301_ (.A1(net5234),
    .A2(net4593),
    .Y(_02891_),
    .B1(_07775_));
 sg13g2_nor2_1 _26302_ (.A(net3045),
    .B(net4594),
    .Y(_07776_));
 sg13g2_a21oi_1 _26303_ (.A1(net5131),
    .A2(net4593),
    .Y(_02892_),
    .B1(_07776_));
 sg13g2_nor2_1 _26304_ (.A(net3077),
    .B(net4593),
    .Y(_07777_));
 sg13g2_a21oi_1 _26305_ (.A1(net5103),
    .A2(net4593),
    .Y(_02893_),
    .B1(_07777_));
 sg13g2_mux2_1 _26306_ (.A0(net3331),
    .A1(net5188),
    .S(net4594),
    .X(_02894_));
 sg13g2_nor2_1 _26307_ (.A(net3671),
    .B(net4593),
    .Y(_07778_));
 sg13g2_a21oi_1 _26308_ (.A1(net5146),
    .A2(net4594),
    .Y(_02895_),
    .B1(_07778_));
 sg13g2_nor2_1 _26309_ (.A(net3093),
    .B(net4594),
    .Y(_07779_));
 sg13g2_a21oi_1 _26310_ (.A1(net5078),
    .A2(net4594),
    .Y(_02896_),
    .B1(_07779_));
 sg13g2_nor2_1 _26311_ (.A(net3579),
    .B(net4594),
    .Y(_07780_));
 sg13g2_a21oi_1 _26312_ (.A1(net5055),
    .A2(net4594),
    .Y(_02897_),
    .B1(_07780_));
 sg13g2_nand2_1 _26313_ (.Y(_07781_),
    .A(_04811_),
    .B(net4733));
 sg13g2_mux2_1 _26314_ (.A0(net5252),
    .A1(net6765),
    .S(net4592),
    .X(_02898_));
 sg13g2_mux2_1 _26315_ (.A0(net5224),
    .A1(net6697),
    .S(net4592),
    .X(_02899_));
 sg13g2_mux2_1 _26316_ (.A0(net5122),
    .A1(net6340),
    .S(net4592),
    .X(_02900_));
 sg13g2_mux2_1 _26317_ (.A0(net5094),
    .A1(net4123),
    .S(net4592),
    .X(_02901_));
 sg13g2_nand2_1 _26318_ (.Y(_07782_),
    .A(net2916),
    .B(net4592));
 sg13g2_o21ai_1 _26319_ (.B1(_07782_),
    .Y(_02902_),
    .A1(net5177),
    .A2(net4592));
 sg13g2_mux2_1 _26320_ (.A0(net5170),
    .A1(net4353),
    .S(net4592),
    .X(_02903_));
 sg13g2_mux2_1 _26321_ (.A0(net5075),
    .A1(net6126),
    .S(net4592),
    .X(_02904_));
 sg13g2_mux2_1 _26322_ (.A0(net5053),
    .A1(net6181),
    .S(_07781_),
    .X(_02905_));
 sg13g2_nand2_1 _26323_ (.Y(_07783_),
    .A(net4737),
    .B(_04811_));
 sg13g2_mux2_1 _26324_ (.A0(net5252),
    .A1(net4219),
    .S(net4591),
    .X(_02906_));
 sg13g2_mux2_1 _26325_ (.A0(net5231),
    .A1(net4013),
    .S(net4591),
    .X(_02907_));
 sg13g2_mux2_1 _26326_ (.A0(net5122),
    .A1(net4342),
    .S(net4591),
    .X(_02908_));
 sg13g2_mux2_1 _26327_ (.A0(net5095),
    .A1(net4070),
    .S(net4591),
    .X(_02909_));
 sg13g2_nand2_1 _26328_ (.Y(_07784_),
    .A(net2932),
    .B(net4591));
 sg13g2_o21ai_1 _26329_ (.B1(_07784_),
    .Y(_02910_),
    .A1(net5183),
    .A2(_07783_));
 sg13g2_mux2_1 _26330_ (.A0(net5170),
    .A1(net4167),
    .S(net4591),
    .X(_02911_));
 sg13g2_mux2_1 _26331_ (.A0(net5075),
    .A1(net4197),
    .S(net4591),
    .X(_02912_));
 sg13g2_mux2_1 _26332_ (.A0(net5053),
    .A1(net4242),
    .S(net4591),
    .X(_02913_));
 sg13g2_nand2_1 _26333_ (.Y(_07785_),
    .A(net5537),
    .B(_10445_));
 sg13g2_nand2_1 _26334_ (.Y(_07786_),
    .A(_07640_),
    .B(_07785_));
 sg13g2_nand2_1 _26335_ (.Y(_07787_),
    .A(\flash_rom.fsm_state[1] ),
    .B(\flash_rom.fsm_state[0] ));
 sg13g2_o21ai_1 _26336_ (.B1(_07642_),
    .Y(_07788_),
    .A1(net5567),
    .A2(_07787_));
 sg13g2_a21oi_1 _26337_ (.A1(_07921_),
    .A2(_08077_),
    .Y(_07789_),
    .B1(\flash_rom.fsm_state[1] ));
 sg13g2_nor4_2 _26338_ (.A(_00137_),
    .B(_08492_),
    .C(_07788_),
    .Y(_07790_),
    .D(_07789_));
 sg13g2_nor2_1 _26339_ (.A(net5537),
    .B(_07639_),
    .Y(_07791_));
 sg13g2_nor3_2 _26340_ (.A(\flash_rom.spi_clk_out ),
    .B(net5537),
    .C(_07639_),
    .Y(_07792_));
 sg13g2_nor2_1 _26341_ (.A(_07639_),
    .B(_07792_),
    .Y(_07793_));
 sg13g2_nor3_2 _26342_ (.A(_07786_),
    .B(_07790_),
    .C(_07792_),
    .Y(_07794_));
 sg13g2_nor2_1 _26343_ (.A(net7174),
    .B(_07794_),
    .Y(_07795_));
 sg13g2_nand2_1 _26344_ (.Y(_07796_),
    .A(\flash_rom.spi_clk_out ),
    .B(_07791_));
 sg13g2_or2_1 _26345_ (.X(_07797_),
    .B(_07796_),
    .A(_07790_));
 sg13g2_nor2_1 _26346_ (.A(_07922_),
    .B(_07797_),
    .Y(_07798_));
 sg13g2_nor3_1 _26347_ (.A(_07638_),
    .B(_07795_),
    .C(_07798_),
    .Y(_02914_));
 sg13g2_nor2_1 _26348_ (.A(net7206),
    .B(_07794_),
    .Y(_07799_));
 sg13g2_xnor2_1 _26349_ (.Y(_07800_),
    .A(net7206),
    .B(net7174));
 sg13g2_a21oi_1 _26350_ (.A1(_07788_),
    .A2(_07800_),
    .Y(_07801_),
    .B1(_07797_));
 sg13g2_nor3_1 _26351_ (.A(net4572),
    .B(_07799_),
    .C(_07801_),
    .Y(_02915_));
 sg13g2_nand3_1 _26352_ (.B(_10352_),
    .C(_07642_),
    .A(_00102_),
    .Y(_07802_));
 sg13g2_nand3b_1 _26353_ (.B(_07802_),
    .C(_10354_),
    .Y(_07803_),
    .A_N(_07797_));
 sg13g2_o21ai_1 _26354_ (.B1(_07803_),
    .Y(_07804_),
    .A1(net7199),
    .A2(_07794_));
 sg13g2_nor2_1 _26355_ (.A(net4572),
    .B(net7200),
    .Y(_02916_));
 sg13g2_or2_1 _26356_ (.X(_07805_),
    .B(_07796_),
    .A(_07642_));
 sg13g2_a21oi_1 _26357_ (.A1(\flash_rom.stall_read ),
    .A2(_07639_),
    .Y(_07806_),
    .B1(_07792_));
 sg13g2_or2_1 _26358_ (.X(_07807_),
    .B(_07643_),
    .A(\flash_rom.stall_read ));
 sg13g2_and4_2 _26359_ (.A(_07785_),
    .B(_07805_),
    .C(_07806_),
    .D(_07807_),
    .X(_07808_));
 sg13g2_nand2_1 _26360_ (.Y(_07809_),
    .A(net7234),
    .B(_07641_));
 sg13g2_and3_1 _26361_ (.X(_07810_),
    .A(_07791_),
    .B(_07808_),
    .C(_07809_));
 sg13g2_nor2_1 _26362_ (.A(net2899),
    .B(_07808_),
    .Y(_07811_));
 sg13g2_nor3_1 _26363_ (.A(net4572),
    .B(_07810_),
    .C(_07811_),
    .Y(_02917_));
 sg13g2_nor2_1 _26364_ (.A(net7246),
    .B(_07808_),
    .Y(_07812_));
 sg13g2_nor2_1 _26365_ (.A(_10351_),
    .B(_10352_),
    .Y(_07813_));
 sg13g2_a21oi_1 _26366_ (.A1(_07808_),
    .A2(_07813_),
    .Y(_07814_),
    .B1(_07638_));
 sg13g2_nor2b_1 _26367_ (.A(_07812_),
    .B_N(_07814_),
    .Y(_02918_));
 sg13g2_o21ai_1 _26368_ (.B1(_07640_),
    .Y(_07815_),
    .A1(net5567),
    .A2(_07787_));
 sg13g2_a21oi_1 _26369_ (.A1(net5567),
    .A2(_07787_),
    .Y(_07816_),
    .B1(_07815_));
 sg13g2_nand2_1 _26370_ (.Y(_07817_),
    .A(_07808_),
    .B(_07816_));
 sg13g2_o21ai_1 _26371_ (.B1(_07817_),
    .Y(_07818_),
    .A1(net5567),
    .A2(_07808_));
 sg13g2_nor2_1 _26372_ (.A(net4572),
    .B(_07818_),
    .Y(_02919_));
 sg13g2_nor2_1 _26373_ (.A(_00137_),
    .B(_07641_),
    .Y(_07819_));
 sg13g2_mux2_1 _26374_ (.A0(net7057),
    .A1(net8),
    .S(net5399),
    .X(_02920_));
 sg13g2_mux2_1 _26375_ (.A0(net4229),
    .A1(net9),
    .S(net5399),
    .X(_02921_));
 sg13g2_mux2_1 _26376_ (.A0(net7045),
    .A1(net10),
    .S(net5399),
    .X(_02922_));
 sg13g2_mux2_1 _26377_ (.A0(net3958),
    .A1(net11),
    .S(net5399),
    .X(_02923_));
 sg13g2_mux2_1 _26378_ (.A0(net3172),
    .A1(\atari2600.rom_data[0] ),
    .S(net5399),
    .X(_02924_));
 sg13g2_mux2_1 _26379_ (.A0(net3001),
    .A1(\atari2600.rom_data[1] ),
    .S(net5399),
    .X(_02925_));
 sg13g2_mux2_1 _26380_ (.A0(net3965),
    .A1(\atari2600.rom_data[2] ),
    .S(net5399),
    .X(_02926_));
 sg13g2_mux2_1 _26381_ (.A0(net3354),
    .A1(\atari2600.rom_data[3] ),
    .S(net5399),
    .X(_02927_));
 sg13g2_a22oi_1 _26382_ (.Y(_07820_),
    .B1(_07791_),
    .B2(net7193),
    .A2(_07786_),
    .A1(\flash_rom.spi_clk_out ));
 sg13g2_nand2b_1 _26383_ (.Y(_02928_),
    .B(net7194),
    .A_N(net4572));
 sg13g2_o21ai_1 _26384_ (.B1(_10350_),
    .Y(_07821_),
    .A1(\flash_rom.fsm_state[1] ),
    .A2(_00138_));
 sg13g2_a21oi_1 _26385_ (.A1(_00102_),
    .A2(net5428),
    .Y(_07822_),
    .B1(_07819_));
 sg13g2_o21ai_1 _26386_ (.B1(_07822_),
    .Y(_07823_),
    .A1(_07796_),
    .A2(_07821_));
 sg13g2_nand2_1 _26387_ (.Y(_07824_),
    .A(_07642_),
    .B(_07823_));
 sg13g2_nand4_1 _26388_ (.B(_07793_),
    .C(_07805_),
    .A(_07785_),
    .Y(_07825_),
    .D(_07824_));
 sg13g2_nor2b_1 _26389_ (.A(_07825_),
    .B_N(_10353_),
    .Y(_07826_));
 sg13g2_nor2b_1 _26390_ (.A(net2900),
    .B_N(_07826_),
    .Y(_07827_));
 sg13g2_nor2b_1 _26391_ (.A(net7081),
    .B_N(_07825_),
    .Y(_07828_));
 sg13g2_nor3_1 _26392_ (.A(net4572),
    .B(_07827_),
    .C(_07828_),
    .Y(_02929_));
 sg13g2_nor2b_1 _26393_ (.A(net7215),
    .B_N(_07825_),
    .Y(_07829_));
 sg13g2_nor3_1 _26394_ (.A(net4572),
    .B(_07826_),
    .C(_07829_),
    .Y(_02930_));
 sg13g2_and3_1 _26395_ (.X(_07830_),
    .A(_08583_),
    .B(_08636_),
    .C(_05408_));
 sg13g2_nand3_1 _26396_ (.B(_08636_),
    .C(_05408_),
    .A(_08583_),
    .Y(_07831_));
 sg13g2_o21ai_1 _26397_ (.B1(net6032),
    .Y(_07832_),
    .A1(_05409_),
    .A2(_07831_));
 sg13g2_a21oi_1 _26398_ (.A1(_07920_),
    .A2(_07831_),
    .Y(_02931_),
    .B1(_07832_));
 sg13g2_o21ai_1 _26399_ (.B1(net6032),
    .Y(_07833_),
    .A1(net7250),
    .A2(_07830_));
 sg13g2_a21oi_1 _26400_ (.A1(_08666_),
    .A2(_07830_),
    .Y(_02932_),
    .B1(_07833_));
 sg13g2_nor2_1 _26401_ (.A(net7104),
    .B(_07830_),
    .Y(_07834_));
 sg13g2_a21oi_1 _26402_ (.A1(_05414_),
    .A2(_07830_),
    .Y(_07835_),
    .B1(net5983));
 sg13g2_nor2b_1 _26403_ (.A(_07834_),
    .B_N(_07835_),
    .Y(_02933_));
 sg13g2_nand2_1 _26404_ (.Y(_07836_),
    .A(net4739),
    .B(_07104_));
 sg13g2_mux2_1 _26405_ (.A0(net5250),
    .A1(net6229),
    .S(_07836_),
    .X(_02934_));
 sg13g2_mux2_1 _26406_ (.A0(net5217),
    .A1(net4367),
    .S(net4590),
    .X(_02935_));
 sg13g2_mux2_1 _26407_ (.A0(net5117),
    .A1(net4402),
    .S(net4590),
    .X(_02936_));
 sg13g2_mux2_1 _26408_ (.A0(net5089),
    .A1(net4198),
    .S(net4590),
    .X(_02937_));
 sg13g2_nand2_1 _26409_ (.Y(_07837_),
    .A(net2946),
    .B(net4590));
 sg13g2_o21ai_1 _26410_ (.B1(_07837_),
    .Y(_02938_),
    .A1(net5173),
    .A2(net4590));
 sg13g2_mux2_1 _26411_ (.A0(net5161),
    .A1(net6610),
    .S(net4590),
    .X(_02939_));
 sg13g2_mux2_1 _26412_ (.A0(net5064),
    .A1(net4156),
    .S(net4590),
    .X(_02940_));
 sg13g2_mux2_1 _26413_ (.A0(net5040),
    .A1(net6189),
    .S(net4590),
    .X(_02941_));
 sg13g2_nand2_1 _26414_ (.Y(_07838_),
    .A(net4735),
    .B(_07104_));
 sg13g2_mux2_1 _26415_ (.A0(net5250),
    .A1(net4072),
    .S(net4589),
    .X(_02942_));
 sg13g2_mux2_1 _26416_ (.A0(net5217),
    .A1(net4018),
    .S(net4589),
    .X(_02943_));
 sg13g2_mux2_1 _26417_ (.A0(net5116),
    .A1(net4131),
    .S(net4589),
    .X(_02944_));
 sg13g2_mux2_1 _26418_ (.A0(net5090),
    .A1(net6410),
    .S(net4589),
    .X(_02945_));
 sg13g2_nand2_1 _26419_ (.Y(_07839_),
    .A(net2917),
    .B(net4589));
 sg13g2_o21ai_1 _26420_ (.B1(_07839_),
    .Y(_02946_),
    .A1(net5173),
    .A2(net4589));
 sg13g2_mux2_1 _26421_ (.A0(net5161),
    .A1(net4419),
    .S(net4589),
    .X(_02947_));
 sg13g2_mux2_1 _26422_ (.A0(net5065),
    .A1(net6369),
    .S(_07838_),
    .X(_02948_));
 sg13g2_mux2_1 _26423_ (.A0(net5040),
    .A1(net6050),
    .S(net4589),
    .X(_02949_));
 sg13g2_and2_1 _26424_ (.A(net4746),
    .B(_04813_),
    .X(_07840_));
 sg13g2_nor2_1 _26425_ (.A(net3743),
    .B(net4573),
    .Y(_07841_));
 sg13g2_a21oi_1 _26426_ (.A1(net5262),
    .A2(net4573),
    .Y(_02950_),
    .B1(_07841_));
 sg13g2_nor2_1 _26427_ (.A(net3289),
    .B(net4573),
    .Y(_07842_));
 sg13g2_a21oi_1 _26428_ (.A1(net5235),
    .A2(net4573),
    .Y(_02951_),
    .B1(_07842_));
 sg13g2_nor2_1 _26429_ (.A(net3006),
    .B(net4573),
    .Y(_07843_));
 sg13g2_a21oi_1 _26430_ (.A1(net5132),
    .A2(net4573),
    .Y(_02952_),
    .B1(_07843_));
 sg13g2_nor2_1 _26431_ (.A(net3915),
    .B(net4573),
    .Y(_07844_));
 sg13g2_a21oi_1 _26432_ (.A1(net5104),
    .A2(net4573),
    .Y(_02953_),
    .B1(_07844_));
 sg13g2_mux2_1 _26433_ (.A0(net3319),
    .A1(net5188),
    .S(net4574),
    .X(_02954_));
 sg13g2_nor2_1 _26434_ (.A(net3869),
    .B(net4574),
    .Y(_07845_));
 sg13g2_a21oi_1 _26435_ (.A1(net5147),
    .A2(net4574),
    .Y(_02955_),
    .B1(_07845_));
 sg13g2_nor2_1 _26436_ (.A(net3038),
    .B(net4574),
    .Y(_07846_));
 sg13g2_a21oi_1 _26437_ (.A1(net5078),
    .A2(net4574),
    .Y(_02956_),
    .B1(_07846_));
 sg13g2_nor2_1 _26438_ (.A(net3760),
    .B(net4574),
    .Y(_07847_));
 sg13g2_a21oi_1 _26439_ (.A1(net5056),
    .A2(net4574),
    .Y(_02957_),
    .B1(_07847_));
 sg13g2_nor2b_1 _26440_ (.A(net4741),
    .B_N(_05071_),
    .Y(_07848_));
 sg13g2_nor2_1 _26441_ (.A(net3657),
    .B(net4588),
    .Y(_07849_));
 sg13g2_a21oi_1 _26442_ (.A1(net5260),
    .A2(net4588),
    .Y(_02958_),
    .B1(_07849_));
 sg13g2_nor2_1 _26443_ (.A(net3007),
    .B(net4588),
    .Y(_07850_));
 sg13g2_a21oi_1 _26444_ (.A1(net5234),
    .A2(net4588),
    .Y(_02959_),
    .B1(_07850_));
 sg13g2_nor2_1 _26445_ (.A(net3525),
    .B(net4587),
    .Y(_07851_));
 sg13g2_a21oi_1 _26446_ (.A1(net5131),
    .A2(net4587),
    .Y(_02960_),
    .B1(_07851_));
 sg13g2_nor2_1 _26447_ (.A(net3404),
    .B(net4587),
    .Y(_07852_));
 sg13g2_a21oi_1 _26448_ (.A1(net5103),
    .A2(net4587),
    .Y(_02961_),
    .B1(_07852_));
 sg13g2_mux2_1 _26449_ (.A0(net3793),
    .A1(net5185),
    .S(net4588),
    .X(_02962_));
 sg13g2_nor2_1 _26450_ (.A(net3984),
    .B(net4587),
    .Y(_07853_));
 sg13g2_a21oi_1 _26451_ (.A1(net5146),
    .A2(net4587),
    .Y(_02963_),
    .B1(_07853_));
 sg13g2_nor2_1 _26452_ (.A(net3110),
    .B(net4588),
    .Y(_07854_));
 sg13g2_a21oi_1 _26453_ (.A1(net5078),
    .A2(net4588),
    .Y(_02964_),
    .B1(_07854_));
 sg13g2_nor2_1 _26454_ (.A(net3073),
    .B(net4587),
    .Y(_07855_));
 sg13g2_a21oi_1 _26455_ (.A1(net5055),
    .A2(net4587),
    .Y(_02965_),
    .B1(_07855_));
 sg13g2_nand2_1 _26456_ (.Y(_07856_),
    .A(net4737),
    .B(_05071_));
 sg13g2_mux2_1 _26457_ (.A0(net5245),
    .A1(net6442),
    .S(_07856_),
    .X(_02966_));
 sg13g2_mux2_1 _26458_ (.A0(net5218),
    .A1(net6090),
    .S(net4586),
    .X(_02967_));
 sg13g2_mux2_1 _26459_ (.A0(net5115),
    .A1(net6941),
    .S(net4586),
    .X(_02968_));
 sg13g2_mux2_1 _26460_ (.A0(net5088),
    .A1(net6196),
    .S(net4586),
    .X(_02969_));
 sg13g2_nand2_1 _26461_ (.Y(_07857_),
    .A(net2906),
    .B(net4586));
 sg13g2_o21ai_1 _26462_ (.B1(_07857_),
    .Y(_02970_),
    .A1(net5173),
    .A2(net4586));
 sg13g2_mux2_1 _26463_ (.A0(net5158),
    .A1(net6399),
    .S(net4586),
    .X(_02971_));
 sg13g2_mux2_1 _26464_ (.A0(net5064),
    .A1(net6598),
    .S(net4586),
    .X(_02972_));
 sg13g2_mux2_1 _26465_ (.A0(net5040),
    .A1(net4298),
    .S(net4586),
    .X(_02973_));
 sg13g2_nand2_1 _26466_ (.Y(_07858_),
    .A(net4733),
    .B(_05071_));
 sg13g2_mux2_1 _26467_ (.A0(net5245),
    .A1(net6686),
    .S(net4585),
    .X(_02974_));
 sg13g2_mux2_1 _26468_ (.A0(net5218),
    .A1(net4507),
    .S(net4585),
    .X(_02975_));
 sg13g2_mux2_1 _26469_ (.A0(net5115),
    .A1(net6828),
    .S(net4585),
    .X(_02976_));
 sg13g2_mux2_1 _26470_ (.A0(net5088),
    .A1(net6615),
    .S(net4585),
    .X(_02977_));
 sg13g2_nand2_1 _26471_ (.Y(_07859_),
    .A(net2945),
    .B(_07858_));
 sg13g2_o21ai_1 _26472_ (.B1(_07859_),
    .Y(_02978_),
    .A1(net5173),
    .A2(net4585));
 sg13g2_mux2_1 _26473_ (.A0(net5158),
    .A1(net6906),
    .S(net4585),
    .X(_02979_));
 sg13g2_mux2_1 _26474_ (.A0(net5064),
    .A1(net6297),
    .S(net4585),
    .X(_02980_));
 sg13g2_mux2_1 _26475_ (.A0(net5040),
    .A1(net6062),
    .S(net4585),
    .X(_02981_));
 sg13g2_nor2b_2 _26476_ (.A(_08592_),
    .B_N(net5211),
    .Y(_07860_));
 sg13g2_nand2b_1 _26477_ (.Y(_07861_),
    .B(net5210),
    .A_N(_08592_));
 sg13g2_nor2_1 _26478_ (.A(net6173),
    .B(_07860_),
    .Y(_07862_));
 sg13g2_a21oi_1 _26479_ (.A1(net5569),
    .A2(_08531_),
    .Y(_07863_),
    .B1(_07861_));
 sg13g2_a22oi_1 _26480_ (.Y(_07864_),
    .B1(_08535_),
    .B2(\atari2600.cpu.PC[13] ),
    .A2(_08528_),
    .A1(net5351));
 sg13g2_a21oi_1 _26481_ (.A1(_07863_),
    .A2(_07864_),
    .Y(_02982_),
    .B1(_07862_));
 sg13g2_a21oi_1 _26482_ (.A1(net5568),
    .A2(net5396),
    .Y(_07865_),
    .B1(_07861_));
 sg13g2_a22oi_1 _26483_ (.Y(_07866_),
    .B1(_08535_),
    .B2(\atari2600.cpu.PC[14] ),
    .A2(_08528_),
    .A1(\atari2600.cpu.DIMUX[6] ));
 sg13g2_a22oi_1 _26484_ (.Y(_02983_),
    .B1(_07865_),
    .B2(_07866_),
    .A2(_07861_),
    .A1(_08071_));
 sg13g2_nor2_1 _26485_ (.A(net6330),
    .B(_07860_),
    .Y(_07867_));
 sg13g2_nand2_1 _26486_ (.Y(_07868_),
    .A(\atari2600.cpu.ADD[7] ),
    .B(net5396));
 sg13g2_a221oi_1 _26487_ (.B2(\atari2600.cpu.PC[15] ),
    .C1(_07861_),
    .B1(_08535_),
    .A1(net5273),
    .Y(_07869_),
    .A2(_08528_));
 sg13g2_a21oi_1 _26488_ (.A1(_07868_),
    .A2(_07869_),
    .Y(_02984_),
    .B1(_07867_));
 sg13g2_or4_1 _26489_ (.A(_08175_),
    .B(net5205),
    .C(_08183_),
    .D(_08217_),
    .X(_07870_));
 sg13g2_nand2_1 _26490_ (.Y(_07871_),
    .A(_08446_),
    .B(_07186_));
 sg13g2_nor4_1 _26491_ (.A(net5275),
    .B(_08183_),
    .C(_08215_),
    .D(_07174_),
    .Y(_07872_));
 sg13g2_and2_1 _26492_ (.A(_08205_),
    .B(_07872_),
    .X(_07873_));
 sg13g2_o21ai_1 _26493_ (.B1(_07870_),
    .Y(_07874_),
    .A1(_08215_),
    .A2(_07228_));
 sg13g2_nor3_1 _26494_ (.A(_07231_),
    .B(_07873_),
    .C(_07874_),
    .Y(_07875_));
 sg13g2_a22oi_1 _26495_ (.Y(_02985_),
    .B1(_07871_),
    .B2(_07875_),
    .A2(net5347),
    .A1(_08054_));
 sg13g2_nor3_1 _26496_ (.A(_08184_),
    .B(_08454_),
    .C(_07212_),
    .Y(_07876_));
 sg13g2_nor4_1 _26497_ (.A(net5349),
    .B(_08405_),
    .C(_07874_),
    .D(_07876_),
    .Y(_07877_));
 sg13g2_a21oi_1 _26498_ (.A1(_08052_),
    .A2(net5349),
    .Y(_02986_),
    .B1(_07877_));
 sg13g2_a21oi_1 _26499_ (.A1(net5202),
    .A2(_07184_),
    .Y(_07878_),
    .B1(_07196_));
 sg13g2_nor3_1 _26500_ (.A(_08175_),
    .B(_08215_),
    .C(_07878_),
    .Y(_07879_));
 sg13g2_a21oi_1 _26501_ (.A1(_08216_),
    .A2(_07213_),
    .Y(_07880_),
    .B1(_07879_));
 sg13g2_and2_1 _26502_ (.A(_07189_),
    .B(_07213_),
    .X(_07881_));
 sg13g2_nor3_1 _26503_ (.A(_07231_),
    .B(_07872_),
    .C(_07881_),
    .Y(_07882_));
 sg13g2_a22oi_1 _26504_ (.Y(_02987_),
    .B1(_07880_),
    .B2(_07882_),
    .A2(net5349),
    .A1(_08053_));
 sg13g2_a22oi_1 _26505_ (.Y(_02988_),
    .B1(_07237_),
    .B2(_07880_),
    .A2(net5347),
    .A1(_08051_));
 sg13g2_nand2_1 _26506_ (.Y(_07883_),
    .A(net5204),
    .B(net5201));
 sg13g2_nor2_1 _26507_ (.A(_08248_),
    .B(_07883_),
    .Y(_07884_));
 sg13g2_a21oi_1 _26508_ (.A1(net5204),
    .A2(_08446_),
    .Y(_07885_),
    .B1(_07884_));
 sg13g2_nor2b_1 _26509_ (.A(_08450_),
    .B_N(_07885_),
    .Y(_07886_));
 sg13g2_nor2_1 _26510_ (.A(net3981),
    .B(net5270),
    .Y(_07887_));
 sg13g2_a21oi_1 _26511_ (.A1(net5270),
    .A2(_07886_),
    .Y(_02989_),
    .B1(_07887_));
 sg13g2_nand2b_1 _26512_ (.Y(_07888_),
    .B(net5199),
    .A_N(_07870_));
 sg13g2_nor2_1 _26513_ (.A(_08447_),
    .B(_07174_),
    .Y(_07889_));
 sg13g2_a22oi_1 _26514_ (.Y(_07890_),
    .B1(_07889_),
    .B2(net5275),
    .A2(_07173_),
    .A1(net5200));
 sg13g2_nand4_1 _26515_ (.B(_07230_),
    .C(_07888_),
    .A(_07197_),
    .Y(_07891_),
    .D(_07890_));
 sg13g2_nor4_1 _26516_ (.A(_08450_),
    .B(_07192_),
    .C(_07884_),
    .D(_07891_),
    .Y(_07892_));
 sg13g2_a21oi_1 _26517_ (.A1(_08060_),
    .A2(net5346),
    .Y(_02990_),
    .B1(_07892_));
 sg13g2_nor2_1 _26518_ (.A(net5346),
    .B(_07891_),
    .Y(_07893_));
 sg13g2_a221oi_1 _26519_ (.B2(_08246_),
    .C1(_07886_),
    .B1(_07884_),
    .A1(net5204),
    .Y(_07894_),
    .A2(_08446_));
 sg13g2_a22oi_1 _26520_ (.Y(_02991_),
    .B1(_07893_),
    .B2(_07894_),
    .A2(net5346),
    .A1(_08059_));
 sg13g2_nand3_1 _26521_ (.B(_07884_),
    .C(_07893_),
    .A(net5274),
    .Y(_07895_));
 sg13g2_o21ai_1 _26522_ (.B1(_07895_),
    .Y(_07896_),
    .A1(net7204),
    .A2(net5270));
 sg13g2_inv_1 _26523_ (.Y(_02992_),
    .A(_07896_));
 sg13g2_nand3_1 _26524_ (.B(_08595_),
    .C(_08634_),
    .A(_08590_),
    .Y(_07897_));
 sg13g2_nand2_1 _26525_ (.Y(_07898_),
    .A(net2972),
    .B(_07897_));
 sg13g2_nor2_2 _26526_ (.A(_08553_),
    .B(net4952),
    .Y(_07899_));
 sg13g2_o21ai_1 _26527_ (.B1(\atari2600.tia.vid_ypos[3] ),
    .Y(_07900_),
    .A1(\atari2600.tia.vid_ypos[2] ),
    .A2(_08136_));
 sg13g2_a21oi_1 _26528_ (.A1(_09823_),
    .A2(_07900_),
    .Y(_07901_),
    .B1(_10306_));
 sg13g2_nand2b_1 _26529_ (.Y(_07902_),
    .B(_00143_),
    .A_N(_07901_));
 sg13g2_a22oi_1 _26530_ (.Y(_07903_),
    .B1(_06442_),
    .B2(\atari2600.tia.cx[1] ),
    .A2(_06430_),
    .A1(\atari2600.tia.cx[2] ));
 sg13g2_a22oi_1 _26531_ (.Y(_07904_),
    .B1(_06614_),
    .B2(\atari2600.tia.cx[14] ),
    .A2(_08583_),
    .A1(\atari2600.tia.cx[4] ));
 sg13g2_a22oi_1 _26532_ (.Y(_07905_),
    .B1(_06807_),
    .B2(\atari2600.tia.cx[8] ),
    .A2(_05257_),
    .A1(\atari2600.tia.cx[12] ));
 sg13g2_nand2_1 _26533_ (.Y(_07906_),
    .A(_07904_),
    .B(_07905_));
 sg13g2_a22oi_1 _26534_ (.Y(_07907_),
    .B1(_07902_),
    .B2(_06454_),
    .A2(_07899_),
    .A1(\atari2600.input_joystick_0[1] ));
 sg13g2_a22oi_1 _26535_ (.Y(_07908_),
    .B1(_05260_),
    .B2(\atari2600.tia.cx[10] ),
    .A2(_08678_),
    .A1(\atari2600.tia.cx[6] ));
 sg13g2_nand3_1 _26536_ (.B(_07907_),
    .C(_07908_),
    .A(_07903_),
    .Y(_07909_));
 sg13g2_nor2_2 _26537_ (.A(_07906_),
    .B(_07909_),
    .Y(_07910_));
 sg13g2_a21oi_1 _26538_ (.A1(_08554_),
    .A2(net5029),
    .Y(_07911_),
    .B1(net5037));
 sg13g2_a21o_1 _26539_ (.A2(_07911_),
    .A1(_08676_),
    .B1(_07897_),
    .X(_07912_));
 sg13g2_o21ai_1 _26540_ (.B1(_07898_),
    .Y(_02993_),
    .A1(_07910_),
    .A2(_07912_));
 sg13g2_nand3_1 _26541_ (.B(net4870),
    .C(_08746_),
    .A(\atari2600.tia.cx[7] ),
    .Y(_07913_));
 sg13g2_nand2_1 _26542_ (.Y(_07914_),
    .A(\atari2600.tia.cx[11] ),
    .B(_05257_));
 sg13g2_a22oi_1 _26543_ (.Y(_07915_),
    .B1(_06614_),
    .B2(\atari2600.tia.cx[13] ),
    .A2(_08583_),
    .A1(\atari2600.tia.cx[3] ));
 sg13g2_a22oi_1 _26544_ (.Y(_07916_),
    .B1(_05260_),
    .B2(\atari2600.tia.cx[9] ),
    .A2(_08678_),
    .A1(\atari2600.tia.cx[5] ));
 sg13g2_nand4_1 _26545_ (.B(_07914_),
    .C(_07915_),
    .A(_07913_),
    .Y(_07917_),
    .D(_07916_));
 sg13g2_a21oi_2 _26546_ (.B1(_07917_),
    .Y(_07918_),
    .A2(_06442_),
    .A1(\atari2600.tia.cx[0] ));
 sg13g2_nand2_1 _26547_ (.Y(_07919_),
    .A(net2956),
    .B(_07897_));
 sg13g2_o21ai_1 _26548_ (.B1(_07919_),
    .Y(_02994_),
    .A1(_07912_),
    .A2(_07918_));
 sg13g2_dfrbp_1 _26549_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1233),
    .D(_00179_),
    .Q_N(_13223_),
    .Q(\scanline[69][0] ));
 sg13g2_dfrbp_1 _26550_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2635),
    .D(_00180_),
    .Q_N(_13222_),
    .Q(\scanline[69][1] ));
 sg13g2_dfrbp_1 _26551_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2634),
    .D(_00181_),
    .Q_N(_13221_),
    .Q(\scanline[69][2] ));
 sg13g2_dfrbp_1 _26552_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2633),
    .D(_00182_),
    .Q_N(_13220_),
    .Q(\scanline[69][3] ));
 sg13g2_dfrbp_1 _26553_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2632),
    .D(_00183_),
    .Q_N(_13219_),
    .Q(\scanline[69][4] ));
 sg13g2_dfrbp_1 _26554_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2631),
    .D(_00184_),
    .Q_N(_13218_),
    .Q(\scanline[69][5] ));
 sg13g2_dfrbp_1 _26555_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2630),
    .D(_00185_),
    .Q_N(_13217_),
    .Q(\scanline[69][6] ));
 sg13g2_dfrbp_1 _26556_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2629),
    .D(_00186_),
    .Q_N(_13216_),
    .Q(\scanline[154][0] ));
 sg13g2_dfrbp_1 _26557_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2628),
    .D(_00187_),
    .Q_N(_13215_),
    .Q(\scanline[154][1] ));
 sg13g2_dfrbp_1 _26558_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2627),
    .D(_00188_),
    .Q_N(_13214_),
    .Q(\scanline[154][2] ));
 sg13g2_dfrbp_1 _26559_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2626),
    .D(_00189_),
    .Q_N(_13213_),
    .Q(\scanline[154][3] ));
 sg13g2_dfrbp_1 _26560_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2625),
    .D(_00190_),
    .Q_N(_13212_),
    .Q(\scanline[154][4] ));
 sg13g2_dfrbp_1 _26561_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2624),
    .D(_00191_),
    .Q_N(_13211_),
    .Q(\scanline[154][5] ));
 sg13g2_dfrbp_1 _26562_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2623),
    .D(_00192_),
    .Q_N(_13210_),
    .Q(\scanline[154][6] ));
 sg13g2_dfrbp_1 _26563_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2622),
    .D(_00193_),
    .Q_N(_13209_),
    .Q(\flash_rom.addr[0] ));
 sg13g2_dfrbp_1 _26564_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2621),
    .D(_00194_),
    .Q_N(_13208_),
    .Q(\flash_rom.addr[1] ));
 sg13g2_dfrbp_1 _26565_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2620),
    .D(_00195_),
    .Q_N(_13207_),
    .Q(\flash_rom.addr[2] ));
 sg13g2_dfrbp_1 _26566_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2619),
    .D(_00196_),
    .Q_N(_13206_),
    .Q(\flash_rom.addr[3] ));
 sg13g2_dfrbp_1 _26567_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2618),
    .D(_00197_),
    .Q_N(_13205_),
    .Q(\flash_rom.addr[4] ));
 sg13g2_dfrbp_1 _26568_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net2617),
    .D(_00198_),
    .Q_N(_13204_),
    .Q(\flash_rom.addr[5] ));
 sg13g2_dfrbp_1 _26569_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net2616),
    .D(_00199_),
    .Q_N(_13203_),
    .Q(\flash_rom.addr[6] ));
 sg13g2_dfrbp_1 _26570_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2615),
    .D(net7141),
    .Q_N(_13202_),
    .Q(\flash_rom.addr[7] ));
 sg13g2_dfrbp_1 _26571_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2614),
    .D(net7112),
    .Q_N(_13201_),
    .Q(\flash_rom.addr[8] ));
 sg13g2_dfrbp_1 _26572_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2613),
    .D(_00202_),
    .Q_N(_13200_),
    .Q(\flash_rom.addr[9] ));
 sg13g2_dfrbp_1 _26573_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net2612),
    .D(_00203_),
    .Q_N(_13199_),
    .Q(\flash_rom.addr[10] ));
 sg13g2_dfrbp_1 _26574_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net2611),
    .D(_00204_),
    .Q_N(_13198_),
    .Q(\flash_rom.addr[11] ));
 sg13g2_dfrbp_1 _26575_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2610),
    .D(_00205_),
    .Q_N(_13197_),
    .Q(\scanline[59][0] ));
 sg13g2_dfrbp_1 _26576_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2609),
    .D(_00206_),
    .Q_N(_13196_),
    .Q(\scanline[59][1] ));
 sg13g2_dfrbp_1 _26577_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2608),
    .D(_00207_),
    .Q_N(_13195_),
    .Q(\scanline[59][2] ));
 sg13g2_dfrbp_1 _26578_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2607),
    .D(_00208_),
    .Q_N(_13194_),
    .Q(\scanline[59][3] ));
 sg13g2_dfrbp_1 _26579_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2606),
    .D(_00209_),
    .Q_N(_13193_),
    .Q(\scanline[59][4] ));
 sg13g2_dfrbp_1 _26580_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2605),
    .D(_00210_),
    .Q_N(_13192_),
    .Q(\scanline[59][5] ));
 sg13g2_dfrbp_1 _26581_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2604),
    .D(_00211_),
    .Q_N(_13191_),
    .Q(\scanline[59][6] ));
 sg13g2_dfrbp_1 _26582_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net2603),
    .D(_00212_),
    .Q_N(_13190_),
    .Q(\flash_rom.addr[16] ));
 sg13g2_dfrbp_1 _26583_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net2601),
    .D(net4010),
    .Q_N(_13189_),
    .Q(\flash_rom.addr[17] ));
 sg13g2_dfrbp_1 _26584_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2599),
    .D(net3647),
    .Q_N(_13188_),
    .Q(\flash_rom.addr[18] ));
 sg13g2_dfrbp_1 _26585_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2597),
    .D(_00215_),
    .Q_N(_13187_),
    .Q(\flash_rom.addr[19] ));
 sg13g2_dfrbp_1 _26586_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net2595),
    .D(_00216_),
    .Q_N(_13186_),
    .Q(\flash_rom.addr[21] ));
 sg13g2_dfrbp_1 _26587_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net2593),
    .D(net3711),
    .Q_N(_13185_),
    .Q(\flash_rom.addr[22] ));
 sg13g2_dfrbp_1 _26588_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net2591),
    .D(net3708),
    .Q_N(_13184_),
    .Q(\flash_rom.addr[23] ));
 sg13g2_dfrbp_1 _26589_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2589),
    .D(_00219_),
    .Q_N(_13183_),
    .Q(\scanline[32][0] ));
 sg13g2_dfrbp_1 _26590_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2588),
    .D(_00220_),
    .Q_N(_13182_),
    .Q(\scanline[32][1] ));
 sg13g2_dfrbp_1 _26591_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2587),
    .D(_00221_),
    .Q_N(_13181_),
    .Q(\scanline[32][2] ));
 sg13g2_dfrbp_1 _26592_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2586),
    .D(_00222_),
    .Q_N(_13180_),
    .Q(\scanline[32][3] ));
 sg13g2_dfrbp_1 _26593_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2585),
    .D(_00223_),
    .Q_N(_13179_),
    .Q(\scanline[32][4] ));
 sg13g2_dfrbp_1 _26594_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2584),
    .D(_00224_),
    .Q_N(_13178_),
    .Q(\scanline[32][5] ));
 sg13g2_dfrbp_1 _26595_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2583),
    .D(_00225_),
    .Q_N(_13177_),
    .Q(\scanline[32][6] ));
 sg13g2_dfrbp_1 _26596_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2582),
    .D(_00226_),
    .Q_N(_13176_),
    .Q(\scanline[31][0] ));
 sg13g2_dfrbp_1 _26597_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2581),
    .D(_00227_),
    .Q_N(_13175_),
    .Q(\scanline[31][1] ));
 sg13g2_dfrbp_1 _26598_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2580),
    .D(_00228_),
    .Q_N(_13174_),
    .Q(\scanline[31][2] ));
 sg13g2_dfrbp_1 _26599_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2579),
    .D(_00229_),
    .Q_N(_13173_),
    .Q(\scanline[31][3] ));
 sg13g2_dfrbp_1 _26600_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2578),
    .D(_00230_),
    .Q_N(_13172_),
    .Q(\scanline[31][4] ));
 sg13g2_dfrbp_1 _26601_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2577),
    .D(_00231_),
    .Q_N(_13171_),
    .Q(\scanline[31][5] ));
 sg13g2_dfrbp_1 _26602_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2576),
    .D(_00232_),
    .Q_N(_13170_),
    .Q(\scanline[31][6] ));
 sg13g2_dfrbp_1 _26603_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2575),
    .D(_00233_),
    .Q_N(_13169_),
    .Q(\scanline[30][0] ));
 sg13g2_dfrbp_1 _26604_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2574),
    .D(_00234_),
    .Q_N(_13168_),
    .Q(\scanline[30][1] ));
 sg13g2_dfrbp_1 _26605_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2573),
    .D(_00235_),
    .Q_N(_13167_),
    .Q(\scanline[30][2] ));
 sg13g2_dfrbp_1 _26606_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2572),
    .D(_00236_),
    .Q_N(_13166_),
    .Q(\scanline[30][3] ));
 sg13g2_dfrbp_1 _26607_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2571),
    .D(_00237_),
    .Q_N(_13165_),
    .Q(\scanline[30][4] ));
 sg13g2_dfrbp_1 _26608_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2570),
    .D(_00238_),
    .Q_N(_13164_),
    .Q(\scanline[30][5] ));
 sg13g2_dfrbp_1 _26609_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2569),
    .D(_00239_),
    .Q_N(_13163_),
    .Q(\scanline[30][6] ));
 sg13g2_dfrbp_1 _26610_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2568),
    .D(_00240_),
    .Q_N(_13162_),
    .Q(\scanline[2][0] ));
 sg13g2_dfrbp_1 _26611_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2567),
    .D(_00241_),
    .Q_N(_13161_),
    .Q(\scanline[2][1] ));
 sg13g2_dfrbp_1 _26612_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2566),
    .D(_00242_),
    .Q_N(_13160_),
    .Q(\scanline[2][2] ));
 sg13g2_dfrbp_1 _26613_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2565),
    .D(_00243_),
    .Q_N(_13159_),
    .Q(\scanline[2][3] ));
 sg13g2_dfrbp_1 _26614_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2564),
    .D(_00244_),
    .Q_N(_13158_),
    .Q(\scanline[2][4] ));
 sg13g2_dfrbp_1 _26615_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2563),
    .D(_00245_),
    .Q_N(_13157_),
    .Q(\scanline[2][5] ));
 sg13g2_dfrbp_1 _26616_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2562),
    .D(_00246_),
    .Q_N(_13156_),
    .Q(\scanline[2][6] ));
 sg13g2_dfrbp_1 _26617_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2561),
    .D(_00247_),
    .Q_N(_13155_),
    .Q(\scanline[28][0] ));
 sg13g2_dfrbp_1 _26618_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2560),
    .D(_00248_),
    .Q_N(_13154_),
    .Q(\scanline[28][1] ));
 sg13g2_dfrbp_1 _26619_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2559),
    .D(_00249_),
    .Q_N(_13153_),
    .Q(\scanline[28][2] ));
 sg13g2_dfrbp_1 _26620_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2558),
    .D(_00250_),
    .Q_N(_13152_),
    .Q(\scanline[28][3] ));
 sg13g2_dfrbp_1 _26621_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2557),
    .D(_00251_),
    .Q_N(_13151_),
    .Q(\scanline[28][4] ));
 sg13g2_dfrbp_1 _26622_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2556),
    .D(_00252_),
    .Q_N(_13150_),
    .Q(\scanline[28][5] ));
 sg13g2_dfrbp_1 _26623_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2555),
    .D(_00253_),
    .Q_N(_13149_),
    .Q(\scanline[28][6] ));
 sg13g2_dfrbp_1 _26624_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2554),
    .D(_00254_),
    .Q_N(_13148_),
    .Q(\scanline[27][0] ));
 sg13g2_dfrbp_1 _26625_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2553),
    .D(_00255_),
    .Q_N(_13147_),
    .Q(\scanline[27][1] ));
 sg13g2_dfrbp_1 _26626_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2552),
    .D(_00256_),
    .Q_N(_13146_),
    .Q(\scanline[27][2] ));
 sg13g2_dfrbp_1 _26627_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2551),
    .D(_00257_),
    .Q_N(_13145_),
    .Q(\scanline[27][3] ));
 sg13g2_dfrbp_1 _26628_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2550),
    .D(_00258_),
    .Q_N(_13144_),
    .Q(\scanline[27][4] ));
 sg13g2_dfrbp_1 _26629_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2549),
    .D(_00259_),
    .Q_N(_13143_),
    .Q(\scanline[27][5] ));
 sg13g2_dfrbp_1 _26630_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2548),
    .D(_00260_),
    .Q_N(_13142_),
    .Q(\scanline[27][6] ));
 sg13g2_dfrbp_1 _26631_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2547),
    .D(_00261_),
    .Q_N(_13141_),
    .Q(\scanline[26][0] ));
 sg13g2_dfrbp_1 _26632_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2546),
    .D(_00262_),
    .Q_N(_13140_),
    .Q(\scanline[26][1] ));
 sg13g2_dfrbp_1 _26633_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2545),
    .D(_00263_),
    .Q_N(_13139_),
    .Q(\scanline[26][2] ));
 sg13g2_dfrbp_1 _26634_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2544),
    .D(_00264_),
    .Q_N(_13138_),
    .Q(\scanline[26][3] ));
 sg13g2_dfrbp_1 _26635_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2543),
    .D(_00265_),
    .Q_N(_13137_),
    .Q(\scanline[26][4] ));
 sg13g2_dfrbp_1 _26636_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2542),
    .D(_00266_),
    .Q_N(_13136_),
    .Q(\scanline[26][5] ));
 sg13g2_dfrbp_1 _26637_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2541),
    .D(_00267_),
    .Q_N(_13135_),
    .Q(\scanline[26][6] ));
 sg13g2_dfrbp_1 _26638_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2540),
    .D(_00268_),
    .Q_N(_13134_),
    .Q(\scanline[25][0] ));
 sg13g2_dfrbp_1 _26639_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2539),
    .D(_00269_),
    .Q_N(_13133_),
    .Q(\scanline[25][1] ));
 sg13g2_dfrbp_1 _26640_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2538),
    .D(_00270_),
    .Q_N(_13132_),
    .Q(\scanline[25][2] ));
 sg13g2_dfrbp_1 _26641_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2537),
    .D(_00271_),
    .Q_N(_13131_),
    .Q(\scanline[25][3] ));
 sg13g2_dfrbp_1 _26642_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2536),
    .D(_00272_),
    .Q_N(_13130_),
    .Q(\scanline[25][4] ));
 sg13g2_dfrbp_1 _26643_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2535),
    .D(_00273_),
    .Q_N(_13129_),
    .Q(\scanline[25][5] ));
 sg13g2_dfrbp_1 _26644_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2534),
    .D(_00274_),
    .Q_N(_13128_),
    .Q(\scanline[25][6] ));
 sg13g2_dfrbp_1 _26645_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2533),
    .D(_00275_),
    .Q_N(_13127_),
    .Q(\scanline[61][0] ));
 sg13g2_dfrbp_1 _26646_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2532),
    .D(_00276_),
    .Q_N(_13126_),
    .Q(\scanline[61][1] ));
 sg13g2_dfrbp_1 _26647_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2531),
    .D(_00277_),
    .Q_N(_13125_),
    .Q(\scanline[61][2] ));
 sg13g2_dfrbp_1 _26648_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2530),
    .D(_00278_),
    .Q_N(_13124_),
    .Q(\scanline[61][3] ));
 sg13g2_dfrbp_1 _26649_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2529),
    .D(_00279_),
    .Q_N(_13123_),
    .Q(\scanline[61][4] ));
 sg13g2_dfrbp_1 _26650_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2528),
    .D(_00280_),
    .Q_N(_13122_),
    .Q(\scanline[61][5] ));
 sg13g2_dfrbp_1 _26651_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2527),
    .D(_00281_),
    .Q_N(_13121_),
    .Q(\scanline[61][6] ));
 sg13g2_dfrbp_1 _26652_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2526),
    .D(_00282_),
    .Q_N(_13120_),
    .Q(\scanline[60][0] ));
 sg13g2_dfrbp_1 _26653_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2525),
    .D(_00283_),
    .Q_N(_13119_),
    .Q(\scanline[60][1] ));
 sg13g2_dfrbp_1 _26654_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2524),
    .D(_00284_),
    .Q_N(_13118_),
    .Q(\scanline[60][2] ));
 sg13g2_dfrbp_1 _26655_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2523),
    .D(_00285_),
    .Q_N(_13117_),
    .Q(\scanline[60][3] ));
 sg13g2_dfrbp_1 _26656_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2522),
    .D(_00286_),
    .Q_N(_13116_),
    .Q(\scanline[60][4] ));
 sg13g2_dfrbp_1 _26657_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2521),
    .D(_00287_),
    .Q_N(_13115_),
    .Q(\scanline[60][5] ));
 sg13g2_dfrbp_1 _26658_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2520),
    .D(_00288_),
    .Q_N(_13114_),
    .Q(\scanline[60][6] ));
 sg13g2_dfrbp_1 _26659_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net2518),
    .D(_00289_),
    .Q_N(_13113_),
    .Q(\atari2600.ram[87][0] ));
 sg13g2_dfrbp_1 _26660_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2517),
    .D(_00290_),
    .Q_N(_13112_),
    .Q(\atari2600.ram[87][1] ));
 sg13g2_dfrbp_1 _26661_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2516),
    .D(_00291_),
    .Q_N(_13111_),
    .Q(\atari2600.ram[87][2] ));
 sg13g2_dfrbp_1 _26662_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net2515),
    .D(_00292_),
    .Q_N(_13110_),
    .Q(\atari2600.ram[87][3] ));
 sg13g2_dfrbp_1 _26663_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net2514),
    .D(_00293_),
    .Q_N(_13109_),
    .Q(\atari2600.ram[87][4] ));
 sg13g2_dfrbp_1 _26664_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2513),
    .D(_00294_),
    .Q_N(_13108_),
    .Q(\atari2600.ram[87][5] ));
 sg13g2_dfrbp_1 _26665_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net2512),
    .D(_00295_),
    .Q_N(_13107_),
    .Q(\atari2600.ram[87][6] ));
 sg13g2_dfrbp_1 _26666_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net2511),
    .D(_00296_),
    .Q_N(_13106_),
    .Q(\atari2600.ram[87][7] ));
 sg13g2_dfrbp_1 _26667_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2509),
    .D(_00297_),
    .Q_N(_13105_),
    .Q(\atari2600.ram[27][0] ));
 sg13g2_dfrbp_1 _26668_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net2508),
    .D(_00298_),
    .Q_N(_13104_),
    .Q(\atari2600.ram[27][1] ));
 sg13g2_dfrbp_1 _26669_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net2507),
    .D(_00299_),
    .Q_N(_13103_),
    .Q(\atari2600.ram[27][2] ));
 sg13g2_dfrbp_1 _26670_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2506),
    .D(_00300_),
    .Q_N(_13102_),
    .Q(\atari2600.ram[27][3] ));
 sg13g2_dfrbp_1 _26671_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net2505),
    .D(_00301_),
    .Q_N(_13101_),
    .Q(\atari2600.ram[27][4] ));
 sg13g2_dfrbp_1 _26672_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net2504),
    .D(_00302_),
    .Q_N(_13100_),
    .Q(\atari2600.ram[27][5] ));
 sg13g2_dfrbp_1 _26673_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2503),
    .D(_00303_),
    .Q_N(_13099_),
    .Q(\atari2600.ram[27][6] ));
 sg13g2_dfrbp_1 _26674_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2502),
    .D(_00304_),
    .Q_N(_13098_),
    .Q(\atari2600.ram[27][7] ));
 sg13g2_dfrbp_1 _26675_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2501),
    .D(_00305_),
    .Q_N(_13097_),
    .Q(\scanline[159][0] ));
 sg13g2_dfrbp_1 _26676_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2500),
    .D(_00306_),
    .Q_N(_13096_),
    .Q(\scanline[159][1] ));
 sg13g2_dfrbp_1 _26677_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2499),
    .D(_00307_),
    .Q_N(_13095_),
    .Q(\scanline[159][2] ));
 sg13g2_dfrbp_1 _26678_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2498),
    .D(_00308_),
    .Q_N(_13094_),
    .Q(\scanline[159][3] ));
 sg13g2_dfrbp_1 _26679_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2497),
    .D(_00309_),
    .Q_N(_13093_),
    .Q(\scanline[159][4] ));
 sg13g2_dfrbp_1 _26680_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2496),
    .D(_00310_),
    .Q_N(_13092_),
    .Q(\scanline[159][5] ));
 sg13g2_dfrbp_1 _26681_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2495),
    .D(_00311_),
    .Q_N(_13091_),
    .Q(\scanline[159][6] ));
 sg13g2_dfrbp_1 _26682_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2494),
    .D(_00312_),
    .Q_N(_13090_),
    .Q(\atari2600.ram[90][0] ));
 sg13g2_dfrbp_1 _26683_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2493),
    .D(_00313_),
    .Q_N(_13089_),
    .Q(\atari2600.ram[90][1] ));
 sg13g2_dfrbp_1 _26684_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net2492),
    .D(_00314_),
    .Q_N(_13088_),
    .Q(\atari2600.ram[90][2] ));
 sg13g2_dfrbp_1 _26685_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net2491),
    .D(_00315_),
    .Q_N(_13087_),
    .Q(\atari2600.ram[90][3] ));
 sg13g2_dfrbp_1 _26686_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2490),
    .D(_00316_),
    .Q_N(_13086_),
    .Q(\atari2600.ram[90][4] ));
 sg13g2_dfrbp_1 _26687_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net2489),
    .D(_00317_),
    .Q_N(_13085_),
    .Q(\atari2600.ram[90][5] ));
 sg13g2_dfrbp_1 _26688_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2488),
    .D(_00318_),
    .Q_N(_13084_),
    .Q(\atari2600.ram[90][6] ));
 sg13g2_dfrbp_1 _26689_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2487),
    .D(_00319_),
    .Q_N(_13083_),
    .Q(\atari2600.ram[90][7] ));
 sg13g2_dfrbp_1 _26690_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2486),
    .D(_00320_),
    .Q_N(_13082_),
    .Q(\atari2600.ram[70][0] ));
 sg13g2_dfrbp_1 _26691_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2485),
    .D(_00321_),
    .Q_N(_13081_),
    .Q(\atari2600.ram[70][1] ));
 sg13g2_dfrbp_1 _26692_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2484),
    .D(_00322_),
    .Q_N(_13080_),
    .Q(\atari2600.ram[70][2] ));
 sg13g2_dfrbp_1 _26693_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2483),
    .D(_00323_),
    .Q_N(_13079_),
    .Q(\atari2600.ram[70][3] ));
 sg13g2_dfrbp_1 _26694_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2482),
    .D(_00324_),
    .Q_N(_13078_),
    .Q(\atari2600.ram[70][4] ));
 sg13g2_dfrbp_1 _26695_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2481),
    .D(_00325_),
    .Q_N(_13077_),
    .Q(\atari2600.ram[70][5] ));
 sg13g2_dfrbp_1 _26696_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2480),
    .D(_00326_),
    .Q_N(_13076_),
    .Q(\atari2600.ram[70][6] ));
 sg13g2_dfrbp_1 _26697_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2479),
    .D(_00327_),
    .Q_N(_13075_),
    .Q(\atari2600.ram[70][7] ));
 sg13g2_dfrbp_1 _26698_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2478),
    .D(_00328_),
    .Q_N(_13074_),
    .Q(\scanline[149][0] ));
 sg13g2_dfrbp_1 _26699_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2477),
    .D(_00329_),
    .Q_N(_13073_),
    .Q(\scanline[149][1] ));
 sg13g2_dfrbp_1 _26700_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2476),
    .D(_00330_),
    .Q_N(_13072_),
    .Q(\scanline[149][2] ));
 sg13g2_dfrbp_1 _26701_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2475),
    .D(_00331_),
    .Q_N(_13071_),
    .Q(\scanline[149][3] ));
 sg13g2_dfrbp_1 _26702_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2474),
    .D(_00332_),
    .Q_N(_13070_),
    .Q(\scanline[149][4] ));
 sg13g2_dfrbp_1 _26703_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2473),
    .D(_00333_),
    .Q_N(_13069_),
    .Q(\scanline[149][5] ));
 sg13g2_dfrbp_1 _26704_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2472),
    .D(_00334_),
    .Q_N(_13068_),
    .Q(\scanline[149][6] ));
 sg13g2_dfrbp_1 _26705_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2471),
    .D(_00335_),
    .Q_N(_13067_),
    .Q(\scanline[139][0] ));
 sg13g2_dfrbp_1 _26706_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2470),
    .D(_00336_),
    .Q_N(_13066_),
    .Q(\scanline[139][1] ));
 sg13g2_dfrbp_1 _26707_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2469),
    .D(_00337_),
    .Q_N(_13065_),
    .Q(\scanline[139][2] ));
 sg13g2_dfrbp_1 _26708_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2468),
    .D(_00338_),
    .Q_N(_13064_),
    .Q(\scanline[139][3] ));
 sg13g2_dfrbp_1 _26709_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2467),
    .D(_00339_),
    .Q_N(_13063_),
    .Q(\scanline[139][4] ));
 sg13g2_dfrbp_1 _26710_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net2466),
    .D(_00340_),
    .Q_N(_13062_),
    .Q(\scanline[139][5] ));
 sg13g2_dfrbp_1 _26711_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2465),
    .D(_00341_),
    .Q_N(_13061_),
    .Q(\scanline[139][6] ));
 sg13g2_dfrbp_1 _26712_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2464),
    .D(_00342_),
    .Q_N(_13060_),
    .Q(\scanline[129][0] ));
 sg13g2_dfrbp_1 _26713_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2463),
    .D(_00343_),
    .Q_N(_13059_),
    .Q(\scanline[129][1] ));
 sg13g2_dfrbp_1 _26714_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2462),
    .D(_00344_),
    .Q_N(_13058_),
    .Q(\scanline[129][2] ));
 sg13g2_dfrbp_1 _26715_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2461),
    .D(_00345_),
    .Q_N(_13057_),
    .Q(\scanline[129][3] ));
 sg13g2_dfrbp_1 _26716_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2460),
    .D(_00346_),
    .Q_N(_13056_),
    .Q(\scanline[129][4] ));
 sg13g2_dfrbp_1 _26717_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2459),
    .D(_00347_),
    .Q_N(_13055_),
    .Q(\scanline[129][5] ));
 sg13g2_dfrbp_1 _26718_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2458),
    .D(_00348_),
    .Q_N(_13054_),
    .Q(\scanline[129][6] ));
 sg13g2_dfrbp_1 _26719_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2457),
    .D(_00349_),
    .Q_N(_13053_),
    .Q(\scanline[119][0] ));
 sg13g2_dfrbp_1 _26720_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2456),
    .D(_00350_),
    .Q_N(_13052_),
    .Q(\scanline[119][1] ));
 sg13g2_dfrbp_1 _26721_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2455),
    .D(_00351_),
    .Q_N(_13051_),
    .Q(\scanline[119][2] ));
 sg13g2_dfrbp_1 _26722_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2454),
    .D(_00352_),
    .Q_N(_13050_),
    .Q(\scanline[119][3] ));
 sg13g2_dfrbp_1 _26723_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2453),
    .D(_00353_),
    .Q_N(_13049_),
    .Q(\scanline[119][4] ));
 sg13g2_dfrbp_1 _26724_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2452),
    .D(_00354_),
    .Q_N(_13048_),
    .Q(\scanline[119][5] ));
 sg13g2_dfrbp_1 _26725_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2451),
    .D(_00355_),
    .Q_N(_13047_),
    .Q(\scanline[119][6] ));
 sg13g2_dfrbp_1 _26726_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2450),
    .D(_00356_),
    .Q_N(_13046_),
    .Q(\scanline[109][0] ));
 sg13g2_dfrbp_1 _26727_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2449),
    .D(_00357_),
    .Q_N(_13045_),
    .Q(\scanline[109][1] ));
 sg13g2_dfrbp_1 _26728_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2448),
    .D(_00358_),
    .Q_N(_13044_),
    .Q(\scanline[109][2] ));
 sg13g2_dfrbp_1 _26729_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net2447),
    .D(_00359_),
    .Q_N(_13043_),
    .Q(\scanline[109][3] ));
 sg13g2_dfrbp_1 _26730_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2446),
    .D(_00360_),
    .Q_N(_13042_),
    .Q(\scanline[109][4] ));
 sg13g2_dfrbp_1 _26731_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2445),
    .D(_00361_),
    .Q_N(_13041_),
    .Q(\scanline[109][5] ));
 sg13g2_dfrbp_1 _26732_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2444),
    .D(_00362_),
    .Q_N(_13040_),
    .Q(\scanline[109][6] ));
 sg13g2_dfrbp_1 _26733_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2442),
    .D(_00363_),
    .Q_N(_13039_),
    .Q(\scanline[126][0] ));
 sg13g2_dfrbp_1 _26734_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2441),
    .D(_00364_),
    .Q_N(_13038_),
    .Q(\scanline[126][1] ));
 sg13g2_dfrbp_1 _26735_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2440),
    .D(_00365_),
    .Q_N(_13037_),
    .Q(\scanline[126][2] ));
 sg13g2_dfrbp_1 _26736_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2439),
    .D(_00366_),
    .Q_N(_13036_),
    .Q(\scanline[126][3] ));
 sg13g2_dfrbp_1 _26737_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2438),
    .D(_00367_),
    .Q_N(_13035_),
    .Q(\scanline[126][4] ));
 sg13g2_dfrbp_1 _26738_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2437),
    .D(_00368_),
    .Q_N(_13034_),
    .Q(\scanline[126][5] ));
 sg13g2_dfrbp_1 _26739_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2436),
    .D(_00369_),
    .Q_N(_13033_),
    .Q(\scanline[126][6] ));
 sg13g2_dfrbp_1 _26740_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2435),
    .D(_00370_),
    .Q_N(_13032_),
    .Q(\scanline[125][0] ));
 sg13g2_dfrbp_1 _26741_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2434),
    .D(_00371_),
    .Q_N(_13031_),
    .Q(\scanline[125][1] ));
 sg13g2_dfrbp_1 _26742_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2433),
    .D(_00372_),
    .Q_N(_13030_),
    .Q(\scanline[125][2] ));
 sg13g2_dfrbp_1 _26743_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2432),
    .D(_00373_),
    .Q_N(_13029_),
    .Q(\scanline[125][3] ));
 sg13g2_dfrbp_1 _26744_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2431),
    .D(_00374_),
    .Q_N(_13028_),
    .Q(\scanline[125][4] ));
 sg13g2_dfrbp_1 _26745_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2430),
    .D(_00375_),
    .Q_N(_13027_),
    .Q(\scanline[125][5] ));
 sg13g2_dfrbp_1 _26746_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2429),
    .D(_00376_),
    .Q_N(_13026_),
    .Q(\scanline[125][6] ));
 sg13g2_dfrbp_1 _26747_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2428),
    .D(_00377_),
    .Q_N(_13025_),
    .Q(\scanline[124][0] ));
 sg13g2_dfrbp_1 _26748_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2427),
    .D(_00378_),
    .Q_N(_13024_),
    .Q(\scanline[124][1] ));
 sg13g2_dfrbp_1 _26749_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2426),
    .D(_00379_),
    .Q_N(_13023_),
    .Q(\scanline[124][2] ));
 sg13g2_dfrbp_1 _26750_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2425),
    .D(_00380_),
    .Q_N(_13022_),
    .Q(\scanline[124][3] ));
 sg13g2_dfrbp_1 _26751_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2424),
    .D(_00381_),
    .Q_N(_13021_),
    .Q(\scanline[124][4] ));
 sg13g2_dfrbp_1 _26752_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2423),
    .D(_00382_),
    .Q_N(_13020_),
    .Q(\scanline[124][5] ));
 sg13g2_dfrbp_1 _26753_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2422),
    .D(_00383_),
    .Q_N(_13019_),
    .Q(\scanline[124][6] ));
 sg13g2_dfrbp_1 _26754_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2421),
    .D(_00384_),
    .Q_N(_13018_),
    .Q(\atari2600.ram[72][0] ));
 sg13g2_dfrbp_1 _26755_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2420),
    .D(_00385_),
    .Q_N(_13017_),
    .Q(\atari2600.ram[72][1] ));
 sg13g2_dfrbp_1 _26756_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2411),
    .D(_00386_),
    .Q_N(_13016_),
    .Q(\atari2600.ram[72][2] ));
 sg13g2_dfrbp_1 _26757_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2410),
    .D(_00387_),
    .Q_N(_13015_),
    .Q(\atari2600.ram[72][3] ));
 sg13g2_dfrbp_1 _26758_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2409),
    .D(_00388_),
    .Q_N(_13014_),
    .Q(\atari2600.ram[72][4] ));
 sg13g2_dfrbp_1 _26759_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2408),
    .D(_00389_),
    .Q_N(_13013_),
    .Q(\atari2600.ram[72][5] ));
 sg13g2_dfrbp_1 _26760_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2407),
    .D(_00390_),
    .Q_N(_13012_),
    .Q(\atari2600.ram[72][6] ));
 sg13g2_dfrbp_1 _26761_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2406),
    .D(_00391_),
    .Q_N(_13011_),
    .Q(\atari2600.ram[72][7] ));
 sg13g2_dfrbp_1 _26762_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2405),
    .D(_00392_),
    .Q_N(_13010_),
    .Q(\scanline[99][0] ));
 sg13g2_dfrbp_1 _26763_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2404),
    .D(_00393_),
    .Q_N(_13009_),
    .Q(\scanline[99][1] ));
 sg13g2_dfrbp_1 _26764_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2403),
    .D(_00394_),
    .Q_N(_13008_),
    .Q(\scanline[99][2] ));
 sg13g2_dfrbp_1 _26765_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2402),
    .D(_00395_),
    .Q_N(_13007_),
    .Q(\scanline[99][3] ));
 sg13g2_dfrbp_1 _26766_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2401),
    .D(_00396_),
    .Q_N(_13006_),
    .Q(\scanline[99][4] ));
 sg13g2_dfrbp_1 _26767_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2400),
    .D(_00397_),
    .Q_N(_13005_),
    .Q(\scanline[99][5] ));
 sg13g2_dfrbp_1 _26768_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2399),
    .D(_00398_),
    .Q_N(_13004_),
    .Q(\scanline[99][6] ));
 sg13g2_dfrbp_1 _26769_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2398),
    .D(_00399_),
    .Q_N(_13003_),
    .Q(\scanline[5][0] ));
 sg13g2_dfrbp_1 _26770_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2397),
    .D(_00400_),
    .Q_N(_13002_),
    .Q(\scanline[5][1] ));
 sg13g2_dfrbp_1 _26771_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2396),
    .D(_00401_),
    .Q_N(_13001_),
    .Q(\scanline[5][2] ));
 sg13g2_dfrbp_1 _26772_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2395),
    .D(_00402_),
    .Q_N(_13000_),
    .Q(\scanline[5][3] ));
 sg13g2_dfrbp_1 _26773_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2394),
    .D(_00403_),
    .Q_N(_12999_),
    .Q(\scanline[5][4] ));
 sg13g2_dfrbp_1 _26774_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2393),
    .D(_00404_),
    .Q_N(_12998_),
    .Q(\scanline[5][5] ));
 sg13g2_dfrbp_1 _26775_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2392),
    .D(_00405_),
    .Q_N(_12997_),
    .Q(\scanline[5][6] ));
 sg13g2_dfrbp_1 _26776_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2391),
    .D(_00406_),
    .Q_N(_12996_),
    .Q(\scanline[89][0] ));
 sg13g2_dfrbp_1 _26777_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2390),
    .D(_00407_),
    .Q_N(_12995_),
    .Q(\scanline[89][1] ));
 sg13g2_dfrbp_1 _26778_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2389),
    .D(_00408_),
    .Q_N(_12994_),
    .Q(\scanline[89][2] ));
 sg13g2_dfrbp_1 _26779_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2388),
    .D(_00409_),
    .Q_N(_12993_),
    .Q(\scanline[89][3] ));
 sg13g2_dfrbp_1 _26780_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2387),
    .D(_00410_),
    .Q_N(_12992_),
    .Q(\scanline[89][4] ));
 sg13g2_dfrbp_1 _26781_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2386),
    .D(_00411_),
    .Q_N(_12991_),
    .Q(\scanline[89][5] ));
 sg13g2_dfrbp_1 _26782_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2385),
    .D(_00412_),
    .Q_N(_12990_),
    .Q(\scanline[89][6] ));
 sg13g2_dfrbp_1 _26783_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2384),
    .D(_00413_),
    .Q_N(_12989_),
    .Q(\scanline[58][0] ));
 sg13g2_dfrbp_1 _26784_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2383),
    .D(_00414_),
    .Q_N(_12988_),
    .Q(\scanline[58][1] ));
 sg13g2_dfrbp_1 _26785_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2382),
    .D(_00415_),
    .Q_N(_12987_),
    .Q(\scanline[58][2] ));
 sg13g2_dfrbp_1 _26786_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2381),
    .D(_00416_),
    .Q_N(_12986_),
    .Q(\scanline[58][3] ));
 sg13g2_dfrbp_1 _26787_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2380),
    .D(_00417_),
    .Q_N(_12985_),
    .Q(\scanline[58][4] ));
 sg13g2_dfrbp_1 _26788_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2379),
    .D(_00418_),
    .Q_N(_12984_),
    .Q(\scanline[58][5] ));
 sg13g2_dfrbp_1 _26789_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2378),
    .D(_00419_),
    .Q_N(_12983_),
    .Q(\scanline[58][6] ));
 sg13g2_dfrbp_1 _26790_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2377),
    .D(_00420_),
    .Q_N(_12982_),
    .Q(\scanline[79][0] ));
 sg13g2_dfrbp_1 _26791_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2376),
    .D(_00421_),
    .Q_N(_12981_),
    .Q(\scanline[79][1] ));
 sg13g2_dfrbp_1 _26792_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2375),
    .D(_00422_),
    .Q_N(_12980_),
    .Q(\scanline[79][2] ));
 sg13g2_dfrbp_1 _26793_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2374),
    .D(_00423_),
    .Q_N(_12979_),
    .Q(\scanline[79][3] ));
 sg13g2_dfrbp_1 _26794_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2373),
    .D(_00424_),
    .Q_N(_12978_),
    .Q(\scanline[79][4] ));
 sg13g2_dfrbp_1 _26795_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2372),
    .D(_00425_),
    .Q_N(_12977_),
    .Q(\scanline[79][5] ));
 sg13g2_dfrbp_1 _26796_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2371),
    .D(_00426_),
    .Q_N(_12976_),
    .Q(\scanline[79][6] ));
 sg13g2_dfrbp_1 _26797_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2370),
    .D(_00427_),
    .Q_N(_12975_),
    .Q(\scanline[123][0] ));
 sg13g2_dfrbp_1 _26798_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2369),
    .D(_00428_),
    .Q_N(_12974_),
    .Q(\scanline[123][1] ));
 sg13g2_dfrbp_1 _26799_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2368),
    .D(_00429_),
    .Q_N(_12973_),
    .Q(\scanline[123][2] ));
 sg13g2_dfrbp_1 _26800_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2367),
    .D(_00430_),
    .Q_N(_12972_),
    .Q(\scanline[123][3] ));
 sg13g2_dfrbp_1 _26801_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2366),
    .D(_00431_),
    .Q_N(_12971_),
    .Q(\scanline[123][4] ));
 sg13g2_dfrbp_1 _26802_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2365),
    .D(_00432_),
    .Q_N(_12970_),
    .Q(\scanline[123][5] ));
 sg13g2_dfrbp_1 _26803_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2364),
    .D(_00433_),
    .Q_N(_12969_),
    .Q(\scanline[123][6] ));
 sg13g2_dfrbp_1 _26804_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2359),
    .D(_00434_),
    .Q_N(_12968_),
    .Q(\scanline[153][0] ));
 sg13g2_dfrbp_1 _26805_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2358),
    .D(_00435_),
    .Q_N(_12967_),
    .Q(\scanline[153][1] ));
 sg13g2_dfrbp_1 _26806_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2357),
    .D(_00436_),
    .Q_N(_12966_),
    .Q(\scanline[153][2] ));
 sg13g2_dfrbp_1 _26807_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2356),
    .D(_00437_),
    .Q_N(_12965_),
    .Q(\scanline[153][3] ));
 sg13g2_dfrbp_1 _26808_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2355),
    .D(_00438_),
    .Q_N(_12964_),
    .Q(\scanline[153][4] ));
 sg13g2_dfrbp_1 _26809_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2354),
    .D(_00439_),
    .Q_N(_12963_),
    .Q(\scanline[153][5] ));
 sg13g2_dfrbp_1 _26810_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2353),
    .D(_00440_),
    .Q_N(_12962_),
    .Q(\scanline[153][6] ));
 sg13g2_dfrbp_1 _26811_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2352),
    .D(_00441_),
    .Q_N(_12961_),
    .Q(\scanline[122][0] ));
 sg13g2_dfrbp_1 _26812_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2351),
    .D(_00442_),
    .Q_N(_12960_),
    .Q(\scanline[122][1] ));
 sg13g2_dfrbp_1 _26813_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2350),
    .D(_00443_),
    .Q_N(_12959_),
    .Q(\scanline[122][2] ));
 sg13g2_dfrbp_1 _26814_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2349),
    .D(_00444_),
    .Q_N(_12958_),
    .Q(\scanline[122][3] ));
 sg13g2_dfrbp_1 _26815_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2348),
    .D(_00445_),
    .Q_N(_12957_),
    .Q(\scanline[122][4] ));
 sg13g2_dfrbp_1 _26816_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2347),
    .D(_00446_),
    .Q_N(_12956_),
    .Q(\scanline[122][5] ));
 sg13g2_dfrbp_1 _26817_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2346),
    .D(_00447_),
    .Q_N(_12955_),
    .Q(\scanline[122][6] ));
 sg13g2_dfrbp_1 _26818_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2345),
    .D(_00448_),
    .Q_N(_12954_),
    .Q(\scanline[121][0] ));
 sg13g2_dfrbp_1 _26819_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2344),
    .D(_00449_),
    .Q_N(_12953_),
    .Q(\scanline[121][1] ));
 sg13g2_dfrbp_1 _26820_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2343),
    .D(_00450_),
    .Q_N(_12952_),
    .Q(\scanline[121][2] ));
 sg13g2_dfrbp_1 _26821_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2342),
    .D(_00451_),
    .Q_N(_12951_),
    .Q(\scanline[121][3] ));
 sg13g2_dfrbp_1 _26822_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2341),
    .D(_00452_),
    .Q_N(_12950_),
    .Q(\scanline[121][4] ));
 sg13g2_dfrbp_1 _26823_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2340),
    .D(_00453_),
    .Q_N(_12949_),
    .Q(\scanline[121][5] ));
 sg13g2_dfrbp_1 _26824_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2339),
    .D(_00454_),
    .Q_N(_12948_),
    .Q(\scanline[121][6] ));
 sg13g2_dfrbp_1 _26825_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2338),
    .D(_00455_),
    .Q_N(_12947_),
    .Q(\scanline[120][0] ));
 sg13g2_dfrbp_1 _26826_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2337),
    .D(_00456_),
    .Q_N(_12946_),
    .Q(\scanline[120][1] ));
 sg13g2_dfrbp_1 _26827_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2336),
    .D(_00457_),
    .Q_N(_12945_),
    .Q(\scanline[120][2] ));
 sg13g2_dfrbp_1 _26828_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2335),
    .D(_00458_),
    .Q_N(_12944_),
    .Q(\scanline[120][3] ));
 sg13g2_dfrbp_1 _26829_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2334),
    .D(_00459_),
    .Q_N(_12943_),
    .Q(\scanline[120][4] ));
 sg13g2_dfrbp_1 _26830_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2333),
    .D(_00460_),
    .Q_N(_12942_),
    .Q(\scanline[120][5] ));
 sg13g2_dfrbp_1 _26831_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2332),
    .D(_00461_),
    .Q_N(_12941_),
    .Q(\scanline[120][6] ));
 sg13g2_dfrbp_1 _26832_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2331),
    .D(_00462_),
    .Q_N(_12940_),
    .Q(\scanline[152][0] ));
 sg13g2_dfrbp_1 _26833_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2330),
    .D(_00463_),
    .Q_N(_12939_),
    .Q(\scanline[152][1] ));
 sg13g2_dfrbp_1 _26834_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2329),
    .D(_00464_),
    .Q_N(_12938_),
    .Q(\scanline[152][2] ));
 sg13g2_dfrbp_1 _26835_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2328),
    .D(_00465_),
    .Q_N(_12937_),
    .Q(\scanline[152][3] ));
 sg13g2_dfrbp_1 _26836_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2327),
    .D(_00466_),
    .Q_N(_12936_),
    .Q(\scanline[152][4] ));
 sg13g2_dfrbp_1 _26837_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2326),
    .D(_00467_),
    .Q_N(_12935_),
    .Q(\scanline[152][5] ));
 sg13g2_dfrbp_1 _26838_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2325),
    .D(_00468_),
    .Q_N(_12934_),
    .Q(\scanline[152][6] ));
 sg13g2_dfrbp_1 _26839_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2324),
    .D(_00469_),
    .Q_N(_12933_),
    .Q(\scanline[11][0] ));
 sg13g2_dfrbp_1 _26840_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2323),
    .D(_00470_),
    .Q_N(_12932_),
    .Q(\scanline[11][1] ));
 sg13g2_dfrbp_1 _26841_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2322),
    .D(_00471_),
    .Q_N(_12931_),
    .Q(\scanline[11][2] ));
 sg13g2_dfrbp_1 _26842_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2321),
    .D(_00472_),
    .Q_N(_12930_),
    .Q(\scanline[11][3] ));
 sg13g2_dfrbp_1 _26843_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2320),
    .D(_00473_),
    .Q_N(_12929_),
    .Q(\scanline[11][4] ));
 sg13g2_dfrbp_1 _26844_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2319),
    .D(_00474_),
    .Q_N(_12928_),
    .Q(\scanline[11][5] ));
 sg13g2_dfrbp_1 _26845_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2318),
    .D(_00475_),
    .Q_N(_12927_),
    .Q(\scanline[11][6] ));
 sg13g2_dfrbp_1 _26846_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2317),
    .D(_00476_),
    .Q_N(_12926_),
    .Q(\scanline[151][0] ));
 sg13g2_dfrbp_1 _26847_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2316),
    .D(_00477_),
    .Q_N(_12925_),
    .Q(\scanline[151][1] ));
 sg13g2_dfrbp_1 _26848_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2315),
    .D(_00478_),
    .Q_N(_12924_),
    .Q(\scanline[151][2] ));
 sg13g2_dfrbp_1 _26849_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2314),
    .D(_00479_),
    .Q_N(_12923_),
    .Q(\scanline[151][3] ));
 sg13g2_dfrbp_1 _26850_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2313),
    .D(_00480_),
    .Q_N(_12922_),
    .Q(\scanline[151][4] ));
 sg13g2_dfrbp_1 _26851_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2312),
    .D(_00481_),
    .Q_N(_12921_),
    .Q(\scanline[151][5] ));
 sg13g2_dfrbp_1 _26852_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2311),
    .D(_00482_),
    .Q_N(_12920_),
    .Q(\scanline[151][6] ));
 sg13g2_dfrbp_1 _26853_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2310),
    .D(_00483_),
    .Q_N(_12919_),
    .Q(\scanline[118][0] ));
 sg13g2_dfrbp_1 _26854_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2309),
    .D(_00484_),
    .Q_N(_12918_),
    .Q(\scanline[118][1] ));
 sg13g2_dfrbp_1 _26855_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2308),
    .D(_00485_),
    .Q_N(_12917_),
    .Q(\scanline[118][2] ));
 sg13g2_dfrbp_1 _26856_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2307),
    .D(_00486_),
    .Q_N(_12916_),
    .Q(\scanline[118][3] ));
 sg13g2_dfrbp_1 _26857_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2306),
    .D(_00487_),
    .Q_N(_12915_),
    .Q(\scanline[118][4] ));
 sg13g2_dfrbp_1 _26858_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2305),
    .D(_00488_),
    .Q_N(_12914_),
    .Q(\scanline[118][5] ));
 sg13g2_dfrbp_1 _26859_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2304),
    .D(_00489_),
    .Q_N(_12913_),
    .Q(\scanline[118][6] ));
 sg13g2_dfrbp_1 _26860_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2303),
    .D(_00490_),
    .Q_N(_12912_),
    .Q(\scanline[150][0] ));
 sg13g2_dfrbp_1 _26861_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2302),
    .D(_00491_),
    .Q_N(_12911_),
    .Q(\scanline[150][1] ));
 sg13g2_dfrbp_1 _26862_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2301),
    .D(_00492_),
    .Q_N(_12910_),
    .Q(\scanline[150][2] ));
 sg13g2_dfrbp_1 _26863_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2300),
    .D(_00493_),
    .Q_N(_12909_),
    .Q(\scanline[150][3] ));
 sg13g2_dfrbp_1 _26864_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2299),
    .D(_00494_),
    .Q_N(_12908_),
    .Q(\scanline[150][4] ));
 sg13g2_dfrbp_1 _26865_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2298),
    .D(_00495_),
    .Q_N(_12907_),
    .Q(\scanline[150][5] ));
 sg13g2_dfrbp_1 _26866_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2297),
    .D(_00496_),
    .Q_N(_12906_),
    .Q(\scanline[150][6] ));
 sg13g2_dfrbp_1 _26867_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2296),
    .D(_00497_),
    .Q_N(_12905_),
    .Q(\scanline[117][0] ));
 sg13g2_dfrbp_1 _26868_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2295),
    .D(_00498_),
    .Q_N(_12904_),
    .Q(\scanline[117][1] ));
 sg13g2_dfrbp_1 _26869_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2294),
    .D(_00499_),
    .Q_N(_12903_),
    .Q(\scanline[117][2] ));
 sg13g2_dfrbp_1 _26870_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2293),
    .D(_00500_),
    .Q_N(_12902_),
    .Q(\scanline[117][3] ));
 sg13g2_dfrbp_1 _26871_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2292),
    .D(_00501_),
    .Q_N(_12901_),
    .Q(\scanline[117][4] ));
 sg13g2_dfrbp_1 _26872_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2291),
    .D(_00502_),
    .Q_N(_12900_),
    .Q(\scanline[117][5] ));
 sg13g2_dfrbp_1 _26873_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2290),
    .D(_00503_),
    .Q_N(_12899_),
    .Q(\scanline[117][6] ));
 sg13g2_dfrbp_1 _26874_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2289),
    .D(_00504_),
    .Q_N(_12898_),
    .Q(\scanline[14][0] ));
 sg13g2_dfrbp_1 _26875_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2288),
    .D(_00505_),
    .Q_N(_12897_),
    .Q(\scanline[14][1] ));
 sg13g2_dfrbp_1 _26876_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2287),
    .D(_00506_),
    .Q_N(_12896_),
    .Q(\scanline[14][2] ));
 sg13g2_dfrbp_1 _26877_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2286),
    .D(_00507_),
    .Q_N(_12895_),
    .Q(\scanline[14][3] ));
 sg13g2_dfrbp_1 _26878_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2285),
    .D(_00508_),
    .Q_N(_12894_),
    .Q(\scanline[14][4] ));
 sg13g2_dfrbp_1 _26879_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2284),
    .D(_00509_),
    .Q_N(_12893_),
    .Q(\scanline[14][5] ));
 sg13g2_dfrbp_1 _26880_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2283),
    .D(_00510_),
    .Q_N(_12892_),
    .Q(\scanline[14][6] ));
 sg13g2_dfrbp_1 _26881_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2282),
    .D(_00511_),
    .Q_N(_12891_),
    .Q(\scanline[116][0] ));
 sg13g2_dfrbp_1 _26882_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2281),
    .D(_00512_),
    .Q_N(_12890_),
    .Q(\scanline[116][1] ));
 sg13g2_dfrbp_1 _26883_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2280),
    .D(_00513_),
    .Q_N(_12889_),
    .Q(\scanline[116][2] ));
 sg13g2_dfrbp_1 _26884_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2279),
    .D(_00514_),
    .Q_N(_12888_),
    .Q(\scanline[116][3] ));
 sg13g2_dfrbp_1 _26885_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2278),
    .D(_00515_),
    .Q_N(_12887_),
    .Q(\scanline[116][4] ));
 sg13g2_dfrbp_1 _26886_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2277),
    .D(_00516_),
    .Q_N(_12886_),
    .Q(\scanline[116][5] ));
 sg13g2_dfrbp_1 _26887_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2276),
    .D(_00517_),
    .Q_N(_12885_),
    .Q(\scanline[116][6] ));
 sg13g2_dfrbp_1 _26888_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2275),
    .D(_00518_),
    .Q_N(_12884_),
    .Q(\scanline[148][0] ));
 sg13g2_dfrbp_1 _26889_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2274),
    .D(_00519_),
    .Q_N(_12883_),
    .Q(\scanline[148][1] ));
 sg13g2_dfrbp_1 _26890_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2273),
    .D(_00520_),
    .Q_N(_12882_),
    .Q(\scanline[148][2] ));
 sg13g2_dfrbp_1 _26891_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2272),
    .D(_00521_),
    .Q_N(_12881_),
    .Q(\scanline[148][3] ));
 sg13g2_dfrbp_1 _26892_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2271),
    .D(_00522_),
    .Q_N(_12880_),
    .Q(\scanline[148][4] ));
 sg13g2_dfrbp_1 _26893_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2270),
    .D(_00523_),
    .Q_N(_12879_),
    .Q(\scanline[148][5] ));
 sg13g2_dfrbp_1 _26894_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2269),
    .D(_00524_),
    .Q_N(_12878_),
    .Q(\scanline[148][6] ));
 sg13g2_dfrbp_1 _26895_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2268),
    .D(_00525_),
    .Q_N(_12877_),
    .Q(\scanline[115][0] ));
 sg13g2_dfrbp_1 _26896_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2267),
    .D(_00526_),
    .Q_N(_12876_),
    .Q(\scanline[115][1] ));
 sg13g2_dfrbp_1 _26897_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2266),
    .D(_00527_),
    .Q_N(_12875_),
    .Q(\scanline[115][2] ));
 sg13g2_dfrbp_1 _26898_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2265),
    .D(_00528_),
    .Q_N(_12874_),
    .Q(\scanline[115][3] ));
 sg13g2_dfrbp_1 _26899_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2264),
    .D(_00529_),
    .Q_N(_12873_),
    .Q(\scanline[115][4] ));
 sg13g2_dfrbp_1 _26900_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2263),
    .D(_00530_),
    .Q_N(_12872_),
    .Q(\scanline[115][5] ));
 sg13g2_dfrbp_1 _26901_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2262),
    .D(_00531_),
    .Q_N(_12871_),
    .Q(\scanline[115][6] ));
 sg13g2_dfrbp_1 _26902_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2261),
    .D(_00532_),
    .Q_N(_12870_),
    .Q(\scanline[147][0] ));
 sg13g2_dfrbp_1 _26903_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2260),
    .D(_00533_),
    .Q_N(_12869_),
    .Q(\scanline[147][1] ));
 sg13g2_dfrbp_1 _26904_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2259),
    .D(_00534_),
    .Q_N(_12868_),
    .Q(\scanline[147][2] ));
 sg13g2_dfrbp_1 _26905_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2258),
    .D(_00535_),
    .Q_N(_12867_),
    .Q(\scanline[147][3] ));
 sg13g2_dfrbp_1 _26906_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2257),
    .D(_00536_),
    .Q_N(_12866_),
    .Q(\scanline[147][4] ));
 sg13g2_dfrbp_1 _26907_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2256),
    .D(_00537_),
    .Q_N(_12865_),
    .Q(\scanline[147][5] ));
 sg13g2_dfrbp_1 _26908_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2255),
    .D(_00538_),
    .Q_N(_12864_),
    .Q(\scanline[147][6] ));
 sg13g2_dfrbp_1 _26909_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2254),
    .D(_00539_),
    .Q_N(_12863_),
    .Q(\scanline[114][0] ));
 sg13g2_dfrbp_1 _26910_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2253),
    .D(_00540_),
    .Q_N(_12862_),
    .Q(\scanline[114][1] ));
 sg13g2_dfrbp_1 _26911_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2252),
    .D(_00541_),
    .Q_N(_12861_),
    .Q(\scanline[114][2] ));
 sg13g2_dfrbp_1 _26912_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2251),
    .D(_00542_),
    .Q_N(_12860_),
    .Q(\scanline[114][3] ));
 sg13g2_dfrbp_1 _26913_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2250),
    .D(_00543_),
    .Q_N(_12859_),
    .Q(\scanline[114][4] ));
 sg13g2_dfrbp_1 _26914_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2249),
    .D(_00544_),
    .Q_N(_12858_),
    .Q(\scanline[114][5] ));
 sg13g2_dfrbp_1 _26915_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2248),
    .D(_00545_),
    .Q_N(_12857_),
    .Q(\scanline[114][6] ));
 sg13g2_dfrbp_1 _26916_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2247),
    .D(_00546_),
    .Q_N(_12856_),
    .Q(\scanline[146][0] ));
 sg13g2_dfrbp_1 _26917_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2246),
    .D(_00547_),
    .Q_N(_12855_),
    .Q(\scanline[146][1] ));
 sg13g2_dfrbp_1 _26918_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2245),
    .D(_00548_),
    .Q_N(_12854_),
    .Q(\scanline[146][2] ));
 sg13g2_dfrbp_1 _26919_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2244),
    .D(_00549_),
    .Q_N(_12853_),
    .Q(\scanline[146][3] ));
 sg13g2_dfrbp_1 _26920_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2243),
    .D(_00550_),
    .Q_N(_12852_),
    .Q(\scanline[146][4] ));
 sg13g2_dfrbp_1 _26921_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2242),
    .D(_00551_),
    .Q_N(_12851_),
    .Q(\scanline[146][5] ));
 sg13g2_dfrbp_1 _26922_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2241),
    .D(_00552_),
    .Q_N(_12850_),
    .Q(\scanline[146][6] ));
 sg13g2_dfrbp_1 _26923_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2240),
    .D(_00553_),
    .Q_N(_12849_),
    .Q(\scanline[113][0] ));
 sg13g2_dfrbp_1 _26924_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2239),
    .D(_00554_),
    .Q_N(_12848_),
    .Q(\scanline[113][1] ));
 sg13g2_dfrbp_1 _26925_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2238),
    .D(_00555_),
    .Q_N(_12847_),
    .Q(\scanline[113][2] ));
 sg13g2_dfrbp_1 _26926_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2237),
    .D(_00556_),
    .Q_N(_12846_),
    .Q(\scanline[113][3] ));
 sg13g2_dfrbp_1 _26927_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2236),
    .D(_00557_),
    .Q_N(_12845_),
    .Q(\scanline[113][4] ));
 sg13g2_dfrbp_1 _26928_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2235),
    .D(_00558_),
    .Q_N(_12844_),
    .Q(\scanline[113][5] ));
 sg13g2_dfrbp_1 _26929_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2234),
    .D(_00559_),
    .Q_N(_12843_),
    .Q(\scanline[113][6] ));
 sg13g2_dfrbp_1 _26930_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2233),
    .D(_00560_),
    .Q_N(_12842_),
    .Q(\scanline[145][0] ));
 sg13g2_dfrbp_1 _26931_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2232),
    .D(_00561_),
    .Q_N(_12841_),
    .Q(\scanline[145][1] ));
 sg13g2_dfrbp_1 _26932_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2231),
    .D(_00562_),
    .Q_N(_12840_),
    .Q(\scanline[145][2] ));
 sg13g2_dfrbp_1 _26933_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2230),
    .D(_00563_),
    .Q_N(_12839_),
    .Q(\scanline[145][3] ));
 sg13g2_dfrbp_1 _26934_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2229),
    .D(_00564_),
    .Q_N(_12838_),
    .Q(\scanline[145][4] ));
 sg13g2_dfrbp_1 _26935_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2228),
    .D(_00565_),
    .Q_N(_12837_),
    .Q(\scanline[145][5] ));
 sg13g2_dfrbp_1 _26936_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2227),
    .D(_00566_),
    .Q_N(_12836_),
    .Q(\scanline[145][6] ));
 sg13g2_dfrbp_1 _26937_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2226),
    .D(_00567_),
    .Q_N(_12835_),
    .Q(\scanline[112][0] ));
 sg13g2_dfrbp_1 _26938_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2225),
    .D(_00568_),
    .Q_N(_12834_),
    .Q(\scanline[112][1] ));
 sg13g2_dfrbp_1 _26939_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2224),
    .D(_00569_),
    .Q_N(_12833_),
    .Q(\scanline[112][2] ));
 sg13g2_dfrbp_1 _26940_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2223),
    .D(_00570_),
    .Q_N(_12832_),
    .Q(\scanline[112][3] ));
 sg13g2_dfrbp_1 _26941_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2222),
    .D(_00571_),
    .Q_N(_12831_),
    .Q(\scanline[112][4] ));
 sg13g2_dfrbp_1 _26942_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2221),
    .D(_00572_),
    .Q_N(_12830_),
    .Q(\scanline[112][5] ));
 sg13g2_dfrbp_1 _26943_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2220),
    .D(_00573_),
    .Q_N(_12829_),
    .Q(\scanline[112][6] ));
 sg13g2_dfrbp_1 _26944_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2219),
    .D(_00574_),
    .Q_N(_12828_),
    .Q(\scanline[144][0] ));
 sg13g2_dfrbp_1 _26945_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2218),
    .D(_00575_),
    .Q_N(_12827_),
    .Q(\scanline[144][1] ));
 sg13g2_dfrbp_1 _26946_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2217),
    .D(_00576_),
    .Q_N(_12826_),
    .Q(\scanline[144][2] ));
 sg13g2_dfrbp_1 _26947_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2216),
    .D(_00577_),
    .Q_N(_12825_),
    .Q(\scanline[144][3] ));
 sg13g2_dfrbp_1 _26948_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2215),
    .D(_00578_),
    .Q_N(_12824_),
    .Q(\scanline[144][4] ));
 sg13g2_dfrbp_1 _26949_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2214),
    .D(_00579_),
    .Q_N(_12823_),
    .Q(\scanline[144][5] ));
 sg13g2_dfrbp_1 _26950_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2213),
    .D(_00580_),
    .Q_N(_12822_),
    .Q(\scanline[144][6] ));
 sg13g2_dfrbp_1 _26951_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2212),
    .D(_00581_),
    .Q_N(_12821_),
    .Q(\scanline[111][0] ));
 sg13g2_dfrbp_1 _26952_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net2211),
    .D(_00582_),
    .Q_N(_12820_),
    .Q(\scanline[111][1] ));
 sg13g2_dfrbp_1 _26953_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2210),
    .D(_00583_),
    .Q_N(_12819_),
    .Q(\scanline[111][2] ));
 sg13g2_dfrbp_1 _26954_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2209),
    .D(_00584_),
    .Q_N(_12818_),
    .Q(\scanline[111][3] ));
 sg13g2_dfrbp_1 _26955_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net2208),
    .D(_00585_),
    .Q_N(_12817_),
    .Q(\scanline[111][4] ));
 sg13g2_dfrbp_1 _26956_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net2207),
    .D(_00586_),
    .Q_N(_12816_),
    .Q(\scanline[111][5] ));
 sg13g2_dfrbp_1 _26957_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2206),
    .D(_00587_),
    .Q_N(_12815_),
    .Q(\scanline[111][6] ));
 sg13g2_dfrbp_1 _26958_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2205),
    .D(_00588_),
    .Q_N(_12814_),
    .Q(\scanline[23][0] ));
 sg13g2_dfrbp_1 _26959_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2204),
    .D(_00589_),
    .Q_N(_12813_),
    .Q(\scanline[23][1] ));
 sg13g2_dfrbp_1 _26960_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2203),
    .D(_00590_),
    .Q_N(_12812_),
    .Q(\scanline[23][2] ));
 sg13g2_dfrbp_1 _26961_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2202),
    .D(_00591_),
    .Q_N(_12811_),
    .Q(\scanline[23][3] ));
 sg13g2_dfrbp_1 _26962_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2201),
    .D(_00592_),
    .Q_N(_12810_),
    .Q(\scanline[23][4] ));
 sg13g2_dfrbp_1 _26963_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2200),
    .D(_00593_),
    .Q_N(_12809_),
    .Q(\scanline[23][5] ));
 sg13g2_dfrbp_1 _26964_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2199),
    .D(_00594_),
    .Q_N(_12808_),
    .Q(\scanline[23][6] ));
 sg13g2_dfrbp_1 _26965_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2183),
    .D(_00595_),
    .Q_N(_12807_),
    .Q(\scanline[22][0] ));
 sg13g2_dfrbp_1 _26966_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2182),
    .D(_00596_),
    .Q_N(_12806_),
    .Q(\scanline[22][1] ));
 sg13g2_dfrbp_1 _26967_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2181),
    .D(_00597_),
    .Q_N(_12805_),
    .Q(\scanline[22][2] ));
 sg13g2_dfrbp_1 _26968_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2180),
    .D(_00598_),
    .Q_N(_12804_),
    .Q(\scanline[22][3] ));
 sg13g2_dfrbp_1 _26969_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2179),
    .D(_00599_),
    .Q_N(_12803_),
    .Q(\scanline[22][4] ));
 sg13g2_dfrbp_1 _26970_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2178),
    .D(_00600_),
    .Q_N(_12802_),
    .Q(\scanline[22][5] ));
 sg13g2_dfrbp_1 _26971_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2177),
    .D(_00601_),
    .Q_N(_12801_),
    .Q(\scanline[22][6] ));
 sg13g2_dfrbp_1 _26972_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2176),
    .D(_00602_),
    .Q_N(_12800_),
    .Q(\scanline[21][0] ));
 sg13g2_dfrbp_1 _26973_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2175),
    .D(_00603_),
    .Q_N(_12799_),
    .Q(\scanline[21][1] ));
 sg13g2_dfrbp_1 _26974_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2174),
    .D(_00604_),
    .Q_N(_12798_),
    .Q(\scanline[21][2] ));
 sg13g2_dfrbp_1 _26975_ (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2173),
    .D(_00605_),
    .Q_N(_12797_),
    .Q(\scanline[21][3] ));
 sg13g2_dfrbp_1 _26976_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2172),
    .D(_00606_),
    .Q_N(_12796_),
    .Q(\scanline[21][4] ));
 sg13g2_dfrbp_1 _26977_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2171),
    .D(_00607_),
    .Q_N(_12795_),
    .Q(\scanline[21][5] ));
 sg13g2_dfrbp_1 _26978_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2170),
    .D(_00608_),
    .Q_N(_12794_),
    .Q(\scanline[21][6] ));
 sg13g2_dfrbp_1 _26979_ (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2153),
    .D(_00609_),
    .Q_N(_12793_),
    .Q(\scanline[20][0] ));
 sg13g2_dfrbp_1 _26980_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2152),
    .D(_00610_),
    .Q_N(_12792_),
    .Q(\scanline[20][1] ));
 sg13g2_dfrbp_1 _26981_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2151),
    .D(_00611_),
    .Q_N(_12791_),
    .Q(\scanline[20][2] ));
 sg13g2_dfrbp_1 _26982_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2150),
    .D(_00612_),
    .Q_N(_12790_),
    .Q(\scanline[20][3] ));
 sg13g2_dfrbp_1 _26983_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2149),
    .D(_00613_),
    .Q_N(_12789_),
    .Q(\scanline[20][4] ));
 sg13g2_dfrbp_1 _26984_ (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2148),
    .D(_00614_),
    .Q_N(_12788_),
    .Q(\scanline[20][5] ));
 sg13g2_dfrbp_1 _26985_ (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2147),
    .D(_00615_),
    .Q_N(_12787_),
    .Q(\scanline[20][6] ));
 sg13g2_dfrbp_1 _26986_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2146),
    .D(_00616_),
    .Q_N(_12786_),
    .Q(\scanline[1][0] ));
 sg13g2_dfrbp_1 _26987_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2145),
    .D(_00617_),
    .Q_N(_12785_),
    .Q(\scanline[1][1] ));
 sg13g2_dfrbp_1 _26988_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2144),
    .D(_00618_),
    .Q_N(_12784_),
    .Q(\scanline[1][2] ));
 sg13g2_dfrbp_1 _26989_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2143),
    .D(_00619_),
    .Q_N(_12783_),
    .Q(\scanline[1][3] ));
 sg13g2_dfrbp_1 _26990_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2142),
    .D(_00620_),
    .Q_N(_12782_),
    .Q(\scanline[1][4] ));
 sg13g2_dfrbp_1 _26991_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2141),
    .D(_00621_),
    .Q_N(_12781_),
    .Q(\scanline[1][5] ));
 sg13g2_dfrbp_1 _26992_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2140),
    .D(_00622_),
    .Q_N(_12780_),
    .Q(\scanline[1][6] ));
 sg13g2_dfrbp_1 _26993_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2139),
    .D(_00623_),
    .Q_N(_12779_),
    .Q(\scanline[24][0] ));
 sg13g2_dfrbp_1 _26994_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2138),
    .D(_00624_),
    .Q_N(_12778_),
    .Q(\scanline[24][1] ));
 sg13g2_dfrbp_1 _26995_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2137),
    .D(_00625_),
    .Q_N(_12777_),
    .Q(\scanline[24][2] ));
 sg13g2_dfrbp_1 _26996_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2136),
    .D(_00626_),
    .Q_N(_12776_),
    .Q(\scanline[24][3] ));
 sg13g2_dfrbp_1 _26997_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2135),
    .D(_00627_),
    .Q_N(_12775_),
    .Q(\scanline[24][4] ));
 sg13g2_dfrbp_1 _26998_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2134),
    .D(_00628_),
    .Q_N(_12774_),
    .Q(\scanline[24][5] ));
 sg13g2_dfrbp_1 _26999_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2133),
    .D(_00629_),
    .Q_N(_12773_),
    .Q(\scanline[24][6] ));
 sg13g2_dfrbp_1 _27000_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2132),
    .D(_00630_),
    .Q_N(_12772_),
    .Q(\scanline[18][0] ));
 sg13g2_dfrbp_1 _27001_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2131),
    .D(_00631_),
    .Q_N(_12771_),
    .Q(\scanline[18][1] ));
 sg13g2_dfrbp_1 _27002_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2130),
    .D(_00632_),
    .Q_N(_12770_),
    .Q(\scanline[18][2] ));
 sg13g2_dfrbp_1 _27003_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2129),
    .D(_00633_),
    .Q_N(_12769_),
    .Q(\scanline[18][3] ));
 sg13g2_dfrbp_1 _27004_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2128),
    .D(_00634_),
    .Q_N(_12768_),
    .Q(\scanline[18][4] ));
 sg13g2_dfrbp_1 _27005_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2127),
    .D(_00635_),
    .Q_N(_12767_),
    .Q(\scanline[18][5] ));
 sg13g2_dfrbp_1 _27006_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2126),
    .D(_00636_),
    .Q_N(_12766_),
    .Q(\scanline[18][6] ));
 sg13g2_dfrbp_1 _27007_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2125),
    .D(_00637_),
    .Q_N(_12765_),
    .Q(\scanline[17][0] ));
 sg13g2_dfrbp_1 _27008_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2124),
    .D(_00638_),
    .Q_N(_12764_),
    .Q(\scanline[17][1] ));
 sg13g2_dfrbp_1 _27009_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2123),
    .D(_00639_),
    .Q_N(_12763_),
    .Q(\scanline[17][2] ));
 sg13g2_dfrbp_1 _27010_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2122),
    .D(_00640_),
    .Q_N(_12762_),
    .Q(\scanline[17][3] ));
 sg13g2_dfrbp_1 _27011_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2121),
    .D(_00641_),
    .Q_N(_12761_),
    .Q(\scanline[17][4] ));
 sg13g2_dfrbp_1 _27012_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2120),
    .D(_00642_),
    .Q_N(_12760_),
    .Q(\scanline[17][5] ));
 sg13g2_dfrbp_1 _27013_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2119),
    .D(_00643_),
    .Q_N(_12759_),
    .Q(\scanline[17][6] ));
 sg13g2_dfrbp_1 _27014_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2118),
    .D(_00644_),
    .Q_N(_12758_),
    .Q(\scanline[16][0] ));
 sg13g2_dfrbp_1 _27015_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2117),
    .D(_00645_),
    .Q_N(_12757_),
    .Q(\scanline[16][1] ));
 sg13g2_dfrbp_1 _27016_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2116),
    .D(_00646_),
    .Q_N(_12756_),
    .Q(\scanline[16][2] ));
 sg13g2_dfrbp_1 _27017_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2115),
    .D(_00647_),
    .Q_N(_12755_),
    .Q(\scanline[16][3] ));
 sg13g2_dfrbp_1 _27018_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2114),
    .D(_00648_),
    .Q_N(_12754_),
    .Q(\scanline[16][4] ));
 sg13g2_dfrbp_1 _27019_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2113),
    .D(_00649_),
    .Q_N(_12753_),
    .Q(\scanline[16][5] ));
 sg13g2_dfrbp_1 _27020_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2112),
    .D(_00650_),
    .Q_N(_12752_),
    .Q(\scanline[16][6] ));
 sg13g2_dfrbp_1 _27021_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2111),
    .D(_00651_),
    .Q_N(_12751_),
    .Q(\scanline[15][0] ));
 sg13g2_dfrbp_1 _27022_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2110),
    .D(_00652_),
    .Q_N(_12750_),
    .Q(\scanline[15][1] ));
 sg13g2_dfrbp_1 _27023_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net2109),
    .D(_00653_),
    .Q_N(_12749_),
    .Q(\scanline[15][2] ));
 sg13g2_dfrbp_1 _27024_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2108),
    .D(_00654_),
    .Q_N(_12748_),
    .Q(\scanline[15][3] ));
 sg13g2_dfrbp_1 _27025_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2107),
    .D(_00655_),
    .Q_N(_12747_),
    .Q(\scanline[15][4] ));
 sg13g2_dfrbp_1 _27026_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2106),
    .D(_00656_),
    .Q_N(_12746_),
    .Q(\scanline[15][5] ));
 sg13g2_dfrbp_1 _27027_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2105),
    .D(_00657_),
    .Q_N(_12745_),
    .Q(\scanline[15][6] ));
 sg13g2_dfrbp_1 _27028_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2104),
    .D(_00658_),
    .Q_N(_12744_),
    .Q(\scanline[158][0] ));
 sg13g2_dfrbp_1 _27029_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2103),
    .D(_00659_),
    .Q_N(_12743_),
    .Q(\scanline[158][1] ));
 sg13g2_dfrbp_1 _27030_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2102),
    .D(_00660_),
    .Q_N(_12742_),
    .Q(\scanline[158][2] ));
 sg13g2_dfrbp_1 _27031_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2101),
    .D(_00661_),
    .Q_N(_12741_),
    .Q(\scanline[158][3] ));
 sg13g2_dfrbp_1 _27032_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2100),
    .D(_00662_),
    .Q_N(_12740_),
    .Q(\scanline[158][4] ));
 sg13g2_dfrbp_1 _27033_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2099),
    .D(_00663_),
    .Q_N(_12739_),
    .Q(\scanline[158][5] ));
 sg13g2_dfrbp_1 _27034_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2098),
    .D(_00664_),
    .Q_N(_12738_),
    .Q(\scanline[158][6] ));
 sg13g2_dfrbp_1 _27035_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2097),
    .D(_00665_),
    .Q_N(_12737_),
    .Q(\scanline[157][0] ));
 sg13g2_dfrbp_1 _27036_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2096),
    .D(_00666_),
    .Q_N(_12736_),
    .Q(\scanline[157][1] ));
 sg13g2_dfrbp_1 _27037_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2095),
    .D(_00667_),
    .Q_N(_12735_),
    .Q(\scanline[157][2] ));
 sg13g2_dfrbp_1 _27038_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2094),
    .D(_00668_),
    .Q_N(_12734_),
    .Q(\scanline[157][3] ));
 sg13g2_dfrbp_1 _27039_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2093),
    .D(net3771),
    .Q_N(_12733_),
    .Q(\scanline[157][4] ));
 sg13g2_dfrbp_1 _27040_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2092),
    .D(_00670_),
    .Q_N(_12732_),
    .Q(\scanline[157][5] ));
 sg13g2_dfrbp_1 _27041_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2091),
    .D(_00671_),
    .Q_N(_12731_),
    .Q(\scanline[157][6] ));
 sg13g2_dfrbp_1 _27042_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2090),
    .D(_00672_),
    .Q_N(_12730_),
    .Q(\scanline[156][0] ));
 sg13g2_dfrbp_1 _27043_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2089),
    .D(_00673_),
    .Q_N(_12729_),
    .Q(\scanline[156][1] ));
 sg13g2_dfrbp_1 _27044_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2088),
    .D(_00674_),
    .Q_N(_12728_),
    .Q(\scanline[156][2] ));
 sg13g2_dfrbp_1 _27045_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2087),
    .D(_00675_),
    .Q_N(_12727_),
    .Q(\scanline[156][3] ));
 sg13g2_dfrbp_1 _27046_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2086),
    .D(_00676_),
    .Q_N(_12726_),
    .Q(\scanline[156][4] ));
 sg13g2_dfrbp_1 _27047_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2085),
    .D(_00677_),
    .Q_N(_12725_),
    .Q(\scanline[156][5] ));
 sg13g2_dfrbp_1 _27048_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2084),
    .D(_00678_),
    .Q_N(_12724_),
    .Q(\scanline[156][6] ));
 sg13g2_dfrbp_1 _27049_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2083),
    .D(_00679_),
    .Q_N(_12723_),
    .Q(\scanline[155][0] ));
 sg13g2_dfrbp_1 _27050_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2082),
    .D(_00680_),
    .Q_N(_12722_),
    .Q(\scanline[155][1] ));
 sg13g2_dfrbp_1 _27051_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2081),
    .D(_00681_),
    .Q_N(_12721_),
    .Q(\scanline[155][2] ));
 sg13g2_dfrbp_1 _27052_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2080),
    .D(_00682_),
    .Q_N(_12720_),
    .Q(\scanline[155][3] ));
 sg13g2_dfrbp_1 _27053_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2079),
    .D(_00683_),
    .Q_N(_12719_),
    .Q(\scanline[155][4] ));
 sg13g2_dfrbp_1 _27054_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2078),
    .D(_00684_),
    .Q_N(_12718_),
    .Q(\scanline[155][5] ));
 sg13g2_dfrbp_1 _27055_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2077),
    .D(_00685_),
    .Q_N(_12717_),
    .Q(\scanline[155][6] ));
 sg13g2_dfrbp_1 _27056_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2076),
    .D(_00686_),
    .Q_N(_12716_),
    .Q(\scanline[72][0] ));
 sg13g2_dfrbp_1 _27057_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2075),
    .D(_00687_),
    .Q_N(_12715_),
    .Q(\scanline[72][1] ));
 sg13g2_dfrbp_1 _27058_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2074),
    .D(_00688_),
    .Q_N(_12714_),
    .Q(\scanline[72][2] ));
 sg13g2_dfrbp_1 _27059_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2073),
    .D(_00689_),
    .Q_N(_12713_),
    .Q(\scanline[72][3] ));
 sg13g2_dfrbp_1 _27060_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net2072),
    .D(_00690_),
    .Q_N(_12712_),
    .Q(\scanline[72][4] ));
 sg13g2_dfrbp_1 _27061_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2071),
    .D(_00691_),
    .Q_N(_12711_),
    .Q(\scanline[72][5] ));
 sg13g2_dfrbp_1 _27062_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2070),
    .D(_00692_),
    .Q_N(_12710_),
    .Q(\scanline[72][6] ));
 sg13g2_dfrbp_1 _27063_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2069),
    .D(_00693_),
    .Q_N(_12709_),
    .Q(\scanline[74][0] ));
 sg13g2_dfrbp_1 _27064_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2068),
    .D(_00694_),
    .Q_N(_12708_),
    .Q(\scanline[74][1] ));
 sg13g2_dfrbp_1 _27065_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2067),
    .D(_00695_),
    .Q_N(_12707_),
    .Q(\scanline[74][2] ));
 sg13g2_dfrbp_1 _27066_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2066),
    .D(_00696_),
    .Q_N(_12706_),
    .Q(\scanline[74][3] ));
 sg13g2_dfrbp_1 _27067_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2065),
    .D(_00697_),
    .Q_N(_12705_),
    .Q(\scanline[74][4] ));
 sg13g2_dfrbp_1 _27068_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2064),
    .D(_00698_),
    .Q_N(_12704_),
    .Q(\scanline[74][5] ));
 sg13g2_dfrbp_1 _27069_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2063),
    .D(_00699_),
    .Q_N(_12703_),
    .Q(\scanline[74][6] ));
 sg13g2_dfrbp_1 _27070_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2062),
    .D(_00700_),
    .Q_N(_12702_),
    .Q(\scanline[81][0] ));
 sg13g2_dfrbp_1 _27071_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2061),
    .D(_00701_),
    .Q_N(_12701_),
    .Q(\scanline[81][1] ));
 sg13g2_dfrbp_1 _27072_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2060),
    .D(_00702_),
    .Q_N(_12700_),
    .Q(\scanline[81][2] ));
 sg13g2_dfrbp_1 _27073_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2059),
    .D(_00703_),
    .Q_N(_12699_),
    .Q(\scanline[81][3] ));
 sg13g2_dfrbp_1 _27074_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2058),
    .D(_00704_),
    .Q_N(_12698_),
    .Q(\scanline[81][4] ));
 sg13g2_dfrbp_1 _27075_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net2057),
    .D(_00705_),
    .Q_N(_12697_),
    .Q(\scanline[81][5] ));
 sg13g2_dfrbp_1 _27076_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2056),
    .D(_00706_),
    .Q_N(_12696_),
    .Q(\scanline[81][6] ));
 sg13g2_dfrbp_1 _27077_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2055),
    .D(_00707_),
    .Q_N(_12695_),
    .Q(\scanline[71][0] ));
 sg13g2_dfrbp_1 _27078_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2054),
    .D(_00708_),
    .Q_N(_12694_),
    .Q(\scanline[71][1] ));
 sg13g2_dfrbp_1 _27079_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2053),
    .D(_00709_),
    .Q_N(_12693_),
    .Q(\scanline[71][2] ));
 sg13g2_dfrbp_1 _27080_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2052),
    .D(_00710_),
    .Q_N(_12692_),
    .Q(\scanline[71][3] ));
 sg13g2_dfrbp_1 _27081_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2051),
    .D(_00711_),
    .Q_N(_12691_),
    .Q(\scanline[71][4] ));
 sg13g2_dfrbp_1 _27082_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2050),
    .D(_00712_),
    .Q_N(_12690_),
    .Q(\scanline[71][5] ));
 sg13g2_dfrbp_1 _27083_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2049),
    .D(_00713_),
    .Q_N(_12689_),
    .Q(\scanline[71][6] ));
 sg13g2_dfrbp_1 _27084_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2048),
    .D(_00714_),
    .Q_N(_12688_),
    .Q(\scanline[76][0] ));
 sg13g2_dfrbp_1 _27085_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2047),
    .D(_00715_),
    .Q_N(_12687_),
    .Q(\scanline[76][1] ));
 sg13g2_dfrbp_1 _27086_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2046),
    .D(_00716_),
    .Q_N(_12686_),
    .Q(\scanline[76][2] ));
 sg13g2_dfrbp_1 _27087_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2045),
    .D(_00717_),
    .Q_N(_12685_),
    .Q(\scanline[76][3] ));
 sg13g2_dfrbp_1 _27088_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2044),
    .D(_00718_),
    .Q_N(_12684_),
    .Q(\scanline[76][4] ));
 sg13g2_dfrbp_1 _27089_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2043),
    .D(_00719_),
    .Q_N(_12683_),
    .Q(\scanline[76][5] ));
 sg13g2_dfrbp_1 _27090_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2042),
    .D(_00720_),
    .Q_N(_12682_),
    .Q(\scanline[76][6] ));
 sg13g2_dfrbp_1 _27091_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2041),
    .D(_00721_),
    .Q_N(_12681_),
    .Q(\scanline[49][0] ));
 sg13g2_dfrbp_1 _27092_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2040),
    .D(_00722_),
    .Q_N(_12680_),
    .Q(\scanline[49][1] ));
 sg13g2_dfrbp_1 _27093_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2039),
    .D(_00723_),
    .Q_N(_12679_),
    .Q(\scanline[49][2] ));
 sg13g2_dfrbp_1 _27094_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net2038),
    .D(_00724_),
    .Q_N(_12678_),
    .Q(\scanline[49][3] ));
 sg13g2_dfrbp_1 _27095_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2037),
    .D(_00725_),
    .Q_N(_12677_),
    .Q(\scanline[49][4] ));
 sg13g2_dfrbp_1 _27096_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2036),
    .D(_00726_),
    .Q_N(_12676_),
    .Q(\scanline[49][5] ));
 sg13g2_dfrbp_1 _27097_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1234),
    .D(_00727_),
    .Q_N(_13224_),
    .Q(\scanline[49][6] ));
 sg13g2_dfrbp_1 _27098_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1235),
    .D(_00001_),
    .Q_N(_13225_),
    .Q(\atari2600.ram_data[0] ));
 sg13g2_dfrbp_1 _27099_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1236),
    .D(_00002_),
    .Q_N(_13226_),
    .Q(\atari2600.ram_data[1] ));
 sg13g2_dfrbp_1 _27100_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1237),
    .D(_00003_),
    .Q_N(_13227_),
    .Q(\atari2600.ram_data[2] ));
 sg13g2_dfrbp_1 _27101_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1238),
    .D(_00004_),
    .Q_N(_13228_),
    .Q(\atari2600.ram_data[3] ));
 sg13g2_dfrbp_1 _27102_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1239),
    .D(_00005_),
    .Q_N(_13229_),
    .Q(\atari2600.ram_data[4] ));
 sg13g2_dfrbp_1 _27103_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1240),
    .D(_00006_),
    .Q_N(_13230_),
    .Q(\atari2600.ram_data[5] ));
 sg13g2_dfrbp_1 _27104_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1635),
    .D(_00007_),
    .Q_N(_13231_),
    .Q(\atari2600.ram_data[6] ));
 sg13g2_dfrbp_1 _27105_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net2035),
    .D(_00008_),
    .Q_N(_12675_),
    .Q(\atari2600.ram_data[7] ));
 sg13g2_dfrbp_1 _27106_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2034),
    .D(_00728_),
    .Q_N(_12674_),
    .Q(\scanline[39][0] ));
 sg13g2_dfrbp_1 _27107_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2033),
    .D(_00729_),
    .Q_N(_12673_),
    .Q(\scanline[39][1] ));
 sg13g2_dfrbp_1 _27108_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2032),
    .D(_00730_),
    .Q_N(_12672_),
    .Q(\scanline[39][2] ));
 sg13g2_dfrbp_1 _27109_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2031),
    .D(_00731_),
    .Q_N(_12671_),
    .Q(\scanline[39][3] ));
 sg13g2_dfrbp_1 _27110_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2030),
    .D(_00732_),
    .Q_N(_12670_),
    .Q(\scanline[39][4] ));
 sg13g2_dfrbp_1 _27111_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2029),
    .D(_00733_),
    .Q_N(_12669_),
    .Q(\scanline[39][5] ));
 sg13g2_dfrbp_1 _27112_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2028),
    .D(_00734_),
    .Q_N(_12668_),
    .Q(\scanline[39][6] ));
 sg13g2_dfrbp_1 _27113_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2027),
    .D(_00735_),
    .Q_N(_12667_),
    .Q(\atari2600.ram[21][0] ));
 sg13g2_dfrbp_1 _27114_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net2026),
    .D(_00736_),
    .Q_N(_12666_),
    .Q(\atari2600.ram[21][1] ));
 sg13g2_dfrbp_1 _27115_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net2025),
    .D(_00737_),
    .Q_N(_12665_),
    .Q(\atari2600.ram[21][2] ));
 sg13g2_dfrbp_1 _27116_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2024),
    .D(_00738_),
    .Q_N(_12664_),
    .Q(\atari2600.ram[21][3] ));
 sg13g2_dfrbp_1 _27117_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2023),
    .D(_00739_),
    .Q_N(_12663_),
    .Q(\atari2600.ram[21][4] ));
 sg13g2_dfrbp_1 _27118_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net2022),
    .D(_00740_),
    .Q_N(_12662_),
    .Q(\atari2600.ram[21][5] ));
 sg13g2_dfrbp_1 _27119_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net2021),
    .D(_00741_),
    .Q_N(_12661_),
    .Q(\atari2600.ram[21][6] ));
 sg13g2_dfrbp_1 _27120_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2020),
    .D(_00742_),
    .Q_N(_12660_),
    .Q(\atari2600.ram[21][7] ));
 sg13g2_dfrbp_1 _27121_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2019),
    .D(_00743_),
    .Q_N(_12659_),
    .Q(\scanline[29][0] ));
 sg13g2_dfrbp_1 _27122_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2018),
    .D(_00744_),
    .Q_N(_12658_),
    .Q(\scanline[29][1] ));
 sg13g2_dfrbp_1 _27123_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2017),
    .D(_00745_),
    .Q_N(_12657_),
    .Q(\scanline[29][2] ));
 sg13g2_dfrbp_1 _27124_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2016),
    .D(_00746_),
    .Q_N(_12656_),
    .Q(\scanline[29][3] ));
 sg13g2_dfrbp_1 _27125_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2015),
    .D(_00747_),
    .Q_N(_12655_),
    .Q(\scanline[29][4] ));
 sg13g2_dfrbp_1 _27126_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2014),
    .D(_00748_),
    .Q_N(_12654_),
    .Q(\scanline[29][5] ));
 sg13g2_dfrbp_1 _27127_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net2013),
    .D(_00749_),
    .Q_N(_12653_),
    .Q(\scanline[29][6] ));
 sg13g2_dfrbp_1 _27128_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2012),
    .D(_00750_),
    .Q_N(_12652_),
    .Q(\scanline[19][0] ));
 sg13g2_dfrbp_1 _27129_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net2011),
    .D(_00751_),
    .Q_N(_12651_),
    .Q(\scanline[19][1] ));
 sg13g2_dfrbp_1 _27130_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net2010),
    .D(_00752_),
    .Q_N(_12650_),
    .Q(\scanline[19][2] ));
 sg13g2_dfrbp_1 _27131_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2009),
    .D(_00753_),
    .Q_N(_12649_),
    .Q(\scanline[19][3] ));
 sg13g2_dfrbp_1 _27132_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net2008),
    .D(_00754_),
    .Q_N(_12648_),
    .Q(\scanline[19][4] ));
 sg13g2_dfrbp_1 _27133_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2007),
    .D(_00755_),
    .Q_N(_12647_),
    .Q(\scanline[19][5] ));
 sg13g2_dfrbp_1 _27134_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net2006),
    .D(_00756_),
    .Q_N(_12646_),
    .Q(\scanline[19][6] ));
 sg13g2_dfrbp_1 _27135_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2005),
    .D(_00757_),
    .Q_N(_12645_),
    .Q(\atari2600.ram[9][0] ));
 sg13g2_dfrbp_1 _27136_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net2004),
    .D(_00758_),
    .Q_N(_12644_),
    .Q(\atari2600.ram[9][1] ));
 sg13g2_dfrbp_1 _27137_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2003),
    .D(_00759_),
    .Q_N(_12643_),
    .Q(\atari2600.ram[9][2] ));
 sg13g2_dfrbp_1 _27138_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net2002),
    .D(_00760_),
    .Q_N(_12642_),
    .Q(\atari2600.ram[9][3] ));
 sg13g2_dfrbp_1 _27139_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2001),
    .D(_00761_),
    .Q_N(_12641_),
    .Q(\atari2600.ram[9][4] ));
 sg13g2_dfrbp_1 _27140_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net2000),
    .D(_00762_),
    .Q_N(_12640_),
    .Q(\atari2600.ram[9][5] ));
 sg13g2_dfrbp_1 _27141_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1999),
    .D(_00763_),
    .Q_N(_12639_),
    .Q(\atari2600.ram[9][6] ));
 sg13g2_dfrbp_1 _27142_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1998),
    .D(_00764_),
    .Q_N(_12638_),
    .Q(\atari2600.ram[9][7] ));
 sg13g2_dfrbp_1 _27143_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1997),
    .D(_00765_),
    .Q_N(_12637_),
    .Q(\scanline[57][0] ));
 sg13g2_dfrbp_1 _27144_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1996),
    .D(_00766_),
    .Q_N(_12636_),
    .Q(\scanline[57][1] ));
 sg13g2_dfrbp_1 _27145_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1995),
    .D(_00767_),
    .Q_N(_12635_),
    .Q(\scanline[57][2] ));
 sg13g2_dfrbp_1 _27146_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1994),
    .D(_00768_),
    .Q_N(_12634_),
    .Q(\scanline[57][3] ));
 sg13g2_dfrbp_1 _27147_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1993),
    .D(_00769_),
    .Q_N(_12633_),
    .Q(\scanline[57][4] ));
 sg13g2_dfrbp_1 _27148_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1992),
    .D(_00770_),
    .Q_N(_12632_),
    .Q(\scanline[57][5] ));
 sg13g2_dfrbp_1 _27149_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1991),
    .D(_00771_),
    .Q_N(_12631_),
    .Q(\scanline[57][6] ));
 sg13g2_dfrbp_1 _27150_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1990),
    .D(_00772_),
    .Q_N(_12630_),
    .Q(\scanline[110][0] ));
 sg13g2_dfrbp_1 _27151_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1989),
    .D(_00773_),
    .Q_N(_12629_),
    .Q(\scanline[110][1] ));
 sg13g2_dfrbp_1 _27152_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1988),
    .D(_00774_),
    .Q_N(_12628_),
    .Q(\scanline[110][2] ));
 sg13g2_dfrbp_1 _27153_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1987),
    .D(_00775_),
    .Q_N(_12627_),
    .Q(\scanline[110][3] ));
 sg13g2_dfrbp_1 _27154_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1986),
    .D(_00776_),
    .Q_N(_12626_),
    .Q(\scanline[110][4] ));
 sg13g2_dfrbp_1 _27155_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1985),
    .D(_00777_),
    .Q_N(_12625_),
    .Q(\scanline[110][5] ));
 sg13g2_dfrbp_1 _27156_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1984),
    .D(_00778_),
    .Q_N(_12624_),
    .Q(\scanline[110][6] ));
 sg13g2_dfrbp_1 _27157_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1983),
    .D(_00779_),
    .Q_N(_12623_),
    .Q(\scanline[143][0] ));
 sg13g2_dfrbp_1 _27158_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1982),
    .D(_00780_),
    .Q_N(_12622_),
    .Q(\scanline[143][1] ));
 sg13g2_dfrbp_1 _27159_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1981),
    .D(_00781_),
    .Q_N(_12621_),
    .Q(\scanline[143][2] ));
 sg13g2_dfrbp_1 _27160_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1980),
    .D(_00782_),
    .Q_N(_12620_),
    .Q(\scanline[143][3] ));
 sg13g2_dfrbp_1 _27161_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1979),
    .D(_00783_),
    .Q_N(_12619_),
    .Q(\scanline[143][4] ));
 sg13g2_dfrbp_1 _27162_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1978),
    .D(_00784_),
    .Q_N(_12618_),
    .Q(\scanline[143][5] ));
 sg13g2_dfrbp_1 _27163_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1977),
    .D(_00785_),
    .Q_N(_12617_),
    .Q(\scanline[143][6] ));
 sg13g2_dfrbp_1 _27164_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1976),
    .D(_00786_),
    .Q_N(_12616_),
    .Q(\scanline[10][0] ));
 sg13g2_dfrbp_1 _27165_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1975),
    .D(_00787_),
    .Q_N(_12615_),
    .Q(\scanline[10][1] ));
 sg13g2_dfrbp_1 _27166_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1974),
    .D(_00788_),
    .Q_N(_12614_),
    .Q(\scanline[10][2] ));
 sg13g2_dfrbp_1 _27167_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1973),
    .D(_00789_),
    .Q_N(_12613_),
    .Q(\scanline[10][3] ));
 sg13g2_dfrbp_1 _27168_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1972),
    .D(_00790_),
    .Q_N(_12612_),
    .Q(\scanline[10][4] ));
 sg13g2_dfrbp_1 _27169_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1971),
    .D(_00791_),
    .Q_N(_12611_),
    .Q(\scanline[10][5] ));
 sg13g2_dfrbp_1 _27170_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1970),
    .D(_00792_),
    .Q_N(_12610_),
    .Q(\scanline[10][6] ));
 sg13g2_dfrbp_1 _27171_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1969),
    .D(_00793_),
    .Q_N(_12609_),
    .Q(\scanline[108][0] ));
 sg13g2_dfrbp_1 _27172_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1968),
    .D(_00794_),
    .Q_N(_12608_),
    .Q(\scanline[108][1] ));
 sg13g2_dfrbp_1 _27173_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1967),
    .D(_00795_),
    .Q_N(_12607_),
    .Q(\scanline[108][2] ));
 sg13g2_dfrbp_1 _27174_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1966),
    .D(_00796_),
    .Q_N(_12606_),
    .Q(\scanline[108][3] ));
 sg13g2_dfrbp_1 _27175_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1965),
    .D(_00797_),
    .Q_N(_12605_),
    .Q(\scanline[108][4] ));
 sg13g2_dfrbp_1 _27176_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1964),
    .D(_00798_),
    .Q_N(_12604_),
    .Q(\scanline[108][5] ));
 sg13g2_dfrbp_1 _27177_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1963),
    .D(_00799_),
    .Q_N(_12603_),
    .Q(\scanline[108][6] ));
 sg13g2_dfrbp_1 _27178_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1962),
    .D(_00800_),
    .Q_N(_12602_),
    .Q(\scanline[142][0] ));
 sg13g2_dfrbp_1 _27179_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1961),
    .D(_00801_),
    .Q_N(_12601_),
    .Q(\scanline[142][1] ));
 sg13g2_dfrbp_1 _27180_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1960),
    .D(_00802_),
    .Q_N(_12600_),
    .Q(\scanline[142][2] ));
 sg13g2_dfrbp_1 _27181_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1959),
    .D(_00803_),
    .Q_N(_12599_),
    .Q(\scanline[142][3] ));
 sg13g2_dfrbp_1 _27182_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1958),
    .D(_00804_),
    .Q_N(_12598_),
    .Q(\scanline[142][4] ));
 sg13g2_dfrbp_1 _27183_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1957),
    .D(_00805_),
    .Q_N(_12597_),
    .Q(\scanline[142][5] ));
 sg13g2_dfrbp_1 _27184_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1956),
    .D(_00806_),
    .Q_N(_12596_),
    .Q(\scanline[142][6] ));
 sg13g2_dfrbp_1 _27185_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1955),
    .D(_00807_),
    .Q_N(_12595_),
    .Q(\scanline[107][0] ));
 sg13g2_dfrbp_1 _27186_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1954),
    .D(_00808_),
    .Q_N(_12594_),
    .Q(\scanline[107][1] ));
 sg13g2_dfrbp_1 _27187_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1953),
    .D(_00809_),
    .Q_N(_12593_),
    .Q(\scanline[107][2] ));
 sg13g2_dfrbp_1 _27188_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1952),
    .D(_00810_),
    .Q_N(_12592_),
    .Q(\scanline[107][3] ));
 sg13g2_dfrbp_1 _27189_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1951),
    .D(_00811_),
    .Q_N(_12591_),
    .Q(\scanline[107][4] ));
 sg13g2_dfrbp_1 _27190_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1950),
    .D(_00812_),
    .Q_N(_12590_),
    .Q(\scanline[107][5] ));
 sg13g2_dfrbp_1 _27191_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1949),
    .D(_00813_),
    .Q_N(_12589_),
    .Q(\scanline[107][6] ));
 sg13g2_dfrbp_1 _27192_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1948),
    .D(_00814_),
    .Q_N(_12588_),
    .Q(\scanline[106][0] ));
 sg13g2_dfrbp_1 _27193_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1947),
    .D(_00815_),
    .Q_N(_12587_),
    .Q(\scanline[106][1] ));
 sg13g2_dfrbp_1 _27194_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1946),
    .D(_00816_),
    .Q_N(_12586_),
    .Q(\scanline[106][2] ));
 sg13g2_dfrbp_1 _27195_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1945),
    .D(_00817_),
    .Q_N(_12585_),
    .Q(\scanline[106][3] ));
 sg13g2_dfrbp_1 _27196_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1944),
    .D(_00818_),
    .Q_N(_12584_),
    .Q(\scanline[106][4] ));
 sg13g2_dfrbp_1 _27197_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1943),
    .D(_00819_),
    .Q_N(_12583_),
    .Q(\scanline[106][5] ));
 sg13g2_dfrbp_1 _27198_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1942),
    .D(_00820_),
    .Q_N(_12582_),
    .Q(\scanline[106][6] ));
 sg13g2_dfrbp_1 _27199_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1941),
    .D(_00821_),
    .Q_N(_12581_),
    .Q(\scanline[141][0] ));
 sg13g2_dfrbp_1 _27200_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1940),
    .D(_00822_),
    .Q_N(_12580_),
    .Q(\scanline[141][1] ));
 sg13g2_dfrbp_1 _27201_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1939),
    .D(_00823_),
    .Q_N(_12579_),
    .Q(\scanline[141][2] ));
 sg13g2_dfrbp_1 _27202_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1938),
    .D(_00824_),
    .Q_N(_12578_),
    .Q(\scanline[141][3] ));
 sg13g2_dfrbp_1 _27203_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1937),
    .D(_00825_),
    .Q_N(_12577_),
    .Q(\scanline[141][4] ));
 sg13g2_dfrbp_1 _27204_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1936),
    .D(_00826_),
    .Q_N(_12576_),
    .Q(\scanline[141][5] ));
 sg13g2_dfrbp_1 _27205_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1935),
    .D(_00827_),
    .Q_N(_12575_),
    .Q(\scanline[141][6] ));
 sg13g2_dfrbp_1 _27206_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1934),
    .D(_00828_),
    .Q_N(_12574_),
    .Q(\scanline[105][0] ));
 sg13g2_dfrbp_1 _27207_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1933),
    .D(_00829_),
    .Q_N(_12573_),
    .Q(\scanline[105][1] ));
 sg13g2_dfrbp_1 _27208_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1932),
    .D(_00830_),
    .Q_N(_12572_),
    .Q(\scanline[105][2] ));
 sg13g2_dfrbp_1 _27209_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1931),
    .D(_00831_),
    .Q_N(_12571_),
    .Q(\scanline[105][3] ));
 sg13g2_dfrbp_1 _27210_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1930),
    .D(_00832_),
    .Q_N(_12570_),
    .Q(\scanline[105][4] ));
 sg13g2_dfrbp_1 _27211_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1929),
    .D(_00833_),
    .Q_N(_12569_),
    .Q(\scanline[105][5] ));
 sg13g2_dfrbp_1 _27212_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1928),
    .D(_00834_),
    .Q_N(_12568_),
    .Q(\scanline[105][6] ));
 sg13g2_dfrbp_1 _27213_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1927),
    .D(_00835_),
    .Q_N(_12567_),
    .Q(\scanline[104][0] ));
 sg13g2_dfrbp_1 _27214_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1926),
    .D(_00836_),
    .Q_N(_12566_),
    .Q(\scanline[104][1] ));
 sg13g2_dfrbp_1 _27215_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1925),
    .D(_00837_),
    .Q_N(_12565_),
    .Q(\scanline[104][2] ));
 sg13g2_dfrbp_1 _27216_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1924),
    .D(_00838_),
    .Q_N(_12564_),
    .Q(\scanline[104][3] ));
 sg13g2_dfrbp_1 _27217_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1923),
    .D(_00839_),
    .Q_N(_12563_),
    .Q(\scanline[104][4] ));
 sg13g2_dfrbp_1 _27218_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1922),
    .D(_00840_),
    .Q_N(_12562_),
    .Q(\scanline[104][5] ));
 sg13g2_dfrbp_1 _27219_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1921),
    .D(_00841_),
    .Q_N(_12561_),
    .Q(\scanline[104][6] ));
 sg13g2_dfrbp_1 _27220_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1920),
    .D(_00842_),
    .Q_N(_12560_),
    .Q(\scanline[140][0] ));
 sg13g2_dfrbp_1 _27221_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1919),
    .D(_00843_),
    .Q_N(_12559_),
    .Q(\scanline[140][1] ));
 sg13g2_dfrbp_1 _27222_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1918),
    .D(_00844_),
    .Q_N(_12558_),
    .Q(\scanline[140][2] ));
 sg13g2_dfrbp_1 _27223_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1917),
    .D(_00845_),
    .Q_N(_12557_),
    .Q(\scanline[140][3] ));
 sg13g2_dfrbp_1 _27224_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1916),
    .D(_00846_),
    .Q_N(_12556_),
    .Q(\scanline[140][4] ));
 sg13g2_dfrbp_1 _27225_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1915),
    .D(_00847_),
    .Q_N(_12555_),
    .Q(\scanline[140][5] ));
 sg13g2_dfrbp_1 _27226_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1914),
    .D(_00848_),
    .Q_N(_12554_),
    .Q(\scanline[140][6] ));
 sg13g2_dfrbp_1 _27227_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1913),
    .D(_00849_),
    .Q_N(_12553_),
    .Q(\scanline[103][0] ));
 sg13g2_dfrbp_1 _27228_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1912),
    .D(_00850_),
    .Q_N(_12552_),
    .Q(\scanline[103][1] ));
 sg13g2_dfrbp_1 _27229_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1911),
    .D(_00851_),
    .Q_N(_12551_),
    .Q(\scanline[103][2] ));
 sg13g2_dfrbp_1 _27230_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1910),
    .D(_00852_),
    .Q_N(_12550_),
    .Q(\scanline[103][3] ));
 sg13g2_dfrbp_1 _27231_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1909),
    .D(_00853_),
    .Q_N(_12549_),
    .Q(\scanline[103][4] ));
 sg13g2_dfrbp_1 _27232_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1908),
    .D(_00854_),
    .Q_N(_12548_),
    .Q(\scanline[103][5] ));
 sg13g2_dfrbp_1 _27233_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1907),
    .D(_00855_),
    .Q_N(_12547_),
    .Q(\scanline[103][6] ));
 sg13g2_dfrbp_1 _27234_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1906),
    .D(_00856_),
    .Q_N(_12546_),
    .Q(\scanline[102][0] ));
 sg13g2_dfrbp_1 _27235_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1905),
    .D(_00857_),
    .Q_N(_12545_),
    .Q(\scanline[102][1] ));
 sg13g2_dfrbp_1 _27236_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1904),
    .D(_00858_),
    .Q_N(_12544_),
    .Q(\scanline[102][2] ));
 sg13g2_dfrbp_1 _27237_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1903),
    .D(_00859_),
    .Q_N(_12543_),
    .Q(\scanline[102][3] ));
 sg13g2_dfrbp_1 _27238_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1902),
    .D(_00860_),
    .Q_N(_12542_),
    .Q(\scanline[102][4] ));
 sg13g2_dfrbp_1 _27239_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1901),
    .D(_00861_),
    .Q_N(_12541_),
    .Q(\scanline[102][5] ));
 sg13g2_dfrbp_1 _27240_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1900),
    .D(_00862_),
    .Q_N(_12540_),
    .Q(\scanline[102][6] ));
 sg13g2_dfrbp_1 _27241_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1899),
    .D(_00863_),
    .Q_N(_12539_),
    .Q(\scanline[13][0] ));
 sg13g2_dfrbp_1 _27242_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1898),
    .D(_00864_),
    .Q_N(_12538_),
    .Q(\scanline[13][1] ));
 sg13g2_dfrbp_1 _27243_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1897),
    .D(_00865_),
    .Q_N(_12537_),
    .Q(\scanline[13][2] ));
 sg13g2_dfrbp_1 _27244_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1896),
    .D(_00866_),
    .Q_N(_12536_),
    .Q(\scanline[13][3] ));
 sg13g2_dfrbp_1 _27245_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1895),
    .D(_00867_),
    .Q_N(_12535_),
    .Q(\scanline[13][4] ));
 sg13g2_dfrbp_1 _27246_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1894),
    .D(_00868_),
    .Q_N(_12534_),
    .Q(\scanline[13][5] ));
 sg13g2_dfrbp_1 _27247_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1893),
    .D(_00869_),
    .Q_N(_12533_),
    .Q(\scanline[13][6] ));
 sg13g2_dfrbp_1 _27248_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1892),
    .D(_00870_),
    .Q_N(_12532_),
    .Q(\scanline[101][0] ));
 sg13g2_dfrbp_1 _27249_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1891),
    .D(_00871_),
    .Q_N(_12531_),
    .Q(\scanline[101][1] ));
 sg13g2_dfrbp_1 _27250_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1890),
    .D(_00872_),
    .Q_N(_12530_),
    .Q(\scanline[101][2] ));
 sg13g2_dfrbp_1 _27251_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1889),
    .D(_00873_),
    .Q_N(_12529_),
    .Q(\scanline[101][3] ));
 sg13g2_dfrbp_1 _27252_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1888),
    .D(_00874_),
    .Q_N(_12528_),
    .Q(\scanline[101][4] ));
 sg13g2_dfrbp_1 _27253_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1887),
    .D(_00875_),
    .Q_N(_12527_),
    .Q(\scanline[101][5] ));
 sg13g2_dfrbp_1 _27254_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1886),
    .D(_00876_),
    .Q_N(_12526_),
    .Q(\scanline[101][6] ));
 sg13g2_dfrbp_1 _27255_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1885),
    .D(_00877_),
    .Q_N(_12525_),
    .Q(\scanline[100][0] ));
 sg13g2_dfrbp_1 _27256_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1884),
    .D(_00878_),
    .Q_N(_12524_),
    .Q(\scanline[100][1] ));
 sg13g2_dfrbp_1 _27257_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1883),
    .D(_00879_),
    .Q_N(_12523_),
    .Q(\scanline[100][2] ));
 sg13g2_dfrbp_1 _27258_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1882),
    .D(_00880_),
    .Q_N(_12522_),
    .Q(\scanline[100][3] ));
 sg13g2_dfrbp_1 _27259_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1881),
    .D(_00881_),
    .Q_N(_12521_),
    .Q(\scanline[100][4] ));
 sg13g2_dfrbp_1 _27260_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1880),
    .D(_00882_),
    .Q_N(_12520_),
    .Q(\scanline[100][5] ));
 sg13g2_dfrbp_1 _27261_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1879),
    .D(_00883_),
    .Q_N(_12519_),
    .Q(\scanline[100][6] ));
 sg13g2_dfrbp_1 _27262_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1878),
    .D(_00884_),
    .Q_N(_12518_),
    .Q(\scanline[138][0] ));
 sg13g2_dfrbp_1 _27263_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1877),
    .D(_00885_),
    .Q_N(_12517_),
    .Q(\scanline[138][1] ));
 sg13g2_dfrbp_1 _27264_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1876),
    .D(_00886_),
    .Q_N(_12516_),
    .Q(\scanline[138][2] ));
 sg13g2_dfrbp_1 _27265_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1875),
    .D(_00887_),
    .Q_N(_12515_),
    .Q(\scanline[138][3] ));
 sg13g2_dfrbp_1 _27266_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1874),
    .D(_00888_),
    .Q_N(_12514_),
    .Q(\scanline[138][4] ));
 sg13g2_dfrbp_1 _27267_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1873),
    .D(_00889_),
    .Q_N(_12513_),
    .Q(\scanline[138][5] ));
 sg13g2_dfrbp_1 _27268_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1872),
    .D(_00890_),
    .Q_N(_12512_),
    .Q(\scanline[138][6] ));
 sg13g2_dfrbp_1 _27269_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1871),
    .D(_00891_),
    .Q_N(_12511_),
    .Q(\scanline[0][0] ));
 sg13g2_dfrbp_1 _27270_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1870),
    .D(_00892_),
    .Q_N(_12510_),
    .Q(\scanline[0][1] ));
 sg13g2_dfrbp_1 _27271_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1869),
    .D(_00893_),
    .Q_N(_12509_),
    .Q(\scanline[0][2] ));
 sg13g2_dfrbp_1 _27272_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1868),
    .D(_00894_),
    .Q_N(_12508_),
    .Q(\scanline[0][3] ));
 sg13g2_dfrbp_1 _27273_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1867),
    .D(_00895_),
    .Q_N(_12507_),
    .Q(\scanline[0][4] ));
 sg13g2_dfrbp_1 _27274_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1866),
    .D(_00896_),
    .Q_N(_12506_),
    .Q(\scanline[0][5] ));
 sg13g2_dfrbp_1 _27275_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1865),
    .D(_00897_),
    .Q_N(_12505_),
    .Q(\scanline[0][6] ));
 sg13g2_dfrbp_1 _27276_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1864),
    .D(_00898_),
    .Q_N(_12504_),
    .Q(\scanline[98][0] ));
 sg13g2_dfrbp_1 _27277_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1863),
    .D(_00899_),
    .Q_N(_12503_),
    .Q(\scanline[98][1] ));
 sg13g2_dfrbp_1 _27278_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1862),
    .D(_00900_),
    .Q_N(_12502_),
    .Q(\scanline[98][2] ));
 sg13g2_dfrbp_1 _27279_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1861),
    .D(_00901_),
    .Q_N(_12501_),
    .Q(\scanline[98][3] ));
 sg13g2_dfrbp_1 _27280_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1860),
    .D(_00902_),
    .Q_N(_12500_),
    .Q(\scanline[98][4] ));
 sg13g2_dfrbp_1 _27281_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1859),
    .D(_00903_),
    .Q_N(_12499_),
    .Q(\scanline[98][5] ));
 sg13g2_dfrbp_1 _27282_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1858),
    .D(_00904_),
    .Q_N(_12498_),
    .Q(\scanline[98][6] ));
 sg13g2_dfrbp_1 _27283_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1857),
    .D(_00905_),
    .Q_N(_12497_),
    .Q(\scanline[137][0] ));
 sg13g2_dfrbp_1 _27284_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1856),
    .D(_00906_),
    .Q_N(_12496_),
    .Q(\scanline[137][1] ));
 sg13g2_dfrbp_1 _27285_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1855),
    .D(_00907_),
    .Q_N(_12495_),
    .Q(\scanline[137][2] ));
 sg13g2_dfrbp_1 _27286_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1854),
    .D(_00908_),
    .Q_N(_12494_),
    .Q(\scanline[137][3] ));
 sg13g2_dfrbp_1 _27287_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1853),
    .D(_00909_),
    .Q_N(_12493_),
    .Q(\scanline[137][4] ));
 sg13g2_dfrbp_1 _27288_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1852),
    .D(_00910_),
    .Q_N(_12492_),
    .Q(\scanline[137][5] ));
 sg13g2_dfrbp_1 _27289_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1851),
    .D(_00911_),
    .Q_N(_12491_),
    .Q(\scanline[137][6] ));
 sg13g2_dfrbp_1 _27290_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1850),
    .D(_00912_),
    .Q_N(_12490_),
    .Q(\scanline[97][0] ));
 sg13g2_dfrbp_1 _27291_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1849),
    .D(_00913_),
    .Q_N(_12489_),
    .Q(\scanline[97][1] ));
 sg13g2_dfrbp_1 _27292_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1848),
    .D(_00914_),
    .Q_N(_12488_),
    .Q(\scanline[97][2] ));
 sg13g2_dfrbp_1 _27293_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1847),
    .D(_00915_),
    .Q_N(_12487_),
    .Q(\scanline[97][3] ));
 sg13g2_dfrbp_1 _27294_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1846),
    .D(_00916_),
    .Q_N(_12486_),
    .Q(\scanline[97][4] ));
 sg13g2_dfrbp_1 _27295_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1845),
    .D(_00917_),
    .Q_N(_12485_),
    .Q(\scanline[97][5] ));
 sg13g2_dfrbp_1 _27296_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1844),
    .D(_00918_),
    .Q_N(_12484_),
    .Q(\scanline[97][6] ));
 sg13g2_dfrbp_1 _27297_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1843),
    .D(_00919_),
    .Q_N(_12483_),
    .Q(\scanline[96][0] ));
 sg13g2_dfrbp_1 _27298_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1842),
    .D(_00920_),
    .Q_N(_12482_),
    .Q(\scanline[96][1] ));
 sg13g2_dfrbp_1 _27299_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1841),
    .D(_00921_),
    .Q_N(_12481_),
    .Q(\scanline[96][2] ));
 sg13g2_dfrbp_1 _27300_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1840),
    .D(_00922_),
    .Q_N(_12480_),
    .Q(\scanline[96][3] ));
 sg13g2_dfrbp_1 _27301_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1839),
    .D(_00923_),
    .Q_N(_12479_),
    .Q(\scanline[96][4] ));
 sg13g2_dfrbp_1 _27302_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1838),
    .D(_00924_),
    .Q_N(_12478_),
    .Q(\scanline[96][5] ));
 sg13g2_dfrbp_1 _27303_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1837),
    .D(_00925_),
    .Q_N(_12477_),
    .Q(\scanline[96][6] ));
 sg13g2_dfrbp_1 _27304_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1836),
    .D(_00926_),
    .Q_N(_12476_),
    .Q(\scanline[136][0] ));
 sg13g2_dfrbp_1 _27305_ (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1835),
    .D(_00927_),
    .Q_N(_12475_),
    .Q(\scanline[136][1] ));
 sg13g2_dfrbp_1 _27306_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1834),
    .D(_00928_),
    .Q_N(_12474_),
    .Q(\scanline[136][2] ));
 sg13g2_dfrbp_1 _27307_ (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1833),
    .D(_00929_),
    .Q_N(_12473_),
    .Q(\scanline[136][3] ));
 sg13g2_dfrbp_1 _27308_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1832),
    .D(_00930_),
    .Q_N(_12472_),
    .Q(\scanline[136][4] ));
 sg13g2_dfrbp_1 _27309_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1831),
    .D(_00931_),
    .Q_N(_12471_),
    .Q(\scanline[136][5] ));
 sg13g2_dfrbp_1 _27310_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1830),
    .D(_00932_),
    .Q_N(_12470_),
    .Q(\scanline[136][6] ));
 sg13g2_dfrbp_1 _27311_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1829),
    .D(_00933_),
    .Q_N(_12469_),
    .Q(\scanline[95][0] ));
 sg13g2_dfrbp_1 _27312_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1828),
    .D(_00934_),
    .Q_N(_12468_),
    .Q(\scanline[95][1] ));
 sg13g2_dfrbp_1 _27313_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1827),
    .D(_00935_),
    .Q_N(_12467_),
    .Q(\scanline[95][2] ));
 sg13g2_dfrbp_1 _27314_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1826),
    .D(_00936_),
    .Q_N(_12466_),
    .Q(\scanline[95][3] ));
 sg13g2_dfrbp_1 _27315_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1825),
    .D(_00937_),
    .Q_N(_12465_),
    .Q(\scanline[95][4] ));
 sg13g2_dfrbp_1 _27316_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1824),
    .D(_00938_),
    .Q_N(_12464_),
    .Q(\scanline[95][5] ));
 sg13g2_dfrbp_1 _27317_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1823),
    .D(_00939_),
    .Q_N(_12463_),
    .Q(\scanline[95][6] ));
 sg13g2_dfrbp_1 _27318_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1822),
    .D(_00940_),
    .Q_N(_12462_),
    .Q(\scanline[94][0] ));
 sg13g2_dfrbp_1 _27319_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1821),
    .D(_00941_),
    .Q_N(_12461_),
    .Q(\scanline[94][1] ));
 sg13g2_dfrbp_1 _27320_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1820),
    .D(_00942_),
    .Q_N(_12460_),
    .Q(\scanline[94][2] ));
 sg13g2_dfrbp_1 _27321_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1819),
    .D(_00943_),
    .Q_N(_12459_),
    .Q(\scanline[94][3] ));
 sg13g2_dfrbp_1 _27322_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1818),
    .D(_00944_),
    .Q_N(_12458_),
    .Q(\scanline[94][4] ));
 sg13g2_dfrbp_1 _27323_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1817),
    .D(_00945_),
    .Q_N(_12457_),
    .Q(\scanline[94][5] ));
 sg13g2_dfrbp_1 _27324_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1816),
    .D(_00946_),
    .Q_N(_12456_),
    .Q(\scanline[94][6] ));
 sg13g2_dfrbp_1 _27325_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1815),
    .D(_00947_),
    .Q_N(_12455_),
    .Q(\scanline[135][0] ));
 sg13g2_dfrbp_1 _27326_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1814),
    .D(_00948_),
    .Q_N(_12454_),
    .Q(\scanline[135][1] ));
 sg13g2_dfrbp_1 _27327_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1813),
    .D(_00949_),
    .Q_N(_12453_),
    .Q(\scanline[135][2] ));
 sg13g2_dfrbp_1 _27328_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1812),
    .D(_00950_),
    .Q_N(_12452_),
    .Q(\scanline[135][3] ));
 sg13g2_dfrbp_1 _27329_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1811),
    .D(_00951_),
    .Q_N(_12451_),
    .Q(\scanline[135][4] ));
 sg13g2_dfrbp_1 _27330_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1810),
    .D(_00952_),
    .Q_N(_12450_),
    .Q(\scanline[135][5] ));
 sg13g2_dfrbp_1 _27331_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1809),
    .D(_00953_),
    .Q_N(_12449_),
    .Q(\scanline[135][6] ));
 sg13g2_dfrbp_1 _27332_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1808),
    .D(_00954_),
    .Q_N(_12448_),
    .Q(\scanline[93][0] ));
 sg13g2_dfrbp_1 _27333_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1807),
    .D(_00955_),
    .Q_N(_12447_),
    .Q(\scanline[93][1] ));
 sg13g2_dfrbp_1 _27334_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1806),
    .D(_00956_),
    .Q_N(_12446_),
    .Q(\scanline[93][2] ));
 sg13g2_dfrbp_1 _27335_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1805),
    .D(_00957_),
    .Q_N(_12445_),
    .Q(\scanline[93][3] ));
 sg13g2_dfrbp_1 _27336_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1804),
    .D(_00958_),
    .Q_N(_12444_),
    .Q(\scanline[93][4] ));
 sg13g2_dfrbp_1 _27337_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1803),
    .D(_00959_),
    .Q_N(_12443_),
    .Q(\scanline[93][5] ));
 sg13g2_dfrbp_1 _27338_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1802),
    .D(_00960_),
    .Q_N(_12442_),
    .Q(\scanline[93][6] ));
 sg13g2_dfrbp_1 _27339_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1801),
    .D(_00961_),
    .Q_N(_12441_),
    .Q(\scanline[92][0] ));
 sg13g2_dfrbp_1 _27340_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1800),
    .D(_00962_),
    .Q_N(_12440_),
    .Q(\scanline[92][1] ));
 sg13g2_dfrbp_1 _27341_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1799),
    .D(_00963_),
    .Q_N(_12439_),
    .Q(\scanline[92][2] ));
 sg13g2_dfrbp_1 _27342_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1798),
    .D(_00964_),
    .Q_N(_12438_),
    .Q(\scanline[92][3] ));
 sg13g2_dfrbp_1 _27343_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1797),
    .D(_00965_),
    .Q_N(_12437_),
    .Q(\scanline[92][4] ));
 sg13g2_dfrbp_1 _27344_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1796),
    .D(_00966_),
    .Q_N(_12436_),
    .Q(\scanline[92][5] ));
 sg13g2_dfrbp_1 _27345_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1795),
    .D(_00967_),
    .Q_N(_12435_),
    .Q(\scanline[92][6] ));
 sg13g2_dfrbp_1 _27346_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1794),
    .D(_00968_),
    .Q_N(_12434_),
    .Q(\scanline[134][0] ));
 sg13g2_dfrbp_1 _27347_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1793),
    .D(_00969_),
    .Q_N(_12433_),
    .Q(\scanline[134][1] ));
 sg13g2_dfrbp_1 _27348_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1792),
    .D(_00970_),
    .Q_N(_12432_),
    .Q(\scanline[134][2] ));
 sg13g2_dfrbp_1 _27349_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1791),
    .D(_00971_),
    .Q_N(_12431_),
    .Q(\scanline[134][3] ));
 sg13g2_dfrbp_1 _27350_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1790),
    .D(_00972_),
    .Q_N(_12430_),
    .Q(\scanline[134][4] ));
 sg13g2_dfrbp_1 _27351_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1789),
    .D(_00973_),
    .Q_N(_12429_),
    .Q(\scanline[134][5] ));
 sg13g2_dfrbp_1 _27352_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1788),
    .D(_00974_),
    .Q_N(_12428_),
    .Q(\scanline[134][6] ));
 sg13g2_dfrbp_1 _27353_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1787),
    .D(_00975_),
    .Q_N(_12427_),
    .Q(\scanline[91][0] ));
 sg13g2_dfrbp_1 _27354_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1786),
    .D(_00976_),
    .Q_N(_12426_),
    .Q(\scanline[91][1] ));
 sg13g2_dfrbp_1 _27355_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1785),
    .D(_00977_),
    .Q_N(_12425_),
    .Q(\scanline[91][2] ));
 sg13g2_dfrbp_1 _27356_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1782),
    .D(_00978_),
    .Q_N(_12424_),
    .Q(\scanline[91][3] ));
 sg13g2_dfrbp_1 _27357_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1781),
    .D(_00979_),
    .Q_N(_12423_),
    .Q(\scanline[91][4] ));
 sg13g2_dfrbp_1 _27358_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1780),
    .D(_00980_),
    .Q_N(_12422_),
    .Q(\scanline[91][5] ));
 sg13g2_dfrbp_1 _27359_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1779),
    .D(_00981_),
    .Q_N(_12421_),
    .Q(\scanline[91][6] ));
 sg13g2_dfrbp_1 _27360_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1778),
    .D(_00982_),
    .Q_N(_12420_),
    .Q(\scanline[90][0] ));
 sg13g2_dfrbp_1 _27361_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1777),
    .D(_00983_),
    .Q_N(_12419_),
    .Q(\scanline[90][1] ));
 sg13g2_dfrbp_1 _27362_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1776),
    .D(_00984_),
    .Q_N(_12418_),
    .Q(\scanline[90][2] ));
 sg13g2_dfrbp_1 _27363_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1775),
    .D(_00985_),
    .Q_N(_12417_),
    .Q(\scanline[90][3] ));
 sg13g2_dfrbp_1 _27364_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1774),
    .D(_00986_),
    .Q_N(_12416_),
    .Q(\scanline[90][4] ));
 sg13g2_dfrbp_1 _27365_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1773),
    .D(_00987_),
    .Q_N(_12415_),
    .Q(\scanline[90][5] ));
 sg13g2_dfrbp_1 _27366_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1772),
    .D(_00988_),
    .Q_N(_12414_),
    .Q(\scanline[90][6] ));
 sg13g2_dfrbp_1 _27367_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1771),
    .D(_00989_),
    .Q_N(_12413_),
    .Q(\scanline[133][0] ));
 sg13g2_dfrbp_1 _27368_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1770),
    .D(_00990_),
    .Q_N(_12412_),
    .Q(\scanline[133][1] ));
 sg13g2_dfrbp_1 _27369_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1769),
    .D(_00991_),
    .Q_N(_12411_),
    .Q(\scanline[133][2] ));
 sg13g2_dfrbp_1 _27370_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1768),
    .D(_00992_),
    .Q_N(_12410_),
    .Q(\scanline[133][3] ));
 sg13g2_dfrbp_1 _27371_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1767),
    .D(_00993_),
    .Q_N(_12409_),
    .Q(\scanline[133][4] ));
 sg13g2_dfrbp_1 _27372_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1766),
    .D(_00994_),
    .Q_N(_12408_),
    .Q(\scanline[133][5] ));
 sg13g2_dfrbp_1 _27373_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1765),
    .D(_00995_),
    .Q_N(_12407_),
    .Q(\scanline[133][6] ));
 sg13g2_dfrbp_1 _27374_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1764),
    .D(_00996_),
    .Q_N(_12406_),
    .Q(\scanline[8][0] ));
 sg13g2_dfrbp_1 _27375_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1763),
    .D(_00997_),
    .Q_N(_12405_),
    .Q(\scanline[8][1] ));
 sg13g2_dfrbp_1 _27376_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1762),
    .D(_00998_),
    .Q_N(_12404_),
    .Q(\scanline[8][2] ));
 sg13g2_dfrbp_1 _27377_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1761),
    .D(_00999_),
    .Q_N(_12403_),
    .Q(\scanline[8][3] ));
 sg13g2_dfrbp_1 _27378_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1760),
    .D(_01000_),
    .Q_N(_12402_),
    .Q(\scanline[8][4] ));
 sg13g2_dfrbp_1 _27379_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1759),
    .D(_01001_),
    .Q_N(_12401_),
    .Q(\scanline[8][5] ));
 sg13g2_dfrbp_1 _27380_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1758),
    .D(_01002_),
    .Q_N(_12400_),
    .Q(\scanline[8][6] ));
 sg13g2_dfrbp_1 _27381_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1757),
    .D(_01003_),
    .Q_N(_12399_),
    .Q(\scanline[88][0] ));
 sg13g2_dfrbp_1 _27382_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1756),
    .D(_01004_),
    .Q_N(_12398_),
    .Q(\scanline[88][1] ));
 sg13g2_dfrbp_1 _27383_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1755),
    .D(_01005_),
    .Q_N(_12397_),
    .Q(\scanline[88][2] ));
 sg13g2_dfrbp_1 _27384_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1754),
    .D(_01006_),
    .Q_N(_12396_),
    .Q(\scanline[88][3] ));
 sg13g2_dfrbp_1 _27385_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1753),
    .D(_01007_),
    .Q_N(_12395_),
    .Q(\scanline[88][4] ));
 sg13g2_dfrbp_1 _27386_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1752),
    .D(_01008_),
    .Q_N(_12394_),
    .Q(\scanline[88][5] ));
 sg13g2_dfrbp_1 _27387_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1751),
    .D(_01009_),
    .Q_N(_12393_),
    .Q(\scanline[88][6] ));
 sg13g2_dfrbp_1 _27388_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1750),
    .D(_01010_),
    .Q_N(_12392_),
    .Q(\scanline[132][0] ));
 sg13g2_dfrbp_1 _27389_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1749),
    .D(_01011_),
    .Q_N(_12391_),
    .Q(\scanline[132][1] ));
 sg13g2_dfrbp_1 _27390_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1748),
    .D(_01012_),
    .Q_N(_12390_),
    .Q(\scanline[132][2] ));
 sg13g2_dfrbp_1 _27391_ (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1747),
    .D(_01013_),
    .Q_N(_12389_),
    .Q(\scanline[132][3] ));
 sg13g2_dfrbp_1 _27392_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1746),
    .D(_01014_),
    .Q_N(_12388_),
    .Q(\scanline[132][4] ));
 sg13g2_dfrbp_1 _27393_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1745),
    .D(_01015_),
    .Q_N(_12387_),
    .Q(\scanline[132][5] ));
 sg13g2_dfrbp_1 _27394_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1744),
    .D(_01016_),
    .Q_N(_12386_),
    .Q(\scanline[132][6] ));
 sg13g2_dfrbp_1 _27395_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1743),
    .D(_01017_),
    .Q_N(_12385_),
    .Q(\scanline[87][0] ));
 sg13g2_dfrbp_1 _27396_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1742),
    .D(_01018_),
    .Q_N(_12384_),
    .Q(\scanline[87][1] ));
 sg13g2_dfrbp_1 _27397_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1741),
    .D(_01019_),
    .Q_N(_12383_),
    .Q(\scanline[87][2] ));
 sg13g2_dfrbp_1 _27398_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1740),
    .D(_01020_),
    .Q_N(_12382_),
    .Q(\scanline[87][3] ));
 sg13g2_dfrbp_1 _27399_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1739),
    .D(_01021_),
    .Q_N(_12381_),
    .Q(\scanline[87][4] ));
 sg13g2_dfrbp_1 _27400_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1738),
    .D(_01022_),
    .Q_N(_12380_),
    .Q(\scanline[87][5] ));
 sg13g2_dfrbp_1 _27401_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1737),
    .D(_01023_),
    .Q_N(_12379_),
    .Q(\scanline[87][6] ));
 sg13g2_dfrbp_1 _27402_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1736),
    .D(_01024_),
    .Q_N(_12378_),
    .Q(\scanline[86][0] ));
 sg13g2_dfrbp_1 _27403_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1735),
    .D(_01025_),
    .Q_N(_12377_),
    .Q(\scanline[86][1] ));
 sg13g2_dfrbp_1 _27404_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1734),
    .D(_01026_),
    .Q_N(_12376_),
    .Q(\scanline[86][2] ));
 sg13g2_dfrbp_1 _27405_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1733),
    .D(_01027_),
    .Q_N(_12375_),
    .Q(\scanline[86][3] ));
 sg13g2_dfrbp_1 _27406_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1732),
    .D(_01028_),
    .Q_N(_12374_),
    .Q(\scanline[86][4] ));
 sg13g2_dfrbp_1 _27407_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1731),
    .D(_01029_),
    .Q_N(_12373_),
    .Q(\scanline[86][5] ));
 sg13g2_dfrbp_1 _27408_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1730),
    .D(_01030_),
    .Q_N(_12372_),
    .Q(\scanline[86][6] ));
 sg13g2_dfrbp_1 _27409_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1729),
    .D(_01031_),
    .Q_N(_12371_),
    .Q(\scanline[131][0] ));
 sg13g2_dfrbp_1 _27410_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1728),
    .D(_01032_),
    .Q_N(_12370_),
    .Q(\scanline[131][1] ));
 sg13g2_dfrbp_1 _27411_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1727),
    .D(_01033_),
    .Q_N(_12369_),
    .Q(\scanline[131][2] ));
 sg13g2_dfrbp_1 _27412_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1726),
    .D(_01034_),
    .Q_N(_12368_),
    .Q(\scanline[131][3] ));
 sg13g2_dfrbp_1 _27413_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1725),
    .D(_01035_),
    .Q_N(_12367_),
    .Q(\scanline[131][4] ));
 sg13g2_dfrbp_1 _27414_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1724),
    .D(_01036_),
    .Q_N(_12366_),
    .Q(\scanline[131][5] ));
 sg13g2_dfrbp_1 _27415_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1723),
    .D(_01037_),
    .Q_N(_12365_),
    .Q(\scanline[131][6] ));
 sg13g2_dfrbp_1 _27416_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1722),
    .D(_01038_),
    .Q_N(_12364_),
    .Q(\scanline[85][0] ));
 sg13g2_dfrbp_1 _27417_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1721),
    .D(_01039_),
    .Q_N(_12363_),
    .Q(\scanline[85][1] ));
 sg13g2_dfrbp_1 _27418_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1720),
    .D(_01040_),
    .Q_N(_12362_),
    .Q(\scanline[85][2] ));
 sg13g2_dfrbp_1 _27419_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1719),
    .D(_01041_),
    .Q_N(_12361_),
    .Q(\scanline[85][3] ));
 sg13g2_dfrbp_1 _27420_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1718),
    .D(_01042_),
    .Q_N(_12360_),
    .Q(\scanline[85][4] ));
 sg13g2_dfrbp_1 _27421_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1716),
    .D(_01043_),
    .Q_N(_12359_),
    .Q(\scanline[85][5] ));
 sg13g2_dfrbp_1 _27422_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1715),
    .D(_01044_),
    .Q_N(_12358_),
    .Q(\scanline[85][6] ));
 sg13g2_dfrbp_1 _27423_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1714),
    .D(_01045_),
    .Q_N(_12357_),
    .Q(\scanline[84][0] ));
 sg13g2_dfrbp_1 _27424_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1713),
    .D(_01046_),
    .Q_N(_12356_),
    .Q(\scanline[84][1] ));
 sg13g2_dfrbp_1 _27425_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1712),
    .D(_01047_),
    .Q_N(_12355_),
    .Q(\scanline[84][2] ));
 sg13g2_dfrbp_1 _27426_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1711),
    .D(_01048_),
    .Q_N(_12354_),
    .Q(\scanline[84][3] ));
 sg13g2_dfrbp_1 _27427_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1710),
    .D(_01049_),
    .Q_N(_12353_),
    .Q(\scanline[84][4] ));
 sg13g2_dfrbp_1 _27428_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1709),
    .D(_01050_),
    .Q_N(_12352_),
    .Q(\scanline[84][5] ));
 sg13g2_dfrbp_1 _27429_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1708),
    .D(_01051_),
    .Q_N(_12351_),
    .Q(\scanline[84][6] ));
 sg13g2_dfrbp_1 _27430_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1707),
    .D(_01052_),
    .Q_N(_12350_),
    .Q(\scanline[130][0] ));
 sg13g2_dfrbp_1 _27431_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1706),
    .D(_01053_),
    .Q_N(_12349_),
    .Q(\scanline[130][1] ));
 sg13g2_dfrbp_1 _27432_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1705),
    .D(_01054_),
    .Q_N(_12348_),
    .Q(\scanline[130][2] ));
 sg13g2_dfrbp_1 _27433_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1704),
    .D(_01055_),
    .Q_N(_12347_),
    .Q(\scanline[130][3] ));
 sg13g2_dfrbp_1 _27434_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1703),
    .D(_01056_),
    .Q_N(_12346_),
    .Q(\scanline[130][4] ));
 sg13g2_dfrbp_1 _27435_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1702),
    .D(_01057_),
    .Q_N(_12345_),
    .Q(\scanline[130][5] ));
 sg13g2_dfrbp_1 _27436_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1701),
    .D(_01058_),
    .Q_N(_12344_),
    .Q(\scanline[130][6] ));
 sg13g2_dfrbp_1 _27437_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1700),
    .D(_01059_),
    .Q_N(_12343_),
    .Q(\scanline[83][0] ));
 sg13g2_dfrbp_1 _27438_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1699),
    .D(_01060_),
    .Q_N(_12342_),
    .Q(\scanline[83][1] ));
 sg13g2_dfrbp_1 _27439_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1698),
    .D(_01061_),
    .Q_N(_12341_),
    .Q(\scanline[83][2] ));
 sg13g2_dfrbp_1 _27440_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1697),
    .D(_01062_),
    .Q_N(_12340_),
    .Q(\scanline[83][3] ));
 sg13g2_dfrbp_1 _27441_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1696),
    .D(_01063_),
    .Q_N(_12339_),
    .Q(\scanline[83][4] ));
 sg13g2_dfrbp_1 _27442_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1695),
    .D(_01064_),
    .Q_N(_12338_),
    .Q(\scanline[83][5] ));
 sg13g2_dfrbp_1 _27443_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1694),
    .D(_01065_),
    .Q_N(_12337_),
    .Q(\scanline[83][6] ));
 sg13g2_dfrbp_1 _27444_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1693),
    .D(_01066_),
    .Q_N(_12336_),
    .Q(\scanline[82][0] ));
 sg13g2_dfrbp_1 _27445_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1692),
    .D(_01067_),
    .Q_N(_12335_),
    .Q(\scanline[82][1] ));
 sg13g2_dfrbp_1 _27446_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1691),
    .D(_01068_),
    .Q_N(_12334_),
    .Q(\scanline[82][2] ));
 sg13g2_dfrbp_1 _27447_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1690),
    .D(_01069_),
    .Q_N(_12333_),
    .Q(\scanline[82][3] ));
 sg13g2_dfrbp_1 _27448_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1689),
    .D(_01070_),
    .Q_N(_12332_),
    .Q(\scanline[82][4] ));
 sg13g2_dfrbp_1 _27449_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1688),
    .D(_01071_),
    .Q_N(_12331_),
    .Q(\scanline[82][5] ));
 sg13g2_dfrbp_1 _27450_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1687),
    .D(_01072_),
    .Q_N(_12330_),
    .Q(\scanline[82][6] ));
 sg13g2_dfrbp_1 _27451_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1686),
    .D(_01073_),
    .Q_N(_12329_),
    .Q(\scanline[12][0] ));
 sg13g2_dfrbp_1 _27452_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1685),
    .D(_01074_),
    .Q_N(_12328_),
    .Q(\scanline[12][1] ));
 sg13g2_dfrbp_1 _27453_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1684),
    .D(_01075_),
    .Q_N(_12327_),
    .Q(\scanline[12][2] ));
 sg13g2_dfrbp_1 _27454_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1683),
    .D(_01076_),
    .Q_N(_12326_),
    .Q(\scanline[12][3] ));
 sg13g2_dfrbp_1 _27455_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1682),
    .D(_01077_),
    .Q_N(_12325_),
    .Q(\scanline[12][4] ));
 sg13g2_dfrbp_1 _27456_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1681),
    .D(_01078_),
    .Q_N(_12324_),
    .Q(\scanline[12][5] ));
 sg13g2_dfrbp_1 _27457_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1680),
    .D(_01079_),
    .Q_N(_12323_),
    .Q(\scanline[12][6] ));
 sg13g2_dfrbp_1 _27458_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1679),
    .D(_01080_),
    .Q_N(_12322_),
    .Q(\scanline[7][0] ));
 sg13g2_dfrbp_1 _27459_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1678),
    .D(_01081_),
    .Q_N(_12321_),
    .Q(\scanline[7][1] ));
 sg13g2_dfrbp_1 _27460_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1677),
    .D(_01082_),
    .Q_N(_12320_),
    .Q(\scanline[7][2] ));
 sg13g2_dfrbp_1 _27461_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1676),
    .D(_01083_),
    .Q_N(_12319_),
    .Q(\scanline[7][3] ));
 sg13g2_dfrbp_1 _27462_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1675),
    .D(_01084_),
    .Q_N(_12318_),
    .Q(\scanline[7][4] ));
 sg13g2_dfrbp_1 _27463_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1674),
    .D(_01085_),
    .Q_N(_12317_),
    .Q(\scanline[7][5] ));
 sg13g2_dfrbp_1 _27464_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1673),
    .D(_01086_),
    .Q_N(_12316_),
    .Q(\scanline[7][6] ));
 sg13g2_dfrbp_1 _27465_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1672),
    .D(_01087_),
    .Q_N(_12315_),
    .Q(\scanline[78][0] ));
 sg13g2_dfrbp_1 _27466_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1671),
    .D(_01088_),
    .Q_N(_12314_),
    .Q(\scanline[78][1] ));
 sg13g2_dfrbp_1 _27467_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1670),
    .D(_01089_),
    .Q_N(_12313_),
    .Q(\scanline[78][2] ));
 sg13g2_dfrbp_1 _27468_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1669),
    .D(_01090_),
    .Q_N(_12312_),
    .Q(\scanline[78][3] ));
 sg13g2_dfrbp_1 _27469_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1668),
    .D(_01091_),
    .Q_N(_12311_),
    .Q(\scanline[78][4] ));
 sg13g2_dfrbp_1 _27470_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1667),
    .D(_01092_),
    .Q_N(_12310_),
    .Q(\scanline[78][5] ));
 sg13g2_dfrbp_1 _27471_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1666),
    .D(_01093_),
    .Q_N(_12309_),
    .Q(\scanline[78][6] ));
 sg13g2_dfrbp_1 _27472_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1665),
    .D(_01094_),
    .Q_N(_12308_),
    .Q(\scanline[75][0] ));
 sg13g2_dfrbp_1 _27473_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1664),
    .D(_01095_),
    .Q_N(_12307_),
    .Q(\scanline[75][1] ));
 sg13g2_dfrbp_1 _27474_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1663),
    .D(_01096_),
    .Q_N(_12306_),
    .Q(\scanline[75][2] ));
 sg13g2_dfrbp_1 _27475_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1662),
    .D(_01097_),
    .Q_N(_12305_),
    .Q(\scanline[75][3] ));
 sg13g2_dfrbp_1 _27476_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1661),
    .D(_01098_),
    .Q_N(_12304_),
    .Q(\scanline[75][4] ));
 sg13g2_dfrbp_1 _27477_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1660),
    .D(_01099_),
    .Q_N(_12303_),
    .Q(\scanline[75][5] ));
 sg13g2_dfrbp_1 _27478_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1659),
    .D(_01100_),
    .Q_N(_12302_),
    .Q(\scanline[75][6] ));
 sg13g2_dfrbp_1 _27479_ (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1658),
    .D(_01101_),
    .Q_N(_12301_),
    .Q(\scanline[77][0] ));
 sg13g2_dfrbp_1 _27480_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1657),
    .D(_01102_),
    .Q_N(_12300_),
    .Q(\scanline[77][1] ));
 sg13g2_dfrbp_1 _27481_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1656),
    .D(_01103_),
    .Q_N(_12299_),
    .Q(\scanline[77][2] ));
 sg13g2_dfrbp_1 _27482_ (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1655),
    .D(_01104_),
    .Q_N(_12298_),
    .Q(\scanline[77][3] ));
 sg13g2_dfrbp_1 _27483_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1654),
    .D(_01105_),
    .Q_N(_12297_),
    .Q(\scanline[77][4] ));
 sg13g2_dfrbp_1 _27484_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1653),
    .D(_01106_),
    .Q_N(_12296_),
    .Q(\scanline[77][5] ));
 sg13g2_dfrbp_1 _27485_ (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1652),
    .D(_01107_),
    .Q_N(_12295_),
    .Q(\scanline[77][6] ));
 sg13g2_dfrbp_1 _27486_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1651),
    .D(_01108_),
    .Q_N(_12294_),
    .Q(\scanline[70][0] ));
 sg13g2_dfrbp_1 _27487_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1650),
    .D(_01109_),
    .Q_N(_12293_),
    .Q(\scanline[70][1] ));
 sg13g2_dfrbp_1 _27488_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1649),
    .D(_01110_),
    .Q_N(_12292_),
    .Q(\scanline[70][2] ));
 sg13g2_dfrbp_1 _27489_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1648),
    .D(_01111_),
    .Q_N(_12291_),
    .Q(\scanline[70][3] ));
 sg13g2_dfrbp_1 _27490_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1647),
    .D(_01112_),
    .Q_N(_12290_),
    .Q(\scanline[70][4] ));
 sg13g2_dfrbp_1 _27491_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1646),
    .D(_01113_),
    .Q_N(_12289_),
    .Q(\scanline[70][5] ));
 sg13g2_dfrbp_1 _27492_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1645),
    .D(_01114_),
    .Q_N(_12288_),
    .Q(\scanline[70][6] ));
 sg13g2_dfrbp_1 _27493_ (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1644),
    .D(_01115_),
    .Q_N(_12287_),
    .Q(\scanline[73][0] ));
 sg13g2_dfrbp_1 _27494_ (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1643),
    .D(_01116_),
    .Q_N(_12286_),
    .Q(\scanline[73][1] ));
 sg13g2_dfrbp_1 _27495_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1642),
    .D(_01117_),
    .Q_N(_12285_),
    .Q(\scanline[73][2] ));
 sg13g2_dfrbp_1 _27496_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1641),
    .D(_01118_),
    .Q_N(_12284_),
    .Q(\scanline[73][3] ));
 sg13g2_dfrbp_1 _27497_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1640),
    .D(_01119_),
    .Q_N(_12283_),
    .Q(\scanline[73][4] ));
 sg13g2_dfrbp_1 _27498_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1639),
    .D(_01120_),
    .Q_N(_12282_),
    .Q(\scanline[73][5] ));
 sg13g2_dfrbp_1 _27499_ (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1638),
    .D(_01121_),
    .Q_N(_12281_),
    .Q(\scanline[73][6] ));
 sg13g2_dfrbp_1 _27500_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1637),
    .D(_01122_),
    .Q_N(_12280_),
    .Q(spi_restart));
 sg13g2_dfrbp_1 _27501_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1636),
    .D(_01123_),
    .Q_N(_13232_),
    .Q(\flash_rom.stall_read ));
 sg13g2_dfrbp_1 _27502_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1717),
    .D(net2892),
    .Q_N(_13233_),
    .Q(spi_data_ready_last));
 sg13g2_dfrbp_1 _27503_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1633),
    .D(_00000_),
    .Q_N(_12279_),
    .Q(rom_data_pending));
 sg13g2_dfrbp_1 _27504_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1631),
    .D(_01124_),
    .Q_N(_00171_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 _27505_ (.CLK(clknet_6_55__leaf_clk),
    .RESET_B(net1630),
    .D(_01125_),
    .Q_N(_12278_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 _27506_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1629),
    .D(_01126_),
    .Q_N(_12277_),
    .Q(\rom_last_read_addr[0] ));
 sg13g2_dfrbp_1 _27507_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1628),
    .D(_01127_),
    .Q_N(_12276_),
    .Q(\rom_last_read_addr[1] ));
 sg13g2_dfrbp_1 _27508_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1627),
    .D(net6934),
    .Q_N(_12275_),
    .Q(\rom_last_read_addr[2] ));
 sg13g2_dfrbp_1 _27509_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1626),
    .D(net6619),
    .Q_N(_12274_),
    .Q(\rom_last_read_addr[3] ));
 sg13g2_dfrbp_1 _27510_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1625),
    .D(net3975),
    .Q_N(_12273_),
    .Q(\rom_last_read_addr[4] ));
 sg13g2_dfrbp_1 _27511_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1624),
    .D(net3978),
    .Q_N(_12272_),
    .Q(\rom_last_read_addr[5] ));
 sg13g2_dfrbp_1 _27512_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1623),
    .D(net6724),
    .Q_N(_12271_),
    .Q(\rom_last_read_addr[6] ));
 sg13g2_dfrbp_1 _27513_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1622),
    .D(net6853),
    .Q_N(_12270_),
    .Q(\rom_last_read_addr[7] ));
 sg13g2_dfrbp_1 _27514_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1621),
    .D(net6985),
    .Q_N(_12269_),
    .Q(\rom_last_read_addr[8] ));
 sg13g2_dfrbp_1 _27515_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1620),
    .D(net7054),
    .Q_N(_12268_),
    .Q(\rom_last_read_addr[9] ));
 sg13g2_dfrbp_1 _27516_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1619),
    .D(net6954),
    .Q_N(_12267_),
    .Q(\rom_last_read_addr[10] ));
 sg13g2_dfrbp_1 _27517_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1618),
    .D(net6768),
    .Q_N(_12266_),
    .Q(\rom_last_read_addr[11] ));
 sg13g2_dfrbp_1 _27518_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1617),
    .D(net7019),
    .Q_N(_00105_),
    .Q(\rom_next_addr_in_queue[0] ));
 sg13g2_dfrbp_1 _27519_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1616),
    .D(_01139_),
    .Q_N(_12265_),
    .Q(\rom_next_addr_in_queue[1] ));
 sg13g2_dfrbp_1 _27520_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1615),
    .D(net7243),
    .Q_N(_12264_),
    .Q(\rom_next_addr_in_queue[2] ));
 sg13g2_dfrbp_1 _27521_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1614),
    .D(_01141_),
    .Q_N(_12263_),
    .Q(\rom_next_addr_in_queue[3] ));
 sg13g2_dfrbp_1 _27522_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1613),
    .D(_01142_),
    .Q_N(_12262_),
    .Q(\rom_next_addr_in_queue[4] ));
 sg13g2_dfrbp_1 _27523_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1612),
    .D(_01143_),
    .Q_N(_12261_),
    .Q(\rom_next_addr_in_queue[5] ));
 sg13g2_dfrbp_1 _27524_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1611),
    .D(_01144_),
    .Q_N(_12260_),
    .Q(\rom_next_addr_in_queue[6] ));
 sg13g2_dfrbp_1 _27525_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1610),
    .D(_01145_),
    .Q_N(_12259_),
    .Q(\rom_next_addr_in_queue[7] ));
 sg13g2_dfrbp_1 _27526_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1609),
    .D(_01146_),
    .Q_N(_12258_),
    .Q(\rom_next_addr_in_queue[8] ));
 sg13g2_dfrbp_1 _27527_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1608),
    .D(_01147_),
    .Q_N(_12257_),
    .Q(\rom_next_addr_in_queue[9] ));
 sg13g2_dfrbp_1 _27528_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1607),
    .D(_01148_),
    .Q_N(_12256_),
    .Q(\rom_next_addr_in_queue[10] ));
 sg13g2_dfrbp_1 _27529_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1606),
    .D(_01149_),
    .Q_N(_12255_),
    .Q(\rom_next_addr_in_queue[11] ));
 sg13g2_dfrbp_1 _27530_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1605),
    .D(net7013),
    .Q_N(_12254_),
    .Q(\audio_pwm_accumulator[0] ));
 sg13g2_dfrbp_1 _27531_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1604),
    .D(_01151_),
    .Q_N(_12253_),
    .Q(\audio_pwm_accumulator[1] ));
 sg13g2_dfrbp_1 _27532_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1603),
    .D(_01152_),
    .Q_N(_12252_),
    .Q(\audio_pwm_accumulator[2] ));
 sg13g2_dfrbp_1 _27533_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1602),
    .D(_01153_),
    .Q_N(_12251_),
    .Q(\audio_pwm_accumulator[3] ));
 sg13g2_dfrbp_1 _27534_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1601),
    .D(_01154_),
    .Q_N(_12250_),
    .Q(\audio_pwm_accumulator[4] ));
 sg13g2_dfrbp_1 _27535_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1600),
    .D(_01155_),
    .Q_N(_12249_),
    .Q(audio_pwm));
 sg13g2_dfrbp_1 _27536_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1599),
    .D(_01156_),
    .Q_N(_12248_),
    .Q(\r_pwm_odd[1] ));
 sg13g2_dfrbp_1 _27537_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1598),
    .D(_01157_),
    .Q_N(_12247_),
    .Q(\r_pwm_odd[2] ));
 sg13g2_dfrbp_1 _27538_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1597),
    .D(_01158_),
    .Q_N(_00063_),
    .Q(\r_pwm_odd[3] ));
 sg13g2_dfrbp_1 _27539_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1596),
    .D(_01159_),
    .Q_N(_12246_),
    .Q(\r_pwm_odd[4] ));
 sg13g2_dfrbp_1 _27540_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1595),
    .D(_01160_),
    .Q_N(_12245_),
    .Q(\r_pwm_odd[5] ));
 sg13g2_dfrbp_1 _27541_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1594),
    .D(_01161_),
    .Q_N(_12244_),
    .Q(\r_pwm_odd[6] ));
 sg13g2_dfrbp_1 _27542_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1593),
    .D(_01162_),
    .Q_N(_12243_),
    .Q(\r_pwm_odd[7] ));
 sg13g2_dfrbp_1 _27543_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1592),
    .D(_01163_),
    .Q_N(_12242_),
    .Q(\r_pwm_odd[8] ));
 sg13g2_dfrbp_1 _27544_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1591),
    .D(_01164_),
    .Q_N(_12241_),
    .Q(\r_pwm_odd[9] ));
 sg13g2_dfrbp_1 _27545_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1590),
    .D(_01165_),
    .Q_N(_12240_),
    .Q(\g_pwm_odd[1] ));
 sg13g2_dfrbp_1 _27546_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1589),
    .D(_01166_),
    .Q_N(_12239_),
    .Q(\g_pwm_odd[2] ));
 sg13g2_dfrbp_1 _27547_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1588),
    .D(_01167_),
    .Q_N(_00062_),
    .Q(\g_pwm_odd[3] ));
 sg13g2_dfrbp_1 _27548_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1587),
    .D(_01168_),
    .Q_N(_12238_),
    .Q(\g_pwm_odd[4] ));
 sg13g2_dfrbp_1 _27549_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1586),
    .D(_01169_),
    .Q_N(_12237_),
    .Q(\g_pwm_odd[5] ));
 sg13g2_dfrbp_1 _27550_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1585),
    .D(_01170_),
    .Q_N(_12236_),
    .Q(\g_pwm_odd[6] ));
 sg13g2_dfrbp_1 _27551_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1584),
    .D(_01171_),
    .Q_N(_12235_),
    .Q(\g_pwm_odd[7] ));
 sg13g2_dfrbp_1 _27552_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1583),
    .D(_01172_),
    .Q_N(_12234_),
    .Q(\g_pwm_odd[8] ));
 sg13g2_dfrbp_1 _27553_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1582),
    .D(_01173_),
    .Q_N(_12233_),
    .Q(\g_pwm_odd[9] ));
 sg13g2_dfrbp_1 _27554_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1581),
    .D(_01174_),
    .Q_N(_12232_),
    .Q(\b_pwm_odd[1] ));
 sg13g2_dfrbp_1 _27555_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1580),
    .D(_01175_),
    .Q_N(_12231_),
    .Q(\b_pwm_odd[2] ));
 sg13g2_dfrbp_1 _27556_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1579),
    .D(_01176_),
    .Q_N(_12230_),
    .Q(\b_pwm_odd[3] ));
 sg13g2_dfrbp_1 _27557_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1578),
    .D(_01177_),
    .Q_N(_12229_),
    .Q(\b_pwm_odd[4] ));
 sg13g2_dfrbp_1 _27558_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1577),
    .D(_01178_),
    .Q_N(_12228_),
    .Q(\b_pwm_odd[5] ));
 sg13g2_dfrbp_1 _27559_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1576),
    .D(_01179_),
    .Q_N(_12227_),
    .Q(\b_pwm_odd[6] ));
 sg13g2_dfrbp_1 _27560_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1575),
    .D(_01180_),
    .Q_N(_12226_),
    .Q(\b_pwm_odd[7] ));
 sg13g2_dfrbp_1 _27561_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1574),
    .D(_01181_),
    .Q_N(_12225_),
    .Q(\b_pwm_odd[8] ));
 sg13g2_dfrbp_1 _27562_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1573),
    .D(_01182_),
    .Q_N(_12224_),
    .Q(\b_pwm_odd[9] ));
 sg13g2_dfrbp_1 _27563_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1572),
    .D(net3735),
    .Q_N(_12223_),
    .Q(\r_pwm_even[1] ));
 sg13g2_dfrbp_1 _27564_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1571),
    .D(_01184_),
    .Q_N(_12222_),
    .Q(\r_pwm_even[2] ));
 sg13g2_dfrbp_1 _27565_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1570),
    .D(_01185_),
    .Q_N(_12221_),
    .Q(\r_pwm_even[3] ));
 sg13g2_dfrbp_1 _27566_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1569),
    .D(_01186_),
    .Q_N(_12220_),
    .Q(\r_pwm_even[4] ));
 sg13g2_dfrbp_1 _27567_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1568),
    .D(_01187_),
    .Q_N(_12219_),
    .Q(\r_pwm_even[5] ));
 sg13g2_dfrbp_1 _27568_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1567),
    .D(_01188_),
    .Q_N(_12218_),
    .Q(\r_pwm_even[6] ));
 sg13g2_dfrbp_1 _27569_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1566),
    .D(_01189_),
    .Q_N(_12217_),
    .Q(\r_pwm_even[7] ));
 sg13g2_dfrbp_1 _27570_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1565),
    .D(_01190_),
    .Q_N(_12216_),
    .Q(\r_pwm_even[8] ));
 sg13g2_dfrbp_1 _27571_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1564),
    .D(_01191_),
    .Q_N(_12215_),
    .Q(\r_pwm_even[9] ));
 sg13g2_dfrbp_1 _27572_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1563),
    .D(net3763),
    .Q_N(_12214_),
    .Q(\g_pwm_even[1] ));
 sg13g2_dfrbp_1 _27573_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1562),
    .D(_01193_),
    .Q_N(_12213_),
    .Q(\g_pwm_even[2] ));
 sg13g2_dfrbp_1 _27574_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1561),
    .D(_01194_),
    .Q_N(_12212_),
    .Q(\g_pwm_even[3] ));
 sg13g2_dfrbp_1 _27575_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1560),
    .D(_01195_),
    .Q_N(_12211_),
    .Q(\g_pwm_even[4] ));
 sg13g2_dfrbp_1 _27576_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1559),
    .D(_01196_),
    .Q_N(_12210_),
    .Q(\g_pwm_even[5] ));
 sg13g2_dfrbp_1 _27577_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1558),
    .D(_01197_),
    .Q_N(_12209_),
    .Q(\g_pwm_even[6] ));
 sg13g2_dfrbp_1 _27578_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1557),
    .D(_01198_),
    .Q_N(_12208_),
    .Q(\g_pwm_even[7] ));
 sg13g2_dfrbp_1 _27579_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1556),
    .D(_01199_),
    .Q_N(_12207_),
    .Q(\g_pwm_even[8] ));
 sg13g2_dfrbp_1 _27580_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1555),
    .D(_01200_),
    .Q_N(_12206_),
    .Q(\g_pwm_even[9] ));
 sg13g2_dfrbp_1 _27581_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1554),
    .D(net2896),
    .Q_N(_00169_),
    .Q(\frame_counter[0] ));
 sg13g2_dfrbp_1 _27582_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1552),
    .D(net3529),
    .Q_N(_12205_),
    .Q(\frame_counter[1] ));
 sg13g2_dfrbp_1 _27583_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1783),
    .D(net6299),
    .Q_N(_13234_),
    .Q(\frame_counter[2] ));
 sg13g2_dfrbp_1 _27584_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1550),
    .D(net6931),
    .Q_N(_12204_),
    .Q(tia_vsync_last));
 sg13g2_dfrbp_1 _27585_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1548),
    .D(_01204_),
    .Q_N(_12203_),
    .Q(\scanline[56][0] ));
 sg13g2_dfrbp_1 _27586_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1547),
    .D(_01205_),
    .Q_N(_12202_),
    .Q(\scanline[56][1] ));
 sg13g2_dfrbp_1 _27587_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1546),
    .D(_01206_),
    .Q_N(_12201_),
    .Q(\scanline[56][2] ));
 sg13g2_dfrbp_1 _27588_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1545),
    .D(_01207_),
    .Q_N(_12200_),
    .Q(\scanline[56][3] ));
 sg13g2_dfrbp_1 _27589_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1544),
    .D(_01208_),
    .Q_N(_12199_),
    .Q(\scanline[56][4] ));
 sg13g2_dfrbp_1 _27590_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1543),
    .D(_01209_),
    .Q_N(_12198_),
    .Q(\scanline[56][5] ));
 sg13g2_dfrbp_1 _27591_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1542),
    .D(_01210_),
    .Q_N(_12197_),
    .Q(\scanline[56][6] ));
 sg13g2_dfrbp_1 _27592_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1541),
    .D(_01211_),
    .Q_N(_12196_),
    .Q(\atari2600.input_joystick_0[0] ));
 sg13g2_dfrbp_1 _27593_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1539),
    .D(_01212_),
    .Q_N(_12195_),
    .Q(\atari2600.input_joystick_0[1] ));
 sg13g2_dfrbp_1 _27594_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1537),
    .D(net2996),
    .Q_N(_12194_),
    .Q(\atari2600.input_joystick_0[2] ));
 sg13g2_dfrbp_1 _27595_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1535),
    .D(_01214_),
    .Q_N(_12193_),
    .Q(\atari2600.input_joystick_0[3] ));
 sg13g2_dfrbp_1 _27596_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1533),
    .D(_01215_),
    .Q_N(_12192_),
    .Q(\atari2600.input_joystick_0[4] ));
 sg13g2_dfrbp_1 _27597_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1531),
    .D(_01216_),
    .Q_N(_12191_),
    .Q(\atari2600.input_joystick_0[5] ));
 sg13g2_dfrbp_1 _27598_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1529),
    .D(_01217_),
    .Q_N(_12190_),
    .Q(\atari2600.input_joystick_0[6] ));
 sg13g2_dfrbp_1 _27599_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1527),
    .D(_01218_),
    .Q_N(_12189_),
    .Q(\joypmod[2] ));
 sg13g2_dfrbp_1 _27600_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1525),
    .D(_01219_),
    .Q_N(_12188_),
    .Q(\atari2600.input_switches[0] ));
 sg13g2_dfrbp_1 _27601_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1523),
    .D(_01220_),
    .Q_N(_12187_),
    .Q(\atari2600.input_switches[1] ));
 sg13g2_dfrbp_1 _27602_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1521),
    .D(_01221_),
    .Q_N(_12186_),
    .Q(\atari2600.input_switches[2] ));
 sg13g2_dfrbp_1 _27603_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1519),
    .D(_01222_),
    .Q_N(_12185_),
    .Q(\atari2600.input_switches[3] ));
 sg13g2_dfrbp_1 _27604_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1517),
    .D(_01223_),
    .Q_N(_12184_),
    .Q(\b_pwm_even[1] ));
 sg13g2_dfrbp_1 _27605_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1516),
    .D(_01224_),
    .Q_N(_12183_),
    .Q(\b_pwm_even[2] ));
 sg13g2_dfrbp_1 _27606_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1515),
    .D(_01225_),
    .Q_N(_12182_),
    .Q(\b_pwm_even[3] ));
 sg13g2_dfrbp_1 _27607_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1514),
    .D(_01226_),
    .Q_N(_12181_),
    .Q(\b_pwm_even[4] ));
 sg13g2_dfrbp_1 _27608_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1513),
    .D(_01227_),
    .Q_N(_12180_),
    .Q(\b_pwm_even[5] ));
 sg13g2_dfrbp_1 _27609_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1512),
    .D(_01228_),
    .Q_N(_12179_),
    .Q(\b_pwm_even[6] ));
 sg13g2_dfrbp_1 _27610_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1511),
    .D(_01229_),
    .Q_N(_12178_),
    .Q(\b_pwm_even[7] ));
 sg13g2_dfrbp_1 _27611_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1510),
    .D(_01230_),
    .Q_N(_12177_),
    .Q(\b_pwm_even[8] ));
 sg13g2_dfrbp_1 _27612_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1509),
    .D(_01231_),
    .Q_N(_12176_),
    .Q(\b_pwm_even[9] ));
 sg13g2_dfrbp_1 _27613_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1508),
    .D(_01232_),
    .Q_N(_12175_),
    .Q(\scanline[128][0] ));
 sg13g2_dfrbp_1 _27614_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1507),
    .D(_01233_),
    .Q_N(_12174_),
    .Q(\scanline[128][1] ));
 sg13g2_dfrbp_1 _27615_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1506),
    .D(_01234_),
    .Q_N(_12173_),
    .Q(\scanline[128][2] ));
 sg13g2_dfrbp_1 _27616_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1505),
    .D(_01235_),
    .Q_N(_12172_),
    .Q(\scanline[128][3] ));
 sg13g2_dfrbp_1 _27617_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1504),
    .D(_01236_),
    .Q_N(_12171_),
    .Q(\scanline[128][4] ));
 sg13g2_dfrbp_1 _27618_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1503),
    .D(_01237_),
    .Q_N(_12170_),
    .Q(\scanline[128][5] ));
 sg13g2_dfrbp_1 _27619_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1502),
    .D(_01238_),
    .Q_N(_12169_),
    .Q(\scanline[128][6] ));
 sg13g2_dfrbp_1 _27620_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1501),
    .D(_01239_),
    .Q_N(_12168_),
    .Q(\scanline[127][0] ));
 sg13g2_dfrbp_1 _27621_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1500),
    .D(_01240_),
    .Q_N(_12167_),
    .Q(\scanline[127][1] ));
 sg13g2_dfrbp_1 _27622_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1499),
    .D(_01241_),
    .Q_N(_12166_),
    .Q(\scanline[127][2] ));
 sg13g2_dfrbp_1 _27623_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1498),
    .D(_01242_),
    .Q_N(_12165_),
    .Q(\scanline[127][3] ));
 sg13g2_dfrbp_1 _27624_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1497),
    .D(_01243_),
    .Q_N(_12164_),
    .Q(\scanline[127][4] ));
 sg13g2_dfrbp_1 _27625_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1496),
    .D(_01244_),
    .Q_N(_12163_),
    .Q(\scanline[127][5] ));
 sg13g2_dfrbp_1 _27626_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1495),
    .D(_01245_),
    .Q_N(_12162_),
    .Q(\scanline[127][6] ));
 sg13g2_dfrbp_1 _27627_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1494),
    .D(_01246_),
    .Q_N(_12161_),
    .Q(\scanline[80][0] ));
 sg13g2_dfrbp_1 _27628_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1493),
    .D(_01247_),
    .Q_N(_12160_),
    .Q(\scanline[80][1] ));
 sg13g2_dfrbp_1 _27629_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1492),
    .D(_01248_),
    .Q_N(_12159_),
    .Q(\scanline[80][2] ));
 sg13g2_dfrbp_1 _27630_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1491),
    .D(_01249_),
    .Q_N(_12158_),
    .Q(\scanline[80][3] ));
 sg13g2_dfrbp_1 _27631_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1490),
    .D(_01250_),
    .Q_N(_12157_),
    .Q(\scanline[80][4] ));
 sg13g2_dfrbp_1 _27632_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1489),
    .D(_01251_),
    .Q_N(_12156_),
    .Q(\scanline[80][5] ));
 sg13g2_dfrbp_1 _27633_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1488),
    .D(_01252_),
    .Q_N(_12155_),
    .Q(\scanline[80][6] ));
 sg13g2_dfrbp_1 _27634_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1487),
    .D(_01253_),
    .Q_N(_12154_),
    .Q(\atari2600.ram[75][0] ));
 sg13g2_dfrbp_1 _27635_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1486),
    .D(_01254_),
    .Q_N(_12153_),
    .Q(\atari2600.ram[75][1] ));
 sg13g2_dfrbp_1 _27636_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1485),
    .D(_01255_),
    .Q_N(_12152_),
    .Q(\atari2600.ram[75][2] ));
 sg13g2_dfrbp_1 _27637_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1484),
    .D(_01256_),
    .Q_N(_12151_),
    .Q(\atari2600.ram[75][3] ));
 sg13g2_dfrbp_1 _27638_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1483),
    .D(_01257_),
    .Q_N(_12150_),
    .Q(\atari2600.ram[75][4] ));
 sg13g2_dfrbp_1 _27639_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1482),
    .D(_01258_),
    .Q_N(_12149_),
    .Q(\atari2600.ram[75][5] ));
 sg13g2_dfrbp_1 _27640_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1481),
    .D(_01259_),
    .Q_N(_12148_),
    .Q(\atari2600.ram[75][6] ));
 sg13g2_dfrbp_1 _27641_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1480),
    .D(_01260_),
    .Q_N(_12147_),
    .Q(\atari2600.ram[75][7] ));
 sg13g2_dfrbp_1 _27642_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1479),
    .D(_01261_),
    .Q_N(_12146_),
    .Q(\atari2600.ram[127][0] ));
 sg13g2_dfrbp_1 _27643_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1478),
    .D(_01262_),
    .Q_N(_12145_),
    .Q(\atari2600.ram[127][1] ));
 sg13g2_dfrbp_1 _27644_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1477),
    .D(_01263_),
    .Q_N(_12144_),
    .Q(\atari2600.ram[127][2] ));
 sg13g2_dfrbp_1 _27645_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1476),
    .D(_01264_),
    .Q_N(_12143_),
    .Q(\atari2600.ram[127][3] ));
 sg13g2_dfrbp_1 _27646_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1475),
    .D(_01265_),
    .Q_N(_12142_),
    .Q(\atari2600.ram[127][4] ));
 sg13g2_dfrbp_1 _27647_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1474),
    .D(_01266_),
    .Q_N(_12141_),
    .Q(\atari2600.ram[127][5] ));
 sg13g2_dfrbp_1 _27648_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1473),
    .D(_01267_),
    .Q_N(_12140_),
    .Q(\atari2600.ram[127][6] ));
 sg13g2_dfrbp_1 _27649_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1784),
    .D(_01268_),
    .Q_N(_13235_),
    .Q(\atari2600.ram[127][7] ));
 sg13g2_dfrbp_1 _27650_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net5997),
    .D(_00173_),
    .Q_N(_13236_),
    .Q(\atari2600.cpu.state[0] ));
 sg13g2_dfrbp_1 _27651_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net5997),
    .D(_00174_),
    .Q_N(_13237_),
    .Q(\atari2600.cpu.state[1] ));
 sg13g2_dfrbp_1 _27652_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net5997),
    .D(_00175_),
    .Q_N(_12139_),
    .Q(\atari2600.cpu.state[2] ));
 sg13g2_dfrbp_1 _27653_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net5997),
    .D(_00178_),
    .Q_N(\atari2600.cpu.state[3] ),
    .Q(_00172_));
 sg13g2_dfrbp_1 _27654_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net5997),
    .D(_00176_),
    .Q_N(_13238_),
    .Q(\atari2600.cpu.state[4] ));
 sg13g2_dfrbp_1 _27655_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net5997),
    .D(_00177_),
    .Q_N(_12138_),
    .Q(\atari2600.cpu.state[5] ));
 sg13g2_dfrbp_1 _27656_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1471),
    .D(_01269_),
    .Q_N(_12137_),
    .Q(\atari2600.ram[7][0] ));
 sg13g2_dfrbp_1 _27657_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1470),
    .D(_01270_),
    .Q_N(_12136_),
    .Q(\atari2600.ram[7][1] ));
 sg13g2_dfrbp_1 _27658_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1469),
    .D(_01271_),
    .Q_N(_12135_),
    .Q(\atari2600.ram[7][2] ));
 sg13g2_dfrbp_1 _27659_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1468),
    .D(_01272_),
    .Q_N(_12134_),
    .Q(\atari2600.ram[7][3] ));
 sg13g2_dfrbp_1 _27660_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1467),
    .D(_01273_),
    .Q_N(_12133_),
    .Q(\atari2600.ram[7][4] ));
 sg13g2_dfrbp_1 _27661_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1466),
    .D(_01274_),
    .Q_N(_12132_),
    .Q(\atari2600.ram[7][5] ));
 sg13g2_dfrbp_1 _27662_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1465),
    .D(_01275_),
    .Q_N(_12131_),
    .Q(\atari2600.ram[7][6] ));
 sg13g2_dfrbp_1 _27663_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1464),
    .D(_01276_),
    .Q_N(_12130_),
    .Q(\atari2600.ram[7][7] ));
 sg13g2_dfrbp_1 _27664_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1463),
    .D(_01277_),
    .Q_N(_12129_),
    .Q(\atari2600.ram[84][0] ));
 sg13g2_dfrbp_1 _27665_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1462),
    .D(_01278_),
    .Q_N(_12128_),
    .Q(\atari2600.ram[84][1] ));
 sg13g2_dfrbp_1 _27666_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1461),
    .D(_01279_),
    .Q_N(_12127_),
    .Q(\atari2600.ram[84][2] ));
 sg13g2_dfrbp_1 _27667_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1460),
    .D(_01280_),
    .Q_N(_12126_),
    .Q(\atari2600.ram[84][3] ));
 sg13g2_dfrbp_1 _27668_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1459),
    .D(_01281_),
    .Q_N(_12125_),
    .Q(\atari2600.ram[84][4] ));
 sg13g2_dfrbp_1 _27669_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1458),
    .D(_01282_),
    .Q_N(_12124_),
    .Q(\atari2600.ram[84][5] ));
 sg13g2_dfrbp_1 _27670_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1457),
    .D(_01283_),
    .Q_N(_12123_),
    .Q(\atari2600.ram[84][6] ));
 sg13g2_dfrbp_1 _27671_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1456),
    .D(_01284_),
    .Q_N(_12122_),
    .Q(\atari2600.ram[84][7] ));
 sg13g2_dfrbp_1 _27672_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1455),
    .D(_01285_),
    .Q_N(_12121_),
    .Q(\atari2600.ram[76][0] ));
 sg13g2_dfrbp_1 _27673_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1454),
    .D(_01286_),
    .Q_N(_12120_),
    .Q(\atari2600.ram[76][1] ));
 sg13g2_dfrbp_1 _27674_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1453),
    .D(_01287_),
    .Q_N(_12119_),
    .Q(\atari2600.ram[76][2] ));
 sg13g2_dfrbp_1 _27675_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1452),
    .D(_01288_),
    .Q_N(_12118_),
    .Q(\atari2600.ram[76][3] ));
 sg13g2_dfrbp_1 _27676_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1451),
    .D(_01289_),
    .Q_N(_12117_),
    .Q(\atari2600.ram[76][4] ));
 sg13g2_dfrbp_1 _27677_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1450),
    .D(_01290_),
    .Q_N(_12116_),
    .Q(\atari2600.ram[76][5] ));
 sg13g2_dfrbp_1 _27678_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1449),
    .D(_01291_),
    .Q_N(_12115_),
    .Q(\atari2600.ram[76][6] ));
 sg13g2_dfrbp_1 _27679_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1448),
    .D(_01292_),
    .Q_N(_12114_),
    .Q(\atari2600.ram[76][7] ));
 sg13g2_dfrbp_1 _27680_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1447),
    .D(_01293_),
    .Q_N(_12113_),
    .Q(\atari2600.ram[81][0] ));
 sg13g2_dfrbp_1 _27681_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1446),
    .D(_01294_),
    .Q_N(_12112_),
    .Q(\atari2600.ram[81][1] ));
 sg13g2_dfrbp_1 _27682_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1445),
    .D(_01295_),
    .Q_N(_12111_),
    .Q(\atari2600.ram[81][2] ));
 sg13g2_dfrbp_1 _27683_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1444),
    .D(_01296_),
    .Q_N(_12110_),
    .Q(\atari2600.ram[81][3] ));
 sg13g2_dfrbp_1 _27684_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1443),
    .D(_01297_),
    .Q_N(_12109_),
    .Q(\atari2600.ram[81][4] ));
 sg13g2_dfrbp_1 _27685_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1442),
    .D(_01298_),
    .Q_N(_12108_),
    .Q(\atari2600.ram[81][5] ));
 sg13g2_dfrbp_1 _27686_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1441),
    .D(_01299_),
    .Q_N(_12107_),
    .Q(\atari2600.ram[81][6] ));
 sg13g2_dfrbp_1 _27687_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1440),
    .D(_01300_),
    .Q_N(_12106_),
    .Q(\atari2600.ram[81][7] ));
 sg13g2_dfrbp_1 _27688_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1439),
    .D(_01301_),
    .Q_N(_12105_),
    .Q(\atari2600.ram[77][0] ));
 sg13g2_dfrbp_1 _27689_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1438),
    .D(_01302_),
    .Q_N(_12104_),
    .Q(\atari2600.ram[77][1] ));
 sg13g2_dfrbp_1 _27690_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1437),
    .D(_01303_),
    .Q_N(_12103_),
    .Q(\atari2600.ram[77][2] ));
 sg13g2_dfrbp_1 _27691_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1436),
    .D(_01304_),
    .Q_N(_12102_),
    .Q(\atari2600.ram[77][3] ));
 sg13g2_dfrbp_1 _27692_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1435),
    .D(_01305_),
    .Q_N(_12101_),
    .Q(\atari2600.ram[77][4] ));
 sg13g2_dfrbp_1 _27693_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1434),
    .D(_01306_),
    .Q_N(_12100_),
    .Q(\atari2600.ram[77][5] ));
 sg13g2_dfrbp_1 _27694_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1433),
    .D(_01307_),
    .Q_N(_12099_),
    .Q(\atari2600.ram[77][6] ));
 sg13g2_dfrbp_1 _27695_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1432),
    .D(_01308_),
    .Q_N(_12098_),
    .Q(\atari2600.ram[77][7] ));
 sg13g2_dfrbp_1 _27696_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1431),
    .D(_01309_),
    .Q_N(_12097_),
    .Q(\atari2600.ram[82][0] ));
 sg13g2_dfrbp_1 _27697_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1430),
    .D(_01310_),
    .Q_N(_12096_),
    .Q(\atari2600.ram[82][1] ));
 sg13g2_dfrbp_1 _27698_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1429),
    .D(_01311_),
    .Q_N(_12095_),
    .Q(\atari2600.ram[82][2] ));
 sg13g2_dfrbp_1 _27699_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1428),
    .D(_01312_),
    .Q_N(_12094_),
    .Q(\atari2600.ram[82][3] ));
 sg13g2_dfrbp_1 _27700_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1427),
    .D(_01313_),
    .Q_N(_12093_),
    .Q(\atari2600.ram[82][4] ));
 sg13g2_dfrbp_1 _27701_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1426),
    .D(_01314_),
    .Q_N(_12092_),
    .Q(\atari2600.ram[82][5] ));
 sg13g2_dfrbp_1 _27702_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1425),
    .D(_01315_),
    .Q_N(_12091_),
    .Q(\atari2600.ram[82][6] ));
 sg13g2_dfrbp_1 _27703_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1424),
    .D(_01316_),
    .Q_N(_12090_),
    .Q(\atari2600.ram[82][7] ));
 sg13g2_dfrbp_1 _27704_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1423),
    .D(_01317_),
    .Q_N(_12089_),
    .Q(\atari2600.ram[80][0] ));
 sg13g2_dfrbp_1 _27705_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1422),
    .D(_01318_),
    .Q_N(_12088_),
    .Q(\atari2600.ram[80][1] ));
 sg13g2_dfrbp_1 _27706_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1421),
    .D(_01319_),
    .Q_N(_12087_),
    .Q(\atari2600.ram[80][2] ));
 sg13g2_dfrbp_1 _27707_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1420),
    .D(_01320_),
    .Q_N(_12086_),
    .Q(\atari2600.ram[80][3] ));
 sg13g2_dfrbp_1 _27708_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1419),
    .D(_01321_),
    .Q_N(_12085_),
    .Q(\atari2600.ram[80][4] ));
 sg13g2_dfrbp_1 _27709_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1418),
    .D(_01322_),
    .Q_N(_12084_),
    .Q(\atari2600.ram[80][5] ));
 sg13g2_dfrbp_1 _27710_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1417),
    .D(_01323_),
    .Q_N(_12083_),
    .Q(\atari2600.ram[80][6] ));
 sg13g2_dfrbp_1 _27711_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1416),
    .D(_01324_),
    .Q_N(_12082_),
    .Q(\atari2600.ram[80][7] ));
 sg13g2_dfrbp_1 _27712_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1415),
    .D(_01325_),
    .Q_N(_12081_),
    .Q(\atari2600.ram[83][0] ));
 sg13g2_dfrbp_1 _27713_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1414),
    .D(_01326_),
    .Q_N(_12080_),
    .Q(\atari2600.ram[83][1] ));
 sg13g2_dfrbp_1 _27714_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1413),
    .D(_01327_),
    .Q_N(_12079_),
    .Q(\atari2600.ram[83][2] ));
 sg13g2_dfrbp_1 _27715_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1412),
    .D(_01328_),
    .Q_N(_12078_),
    .Q(\atari2600.ram[83][3] ));
 sg13g2_dfrbp_1 _27716_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1411),
    .D(_01329_),
    .Q_N(_12077_),
    .Q(\atari2600.ram[83][4] ));
 sg13g2_dfrbp_1 _27717_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1410),
    .D(_01330_),
    .Q_N(_12076_),
    .Q(\atari2600.ram[83][5] ));
 sg13g2_dfrbp_1 _27718_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1409),
    .D(_01331_),
    .Q_N(_12075_),
    .Q(\atari2600.ram[83][6] ));
 sg13g2_dfrbp_1 _27719_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1408),
    .D(_01332_),
    .Q_N(_12074_),
    .Q(\atari2600.ram[83][7] ));
 sg13g2_dfrbp_1 _27720_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1407),
    .D(_01333_),
    .Q_N(_12073_),
    .Q(\atari2600.ram[78][0] ));
 sg13g2_dfrbp_1 _27721_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1406),
    .D(_01334_),
    .Q_N(_12072_),
    .Q(\atari2600.ram[78][1] ));
 sg13g2_dfrbp_1 _27722_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1405),
    .D(_01335_),
    .Q_N(_12071_),
    .Q(\atari2600.ram[78][2] ));
 sg13g2_dfrbp_1 _27723_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1404),
    .D(_01336_),
    .Q_N(_12070_),
    .Q(\atari2600.ram[78][3] ));
 sg13g2_dfrbp_1 _27724_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1403),
    .D(_01337_),
    .Q_N(_12069_),
    .Q(\atari2600.ram[78][4] ));
 sg13g2_dfrbp_1 _27725_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1402),
    .D(_01338_),
    .Q_N(_12068_),
    .Q(\atari2600.ram[78][5] ));
 sg13g2_dfrbp_1 _27726_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1401),
    .D(_01339_),
    .Q_N(_12067_),
    .Q(\atari2600.ram[78][6] ));
 sg13g2_dfrbp_1 _27727_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1400),
    .D(_01340_),
    .Q_N(_12066_),
    .Q(\atari2600.ram[78][7] ));
 sg13g2_dfrbp_1 _27728_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1399),
    .D(_01341_),
    .Q_N(_12065_),
    .Q(\atari2600.ram[12][0] ));
 sg13g2_dfrbp_1 _27729_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1398),
    .D(_01342_),
    .Q_N(_12064_),
    .Q(\atari2600.ram[12][1] ));
 sg13g2_dfrbp_1 _27730_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1397),
    .D(_01343_),
    .Q_N(_12063_),
    .Q(\atari2600.ram[12][2] ));
 sg13g2_dfrbp_1 _27731_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1396),
    .D(_01344_),
    .Q_N(_12062_),
    .Q(\atari2600.ram[12][3] ));
 sg13g2_dfrbp_1 _27732_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1395),
    .D(_01345_),
    .Q_N(_12061_),
    .Q(\atari2600.ram[12][4] ));
 sg13g2_dfrbp_1 _27733_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1394),
    .D(_01346_),
    .Q_N(_12060_),
    .Q(\atari2600.ram[12][5] ));
 sg13g2_dfrbp_1 _27734_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1393),
    .D(_01347_),
    .Q_N(_12059_),
    .Q(\atari2600.ram[12][6] ));
 sg13g2_dfrbp_1 _27735_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1392),
    .D(_01348_),
    .Q_N(_12058_),
    .Q(\atari2600.ram[12][7] ));
 sg13g2_dfrbp_1 _27736_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1391),
    .D(net7181),
    .Q_N(_12057_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 _27737_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1390),
    .D(_01350_),
    .Q_N(_12056_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 _27738_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1389),
    .D(_01351_),
    .Q_N(_00061_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 _27739_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1388),
    .D(_01352_),
    .Q_N(_12055_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 _27740_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1387),
    .D(_01353_),
    .Q_N(_00060_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 _27741_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1386),
    .D(_01354_),
    .Q_N(_12054_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 _27742_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1385),
    .D(_01355_),
    .Q_N(_00059_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 _27743_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1384),
    .D(_01356_),
    .Q_N(_00146_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _27744_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1383),
    .D(_01357_),
    .Q_N(_12053_),
    .Q(\atari2600.ram[8][0] ));
 sg13g2_dfrbp_1 _27745_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1382),
    .D(_01358_),
    .Q_N(_12052_),
    .Q(\atari2600.ram[8][1] ));
 sg13g2_dfrbp_1 _27746_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1381),
    .D(_01359_),
    .Q_N(_12051_),
    .Q(\atari2600.ram[8][2] ));
 sg13g2_dfrbp_1 _27747_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1380),
    .D(_01360_),
    .Q_N(_12050_),
    .Q(\atari2600.ram[8][3] ));
 sg13g2_dfrbp_1 _27748_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1379),
    .D(_01361_),
    .Q_N(_12049_),
    .Q(\atari2600.ram[8][4] ));
 sg13g2_dfrbp_1 _27749_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1378),
    .D(_01362_),
    .Q_N(_12048_),
    .Q(\atari2600.ram[8][5] ));
 sg13g2_dfrbp_1 _27750_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1377),
    .D(_01363_),
    .Q_N(_12047_),
    .Q(\atari2600.ram[8][6] ));
 sg13g2_dfrbp_1 _27751_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1376),
    .D(_01364_),
    .Q_N(_12046_),
    .Q(\atari2600.ram[8][7] ));
 sg13g2_dfrbp_1 _27752_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1375),
    .D(_01365_),
    .Q_N(_12045_),
    .Q(\atari2600.cpu.ABH[0] ));
 sg13g2_dfrbp_1 _27753_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1374),
    .D(_01366_),
    .Q_N(_12044_),
    .Q(\atari2600.cpu.ABH[1] ));
 sg13g2_dfrbp_1 _27754_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1373),
    .D(_01367_),
    .Q_N(_12043_),
    .Q(\atari2600.cpu.ABH[2] ));
 sg13g2_dfrbp_1 _27755_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1372),
    .D(_01368_),
    .Q_N(_12042_),
    .Q(\atari2600.cpu.ABH[3] ));
 sg13g2_dfrbp_1 _27756_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1371),
    .D(_01369_),
    .Q_N(_12041_),
    .Q(\atari2600.cpu.ABH[4] ));
 sg13g2_dfrbp_1 _27757_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1370),
    .D(_01370_),
    .Q_N(_12040_),
    .Q(\atari2600.ram[92][0] ));
 sg13g2_dfrbp_1 _27758_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1369),
    .D(_01371_),
    .Q_N(_12039_),
    .Q(\atari2600.ram[92][1] ));
 sg13g2_dfrbp_1 _27759_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1368),
    .D(_01372_),
    .Q_N(_12038_),
    .Q(\atari2600.ram[92][2] ));
 sg13g2_dfrbp_1 _27760_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1367),
    .D(_01373_),
    .Q_N(_12037_),
    .Q(\atari2600.ram[92][3] ));
 sg13g2_dfrbp_1 _27761_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1366),
    .D(_01374_),
    .Q_N(_12036_),
    .Q(\atari2600.ram[92][4] ));
 sg13g2_dfrbp_1 _27762_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1365),
    .D(_01375_),
    .Q_N(_12035_),
    .Q(\atari2600.ram[92][5] ));
 sg13g2_dfrbp_1 _27763_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1364),
    .D(_01376_),
    .Q_N(_12034_),
    .Q(\atari2600.ram[92][6] ));
 sg13g2_dfrbp_1 _27764_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1363),
    .D(_01377_),
    .Q_N(_12033_),
    .Q(\atari2600.ram[92][7] ));
 sg13g2_dfrbp_1 _27765_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1362),
    .D(_01378_),
    .Q_N(_12032_),
    .Q(\atari2600.ram[13][0] ));
 sg13g2_dfrbp_1 _27766_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1361),
    .D(_01379_),
    .Q_N(_12031_),
    .Q(\atari2600.ram[13][1] ));
 sg13g2_dfrbp_1 _27767_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1360),
    .D(_01380_),
    .Q_N(_12030_),
    .Q(\atari2600.ram[13][2] ));
 sg13g2_dfrbp_1 _27768_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1359),
    .D(_01381_),
    .Q_N(_12029_),
    .Q(\atari2600.ram[13][3] ));
 sg13g2_dfrbp_1 _27769_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1358),
    .D(_01382_),
    .Q_N(_12028_),
    .Q(\atari2600.ram[13][4] ));
 sg13g2_dfrbp_1 _27770_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1357),
    .D(_01383_),
    .Q_N(_12027_),
    .Q(\atari2600.ram[13][5] ));
 sg13g2_dfrbp_1 _27771_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1356),
    .D(_01384_),
    .Q_N(_12026_),
    .Q(\atari2600.ram[13][6] ));
 sg13g2_dfrbp_1 _27772_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1355),
    .D(_01385_),
    .Q_N(_12025_),
    .Q(\atari2600.ram[13][7] ));
 sg13g2_dfrbp_1 _27773_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1354),
    .D(_01386_),
    .Q_N(_12024_),
    .Q(\atari2600.ram[93][0] ));
 sg13g2_dfrbp_1 _27774_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1353),
    .D(_01387_),
    .Q_N(_12023_),
    .Q(\atari2600.ram[93][1] ));
 sg13g2_dfrbp_1 _27775_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1352),
    .D(_01388_),
    .Q_N(_12022_),
    .Q(\atari2600.ram[93][2] ));
 sg13g2_dfrbp_1 _27776_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1351),
    .D(_01389_),
    .Q_N(_12021_),
    .Q(\atari2600.ram[93][3] ));
 sg13g2_dfrbp_1 _27777_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1350),
    .D(_01390_),
    .Q_N(_12020_),
    .Q(\atari2600.ram[93][4] ));
 sg13g2_dfrbp_1 _27778_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1349),
    .D(_01391_),
    .Q_N(_12019_),
    .Q(\atari2600.ram[93][5] ));
 sg13g2_dfrbp_1 _27779_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1348),
    .D(_01392_),
    .Q_N(_12018_),
    .Q(\atari2600.ram[93][6] ));
 sg13g2_dfrbp_1 _27780_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1347),
    .D(_01393_),
    .Q_N(_12017_),
    .Q(\atari2600.ram[93][7] ));
 sg13g2_dfrbp_1 _27781_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1346),
    .D(_01394_),
    .Q_N(_12016_),
    .Q(\atari2600.ram[94][0] ));
 sg13g2_dfrbp_1 _27782_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1345),
    .D(_01395_),
    .Q_N(_12015_),
    .Q(\atari2600.ram[94][1] ));
 sg13g2_dfrbp_1 _27783_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1344),
    .D(_01396_),
    .Q_N(_12014_),
    .Q(\atari2600.ram[94][2] ));
 sg13g2_dfrbp_1 _27784_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1343),
    .D(_01397_),
    .Q_N(_12013_),
    .Q(\atari2600.ram[94][3] ));
 sg13g2_dfrbp_1 _27785_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1342),
    .D(_01398_),
    .Q_N(_12012_),
    .Q(\atari2600.ram[94][4] ));
 sg13g2_dfrbp_1 _27786_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1341),
    .D(_01399_),
    .Q_N(_12011_),
    .Q(\atari2600.ram[94][5] ));
 sg13g2_dfrbp_1 _27787_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1340),
    .D(_01400_),
    .Q_N(_12010_),
    .Q(\atari2600.ram[94][6] ));
 sg13g2_dfrbp_1 _27788_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1339),
    .D(_01401_),
    .Q_N(_12009_),
    .Q(\atari2600.ram[94][7] ));
 sg13g2_dfrbp_1 _27789_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1338),
    .D(_01402_),
    .Q_N(_12008_),
    .Q(\atari2600.ram[95][0] ));
 sg13g2_dfrbp_1 _27790_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1337),
    .D(_01403_),
    .Q_N(_12007_),
    .Q(\atari2600.ram[95][1] ));
 sg13g2_dfrbp_1 _27791_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1336),
    .D(_01404_),
    .Q_N(_12006_),
    .Q(\atari2600.ram[95][2] ));
 sg13g2_dfrbp_1 _27792_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1335),
    .D(_01405_),
    .Q_N(_12005_),
    .Q(\atari2600.ram[95][3] ));
 sg13g2_dfrbp_1 _27793_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1334),
    .D(_01406_),
    .Q_N(_12004_),
    .Q(\atari2600.ram[95][4] ));
 sg13g2_dfrbp_1 _27794_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1333),
    .D(_01407_),
    .Q_N(_12003_),
    .Q(\atari2600.ram[95][5] ));
 sg13g2_dfrbp_1 _27795_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1332),
    .D(_01408_),
    .Q_N(_12002_),
    .Q(\atari2600.ram[95][6] ));
 sg13g2_dfrbp_1 _27796_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1331),
    .D(_01409_),
    .Q_N(_12001_),
    .Q(\atari2600.ram[95][7] ));
 sg13g2_dfrbp_1 _27797_ (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1330),
    .D(_01410_),
    .Q_N(_12000_),
    .Q(\atari2600.ram[96][0] ));
 sg13g2_dfrbp_1 _27798_ (.CLK(clknet_leaf_339_clk),
    .RESET_B(net1329),
    .D(_01411_),
    .Q_N(_11999_),
    .Q(\atari2600.ram[96][1] ));
 sg13g2_dfrbp_1 _27799_ (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1328),
    .D(_01412_),
    .Q_N(_11998_),
    .Q(\atari2600.ram[96][2] ));
 sg13g2_dfrbp_1 _27800_ (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1327),
    .D(_01413_),
    .Q_N(_11997_),
    .Q(\atari2600.ram[96][3] ));
 sg13g2_dfrbp_1 _27801_ (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1326),
    .D(_01414_),
    .Q_N(_11996_),
    .Q(\atari2600.ram[96][4] ));
 sg13g2_dfrbp_1 _27802_ (.CLK(clknet_leaf_339_clk),
    .RESET_B(net1325),
    .D(_01415_),
    .Q_N(_11995_),
    .Q(\atari2600.ram[96][5] ));
 sg13g2_dfrbp_1 _27803_ (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1324),
    .D(_01416_),
    .Q_N(_11994_),
    .Q(\atari2600.ram[96][6] ));
 sg13g2_dfrbp_1 _27804_ (.CLK(clknet_leaf_333_clk),
    .RESET_B(net1323),
    .D(_01417_),
    .Q_N(_11993_),
    .Q(\atari2600.ram[96][7] ));
 sg13g2_dfrbp_1 _27805_ (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1322),
    .D(_01418_),
    .Q_N(_11992_),
    .Q(\atari2600.ram[97][0] ));
 sg13g2_dfrbp_1 _27806_ (.CLK(clknet_leaf_338_clk),
    .RESET_B(net1321),
    .D(_01419_),
    .Q_N(_11991_),
    .Q(\atari2600.ram[97][1] ));
 sg13g2_dfrbp_1 _27807_ (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1320),
    .D(_01420_),
    .Q_N(_11990_),
    .Q(\atari2600.ram[97][2] ));
 sg13g2_dfrbp_1 _27808_ (.CLK(clknet_leaf_336_clk),
    .RESET_B(net1319),
    .D(_01421_),
    .Q_N(_11989_),
    .Q(\atari2600.ram[97][3] ));
 sg13g2_dfrbp_1 _27809_ (.CLK(clknet_leaf_330_clk),
    .RESET_B(net1318),
    .D(_01422_),
    .Q_N(_11988_),
    .Q(\atari2600.ram[97][4] ));
 sg13g2_dfrbp_1 _27810_ (.CLK(clknet_leaf_337_clk),
    .RESET_B(net1317),
    .D(_01423_),
    .Q_N(_11987_),
    .Q(\atari2600.ram[97][5] ));
 sg13g2_dfrbp_1 _27811_ (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1316),
    .D(_01424_),
    .Q_N(_11986_),
    .Q(\atari2600.ram[97][6] ));
 sg13g2_dfrbp_1 _27812_ (.CLK(clknet_leaf_336_clk),
    .RESET_B(net1315),
    .D(_01425_),
    .Q_N(_11985_),
    .Q(\atari2600.ram[97][7] ));
 sg13g2_dfrbp_1 _27813_ (.CLK(clknet_leaf_336_clk),
    .RESET_B(net1314),
    .D(_01426_),
    .Q_N(_11984_),
    .Q(\atari2600.ram[98][0] ));
 sg13g2_dfrbp_1 _27814_ (.CLK(clknet_leaf_337_clk),
    .RESET_B(net1313),
    .D(_01427_),
    .Q_N(_11983_),
    .Q(\atari2600.ram[98][1] ));
 sg13g2_dfrbp_1 _27815_ (.CLK(clknet_leaf_336_clk),
    .RESET_B(net1312),
    .D(_01428_),
    .Q_N(_11982_),
    .Q(\atari2600.ram[98][2] ));
 sg13g2_dfrbp_1 _27816_ (.CLK(clknet_leaf_336_clk),
    .RESET_B(net1311),
    .D(_01429_),
    .Q_N(_11981_),
    .Q(\atari2600.ram[98][3] ));
 sg13g2_dfrbp_1 _27817_ (.CLK(clknet_leaf_329_clk),
    .RESET_B(net1310),
    .D(_01430_),
    .Q_N(_11980_),
    .Q(\atari2600.ram[98][4] ));
 sg13g2_dfrbp_1 _27818_ (.CLK(clknet_leaf_337_clk),
    .RESET_B(net1309),
    .D(_01431_),
    .Q_N(_11979_),
    .Q(\atari2600.ram[98][5] ));
 sg13g2_dfrbp_1 _27819_ (.CLK(clknet_leaf_336_clk),
    .RESET_B(net1308),
    .D(_01432_),
    .Q_N(_11978_),
    .Q(\atari2600.ram[98][6] ));
 sg13g2_dfrbp_1 _27820_ (.CLK(clknet_leaf_336_clk),
    .RESET_B(net1307),
    .D(_01433_),
    .Q_N(_11977_),
    .Q(\atari2600.ram[98][7] ));
 sg13g2_dfrbp_1 _27821_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1306),
    .D(_01434_),
    .Q_N(_11976_),
    .Q(\atari2600.ram[0][0] ));
 sg13g2_dfrbp_1 _27822_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1305),
    .D(_01435_),
    .Q_N(_11975_),
    .Q(\atari2600.ram[0][1] ));
 sg13g2_dfrbp_1 _27823_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1304),
    .D(_01436_),
    .Q_N(_11974_),
    .Q(\atari2600.ram[0][2] ));
 sg13g2_dfrbp_1 _27824_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1303),
    .D(_01437_),
    .Q_N(_11973_),
    .Q(\atari2600.ram[0][3] ));
 sg13g2_dfrbp_1 _27825_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1302),
    .D(_01438_),
    .Q_N(_11972_),
    .Q(\atari2600.ram[0][4] ));
 sg13g2_dfrbp_1 _27826_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1301),
    .D(_01439_),
    .Q_N(_11971_),
    .Q(\atari2600.ram[0][5] ));
 sg13g2_dfrbp_1 _27827_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1300),
    .D(_01440_),
    .Q_N(_11970_),
    .Q(\atari2600.ram[0][6] ));
 sg13g2_dfrbp_1 _27828_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1299),
    .D(_01441_),
    .Q_N(_11969_),
    .Q(\atari2600.ram[0][7] ));
 sg13g2_dfrbp_1 _27829_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1298),
    .D(_01442_),
    .Q_N(_11968_),
    .Q(\atari2600.ram[100][0] ));
 sg13g2_dfrbp_1 _27830_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1297),
    .D(_01443_),
    .Q_N(_11967_),
    .Q(\atari2600.ram[100][1] ));
 sg13g2_dfrbp_1 _27831_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1296),
    .D(_01444_),
    .Q_N(_11966_),
    .Q(\atari2600.ram[100][2] ));
 sg13g2_dfrbp_1 _27832_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1295),
    .D(_01445_),
    .Q_N(_11965_),
    .Q(\atari2600.ram[100][3] ));
 sg13g2_dfrbp_1 _27833_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1294),
    .D(_01446_),
    .Q_N(_11964_),
    .Q(\atari2600.ram[100][4] ));
 sg13g2_dfrbp_1 _27834_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1293),
    .D(_01447_),
    .Q_N(_11963_),
    .Q(\atari2600.ram[100][5] ));
 sg13g2_dfrbp_1 _27835_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1292),
    .D(_01448_),
    .Q_N(_11962_),
    .Q(\atari2600.ram[100][6] ));
 sg13g2_dfrbp_1 _27836_ (.CLK(clknet_leaf_329_clk),
    .RESET_B(net1291),
    .D(_01449_),
    .Q_N(_11961_),
    .Q(\atari2600.ram[100][7] ));
 sg13g2_dfrbp_1 _27837_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1290),
    .D(_01450_),
    .Q_N(_11960_),
    .Q(\atari2600.ram[101][0] ));
 sg13g2_dfrbp_1 _27838_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1289),
    .D(_01451_),
    .Q_N(_11959_),
    .Q(\atari2600.ram[101][1] ));
 sg13g2_dfrbp_1 _27839_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1288),
    .D(_01452_),
    .Q_N(_11958_),
    .Q(\atari2600.ram[101][2] ));
 sg13g2_dfrbp_1 _27840_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1287),
    .D(_01453_),
    .Q_N(_11957_),
    .Q(\atari2600.ram[101][3] ));
 sg13g2_dfrbp_1 _27841_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1286),
    .D(_01454_),
    .Q_N(_11956_),
    .Q(\atari2600.ram[101][4] ));
 sg13g2_dfrbp_1 _27842_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1285),
    .D(_01455_),
    .Q_N(_11955_),
    .Q(\atari2600.ram[101][5] ));
 sg13g2_dfrbp_1 _27843_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1284),
    .D(_01456_),
    .Q_N(_11954_),
    .Q(\atari2600.ram[101][6] ));
 sg13g2_dfrbp_1 _27844_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1283),
    .D(_01457_),
    .Q_N(_11953_),
    .Q(\atari2600.ram[101][7] ));
 sg13g2_dfrbp_1 _27845_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1282),
    .D(_01458_),
    .Q_N(_11952_),
    .Q(\atari2600.ram[102][0] ));
 sg13g2_dfrbp_1 _27846_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1281),
    .D(_01459_),
    .Q_N(_11951_),
    .Q(\atari2600.ram[102][1] ));
 sg13g2_dfrbp_1 _27847_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1280),
    .D(_01460_),
    .Q_N(_11950_),
    .Q(\atari2600.ram[102][2] ));
 sg13g2_dfrbp_1 _27848_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1279),
    .D(_01461_),
    .Q_N(_11949_),
    .Q(\atari2600.ram[102][3] ));
 sg13g2_dfrbp_1 _27849_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1278),
    .D(_01462_),
    .Q_N(_11948_),
    .Q(\atari2600.ram[102][4] ));
 sg13g2_dfrbp_1 _27850_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1277),
    .D(_01463_),
    .Q_N(_11947_),
    .Q(\atari2600.ram[102][5] ));
 sg13g2_dfrbp_1 _27851_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1276),
    .D(_01464_),
    .Q_N(_11946_),
    .Q(\atari2600.ram[102][6] ));
 sg13g2_dfrbp_1 _27852_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1275),
    .D(_01465_),
    .Q_N(_11945_),
    .Q(\atari2600.ram[102][7] ));
 sg13g2_dfrbp_1 _27853_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1274),
    .D(_01466_),
    .Q_N(_11944_),
    .Q(\atari2600.ram[103][0] ));
 sg13g2_dfrbp_1 _27854_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1273),
    .D(_01467_),
    .Q_N(_11943_),
    .Q(\atari2600.ram[103][1] ));
 sg13g2_dfrbp_1 _27855_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1272),
    .D(_01468_),
    .Q_N(_11942_),
    .Q(\atari2600.ram[103][2] ));
 sg13g2_dfrbp_1 _27856_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1271),
    .D(_01469_),
    .Q_N(_11941_),
    .Q(\atari2600.ram[103][3] ));
 sg13g2_dfrbp_1 _27857_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1270),
    .D(_01470_),
    .Q_N(_11940_),
    .Q(\atari2600.ram[103][4] ));
 sg13g2_dfrbp_1 _27858_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1269),
    .D(_01471_),
    .Q_N(_11939_),
    .Q(\atari2600.ram[103][5] ));
 sg13g2_dfrbp_1 _27859_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1268),
    .D(_01472_),
    .Q_N(_11938_),
    .Q(\atari2600.ram[103][6] ));
 sg13g2_dfrbp_1 _27860_ (.CLK(clknet_leaf_329_clk),
    .RESET_B(net1267),
    .D(_01473_),
    .Q_N(_11937_),
    .Q(\atari2600.ram[103][7] ));
 sg13g2_dfrbp_1 _27861_ (.CLK(clknet_leaf_337_clk),
    .RESET_B(net1266),
    .D(_01474_),
    .Q_N(_11936_),
    .Q(\atari2600.ram[104][0] ));
 sg13g2_dfrbp_1 _27862_ (.CLK(clknet_leaf_332_clk),
    .RESET_B(net1265),
    .D(_01475_),
    .Q_N(_11935_),
    .Q(\atari2600.ram[104][1] ));
 sg13g2_dfrbp_1 _27863_ (.CLK(clknet_leaf_337_clk),
    .RESET_B(net1264),
    .D(_01476_),
    .Q_N(_11934_),
    .Q(\atari2600.ram[104][2] ));
 sg13g2_dfrbp_1 _27864_ (.CLK(clknet_leaf_330_clk),
    .RESET_B(net1263),
    .D(_01477_),
    .Q_N(_11933_),
    .Q(\atari2600.ram[104][3] ));
 sg13g2_dfrbp_1 _27865_ (.CLK(clknet_leaf_329_clk),
    .RESET_B(net1262),
    .D(_01478_),
    .Q_N(_11932_),
    .Q(\atari2600.ram[104][4] ));
 sg13g2_dfrbp_1 _27866_ (.CLK(clknet_leaf_329_clk),
    .RESET_B(net1261),
    .D(_01479_),
    .Q_N(_11931_),
    .Q(\atari2600.ram[104][5] ));
 sg13g2_dfrbp_1 _27867_ (.CLK(clknet_leaf_330_clk),
    .RESET_B(net1260),
    .D(_01480_),
    .Q_N(_11930_),
    .Q(\atari2600.ram[104][6] ));
 sg13g2_dfrbp_1 _27868_ (.CLK(clknet_leaf_330_clk),
    .RESET_B(net1259),
    .D(_01481_),
    .Q_N(_11929_),
    .Q(\atari2600.ram[104][7] ));
 sg13g2_dfrbp_1 _27869_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1258),
    .D(_01482_),
    .Q_N(_11928_),
    .Q(\atari2600.ram[105][0] ));
 sg13g2_dfrbp_1 _27870_ (.CLK(clknet_leaf_328_clk),
    .RESET_B(net1257),
    .D(_01483_),
    .Q_N(_11927_),
    .Q(\atari2600.ram[105][1] ));
 sg13g2_dfrbp_1 _27871_ (.CLK(clknet_leaf_329_clk),
    .RESET_B(net1256),
    .D(_01484_),
    .Q_N(_11926_),
    .Q(\atari2600.ram[105][2] ));
 sg13g2_dfrbp_1 _27872_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1255),
    .D(_01485_),
    .Q_N(_11925_),
    .Q(\atari2600.ram[105][3] ));
 sg13g2_dfrbp_1 _27873_ (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1254),
    .D(_01486_),
    .Q_N(_11924_),
    .Q(\atari2600.ram[105][4] ));
 sg13g2_dfrbp_1 _27874_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1253),
    .D(_01487_),
    .Q_N(_11923_),
    .Q(\atari2600.ram[105][5] ));
 sg13g2_dfrbp_1 _27875_ (.CLK(clknet_leaf_330_clk),
    .RESET_B(net1252),
    .D(_01488_),
    .Q_N(_11922_),
    .Q(\atari2600.ram[105][6] ));
 sg13g2_dfrbp_1 _27876_ (.CLK(clknet_leaf_327_clk),
    .RESET_B(net1251),
    .D(_01489_),
    .Q_N(_11921_),
    .Q(\atari2600.ram[105][7] ));
 sg13g2_dfrbp_1 _27877_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1250),
    .D(_01490_),
    .Q_N(_11920_),
    .Q(\atari2600.ram[106][0] ));
 sg13g2_dfrbp_1 _27878_ (.CLK(clknet_leaf_328_clk),
    .RESET_B(net1249),
    .D(_01491_),
    .Q_N(_11919_),
    .Q(\atari2600.ram[106][1] ));
 sg13g2_dfrbp_1 _27879_ (.CLK(clknet_leaf_329_clk),
    .RESET_B(net1248),
    .D(_01492_),
    .Q_N(_11918_),
    .Q(\atari2600.ram[106][2] ));
 sg13g2_dfrbp_1 _27880_ (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1247),
    .D(_01493_),
    .Q_N(_11917_),
    .Q(\atari2600.ram[106][3] ));
 sg13g2_dfrbp_1 _27881_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1246),
    .D(_01494_),
    .Q_N(_11916_),
    .Q(\atari2600.ram[106][4] ));
 sg13g2_dfrbp_1 _27882_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1245),
    .D(_01495_),
    .Q_N(_11915_),
    .Q(\atari2600.ram[106][5] ));
 sg13g2_dfrbp_1 _27883_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1244),
    .D(_01496_),
    .Q_N(_11914_),
    .Q(\atari2600.ram[106][6] ));
 sg13g2_dfrbp_1 _27884_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1243),
    .D(_01497_),
    .Q_N(_11913_),
    .Q(\atari2600.ram[106][7] ));
 sg13g2_dfrbp_1 _27885_ (.CLK(clknet_leaf_337_clk),
    .RESET_B(net1242),
    .D(_01498_),
    .Q_N(_11912_),
    .Q(\atari2600.ram[107][0] ));
 sg13g2_dfrbp_1 _27886_ (.CLK(clknet_leaf_332_clk),
    .RESET_B(net1241),
    .D(_01499_),
    .Q_N(_11911_),
    .Q(\atari2600.ram[107][1] ));
 sg13g2_dfrbp_1 _27887_ (.CLK(clknet_leaf_336_clk),
    .RESET_B(net1232),
    .D(_01500_),
    .Q_N(_11910_),
    .Q(\atari2600.ram[107][2] ));
 sg13g2_dfrbp_1 _27888_ (.CLK(clknet_leaf_330_clk),
    .RESET_B(net1231),
    .D(_01501_),
    .Q_N(_11909_),
    .Q(\atari2600.ram[107][3] ));
 sg13g2_dfrbp_1 _27889_ (.CLK(clknet_leaf_328_clk),
    .RESET_B(net1230),
    .D(_01502_),
    .Q_N(_11908_),
    .Q(\atari2600.ram[107][4] ));
 sg13g2_dfrbp_1 _27890_ (.CLK(clknet_leaf_337_clk),
    .RESET_B(net1229),
    .D(_01503_),
    .Q_N(_11907_),
    .Q(\atari2600.ram[107][5] ));
 sg13g2_dfrbp_1 _27891_ (.CLK(clknet_leaf_330_clk),
    .RESET_B(net1228),
    .D(_01504_),
    .Q_N(_11906_),
    .Q(\atari2600.ram[107][6] ));
 sg13g2_dfrbp_1 _27892_ (.CLK(clknet_leaf_331_clk),
    .RESET_B(net1227),
    .D(_01505_),
    .Q_N(_11905_),
    .Q(\atari2600.ram[107][7] ));
 sg13g2_dfrbp_1 _27893_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1226),
    .D(_01506_),
    .Q_N(_11904_),
    .Q(\atari2600.ram[108][0] ));
 sg13g2_dfrbp_1 _27894_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1225),
    .D(_01507_),
    .Q_N(_11903_),
    .Q(\atari2600.ram[108][1] ));
 sg13g2_dfrbp_1 _27895_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1224),
    .D(_01508_),
    .Q_N(_11902_),
    .Q(\atari2600.ram[108][2] ));
 sg13g2_dfrbp_1 _27896_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1223),
    .D(_01509_),
    .Q_N(_11901_),
    .Q(\atari2600.ram[108][3] ));
 sg13g2_dfrbp_1 _27897_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1222),
    .D(_01510_),
    .Q_N(_11900_),
    .Q(\atari2600.ram[108][4] ));
 sg13g2_dfrbp_1 _27898_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1221),
    .D(_01511_),
    .Q_N(_11899_),
    .Q(\atari2600.ram[108][5] ));
 sg13g2_dfrbp_1 _27899_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1220),
    .D(_01512_),
    .Q_N(_11898_),
    .Q(\atari2600.ram[108][6] ));
 sg13g2_dfrbp_1 _27900_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1219),
    .D(_01513_),
    .Q_N(_11897_),
    .Q(\atari2600.ram[108][7] ));
 sg13g2_dfrbp_1 _27901_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1218),
    .D(_01514_),
    .Q_N(_11896_),
    .Q(\atari2600.ram[10][0] ));
 sg13g2_dfrbp_1 _27902_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1217),
    .D(_01515_),
    .Q_N(_11895_),
    .Q(\atari2600.ram[10][1] ));
 sg13g2_dfrbp_1 _27903_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1216),
    .D(_01516_),
    .Q_N(_11894_),
    .Q(\atari2600.ram[10][2] ));
 sg13g2_dfrbp_1 _27904_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1215),
    .D(_01517_),
    .Q_N(_11893_),
    .Q(\atari2600.ram[10][3] ));
 sg13g2_dfrbp_1 _27905_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1214),
    .D(_01518_),
    .Q_N(_11892_),
    .Q(\atari2600.ram[10][4] ));
 sg13g2_dfrbp_1 _27906_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1213),
    .D(_01519_),
    .Q_N(_11891_),
    .Q(\atari2600.ram[10][5] ));
 sg13g2_dfrbp_1 _27907_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1212),
    .D(_01520_),
    .Q_N(_11890_),
    .Q(\atari2600.ram[10][6] ));
 sg13g2_dfrbp_1 _27908_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1211),
    .D(_01521_),
    .Q_N(_11889_),
    .Q(\atari2600.ram[10][7] ));
 sg13g2_dfrbp_1 _27909_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1210),
    .D(_01522_),
    .Q_N(_11888_),
    .Q(\atari2600.ram[110][0] ));
 sg13g2_dfrbp_1 _27910_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1209),
    .D(_01523_),
    .Q_N(_11887_),
    .Q(\atari2600.ram[110][1] ));
 sg13g2_dfrbp_1 _27911_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1208),
    .D(_01524_),
    .Q_N(_11886_),
    .Q(\atari2600.ram[110][2] ));
 sg13g2_dfrbp_1 _27912_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1207),
    .D(_01525_),
    .Q_N(_11885_),
    .Q(\atari2600.ram[110][3] ));
 sg13g2_dfrbp_1 _27913_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1206),
    .D(_01526_),
    .Q_N(_11884_),
    .Q(\atari2600.ram[110][4] ));
 sg13g2_dfrbp_1 _27914_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1205),
    .D(_01527_),
    .Q_N(_11883_),
    .Q(\atari2600.ram[110][5] ));
 sg13g2_dfrbp_1 _27915_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1204),
    .D(_01528_),
    .Q_N(_11882_),
    .Q(\atari2600.ram[110][6] ));
 sg13g2_dfrbp_1 _27916_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1203),
    .D(_01529_),
    .Q_N(_11881_),
    .Q(\atari2600.ram[110][7] ));
 sg13g2_dfrbp_1 _27917_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1202),
    .D(_01530_),
    .Q_N(_11880_),
    .Q(\atari2600.ram[111][0] ));
 sg13g2_dfrbp_1 _27918_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1201),
    .D(_01531_),
    .Q_N(_11879_),
    .Q(\atari2600.ram[111][1] ));
 sg13g2_dfrbp_1 _27919_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1200),
    .D(_01532_),
    .Q_N(_11878_),
    .Q(\atari2600.ram[111][2] ));
 sg13g2_dfrbp_1 _27920_ (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1199),
    .D(_01533_),
    .Q_N(_11877_),
    .Q(\atari2600.ram[111][3] ));
 sg13g2_dfrbp_1 _27921_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1198),
    .D(_01534_),
    .Q_N(_11876_),
    .Q(\atari2600.ram[111][4] ));
 sg13g2_dfrbp_1 _27922_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1197),
    .D(_01535_),
    .Q_N(_11875_),
    .Q(\atari2600.ram[111][5] ));
 sg13g2_dfrbp_1 _27923_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1196),
    .D(_01536_),
    .Q_N(_11874_),
    .Q(\atari2600.ram[111][6] ));
 sg13g2_dfrbp_1 _27924_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1195),
    .D(_01537_),
    .Q_N(_11873_),
    .Q(\atari2600.ram[111][7] ));
 sg13g2_dfrbp_1 _27925_ (.CLK(clknet_leaf_339_clk),
    .RESET_B(net1194),
    .D(_01538_),
    .Q_N(_11872_),
    .Q(\atari2600.ram[112][0] ));
 sg13g2_dfrbp_1 _27926_ (.CLK(clknet_leaf_339_clk),
    .RESET_B(net1193),
    .D(_01539_),
    .Q_N(_11871_),
    .Q(\atari2600.ram[112][1] ));
 sg13g2_dfrbp_1 _27927_ (.CLK(clknet_leaf_339_clk),
    .RESET_B(net1192),
    .D(_01540_),
    .Q_N(_11870_),
    .Q(\atari2600.ram[112][2] ));
 sg13g2_dfrbp_1 _27928_ (.CLK(clknet_leaf_345_clk),
    .RESET_B(net1191),
    .D(_01541_),
    .Q_N(_11869_),
    .Q(\atari2600.ram[112][3] ));
 sg13g2_dfrbp_1 _27929_ (.CLK(clknet_leaf_338_clk),
    .RESET_B(net1190),
    .D(_01542_),
    .Q_N(_11868_),
    .Q(\atari2600.ram[112][4] ));
 sg13g2_dfrbp_1 _27930_ (.CLK(clknet_leaf_344_clk),
    .RESET_B(net1189),
    .D(_01543_),
    .Q_N(_11867_),
    .Q(\atari2600.ram[112][5] ));
 sg13g2_dfrbp_1 _27931_ (.CLK(clknet_leaf_344_clk),
    .RESET_B(net1188),
    .D(_01544_),
    .Q_N(_11866_),
    .Q(\atari2600.ram[112][6] ));
 sg13g2_dfrbp_1 _27932_ (.CLK(clknet_leaf_338_clk),
    .RESET_B(net1187),
    .D(_01545_),
    .Q_N(_11865_),
    .Q(\atari2600.ram[112][7] ));
 sg13g2_dfrbp_1 _27933_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1186),
    .D(_01546_),
    .Q_N(_11864_),
    .Q(\atari2600.ram[113][0] ));
 sg13g2_dfrbp_1 _27934_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1185),
    .D(_01547_),
    .Q_N(_11863_),
    .Q(\atari2600.ram[113][1] ));
 sg13g2_dfrbp_1 _27935_ (.CLK(clknet_leaf_338_clk),
    .RESET_B(net1184),
    .D(_01548_),
    .Q_N(_11862_),
    .Q(\atari2600.ram[113][2] ));
 sg13g2_dfrbp_1 _27936_ (.CLK(clknet_leaf_345_clk),
    .RESET_B(net1183),
    .D(_01549_),
    .Q_N(_11861_),
    .Q(\atari2600.ram[113][3] ));
 sg13g2_dfrbp_1 _27937_ (.CLK(clknet_leaf_345_clk),
    .RESET_B(net1182),
    .D(_01550_),
    .Q_N(_11860_),
    .Q(\atari2600.ram[113][4] ));
 sg13g2_dfrbp_1 _27938_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1181),
    .D(_01551_),
    .Q_N(_11859_),
    .Q(\atari2600.ram[113][5] ));
 sg13g2_dfrbp_1 _27939_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1180),
    .D(_01552_),
    .Q_N(_11858_),
    .Q(\atari2600.ram[113][6] ));
 sg13g2_dfrbp_1 _27940_ (.CLK(clknet_leaf_337_clk),
    .RESET_B(net1179),
    .D(_01553_),
    .Q_N(_11857_),
    .Q(\atari2600.ram[113][7] ));
 sg13g2_dfrbp_1 _27941_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1178),
    .D(_01554_),
    .Q_N(_11856_),
    .Q(\atari2600.ram[114][0] ));
 sg13g2_dfrbp_1 _27942_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1177),
    .D(_01555_),
    .Q_N(_11855_),
    .Q(\atari2600.ram[114][1] ));
 sg13g2_dfrbp_1 _27943_ (.CLK(clknet_leaf_344_clk),
    .RESET_B(net1176),
    .D(_01556_),
    .Q_N(_11854_),
    .Q(\atari2600.ram[114][2] ));
 sg13g2_dfrbp_1 _27944_ (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1175),
    .D(_01557_),
    .Q_N(_11853_),
    .Q(\atari2600.ram[114][3] ));
 sg13g2_dfrbp_1 _27945_ (.CLK(clknet_leaf_345_clk),
    .RESET_B(net1174),
    .D(_01558_),
    .Q_N(_11852_),
    .Q(\atari2600.ram[114][4] ));
 sg13g2_dfrbp_1 _27946_ (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1173),
    .D(_01559_),
    .Q_N(_11851_),
    .Q(\atari2600.ram[114][5] ));
 sg13g2_dfrbp_1 _27947_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1172),
    .D(_01560_),
    .Q_N(_11850_),
    .Q(\atari2600.ram[114][6] ));
 sg13g2_dfrbp_1 _27948_ (.CLK(clknet_leaf_345_clk),
    .RESET_B(net1171),
    .D(_01561_),
    .Q_N(_11849_),
    .Q(\atari2600.ram[114][7] ));
 sg13g2_dfrbp_1 _27949_ (.CLK(clknet_leaf_339_clk),
    .RESET_B(net1170),
    .D(_01562_),
    .Q_N(_11848_),
    .Q(\atari2600.ram[115][0] ));
 sg13g2_dfrbp_1 _27950_ (.CLK(clknet_leaf_339_clk),
    .RESET_B(net1169),
    .D(_01563_),
    .Q_N(_11847_),
    .Q(\atari2600.ram[115][1] ));
 sg13g2_dfrbp_1 _27951_ (.CLK(clknet_leaf_338_clk),
    .RESET_B(net1168),
    .D(_01564_),
    .Q_N(_11846_),
    .Q(\atari2600.ram[115][2] ));
 sg13g2_dfrbp_1 _27952_ (.CLK(clknet_leaf_344_clk),
    .RESET_B(net1167),
    .D(_01565_),
    .Q_N(_11845_),
    .Q(\atari2600.ram[115][3] ));
 sg13g2_dfrbp_1 _27953_ (.CLK(clknet_leaf_338_clk),
    .RESET_B(net1166),
    .D(_01566_),
    .Q_N(_11844_),
    .Q(\atari2600.ram[115][4] ));
 sg13g2_dfrbp_1 _27954_ (.CLK(clknet_leaf_345_clk),
    .RESET_B(net1165),
    .D(_01567_),
    .Q_N(_11843_),
    .Q(\atari2600.ram[115][5] ));
 sg13g2_dfrbp_1 _27955_ (.CLK(clknet_leaf_344_clk),
    .RESET_B(net1164),
    .D(_01568_),
    .Q_N(_11842_),
    .Q(\atari2600.ram[115][6] ));
 sg13g2_dfrbp_1 _27956_ (.CLK(clknet_leaf_338_clk),
    .RESET_B(net1163),
    .D(_01569_),
    .Q_N(_11841_),
    .Q(\atari2600.ram[115][7] ));
 sg13g2_dfrbp_1 _27957_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1162),
    .D(_01570_),
    .Q_N(_11840_),
    .Q(\atari2600.ram[116][0] ));
 sg13g2_dfrbp_1 _27958_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1161),
    .D(_01571_),
    .Q_N(_11839_),
    .Q(\atari2600.ram[116][1] ));
 sg13g2_dfrbp_1 _27959_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1160),
    .D(_01572_),
    .Q_N(_11838_),
    .Q(\atari2600.ram[116][2] ));
 sg13g2_dfrbp_1 _27960_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1159),
    .D(_01573_),
    .Q_N(_11837_),
    .Q(\atari2600.ram[116][3] ));
 sg13g2_dfrbp_1 _27961_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1158),
    .D(_01574_),
    .Q_N(_11836_),
    .Q(\atari2600.ram[116][4] ));
 sg13g2_dfrbp_1 _27962_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1157),
    .D(_01575_),
    .Q_N(_11835_),
    .Q(\atari2600.ram[116][5] ));
 sg13g2_dfrbp_1 _27963_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1156),
    .D(_01576_),
    .Q_N(_11834_),
    .Q(\atari2600.ram[116][6] ));
 sg13g2_dfrbp_1 _27964_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1155),
    .D(_01577_),
    .Q_N(_11833_),
    .Q(\atari2600.ram[116][7] ));
 sg13g2_dfrbp_1 _27965_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1154),
    .D(_01578_),
    .Q_N(_11832_),
    .Q(\atari2600.ram[117][0] ));
 sg13g2_dfrbp_1 _27966_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1153),
    .D(_01579_),
    .Q_N(_11831_),
    .Q(\atari2600.ram[117][1] ));
 sg13g2_dfrbp_1 _27967_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1152),
    .D(_01580_),
    .Q_N(_11830_),
    .Q(\atari2600.ram[117][2] ));
 sg13g2_dfrbp_1 _27968_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1151),
    .D(_01581_),
    .Q_N(_11829_),
    .Q(\atari2600.ram[117][3] ));
 sg13g2_dfrbp_1 _27969_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1150),
    .D(_01582_),
    .Q_N(_11828_),
    .Q(\atari2600.ram[117][4] ));
 sg13g2_dfrbp_1 _27970_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1149),
    .D(_01583_),
    .Q_N(_11827_),
    .Q(\atari2600.ram[117][5] ));
 sg13g2_dfrbp_1 _27971_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1148),
    .D(_01584_),
    .Q_N(_11826_),
    .Q(\atari2600.ram[117][6] ));
 sg13g2_dfrbp_1 _27972_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1147),
    .D(_01585_),
    .Q_N(_11825_),
    .Q(\atari2600.ram[117][7] ));
 sg13g2_dfrbp_1 _27973_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1146),
    .D(_01586_),
    .Q_N(_11824_),
    .Q(\atari2600.ram[118][0] ));
 sg13g2_dfrbp_1 _27974_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1145),
    .D(_01587_),
    .Q_N(_11823_),
    .Q(\atari2600.ram[118][1] ));
 sg13g2_dfrbp_1 _27975_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1144),
    .D(_01588_),
    .Q_N(_11822_),
    .Q(\atari2600.ram[118][2] ));
 sg13g2_dfrbp_1 _27976_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1143),
    .D(_01589_),
    .Q_N(_11821_),
    .Q(\atari2600.ram[118][3] ));
 sg13g2_dfrbp_1 _27977_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1142),
    .D(_01590_),
    .Q_N(_11820_),
    .Q(\atari2600.ram[118][4] ));
 sg13g2_dfrbp_1 _27978_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1141),
    .D(_01591_),
    .Q_N(_11819_),
    .Q(\atari2600.ram[118][5] ));
 sg13g2_dfrbp_1 _27979_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1140),
    .D(_01592_),
    .Q_N(_11818_),
    .Q(\atari2600.ram[118][6] ));
 sg13g2_dfrbp_1 _27980_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1139),
    .D(_01593_),
    .Q_N(_11817_),
    .Q(\atari2600.ram[118][7] ));
 sg13g2_dfrbp_1 _27981_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1138),
    .D(_01594_),
    .Q_N(_11816_),
    .Q(\atari2600.ram[11][0] ));
 sg13g2_dfrbp_1 _27982_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1137),
    .D(_01595_),
    .Q_N(_11815_),
    .Q(\atari2600.ram[11][1] ));
 sg13g2_dfrbp_1 _27983_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1136),
    .D(_01596_),
    .Q_N(_11814_),
    .Q(\atari2600.ram[11][2] ));
 sg13g2_dfrbp_1 _27984_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1135),
    .D(_01597_),
    .Q_N(_11813_),
    .Q(\atari2600.ram[11][3] ));
 sg13g2_dfrbp_1 _27985_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1134),
    .D(_01598_),
    .Q_N(_11812_),
    .Q(\atari2600.ram[11][4] ));
 sg13g2_dfrbp_1 _27986_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1133),
    .D(_01599_),
    .Q_N(_11811_),
    .Q(\atari2600.ram[11][5] ));
 sg13g2_dfrbp_1 _27987_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1132),
    .D(_01600_),
    .Q_N(_11810_),
    .Q(\atari2600.ram[11][6] ));
 sg13g2_dfrbp_1 _27988_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1131),
    .D(_01601_),
    .Q_N(_11809_),
    .Q(\atari2600.ram[11][7] ));
 sg13g2_dfrbp_1 _27989_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1130),
    .D(_01602_),
    .Q_N(_11808_),
    .Q(\atari2600.ram[120][0] ));
 sg13g2_dfrbp_1 _27990_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1129),
    .D(_01603_),
    .Q_N(_11807_),
    .Q(\atari2600.ram[120][1] ));
 sg13g2_dfrbp_1 _27991_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1128),
    .D(_01604_),
    .Q_N(_11806_),
    .Q(\atari2600.ram[120][2] ));
 sg13g2_dfrbp_1 _27992_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1127),
    .D(_01605_),
    .Q_N(_11805_),
    .Q(\atari2600.ram[120][3] ));
 sg13g2_dfrbp_1 _27993_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1126),
    .D(_01606_),
    .Q_N(_11804_),
    .Q(\atari2600.ram[120][4] ));
 sg13g2_dfrbp_1 _27994_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1125),
    .D(_01607_),
    .Q_N(_11803_),
    .Q(\atari2600.ram[120][5] ));
 sg13g2_dfrbp_1 _27995_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1124),
    .D(_01608_),
    .Q_N(_11802_),
    .Q(\atari2600.ram[120][6] ));
 sg13g2_dfrbp_1 _27996_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1123),
    .D(_01609_),
    .Q_N(_11801_),
    .Q(\atari2600.ram[120][7] ));
 sg13g2_dfrbp_1 _27997_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1122),
    .D(_01610_),
    .Q_N(_11800_),
    .Q(\atari2600.ram[123][0] ));
 sg13g2_dfrbp_1 _27998_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1121),
    .D(_01611_),
    .Q_N(_11799_),
    .Q(\atari2600.ram[123][1] ));
 sg13g2_dfrbp_1 _27999_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1120),
    .D(_01612_),
    .Q_N(_11798_),
    .Q(\atari2600.ram[123][2] ));
 sg13g2_dfrbp_1 _28000_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1119),
    .D(_01613_),
    .Q_N(_11797_),
    .Q(\atari2600.ram[123][3] ));
 sg13g2_dfrbp_1 _28001_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1118),
    .D(_01614_),
    .Q_N(_11796_),
    .Q(\atari2600.ram[123][4] ));
 sg13g2_dfrbp_1 _28002_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1117),
    .D(_01615_),
    .Q_N(_11795_),
    .Q(\atari2600.ram[123][5] ));
 sg13g2_dfrbp_1 _28003_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1116),
    .D(_01616_),
    .Q_N(_11794_),
    .Q(\atari2600.ram[123][6] ));
 sg13g2_dfrbp_1 _28004_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1115),
    .D(_01617_),
    .Q_N(_11793_),
    .Q(\atari2600.ram[123][7] ));
 sg13g2_dfrbp_1 _28005_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1114),
    .D(_01618_),
    .Q_N(_11792_),
    .Q(\atari2600.ram[121][0] ));
 sg13g2_dfrbp_1 _28006_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1113),
    .D(_01619_),
    .Q_N(_11791_),
    .Q(\atari2600.ram[121][1] ));
 sg13g2_dfrbp_1 _28007_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1112),
    .D(_01620_),
    .Q_N(_11790_),
    .Q(\atari2600.ram[121][2] ));
 sg13g2_dfrbp_1 _28008_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1111),
    .D(_01621_),
    .Q_N(_11789_),
    .Q(\atari2600.ram[121][3] ));
 sg13g2_dfrbp_1 _28009_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1110),
    .D(_01622_),
    .Q_N(_11788_),
    .Q(\atari2600.ram[121][4] ));
 sg13g2_dfrbp_1 _28010_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1109),
    .D(_01623_),
    .Q_N(_11787_),
    .Q(\atari2600.ram[121][5] ));
 sg13g2_dfrbp_1 _28011_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1108),
    .D(_01624_),
    .Q_N(_11786_),
    .Q(\atari2600.ram[121][6] ));
 sg13g2_dfrbp_1 _28012_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1107),
    .D(_01625_),
    .Q_N(_11785_),
    .Q(\atari2600.ram[121][7] ));
 sg13g2_dfrbp_1 _28013_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1106),
    .D(_01626_),
    .Q_N(_11784_),
    .Q(\atari2600.ram[122][0] ));
 sg13g2_dfrbp_1 _28014_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1105),
    .D(_01627_),
    .Q_N(_11783_),
    .Q(\atari2600.ram[122][1] ));
 sg13g2_dfrbp_1 _28015_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1104),
    .D(_01628_),
    .Q_N(_11782_),
    .Q(\atari2600.ram[122][2] ));
 sg13g2_dfrbp_1 _28016_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1103),
    .D(_01629_),
    .Q_N(_11781_),
    .Q(\atari2600.ram[122][3] ));
 sg13g2_dfrbp_1 _28017_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1102),
    .D(_01630_),
    .Q_N(_11780_),
    .Q(\atari2600.ram[122][4] ));
 sg13g2_dfrbp_1 _28018_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1101),
    .D(_01631_),
    .Q_N(_11779_),
    .Q(\atari2600.ram[122][5] ));
 sg13g2_dfrbp_1 _28019_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1100),
    .D(_01632_),
    .Q_N(_11778_),
    .Q(\atari2600.ram[122][6] ));
 sg13g2_dfrbp_1 _28020_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1099),
    .D(_01633_),
    .Q_N(_11777_),
    .Q(\atari2600.ram[122][7] ));
 sg13g2_dfrbp_1 _28021_ (.CLK(clknet_leaf_362_clk),
    .RESET_B(net1098),
    .D(_01634_),
    .Q_N(_00092_),
    .Q(\atari2600.cpu.AXYS[3][0] ));
 sg13g2_dfrbp_1 _28022_ (.CLK(clknet_leaf_361_clk),
    .RESET_B(net1097),
    .D(_01635_),
    .Q_N(_00086_),
    .Q(\atari2600.cpu.AXYS[3][1] ));
 sg13g2_dfrbp_1 _28023_ (.CLK(clknet_leaf_359_clk),
    .RESET_B(net1096),
    .D(_01636_),
    .Q_N(_11776_),
    .Q(\atari2600.cpu.AXYS[3][2] ));
 sg13g2_dfrbp_1 _28024_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1095),
    .D(_01637_),
    .Q_N(_11775_),
    .Q(\atari2600.cpu.AXYS[3][3] ));
 sg13g2_dfrbp_1 _28025_ (.CLK(clknet_leaf_359_clk),
    .RESET_B(net1094),
    .D(_01638_),
    .Q_N(_11774_),
    .Q(\atari2600.cpu.AXYS[3][4] ));
 sg13g2_dfrbp_1 _28026_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1093),
    .D(_01639_),
    .Q_N(_11773_),
    .Q(\atari2600.cpu.AXYS[3][5] ));
 sg13g2_dfrbp_1 _28027_ (.CLK(clknet_leaf_360_clk),
    .RESET_B(net1092),
    .D(_01640_),
    .Q_N(_11772_),
    .Q(\atari2600.cpu.AXYS[3][6] ));
 sg13g2_dfrbp_1 _28028_ (.CLK(clknet_leaf_361_clk),
    .RESET_B(net1091),
    .D(_01641_),
    .Q_N(_11771_),
    .Q(\atari2600.cpu.AXYS[3][7] ));
 sg13g2_dfrbp_1 _28029_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1090),
    .D(_01642_),
    .Q_N(_11770_),
    .Q(\atari2600.ram[19][0] ));
 sg13g2_dfrbp_1 _28030_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1089),
    .D(_01643_),
    .Q_N(_11769_),
    .Q(\atari2600.ram[19][1] ));
 sg13g2_dfrbp_1 _28031_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1088),
    .D(_01644_),
    .Q_N(_11768_),
    .Q(\atari2600.ram[19][2] ));
 sg13g2_dfrbp_1 _28032_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1087),
    .D(_01645_),
    .Q_N(_11767_),
    .Q(\atari2600.ram[19][3] ));
 sg13g2_dfrbp_1 _28033_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1086),
    .D(_01646_),
    .Q_N(_11766_),
    .Q(\atari2600.ram[19][4] ));
 sg13g2_dfrbp_1 _28034_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1085),
    .D(_01647_),
    .Q_N(_11765_),
    .Q(\atari2600.ram[19][5] ));
 sg13g2_dfrbp_1 _28035_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1084),
    .D(_01648_),
    .Q_N(_11764_),
    .Q(\atari2600.ram[19][6] ));
 sg13g2_dfrbp_1 _28036_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1083),
    .D(_01649_),
    .Q_N(_11763_),
    .Q(\atari2600.ram[19][7] ));
 sg13g2_dfrbp_1 _28037_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1082),
    .D(_01650_),
    .Q_N(_11762_),
    .Q(\atari2600.ram[29][0] ));
 sg13g2_dfrbp_1 _28038_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1081),
    .D(_01651_),
    .Q_N(_11761_),
    .Q(\atari2600.ram[29][1] ));
 sg13g2_dfrbp_1 _28039_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1080),
    .D(_01652_),
    .Q_N(_11760_),
    .Q(\atari2600.ram[29][2] ));
 sg13g2_dfrbp_1 _28040_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1079),
    .D(_01653_),
    .Q_N(_11759_),
    .Q(\atari2600.ram[29][3] ));
 sg13g2_dfrbp_1 _28041_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1078),
    .D(_01654_),
    .Q_N(_11758_),
    .Q(\atari2600.ram[29][4] ));
 sg13g2_dfrbp_1 _28042_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1077),
    .D(_01655_),
    .Q_N(_11757_),
    .Q(\atari2600.ram[29][5] ));
 sg13g2_dfrbp_1 _28043_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1076),
    .D(_01656_),
    .Q_N(_11756_),
    .Q(\atari2600.ram[29][6] ));
 sg13g2_dfrbp_1 _28044_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1075),
    .D(_01657_),
    .Q_N(_11755_),
    .Q(\atari2600.ram[29][7] ));
 sg13g2_dfrbp_1 _28045_ (.CLK(clknet_leaf_358_clk),
    .RESET_B(net1074),
    .D(_01658_),
    .Q_N(_11754_),
    .Q(\atari2600.ram[39][0] ));
 sg13g2_dfrbp_1 _28046_ (.CLK(clknet_leaf_358_clk),
    .RESET_B(net1073),
    .D(_01659_),
    .Q_N(_11753_),
    .Q(\atari2600.ram[39][1] ));
 sg13g2_dfrbp_1 _28047_ (.CLK(clknet_leaf_358_clk),
    .RESET_B(net1072),
    .D(_01660_),
    .Q_N(_11752_),
    .Q(\atari2600.ram[39][2] ));
 sg13g2_dfrbp_1 _28048_ (.CLK(clknet_leaf_359_clk),
    .RESET_B(net1071),
    .D(_01661_),
    .Q_N(_11751_),
    .Q(\atari2600.ram[39][3] ));
 sg13g2_dfrbp_1 _28049_ (.CLK(clknet_leaf_351_clk),
    .RESET_B(net1070),
    .D(_01662_),
    .Q_N(_11750_),
    .Q(\atari2600.ram[39][4] ));
 sg13g2_dfrbp_1 _28050_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1069),
    .D(_01663_),
    .Q_N(_11749_),
    .Q(\atari2600.ram[39][5] ));
 sg13g2_dfrbp_1 _28051_ (.CLK(clknet_leaf_356_clk),
    .RESET_B(net1068),
    .D(_01664_),
    .Q_N(_11748_),
    .Q(\atari2600.ram[39][6] ));
 sg13g2_dfrbp_1 _28052_ (.CLK(clknet_leaf_357_clk),
    .RESET_B(net1067),
    .D(_01665_),
    .Q_N(_11747_),
    .Q(\atari2600.ram[39][7] ));
 sg13g2_dfrbp_1 _28053_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1066),
    .D(_01666_),
    .Q_N(_11746_),
    .Q(\atari2600.ram[49][0] ));
 sg13g2_dfrbp_1 _28054_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1065),
    .D(_01667_),
    .Q_N(_11745_),
    .Q(\atari2600.ram[49][1] ));
 sg13g2_dfrbp_1 _28055_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1064),
    .D(_01668_),
    .Q_N(_11744_),
    .Q(\atari2600.ram[49][2] ));
 sg13g2_dfrbp_1 _28056_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1063),
    .D(_01669_),
    .Q_N(_11743_),
    .Q(\atari2600.ram[49][3] ));
 sg13g2_dfrbp_1 _28057_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1062),
    .D(_01670_),
    .Q_N(_11742_),
    .Q(\atari2600.ram[49][4] ));
 sg13g2_dfrbp_1 _28058_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1061),
    .D(_01671_),
    .Q_N(_11741_),
    .Q(\atari2600.ram[49][5] ));
 sg13g2_dfrbp_1 _28059_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1060),
    .D(_01672_),
    .Q_N(_11740_),
    .Q(\atari2600.ram[49][6] ));
 sg13g2_dfrbp_1 _28060_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1059),
    .D(_01673_),
    .Q_N(_11739_),
    .Q(\atari2600.ram[49][7] ));
 sg13g2_dfrbp_1 _28061_ (.CLK(clknet_leaf_340_clk),
    .RESET_B(net1058),
    .D(_01674_),
    .Q_N(_11738_),
    .Q(\atari2600.ram[59][0] ));
 sg13g2_dfrbp_1 _28062_ (.CLK(clknet_leaf_354_clk),
    .RESET_B(net1057),
    .D(_01675_),
    .Q_N(_11737_),
    .Q(\atari2600.ram[59][1] ));
 sg13g2_dfrbp_1 _28063_ (.CLK(clknet_leaf_354_clk),
    .RESET_B(net1056),
    .D(_01676_),
    .Q_N(_11736_),
    .Q(\atari2600.ram[59][2] ));
 sg13g2_dfrbp_1 _28064_ (.CLK(clknet_leaf_341_clk),
    .RESET_B(net1055),
    .D(_01677_),
    .Q_N(_11735_),
    .Q(\atari2600.ram[59][3] ));
 sg13g2_dfrbp_1 _28065_ (.CLK(clknet_leaf_354_clk),
    .RESET_B(net1054),
    .D(_01678_),
    .Q_N(_11734_),
    .Q(\atari2600.ram[59][4] ));
 sg13g2_dfrbp_1 _28066_ (.CLK(clknet_leaf_340_clk),
    .RESET_B(net1053),
    .D(_01679_),
    .Q_N(_11733_),
    .Q(\atari2600.ram[59][5] ));
 sg13g2_dfrbp_1 _28067_ (.CLK(clknet_leaf_341_clk),
    .RESET_B(net1052),
    .D(_01680_),
    .Q_N(_11732_),
    .Q(\atari2600.ram[59][6] ));
 sg13g2_dfrbp_1 _28068_ (.CLK(clknet_leaf_341_clk),
    .RESET_B(net1051),
    .D(_01681_),
    .Q_N(_11731_),
    .Q(\atari2600.ram[59][7] ));
 sg13g2_dfrbp_1 _28069_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1050),
    .D(_01682_),
    .Q_N(_11730_),
    .Q(\atari2600.ram[69][0] ));
 sg13g2_dfrbp_1 _28070_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1049),
    .D(_01683_),
    .Q_N(_11729_),
    .Q(\atari2600.ram[69][1] ));
 sg13g2_dfrbp_1 _28071_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1048),
    .D(_01684_),
    .Q_N(_11728_),
    .Q(\atari2600.ram[69][2] ));
 sg13g2_dfrbp_1 _28072_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1047),
    .D(_01685_),
    .Q_N(_11727_),
    .Q(\atari2600.ram[69][3] ));
 sg13g2_dfrbp_1 _28073_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1046),
    .D(_01686_),
    .Q_N(_11726_),
    .Q(\atari2600.ram[69][4] ));
 sg13g2_dfrbp_1 _28074_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1045),
    .D(_01687_),
    .Q_N(_11725_),
    .Q(\atari2600.ram[69][5] ));
 sg13g2_dfrbp_1 _28075_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1044),
    .D(_01688_),
    .Q_N(_11724_),
    .Q(\atari2600.ram[69][6] ));
 sg13g2_dfrbp_1 _28076_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1043),
    .D(_01689_),
    .Q_N(_11723_),
    .Q(\atari2600.ram[69][7] ));
 sg13g2_dfrbp_1 _28077_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1042),
    .D(_01690_),
    .Q_N(_11722_),
    .Q(\atari2600.ram[79][0] ));
 sg13g2_dfrbp_1 _28078_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1041),
    .D(_01691_),
    .Q_N(_11721_),
    .Q(\atari2600.ram[79][1] ));
 sg13g2_dfrbp_1 _28079_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1040),
    .D(_01692_),
    .Q_N(_11720_),
    .Q(\atari2600.ram[79][2] ));
 sg13g2_dfrbp_1 _28080_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1039),
    .D(_01693_),
    .Q_N(_11719_),
    .Q(\atari2600.ram[79][3] ));
 sg13g2_dfrbp_1 _28081_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1038),
    .D(_01694_),
    .Q_N(_11718_),
    .Q(\atari2600.ram[79][4] ));
 sg13g2_dfrbp_1 _28082_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1037),
    .D(_01695_),
    .Q_N(_11717_),
    .Q(\atari2600.ram[79][5] ));
 sg13g2_dfrbp_1 _28083_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1036),
    .D(_01696_),
    .Q_N(_11716_),
    .Q(\atari2600.ram[79][6] ));
 sg13g2_dfrbp_1 _28084_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1035),
    .D(_01697_),
    .Q_N(_11715_),
    .Q(\atari2600.ram[79][7] ));
 sg13g2_dfrbp_1 _28085_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1034),
    .D(_01698_),
    .Q_N(_11714_),
    .Q(\atari2600.ram[89][0] ));
 sg13g2_dfrbp_1 _28086_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1033),
    .D(_01699_),
    .Q_N(_11713_),
    .Q(\atari2600.ram[89][1] ));
 sg13g2_dfrbp_1 _28087_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1032),
    .D(_01700_),
    .Q_N(_11712_),
    .Q(\atari2600.ram[89][2] ));
 sg13g2_dfrbp_1 _28088_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1031),
    .D(_01701_),
    .Q_N(_11711_),
    .Q(\atari2600.ram[89][3] ));
 sg13g2_dfrbp_1 _28089_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1030),
    .D(_01702_),
    .Q_N(_11710_),
    .Q(\atari2600.ram[89][4] ));
 sg13g2_dfrbp_1 _28090_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1029),
    .D(_01703_),
    .Q_N(_11709_),
    .Q(\atari2600.ram[89][5] ));
 sg13g2_dfrbp_1 _28091_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1028),
    .D(_01704_),
    .Q_N(_11708_),
    .Q(\atari2600.ram[89][6] ));
 sg13g2_dfrbp_1 _28092_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1027),
    .D(_01705_),
    .Q_N(_11707_),
    .Q(\atari2600.ram[89][7] ));
 sg13g2_dfrbp_1 _28093_ (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1026),
    .D(_01706_),
    .Q_N(_11706_),
    .Q(\atari2600.ram[99][0] ));
 sg13g2_dfrbp_1 _28094_ (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1025),
    .D(_01707_),
    .Q_N(_11705_),
    .Q(\atari2600.ram[99][1] ));
 sg13g2_dfrbp_1 _28095_ (.CLK(clknet_leaf_335_clk),
    .RESET_B(net1024),
    .D(_01708_),
    .Q_N(_11704_),
    .Q(\atari2600.ram[99][2] ));
 sg13g2_dfrbp_1 _28096_ (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1023),
    .D(_01709_),
    .Q_N(_11703_),
    .Q(\atari2600.ram[99][3] ));
 sg13g2_dfrbp_1 _28097_ (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1022),
    .D(_01710_),
    .Q_N(_11702_),
    .Q(\atari2600.ram[99][4] ));
 sg13g2_dfrbp_1 _28098_ (.CLK(clknet_leaf_339_clk),
    .RESET_B(net1021),
    .D(_01711_),
    .Q_N(_11701_),
    .Q(\atari2600.ram[99][5] ));
 sg13g2_dfrbp_1 _28099_ (.CLK(clknet_leaf_334_clk),
    .RESET_B(net1020),
    .D(_01712_),
    .Q_N(_11700_),
    .Q(\atari2600.ram[99][6] ));
 sg13g2_dfrbp_1 _28100_ (.CLK(clknet_leaf_333_clk),
    .RESET_B(net1019),
    .D(_01713_),
    .Q_N(_11699_),
    .Q(\atari2600.ram[99][7] ));
 sg13g2_dfrbp_1 _28101_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1018),
    .D(_01714_),
    .Q_N(_11698_),
    .Q(\atari2600.ram[109][0] ));
 sg13g2_dfrbp_1 _28102_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1017),
    .D(_01715_),
    .Q_N(_11697_),
    .Q(\atari2600.ram[109][1] ));
 sg13g2_dfrbp_1 _28103_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1016),
    .D(_01716_),
    .Q_N(_11696_),
    .Q(\atari2600.ram[109][2] ));
 sg13g2_dfrbp_1 _28104_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1015),
    .D(_01717_),
    .Q_N(_11695_),
    .Q(\atari2600.ram[109][3] ));
 sg13g2_dfrbp_1 _28105_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1014),
    .D(_01718_),
    .Q_N(_11694_),
    .Q(\atari2600.ram[109][4] ));
 sg13g2_dfrbp_1 _28106_ (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1013),
    .D(_01719_),
    .Q_N(_11693_),
    .Q(\atari2600.ram[109][5] ));
 sg13g2_dfrbp_1 _28107_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1012),
    .D(_01720_),
    .Q_N(_11692_),
    .Q(\atari2600.ram[109][6] ));
 sg13g2_dfrbp_1 _28108_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1011),
    .D(_01721_),
    .Q_N(_11691_),
    .Q(\atari2600.ram[109][7] ));
 sg13g2_dfrbp_1 _28109_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1010),
    .D(_01722_),
    .Q_N(_11690_),
    .Q(\atari2600.ram[119][0] ));
 sg13g2_dfrbp_1 _28110_ (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1009),
    .D(_01723_),
    .Q_N(_11689_),
    .Q(\atari2600.ram[119][1] ));
 sg13g2_dfrbp_1 _28111_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1008),
    .D(_01724_),
    .Q_N(_11688_),
    .Q(\atari2600.ram[119][2] ));
 sg13g2_dfrbp_1 _28112_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1007),
    .D(_01725_),
    .Q_N(_11687_),
    .Q(\atari2600.ram[119][3] ));
 sg13g2_dfrbp_1 _28113_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1006),
    .D(_01726_),
    .Q_N(_11686_),
    .Q(\atari2600.ram[119][4] ));
 sg13g2_dfrbp_1 _28114_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1005),
    .D(_01727_),
    .Q_N(_11685_),
    .Q(\atari2600.ram[119][5] ));
 sg13g2_dfrbp_1 _28115_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1004),
    .D(_01728_),
    .Q_N(_11684_),
    .Q(\atari2600.ram[119][6] ));
 sg13g2_dfrbp_1 _28116_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1003),
    .D(_01729_),
    .Q_N(_11683_),
    .Q(\atari2600.ram[119][7] ));
 sg13g2_dfrbp_1 _28117_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1002),
    .D(_01730_),
    .Q_N(_11682_),
    .Q(\atari2600.ram[74][0] ));
 sg13g2_dfrbp_1 _28118_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1001),
    .D(_01731_),
    .Q_N(_11681_),
    .Q(\atari2600.ram[74][1] ));
 sg13g2_dfrbp_1 _28119_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1000),
    .D(_01732_),
    .Q_N(_11680_),
    .Q(\atari2600.ram[74][2] ));
 sg13g2_dfrbp_1 _28120_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net999),
    .D(_01733_),
    .Q_N(_11679_),
    .Q(\atari2600.ram[74][3] ));
 sg13g2_dfrbp_1 _28121_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net998),
    .D(_01734_),
    .Q_N(_11678_),
    .Q(\atari2600.ram[74][4] ));
 sg13g2_dfrbp_1 _28122_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net997),
    .D(_01735_),
    .Q_N(_11677_),
    .Q(\atari2600.ram[74][5] ));
 sg13g2_dfrbp_1 _28123_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net996),
    .D(_01736_),
    .Q_N(_11676_),
    .Q(\atari2600.ram[74][6] ));
 sg13g2_dfrbp_1 _28124_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net995),
    .D(_01737_),
    .Q_N(_11675_),
    .Q(\atari2600.ram[74][7] ));
 sg13g2_dfrbp_1 _28125_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net994),
    .D(_01738_),
    .Q_N(_11674_),
    .Q(\atari2600.ram[85][0] ));
 sg13g2_dfrbp_1 _28126_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net993),
    .D(_01739_),
    .Q_N(_11673_),
    .Q(\atari2600.ram[85][1] ));
 sg13g2_dfrbp_1 _28127_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net992),
    .D(_01740_),
    .Q_N(_11672_),
    .Q(\atari2600.ram[85][2] ));
 sg13g2_dfrbp_1 _28128_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net991),
    .D(_01741_),
    .Q_N(_11671_),
    .Q(\atari2600.ram[85][3] ));
 sg13g2_dfrbp_1 _28129_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net990),
    .D(_01742_),
    .Q_N(_11670_),
    .Q(\atari2600.ram[85][4] ));
 sg13g2_dfrbp_1 _28130_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net989),
    .D(_01743_),
    .Q_N(_11669_),
    .Q(\atari2600.ram[85][5] ));
 sg13g2_dfrbp_1 _28131_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net988),
    .D(_01744_),
    .Q_N(_11668_),
    .Q(\atari2600.ram[85][6] ));
 sg13g2_dfrbp_1 _28132_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net987),
    .D(_01745_),
    .Q_N(_11667_),
    .Q(\atari2600.ram[85][7] ));
 sg13g2_dfrbp_1 _28133_ (.CLK(clknet_leaf_352_clk),
    .RESET_B(net986),
    .D(_01746_),
    .Q_N(_11666_),
    .Q(\atari2600.ram[34][0] ));
 sg13g2_dfrbp_1 _28134_ (.CLK(clknet_leaf_350_clk),
    .RESET_B(net985),
    .D(_01747_),
    .Q_N(_11665_),
    .Q(\atari2600.ram[34][1] ));
 sg13g2_dfrbp_1 _28135_ (.CLK(clknet_leaf_351_clk),
    .RESET_B(net984),
    .D(_01748_),
    .Q_N(_11664_),
    .Q(\atari2600.ram[34][2] ));
 sg13g2_dfrbp_1 _28136_ (.CLK(clknet_leaf_352_clk),
    .RESET_B(net983),
    .D(_01749_),
    .Q_N(_11663_),
    .Q(\atari2600.ram[34][3] ));
 sg13g2_dfrbp_1 _28137_ (.CLK(clknet_leaf_352_clk),
    .RESET_B(net982),
    .D(_01750_),
    .Q_N(_11662_),
    .Q(\atari2600.ram[34][4] ));
 sg13g2_dfrbp_1 _28138_ (.CLK(clknet_leaf_351_clk),
    .RESET_B(net981),
    .D(_01751_),
    .Q_N(_11661_),
    .Q(\atari2600.ram[34][5] ));
 sg13g2_dfrbp_1 _28139_ (.CLK(clknet_leaf_352_clk),
    .RESET_B(net980),
    .D(_01752_),
    .Q_N(_11660_),
    .Q(\atari2600.ram[34][6] ));
 sg13g2_dfrbp_1 _28140_ (.CLK(clknet_leaf_352_clk),
    .RESET_B(net979),
    .D(_01753_),
    .Q_N(_11659_),
    .Q(\atari2600.ram[34][7] ));
 sg13g2_dfrbp_1 _28141_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net978),
    .D(_01754_),
    .Q_N(_11658_),
    .Q(\atari2600.cpu.ALU.BI7 ));
 sg13g2_dfrbp_1 _28142_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net977),
    .D(_01755_),
    .Q_N(_11657_),
    .Q(\atari2600.pia.diag[0] ));
 sg13g2_dfrbp_1 _28143_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net975),
    .D(net7088),
    .Q_N(_11656_),
    .Q(\atari2600.pia.diag[1] ));
 sg13g2_dfrbp_1 _28144_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net973),
    .D(_01757_),
    .Q_N(_11655_),
    .Q(\atari2600.pia.diag[2] ));
 sg13g2_dfrbp_1 _28145_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net971),
    .D(_01758_),
    .Q_N(_11654_),
    .Q(\atari2600.pia.diag[3] ));
 sg13g2_dfrbp_1 _28146_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net969),
    .D(net3830),
    .Q_N(_11653_),
    .Q(\atari2600.pia.diag[4] ));
 sg13g2_dfrbp_1 _28147_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net967),
    .D(_01760_),
    .Q_N(_11652_),
    .Q(\atari2600.pia.diag[5] ));
 sg13g2_dfrbp_1 _28148_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net965),
    .D(net7061),
    .Q_N(_11651_),
    .Q(\atari2600.pia.diag[6] ));
 sg13g2_dfrbp_1 _28149_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net963),
    .D(net6952),
    .Q_N(_11650_),
    .Q(\atari2600.pia.diag[7] ));
 sg13g2_dfrbp_1 _28150_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net961),
    .D(_01763_),
    .Q_N(_11649_),
    .Q(\atari2600.pia.instat[1] ));
 sg13g2_dfrbp_1 _28151_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net959),
    .D(net4020),
    .Q_N(_11648_),
    .Q(\atari2600.pia.dat_o[0] ));
 sg13g2_dfrbp_1 _28152_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net958),
    .D(net3988),
    .Q_N(_11647_),
    .Q(\atari2600.pia.dat_o[1] ));
 sg13g2_dfrbp_1 _28153_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net957),
    .D(net3314),
    .Q_N(_11646_),
    .Q(\atari2600.pia.dat_o[2] ));
 sg13g2_dfrbp_1 _28154_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net956),
    .D(net6224),
    .Q_N(_11645_),
    .Q(\atari2600.pia.dat_o[3] ));
 sg13g2_dfrbp_1 _28155_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net955),
    .D(_01768_),
    .Q_N(_11644_),
    .Q(\atari2600.pia.dat_o[4] ));
 sg13g2_dfrbp_1 _28156_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net954),
    .D(_01769_),
    .Q_N(_11643_),
    .Q(\atari2600.pia.dat_o[5] ));
 sg13g2_dfrbp_1 _28157_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net953),
    .D(net3066),
    .Q_N(_11642_),
    .Q(\atari2600.pia.dat_o[6] ));
 sg13g2_dfrbp_1 _28158_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net952),
    .D(net3410),
    .Q_N(_11641_),
    .Q(\atari2600.pia.dat_o[7] ));
 sg13g2_dfrbp_1 _28159_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net951),
    .D(_01772_),
    .Q_N(_11640_),
    .Q(\atari2600.pia.time_counter[0] ));
 sg13g2_dfrbp_1 _28160_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net949),
    .D(_01773_),
    .Q_N(_11639_),
    .Q(\atari2600.pia.time_counter[1] ));
 sg13g2_dfrbp_1 _28161_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net947),
    .D(net6991),
    .Q_N(_11638_),
    .Q(\atari2600.pia.time_counter[2] ));
 sg13g2_dfrbp_1 _28162_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net945),
    .D(net7073),
    .Q_N(_11637_),
    .Q(\atari2600.pia.time_counter[3] ));
 sg13g2_dfrbp_1 _28163_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net943),
    .D(_01776_),
    .Q_N(_11636_),
    .Q(\atari2600.pia.time_counter[4] ));
 sg13g2_dfrbp_1 _28164_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net941),
    .D(_01777_),
    .Q_N(_11635_),
    .Q(\atari2600.pia.time_counter[5] ));
 sg13g2_dfrbp_1 _28165_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net939),
    .D(_01778_),
    .Q_N(_00078_),
    .Q(\atari2600.pia.time_counter[6] ));
 sg13g2_dfrbp_1 _28166_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net937),
    .D(_01779_),
    .Q_N(_11634_),
    .Q(\atari2600.pia.time_counter[7] ));
 sg13g2_dfrbp_1 _28167_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net935),
    .D(net6151),
    .Q_N(_11633_),
    .Q(\atari2600.pia.time_counter[8] ));
 sg13g2_dfrbp_1 _28168_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net933),
    .D(net3872),
    .Q_N(_11632_),
    .Q(\atari2600.pia.time_counter[9] ));
 sg13g2_dfrbp_1 _28169_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net931),
    .D(_01782_),
    .Q_N(_00079_),
    .Q(\atari2600.pia.time_counter[10] ));
 sg13g2_dfrbp_1 _28170_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net929),
    .D(net4024),
    .Q_N(_11631_),
    .Q(\atari2600.pia.time_counter[11] ));
 sg13g2_dfrbp_1 _28171_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net927),
    .D(_01784_),
    .Q_N(_11630_),
    .Q(\atari2600.pia.time_counter[12] ));
 sg13g2_dfrbp_1 _28172_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net925),
    .D(_01785_),
    .Q_N(_11629_),
    .Q(\atari2600.pia.time_counter[13] ));
 sg13g2_dfrbp_1 _28173_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net923),
    .D(net3796),
    .Q_N(_11628_),
    .Q(\atari2600.pia.time_counter[14] ));
 sg13g2_dfrbp_1 _28174_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net921),
    .D(_01787_),
    .Q_N(_11627_),
    .Q(\atari2600.pia.time_counter[15] ));
 sg13g2_dfrbp_1 _28175_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net919),
    .D(_01788_),
    .Q_N(_11626_),
    .Q(\atari2600.pia.time_counter[16] ));
 sg13g2_dfrbp_1 _28176_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net917),
    .D(_01789_),
    .Q_N(_11625_),
    .Q(\atari2600.pia.time_counter[17] ));
 sg13g2_dfrbp_1 _28177_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net915),
    .D(net3416),
    .Q_N(_11624_),
    .Q(\atari2600.pia.time_counter[18] ));
 sg13g2_dfrbp_1 _28178_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net913),
    .D(net6535),
    .Q_N(_11623_),
    .Q(\atari2600.pia.time_counter[19] ));
 sg13g2_dfrbp_1 _28179_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net911),
    .D(net3582),
    .Q_N(_11622_),
    .Q(\atari2600.pia.time_counter[20] ));
 sg13g2_dfrbp_1 _28180_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net909),
    .D(_01793_),
    .Q_N(_11621_),
    .Q(\atari2600.pia.time_counter[21] ));
 sg13g2_dfrbp_1 _28181_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net907),
    .D(_01794_),
    .Q_N(_11620_),
    .Q(\atari2600.pia.time_counter[22] ));
 sg13g2_dfrbp_1 _28182_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net905),
    .D(_01795_),
    .Q_N(_11619_),
    .Q(\atari2600.pia.time_counter[23] ));
 sg13g2_dfrbp_1 _28183_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net903),
    .D(net7332),
    .Q_N(_11618_),
    .Q(\atari2600.pia.underflow ));
 sg13g2_dfrbp_1 _28184_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net902),
    .D(_01797_),
    .Q_N(_11617_),
    .Q(\atari2600.pia.reset_timer[0] ));
 sg13g2_dfrbp_1 _28185_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net901),
    .D(_01798_),
    .Q_N(_11616_),
    .Q(\atari2600.pia.reset_timer[1] ));
 sg13g2_dfrbp_1 _28186_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net900),
    .D(_01799_),
    .Q_N(_11615_),
    .Q(\atari2600.pia.reset_timer[2] ));
 sg13g2_dfrbp_1 _28187_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net899),
    .D(_01800_),
    .Q_N(_11614_),
    .Q(\atari2600.pia.reset_timer[3] ));
 sg13g2_dfrbp_1 _28188_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net898),
    .D(_01801_),
    .Q_N(_11613_),
    .Q(\atari2600.pia.reset_timer[4] ));
 sg13g2_dfrbp_1 _28189_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net897),
    .D(_01802_),
    .Q_N(_11612_),
    .Q(\atari2600.pia.reset_timer[5] ));
 sg13g2_dfrbp_1 _28190_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net896),
    .D(_01803_),
    .Q_N(_11611_),
    .Q(\atari2600.pia.reset_timer[6] ));
 sg13g2_dfrbp_1 _28191_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net895),
    .D(_01804_),
    .Q_N(_11610_),
    .Q(\atari2600.pia.reset_timer[7] ));
 sg13g2_dfrbp_1 _28192_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net894),
    .D(_01805_),
    .Q_N(_11609_),
    .Q(\atari2600.pia.swa_dir[0] ));
 sg13g2_dfrbp_1 _28193_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net893),
    .D(_01806_),
    .Q_N(_11608_),
    .Q(\atari2600.pia.swa_dir[1] ));
 sg13g2_dfrbp_1 _28194_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net892),
    .D(_01807_),
    .Q_N(_11607_),
    .Q(\atari2600.pia.swa_dir[2] ));
 sg13g2_dfrbp_1 _28195_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net891),
    .D(_01808_),
    .Q_N(_11606_),
    .Q(\atari2600.pia.swa_dir[3] ));
 sg13g2_dfrbp_1 _28196_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net890),
    .D(_01809_),
    .Q_N(_11605_),
    .Q(\atari2600.pia.swa_dir[4] ));
 sg13g2_dfrbp_1 _28197_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net889),
    .D(_01810_),
    .Q_N(_11604_),
    .Q(\atari2600.pia.swa_dir[5] ));
 sg13g2_dfrbp_1 _28198_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net888),
    .D(_01811_),
    .Q_N(_11603_),
    .Q(\atari2600.pia.swa_dir[6] ));
 sg13g2_dfrbp_1 _28199_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net887),
    .D(_01812_),
    .Q_N(_11602_),
    .Q(\atari2600.pia.swa_dir[7] ));
 sg13g2_dfrbp_1 _28200_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net886),
    .D(_01813_),
    .Q_N(_11601_),
    .Q(\scanline[55][0] ));
 sg13g2_dfrbp_1 _28201_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net885),
    .D(_01814_),
    .Q_N(_11600_),
    .Q(\scanline[55][1] ));
 sg13g2_dfrbp_1 _28202_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net884),
    .D(_01815_),
    .Q_N(_11599_),
    .Q(\scanline[55][2] ));
 sg13g2_dfrbp_1 _28203_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net883),
    .D(_01816_),
    .Q_N(_11598_),
    .Q(\scanline[55][3] ));
 sg13g2_dfrbp_1 _28204_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net882),
    .D(_01817_),
    .Q_N(_11597_),
    .Q(\scanline[55][4] ));
 sg13g2_dfrbp_1 _28205_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net881),
    .D(_01818_),
    .Q_N(_11596_),
    .Q(\scanline[55][5] ));
 sg13g2_dfrbp_1 _28206_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net880),
    .D(_01819_),
    .Q_N(_11595_),
    .Q(\scanline[55][6] ));
 sg13g2_dfrbp_1 _28207_ (.CLK(clknet_leaf_333_clk),
    .RESET_B(net879),
    .D(net2948),
    .Q_N(_11594_),
    .Q(\atari2600.tia.old_grp1[0] ));
 sg13g2_dfrbp_1 _28208_ (.CLK(clknet_leaf_333_clk),
    .RESET_B(net878),
    .D(net2990),
    .Q_N(_11593_),
    .Q(\atari2600.tia.old_grp1[1] ));
 sg13g2_dfrbp_1 _28209_ (.CLK(clknet_leaf_334_clk),
    .RESET_B(net877),
    .D(net2941),
    .Q_N(_11592_),
    .Q(\atari2600.tia.old_grp1[2] ));
 sg13g2_dfrbp_1 _28210_ (.CLK(clknet_leaf_332_clk),
    .RESET_B(net876),
    .D(net3055),
    .Q_N(_11591_),
    .Q(\atari2600.tia.old_grp1[3] ));
 sg13g2_dfrbp_1 _28211_ (.CLK(clknet_leaf_331_clk),
    .RESET_B(net875),
    .D(net4318),
    .Q_N(_11590_),
    .Q(\atari2600.tia.old_grp1[4] ));
 sg13g2_dfrbp_1 _28212_ (.CLK(clknet_leaf_331_clk),
    .RESET_B(net874),
    .D(net6660),
    .Q_N(_11589_),
    .Q(\atari2600.tia.old_grp1[5] ));
 sg13g2_dfrbp_1 _28213_ (.CLK(clknet_leaf_330_clk),
    .RESET_B(net873),
    .D(net2965),
    .Q_N(_11588_),
    .Q(\atari2600.tia.old_grp1[6] ));
 sg13g2_dfrbp_1 _28214_ (.CLK(clknet_leaf_331_clk),
    .RESET_B(net872),
    .D(net2935),
    .Q_N(_11587_),
    .Q(\atari2600.tia.old_grp1[7] ));
 sg13g2_dfrbp_1 _28215_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net871),
    .D(_01828_),
    .Q_N(_11586_),
    .Q(\scanline[54][0] ));
 sg13g2_dfrbp_1 _28216_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net870),
    .D(_01829_),
    .Q_N(_11585_),
    .Q(\scanline[54][1] ));
 sg13g2_dfrbp_1 _28217_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net869),
    .D(_01830_),
    .Q_N(_11584_),
    .Q(\scanline[54][2] ));
 sg13g2_dfrbp_1 _28218_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net868),
    .D(_01831_),
    .Q_N(_11583_),
    .Q(\scanline[54][3] ));
 sg13g2_dfrbp_1 _28219_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net867),
    .D(_01832_),
    .Q_N(_11582_),
    .Q(\scanline[54][4] ));
 sg13g2_dfrbp_1 _28220_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net866),
    .D(_01833_),
    .Q_N(_11581_),
    .Q(\scanline[54][5] ));
 sg13g2_dfrbp_1 _28221_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net865),
    .D(_01834_),
    .Q_N(_11580_),
    .Q(\scanline[54][6] ));
 sg13g2_dfrbp_1 _28222_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net864),
    .D(_01835_),
    .Q_N(_11579_),
    .Q(\atari2600.tia.p0_spacing[4] ));
 sg13g2_dfrbp_1 _28223_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net862),
    .D(_01836_),
    .Q_N(_11578_),
    .Q(\atari2600.tia.p0_spacing[5] ));
 sg13g2_dfrbp_1 _28224_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net860),
    .D(_01837_),
    .Q_N(_11577_),
    .Q(\atari2600.tia.p0_spacing[6] ));
 sg13g2_dfrbp_1 _28225_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net858),
    .D(_01838_),
    .Q_N(_11576_),
    .Q(\atari2600.tia.p1_w[3] ));
 sg13g2_dfrbp_1 _28226_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net856),
    .D(_01839_),
    .Q_N(_11575_),
    .Q(\atari2600.tia.p1_w[4] ));
 sg13g2_dfrbp_1 _28227_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net854),
    .D(_01840_),
    .Q_N(_11574_),
    .Q(\atari2600.tia.p1_w[5] ));
 sg13g2_dfrbp_1 _28228_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net852),
    .D(_01841_),
    .Q_N(_11573_),
    .Q(\atari2600.tia.p1_scale[0] ));
 sg13g2_dfrbp_1 _28229_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net850),
    .D(_01842_),
    .Q_N(_11572_),
    .Q(\atari2600.tia.p1_scale[1] ));
 sg13g2_dfrbp_1 _28230_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net848),
    .D(_01843_),
    .Q_N(_11571_),
    .Q(\atari2600.tia.p0_scale[0] ));
 sg13g2_dfrbp_1 _28231_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net846),
    .D(_01844_),
    .Q_N(_11570_),
    .Q(\atari2600.tia.p0_scale[1] ));
 sg13g2_dfrbp_1 _28232_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net844),
    .D(_01845_),
    .Q_N(_11569_),
    .Q(\atari2600.tia.p0_w[3] ));
 sg13g2_dfrbp_1 _28233_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net842),
    .D(_01846_),
    .Q_N(_11568_),
    .Q(\atari2600.tia.p0_w[4] ));
 sg13g2_dfrbp_1 _28234_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net840),
    .D(_01847_),
    .Q_N(_11567_),
    .Q(\atari2600.tia.p0_w[5] ));
 sg13g2_dfrbp_1 _28235_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net838),
    .D(_01848_),
    .Q_N(_11566_),
    .Q(\atari2600.pia.interval[3] ));
 sg13g2_dfrbp_1 _28236_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net836),
    .D(_01849_),
    .Q_N(_11565_),
    .Q(\atari2600.pia.interval[6] ));
 sg13g2_dfrbp_1 _28237_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net834),
    .D(_01850_),
    .Q_N(_11564_),
    .Q(\atari2600.pia.interval[10] ));
 sg13g2_dfrbp_1 _28238_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net832),
    .D(_01851_),
    .Q_N(_11563_),
    .Q(\atari2600.tia.m1_w[0] ));
 sg13g2_dfrbp_1 _28239_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net830),
    .D(_01852_),
    .Q_N(_11562_),
    .Q(\atari2600.tia.m1_w[1] ));
 sg13g2_dfrbp_1 _28240_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net828),
    .D(_01853_),
    .Q_N(_11561_),
    .Q(\atari2600.tia.m1_w[2] ));
 sg13g2_dfrbp_1 _28241_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net826),
    .D(_01854_),
    .Q_N(_11560_),
    .Q(\atari2600.tia.m1_w[3] ));
 sg13g2_dfrbp_1 _28242_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net824),
    .D(_01855_),
    .Q_N(_11559_),
    .Q(\atari2600.tia.m0_w[0] ));
 sg13g2_dfrbp_1 _28243_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net822),
    .D(_01856_),
    .Q_N(_11558_),
    .Q(\atari2600.tia.m0_w[1] ));
 sg13g2_dfrbp_1 _28244_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net820),
    .D(_01857_),
    .Q_N(_11557_),
    .Q(\atari2600.tia.m0_w[2] ));
 sg13g2_dfrbp_1 _28245_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net818),
    .D(_01858_),
    .Q_N(_11556_),
    .Q(\atari2600.tia.m0_w[3] ));
 sg13g2_dfrbp_1 _28246_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net816),
    .D(_01859_),
    .Q_N(_11555_),
    .Q(\atari2600.tia.ball_w[0] ));
 sg13g2_dfrbp_1 _28247_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net814),
    .D(_01860_),
    .Q_N(_11554_),
    .Q(\atari2600.tia.ball_w[1] ));
 sg13g2_dfrbp_1 _28248_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net812),
    .D(_01861_),
    .Q_N(_11553_),
    .Q(\atari2600.tia.ball_w[2] ));
 sg13g2_dfrbp_1 _28249_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net810),
    .D(_01862_),
    .Q_N(_11552_),
    .Q(\atari2600.tia.ball_w[3] ));
 sg13g2_dfrbp_1 _28250_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net808),
    .D(_01863_),
    .Q_N(_11551_),
    .Q(\scanline[53][0] ));
 sg13g2_dfrbp_1 _28251_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net807),
    .D(_01864_),
    .Q_N(_11550_),
    .Q(\scanline[53][1] ));
 sg13g2_dfrbp_1 _28252_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net806),
    .D(_01865_),
    .Q_N(_11549_),
    .Q(\scanline[53][2] ));
 sg13g2_dfrbp_1 _28253_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net805),
    .D(_01866_),
    .Q_N(_11548_),
    .Q(\scanline[53][3] ));
 sg13g2_dfrbp_1 _28254_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net804),
    .D(_01867_),
    .Q_N(_11547_),
    .Q(\scanline[53][4] ));
 sg13g2_dfrbp_1 _28255_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net803),
    .D(_01868_),
    .Q_N(_11546_),
    .Q(\scanline[53][5] ));
 sg13g2_dfrbp_1 _28256_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net802),
    .D(_01869_),
    .Q_N(_11545_),
    .Q(\scanline[53][6] ));
 sg13g2_dfrbp_1 _28257_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net801),
    .D(_01870_),
    .Q_N(_11544_),
    .Q(\scanline[68][0] ));
 sg13g2_dfrbp_1 _28258_ (.CLK(clknet_leaf_285_clk),
    .RESET_B(net800),
    .D(_01871_),
    .Q_N(_11543_),
    .Q(\scanline[68][1] ));
 sg13g2_dfrbp_1 _28259_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net799),
    .D(_01872_),
    .Q_N(_11542_),
    .Q(\scanline[68][2] ));
 sg13g2_dfrbp_1 _28260_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net798),
    .D(_01873_),
    .Q_N(_11541_),
    .Q(\scanline[68][3] ));
 sg13g2_dfrbp_1 _28261_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net797),
    .D(_01874_),
    .Q_N(_11540_),
    .Q(\scanline[68][4] ));
 sg13g2_dfrbp_1 _28262_ (.CLK(clknet_leaf_287_clk),
    .RESET_B(net796),
    .D(_01875_),
    .Q_N(_11539_),
    .Q(\scanline[68][5] ));
 sg13g2_dfrbp_1 _28263_ (.CLK(clknet_leaf_275_clk),
    .RESET_B(net795),
    .D(_01876_),
    .Q_N(_11538_),
    .Q(\scanline[68][6] ));
 sg13g2_dfrbp_1 _28264_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net794),
    .D(_01877_),
    .Q_N(_11537_),
    .Q(\scanline[52][0] ));
 sg13g2_dfrbp_1 _28265_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net793),
    .D(_01878_),
    .Q_N(_11536_),
    .Q(\scanline[52][1] ));
 sg13g2_dfrbp_1 _28266_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net792),
    .D(_01879_),
    .Q_N(_11535_),
    .Q(\scanline[52][2] ));
 sg13g2_dfrbp_1 _28267_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net791),
    .D(_01880_),
    .Q_N(_11534_),
    .Q(\scanline[52][3] ));
 sg13g2_dfrbp_1 _28268_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net790),
    .D(_01881_),
    .Q_N(_11533_),
    .Q(\scanline[52][4] ));
 sg13g2_dfrbp_1 _28269_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net789),
    .D(_01882_),
    .Q_N(_11532_),
    .Q(\scanline[52][5] ));
 sg13g2_dfrbp_1 _28270_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net788),
    .D(_01883_),
    .Q_N(_11531_),
    .Q(\scanline[52][6] ));
 sg13g2_dfrbp_1 _28271_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net787),
    .D(_01884_),
    .Q_N(_11530_),
    .Q(\scanline[51][0] ));
 sg13g2_dfrbp_1 _28272_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net786),
    .D(_01885_),
    .Q_N(_11529_),
    .Q(\scanline[51][1] ));
 sg13g2_dfrbp_1 _28273_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net785),
    .D(_01886_),
    .Q_N(_11528_),
    .Q(\scanline[51][2] ));
 sg13g2_dfrbp_1 _28274_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net784),
    .D(_01887_),
    .Q_N(_11527_),
    .Q(\scanline[51][3] ));
 sg13g2_dfrbp_1 _28275_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net783),
    .D(_01888_),
    .Q_N(_11526_),
    .Q(\scanline[51][4] ));
 sg13g2_dfrbp_1 _28276_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net782),
    .D(_01889_),
    .Q_N(_11525_),
    .Q(\scanline[51][5] ));
 sg13g2_dfrbp_1 _28277_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net781),
    .D(_01890_),
    .Q_N(_11524_),
    .Q(\scanline[51][6] ));
 sg13g2_dfrbp_1 _28278_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net780),
    .D(_01891_),
    .Q_N(_11523_),
    .Q(\scanline[50][0] ));
 sg13g2_dfrbp_1 _28279_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net779),
    .D(_01892_),
    .Q_N(_11522_),
    .Q(\scanline[50][1] ));
 sg13g2_dfrbp_1 _28280_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net778),
    .D(_01893_),
    .Q_N(_11521_),
    .Q(\scanline[50][2] ));
 sg13g2_dfrbp_1 _28281_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net777),
    .D(_01894_),
    .Q_N(_11520_),
    .Q(\scanline[50][3] ));
 sg13g2_dfrbp_1 _28282_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net776),
    .D(_01895_),
    .Q_N(_11519_),
    .Q(\scanline[50][4] ));
 sg13g2_dfrbp_1 _28283_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net775),
    .D(_01896_),
    .Q_N(_11518_),
    .Q(\scanline[50][5] ));
 sg13g2_dfrbp_1 _28284_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net774),
    .D(_01897_),
    .Q_N(_11517_),
    .Q(\scanline[50][6] ));
 sg13g2_dfrbp_1 _28285_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net773),
    .D(_01898_),
    .Q_N(_11516_),
    .Q(\scanline[4][0] ));
 sg13g2_dfrbp_1 _28286_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net772),
    .D(_01899_),
    .Q_N(_11515_),
    .Q(\scanline[4][1] ));
 sg13g2_dfrbp_1 _28287_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net771),
    .D(_01900_),
    .Q_N(_11514_),
    .Q(\scanline[4][2] ));
 sg13g2_dfrbp_1 _28288_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net770),
    .D(_01901_),
    .Q_N(_11513_),
    .Q(\scanline[4][3] ));
 sg13g2_dfrbp_1 _28289_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net769),
    .D(_01902_),
    .Q_N(_11512_),
    .Q(\scanline[4][4] ));
 sg13g2_dfrbp_1 _28290_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net768),
    .D(_01903_),
    .Q_N(_11511_),
    .Q(\scanline[4][5] ));
 sg13g2_dfrbp_1 _28291_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net767),
    .D(_01904_),
    .Q_N(_11510_),
    .Q(\scanline[4][6] ));
 sg13g2_dfrbp_1 _28292_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net766),
    .D(_01905_),
    .Q_N(_11509_),
    .Q(\scanline[48][0] ));
 sg13g2_dfrbp_1 _28293_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net765),
    .D(_01906_),
    .Q_N(_11508_),
    .Q(\scanline[48][1] ));
 sg13g2_dfrbp_1 _28294_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net764),
    .D(_01907_),
    .Q_N(_11507_),
    .Q(\scanline[48][2] ));
 sg13g2_dfrbp_1 _28295_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net763),
    .D(_01908_),
    .Q_N(_11506_),
    .Q(\scanline[48][3] ));
 sg13g2_dfrbp_1 _28296_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net762),
    .D(_01909_),
    .Q_N(_11505_),
    .Q(\scanline[48][4] ));
 sg13g2_dfrbp_1 _28297_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net761),
    .D(_01910_),
    .Q_N(_11504_),
    .Q(\scanline[48][5] ));
 sg13g2_dfrbp_1 _28298_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net760),
    .D(_01911_),
    .Q_N(_11503_),
    .Q(\scanline[48][6] ));
 sg13g2_dfrbp_1 _28299_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net759),
    .D(_01912_),
    .Q_N(_11502_),
    .Q(\atari2600.ram[71][0] ));
 sg13g2_dfrbp_1 _28300_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net758),
    .D(_01913_),
    .Q_N(_11501_),
    .Q(\atari2600.ram[71][1] ));
 sg13g2_dfrbp_1 _28301_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net757),
    .D(_01914_),
    .Q_N(_11500_),
    .Q(\atari2600.ram[71][2] ));
 sg13g2_dfrbp_1 _28302_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net756),
    .D(_01915_),
    .Q_N(_11499_),
    .Q(\atari2600.ram[71][3] ));
 sg13g2_dfrbp_1 _28303_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net755),
    .D(_01916_),
    .Q_N(_11498_),
    .Q(\atari2600.ram[71][4] ));
 sg13g2_dfrbp_1 _28304_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net754),
    .D(_01917_),
    .Q_N(_11497_),
    .Q(\atari2600.ram[71][5] ));
 sg13g2_dfrbp_1 _28305_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net753),
    .D(_01918_),
    .Q_N(_11496_),
    .Q(\atari2600.ram[71][6] ));
 sg13g2_dfrbp_1 _28306_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net752),
    .D(_01919_),
    .Q_N(_11495_),
    .Q(\atari2600.ram[71][7] ));
 sg13g2_dfrbp_1 _28307_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net751),
    .D(net4166),
    .Q_N(_11494_),
    .Q(\flash_rom.addr[12] ));
 sg13g2_dfrbp_1 _28308_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net749),
    .D(net3022),
    .Q_N(_11493_),
    .Q(\flash_rom.addr[13] ));
 sg13g2_dfrbp_1 _28309_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net747),
    .D(_01922_),
    .Q_N(_11492_),
    .Q(\flash_rom.addr[14] ));
 sg13g2_dfrbp_1 _28310_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net745),
    .D(net3847),
    .Q_N(_11491_),
    .Q(\flash_rom.addr[15] ));
 sg13g2_dfrbp_1 _28311_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net743),
    .D(_01924_),
    .Q_N(_11490_),
    .Q(\flash_rom.addr[20] ));
 sg13g2_dfrbp_1 _28312_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net741),
    .D(_01925_),
    .Q_N(_11489_),
    .Q(\scanline[47][0] ));
 sg13g2_dfrbp_1 _28313_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net740),
    .D(_01926_),
    .Q_N(_11488_),
    .Q(\scanline[47][1] ));
 sg13g2_dfrbp_1 _28314_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net739),
    .D(_01927_),
    .Q_N(_11487_),
    .Q(\scanline[47][2] ));
 sg13g2_dfrbp_1 _28315_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net738),
    .D(_01928_),
    .Q_N(_11486_),
    .Q(\scanline[47][3] ));
 sg13g2_dfrbp_1 _28316_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net737),
    .D(_01929_),
    .Q_N(_11485_),
    .Q(\scanline[47][4] ));
 sg13g2_dfrbp_1 _28317_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net736),
    .D(_01930_),
    .Q_N(_11484_),
    .Q(\scanline[47][5] ));
 sg13g2_dfrbp_1 _28318_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net735),
    .D(_01931_),
    .Q_N(_11483_),
    .Q(\scanline[47][6] ));
 sg13g2_dfrbp_1 _28319_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net734),
    .D(_01932_),
    .Q_N(_11482_),
    .Q(\scanline[46][0] ));
 sg13g2_dfrbp_1 _28320_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net733),
    .D(_01933_),
    .Q_N(_11481_),
    .Q(\scanline[46][1] ));
 sg13g2_dfrbp_1 _28321_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net732),
    .D(_01934_),
    .Q_N(_11480_),
    .Q(\scanline[46][2] ));
 sg13g2_dfrbp_1 _28322_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net731),
    .D(_01935_),
    .Q_N(_11479_),
    .Q(\scanline[46][3] ));
 sg13g2_dfrbp_1 _28323_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net730),
    .D(_01936_),
    .Q_N(_11478_),
    .Q(\scanline[46][4] ));
 sg13g2_dfrbp_1 _28324_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net729),
    .D(_01937_),
    .Q_N(_11477_),
    .Q(\scanline[46][5] ));
 sg13g2_dfrbp_1 _28325_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net728),
    .D(_01938_),
    .Q_N(_11476_),
    .Q(\scanline[46][6] ));
 sg13g2_dfrbp_1 _28326_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net727),
    .D(_01939_),
    .Q_N(_11475_),
    .Q(\scanline[45][0] ));
 sg13g2_dfrbp_1 _28327_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net726),
    .D(_01940_),
    .Q_N(_11474_),
    .Q(\scanline[45][1] ));
 sg13g2_dfrbp_1 _28328_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net725),
    .D(_01941_),
    .Q_N(_11473_),
    .Q(\scanline[45][2] ));
 sg13g2_dfrbp_1 _28329_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net724),
    .D(_01942_),
    .Q_N(_11472_),
    .Q(\scanline[45][3] ));
 sg13g2_dfrbp_1 _28330_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net723),
    .D(_01943_),
    .Q_N(_11471_),
    .Q(\scanline[45][4] ));
 sg13g2_dfrbp_1 _28331_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net722),
    .D(_01944_),
    .Q_N(_11470_),
    .Q(\scanline[45][5] ));
 sg13g2_dfrbp_1 _28332_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net721),
    .D(_01945_),
    .Q_N(_11469_),
    .Q(\scanline[45][6] ));
 sg13g2_dfrbp_1 _28333_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net720),
    .D(_01946_),
    .Q_N(_11468_),
    .Q(\scanline[44][0] ));
 sg13g2_dfrbp_1 _28334_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net719),
    .D(_01947_),
    .Q_N(_11467_),
    .Q(\scanline[44][1] ));
 sg13g2_dfrbp_1 _28335_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net718),
    .D(_01948_),
    .Q_N(_11466_),
    .Q(\scanline[44][2] ));
 sg13g2_dfrbp_1 _28336_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net717),
    .D(_01949_),
    .Q_N(_11465_),
    .Q(\scanline[44][3] ));
 sg13g2_dfrbp_1 _28337_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net716),
    .D(_01950_),
    .Q_N(_11464_),
    .Q(\scanline[44][4] ));
 sg13g2_dfrbp_1 _28338_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net715),
    .D(_01951_),
    .Q_N(_11463_),
    .Q(\scanline[44][5] ));
 sg13g2_dfrbp_1 _28339_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net714),
    .D(_01952_),
    .Q_N(_11462_),
    .Q(\scanline[44][6] ));
 sg13g2_dfrbp_1 _28340_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net713),
    .D(_01953_),
    .Q_N(_11461_),
    .Q(\atari2600.ram[48][0] ));
 sg13g2_dfrbp_1 _28341_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net712),
    .D(_01954_),
    .Q_N(_11460_),
    .Q(\atari2600.ram[48][1] ));
 sg13g2_dfrbp_1 _28342_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net711),
    .D(_01955_),
    .Q_N(_11459_),
    .Q(\atari2600.ram[48][2] ));
 sg13g2_dfrbp_1 _28343_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net710),
    .D(_01956_),
    .Q_N(_11458_),
    .Q(\atari2600.ram[48][3] ));
 sg13g2_dfrbp_1 _28344_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net709),
    .D(_01957_),
    .Q_N(_11457_),
    .Q(\atari2600.ram[48][4] ));
 sg13g2_dfrbp_1 _28345_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net708),
    .D(_01958_),
    .Q_N(_11456_),
    .Q(\atari2600.ram[48][5] ));
 sg13g2_dfrbp_1 _28346_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net707),
    .D(_01959_),
    .Q_N(_11455_),
    .Q(\atari2600.ram[48][6] ));
 sg13g2_dfrbp_1 _28347_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net706),
    .D(_01960_),
    .Q_N(_11454_),
    .Q(\atari2600.ram[48][7] ));
 sg13g2_dfrbp_1 _28348_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net705),
    .D(_01961_),
    .Q_N(_11453_),
    .Q(\atari2600.ram[2][0] ));
 sg13g2_dfrbp_1 _28349_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net704),
    .D(_01962_),
    .Q_N(_11452_),
    .Q(\atari2600.ram[2][1] ));
 sg13g2_dfrbp_1 _28350_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net703),
    .D(_01963_),
    .Q_N(_11451_),
    .Q(\atari2600.ram[2][2] ));
 sg13g2_dfrbp_1 _28351_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net702),
    .D(_01964_),
    .Q_N(_11450_),
    .Q(\atari2600.ram[2][3] ));
 sg13g2_dfrbp_1 _28352_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net701),
    .D(_01965_),
    .Q_N(_11449_),
    .Q(\atari2600.ram[2][4] ));
 sg13g2_dfrbp_1 _28353_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net700),
    .D(_01966_),
    .Q_N(_11448_),
    .Q(\atari2600.ram[2][5] ));
 sg13g2_dfrbp_1 _28354_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net699),
    .D(_01967_),
    .Q_N(_11447_),
    .Q(\atari2600.ram[2][6] ));
 sg13g2_dfrbp_1 _28355_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net698),
    .D(_01968_),
    .Q_N(_11446_),
    .Q(\atari2600.ram[2][7] ));
 sg13g2_dfrbp_1 _28356_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net697),
    .D(_01969_),
    .Q_N(_11445_),
    .Q(\atari2600.ram[28][0] ));
 sg13g2_dfrbp_1 _28357_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net696),
    .D(_01970_),
    .Q_N(_11444_),
    .Q(\atari2600.ram[28][1] ));
 sg13g2_dfrbp_1 _28358_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net695),
    .D(_01971_),
    .Q_N(_11443_),
    .Q(\atari2600.ram[28][2] ));
 sg13g2_dfrbp_1 _28359_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net694),
    .D(_01972_),
    .Q_N(_11442_),
    .Q(\atari2600.ram[28][3] ));
 sg13g2_dfrbp_1 _28360_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net693),
    .D(_01973_),
    .Q_N(_11441_),
    .Q(\atari2600.ram[28][4] ));
 sg13g2_dfrbp_1 _28361_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net692),
    .D(_01974_),
    .Q_N(_11440_),
    .Q(\atari2600.ram[28][5] ));
 sg13g2_dfrbp_1 _28362_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net691),
    .D(_01975_),
    .Q_N(_11439_),
    .Q(\atari2600.ram[28][6] ));
 sg13g2_dfrbp_1 _28363_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net690),
    .D(_01976_),
    .Q_N(_11438_),
    .Q(\atari2600.ram[28][7] ));
 sg13g2_dfrbp_1 _28364_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net689),
    .D(_01977_),
    .Q_N(_11437_),
    .Q(\scanline[43][0] ));
 sg13g2_dfrbp_1 _28365_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net688),
    .D(_01978_),
    .Q_N(_11436_),
    .Q(\scanline[43][1] ));
 sg13g2_dfrbp_1 _28366_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net687),
    .D(_01979_),
    .Q_N(_11435_),
    .Q(\scanline[43][2] ));
 sg13g2_dfrbp_1 _28367_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net686),
    .D(_01980_),
    .Q_N(_11434_),
    .Q(\scanline[43][3] ));
 sg13g2_dfrbp_1 _28368_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net685),
    .D(_01981_),
    .Q_N(_11433_),
    .Q(\scanline[43][4] ));
 sg13g2_dfrbp_1 _28369_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net684),
    .D(_01982_),
    .Q_N(_11432_),
    .Q(\scanline[43][5] ));
 sg13g2_dfrbp_1 _28370_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net683),
    .D(_01983_),
    .Q_N(_11431_),
    .Q(\scanline[43][6] ));
 sg13g2_dfrbp_1 _28371_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net682),
    .D(_01984_),
    .Q_N(_11430_),
    .Q(\scanline[42][0] ));
 sg13g2_dfrbp_1 _28372_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net681),
    .D(_01985_),
    .Q_N(_11429_),
    .Q(\scanline[42][1] ));
 sg13g2_dfrbp_1 _28373_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net680),
    .D(_01986_),
    .Q_N(_11428_),
    .Q(\scanline[42][2] ));
 sg13g2_dfrbp_1 _28374_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net679),
    .D(_01987_),
    .Q_N(_11427_),
    .Q(\scanline[42][3] ));
 sg13g2_dfrbp_1 _28375_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net678),
    .D(_01988_),
    .Q_N(_11426_),
    .Q(\scanline[42][4] ));
 sg13g2_dfrbp_1 _28376_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net677),
    .D(_01989_),
    .Q_N(_11425_),
    .Q(\scanline[42][5] ));
 sg13g2_dfrbp_1 _28377_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net676),
    .D(_01990_),
    .Q_N(_11424_),
    .Q(\scanline[42][6] ));
 sg13g2_dfrbp_1 _28378_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net675),
    .D(_01991_),
    .Q_N(_11423_),
    .Q(\scanline[41][0] ));
 sg13g2_dfrbp_1 _28379_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net674),
    .D(_01992_),
    .Q_N(_11422_),
    .Q(\scanline[41][1] ));
 sg13g2_dfrbp_1 _28380_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net673),
    .D(_01993_),
    .Q_N(_11421_),
    .Q(\scanline[41][2] ));
 sg13g2_dfrbp_1 _28381_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net672),
    .D(_01994_),
    .Q_N(_11420_),
    .Q(\scanline[41][3] ));
 sg13g2_dfrbp_1 _28382_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net671),
    .D(_01995_),
    .Q_N(_11419_),
    .Q(\scanline[41][4] ));
 sg13g2_dfrbp_1 _28383_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net670),
    .D(_01996_),
    .Q_N(_11418_),
    .Q(\scanline[41][5] ));
 sg13g2_dfrbp_1 _28384_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net669),
    .D(_01997_),
    .Q_N(_11417_),
    .Q(\scanline[41][6] ));
 sg13g2_dfrbp_1 _28385_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net668),
    .D(_01998_),
    .Q_N(_11416_),
    .Q(\scanline[40][0] ));
 sg13g2_dfrbp_1 _28386_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net667),
    .D(_01999_),
    .Q_N(_11415_),
    .Q(\scanline[40][1] ));
 sg13g2_dfrbp_1 _28387_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net666),
    .D(_02000_),
    .Q_N(_11414_),
    .Q(\scanline[40][2] ));
 sg13g2_dfrbp_1 _28388_ (.CLK(clknet_leaf_273_clk),
    .RESET_B(net665),
    .D(_02001_),
    .Q_N(_11413_),
    .Q(\scanline[40][3] ));
 sg13g2_dfrbp_1 _28389_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net664),
    .D(_02002_),
    .Q_N(_11412_),
    .Q(\scanline[40][4] ));
 sg13g2_dfrbp_1 _28390_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net663),
    .D(_02003_),
    .Q_N(_11411_),
    .Q(\scanline[40][5] ));
 sg13g2_dfrbp_1 _28391_ (.CLK(clknet_leaf_274_clk),
    .RESET_B(net662),
    .D(_02004_),
    .Q_N(_11410_),
    .Q(\scanline[40][6] ));
 sg13g2_dfrbp_1 _28392_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net661),
    .D(_02005_),
    .Q_N(_11409_),
    .Q(\scanline[3][0] ));
 sg13g2_dfrbp_1 _28393_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net660),
    .D(_02006_),
    .Q_N(_11408_),
    .Q(\scanline[3][1] ));
 sg13g2_dfrbp_1 _28394_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net659),
    .D(_02007_),
    .Q_N(_11407_),
    .Q(\scanline[3][2] ));
 sg13g2_dfrbp_1 _28395_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net658),
    .D(_02008_),
    .Q_N(_11406_),
    .Q(\scanline[3][3] ));
 sg13g2_dfrbp_1 _28396_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net657),
    .D(_02009_),
    .Q_N(_11405_),
    .Q(\scanline[3][4] ));
 sg13g2_dfrbp_1 _28397_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net656),
    .D(_02010_),
    .Q_N(_11404_),
    .Q(\scanline[3][5] ));
 sg13g2_dfrbp_1 _28398_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net655),
    .D(_02011_),
    .Q_N(_11403_),
    .Q(\scanline[3][6] ));
 sg13g2_dfrbp_1 _28399_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net654),
    .D(net3466),
    .Q_N(_00106_),
    .Q(\atari2600.tia.audio_left_counter[0] ));
 sg13g2_dfrbp_1 _28400_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net652),
    .D(net7022),
    .Q_N(_11402_),
    .Q(\atari2600.tia.audio_left_counter[1] ));
 sg13g2_dfrbp_1 _28401_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net650),
    .D(net3934),
    .Q_N(_00108_),
    .Q(\atari2600.tia.audio_left_counter[2] ));
 sg13g2_dfrbp_1 _28402_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net648),
    .D(_02015_),
    .Q_N(_00109_),
    .Q(\atari2600.tia.audio_left_counter[3] ));
 sg13g2_dfrbp_1 _28403_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net646),
    .D(net3134),
    .Q_N(_00110_),
    .Q(\atari2600.tia.audio_left_counter[4] ));
 sg13g2_dfrbp_1 _28404_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net644),
    .D(_02017_),
    .Q_N(_00111_),
    .Q(\atari2600.tia.audio_left_counter[5] ));
 sg13g2_dfrbp_1 _28405_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net642),
    .D(net3993),
    .Q_N(_00113_),
    .Q(\atari2600.tia.audio_left_counter[6] ));
 sg13g2_dfrbp_1 _28406_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net640),
    .D(_02019_),
    .Q_N(_00114_),
    .Q(\atari2600.tia.audio_left_counter[7] ));
 sg13g2_dfrbp_1 _28407_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net638),
    .D(net3146),
    .Q_N(_00115_),
    .Q(\atari2600.tia.audio_left_counter[8] ));
 sg13g2_dfrbp_1 _28408_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net636),
    .D(_02021_),
    .Q_N(_00116_),
    .Q(\atari2600.tia.audio_left_counter[9] ));
 sg13g2_dfrbp_1 _28409_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net634),
    .D(net3806),
    .Q_N(_00117_),
    .Q(\atari2600.tia.audio_left_counter[10] ));
 sg13g2_dfrbp_1 _28410_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net632),
    .D(_02023_),
    .Q_N(_00118_),
    .Q(\atari2600.tia.audio_left_counter[11] ));
 sg13g2_dfrbp_1 _28411_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net630),
    .D(net3119),
    .Q_N(_00119_),
    .Q(\atari2600.tia.audio_left_counter[12] ));
 sg13g2_dfrbp_1 _28412_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net628),
    .D(_02025_),
    .Q_N(_00120_),
    .Q(\atari2600.tia.audio_left_counter[13] ));
 sg13g2_dfrbp_1 _28413_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net626),
    .D(net2975),
    .Q_N(_00121_),
    .Q(\atari2600.tia.audio_left_counter[14] ));
 sg13g2_dfrbp_1 _28414_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net624),
    .D(_02027_),
    .Q_N(_00122_),
    .Q(\atari2600.tia.audio_left_counter[15] ));
 sg13g2_dfrbp_1 _28415_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net622),
    .D(net2905),
    .Q_N(_00168_),
    .Q(\atari2600.tia.audio_right_counter[0] ));
 sg13g2_dfrbp_1 _28416_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net620),
    .D(net7245),
    .Q_N(_11401_),
    .Q(\atari2600.tia.audio_right_counter[1] ));
 sg13g2_dfrbp_1 _28417_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net618),
    .D(net6890),
    .Q_N(_00123_),
    .Q(\atari2600.tia.audio_right_counter[2] ));
 sg13g2_dfrbp_1 _28418_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net616),
    .D(net3839),
    .Q_N(_00124_),
    .Q(\atari2600.tia.audio_right_counter[3] ));
 sg13g2_dfrbp_1 _28419_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net614),
    .D(net6285),
    .Q_N(_00125_),
    .Q(\atari2600.tia.audio_right_counter[4] ));
 sg13g2_dfrbp_1 _28420_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net612),
    .D(net4136),
    .Q_N(_00126_),
    .Q(\atari2600.tia.audio_right_counter[5] ));
 sg13g2_dfrbp_1 _28421_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net610),
    .D(_02034_),
    .Q_N(_00127_),
    .Q(\atari2600.tia.audio_right_counter[6] ));
 sg13g2_dfrbp_1 _28422_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net608),
    .D(net3927),
    .Q_N(_00128_),
    .Q(\atari2600.tia.audio_right_counter[7] ));
 sg13g2_dfrbp_1 _28423_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net606),
    .D(net6792),
    .Q_N(_00129_),
    .Q(\atari2600.tia.audio_right_counter[8] ));
 sg13g2_dfrbp_1 _28424_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net604),
    .D(net3983),
    .Q_N(_00130_),
    .Q(\atari2600.tia.audio_right_counter[9] ));
 sg13g2_dfrbp_1 _28425_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net602),
    .D(net6204),
    .Q_N(_00131_),
    .Q(\atari2600.tia.audio_right_counter[10] ));
 sg13g2_dfrbp_1 _28426_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net600),
    .D(net3755),
    .Q_N(_00132_),
    .Q(\atari2600.tia.audio_right_counter[11] ));
 sg13g2_dfrbp_1 _28427_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net598),
    .D(_02040_),
    .Q_N(_00133_),
    .Q(\atari2600.tia.audio_right_counter[12] ));
 sg13g2_dfrbp_1 _28428_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net596),
    .D(net3857),
    .Q_N(_00134_),
    .Q(\atari2600.tia.audio_right_counter[13] ));
 sg13g2_dfrbp_1 _28429_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net594),
    .D(net4008),
    .Q_N(_00135_),
    .Q(\atari2600.tia.audio_right_counter[14] ));
 sg13g2_dfrbp_1 _28430_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net592),
    .D(_02043_),
    .Q_N(_00136_),
    .Q(\atari2600.tia.audio_right_counter[15] ));
 sg13g2_dfrbp_1 _28431_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net590),
    .D(_02044_),
    .Q_N(_00167_),
    .Q(\atari2600.tia.audio_l ));
 sg13g2_dfrbp_1 _28432_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net588),
    .D(net7307),
    .Q_N(_00166_),
    .Q(\atari2600.tia.audio_r ));
 sg13g2_dfrbp_1 _28433_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2154),
    .D(_02046_),
    .Q_N(_13239_),
    .Q(\atari2600.tia.vid_vsync ));
 sg13g2_dfrbp_1 _28434_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2155),
    .D(_00030_),
    .Q_N(_00165_),
    .Q(\atari2600.tia.vid_xpos[0] ));
 sg13g2_dfrbp_1 _28435_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2156),
    .D(_00031_),
    .Q_N(_00164_),
    .Q(\atari2600.tia.vid_xpos[1] ));
 sg13g2_dfrbp_1 _28436_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2157),
    .D(_00032_),
    .Q_N(_00151_),
    .Q(\atari2600.tia.vid_xpos[2] ));
 sg13g2_dfrbp_1 _28437_ (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2158),
    .D(_00033_),
    .Q_N(_00152_),
    .Q(\atari2600.tia.vid_xpos[3] ));
 sg13g2_dfrbp_1 _28438_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net2159),
    .D(_00034_),
    .Q_N(_00156_),
    .Q(\atari2600.tia.vid_xpos[4] ));
 sg13g2_dfrbp_1 _28439_ (.CLK(clknet_leaf_304_clk),
    .RESET_B(net2160),
    .D(_00035_),
    .Q_N(_00153_),
    .Q(\atari2600.tia.vid_xpos[5] ));
 sg13g2_dfrbp_1 _28440_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net2161),
    .D(_00036_),
    .Q_N(_00154_),
    .Q(\atari2600.tia.vid_xpos[6] ));
 sg13g2_dfrbp_1 _28441_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net2162),
    .D(_00037_),
    .Q_N(_00150_),
    .Q(\atari2600.tia.vid_xpos[7] ));
 sg13g2_dfrbp_1 _28442_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2163),
    .D(_00038_),
    .Q_N(_00048_),
    .Q(\atari2600.tia.vid_ypos[0] ));
 sg13g2_dfrbp_1 _28443_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2164),
    .D(_00039_),
    .Q_N(_00049_),
    .Q(\atari2600.tia.vid_ypos[1] ));
 sg13g2_dfrbp_1 _28444_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2165),
    .D(_00040_),
    .Q_N(_00050_),
    .Q(\atari2600.tia.vid_ypos[2] ));
 sg13g2_dfrbp_1 _28445_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2166),
    .D(_00041_),
    .Q_N(_00144_),
    .Q(\atari2600.tia.vid_ypos[3] ));
 sg13g2_dfrbp_1 _28446_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net2167),
    .D(net6757),
    .Q_N(_00051_),
    .Q(\atari2600.tia.vid_ypos[4] ));
 sg13g2_dfrbp_1 _28447_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2168),
    .D(net3680),
    .Q_N(_00077_),
    .Q(\atari2600.tia.vid_ypos[5] ));
 sg13g2_dfrbp_1 _28448_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2169),
    .D(net6883),
    .Q_N(_00052_),
    .Q(\atari2600.tia.vid_ypos[6] ));
 sg13g2_dfrbp_1 _28449_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2184),
    .D(net2931),
    .Q_N(_00053_),
    .Q(\atari2600.tia.vid_ypos[7] ));
 sg13g2_dfrbp_1 _28450_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net586),
    .D(_00046_),
    .Q_N(_00143_),
    .Q(\atari2600.tia.vid_ypos[8] ));
 sg13g2_dfrbp_1 _28451_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net584),
    .D(_02047_),
    .Q_N(_11400_),
    .Q(\atari2600.tia.vblank ));
 sg13g2_dfrbp_1 _28452_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net582),
    .D(_02048_),
    .Q_N(_11399_),
    .Q(\atari2600.stall_cpu ));
 sg13g2_dfrbp_1 _28453_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net580),
    .D(_02049_),
    .Q_N(_11398_),
    .Q(\atari2600.pia.swb_dir[2] ));
 sg13g2_dfrbp_1 _28454_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net579),
    .D(_02050_),
    .Q_N(_11397_),
    .Q(\atari2600.pia.swb_dir[4] ));
 sg13g2_dfrbp_1 _28455_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net578),
    .D(_02051_),
    .Q_N(_11396_),
    .Q(\atari2600.pia.swb_dir[5] ));
 sg13g2_dfrbp_1 _28456_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net577),
    .D(_02052_),
    .Q_N(_11395_),
    .Q(\atari2600.tia.colubk[0] ));
 sg13g2_dfrbp_1 _28457_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net575),
    .D(_02053_),
    .Q_N(_11394_),
    .Q(\atari2600.tia.colubk[1] ));
 sg13g2_dfrbp_1 _28458_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net573),
    .D(_02054_),
    .Q_N(_11393_),
    .Q(\atari2600.tia.colubk[2] ));
 sg13g2_dfrbp_1 _28459_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net571),
    .D(_02055_),
    .Q_N(_11392_),
    .Q(\atari2600.tia.colubk[3] ));
 sg13g2_dfrbp_1 _28460_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net569),
    .D(_02056_),
    .Q_N(_11391_),
    .Q(\atari2600.tia.colubk[4] ));
 sg13g2_dfrbp_1 _28461_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net567),
    .D(_02057_),
    .Q_N(_11390_),
    .Q(\atari2600.tia.colubk[5] ));
 sg13g2_dfrbp_1 _28462_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net565),
    .D(_02058_),
    .Q_N(_11389_),
    .Q(\atari2600.tia.colubk[6] ));
 sg13g2_dfrbp_1 _28463_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net563),
    .D(_02059_),
    .Q_N(_11388_),
    .Q(\atari2600.tia.colup0[0] ));
 sg13g2_dfrbp_1 _28464_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net561),
    .D(_02060_),
    .Q_N(_11387_),
    .Q(\atari2600.tia.colup0[1] ));
 sg13g2_dfrbp_1 _28465_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net559),
    .D(_02061_),
    .Q_N(_11386_),
    .Q(\atari2600.tia.colup0[2] ));
 sg13g2_dfrbp_1 _28466_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net557),
    .D(_02062_),
    .Q_N(_11385_),
    .Q(\atari2600.tia.colup0[3] ));
 sg13g2_dfrbp_1 _28467_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net555),
    .D(_02063_),
    .Q_N(_11384_),
    .Q(\atari2600.tia.colup0[4] ));
 sg13g2_dfrbp_1 _28468_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net553),
    .D(_02064_),
    .Q_N(_11383_),
    .Q(\atari2600.tia.colup0[5] ));
 sg13g2_dfrbp_1 _28469_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net551),
    .D(_02065_),
    .Q_N(_11382_),
    .Q(\atari2600.tia.colup0[6] ));
 sg13g2_dfrbp_1 _28470_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net549),
    .D(_02066_),
    .Q_N(_11381_),
    .Q(\atari2600.tia.colup1[0] ));
 sg13g2_dfrbp_1 _28471_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net547),
    .D(_02067_),
    .Q_N(_11380_),
    .Q(\atari2600.tia.colup1[1] ));
 sg13g2_dfrbp_1 _28472_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net545),
    .D(_02068_),
    .Q_N(_11379_),
    .Q(\atari2600.tia.colup1[2] ));
 sg13g2_dfrbp_1 _28473_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net543),
    .D(_02069_),
    .Q_N(_11378_),
    .Q(\atari2600.tia.colup1[3] ));
 sg13g2_dfrbp_1 _28474_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net541),
    .D(_02070_),
    .Q_N(_11377_),
    .Q(\atari2600.tia.colup1[4] ));
 sg13g2_dfrbp_1 _28475_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net539),
    .D(_02071_),
    .Q_N(_11376_),
    .Q(\atari2600.tia.colup1[5] ));
 sg13g2_dfrbp_1 _28476_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net537),
    .D(_02072_),
    .Q_N(_11375_),
    .Q(\atari2600.tia.colup1[6] ));
 sg13g2_dfrbp_1 _28477_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net535),
    .D(_02073_),
    .Q_N(_11374_),
    .Q(\atari2600.tia.colupf[0] ));
 sg13g2_dfrbp_1 _28478_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net533),
    .D(_02074_),
    .Q_N(_11373_),
    .Q(\atari2600.tia.colupf[1] ));
 sg13g2_dfrbp_1 _28479_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net531),
    .D(_02075_),
    .Q_N(_11372_),
    .Q(\atari2600.tia.colupf[2] ));
 sg13g2_dfrbp_1 _28480_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net529),
    .D(_02076_),
    .Q_N(_11371_),
    .Q(\atari2600.tia.colupf[3] ));
 sg13g2_dfrbp_1 _28481_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net527),
    .D(_02077_),
    .Q_N(_11370_),
    .Q(\atari2600.tia.colupf[4] ));
 sg13g2_dfrbp_1 _28482_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net525),
    .D(_02078_),
    .Q_N(_11369_),
    .Q(\atari2600.tia.colupf[5] ));
 sg13g2_dfrbp_1 _28483_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net523),
    .D(_02079_),
    .Q_N(_11368_),
    .Q(\atari2600.tia.colupf[6] ));
 sg13g2_dfrbp_1 _28484_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net521),
    .D(_02080_),
    .Q_N(_11367_),
    .Q(\atari2600.tia.enam0 ));
 sg13g2_dfrbp_1 _28485_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net519),
    .D(_02081_),
    .Q_N(_11366_),
    .Q(\atari2600.tia.enam1 ));
 sg13g2_dfrbp_1 _28486_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net517),
    .D(_02082_),
    .Q_N(_11365_),
    .Q(\atari2600.tia.enabl ));
 sg13g2_dfrbp_1 _28487_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net515),
    .D(_02083_),
    .Q_N(_11364_),
    .Q(\scanline[38][0] ));
 sg13g2_dfrbp_1 _28488_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net514),
    .D(_02084_),
    .Q_N(_11363_),
    .Q(\scanline[38][1] ));
 sg13g2_dfrbp_1 _28489_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net513),
    .D(_02085_),
    .Q_N(_11362_),
    .Q(\scanline[38][2] ));
 sg13g2_dfrbp_1 _28490_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net512),
    .D(_02086_),
    .Q_N(_11361_),
    .Q(\scanline[38][3] ));
 sg13g2_dfrbp_1 _28491_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net511),
    .D(_02087_),
    .Q_N(_11360_),
    .Q(\scanline[38][4] ));
 sg13g2_dfrbp_1 _28492_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net510),
    .D(_02088_),
    .Q_N(_11359_),
    .Q(\scanline[38][5] ));
 sg13g2_dfrbp_1 _28493_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net509),
    .D(_02089_),
    .Q_N(_11358_),
    .Q(\scanline[38][6] ));
 sg13g2_dfrbp_1 _28494_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net508),
    .D(_02090_),
    .Q_N(_11357_),
    .Q(\atari2600.tia.vdelp0 ));
 sg13g2_dfrbp_1 _28495_ (.CLK(clknet_leaf_331_clk),
    .RESET_B(net506),
    .D(_02091_),
    .Q_N(_11356_),
    .Q(\atari2600.tia.vdelp1 ));
 sg13g2_dfrbp_1 _28496_ (.CLK(clknet_leaf_326_clk),
    .RESET_B(net504),
    .D(_02092_),
    .Q_N(_00163_),
    .Q(\atari2600.tia.refp0 ));
 sg13g2_dfrbp_1 _28497_ (.CLK(clknet_leaf_328_clk),
    .RESET_B(net502),
    .D(_02093_),
    .Q_N(_00159_),
    .Q(\atari2600.tia.refp1 ));
 sg13g2_dfrbp_1 _28498_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net500),
    .D(_02094_),
    .Q_N(_11355_),
    .Q(\atari2600.tia.refpf ));
 sg13g2_dfrbp_1 _28499_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net498),
    .D(_02095_),
    .Q_N(_11354_),
    .Q(\atari2600.tia.scorepf ));
 sg13g2_dfrbp_1 _28500_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net496),
    .D(_02096_),
    .Q_N(_11353_),
    .Q(\atari2600.tia.pf_priority ));
 sg13g2_dfrbp_1 _28501_ (.CLK(clknet_leaf_327_clk),
    .RESET_B(net494),
    .D(_02097_),
    .Q_N(_11352_),
    .Q(\atari2600.tia.diag[104] ));
 sg13g2_dfrbp_1 _28502_ (.CLK(clknet_leaf_327_clk),
    .RESET_B(net492),
    .D(_02098_),
    .Q_N(_11351_),
    .Q(\atari2600.tia.diag[105] ));
 sg13g2_dfrbp_1 _28503_ (.CLK(clknet_leaf_329_clk),
    .RESET_B(net490),
    .D(_02099_),
    .Q_N(_11350_),
    .Q(\atari2600.tia.diag[106] ));
 sg13g2_dfrbp_1 _28504_ (.CLK(clknet_leaf_327_clk),
    .RESET_B(net488),
    .D(_02100_),
    .Q_N(_11349_),
    .Q(\atari2600.tia.diag[107] ));
 sg13g2_dfrbp_1 _28505_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net486),
    .D(_02101_),
    .Q_N(_11348_),
    .Q(\atari2600.tia.diag[108] ));
 sg13g2_dfrbp_1 _28506_ (.CLK(clknet_leaf_326_clk),
    .RESET_B(net484),
    .D(_02102_),
    .Q_N(_11347_),
    .Q(\atari2600.tia.diag[109] ));
 sg13g2_dfrbp_1 _28507_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net482),
    .D(_02103_),
    .Q_N(_11346_),
    .Q(\atari2600.tia.diag[110] ));
 sg13g2_dfrbp_1 _28508_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net480),
    .D(_02104_),
    .Q_N(_11345_),
    .Q(\atari2600.tia.diag[111] ));
 sg13g2_dfrbp_1 _28509_ (.CLK(clknet_leaf_333_clk),
    .RESET_B(net478),
    .D(_02105_),
    .Q_N(_11344_),
    .Q(\atari2600.tia.diag[96] ));
 sg13g2_dfrbp_1 _28510_ (.CLK(clknet_leaf_333_clk),
    .RESET_B(net476),
    .D(_02106_),
    .Q_N(_11343_),
    .Q(\atari2600.tia.diag[97] ));
 sg13g2_dfrbp_1 _28511_ (.CLK(clknet_leaf_334_clk),
    .RESET_B(net474),
    .D(_02107_),
    .Q_N(_11342_),
    .Q(\atari2600.tia.diag[98] ));
 sg13g2_dfrbp_1 _28512_ (.CLK(clknet_leaf_332_clk),
    .RESET_B(net472),
    .D(_02108_),
    .Q_N(_11341_),
    .Q(\atari2600.tia.diag[99] ));
 sg13g2_dfrbp_1 _28513_ (.CLK(clknet_leaf_328_clk),
    .RESET_B(net470),
    .D(_02109_),
    .Q_N(_11340_),
    .Q(\atari2600.tia.diag[100] ));
 sg13g2_dfrbp_1 _28514_ (.CLK(clknet_leaf_328_clk),
    .RESET_B(net468),
    .D(_02110_),
    .Q_N(_11339_),
    .Q(\atari2600.tia.diag[101] ));
 sg13g2_dfrbp_1 _28515_ (.CLK(clknet_leaf_331_clk),
    .RESET_B(net466),
    .D(_02111_),
    .Q_N(_11338_),
    .Q(\atari2600.tia.diag[102] ));
 sg13g2_dfrbp_1 _28516_ (.CLK(clknet_leaf_332_clk),
    .RESET_B(net464),
    .D(_02112_),
    .Q_N(_11337_),
    .Q(\atari2600.tia.diag[103] ));
 sg13g2_dfrbp_1 _28517_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net462),
    .D(_02113_),
    .Q_N(_11336_),
    .Q(\atari2600.tia.vid_out[0] ));
 sg13g2_dfrbp_1 _28518_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net461),
    .D(_02114_),
    .Q_N(_11335_),
    .Q(\atari2600.tia.vid_out[1] ));
 sg13g2_dfrbp_1 _28519_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net460),
    .D(_02115_),
    .Q_N(_11334_),
    .Q(\atari2600.tia.vid_out[2] ));
 sg13g2_dfrbp_1 _28520_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net459),
    .D(_02116_),
    .Q_N(_11333_),
    .Q(\atari2600.tia.vid_out[3] ));
 sg13g2_dfrbp_1 _28521_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net458),
    .D(_02117_),
    .Q_N(_11332_),
    .Q(\atari2600.tia.vid_out[4] ));
 sg13g2_dfrbp_1 _28522_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net457),
    .D(_02118_),
    .Q_N(_11331_),
    .Q(\atari2600.tia.vid_out[5] ));
 sg13g2_dfrbp_1 _28523_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net456),
    .D(_02119_),
    .Q_N(_11330_),
    .Q(\atari2600.tia.vid_out[6] ));
 sg13g2_dfrbp_1 _28524_ (.CLK(clknet_leaf_327_clk),
    .RESET_B(net455),
    .D(net3462),
    .Q_N(_11329_),
    .Q(\atari2600.tia.old_grp0[0] ));
 sg13g2_dfrbp_1 _28525_ (.CLK(clknet_leaf_325_clk),
    .RESET_B(net454),
    .D(net3370),
    .Q_N(_11328_),
    .Q(\atari2600.tia.old_grp0[1] ));
 sg13g2_dfrbp_1 _28526_ (.CLK(clknet_leaf_327_clk),
    .RESET_B(net453),
    .D(net3628),
    .Q_N(_11327_),
    .Q(\atari2600.tia.old_grp0[2] ));
 sg13g2_dfrbp_1 _28527_ (.CLK(clknet_leaf_327_clk),
    .RESET_B(net452),
    .D(net3202),
    .Q_N(_11326_),
    .Q(\atari2600.tia.old_grp0[3] ));
 sg13g2_dfrbp_1 _28528_ (.CLK(clknet_leaf_326_clk),
    .RESET_B(net451),
    .D(net3365),
    .Q_N(_11325_),
    .Q(\atari2600.tia.old_grp0[4] ));
 sg13g2_dfrbp_1 _28529_ (.CLK(clknet_leaf_326_clk),
    .RESET_B(net450),
    .D(net3219),
    .Q_N(_11324_),
    .Q(\atari2600.tia.old_grp0[5] ));
 sg13g2_dfrbp_1 _28530_ (.CLK(clknet_leaf_326_clk),
    .RESET_B(net449),
    .D(net3240),
    .Q_N(_11323_),
    .Q(\atari2600.tia.old_grp0[6] ));
 sg13g2_dfrbp_1 _28531_ (.CLK(clknet_leaf_326_clk),
    .RESET_B(net448),
    .D(net3272),
    .Q_N(_11322_),
    .Q(\atari2600.tia.old_grp0[7] ));
 sg13g2_dfrbp_1 _28532_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net447),
    .D(net7286),
    .Q_N(_11321_),
    .Q(\atari2600.tia.diag[64] ));
 sg13g2_dfrbp_1 _28533_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net445),
    .D(net7297),
    .Q_N(_11320_),
    .Q(\atari2600.tia.diag[65] ));
 sg13g2_dfrbp_1 _28534_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net443),
    .D(_02130_),
    .Q_N(_11319_),
    .Q(\atari2600.tia.diag[66] ));
 sg13g2_dfrbp_1 _28535_ (.CLK(clknet_leaf_326_clk),
    .RESET_B(net441),
    .D(_02131_),
    .Q_N(_11318_),
    .Q(\atari2600.tia.diag[67] ));
 sg13g2_dfrbp_1 _28536_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net439),
    .D(_02132_),
    .Q_N(_11317_),
    .Q(\atari2600.tia.diag[68] ));
 sg13g2_dfrbp_1 _28537_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net437),
    .D(_02133_),
    .Q_N(_00161_),
    .Q(\atari2600.tia.diag[69] ));
 sg13g2_dfrbp_1 _28538_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net435),
    .D(_02134_),
    .Q_N(_00160_),
    .Q(\atari2600.tia.diag[70] ));
 sg13g2_dfrbp_1 _28539_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net433),
    .D(_02135_),
    .Q_N(_00162_),
    .Q(\atari2600.tia.diag[71] ));
 sg13g2_dfrbp_1 _28540_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net431),
    .D(net7248),
    .Q_N(_11316_),
    .Q(\atari2600.tia.diag[56] ));
 sg13g2_dfrbp_1 _28541_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net429),
    .D(net7290),
    .Q_N(_11315_),
    .Q(\atari2600.tia.diag[57] ));
 sg13g2_dfrbp_1 _28542_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net427),
    .D(_02138_),
    .Q_N(_11314_),
    .Q(\atari2600.tia.diag[58] ));
 sg13g2_dfrbp_1 _28543_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net425),
    .D(_02139_),
    .Q_N(_11313_),
    .Q(\atari2600.tia.diag[59] ));
 sg13g2_dfrbp_1 _28544_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net423),
    .D(_02140_),
    .Q_N(_11312_),
    .Q(\atari2600.tia.diag[60] ));
 sg13g2_dfrbp_1 _28545_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net421),
    .D(_02141_),
    .Q_N(_00157_),
    .Q(\atari2600.tia.diag[61] ));
 sg13g2_dfrbp_1 _28546_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net419),
    .D(_02142_),
    .Q_N(_00155_),
    .Q(\atari2600.tia.diag[62] ));
 sg13g2_dfrbp_1 _28547_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net417),
    .D(_02143_),
    .Q_N(_00158_),
    .Q(\atari2600.tia.diag[63] ));
 sg13g2_dfrbp_1 _28548_ (.CLK(clknet_leaf_331_clk),
    .RESET_B(net415),
    .D(_02144_),
    .Q_N(_11311_),
    .Q(\atari2600.tia.diag[48] ));
 sg13g2_dfrbp_1 _28549_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net413),
    .D(_02145_),
    .Q_N(_11310_),
    .Q(\atari2600.tia.diag[49] ));
 sg13g2_dfrbp_1 _28550_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net411),
    .D(_02146_),
    .Q_N(_11309_),
    .Q(\atari2600.tia.diag[50] ));
 sg13g2_dfrbp_1 _28551_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net409),
    .D(net7310),
    .Q_N(_11308_),
    .Q(\atari2600.tia.diag[51] ));
 sg13g2_dfrbp_1 _28552_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net407),
    .D(_02148_),
    .Q_N(_11307_),
    .Q(\atari2600.tia.diag[52] ));
 sg13g2_dfrbp_1 _28553_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net405),
    .D(_02149_),
    .Q_N(_11306_),
    .Q(\atari2600.tia.diag[53] ));
 sg13g2_dfrbp_1 _28554_ (.CLK(clknet_leaf_297_clk),
    .RESET_B(net403),
    .D(_02150_),
    .Q_N(_11305_),
    .Q(\atari2600.tia.diag[54] ));
 sg13g2_dfrbp_1 _28555_ (.CLK(clknet_leaf_327_clk),
    .RESET_B(net401),
    .D(_02151_),
    .Q_N(_11304_),
    .Q(\atari2600.tia.diag[55] ));
 sg13g2_dfrbp_1 _28556_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net399),
    .D(_02152_),
    .Q_N(_11303_),
    .Q(\atari2600.tia.diag[40] ));
 sg13g2_dfrbp_1 _28557_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net397),
    .D(net7274),
    .Q_N(_11302_),
    .Q(\atari2600.tia.diag[41] ));
 sg13g2_dfrbp_1 _28558_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net395),
    .D(_02154_),
    .Q_N(_11301_),
    .Q(\atari2600.tia.diag[42] ));
 sg13g2_dfrbp_1 _28559_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net393),
    .D(_02155_),
    .Q_N(_11300_),
    .Q(\atari2600.tia.diag[43] ));
 sg13g2_dfrbp_1 _28560_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net391),
    .D(_02156_),
    .Q_N(_11299_),
    .Q(\atari2600.tia.diag[44] ));
 sg13g2_dfrbp_1 _28561_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net389),
    .D(_02157_),
    .Q_N(_11298_),
    .Q(\atari2600.tia.diag[45] ));
 sg13g2_dfrbp_1 _28562_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net387),
    .D(_02158_),
    .Q_N(_11297_),
    .Q(\atari2600.tia.diag[46] ));
 sg13g2_dfrbp_1 _28563_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net385),
    .D(_02159_),
    .Q_N(_11296_),
    .Q(\atari2600.tia.diag[47] ));
 sg13g2_dfrbp_1 _28564_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net383),
    .D(_02160_),
    .Q_N(_11295_),
    .Q(\atari2600.tia.diag[32] ));
 sg13g2_dfrbp_1 _28565_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net381),
    .D(net7299),
    .Q_N(_11294_),
    .Q(\atari2600.tia.diag[33] ));
 sg13g2_dfrbp_1 _28566_ (.CLK(clknet_leaf_292_clk),
    .RESET_B(net379),
    .D(_02162_),
    .Q_N(_11293_),
    .Q(\atari2600.tia.diag[34] ));
 sg13g2_dfrbp_1 _28567_ (.CLK(clknet_leaf_296_clk),
    .RESET_B(net377),
    .D(_02163_),
    .Q_N(_11292_),
    .Q(\atari2600.tia.diag[35] ));
 sg13g2_dfrbp_1 _28568_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net375),
    .D(_02164_),
    .Q_N(_11291_),
    .Q(\atari2600.tia.diag[36] ));
 sg13g2_dfrbp_1 _28569_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net373),
    .D(_02165_),
    .Q_N(_11290_),
    .Q(\atari2600.tia.diag[37] ));
 sg13g2_dfrbp_1 _28570_ (.CLK(clknet_leaf_298_clk),
    .RESET_B(net371),
    .D(_02166_),
    .Q_N(_11289_),
    .Q(\atari2600.tia.diag[38] ));
 sg13g2_dfrbp_1 _28571_ (.CLK(clknet_leaf_305_clk),
    .RESET_B(net369),
    .D(_02167_),
    .Q_N(_11288_),
    .Q(\atari2600.tia.diag[39] ));
 sg13g2_dfrbp_1 _28572_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net367),
    .D(_02168_),
    .Q_N(_11287_),
    .Q(\atari2600.tia.diag[88] ));
 sg13g2_dfrbp_1 _28573_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net365),
    .D(_02169_),
    .Q_N(_11286_),
    .Q(\atari2600.tia.diag[89] ));
 sg13g2_dfrbp_1 _28574_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net363),
    .D(_02170_),
    .Q_N(_11285_),
    .Q(\atari2600.tia.diag[90] ));
 sg13g2_dfrbp_1 _28575_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net361),
    .D(_02171_),
    .Q_N(_11284_),
    .Q(\atari2600.tia.diag[91] ));
 sg13g2_dfrbp_1 _28576_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net359),
    .D(_02172_),
    .Q_N(_11283_),
    .Q(\atari2600.tia.diag[92] ));
 sg13g2_dfrbp_1 _28577_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net357),
    .D(_02173_),
    .Q_N(_11282_),
    .Q(\atari2600.tia.diag[93] ));
 sg13g2_dfrbp_1 _28578_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net355),
    .D(_02174_),
    .Q_N(_11281_),
    .Q(\atari2600.tia.diag[94] ));
 sg13g2_dfrbp_1 _28579_ (.CLK(clknet_leaf_314_clk),
    .RESET_B(net353),
    .D(_02175_),
    .Q_N(_11280_),
    .Q(\atari2600.tia.diag[95] ));
 sg13g2_dfrbp_1 _28580_ (.CLK(clknet_leaf_333_clk),
    .RESET_B(net351),
    .D(_02176_),
    .Q_N(_11279_),
    .Q(\atari2600.tia.hmp0[0] ));
 sg13g2_dfrbp_1 _28581_ (.CLK(clknet_leaf_332_clk),
    .RESET_B(net349),
    .D(_02177_),
    .Q_N(_11278_),
    .Q(\atari2600.tia.hmp0[1] ));
 sg13g2_dfrbp_1 _28582_ (.CLK(clknet_leaf_333_clk),
    .RESET_B(net347),
    .D(_02178_),
    .Q_N(_11277_),
    .Q(\atari2600.tia.hmp0[2] ));
 sg13g2_dfrbp_1 _28583_ (.CLK(clknet_leaf_328_clk),
    .RESET_B(net345),
    .D(_02179_),
    .Q_N(_11276_),
    .Q(\atari2600.tia.hmp0[3] ));
 sg13g2_dfrbp_1 _28584_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net343),
    .D(_02180_),
    .Q_N(_11275_),
    .Q(\atari2600.tia.hmp1[0] ));
 sg13g2_dfrbp_1 _28585_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net341),
    .D(_02181_),
    .Q_N(_11274_),
    .Q(\atari2600.tia.hmp1[1] ));
 sg13g2_dfrbp_1 _28586_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net339),
    .D(_02182_),
    .Q_N(_11273_),
    .Q(\atari2600.tia.hmp1[2] ));
 sg13g2_dfrbp_1 _28587_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net337),
    .D(_02183_),
    .Q_N(_11272_),
    .Q(\atari2600.tia.hmp1[3] ));
 sg13g2_dfrbp_1 _28588_ (.CLK(clknet_leaf_332_clk),
    .RESET_B(net335),
    .D(_02184_),
    .Q_N(_11271_),
    .Q(\atari2600.tia.hmm0[0] ));
 sg13g2_dfrbp_1 _28589_ (.CLK(clknet_leaf_332_clk),
    .RESET_B(net333),
    .D(_02185_),
    .Q_N(_11270_),
    .Q(\atari2600.tia.hmm0[1] ));
 sg13g2_dfrbp_1 _28590_ (.CLK(clknet_leaf_331_clk),
    .RESET_B(net331),
    .D(_02186_),
    .Q_N(_11269_),
    .Q(\atari2600.tia.hmm0[2] ));
 sg13g2_dfrbp_1 _28591_ (.CLK(clknet_leaf_328_clk),
    .RESET_B(net329),
    .D(_02187_),
    .Q_N(_11268_),
    .Q(\atari2600.tia.hmm0[3] ));
 sg13g2_dfrbp_1 _28592_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net327),
    .D(_02188_),
    .Q_N(_11267_),
    .Q(\atari2600.tia.hmm1[0] ));
 sg13g2_dfrbp_1 _28593_ (.CLK(clknet_leaf_294_clk),
    .RESET_B(net325),
    .D(_02189_),
    .Q_N(_11266_),
    .Q(\atari2600.tia.hmm1[1] ));
 sg13g2_dfrbp_1 _28594_ (.CLK(clknet_leaf_291_clk),
    .RESET_B(net323),
    .D(_02190_),
    .Q_N(_11265_),
    .Q(\atari2600.tia.hmm1[2] ));
 sg13g2_dfrbp_1 _28595_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net321),
    .D(_02191_),
    .Q_N(_11264_),
    .Q(\atari2600.tia.hmm1[3] ));
 sg13g2_dfrbp_1 _28596_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net319),
    .D(_02192_),
    .Q_N(_11263_),
    .Q(\atari2600.tia.hmbl[0] ));
 sg13g2_dfrbp_1 _28597_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net317),
    .D(_02193_),
    .Q_N(_11262_),
    .Q(\atari2600.tia.hmbl[1] ));
 sg13g2_dfrbp_1 _28598_ (.CLK(clknet_leaf_293_clk),
    .RESET_B(net315),
    .D(_02194_),
    .Q_N(_11261_),
    .Q(\atari2600.tia.hmbl[2] ));
 sg13g2_dfrbp_1 _28599_ (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2185),
    .D(_02195_),
    .Q_N(_13240_),
    .Q(\atari2600.tia.hmbl[3] ));
 sg13g2_dfrbp_1 _28600_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2186),
    .D(_00015_),
    .Q_N(_13241_),
    .Q(\atari2600.tia.cx[0] ));
 sg13g2_dfrbp_1 _28601_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2187),
    .D(_00021_),
    .Q_N(_13242_),
    .Q(\atari2600.tia.cx[1] ));
 sg13g2_dfrbp_1 _28602_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2188),
    .D(_00022_),
    .Q_N(_13243_),
    .Q(\atari2600.tia.cx[2] ));
 sg13g2_dfrbp_1 _28603_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2189),
    .D(_00023_),
    .Q_N(_13244_),
    .Q(\atari2600.tia.cx[3] ));
 sg13g2_dfrbp_1 _28604_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2190),
    .D(_00024_),
    .Q_N(_13245_),
    .Q(\atari2600.tia.cx[4] ));
 sg13g2_dfrbp_1 _28605_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2191),
    .D(_00025_),
    .Q_N(_13246_),
    .Q(\atari2600.tia.cx[5] ));
 sg13g2_dfrbp_1 _28606_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2192),
    .D(_00026_),
    .Q_N(_13247_),
    .Q(\atari2600.tia.cx[6] ));
 sg13g2_dfrbp_1 _28607_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2193),
    .D(_00027_),
    .Q_N(_13248_),
    .Q(\atari2600.tia.cx[7] ));
 sg13g2_dfrbp_1 _28608_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2194),
    .D(_00028_),
    .Q_N(_13249_),
    .Q(\atari2600.tia.cx[8] ));
 sg13g2_dfrbp_1 _28609_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2195),
    .D(_00029_),
    .Q_N(_13250_),
    .Q(\atari2600.tia.cx[9] ));
 sg13g2_dfrbp_1 _28610_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2196),
    .D(_00016_),
    .Q_N(_13251_),
    .Q(\atari2600.tia.cx[10] ));
 sg13g2_dfrbp_1 _28611_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2197),
    .D(_00017_),
    .Q_N(_13252_),
    .Q(\atari2600.tia.cx[11] ));
 sg13g2_dfrbp_1 _28612_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2198),
    .D(_00018_),
    .Q_N(_13253_),
    .Q(\atari2600.tia.cx[12] ));
 sg13g2_dfrbp_1 _28613_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2360),
    .D(_00019_),
    .Q_N(_13254_),
    .Q(\atari2600.tia.cx[13] ));
 sg13g2_dfrbp_1 _28614_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net313),
    .D(_00020_),
    .Q_N(_11260_),
    .Q(\atari2600.tia.cx[14] ));
 sg13g2_dfrbp_1 _28615_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net311),
    .D(_02196_),
    .Q_N(_11259_),
    .Q(\atari2600.tia.cx_clr ));
 sg13g2_dfrbp_1 _28616_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net309),
    .D(_02197_),
    .Q_N(_11258_),
    .Q(\atari2600.tia.audc0[0] ));
 sg13g2_dfrbp_1 _28617_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net307),
    .D(_02198_),
    .Q_N(_11257_),
    .Q(\atari2600.tia.audc0[1] ));
 sg13g2_dfrbp_1 _28618_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net305),
    .D(_02199_),
    .Q_N(_11256_),
    .Q(\atari2600.tia.audc0[2] ));
 sg13g2_dfrbp_1 _28619_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net303),
    .D(_02200_),
    .Q_N(_11255_),
    .Q(\atari2600.tia.audc0[3] ));
 sg13g2_dfrbp_1 _28620_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net301),
    .D(_02201_),
    .Q_N(_11254_),
    .Q(\atari2600.tia.audc1[0] ));
 sg13g2_dfrbp_1 _28621_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net299),
    .D(_02202_),
    .Q_N(_11253_),
    .Q(\atari2600.tia.audc1[1] ));
 sg13g2_dfrbp_1 _28622_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net297),
    .D(_02203_),
    .Q_N(_11252_),
    .Q(\atari2600.tia.audc1[2] ));
 sg13g2_dfrbp_1 _28623_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net295),
    .D(_02204_),
    .Q_N(_11251_),
    .Q(\atari2600.tia.audc1[3] ));
 sg13g2_dfrbp_1 _28624_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net293),
    .D(_02205_),
    .Q_N(_11250_),
    .Q(\atari2600.tia.audv0[0] ));
 sg13g2_dfrbp_1 _28625_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net291),
    .D(_02206_),
    .Q_N(_11249_),
    .Q(\atari2600.tia.audv0[1] ));
 sg13g2_dfrbp_1 _28626_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net289),
    .D(_02207_),
    .Q_N(_11248_),
    .Q(\atari2600.tia.audv0[2] ));
 sg13g2_dfrbp_1 _28627_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net287),
    .D(_02208_),
    .Q_N(_11247_),
    .Q(\atari2600.tia.audv0[3] ));
 sg13g2_dfrbp_1 _28628_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net285),
    .D(_02209_),
    .Q_N(_11246_),
    .Q(\atari2600.tia.audv1[0] ));
 sg13g2_dfrbp_1 _28629_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net283),
    .D(_02210_),
    .Q_N(_11245_),
    .Q(\atari2600.tia.audv1[1] ));
 sg13g2_dfrbp_1 _28630_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net281),
    .D(_02211_),
    .Q_N(_11244_),
    .Q(\atari2600.tia.audv1[2] ));
 sg13g2_dfrbp_1 _28631_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net279),
    .D(_02212_),
    .Q_N(_11243_),
    .Q(\atari2600.tia.audv1[3] ));
 sg13g2_dfrbp_1 _28632_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net277),
    .D(_02213_),
    .Q_N(_00107_),
    .Q(\atari2600.tia.audf0[0] ));
 sg13g2_dfrbp_1 _28633_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net275),
    .D(_02214_),
    .Q_N(_11242_),
    .Q(\atari2600.tia.audf0[1] ));
 sg13g2_dfrbp_1 _28634_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net273),
    .D(_02215_),
    .Q_N(_11241_),
    .Q(\atari2600.tia.audf0[2] ));
 sg13g2_dfrbp_1 _28635_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net271),
    .D(_02216_),
    .Q_N(_11240_),
    .Q(\atari2600.tia.audf0[3] ));
 sg13g2_dfrbp_1 _28636_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net269),
    .D(_02217_),
    .Q_N(_00112_),
    .Q(\atari2600.tia.audf0[4] ));
 sg13g2_dfrbp_1 _28637_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net267),
    .D(_02218_),
    .Q_N(_00139_),
    .Q(\atari2600.tia.audf1[0] ));
 sg13g2_dfrbp_1 _28638_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net265),
    .D(_02219_),
    .Q_N(_11239_),
    .Q(\atari2600.tia.audf1[1] ));
 sg13g2_dfrbp_1 _28639_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net263),
    .D(_02220_),
    .Q_N(_11238_),
    .Q(\atari2600.tia.audf1[2] ));
 sg13g2_dfrbp_1 _28640_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net261),
    .D(_02221_),
    .Q_N(_11237_),
    .Q(\atari2600.tia.audf1[3] ));
 sg13g2_dfrbp_1 _28641_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net259),
    .D(_02222_),
    .Q_N(_00140_),
    .Q(\atari2600.tia.audf1[4] ));
 sg13g2_dfrbp_1 _28642_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net257),
    .D(_02223_),
    .Q_N(_11236_),
    .Q(\atari2600.tia.p4_l ));
 sg13g2_dfrbp_1 _28643_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net255),
    .D(_02224_),
    .Q_N(_11235_),
    .Q(\atari2600.tia.poly4_l.x[1] ));
 sg13g2_dfrbp_1 _28644_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net253),
    .D(net3506),
    .Q_N(_11234_),
    .Q(\atari2600.tia.poly4_l.x[2] ));
 sg13g2_dfrbp_1 _28645_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net251),
    .D(_02226_),
    .Q_N(_11233_),
    .Q(\atari2600.tia.poly4_l.x[3] ));
 sg13g2_dfrbp_1 _28646_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net249),
    .D(net3233),
    .Q_N(_11232_),
    .Q(\atari2600.tia.p5_l ));
 sg13g2_dfrbp_1 _28647_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net247),
    .D(_02228_),
    .Q_N(_11231_),
    .Q(\atari2600.tia.poly5_l.x[1] ));
 sg13g2_dfrbp_1 _28648_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net245),
    .D(_02229_),
    .Q_N(_11230_),
    .Q(\atari2600.tia.poly5_l.x[2] ));
 sg13g2_dfrbp_1 _28649_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net243),
    .D(net3914),
    .Q_N(_11229_),
    .Q(\atari2600.tia.poly5_l.x[3] ));
 sg13g2_dfrbp_1 _28650_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net241),
    .D(net6855),
    .Q_N(_11228_),
    .Q(\atari2600.tia.poly5_l.x[4] ));
 sg13g2_dfrbp_1 _28651_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net239),
    .D(net3802),
    .Q_N(_11227_),
    .Q(\atari2600.tia.p9_l ));
 sg13g2_dfrbp_1 _28652_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net237),
    .D(net3242),
    .Q_N(_11226_),
    .Q(\atari2600.tia.poly9_l.x[1] ));
 sg13g2_dfrbp_1 _28653_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net235),
    .D(_02234_),
    .Q_N(_11225_),
    .Q(\atari2600.tia.poly9_l.x[2] ));
 sg13g2_dfrbp_1 _28654_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net233),
    .D(_02235_),
    .Q_N(_11224_),
    .Q(\atari2600.tia.poly9_l.x[3] ));
 sg13g2_dfrbp_1 _28655_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net231),
    .D(_02236_),
    .Q_N(_11223_),
    .Q(\atari2600.tia.poly9_l.x[4] ));
 sg13g2_dfrbp_1 _28656_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net229),
    .D(_02237_),
    .Q_N(_11222_),
    .Q(\atari2600.tia.poly9_l.x[5] ));
 sg13g2_dfrbp_1 _28657_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net227),
    .D(_02238_),
    .Q_N(_11221_),
    .Q(\atari2600.tia.poly9_l.x[6] ));
 sg13g2_dfrbp_1 _28658_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net225),
    .D(net3943),
    .Q_N(_11220_),
    .Q(\atari2600.tia.poly9_l.x[7] ));
 sg13g2_dfrbp_1 _28659_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net223),
    .D(_02240_),
    .Q_N(_11219_),
    .Q(\atari2600.tia.poly9_l.x[8] ));
 sg13g2_dfrbp_1 _28660_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net221),
    .D(net6878),
    .Q_N(_11218_),
    .Q(\atari2600.tia.p4_r ));
 sg13g2_dfrbp_1 _28661_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net219),
    .D(_02242_),
    .Q_N(_11217_),
    .Q(\atari2600.tia.poly4_r.x[1] ));
 sg13g2_dfrbp_1 _28662_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net217),
    .D(_02243_),
    .Q_N(_11216_),
    .Q(\atari2600.tia.poly4_r.x[2] ));
 sg13g2_dfrbp_1 _28663_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net215),
    .D(net6749),
    .Q_N(_11215_),
    .Q(\atari2600.tia.poly4_r.x[3] ));
 sg13g2_dfrbp_1 _28664_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net213),
    .D(net7168),
    .Q_N(_11214_),
    .Q(\atari2600.tia.p5_r ));
 sg13g2_dfrbp_1 _28665_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net211),
    .D(net3057),
    .Q_N(_11213_),
    .Q(\atari2600.tia.poly5_r.x[1] ));
 sg13g2_dfrbp_1 _28666_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net209),
    .D(_02247_),
    .Q_N(_11212_),
    .Q(\atari2600.tia.poly5_r.x[2] ));
 sg13g2_dfrbp_1 _28667_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net207),
    .D(_02248_),
    .Q_N(_11211_),
    .Q(\atari2600.tia.poly5_r.x[3] ));
 sg13g2_dfrbp_1 _28668_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net205),
    .D(_02249_),
    .Q_N(_11210_),
    .Q(\atari2600.tia.poly5_r.x[4] ));
 sg13g2_dfrbp_1 _28669_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net203),
    .D(net7241),
    .Q_N(_11209_),
    .Q(\atari2600.tia.p9_r ));
 sg13g2_dfrbp_1 _28670_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net201),
    .D(_02251_),
    .Q_N(_11208_),
    .Q(\atari2600.tia.poly9_r.x[1] ));
 sg13g2_dfrbp_1 _28671_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net199),
    .D(_02252_),
    .Q_N(_11207_),
    .Q(\atari2600.tia.poly9_r.x[2] ));
 sg13g2_dfrbp_1 _28672_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net197),
    .D(net4415),
    .Q_N(_11206_),
    .Q(\atari2600.tia.poly9_r.x[3] ));
 sg13g2_dfrbp_1 _28673_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net195),
    .D(net6940),
    .Q_N(_11205_),
    .Q(\atari2600.tia.poly9_r.x[4] ));
 sg13g2_dfrbp_1 _28674_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net193),
    .D(_02255_),
    .Q_N(_11204_),
    .Q(\atari2600.tia.poly9_r.x[5] ));
 sg13g2_dfrbp_1 _28675_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net191),
    .D(_02256_),
    .Q_N(_11203_),
    .Q(\atari2600.tia.poly9_r.x[6] ));
 sg13g2_dfrbp_1 _28676_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net189),
    .D(_02257_),
    .Q_N(_11202_),
    .Q(\atari2600.tia.poly9_r.x[7] ));
 sg13g2_dfrbp_1 _28677_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net187),
    .D(net4358),
    .Q_N(_11201_),
    .Q(\atari2600.tia.poly9_r.x[8] ));
 sg13g2_dfrbp_1 _28678_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net185),
    .D(_02259_),
    .Q_N(_11200_),
    .Q(\scanline[67][0] ));
 sg13g2_dfrbp_1 _28679_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net184),
    .D(_02260_),
    .Q_N(_11199_),
    .Q(\scanline[67][1] ));
 sg13g2_dfrbp_1 _28680_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net183),
    .D(_02261_),
    .Q_N(_11198_),
    .Q(\scanline[67][2] ));
 sg13g2_dfrbp_1 _28681_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net182),
    .D(_02262_),
    .Q_N(_11197_),
    .Q(\scanline[67][3] ));
 sg13g2_dfrbp_1 _28682_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net181),
    .D(_02263_),
    .Q_N(_11196_),
    .Q(\scanline[67][4] ));
 sg13g2_dfrbp_1 _28683_ (.CLK(clknet_leaf_282_clk),
    .RESET_B(net180),
    .D(_02264_),
    .Q_N(_11195_),
    .Q(\scanline[67][5] ));
 sg13g2_dfrbp_1 _28684_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net179),
    .D(_02265_),
    .Q_N(_11194_),
    .Q(\scanline[67][6] ));
 sg13g2_dfrbp_1 _28685_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net178),
    .D(_02266_),
    .Q_N(_11193_),
    .Q(\scanline[9][0] ));
 sg13g2_dfrbp_1 _28686_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net177),
    .D(_02267_),
    .Q_N(_11192_),
    .Q(\scanline[9][1] ));
 sg13g2_dfrbp_1 _28687_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net176),
    .D(_02268_),
    .Q_N(_11191_),
    .Q(\scanline[9][2] ));
 sg13g2_dfrbp_1 _28688_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net175),
    .D(_02269_),
    .Q_N(_11190_),
    .Q(\scanline[9][3] ));
 sg13g2_dfrbp_1 _28689_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net174),
    .D(_02270_),
    .Q_N(_11189_),
    .Q(\scanline[9][4] ));
 sg13g2_dfrbp_1 _28690_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net173),
    .D(_02271_),
    .Q_N(_11188_),
    .Q(\scanline[9][5] ));
 sg13g2_dfrbp_1 _28691_ (.CLK(clknet_leaf_272_clk),
    .RESET_B(net172),
    .D(_02272_),
    .Q_N(_11187_),
    .Q(\scanline[9][6] ));
 sg13g2_dfrbp_1 _28692_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net171),
    .D(_02273_),
    .Q_N(_11186_),
    .Q(\scanline[66][0] ));
 sg13g2_dfrbp_1 _28693_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net170),
    .D(_02274_),
    .Q_N(_11185_),
    .Q(\scanline[66][1] ));
 sg13g2_dfrbp_1 _28694_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net169),
    .D(_02275_),
    .Q_N(_11184_),
    .Q(\scanline[66][2] ));
 sg13g2_dfrbp_1 _28695_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net168),
    .D(_02276_),
    .Q_N(_11183_),
    .Q(\scanline[66][3] ));
 sg13g2_dfrbp_1 _28696_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net167),
    .D(_02277_),
    .Q_N(_11182_),
    .Q(\scanline[66][4] ));
 sg13g2_dfrbp_1 _28697_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net166),
    .D(_02278_),
    .Q_N(_11181_),
    .Q(\scanline[66][5] ));
 sg13g2_dfrbp_1 _28698_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net165),
    .D(_02279_),
    .Q_N(_11180_),
    .Q(\scanline[66][6] ));
 sg13g2_dfrbp_1 _28699_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net164),
    .D(_02280_),
    .Q_N(_11179_),
    .Q(\scanline[6][0] ));
 sg13g2_dfrbp_1 _28700_ (.CLK(clknet_leaf_270_clk),
    .RESET_B(net163),
    .D(_02281_),
    .Q_N(_11178_),
    .Q(\scanline[6][1] ));
 sg13g2_dfrbp_1 _28701_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net162),
    .D(_02282_),
    .Q_N(_11177_),
    .Q(\scanline[6][2] ));
 sg13g2_dfrbp_1 _28702_ (.CLK(clknet_leaf_268_clk),
    .RESET_B(net161),
    .D(_02283_),
    .Q_N(_11176_),
    .Q(\scanline[6][3] ));
 sg13g2_dfrbp_1 _28703_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net160),
    .D(_02284_),
    .Q_N(_11175_),
    .Q(\scanline[6][4] ));
 sg13g2_dfrbp_1 _28704_ (.CLK(clknet_leaf_263_clk),
    .RESET_B(net159),
    .D(_02285_),
    .Q_N(_11174_),
    .Q(\scanline[6][5] ));
 sg13g2_dfrbp_1 _28705_ (.CLK(clknet_leaf_269_clk),
    .RESET_B(net158),
    .D(_02286_),
    .Q_N(_11173_),
    .Q(\scanline[6][6] ));
 sg13g2_dfrbp_1 _28706_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net157),
    .D(_02287_),
    .Q_N(_11172_),
    .Q(\scanline[62][0] ));
 sg13g2_dfrbp_1 _28707_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net156),
    .D(_02288_),
    .Q_N(_11171_),
    .Q(\scanline[62][1] ));
 sg13g2_dfrbp_1 _28708_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net155),
    .D(_02289_),
    .Q_N(_11170_),
    .Q(\scanline[62][2] ));
 sg13g2_dfrbp_1 _28709_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net154),
    .D(_02290_),
    .Q_N(_11169_),
    .Q(\scanline[62][3] ));
 sg13g2_dfrbp_1 _28710_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net153),
    .D(_02291_),
    .Q_N(_11168_),
    .Q(\scanline[62][4] ));
 sg13g2_dfrbp_1 _28711_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net152),
    .D(_02292_),
    .Q_N(_11167_),
    .Q(\scanline[62][5] ));
 sg13g2_dfrbp_1 _28712_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net151),
    .D(_02293_),
    .Q_N(_11166_),
    .Q(\scanline[62][6] ));
 sg13g2_dfrbp_1 _28713_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net150),
    .D(_02294_),
    .Q_N(_11165_),
    .Q(\scanline[63][0] ));
 sg13g2_dfrbp_1 _28714_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net149),
    .D(_02295_),
    .Q_N(_11164_),
    .Q(\scanline[63][1] ));
 sg13g2_dfrbp_1 _28715_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net148),
    .D(_02296_),
    .Q_N(_11163_),
    .Q(\scanline[63][2] ));
 sg13g2_dfrbp_1 _28716_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net147),
    .D(_02297_),
    .Q_N(_11162_),
    .Q(\scanline[63][3] ));
 sg13g2_dfrbp_1 _28717_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net146),
    .D(_02298_),
    .Q_N(_11161_),
    .Q(\scanline[63][4] ));
 sg13g2_dfrbp_1 _28718_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net145),
    .D(_02299_),
    .Q_N(_11160_),
    .Q(\scanline[63][5] ));
 sg13g2_dfrbp_1 _28719_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net144),
    .D(_02300_),
    .Q_N(_11159_),
    .Q(\scanline[63][6] ));
 sg13g2_dfrbp_1 _28720_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net143),
    .D(net6324),
    .Q_N(_11158_),
    .Q(\atari2600.pia.interval[0] ));
 sg13g2_dfrbp_1 _28721_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net142),
    .D(_02302_),
    .Q_N(_11157_),
    .Q(\scanline[37][0] ));
 sg13g2_dfrbp_1 _28722_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net141),
    .D(_02303_),
    .Q_N(_11156_),
    .Q(\scanline[37][1] ));
 sg13g2_dfrbp_1 _28723_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net140),
    .D(_02304_),
    .Q_N(_11155_),
    .Q(\scanline[37][2] ));
 sg13g2_dfrbp_1 _28724_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net139),
    .D(_02305_),
    .Q_N(_11154_),
    .Q(\scanline[37][3] ));
 sg13g2_dfrbp_1 _28725_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net138),
    .D(_02306_),
    .Q_N(_11153_),
    .Q(\scanline[37][4] ));
 sg13g2_dfrbp_1 _28726_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net137),
    .D(_02307_),
    .Q_N(_11152_),
    .Q(\scanline[37][5] ));
 sg13g2_dfrbp_1 _28727_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net136),
    .D(_02308_),
    .Q_N(_11151_),
    .Q(\scanline[37][6] ));
 sg13g2_dfrbp_1 _28728_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net135),
    .D(net3156),
    .Q_N(_11150_),
    .Q(\atari2600.pia.instat[0] ));
 sg13g2_dfrbp_1 _28729_ (.CLK(clknet_leaf_271_clk),
    .RESET_B(net134),
    .D(_02310_),
    .Q_N(_11149_),
    .Q(\scanline[36][0] ));
 sg13g2_dfrbp_1 _28730_ (.CLK(clknet_leaf_276_clk),
    .RESET_B(net133),
    .D(_02311_),
    .Q_N(_11148_),
    .Q(\scanline[36][1] ));
 sg13g2_dfrbp_1 _28731_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net132),
    .D(_02312_),
    .Q_N(_11147_),
    .Q(\scanline[36][2] ));
 sg13g2_dfrbp_1 _28732_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net131),
    .D(_02313_),
    .Q_N(_11146_),
    .Q(\scanline[36][3] ));
 sg13g2_dfrbp_1 _28733_ (.CLK(clknet_leaf_278_clk),
    .RESET_B(net130),
    .D(_02314_),
    .Q_N(_11145_),
    .Q(\scanline[36][4] ));
 sg13g2_dfrbp_1 _28734_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net129),
    .D(_02315_),
    .Q_N(_11144_),
    .Q(\scanline[36][5] ));
 sg13g2_dfrbp_1 _28735_ (.CLK(clknet_leaf_277_clk),
    .RESET_B(net128),
    .D(_02316_),
    .Q_N(_11143_),
    .Q(\scanline[36][6] ));
 sg13g2_dfrbp_1 _28736_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net127),
    .D(_02317_),
    .Q_N(_11142_),
    .Q(\scanline[65][0] ));
 sg13g2_dfrbp_1 _28737_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net126),
    .D(_02318_),
    .Q_N(_11141_),
    .Q(\scanline[65][1] ));
 sg13g2_dfrbp_1 _28738_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net125),
    .D(_02319_),
    .Q_N(_11140_),
    .Q(\scanline[65][2] ));
 sg13g2_dfrbp_1 _28739_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net124),
    .D(_02320_),
    .Q_N(_11139_),
    .Q(\scanline[65][3] ));
 sg13g2_dfrbp_1 _28740_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net123),
    .D(_02321_),
    .Q_N(_11138_),
    .Q(\scanline[65][4] ));
 sg13g2_dfrbp_1 _28741_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net122),
    .D(_02322_),
    .Q_N(_11137_),
    .Q(\scanline[65][5] ));
 sg13g2_dfrbp_1 _28742_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net121),
    .D(_02323_),
    .Q_N(_11136_),
    .Q(\scanline[65][6] ));
 sg13g2_dfrbp_1 _28743_ (.CLK(clknet_leaf_302_clk),
    .RESET_B(net120),
    .D(_02324_),
    .Q_N(_11135_),
    .Q(\scanline[64][0] ));
 sg13g2_dfrbp_1 _28744_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net119),
    .D(_02325_),
    .Q_N(_11134_),
    .Q(\scanline[64][1] ));
 sg13g2_dfrbp_1 _28745_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net118),
    .D(_02326_),
    .Q_N(_11133_),
    .Q(\scanline[64][2] ));
 sg13g2_dfrbp_1 _28746_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net117),
    .D(_02327_),
    .Q_N(_11132_),
    .Q(\scanline[64][3] ));
 sg13g2_dfrbp_1 _28747_ (.CLK(clknet_leaf_280_clk),
    .RESET_B(net116),
    .D(_02328_),
    .Q_N(_11131_),
    .Q(\scanline[64][4] ));
 sg13g2_dfrbp_1 _28748_ (.CLK(clknet_leaf_281_clk),
    .RESET_B(net115),
    .D(_02329_),
    .Q_N(_11130_),
    .Q(\scanline[64][5] ));
 sg13g2_dfrbp_1 _28749_ (.CLK(clknet_leaf_279_clk),
    .RESET_B(net114),
    .D(_02330_),
    .Q_N(_11129_),
    .Q(\scanline[64][6] ));
 sg13g2_dfrbp_1 _28750_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net113),
    .D(_02331_),
    .Q_N(_11128_),
    .Q(\atari2600.ram[47][0] ));
 sg13g2_dfrbp_1 _28751_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net112),
    .D(_02332_),
    .Q_N(_11127_),
    .Q(\atari2600.ram[47][1] ));
 sg13g2_dfrbp_1 _28752_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net111),
    .D(_02333_),
    .Q_N(_11126_),
    .Q(\atari2600.ram[47][2] ));
 sg13g2_dfrbp_1 _28753_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net110),
    .D(_02334_),
    .Q_N(_11125_),
    .Q(\atari2600.ram[47][3] ));
 sg13g2_dfrbp_1 _28754_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net109),
    .D(_02335_),
    .Q_N(_11124_),
    .Q(\atari2600.ram[47][4] ));
 sg13g2_dfrbp_1 _28755_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net108),
    .D(_02336_),
    .Q_N(_11123_),
    .Q(\atari2600.ram[47][5] ));
 sg13g2_dfrbp_1 _28756_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net107),
    .D(_02337_),
    .Q_N(_11122_),
    .Q(\atari2600.ram[47][6] ));
 sg13g2_dfrbp_1 _28757_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net106),
    .D(_02338_),
    .Q_N(_11121_),
    .Q(\atari2600.ram[47][7] ));
 sg13g2_dfrbp_1 _28758_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net105),
    .D(_02339_),
    .Q_N(_11120_),
    .Q(\atari2600.ram[46][0] ));
 sg13g2_dfrbp_1 _28759_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net104),
    .D(_02340_),
    .Q_N(_11119_),
    .Q(\atari2600.ram[46][1] ));
 sg13g2_dfrbp_1 _28760_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net103),
    .D(_02341_),
    .Q_N(_11118_),
    .Q(\atari2600.ram[46][2] ));
 sg13g2_dfrbp_1 _28761_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net102),
    .D(_02342_),
    .Q_N(_11117_),
    .Q(\atari2600.ram[46][3] ));
 sg13g2_dfrbp_1 _28762_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net101),
    .D(_02343_),
    .Q_N(_11116_),
    .Q(\atari2600.ram[46][4] ));
 sg13g2_dfrbp_1 _28763_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net100),
    .D(_02344_),
    .Q_N(_11115_),
    .Q(\atari2600.ram[46][5] ));
 sg13g2_dfrbp_1 _28764_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net99),
    .D(_02345_),
    .Q_N(_11114_),
    .Q(\atari2600.ram[46][6] ));
 sg13g2_dfrbp_1 _28765_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net98),
    .D(_02346_),
    .Q_N(_11113_),
    .Q(\atari2600.ram[46][7] ));
 sg13g2_dfrbp_1 _28766_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net97),
    .D(_02347_),
    .Q_N(_11112_),
    .Q(\atari2600.ram[45][0] ));
 sg13g2_dfrbp_1 _28767_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net96),
    .D(_02348_),
    .Q_N(_11111_),
    .Q(\atari2600.ram[45][1] ));
 sg13g2_dfrbp_1 _28768_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net95),
    .D(_02349_),
    .Q_N(_11110_),
    .Q(\atari2600.ram[45][2] ));
 sg13g2_dfrbp_1 _28769_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net94),
    .D(_02350_),
    .Q_N(_11109_),
    .Q(\atari2600.ram[45][3] ));
 sg13g2_dfrbp_1 _28770_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net93),
    .D(_02351_),
    .Q_N(_11108_),
    .Q(\atari2600.ram[45][4] ));
 sg13g2_dfrbp_1 _28771_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net92),
    .D(_02352_),
    .Q_N(_11107_),
    .Q(\atari2600.ram[45][5] ));
 sg13g2_dfrbp_1 _28772_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net91),
    .D(_02353_),
    .Q_N(_11106_),
    .Q(\atari2600.ram[45][6] ));
 sg13g2_dfrbp_1 _28773_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net90),
    .D(_02354_),
    .Q_N(_11105_),
    .Q(\atari2600.ram[45][7] ));
 sg13g2_dfrbp_1 _28774_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net89),
    .D(_02355_),
    .Q_N(_11104_),
    .Q(\atari2600.ram[44][0] ));
 sg13g2_dfrbp_1 _28775_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net88),
    .D(_02356_),
    .Q_N(_11103_),
    .Q(\atari2600.ram[44][1] ));
 sg13g2_dfrbp_1 _28776_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net87),
    .D(_02357_),
    .Q_N(_11102_),
    .Q(\atari2600.ram[44][2] ));
 sg13g2_dfrbp_1 _28777_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net86),
    .D(_02358_),
    .Q_N(_11101_),
    .Q(\atari2600.ram[44][3] ));
 sg13g2_dfrbp_1 _28778_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net85),
    .D(_02359_),
    .Q_N(_11100_),
    .Q(\atari2600.ram[44][4] ));
 sg13g2_dfrbp_1 _28779_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net84),
    .D(_02360_),
    .Q_N(_11099_),
    .Q(\atari2600.ram[44][5] ));
 sg13g2_dfrbp_1 _28780_ (.CLK(clknet_leaf_350_clk),
    .RESET_B(net83),
    .D(_02361_),
    .Q_N(_11098_),
    .Q(\atari2600.ram[44][6] ));
 sg13g2_dfrbp_1 _28781_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net82),
    .D(_02362_),
    .Q_N(_11097_),
    .Q(\atari2600.ram[44][7] ));
 sg13g2_dfrbp_1 _28782_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net81),
    .D(_02363_),
    .Q_N(_11096_),
    .Q(\atari2600.ram[30][0] ));
 sg13g2_dfrbp_1 _28783_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net80),
    .D(_02364_),
    .Q_N(_11095_),
    .Q(\atari2600.ram[30][1] ));
 sg13g2_dfrbp_1 _28784_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net79),
    .D(_02365_),
    .Q_N(_11094_),
    .Q(\atari2600.ram[30][2] ));
 sg13g2_dfrbp_1 _28785_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net78),
    .D(_02366_),
    .Q_N(_11093_),
    .Q(\atari2600.ram[30][3] ));
 sg13g2_dfrbp_1 _28786_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net77),
    .D(_02367_),
    .Q_N(_11092_),
    .Q(\atari2600.ram[30][4] ));
 sg13g2_dfrbp_1 _28787_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net76),
    .D(_02368_),
    .Q_N(_11091_),
    .Q(\atari2600.ram[30][5] ));
 sg13g2_dfrbp_1 _28788_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net75),
    .D(_02369_),
    .Q_N(_11090_),
    .Q(\atari2600.ram[30][6] ));
 sg13g2_dfrbp_1 _28789_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net74),
    .D(_02370_),
    .Q_N(_11089_),
    .Q(\atari2600.ram[30][7] ));
 sg13g2_dfrbp_1 _28790_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net73),
    .D(_02371_),
    .Q_N(_00090_),
    .Q(\atari2600.cpu.AXYS[1][0] ));
 sg13g2_dfrbp_1 _28791_ (.CLK(clknet_leaf_361_clk),
    .RESET_B(net72),
    .D(_02372_),
    .Q_N(_00084_),
    .Q(\atari2600.cpu.AXYS[1][1] ));
 sg13g2_dfrbp_1 _28792_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net71),
    .D(_02373_),
    .Q_N(_11088_),
    .Q(\atari2600.cpu.AXYS[1][2] ));
 sg13g2_dfrbp_1 _28793_ (.CLK(clknet_leaf_362_clk),
    .RESET_B(net70),
    .D(_02374_),
    .Q_N(_11087_),
    .Q(\atari2600.cpu.AXYS[1][3] ));
 sg13g2_dfrbp_1 _28794_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net69),
    .D(_02375_),
    .Q_N(_11086_),
    .Q(\atari2600.cpu.AXYS[1][4] ));
 sg13g2_dfrbp_1 _28795_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net68),
    .D(_02376_),
    .Q_N(_11085_),
    .Q(\atari2600.cpu.AXYS[1][5] ));
 sg13g2_dfrbp_1 _28796_ (.CLK(clknet_leaf_360_clk),
    .RESET_B(net67),
    .D(_02377_),
    .Q_N(_11084_),
    .Q(\atari2600.cpu.AXYS[1][6] ));
 sg13g2_dfrbp_1 _28797_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net66),
    .D(_02378_),
    .Q_N(_11083_),
    .Q(\atari2600.cpu.AXYS[1][7] ));
 sg13g2_dfrbp_1 _28798_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net65),
    .D(_02379_),
    .Q_N(_11082_),
    .Q(\atari2600.tia.diag[76] ));
 sg13g2_dfrbp_1 _28799_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net63),
    .D(_02380_),
    .Q_N(_11081_),
    .Q(\atari2600.tia.diag[77] ));
 sg13g2_dfrbp_1 _28800_ (.CLK(clknet_leaf_311_clk),
    .RESET_B(net61),
    .D(_02381_),
    .Q_N(_11080_),
    .Q(\atari2600.tia.diag[78] ));
 sg13g2_dfrbp_1 _28801_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net59),
    .D(_02382_),
    .Q_N(_11079_),
    .Q(\atari2600.tia.diag[79] ));
 sg13g2_dfrbp_1 _28802_ (.CLK(clknet_leaf_315_clk),
    .RESET_B(net57),
    .D(_02383_),
    .Q_N(_11078_),
    .Q(\atari2600.tia.diag[80] ));
 sg13g2_dfrbp_1 _28803_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net55),
    .D(_02384_),
    .Q_N(_11077_),
    .Q(\atari2600.tia.diag[81] ));
 sg13g2_dfrbp_1 _28804_ (.CLK(clknet_leaf_310_clk),
    .RESET_B(net53),
    .D(_02385_),
    .Q_N(_11076_),
    .Q(\atari2600.tia.diag[82] ));
 sg13g2_dfrbp_1 _28805_ (.CLK(clknet_leaf_309_clk),
    .RESET_B(net51),
    .D(_02386_),
    .Q_N(_11075_),
    .Q(\atari2600.tia.diag[83] ));
 sg13g2_dfrbp_1 _28806_ (.CLK(clknet_leaf_312_clk),
    .RESET_B(net49),
    .D(_02387_),
    .Q_N(_11074_),
    .Q(\atari2600.tia.diag[84] ));
 sg13g2_dfrbp_1 _28807_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net47),
    .D(_02388_),
    .Q_N(_11073_),
    .Q(\atari2600.tia.diag[85] ));
 sg13g2_dfrbp_1 _28808_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net45),
    .D(_02389_),
    .Q_N(_11072_),
    .Q(\atari2600.tia.diag[86] ));
 sg13g2_dfrbp_1 _28809_ (.CLK(clknet_leaf_313_clk),
    .RESET_B(net43),
    .D(_02390_),
    .Q_N(_11071_),
    .Q(\atari2600.tia.diag[87] ));
 sg13g2_dfrbp_1 _28810_ (.CLK(clknet_leaf_362_clk),
    .RESET_B(net41),
    .D(_02391_),
    .Q_N(_00089_),
    .Q(\atari2600.cpu.AXYS[0][0] ));
 sg13g2_dfrbp_1 _28811_ (.CLK(clknet_leaf_361_clk),
    .RESET_B(net40),
    .D(_02392_),
    .Q_N(_00083_),
    .Q(\atari2600.cpu.AXYS[0][1] ));
 sg13g2_dfrbp_1 _28812_ (.CLK(clknet_leaf_361_clk),
    .RESET_B(net39),
    .D(_02393_),
    .Q_N(_11070_),
    .Q(\atari2600.cpu.AXYS[0][2] ));
 sg13g2_dfrbp_1 _28813_ (.CLK(clknet_leaf_362_clk),
    .RESET_B(net38),
    .D(_02394_),
    .Q_N(_11069_),
    .Q(\atari2600.cpu.AXYS[0][3] ));
 sg13g2_dfrbp_1 _28814_ (.CLK(clknet_leaf_359_clk),
    .RESET_B(net37),
    .D(_02395_),
    .Q_N(_11068_),
    .Q(\atari2600.cpu.AXYS[0][4] ));
 sg13g2_dfrbp_1 _28815_ (.CLK(clknet_leaf_359_clk),
    .RESET_B(net36),
    .D(_02396_),
    .Q_N(_11067_),
    .Q(\atari2600.cpu.AXYS[0][5] ));
 sg13g2_dfrbp_1 _28816_ (.CLK(clknet_leaf_360_clk),
    .RESET_B(net35),
    .D(_02397_),
    .Q_N(_11066_),
    .Q(\atari2600.cpu.AXYS[0][6] ));
 sg13g2_dfrbp_1 _28817_ (.CLK(clknet_leaf_360_clk),
    .RESET_B(net34),
    .D(_02398_),
    .Q_N(_11065_),
    .Q(\atari2600.cpu.AXYS[0][7] ));
 sg13g2_dfrbp_1 _28818_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net33),
    .D(_02399_),
    .Q_N(_11064_),
    .Q(\atari2600.ram[24][0] ));
 sg13g2_dfrbp_1 _28819_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net32),
    .D(_02400_),
    .Q_N(_11063_),
    .Q(\atari2600.ram[24][1] ));
 sg13g2_dfrbp_1 _28820_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net31),
    .D(_02401_),
    .Q_N(_11062_),
    .Q(\atari2600.ram[24][2] ));
 sg13g2_dfrbp_1 _28821_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net30),
    .D(_02402_),
    .Q_N(_11061_),
    .Q(\atari2600.ram[24][3] ));
 sg13g2_dfrbp_1 _28822_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net29),
    .D(_02403_),
    .Q_N(_11060_),
    .Q(\atari2600.ram[24][4] ));
 sg13g2_dfrbp_1 _28823_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net28),
    .D(_02404_),
    .Q_N(_11059_),
    .Q(\atari2600.ram[24][5] ));
 sg13g2_dfrbp_1 _28824_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net27),
    .D(_02405_),
    .Q_N(_11058_),
    .Q(\atari2600.ram[24][6] ));
 sg13g2_dfrbp_1 _28825_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2361),
    .D(_02406_),
    .Q_N(_13255_),
    .Q(\atari2600.ram[24][7] ));
 sg13g2_dfrbp_1 _28826_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net2362),
    .D(_00011_),
    .Q_N(_13256_),
    .Q(\atari2600.tia.p1_copies[1] ));
 sg13g2_dfrbp_1 _28827_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2363),
    .D(_00012_),
    .Q_N(_13257_),
    .Q(\atari2600.tia.p1_copies[2] ));
 sg13g2_dfrbp_1 _28828_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net2412),
    .D(_00009_),
    .Q_N(_13258_),
    .Q(\atari2600.tia.p0_copies[1] ));
 sg13g2_dfrbp_1 _28829_ (.CLK(clknet_leaf_306_clk),
    .RESET_B(net26),
    .D(_00010_),
    .Q_N(_11057_),
    .Q(\atari2600.tia.p0_copies[2] ));
 sg13g2_dfrbp_1 _28830_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net25),
    .D(_02407_),
    .Q_N(_00094_),
    .Q(\atari2600.cpu.DI[0] ));
 sg13g2_dfrbp_1 _28831_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net24),
    .D(_02408_),
    .Q_N(_00088_),
    .Q(\atari2600.cpu.DI[1] ));
 sg13g2_dfrbp_1 _28832_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net23),
    .D(_02409_),
    .Q_N(_11056_),
    .Q(\atari2600.cpu.DI[2] ));
 sg13g2_dfrbp_1 _28833_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net22),
    .D(_02410_),
    .Q_N(_11055_),
    .Q(\atari2600.cpu.DI[3] ));
 sg13g2_dfrbp_1 _28834_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net21),
    .D(_02411_),
    .Q_N(_11054_),
    .Q(\atari2600.cpu.DI[4] ));
 sg13g2_dfrbp_1 _28835_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net20),
    .D(_02412_),
    .Q_N(_11053_),
    .Q(\atari2600.cpu.DI[5] ));
 sg13g2_dfrbp_1 _28836_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net19),
    .D(_02413_),
    .Q_N(_11052_),
    .Q(\atari2600.cpu.DI[6] ));
 sg13g2_dfrbp_1 _28837_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net18),
    .D(_02414_),
    .Q_N(_11051_),
    .Q(\atari2600.cpu.DI[7] ));
 sg13g2_dfrbp_1 _28838_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net17),
    .D(_02415_),
    .Q_N(_11050_),
    .Q(\atari2600.cpu.cond_code[0] ));
 sg13g2_dfrbp_1 _28839_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net16),
    .D(_02416_),
    .Q_N(_11049_),
    .Q(\atari2600.cpu.cond_code[1] ));
 sg13g2_dfrbp_1 _28840_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net15),
    .D(_02417_),
    .Q_N(_00058_),
    .Q(\atari2600.cpu.cond_code[2] ));
 sg13g2_dfrbp_1 _28841_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net14),
    .D(_02418_),
    .Q_N(_00145_),
    .Q(\atari2600.cpu.plp ));
 sg13g2_dfrbp_1 _28842_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net13),
    .D(_02419_),
    .Q_N(_11048_),
    .Q(\atari2600.cpu.php ));
 sg13g2_dfrbp_1 _28843_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net12),
    .D(_02420_),
    .Q_N(_00057_),
    .Q(\atari2600.cpu.clc ));
 sg13g2_dfrbp_1 _28844_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2885),
    .D(_02421_),
    .Q_N(_11047_),
    .Q(\atari2600.cpu.sec ));
 sg13g2_dfrbp_1 _28845_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2884),
    .D(_02422_),
    .Q_N(_00055_),
    .Q(\atari2600.cpu.cld ));
 sg13g2_dfrbp_1 _28846_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2883),
    .D(_02423_),
    .Q_N(_11046_),
    .Q(\atari2600.cpu.sed ));
 sg13g2_dfrbp_1 _28847_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2882),
    .D(_02424_),
    .Q_N(_00056_),
    .Q(\atari2600.cpu.cli ));
 sg13g2_dfrbp_1 _28848_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2881),
    .D(_02425_),
    .Q_N(_11045_),
    .Q(\atari2600.cpu.sei ));
 sg13g2_dfrbp_1 _28849_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2880),
    .D(_02426_),
    .Q_N(_11044_),
    .Q(\scanline[35][0] ));
 sg13g2_dfrbp_1 _28850_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2879),
    .D(_02427_),
    .Q_N(_11043_),
    .Q(\scanline[35][1] ));
 sg13g2_dfrbp_1 _28851_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2878),
    .D(_02428_),
    .Q_N(_11042_),
    .Q(\scanline[35][2] ));
 sg13g2_dfrbp_1 _28852_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2877),
    .D(_02429_),
    .Q_N(_11041_),
    .Q(\scanline[35][3] ));
 sg13g2_dfrbp_1 _28853_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2876),
    .D(_02430_),
    .Q_N(_11040_),
    .Q(\scanline[35][4] ));
 sg13g2_dfrbp_1 _28854_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2875),
    .D(_02431_),
    .Q_N(_11039_),
    .Q(\scanline[35][5] ));
 sg13g2_dfrbp_1 _28855_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2874),
    .D(_02432_),
    .Q_N(_11038_),
    .Q(\scanline[35][6] ));
 sg13g2_dfrbp_1 _28856_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2873),
    .D(_02433_),
    .Q_N(_11037_),
    .Q(\atari2600.cpu.clv ));
 sg13g2_dfrbp_1 _28857_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net2872),
    .D(_02434_),
    .Q_N(_11036_),
    .Q(\atari2600.cpu.bit_ins ));
 sg13g2_dfrbp_1 _28858_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2871),
    .D(_02435_),
    .Q_N(_11035_),
    .Q(\atari2600.cpu.rotate ));
 sg13g2_dfrbp_1 _28859_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net2870),
    .D(_02436_),
    .Q_N(_11034_),
    .Q(\atari2600.cpu.shift_right ));
 sg13g2_dfrbp_1 _28860_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net2869),
    .D(_02437_),
    .Q_N(_11033_),
    .Q(\atari2600.cpu.compare ));
 sg13g2_dfrbp_1 _28861_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net2868),
    .D(_02438_),
    .Q_N(_11032_),
    .Q(\atari2600.cpu.adc_bcd ));
 sg13g2_dfrbp_1 _28862_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2866),
    .D(_02439_),
    .Q_N(_11031_),
    .Q(\atari2600.cpu.shift ));
 sg13g2_dfrbp_1 _28863_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net2865),
    .D(_02440_),
    .Q_N(_11030_),
    .Q(\atari2600.cpu.adc_sbc ));
 sg13g2_dfrbp_1 _28864_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2864),
    .D(_02441_),
    .Q_N(_11029_),
    .Q(\atari2600.cpu.inc ));
 sg13g2_dfrbp_1 _28865_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2863),
    .D(_02442_),
    .Q_N(_11028_),
    .Q(\atari2600.cpu.load_only ));
 sg13g2_dfrbp_1 _28866_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2862),
    .D(_02443_),
    .Q_N(_00141_),
    .Q(\atari2600.cpu.write_back ));
 sg13g2_dfrbp_1 _28867_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net2861),
    .D(_02444_),
    .Q_N(_11027_),
    .Q(\atari2600.cpu.store ));
 sg13g2_dfrbp_1 _28868_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2860),
    .D(_02445_),
    .Q_N(_11026_),
    .Q(\atari2600.cpu.index_y ));
 sg13g2_dfrbp_1 _28869_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net2859),
    .D(_02446_),
    .Q_N(_11025_),
    .Q(\atari2600.cpu.res ));
 sg13g2_dfrbp_1 _28870_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2857),
    .D(_02447_),
    .Q_N(_11024_),
    .Q(\atari2600.ram[91][0] ));
 sg13g2_dfrbp_1 _28871_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2856),
    .D(_02448_),
    .Q_N(_11023_),
    .Q(\atari2600.ram[91][1] ));
 sg13g2_dfrbp_1 _28872_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2855),
    .D(_02449_),
    .Q_N(_11022_),
    .Q(\atari2600.ram[91][2] ));
 sg13g2_dfrbp_1 _28873_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2854),
    .D(_02450_),
    .Q_N(_11021_),
    .Q(\atari2600.ram[91][3] ));
 sg13g2_dfrbp_1 _28874_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2853),
    .D(_02451_),
    .Q_N(_11020_),
    .Q(\atari2600.ram[91][4] ));
 sg13g2_dfrbp_1 _28875_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net2852),
    .D(_02452_),
    .Q_N(_11019_),
    .Q(\atari2600.ram[91][5] ));
 sg13g2_dfrbp_1 _28876_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2851),
    .D(_02453_),
    .Q_N(_11018_),
    .Q(\atari2600.ram[91][6] ));
 sg13g2_dfrbp_1 _28877_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2413),
    .D(_02454_),
    .Q_N(_13259_),
    .Q(\atari2600.ram[91][7] ));
 sg13g2_dfrbp_1 _28878_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2414),
    .D(\atari2600.cpu.DIMUX[0] ),
    .Q_N(_00093_),
    .Q(\atari2600.cpu.DIHOLD[0] ));
 sg13g2_dfrbp_1 _28879_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2415),
    .D(\atari2600.cpu.DIMUX[1] ),
    .Q_N(_00087_),
    .Q(\atari2600.cpu.DIHOLD[1] ));
 sg13g2_dfrbp_1 _28880_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2416),
    .D(\atari2600.cpu.DIMUX[2] ),
    .Q_N(_13260_),
    .Q(\atari2600.cpu.DIHOLD[2] ));
 sg13g2_dfrbp_1 _28881_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2417),
    .D(\atari2600.cpu.DIMUX[3] ),
    .Q_N(_13261_),
    .Q(\atari2600.cpu.DIHOLD[3] ));
 sg13g2_dfrbp_1 _28882_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2418),
    .D(\atari2600.cpu.DIMUX[4] ),
    .Q_N(_13262_),
    .Q(\atari2600.cpu.DIHOLD[4] ));
 sg13g2_dfrbp_1 _28883_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2419),
    .D(net5351),
    .Q_N(_13263_),
    .Q(\atari2600.cpu.DIHOLD[5] ));
 sg13g2_dfrbp_1 _28884_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2443),
    .D(\atari2600.cpu.DIMUX[6] ),
    .Q_N(_13264_),
    .Q(\atari2600.cpu.DIHOLD[6] ));
 sg13g2_dfrbp_1 _28885_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2850),
    .D(net5273),
    .Q_N(_11017_),
    .Q(\atari2600.cpu.DIHOLD[7] ));
 sg13g2_dfrbp_1 _28886_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net2849),
    .D(_02455_),
    .Q_N(_11016_),
    .Q(\atari2600.cpu.load_reg ));
 sg13g2_dfrbp_1 _28887_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2848),
    .D(_02456_),
    .Q_N(_11015_),
    .Q(\atari2600.cpu.IRHOLD_valid ));
 sg13g2_dfrbp_1 _28888_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2846),
    .D(net6972),
    .Q_N(_11014_),
    .Q(\atari2600.cpu.IRHOLD[0] ));
 sg13g2_dfrbp_1 _28889_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2845),
    .D(net7033),
    .Q_N(_11013_),
    .Q(\atari2600.cpu.IRHOLD[1] ));
 sg13g2_dfrbp_1 _28890_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2844),
    .D(_02459_),
    .Q_N(_11012_),
    .Q(\atari2600.cpu.IRHOLD[2] ));
 sg13g2_dfrbp_1 _28891_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2843),
    .D(_02460_),
    .Q_N(_11011_),
    .Q(\atari2600.cpu.IRHOLD[3] ));
 sg13g2_dfrbp_1 _28892_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2842),
    .D(_02461_),
    .Q_N(_11010_),
    .Q(\atari2600.cpu.IRHOLD[4] ));
 sg13g2_dfrbp_1 _28893_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net2841),
    .D(_02462_),
    .Q_N(_11009_),
    .Q(\atari2600.cpu.IRHOLD[5] ));
 sg13g2_dfrbp_1 _28894_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2840),
    .D(_02463_),
    .Q_N(_11008_),
    .Q(\atari2600.cpu.IRHOLD[6] ));
 sg13g2_dfrbp_1 _28895_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net2839),
    .D(net3072),
    .Q_N(_11007_),
    .Q(\atari2600.cpu.IRHOLD[7] ));
 sg13g2_dfrbp_1 _28896_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2838),
    .D(_02465_),
    .Q_N(_00147_),
    .Q(\atari2600.cpu.D ));
 sg13g2_dfrbp_1 _28897_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2836),
    .D(net4148),
    .Q_N(_00098_),
    .Q(\atari2600.cpu.I ));
 sg13g2_dfrbp_1 _28898_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2834),
    .D(net3685),
    .Q_N(_00148_),
    .Q(\atari2600.cpu.V ));
 sg13g2_dfrbp_1 _28899_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2833),
    .D(net4090),
    .Q_N(_00149_),
    .Q(\atari2600.cpu.N ));
 sg13g2_dfrbp_1 _28900_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2832),
    .D(_02469_),
    .Q_N(_00096_),
    .Q(\atari2600.cpu.Z ));
 sg13g2_dfrbp_1 _28901_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net2831),
    .D(net7282),
    .Q_N(_00095_),
    .Q(\atari2600.cpu.C ));
 sg13g2_dfrbp_1 _28902_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2830),
    .D(_02471_),
    .Q_N(_11006_),
    .Q(\scanline[34][0] ));
 sg13g2_dfrbp_1 _28903_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2829),
    .D(_02472_),
    .Q_N(_11005_),
    .Q(\scanline[34][1] ));
 sg13g2_dfrbp_1 _28904_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2828),
    .D(_02473_),
    .Q_N(_11004_),
    .Q(\scanline[34][2] ));
 sg13g2_dfrbp_1 _28905_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2827),
    .D(_02474_),
    .Q_N(_11003_),
    .Q(\scanline[34][3] ));
 sg13g2_dfrbp_1 _28906_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2826),
    .D(_02475_),
    .Q_N(_11002_),
    .Q(\scanline[34][4] ));
 sg13g2_dfrbp_1 _28907_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2825),
    .D(_02476_),
    .Q_N(_11001_),
    .Q(\scanline[34][5] ));
 sg13g2_dfrbp_1 _28908_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2510),
    .D(_02477_),
    .Q_N(_13265_),
    .Q(\scanline[34][6] ));
 sg13g2_dfrbp_1 _28909_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net2824),
    .D(net6734),
    .Q_N(_00054_),
    .Q(\atari2600.cpu.adj_bcd ));
 sg13g2_dfrbp_1 _28910_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2823),
    .D(net7203),
    .Q_N(_11000_),
    .Q(\atari2600.cpu.backwards ));
 sg13g2_dfrbp_1 _28911_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2822),
    .D(_02479_),
    .Q_N(_10999_),
    .Q(\atari2600.cpu.ABL[0] ));
 sg13g2_dfrbp_1 _28912_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net2821),
    .D(_02480_),
    .Q_N(_10998_),
    .Q(\atari2600.cpu.ABL[1] ));
 sg13g2_dfrbp_1 _28913_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net2820),
    .D(net4292),
    .Q_N(_10997_),
    .Q(\atari2600.cpu.ABL[2] ));
 sg13g2_dfrbp_1 _28914_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net2819),
    .D(net3431),
    .Q_N(_10996_),
    .Q(\atari2600.cpu.ABL[3] ));
 sg13g2_dfrbp_1 _28915_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net2818),
    .D(_02483_),
    .Q_N(_10995_),
    .Q(\atari2600.cpu.ABL[4] ));
 sg13g2_dfrbp_1 _28916_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net2817),
    .D(_02484_),
    .Q_N(_10994_),
    .Q(\atari2600.cpu.ABL[5] ));
 sg13g2_dfrbp_1 _28917_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net2816),
    .D(_02485_),
    .Q_N(_10993_),
    .Q(\atari2600.cpu.ABL[6] ));
 sg13g2_dfrbp_1 _28918_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net2815),
    .D(_02486_),
    .Q_N(_10992_),
    .Q(\atari2600.cpu.ABL[7] ));
 sg13g2_dfrbp_1 _28919_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2814),
    .D(net6092),
    .Q_N(_10991_),
    .Q(\atari2600.cpu.ALU.AI7 ));
 sg13g2_dfrbp_1 _28920_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net2813),
    .D(_02488_),
    .Q_N(_10990_),
    .Q(\atari2600.cpu.ADD[0] ));
 sg13g2_dfrbp_1 _28921_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net2812),
    .D(_02489_),
    .Q_N(_00097_),
    .Q(\atari2600.cpu.ADD[1] ));
 sg13g2_dfrbp_1 _28922_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net2811),
    .D(_02490_),
    .Q_N(_00099_),
    .Q(\atari2600.cpu.ADD[2] ));
 sg13g2_dfrbp_1 _28923_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net2810),
    .D(_02491_),
    .Q_N(_00101_),
    .Q(\atari2600.cpu.ADD[3] ));
 sg13g2_dfrbp_1 _28924_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2809),
    .D(_02492_),
    .Q_N(_10989_),
    .Q(\atari2600.cpu.ADD[4] ));
 sg13g2_dfrbp_1 _28925_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2808),
    .D(_02493_),
    .Q_N(_00100_),
    .Q(\atari2600.cpu.ADD[5] ));
 sg13g2_dfrbp_1 _28926_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2807),
    .D(_02494_),
    .Q_N(_00103_),
    .Q(\atari2600.cpu.ADD[6] ));
 sg13g2_dfrbp_1 _28927_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net2806),
    .D(_02495_),
    .Q_N(_00104_),
    .Q(\atari2600.cpu.ADD[7] ));
 sg13g2_dfrbp_1 _28928_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net2805),
    .D(_02496_),
    .Q_N(_10988_),
    .Q(\atari2600.cpu.ALU.HC ));
 sg13g2_dfrbp_1 _28929_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net2804),
    .D(_02497_),
    .Q_N(_10987_),
    .Q(\atari2600.cpu.ALU.CO ));
 sg13g2_dfrbp_1 _28930_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2803),
    .D(net7124),
    .Q_N(_00065_),
    .Q(\atari2600.cpu.PC[0] ));
 sg13g2_dfrbp_1 _28931_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2802),
    .D(net7056),
    .Q_N(_00064_),
    .Q(\atari2600.cpu.PC[1] ));
 sg13g2_dfrbp_1 _28932_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net2801),
    .D(net6981),
    .Q_N(_00082_),
    .Q(\atari2600.cpu.PC[2] ));
 sg13g2_dfrbp_1 _28933_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net2800),
    .D(net7156),
    .Q_N(_00066_),
    .Q(\atari2600.cpu.PC[3] ));
 sg13g2_dfrbp_1 _28934_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net2799),
    .D(_02502_),
    .Q_N(_00067_),
    .Q(\atari2600.cpu.PC[4] ));
 sg13g2_dfrbp_1 _28935_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net2798),
    .D(net7133),
    .Q_N(_00068_),
    .Q(\atari2600.cpu.PC[5] ));
 sg13g2_dfrbp_1 _28936_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2797),
    .D(net7080),
    .Q_N(_00069_),
    .Q(\atari2600.cpu.PC[6] ));
 sg13g2_dfrbp_1 _28937_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2796),
    .D(net7069),
    .Q_N(_00070_),
    .Q(\atari2600.cpu.PC[7] ));
 sg13g2_dfrbp_1 _28938_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2795),
    .D(_02506_),
    .Q_N(_00071_),
    .Q(\atari2600.cpu.PC[8] ));
 sg13g2_dfrbp_1 _28939_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2794),
    .D(net4059),
    .Q_N(_00072_),
    .Q(\atari2600.cpu.PC[9] ));
 sg13g2_dfrbp_1 _28940_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net2793),
    .D(net7000),
    .Q_N(_00073_),
    .Q(\atari2600.cpu.PC[10] ));
 sg13g2_dfrbp_1 _28941_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net2792),
    .D(net7090),
    .Q_N(_00074_),
    .Q(\atari2600.cpu.PC[11] ));
 sg13g2_dfrbp_1 _28942_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net2791),
    .D(net6920),
    .Q_N(_00075_),
    .Q(\atari2600.cpu.PC[12] ));
 sg13g2_dfrbp_1 _28943_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2790),
    .D(net6582),
    .Q_N(_00076_),
    .Q(\atari2600.cpu.PC[13] ));
 sg13g2_dfrbp_1 _28944_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2789),
    .D(_02512_),
    .Q_N(_10986_),
    .Q(\atari2600.cpu.PC[14] ));
 sg13g2_dfrbp_1 _28945_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net2788),
    .D(net7084),
    .Q_N(_10985_),
    .Q(\atari2600.cpu.PC[15] ));
 sg13g2_dfrbp_1 _28946_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net2787),
    .D(_02514_),
    .Q_N(_10984_),
    .Q(\atari2600.ram[23][0] ));
 sg13g2_dfrbp_1 _28947_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2786),
    .D(_02515_),
    .Q_N(_10983_),
    .Q(\atari2600.ram[23][1] ));
 sg13g2_dfrbp_1 _28948_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net2785),
    .D(_02516_),
    .Q_N(_10982_),
    .Q(\atari2600.ram[23][2] ));
 sg13g2_dfrbp_1 _28949_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2784),
    .D(_02517_),
    .Q_N(_10981_),
    .Q(\atari2600.ram[23][3] ));
 sg13g2_dfrbp_1 _28950_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2783),
    .D(_02518_),
    .Q_N(_10980_),
    .Q(\atari2600.ram[23][4] ));
 sg13g2_dfrbp_1 _28951_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net2782),
    .D(_02519_),
    .Q_N(_10979_),
    .Q(\atari2600.ram[23][5] ));
 sg13g2_dfrbp_1 _28952_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net2781),
    .D(_02520_),
    .Q_N(_10978_),
    .Q(\atari2600.ram[23][6] ));
 sg13g2_dfrbp_1 _28953_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net2780),
    .D(_02521_),
    .Q_N(_10977_),
    .Q(\atari2600.ram[23][7] ));
 sg13g2_dfrbp_1 _28954_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2779),
    .D(_02522_),
    .Q_N(_10976_),
    .Q(\atari2600.ram[88][0] ));
 sg13g2_dfrbp_1 _28955_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net2778),
    .D(_02523_),
    .Q_N(_10975_),
    .Q(\atari2600.ram[88][1] ));
 sg13g2_dfrbp_1 _28956_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2777),
    .D(_02524_),
    .Q_N(_10974_),
    .Q(\atari2600.ram[88][2] ));
 sg13g2_dfrbp_1 _28957_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2776),
    .D(_02525_),
    .Q_N(_10973_),
    .Q(\atari2600.ram[88][3] ));
 sg13g2_dfrbp_1 _28958_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2775),
    .D(_02526_),
    .Q_N(_10972_),
    .Q(\atari2600.ram[88][4] ));
 sg13g2_dfrbp_1 _28959_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2774),
    .D(_02527_),
    .Q_N(_10971_),
    .Q(\atari2600.ram[88][5] ));
 sg13g2_dfrbp_1 _28960_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2773),
    .D(_02528_),
    .Q_N(_10970_),
    .Q(\atari2600.ram[88][6] ));
 sg13g2_dfrbp_1 _28961_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2772),
    .D(_02529_),
    .Q_N(_10969_),
    .Q(\atari2600.ram[88][7] ));
 sg13g2_dfrbp_1 _28962_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2771),
    .D(_02530_),
    .Q_N(_10968_),
    .Q(\scanline[33][0] ));
 sg13g2_dfrbp_1 _28963_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2770),
    .D(_02531_),
    .Q_N(_10967_),
    .Q(\scanline[33][1] ));
 sg13g2_dfrbp_1 _28964_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2769),
    .D(_02532_),
    .Q_N(_10966_),
    .Q(\scanline[33][2] ));
 sg13g2_dfrbp_1 _28965_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net2768),
    .D(_02533_),
    .Q_N(_10965_),
    .Q(\scanline[33][3] ));
 sg13g2_dfrbp_1 _28966_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2767),
    .D(_02534_),
    .Q_N(_10964_),
    .Q(\scanline[33][4] ));
 sg13g2_dfrbp_1 _28967_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2766),
    .D(_02535_),
    .Q_N(_10963_),
    .Q(\scanline[33][5] ));
 sg13g2_dfrbp_1 _28968_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net2765),
    .D(_02536_),
    .Q_N(_10962_),
    .Q(\scanline[33][6] ));
 sg13g2_dfrbp_1 _28969_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2764),
    .D(_02537_),
    .Q_N(_10961_),
    .Q(\atari2600.ram[43][0] ));
 sg13g2_dfrbp_1 _28970_ (.CLK(clknet_leaf_349_clk),
    .RESET_B(net2763),
    .D(_02538_),
    .Q_N(_10960_),
    .Q(\atari2600.ram[43][1] ));
 sg13g2_dfrbp_1 _28971_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2762),
    .D(_02539_),
    .Q_N(_10959_),
    .Q(\atari2600.ram[43][2] ));
 sg13g2_dfrbp_1 _28972_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net2761),
    .D(_02540_),
    .Q_N(_10958_),
    .Q(\atari2600.ram[43][3] ));
 sg13g2_dfrbp_1 _28973_ (.CLK(clknet_leaf_350_clk),
    .RESET_B(net2760),
    .D(_02541_),
    .Q_N(_10957_),
    .Q(\atari2600.ram[43][4] ));
 sg13g2_dfrbp_1 _28974_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net2759),
    .D(_02542_),
    .Q_N(_10956_),
    .Q(\atari2600.ram[43][5] ));
 sg13g2_dfrbp_1 _28975_ (.CLK(clknet_leaf_349_clk),
    .RESET_B(net2758),
    .D(_02543_),
    .Q_N(_10955_),
    .Q(\atari2600.ram[43][6] ));
 sg13g2_dfrbp_1 _28976_ (.CLK(clknet_leaf_349_clk),
    .RESET_B(net2757),
    .D(_02544_),
    .Q_N(_10954_),
    .Q(\atari2600.ram[43][7] ));
 sg13g2_dfrbp_1 _28977_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net2756),
    .D(_02545_),
    .Q_N(_10953_),
    .Q(\atari2600.ram[42][0] ));
 sg13g2_dfrbp_1 _28978_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net2755),
    .D(_02546_),
    .Q_N(_10952_),
    .Q(\atari2600.ram[42][1] ));
 sg13g2_dfrbp_1 _28979_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net2754),
    .D(_02547_),
    .Q_N(_10951_),
    .Q(\atari2600.ram[42][2] ));
 sg13g2_dfrbp_1 _28980_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net2753),
    .D(_02548_),
    .Q_N(_10950_),
    .Q(\atari2600.ram[42][3] ));
 sg13g2_dfrbp_1 _28981_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2752),
    .D(_02549_),
    .Q_N(_10949_),
    .Q(\atari2600.ram[42][4] ));
 sg13g2_dfrbp_1 _28982_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2751),
    .D(_02550_),
    .Q_N(_10948_),
    .Q(\atari2600.ram[42][5] ));
 sg13g2_dfrbp_1 _28983_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2750),
    .D(_02551_),
    .Q_N(_10947_),
    .Q(\atari2600.ram[42][6] ));
 sg13g2_dfrbp_1 _28984_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net2749),
    .D(_02552_),
    .Q_N(_10946_),
    .Q(\atari2600.ram[42][7] ));
 sg13g2_dfrbp_1 _28985_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2748),
    .D(_02553_),
    .Q_N(_10945_),
    .Q(\atari2600.ram[73][0] ));
 sg13g2_dfrbp_1 _28986_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2747),
    .D(_02554_),
    .Q_N(_10944_),
    .Q(\atari2600.ram[73][1] ));
 sg13g2_dfrbp_1 _28987_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net2746),
    .D(_02555_),
    .Q_N(_10943_),
    .Q(\atari2600.ram[73][2] ));
 sg13g2_dfrbp_1 _28988_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2745),
    .D(_02556_),
    .Q_N(_10942_),
    .Q(\atari2600.ram[73][3] ));
 sg13g2_dfrbp_1 _28989_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2744),
    .D(_02557_),
    .Q_N(_10941_),
    .Q(\atari2600.ram[73][4] ));
 sg13g2_dfrbp_1 _28990_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2743),
    .D(_02558_),
    .Q_N(_10940_),
    .Q(\atari2600.ram[73][5] ));
 sg13g2_dfrbp_1 _28991_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2742),
    .D(_02559_),
    .Q_N(_10939_),
    .Q(\atari2600.ram[73][6] ));
 sg13g2_dfrbp_1 _28992_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2741),
    .D(_02560_),
    .Q_N(_10938_),
    .Q(\atari2600.ram[73][7] ));
 sg13g2_dfrbp_1 _28993_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2740),
    .D(_02561_),
    .Q_N(_10937_),
    .Q(\atari2600.clk_counter[0] ));
 sg13g2_dfrbp_1 _28994_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2738),
    .D(_02562_),
    .Q_N(_10936_),
    .Q(\atari2600.clk_counter[1] ));
 sg13g2_dfrbp_1 _28995_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2736),
    .D(_02563_),
    .Q_N(_10935_),
    .Q(\atari2600.clk_counter[2] ));
 sg13g2_dfrbp_1 _28996_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2734),
    .D(_02564_),
    .Q_N(_10934_),
    .Q(\atari2600.clk_counter[3] ));
 sg13g2_dfrbp_1 _28997_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2732),
    .D(_02565_),
    .Q_N(_10933_),
    .Q(\atari2600.clk_counter[4] ));
 sg13g2_dfrbp_1 _28998_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2730),
    .D(_02566_),
    .Q_N(_10932_),
    .Q(\atari2600.clk_counter[5] ));
 sg13g2_dfrbp_1 _28999_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2728),
    .D(_02567_),
    .Q_N(_10931_),
    .Q(\atari2600.clk_counter[6] ));
 sg13g2_dfrbp_1 _29000_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2726),
    .D(_02568_),
    .Q_N(_10930_),
    .Q(\atari2600.clk_counter[7] ));
 sg13g2_dfrbp_1 _29001_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2724),
    .D(_02569_),
    .Q_N(_00142_),
    .Q(\atari2600.clk_counter[8] ));
 sg13g2_dfrbp_1 _29002_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2722),
    .D(_02570_),
    .Q_N(_10929_),
    .Q(\atari2600.ram[6][0] ));
 sg13g2_dfrbp_1 _29003_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2721),
    .D(_02571_),
    .Q_N(_10928_),
    .Q(\atari2600.ram[6][1] ));
 sg13g2_dfrbp_1 _29004_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2720),
    .D(_02572_),
    .Q_N(_10927_),
    .Q(\atari2600.ram[6][2] ));
 sg13g2_dfrbp_1 _29005_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2719),
    .D(_02573_),
    .Q_N(_10926_),
    .Q(\atari2600.ram[6][3] ));
 sg13g2_dfrbp_1 _29006_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2718),
    .D(_02574_),
    .Q_N(_10925_),
    .Q(\atari2600.ram[6][4] ));
 sg13g2_dfrbp_1 _29007_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2717),
    .D(_02575_),
    .Q_N(_10924_),
    .Q(\atari2600.ram[6][5] ));
 sg13g2_dfrbp_1 _29008_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2716),
    .D(_02576_),
    .Q_N(_10923_),
    .Q(\atari2600.ram[6][6] ));
 sg13g2_dfrbp_1 _29009_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2715),
    .D(_02577_),
    .Q_N(_10922_),
    .Q(\atari2600.ram[6][7] ));
 sg13g2_dfrbp_1 _29010_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net2714),
    .D(_02578_),
    .Q_N(_10921_),
    .Q(\atari2600.ram[86][0] ));
 sg13g2_dfrbp_1 _29011_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2713),
    .D(_02579_),
    .Q_N(_10920_),
    .Q(\atari2600.ram[86][1] ));
 sg13g2_dfrbp_1 _29012_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2712),
    .D(_02580_),
    .Q_N(_10919_),
    .Q(\atari2600.ram[86][2] ));
 sg13g2_dfrbp_1 _29013_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2711),
    .D(_02581_),
    .Q_N(_10918_),
    .Q(\atari2600.ram[86][3] ));
 sg13g2_dfrbp_1 _29014_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net2710),
    .D(_02582_),
    .Q_N(_10917_),
    .Q(\atari2600.ram[86][4] ));
 sg13g2_dfrbp_1 _29015_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net2709),
    .D(_02583_),
    .Q_N(_10916_),
    .Q(\atari2600.ram[86][5] ));
 sg13g2_dfrbp_1 _29016_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2708),
    .D(_02584_),
    .Q_N(_10915_),
    .Q(\atari2600.ram[86][6] ));
 sg13g2_dfrbp_1 _29017_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2519),
    .D(_02585_),
    .Q_N(_13266_),
    .Q(\atari2600.ram[86][7] ));
 sg13g2_dfrbp_1 _29018_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net2707),
    .D(_00013_),
    .Q_N(_10914_),
    .Q(\hvsync_gen.vga.vsync ));
 sg13g2_dfrbp_1 _29019_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2706),
    .D(_02586_),
    .Q_N(_00170_),
    .Q(\hvsync_gen.vga.vpos[0] ));
 sg13g2_dfrbp_1 _29020_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2704),
    .D(_02587_),
    .Q_N(_10913_),
    .Q(\hvsync_gen.vga.vpos[1] ));
 sg13g2_dfrbp_1 _29021_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2702),
    .D(_02588_),
    .Q_N(_10912_),
    .Q(\hvsync_gen.vga.vpos[2] ));
 sg13g2_dfrbp_1 _29022_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2700),
    .D(_02589_),
    .Q_N(_10911_),
    .Q(\hvsync_gen.vga.vpos[3] ));
 sg13g2_dfrbp_1 _29023_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2698),
    .D(_02590_),
    .Q_N(_10910_),
    .Q(\hvsync_gen.vga.vpos[4] ));
 sg13g2_dfrbp_1 _29024_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2696),
    .D(_02591_),
    .Q_N(_10909_),
    .Q(\hvsync_gen.vga.vpos[5] ));
 sg13g2_dfrbp_1 _29025_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2694),
    .D(_02592_),
    .Q_N(_10908_),
    .Q(\hvsync_gen.vga.vpos[6] ));
 sg13g2_dfrbp_1 _29026_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2692),
    .D(_02593_),
    .Q_N(_10907_),
    .Q(\hvsync_gen.vga.vpos[7] ));
 sg13g2_dfrbp_1 _29027_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2690),
    .D(_02594_),
    .Q_N(_10906_),
    .Q(\hvsync_gen.vga.vpos[8] ));
 sg13g2_dfrbp_1 _29028_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net234),
    .D(net7143),
    .Q_N(_13267_),
    .Q(\hvsync_gen.vga.vpos[9] ));
 sg13g2_dfrbp_1 _29029_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net2688),
    .D(_00047_),
    .Q_N(_10905_),
    .Q(hsync));
 sg13g2_dfrbp_1 _29030_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net2686),
    .D(net7231),
    .Q_N(_10904_),
    .Q(\flash_rom.data_ready ));
 sg13g2_dfrbp_1 _29031_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2685),
    .D(_02597_),
    .Q_N(_10903_),
    .Q(\atari2600.ram[31][0] ));
 sg13g2_dfrbp_1 _29032_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2684),
    .D(_02598_),
    .Q_N(_10902_),
    .Q(\atari2600.ram[31][1] ));
 sg13g2_dfrbp_1 _29033_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2683),
    .D(_02599_),
    .Q_N(_10901_),
    .Q(\atari2600.ram[31][2] ));
 sg13g2_dfrbp_1 _29034_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2682),
    .D(_02600_),
    .Q_N(_10900_),
    .Q(\atari2600.ram[31][3] ));
 sg13g2_dfrbp_1 _29035_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2681),
    .D(_02601_),
    .Q_N(_10899_),
    .Q(\atari2600.ram[31][4] ));
 sg13g2_dfrbp_1 _29036_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net2680),
    .D(_02602_),
    .Q_N(_10898_),
    .Q(\atari2600.ram[31][5] ));
 sg13g2_dfrbp_1 _29037_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net2679),
    .D(_02603_),
    .Q_N(_10897_),
    .Q(\atari2600.ram[31][6] ));
 sg13g2_dfrbp_1 _29038_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net2678),
    .D(_02604_),
    .Q_N(_10896_),
    .Q(\atari2600.ram[31][7] ));
 sg13g2_dfrbp_1 _29039_ (.CLK(clknet_leaf_356_clk),
    .RESET_B(net2677),
    .D(_02605_),
    .Q_N(_10895_),
    .Q(\atari2600.ram[32][0] ));
 sg13g2_dfrbp_1 _29040_ (.CLK(clknet_leaf_355_clk),
    .RESET_B(net2676),
    .D(_02606_),
    .Q_N(_10894_),
    .Q(\atari2600.ram[32][1] ));
 sg13g2_dfrbp_1 _29041_ (.CLK(clknet_leaf_356_clk),
    .RESET_B(net2675),
    .D(_02607_),
    .Q_N(_10893_),
    .Q(\atari2600.ram[32][2] ));
 sg13g2_dfrbp_1 _29042_ (.CLK(clknet_leaf_356_clk),
    .RESET_B(net2674),
    .D(_02608_),
    .Q_N(_10892_),
    .Q(\atari2600.ram[32][3] ));
 sg13g2_dfrbp_1 _29043_ (.CLK(clknet_leaf_353_clk),
    .RESET_B(net2673),
    .D(_02609_),
    .Q_N(_10891_),
    .Q(\atari2600.ram[32][4] ));
 sg13g2_dfrbp_1 _29044_ (.CLK(clknet_leaf_355_clk),
    .RESET_B(net2672),
    .D(_02610_),
    .Q_N(_10890_),
    .Q(\atari2600.ram[32][5] ));
 sg13g2_dfrbp_1 _29045_ (.CLK(clknet_leaf_355_clk),
    .RESET_B(net2671),
    .D(_02611_),
    .Q_N(_10889_),
    .Q(\atari2600.ram[32][6] ));
 sg13g2_dfrbp_1 _29046_ (.CLK(clknet_leaf_355_clk),
    .RESET_B(net2670),
    .D(_02612_),
    .Q_N(_10888_),
    .Q(\atari2600.ram[32][7] ));
 sg13g2_dfrbp_1 _29047_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2669),
    .D(_02613_),
    .Q_N(_10887_),
    .Q(\atari2600.ram[22][0] ));
 sg13g2_dfrbp_1 _29048_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2668),
    .D(_02614_),
    .Q_N(_10886_),
    .Q(\atari2600.ram[22][1] ));
 sg13g2_dfrbp_1 _29049_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net2667),
    .D(_02615_),
    .Q_N(_10885_),
    .Q(\atari2600.ram[22][2] ));
 sg13g2_dfrbp_1 _29050_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net2666),
    .D(_02616_),
    .Q_N(_10884_),
    .Q(\atari2600.ram[22][3] ));
 sg13g2_dfrbp_1 _29051_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2665),
    .D(_02617_),
    .Q_N(_10883_),
    .Q(\atari2600.ram[22][4] ));
 sg13g2_dfrbp_1 _29052_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2664),
    .D(_02618_),
    .Q_N(_10882_),
    .Q(\atari2600.ram[22][5] ));
 sg13g2_dfrbp_1 _29053_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2663),
    .D(_02619_),
    .Q_N(_10881_),
    .Q(\atari2600.ram[22][6] ));
 sg13g2_dfrbp_1 _29054_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net2662),
    .D(_02620_),
    .Q_N(_10880_),
    .Q(\atari2600.ram[22][7] ));
 sg13g2_dfrbp_1 _29055_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2661),
    .D(_02621_),
    .Q_N(_10879_),
    .Q(\atari2600.ram[26][0] ));
 sg13g2_dfrbp_1 _29056_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2660),
    .D(_02622_),
    .Q_N(_10878_),
    .Q(\atari2600.ram[26][1] ));
 sg13g2_dfrbp_1 _29057_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2659),
    .D(_02623_),
    .Q_N(_10877_),
    .Q(\atari2600.ram[26][2] ));
 sg13g2_dfrbp_1 _29058_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2658),
    .D(_02624_),
    .Q_N(_10876_),
    .Q(\atari2600.ram[26][3] ));
 sg13g2_dfrbp_1 _29059_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2657),
    .D(_02625_),
    .Q_N(_10875_),
    .Q(\atari2600.ram[26][4] ));
 sg13g2_dfrbp_1 _29060_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net2656),
    .D(_02626_),
    .Q_N(_10874_),
    .Q(\atari2600.ram[26][5] ));
 sg13g2_dfrbp_1 _29061_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2655),
    .D(_02627_),
    .Q_N(_10873_),
    .Q(\atari2600.ram[26][6] ));
 sg13g2_dfrbp_1 _29062_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2654),
    .D(_02628_),
    .Q_N(_10872_),
    .Q(\atari2600.ram[26][7] ));
 sg13g2_dfrbp_1 _29063_ (.CLK(clknet_leaf_352_clk),
    .RESET_B(net2653),
    .D(_02629_),
    .Q_N(_10871_),
    .Q(\atari2600.ram[33][0] ));
 sg13g2_dfrbp_1 _29064_ (.CLK(clknet_leaf_353_clk),
    .RESET_B(net2652),
    .D(_02630_),
    .Q_N(_10870_),
    .Q(\atari2600.ram[33][1] ));
 sg13g2_dfrbp_1 _29065_ (.CLK(clknet_leaf_351_clk),
    .RESET_B(net2651),
    .D(_02631_),
    .Q_N(_10869_),
    .Q(\atari2600.ram[33][2] ));
 sg13g2_dfrbp_1 _29066_ (.CLK(clknet_leaf_357_clk),
    .RESET_B(net2650),
    .D(_02632_),
    .Q_N(_10868_),
    .Q(\atari2600.ram[33][3] ));
 sg13g2_dfrbp_1 _29067_ (.CLK(clknet_leaf_353_clk),
    .RESET_B(net2649),
    .D(_02633_),
    .Q_N(_10867_),
    .Q(\atari2600.ram[33][4] ));
 sg13g2_dfrbp_1 _29068_ (.CLK(clknet_leaf_357_clk),
    .RESET_B(net2648),
    .D(_02634_),
    .Q_N(_10866_),
    .Q(\atari2600.ram[33][5] ));
 sg13g2_dfrbp_1 _29069_ (.CLK(clknet_leaf_353_clk),
    .RESET_B(net2647),
    .D(_02635_),
    .Q_N(_10865_),
    .Q(\atari2600.ram[33][6] ));
 sg13g2_dfrbp_1 _29070_ (.CLK(clknet_leaf_352_clk),
    .RESET_B(net2646),
    .D(_02636_),
    .Q_N(_10864_),
    .Q(\atari2600.ram[33][7] ));
 sg13g2_dfrbp_1 _29071_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2645),
    .D(_02637_),
    .Q_N(_10863_),
    .Q(\atari2600.ram[25][0] ));
 sg13g2_dfrbp_1 _29072_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net2644),
    .D(_02638_),
    .Q_N(_10862_),
    .Q(\atari2600.ram[25][1] ));
 sg13g2_dfrbp_1 _29073_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2643),
    .D(_02639_),
    .Q_N(_10861_),
    .Q(\atari2600.ram[25][2] ));
 sg13g2_dfrbp_1 _29074_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2642),
    .D(_02640_),
    .Q_N(_10860_),
    .Q(\atari2600.ram[25][3] ));
 sg13g2_dfrbp_1 _29075_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2641),
    .D(_02641_),
    .Q_N(_10859_),
    .Q(\atari2600.ram[25][4] ));
 sg13g2_dfrbp_1 _29076_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2640),
    .D(_02642_),
    .Q_N(_10858_),
    .Q(\atari2600.ram[25][5] ));
 sg13g2_dfrbp_1 _29077_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net2639),
    .D(_02643_),
    .Q_N(_10857_),
    .Q(\atari2600.ram[25][6] ));
 sg13g2_dfrbp_1 _29078_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2638),
    .D(_02644_),
    .Q_N(_10856_),
    .Q(\atari2600.ram[25][7] ));
 sg13g2_dfrbp_1 _29079_ (.CLK(clknet_leaf_355_clk),
    .RESET_B(net2637),
    .D(_02645_),
    .Q_N(_10855_),
    .Q(\atari2600.ram[35][0] ));
 sg13g2_dfrbp_1 _29080_ (.CLK(clknet_leaf_354_clk),
    .RESET_B(net2636),
    .D(_02646_),
    .Q_N(_10854_),
    .Q(\atari2600.ram[35][1] ));
 sg13g2_dfrbp_1 _29081_ (.CLK(clknet_leaf_356_clk),
    .RESET_B(net2602),
    .D(_02647_),
    .Q_N(_10853_),
    .Q(\atari2600.ram[35][2] ));
 sg13g2_dfrbp_1 _29082_ (.CLK(clknet_leaf_356_clk),
    .RESET_B(net2600),
    .D(_02648_),
    .Q_N(_10852_),
    .Q(\atari2600.ram[35][3] ));
 sg13g2_dfrbp_1 _29083_ (.CLK(clknet_leaf_354_clk),
    .RESET_B(net2598),
    .D(_02649_),
    .Q_N(_10851_),
    .Q(\atari2600.ram[35][4] ));
 sg13g2_dfrbp_1 _29084_ (.CLK(clknet_leaf_355_clk),
    .RESET_B(net2596),
    .D(_02650_),
    .Q_N(_10850_),
    .Q(\atari2600.ram[35][5] ));
 sg13g2_dfrbp_1 _29085_ (.CLK(clknet_leaf_355_clk),
    .RESET_B(net2594),
    .D(_02651_),
    .Q_N(_10849_),
    .Q(\atari2600.ram[35][6] ));
 sg13g2_dfrbp_1 _29086_ (.CLK(clknet_leaf_355_clk),
    .RESET_B(net2592),
    .D(_02652_),
    .Q_N(_10848_),
    .Q(\atari2600.ram[35][7] ));
 sg13g2_dfrbp_1 _29087_ (.CLK(clknet_leaf_362_clk),
    .RESET_B(net2590),
    .D(_02653_),
    .Q_N(_00091_),
    .Q(\atari2600.cpu.AXYS[2][0] ));
 sg13g2_dfrbp_1 _29088_ (.CLK(clknet_leaf_361_clk),
    .RESET_B(net1634),
    .D(_02654_),
    .Q_N(_00085_),
    .Q(\atari2600.cpu.AXYS[2][1] ));
 sg13g2_dfrbp_1 _29089_ (.CLK(clknet_leaf_361_clk),
    .RESET_B(net1632),
    .D(_02655_),
    .Q_N(_10847_),
    .Q(\atari2600.cpu.AXYS[2][2] ));
 sg13g2_dfrbp_1 _29090_ (.CLK(clknet_leaf_361_clk),
    .RESET_B(net1553),
    .D(_02656_),
    .Q_N(_10846_),
    .Q(\atari2600.cpu.AXYS[2][3] ));
 sg13g2_dfrbp_1 _29091_ (.CLK(clknet_leaf_359_clk),
    .RESET_B(net1551),
    .D(_02657_),
    .Q_N(_10845_),
    .Q(\atari2600.cpu.AXYS[2][4] ));
 sg13g2_dfrbp_1 _29092_ (.CLK(clknet_leaf_359_clk),
    .RESET_B(net1549),
    .D(_02658_),
    .Q_N(_10844_),
    .Q(\atari2600.cpu.AXYS[2][5] ));
 sg13g2_dfrbp_1 _29093_ (.CLK(clknet_leaf_360_clk),
    .RESET_B(net1540),
    .D(_02659_),
    .Q_N(_10843_),
    .Q(\atari2600.cpu.AXYS[2][6] ));
 sg13g2_dfrbp_1 _29094_ (.CLK(clknet_leaf_360_clk),
    .RESET_B(net1538),
    .D(_02660_),
    .Q_N(_10842_),
    .Q(\atari2600.cpu.AXYS[2][7] ));
 sg13g2_dfrbp_1 _29095_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1536),
    .D(_02661_),
    .Q_N(_10841_),
    .Q(\atari2600.ram[4][0] ));
 sg13g2_dfrbp_1 _29096_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1534),
    .D(_02662_),
    .Q_N(_10840_),
    .Q(\atari2600.ram[4][1] ));
 sg13g2_dfrbp_1 _29097_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1532),
    .D(_02663_),
    .Q_N(_10839_),
    .Q(\atari2600.ram[4][2] ));
 sg13g2_dfrbp_1 _29098_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1530),
    .D(_02664_),
    .Q_N(_10838_),
    .Q(\atari2600.ram[4][3] ));
 sg13g2_dfrbp_1 _29099_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1528),
    .D(_02665_),
    .Q_N(_10837_),
    .Q(\atari2600.ram[4][4] ));
 sg13g2_dfrbp_1 _29100_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1526),
    .D(_02666_),
    .Q_N(_10836_),
    .Q(\atari2600.ram[4][5] ));
 sg13g2_dfrbp_1 _29101_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1524),
    .D(_02667_),
    .Q_N(_10835_),
    .Q(\atari2600.ram[4][6] ));
 sg13g2_dfrbp_1 _29102_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1522),
    .D(_02668_),
    .Q_N(_10834_),
    .Q(\atari2600.ram[4][7] ));
 sg13g2_dfrbp_1 _29103_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1520),
    .D(_02669_),
    .Q_N(_10833_),
    .Q(\atari2600.ram[50][0] ));
 sg13g2_dfrbp_1 _29104_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1518),
    .D(_02670_),
    .Q_N(_10832_),
    .Q(\atari2600.ram[50][1] ));
 sg13g2_dfrbp_1 _29105_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1472),
    .D(_02671_),
    .Q_N(_10831_),
    .Q(\atari2600.ram[50][2] ));
 sg13g2_dfrbp_1 _29106_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net976),
    .D(_02672_),
    .Q_N(_10830_),
    .Q(\atari2600.ram[50][3] ));
 sg13g2_dfrbp_1 _29107_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net974),
    .D(_02673_),
    .Q_N(_10829_),
    .Q(\atari2600.ram[50][4] ));
 sg13g2_dfrbp_1 _29108_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net972),
    .D(_02674_),
    .Q_N(_10828_),
    .Q(\atari2600.ram[50][5] ));
 sg13g2_dfrbp_1 _29109_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net970),
    .D(_02675_),
    .Q_N(_10827_),
    .Q(\atari2600.ram[50][6] ));
 sg13g2_dfrbp_1 _29110_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net968),
    .D(_02676_),
    .Q_N(_10826_),
    .Q(\atari2600.ram[50][7] ));
 sg13g2_dfrbp_1 _29111_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net966),
    .D(_02677_),
    .Q_N(_10825_),
    .Q(\atari2600.ram[51][0] ));
 sg13g2_dfrbp_1 _29112_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net964),
    .D(_02678_),
    .Q_N(_10824_),
    .Q(\atari2600.ram[51][1] ));
 sg13g2_dfrbp_1 _29113_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net962),
    .D(_02679_),
    .Q_N(_10823_),
    .Q(\atari2600.ram[51][2] ));
 sg13g2_dfrbp_1 _29114_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net960),
    .D(_02680_),
    .Q_N(_10822_),
    .Q(\atari2600.ram[51][3] ));
 sg13g2_dfrbp_1 _29115_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net950),
    .D(_02681_),
    .Q_N(_10821_),
    .Q(\atari2600.ram[51][4] ));
 sg13g2_dfrbp_1 _29116_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net948),
    .D(_02682_),
    .Q_N(_10820_),
    .Q(\atari2600.ram[51][5] ));
 sg13g2_dfrbp_1 _29117_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net946),
    .D(_02683_),
    .Q_N(_10819_),
    .Q(\atari2600.ram[51][6] ));
 sg13g2_dfrbp_1 _29118_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net944),
    .D(_02684_),
    .Q_N(_10818_),
    .Q(\atari2600.ram[51][7] ));
 sg13g2_dfrbp_1 _29119_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net942),
    .D(_02685_),
    .Q_N(_10817_),
    .Q(\atari2600.ram[52][0] ));
 sg13g2_dfrbp_1 _29120_ (.CLK(clknet_leaf_340_clk),
    .RESET_B(net940),
    .D(_02686_),
    .Q_N(_10816_),
    .Q(\atari2600.ram[52][1] ));
 sg13g2_dfrbp_1 _29121_ (.CLK(clknet_leaf_340_clk),
    .RESET_B(net938),
    .D(_02687_),
    .Q_N(_10815_),
    .Q(\atari2600.ram[52][2] ));
 sg13g2_dfrbp_1 _29122_ (.CLK(clknet_leaf_345_clk),
    .RESET_B(net936),
    .D(_02688_),
    .Q_N(_10814_),
    .Q(\atari2600.ram[52][3] ));
 sg13g2_dfrbp_1 _29123_ (.CLK(clknet_leaf_346_clk),
    .RESET_B(net934),
    .D(_02689_),
    .Q_N(_10813_),
    .Q(\atari2600.ram[52][4] ));
 sg13g2_dfrbp_1 _29124_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net932),
    .D(_02690_),
    .Q_N(_10812_),
    .Q(\atari2600.ram[52][5] ));
 sg13g2_dfrbp_1 _29125_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net930),
    .D(_02691_),
    .Q_N(_10811_),
    .Q(\atari2600.ram[52][6] ));
 sg13g2_dfrbp_1 _29126_ (.CLK(clknet_leaf_340_clk),
    .RESET_B(net928),
    .D(_02692_),
    .Q_N(_10810_),
    .Q(\atari2600.ram[52][7] ));
 sg13g2_dfrbp_1 _29127_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net926),
    .D(_02693_),
    .Q_N(_10809_),
    .Q(\atari2600.ram[53][0] ));
 sg13g2_dfrbp_1 _29128_ (.CLK(clknet_leaf_340_clk),
    .RESET_B(net924),
    .D(_02694_),
    .Q_N(_10808_),
    .Q(\atari2600.ram[53][1] ));
 sg13g2_dfrbp_1 _29129_ (.CLK(clknet_leaf_340_clk),
    .RESET_B(net922),
    .D(_02695_),
    .Q_N(_10807_),
    .Q(\atari2600.ram[53][2] ));
 sg13g2_dfrbp_1 _29130_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net920),
    .D(_02696_),
    .Q_N(_10806_),
    .Q(\atari2600.ram[53][3] ));
 sg13g2_dfrbp_1 _29131_ (.CLK(clknet_leaf_346_clk),
    .RESET_B(net918),
    .D(_02697_),
    .Q_N(_10805_),
    .Q(\atari2600.ram[53][4] ));
 sg13g2_dfrbp_1 _29132_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net916),
    .D(_02698_),
    .Q_N(_10804_),
    .Q(\atari2600.ram[53][5] ));
 sg13g2_dfrbp_1 _29133_ (.CLK(clknet_leaf_347_clk),
    .RESET_B(net914),
    .D(_02699_),
    .Q_N(_10803_),
    .Q(\atari2600.ram[53][6] ));
 sg13g2_dfrbp_1 _29134_ (.CLK(clknet_leaf_344_clk),
    .RESET_B(net912),
    .D(_02700_),
    .Q_N(_10802_),
    .Q(\atari2600.ram[53][7] ));
 sg13g2_dfrbp_1 _29135_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net910),
    .D(_02701_),
    .Q_N(_10801_),
    .Q(\atari2600.ram[54][0] ));
 sg13g2_dfrbp_1 _29136_ (.CLK(clknet_leaf_343_clk),
    .RESET_B(net908),
    .D(_02702_),
    .Q_N(_10800_),
    .Q(\atari2600.ram[54][1] ));
 sg13g2_dfrbp_1 _29137_ (.CLK(clknet_leaf_343_clk),
    .RESET_B(net906),
    .D(_02703_),
    .Q_N(_10799_),
    .Q(\atari2600.ram[54][2] ));
 sg13g2_dfrbp_1 _29138_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net904),
    .D(_02704_),
    .Q_N(_10798_),
    .Q(\atari2600.ram[54][3] ));
 sg13g2_dfrbp_1 _29139_ (.CLK(clknet_leaf_345_clk),
    .RESET_B(net863),
    .D(_02705_),
    .Q_N(_10797_),
    .Q(\atari2600.ram[54][4] ));
 sg13g2_dfrbp_1 _29140_ (.CLK(clknet_leaf_321_clk),
    .RESET_B(net861),
    .D(_02706_),
    .Q_N(_10796_),
    .Q(\atari2600.ram[54][5] ));
 sg13g2_dfrbp_1 _29141_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net859),
    .D(_02707_),
    .Q_N(_10795_),
    .Q(\atari2600.ram[54][6] ));
 sg13g2_dfrbp_1 _29142_ (.CLK(clknet_leaf_344_clk),
    .RESET_B(net857),
    .D(_02708_),
    .Q_N(_10794_),
    .Q(\atari2600.ram[54][7] ));
 sg13g2_dfrbp_1 _29143_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net855),
    .D(_02709_),
    .Q_N(_10793_),
    .Q(\atari2600.ram[55][0] ));
 sg13g2_dfrbp_1 _29144_ (.CLK(clknet_leaf_342_clk),
    .RESET_B(net853),
    .D(_02710_),
    .Q_N(_10792_),
    .Q(\atari2600.ram[55][1] ));
 sg13g2_dfrbp_1 _29145_ (.CLK(clknet_leaf_344_clk),
    .RESET_B(net851),
    .D(_02711_),
    .Q_N(_10791_),
    .Q(\atari2600.ram[55][2] ));
 sg13g2_dfrbp_1 _29146_ (.CLK(clknet_leaf_347_clk),
    .RESET_B(net849),
    .D(_02712_),
    .Q_N(_10790_),
    .Q(\atari2600.ram[55][3] ));
 sg13g2_dfrbp_1 _29147_ (.CLK(clknet_leaf_347_clk),
    .RESET_B(net847),
    .D(_02713_),
    .Q_N(_10789_),
    .Q(\atari2600.ram[55][4] ));
 sg13g2_dfrbp_1 _29148_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net845),
    .D(_02714_),
    .Q_N(_10788_),
    .Q(\atari2600.ram[55][5] ));
 sg13g2_dfrbp_1 _29149_ (.CLK(clknet_leaf_319_clk),
    .RESET_B(net843),
    .D(_02715_),
    .Q_N(_10787_),
    .Q(\atari2600.ram[55][6] ));
 sg13g2_dfrbp_1 _29150_ (.CLK(clknet_leaf_338_clk),
    .RESET_B(net841),
    .D(_02716_),
    .Q_N(_10786_),
    .Q(\atari2600.ram[55][7] ));
 sg13g2_dfrbp_1 _29151_ (.CLK(clknet_leaf_340_clk),
    .RESET_B(net839),
    .D(_02717_),
    .Q_N(_10785_),
    .Q(\atari2600.ram[56][0] ));
 sg13g2_dfrbp_1 _29152_ (.CLK(clknet_leaf_354_clk),
    .RESET_B(net837),
    .D(_02718_),
    .Q_N(_10784_),
    .Q(\atari2600.ram[56][1] ));
 sg13g2_dfrbp_1 _29153_ (.CLK(clknet_leaf_354_clk),
    .RESET_B(net835),
    .D(_02719_),
    .Q_N(_10783_),
    .Q(\atari2600.ram[56][2] ));
 sg13g2_dfrbp_1 _29154_ (.CLK(clknet_leaf_341_clk),
    .RESET_B(net833),
    .D(_02720_),
    .Q_N(_10782_),
    .Q(\atari2600.ram[56][3] ));
 sg13g2_dfrbp_1 _29155_ (.CLK(clknet_leaf_354_clk),
    .RESET_B(net831),
    .D(_02721_),
    .Q_N(_10781_),
    .Q(\atari2600.ram[56][4] ));
 sg13g2_dfrbp_1 _29156_ (.CLK(clknet_leaf_341_clk),
    .RESET_B(net829),
    .D(_02722_),
    .Q_N(_10780_),
    .Q(\atari2600.ram[56][5] ));
 sg13g2_dfrbp_1 _29157_ (.CLK(clknet_leaf_341_clk),
    .RESET_B(net827),
    .D(_02723_),
    .Q_N(_10779_),
    .Q(\atari2600.ram[56][6] ));
 sg13g2_dfrbp_1 _29158_ (.CLK(clknet_leaf_341_clk),
    .RESET_B(net825),
    .D(_02724_),
    .Q_N(_10778_),
    .Q(\atari2600.ram[56][7] ));
 sg13g2_dfrbp_1 _29159_ (.CLK(clknet_leaf_342_clk),
    .RESET_B(net823),
    .D(_02725_),
    .Q_N(_10777_),
    .Q(\atari2600.ram[57][0] ));
 sg13g2_dfrbp_1 _29160_ (.CLK(clknet_leaf_342_clk),
    .RESET_B(net821),
    .D(_02726_),
    .Q_N(_10776_),
    .Q(\atari2600.ram[57][1] ));
 sg13g2_dfrbp_1 _29161_ (.CLK(clknet_leaf_353_clk),
    .RESET_B(net819),
    .D(_02727_),
    .Q_N(_10775_),
    .Q(\atari2600.ram[57][2] ));
 sg13g2_dfrbp_1 _29162_ (.CLK(clknet_leaf_342_clk),
    .RESET_B(net817),
    .D(_02728_),
    .Q_N(_10774_),
    .Q(\atari2600.ram[57][3] ));
 sg13g2_dfrbp_1 _29163_ (.CLK(clknet_leaf_353_clk),
    .RESET_B(net815),
    .D(_02729_),
    .Q_N(_10773_),
    .Q(\atari2600.ram[57][4] ));
 sg13g2_dfrbp_1 _29164_ (.CLK(clknet_leaf_342_clk),
    .RESET_B(net813),
    .D(_02730_),
    .Q_N(_10772_),
    .Q(\atari2600.ram[57][5] ));
 sg13g2_dfrbp_1 _29165_ (.CLK(clknet_leaf_342_clk),
    .RESET_B(net811),
    .D(_02731_),
    .Q_N(_10771_),
    .Q(\atari2600.ram[57][6] ));
 sg13g2_dfrbp_1 _29166_ (.CLK(clknet_leaf_341_clk),
    .RESET_B(net809),
    .D(_02732_),
    .Q_N(_10770_),
    .Q(\atari2600.ram[57][7] ));
 sg13g2_dfrbp_1 _29167_ (.CLK(clknet_leaf_343_clk),
    .RESET_B(net750),
    .D(_02733_),
    .Q_N(_10769_),
    .Q(\atari2600.ram[58][0] ));
 sg13g2_dfrbp_1 _29168_ (.CLK(clknet_leaf_353_clk),
    .RESET_B(net748),
    .D(_02734_),
    .Q_N(_10768_),
    .Q(\atari2600.ram[58][1] ));
 sg13g2_dfrbp_1 _29169_ (.CLK(clknet_leaf_353_clk),
    .RESET_B(net746),
    .D(_02735_),
    .Q_N(_10767_),
    .Q(\atari2600.ram[58][2] ));
 sg13g2_dfrbp_1 _29170_ (.CLK(clknet_leaf_343_clk),
    .RESET_B(net744),
    .D(_02736_),
    .Q_N(_10766_),
    .Q(\atari2600.ram[58][3] ));
 sg13g2_dfrbp_1 _29171_ (.CLK(clknet_leaf_342_clk),
    .RESET_B(net742),
    .D(_02737_),
    .Q_N(_10765_),
    .Q(\atari2600.ram[58][4] ));
 sg13g2_dfrbp_1 _29172_ (.CLK(clknet_leaf_343_clk),
    .RESET_B(net653),
    .D(_02738_),
    .Q_N(_10764_),
    .Q(\atari2600.ram[58][5] ));
 sg13g2_dfrbp_1 _29173_ (.CLK(clknet_leaf_343_clk),
    .RESET_B(net651),
    .D(_02739_),
    .Q_N(_10763_),
    .Q(\atari2600.ram[58][6] ));
 sg13g2_dfrbp_1 _29174_ (.CLK(clknet_leaf_342_clk),
    .RESET_B(net649),
    .D(_02740_),
    .Q_N(_10762_),
    .Q(\atari2600.ram[58][7] ));
 sg13g2_dfrbp_1 _29175_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net647),
    .D(_02741_),
    .Q_N(_10761_),
    .Q(\atari2600.ram[5][0] ));
 sg13g2_dfrbp_1 _29176_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net645),
    .D(_02742_),
    .Q_N(_10760_),
    .Q(\atari2600.ram[5][1] ));
 sg13g2_dfrbp_1 _29177_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net643),
    .D(_02743_),
    .Q_N(_10759_),
    .Q(\atari2600.ram[5][2] ));
 sg13g2_dfrbp_1 _29178_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net641),
    .D(_02744_),
    .Q_N(_10758_),
    .Q(\atari2600.ram[5][3] ));
 sg13g2_dfrbp_1 _29179_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net639),
    .D(_02745_),
    .Q_N(_10757_),
    .Q(\atari2600.ram[5][4] ));
 sg13g2_dfrbp_1 _29180_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net637),
    .D(_02746_),
    .Q_N(_10756_),
    .Q(\atari2600.ram[5][5] ));
 sg13g2_dfrbp_1 _29181_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net635),
    .D(_02747_),
    .Q_N(_10755_),
    .Q(\atari2600.ram[5][6] ));
 sg13g2_dfrbp_1 _29182_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net633),
    .D(_02748_),
    .Q_N(_10754_),
    .Q(\atari2600.ram[5][7] ));
 sg13g2_dfrbp_1 _29183_ (.CLK(clknet_leaf_346_clk),
    .RESET_B(net631),
    .D(_02749_),
    .Q_N(_10753_),
    .Q(\atari2600.ram[60][0] ));
 sg13g2_dfrbp_1 _29184_ (.CLK(clknet_leaf_350_clk),
    .RESET_B(net629),
    .D(_02750_),
    .Q_N(_10752_),
    .Q(\atari2600.ram[60][1] ));
 sg13g2_dfrbp_1 _29185_ (.CLK(clknet_leaf_352_clk),
    .RESET_B(net627),
    .D(_02751_),
    .Q_N(_10751_),
    .Q(\atari2600.ram[60][2] ));
 sg13g2_dfrbp_1 _29186_ (.CLK(clknet_leaf_348_clk),
    .RESET_B(net625),
    .D(_02752_),
    .Q_N(_10750_),
    .Q(\atari2600.ram[60][3] ));
 sg13g2_dfrbp_1 _29187_ (.CLK(clknet_leaf_343_clk),
    .RESET_B(net623),
    .D(_02753_),
    .Q_N(_10749_),
    .Q(\atari2600.ram[60][4] ));
 sg13g2_dfrbp_1 _29188_ (.CLK(clknet_leaf_347_clk),
    .RESET_B(net621),
    .D(_02754_),
    .Q_N(_10748_),
    .Q(\atari2600.ram[60][5] ));
 sg13g2_dfrbp_1 _29189_ (.CLK(clknet_leaf_347_clk),
    .RESET_B(net619),
    .D(_02755_),
    .Q_N(_10747_),
    .Q(\atari2600.ram[60][6] ));
 sg13g2_dfrbp_1 _29190_ (.CLK(clknet_leaf_343_clk),
    .RESET_B(net617),
    .D(_02756_),
    .Q_N(_10746_),
    .Q(\atari2600.ram[60][7] ));
 sg13g2_dfrbp_1 _29191_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net615),
    .D(_02757_),
    .Q_N(_10745_),
    .Q(\atari2600.ram[61][0] ));
 sg13g2_dfrbp_1 _29192_ (.CLK(clknet_leaf_348_clk),
    .RESET_B(net613),
    .D(_02758_),
    .Q_N(_10744_),
    .Q(\atari2600.ram[61][1] ));
 sg13g2_dfrbp_1 _29193_ (.CLK(clknet_leaf_349_clk),
    .RESET_B(net611),
    .D(_02759_),
    .Q_N(_10743_),
    .Q(\atari2600.ram[61][2] ));
 sg13g2_dfrbp_1 _29194_ (.CLK(clknet_leaf_348_clk),
    .RESET_B(net609),
    .D(_02760_),
    .Q_N(_10742_),
    .Q(\atari2600.ram[61][3] ));
 sg13g2_dfrbp_1 _29195_ (.CLK(clknet_leaf_348_clk),
    .RESET_B(net607),
    .D(_02761_),
    .Q_N(_10741_),
    .Q(\atari2600.ram[61][4] ));
 sg13g2_dfrbp_1 _29196_ (.CLK(clknet_leaf_348_clk),
    .RESET_B(net605),
    .D(_02762_),
    .Q_N(_10740_),
    .Q(\atari2600.ram[61][5] ));
 sg13g2_dfrbp_1 _29197_ (.CLK(clknet_leaf_348_clk),
    .RESET_B(net603),
    .D(_02763_),
    .Q_N(_10739_),
    .Q(\atari2600.ram[61][6] ));
 sg13g2_dfrbp_1 _29198_ (.CLK(clknet_leaf_346_clk),
    .RESET_B(net601),
    .D(_02764_),
    .Q_N(_10738_),
    .Q(\atari2600.ram[61][7] ));
 sg13g2_dfrbp_1 _29199_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net599),
    .D(_02765_),
    .Q_N(_10737_),
    .Q(\atari2600.ram[62][0] ));
 sg13g2_dfrbp_1 _29200_ (.CLK(clknet_leaf_348_clk),
    .RESET_B(net597),
    .D(_02766_),
    .Q_N(_10736_),
    .Q(\atari2600.ram[62][1] ));
 sg13g2_dfrbp_1 _29201_ (.CLK(clknet_leaf_349_clk),
    .RESET_B(net595),
    .D(_02767_),
    .Q_N(_10735_),
    .Q(\atari2600.ram[62][2] ));
 sg13g2_dfrbp_1 _29202_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net593),
    .D(_02768_),
    .Q_N(_10734_),
    .Q(\atari2600.ram[62][3] ));
 sg13g2_dfrbp_1 _29203_ (.CLK(clknet_leaf_347_clk),
    .RESET_B(net591),
    .D(_02769_),
    .Q_N(_10733_),
    .Q(\atari2600.ram[62][4] ));
 sg13g2_dfrbp_1 _29204_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net589),
    .D(_02770_),
    .Q_N(_10732_),
    .Q(\atari2600.ram[62][5] ));
 sg13g2_dfrbp_1 _29205_ (.CLK(clknet_leaf_320_clk),
    .RESET_B(net587),
    .D(_02771_),
    .Q_N(_10731_),
    .Q(\atari2600.ram[62][6] ));
 sg13g2_dfrbp_1 _29206_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net585),
    .D(_02772_),
    .Q_N(_10730_),
    .Q(\atari2600.ram[62][7] ));
 sg13g2_dfrbp_1 _29207_ (.CLK(clknet_leaf_346_clk),
    .RESET_B(net583),
    .D(_02773_),
    .Q_N(_10729_),
    .Q(\atari2600.ram[63][0] ));
 sg13g2_dfrbp_1 _29208_ (.CLK(clknet_leaf_349_clk),
    .RESET_B(net581),
    .D(_02774_),
    .Q_N(_10728_),
    .Q(\atari2600.ram[63][1] ));
 sg13g2_dfrbp_1 _29209_ (.CLK(clknet_leaf_346_clk),
    .RESET_B(net576),
    .D(_02775_),
    .Q_N(_10727_),
    .Q(\atari2600.ram[63][2] ));
 sg13g2_dfrbp_1 _29210_ (.CLK(clknet_leaf_348_clk),
    .RESET_B(net574),
    .D(_02776_),
    .Q_N(_10726_),
    .Q(\atari2600.ram[63][3] ));
 sg13g2_dfrbp_1 _29211_ (.CLK(clknet_leaf_346_clk),
    .RESET_B(net572),
    .D(_02777_),
    .Q_N(_10725_),
    .Q(\atari2600.ram[63][4] ));
 sg13g2_dfrbp_1 _29212_ (.CLK(clknet_leaf_347_clk),
    .RESET_B(net570),
    .D(_02778_),
    .Q_N(_10724_),
    .Q(\atari2600.ram[63][5] ));
 sg13g2_dfrbp_1 _29213_ (.CLK(clknet_leaf_347_clk),
    .RESET_B(net568),
    .D(_02779_),
    .Q_N(_10723_),
    .Q(\atari2600.ram[63][6] ));
 sg13g2_dfrbp_1 _29214_ (.CLK(clknet_leaf_346_clk),
    .RESET_B(net566),
    .D(_02780_),
    .Q_N(_10722_),
    .Q(\atari2600.ram[63][7] ));
 sg13g2_dfrbp_1 _29215_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net564),
    .D(_02781_),
    .Q_N(_10721_),
    .Q(\atari2600.ram[64][0] ));
 sg13g2_dfrbp_1 _29216_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net562),
    .D(_02782_),
    .Q_N(_10720_),
    .Q(\atari2600.ram[64][1] ));
 sg13g2_dfrbp_1 _29217_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net560),
    .D(_02783_),
    .Q_N(_10719_),
    .Q(\atari2600.ram[64][2] ));
 sg13g2_dfrbp_1 _29218_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net558),
    .D(_02784_),
    .Q_N(_10718_),
    .Q(\atari2600.ram[64][3] ));
 sg13g2_dfrbp_1 _29219_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net556),
    .D(_02785_),
    .Q_N(_10717_),
    .Q(\atari2600.ram[64][4] ));
 sg13g2_dfrbp_1 _29220_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net554),
    .D(_02786_),
    .Q_N(_10716_),
    .Q(\atari2600.ram[64][5] ));
 sg13g2_dfrbp_1 _29221_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net552),
    .D(_02787_),
    .Q_N(_10715_),
    .Q(\atari2600.ram[64][6] ));
 sg13g2_dfrbp_1 _29222_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net550),
    .D(_02788_),
    .Q_N(_10714_),
    .Q(\atari2600.ram[64][7] ));
 sg13g2_dfrbp_1 _29223_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net548),
    .D(_02789_),
    .Q_N(_10713_),
    .Q(\atari2600.ram[65][0] ));
 sg13g2_dfrbp_1 _29224_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net546),
    .D(_02790_),
    .Q_N(_10712_),
    .Q(\atari2600.ram[65][1] ));
 sg13g2_dfrbp_1 _29225_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net544),
    .D(_02791_),
    .Q_N(_10711_),
    .Q(\atari2600.ram[65][2] ));
 sg13g2_dfrbp_1 _29226_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net542),
    .D(_02792_),
    .Q_N(_10710_),
    .Q(\atari2600.ram[65][3] ));
 sg13g2_dfrbp_1 _29227_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net540),
    .D(_02793_),
    .Q_N(_10709_),
    .Q(\atari2600.ram[65][4] ));
 sg13g2_dfrbp_1 _29228_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net538),
    .D(_02794_),
    .Q_N(_10708_),
    .Q(\atari2600.ram[65][5] ));
 sg13g2_dfrbp_1 _29229_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net536),
    .D(_02795_),
    .Q_N(_10707_),
    .Q(\atari2600.ram[65][6] ));
 sg13g2_dfrbp_1 _29230_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net534),
    .D(_02796_),
    .Q_N(_10706_),
    .Q(\atari2600.ram[65][7] ));
 sg13g2_dfrbp_1 _29231_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net532),
    .D(_02797_),
    .Q_N(_10705_),
    .Q(\atari2600.ram[66][0] ));
 sg13g2_dfrbp_1 _29232_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net530),
    .D(_02798_),
    .Q_N(_10704_),
    .Q(\atari2600.ram[66][1] ));
 sg13g2_dfrbp_1 _29233_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net528),
    .D(_02799_),
    .Q_N(_10703_),
    .Q(\atari2600.ram[66][2] ));
 sg13g2_dfrbp_1 _29234_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net526),
    .D(_02800_),
    .Q_N(_10702_),
    .Q(\atari2600.ram[66][3] ));
 sg13g2_dfrbp_1 _29235_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net524),
    .D(_02801_),
    .Q_N(_10701_),
    .Q(\atari2600.ram[66][4] ));
 sg13g2_dfrbp_1 _29236_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net522),
    .D(_02802_),
    .Q_N(_10700_),
    .Q(\atari2600.ram[66][5] ));
 sg13g2_dfrbp_1 _29237_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net520),
    .D(_02803_),
    .Q_N(_10699_),
    .Q(\atari2600.ram[66][6] ));
 sg13g2_dfrbp_1 _29238_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net518),
    .D(_02804_),
    .Q_N(_10698_),
    .Q(\atari2600.ram[66][7] ));
 sg13g2_dfrbp_1 _29239_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net516),
    .D(_02805_),
    .Q_N(_10697_),
    .Q(\atari2600.ram[67][0] ));
 sg13g2_dfrbp_1 _29240_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net507),
    .D(_02806_),
    .Q_N(_10696_),
    .Q(\atari2600.ram[67][1] ));
 sg13g2_dfrbp_1 _29241_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net505),
    .D(_02807_),
    .Q_N(_10695_),
    .Q(\atari2600.ram[67][2] ));
 sg13g2_dfrbp_1 _29242_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net503),
    .D(_02808_),
    .Q_N(_10694_),
    .Q(\atari2600.ram[67][3] ));
 sg13g2_dfrbp_1 _29243_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net501),
    .D(_02809_),
    .Q_N(_10693_),
    .Q(\atari2600.ram[67][4] ));
 sg13g2_dfrbp_1 _29244_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net499),
    .D(_02810_),
    .Q_N(_10692_),
    .Q(\atari2600.ram[67][5] ));
 sg13g2_dfrbp_1 _29245_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net497),
    .D(_02811_),
    .Q_N(_10691_),
    .Q(\atari2600.ram[67][6] ));
 sg13g2_dfrbp_1 _29246_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net495),
    .D(_02812_),
    .Q_N(_10690_),
    .Q(\atari2600.ram[67][7] ));
 sg13g2_dfrbp_1 _29247_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net493),
    .D(_02813_),
    .Q_N(_10689_),
    .Q(\atari2600.ram[68][0] ));
 sg13g2_dfrbp_1 _29248_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net491),
    .D(_02814_),
    .Q_N(_10688_),
    .Q(\atari2600.ram[68][1] ));
 sg13g2_dfrbp_1 _29249_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net489),
    .D(_02815_),
    .Q_N(_10687_),
    .Q(\atari2600.ram[68][2] ));
 sg13g2_dfrbp_1 _29250_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net487),
    .D(_02816_),
    .Q_N(_10686_),
    .Q(\atari2600.ram[68][3] ));
 sg13g2_dfrbp_1 _29251_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net485),
    .D(_02817_),
    .Q_N(_10685_),
    .Q(\atari2600.ram[68][4] ));
 sg13g2_dfrbp_1 _29252_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net483),
    .D(_02818_),
    .Q_N(_10684_),
    .Q(\atari2600.ram[68][5] ));
 sg13g2_dfrbp_1 _29253_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net481),
    .D(_02819_),
    .Q_N(_10683_),
    .Q(\atari2600.ram[68][6] ));
 sg13g2_dfrbp_1 _29254_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net479),
    .D(_02820_),
    .Q_N(_10682_),
    .Q(\atari2600.ram[68][7] ));
 sg13g2_dfrbp_1 _29255_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net477),
    .D(_02821_),
    .Q_N(_10681_),
    .Q(\atari2600.ram[20][0] ));
 sg13g2_dfrbp_1 _29256_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net475),
    .D(_02822_),
    .Q_N(_10680_),
    .Q(\atari2600.ram[20][1] ));
 sg13g2_dfrbp_1 _29257_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net473),
    .D(_02823_),
    .Q_N(_10679_),
    .Q(\atari2600.ram[20][2] ));
 sg13g2_dfrbp_1 _29258_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net471),
    .D(_02824_),
    .Q_N(_10678_),
    .Q(\atari2600.ram[20][3] ));
 sg13g2_dfrbp_1 _29259_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net469),
    .D(_02825_),
    .Q_N(_10677_),
    .Q(\atari2600.ram[20][4] ));
 sg13g2_dfrbp_1 _29260_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net467),
    .D(_02826_),
    .Q_N(_10676_),
    .Q(\atari2600.ram[20][5] ));
 sg13g2_dfrbp_1 _29261_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net465),
    .D(_02827_),
    .Q_N(_10675_),
    .Q(\atari2600.ram[20][6] ));
 sg13g2_dfrbp_1 _29262_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net463),
    .D(_02828_),
    .Q_N(_10674_),
    .Q(\atari2600.ram[20][7] ));
 sg13g2_dfrbp_1 _29263_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net446),
    .D(_02829_),
    .Q_N(_10673_),
    .Q(\atari2600.ram[1][0] ));
 sg13g2_dfrbp_1 _29264_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net444),
    .D(_02830_),
    .Q_N(_10672_),
    .Q(\atari2600.ram[1][1] ));
 sg13g2_dfrbp_1 _29265_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net442),
    .D(_02831_),
    .Q_N(_10671_),
    .Q(\atari2600.ram[1][2] ));
 sg13g2_dfrbp_1 _29266_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net440),
    .D(_02832_),
    .Q_N(_10670_),
    .Q(\atari2600.ram[1][3] ));
 sg13g2_dfrbp_1 _29267_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net438),
    .D(_02833_),
    .Q_N(_10669_),
    .Q(\atari2600.ram[1][4] ));
 sg13g2_dfrbp_1 _29268_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net436),
    .D(_02834_),
    .Q_N(_10668_),
    .Q(\atari2600.ram[1][5] ));
 sg13g2_dfrbp_1 _29269_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net434),
    .D(_02835_),
    .Q_N(_10667_),
    .Q(\atari2600.ram[1][6] ));
 sg13g2_dfrbp_1 _29270_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net432),
    .D(_02836_),
    .Q_N(_10666_),
    .Q(\atari2600.ram[1][7] ));
 sg13g2_dfrbp_1 _29271_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net430),
    .D(_02837_),
    .Q_N(_10665_),
    .Q(\atari2600.ram[18][0] ));
 sg13g2_dfrbp_1 _29272_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net428),
    .D(_02838_),
    .Q_N(_10664_),
    .Q(\atari2600.ram[18][1] ));
 sg13g2_dfrbp_1 _29273_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net426),
    .D(_02839_),
    .Q_N(_10663_),
    .Q(\atari2600.ram[18][2] ));
 sg13g2_dfrbp_1 _29274_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net424),
    .D(_02840_),
    .Q_N(_10662_),
    .Q(\atari2600.ram[18][3] ));
 sg13g2_dfrbp_1 _29275_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net422),
    .D(_02841_),
    .Q_N(_10661_),
    .Q(\atari2600.ram[18][4] ));
 sg13g2_dfrbp_1 _29276_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net420),
    .D(_02842_),
    .Q_N(_10660_),
    .Q(\atari2600.ram[18][5] ));
 sg13g2_dfrbp_1 _29277_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net418),
    .D(_02843_),
    .Q_N(_10659_),
    .Q(\atari2600.ram[18][6] ));
 sg13g2_dfrbp_1 _29278_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net416),
    .D(_02844_),
    .Q_N(_10658_),
    .Q(\atari2600.ram[18][7] ));
 sg13g2_dfrbp_1 _29279_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net414),
    .D(_02845_),
    .Q_N(_10657_),
    .Q(\atari2600.ram[17][0] ));
 sg13g2_dfrbp_1 _29280_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net412),
    .D(_02846_),
    .Q_N(_10656_),
    .Q(\atari2600.ram[17][1] ));
 sg13g2_dfrbp_1 _29281_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net410),
    .D(_02847_),
    .Q_N(_10655_),
    .Q(\atari2600.ram[17][2] ));
 sg13g2_dfrbp_1 _29282_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net408),
    .D(_02848_),
    .Q_N(_10654_),
    .Q(\atari2600.ram[17][3] ));
 sg13g2_dfrbp_1 _29283_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net406),
    .D(_02849_),
    .Q_N(_10653_),
    .Q(\atari2600.ram[17][4] ));
 sg13g2_dfrbp_1 _29284_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net404),
    .D(_02850_),
    .Q_N(_10652_),
    .Q(\atari2600.ram[17][5] ));
 sg13g2_dfrbp_1 _29285_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net402),
    .D(_02851_),
    .Q_N(_10651_),
    .Q(\atari2600.ram[17][6] ));
 sg13g2_dfrbp_1 _29286_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net400),
    .D(_02852_),
    .Q_N(_10650_),
    .Q(\atari2600.ram[17][7] ));
 sg13g2_dfrbp_1 _29287_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net398),
    .D(_02853_),
    .Q_N(_10649_),
    .Q(\atari2600.address_bus_r[0] ));
 sg13g2_dfrbp_1 _29288_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net396),
    .D(_02854_),
    .Q_N(_10648_),
    .Q(\atari2600.address_bus_r[1] ));
 sg13g2_dfrbp_1 _29289_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net394),
    .D(_02855_),
    .Q_N(_10647_),
    .Q(\atari2600.address_bus_r[2] ));
 sg13g2_dfrbp_1 _29290_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net392),
    .D(_02856_),
    .Q_N(_10646_),
    .Q(\atari2600.address_bus_r[3] ));
 sg13g2_dfrbp_1 _29291_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net390),
    .D(_02857_),
    .Q_N(_10645_),
    .Q(\atari2600.address_bus_r[4] ));
 sg13g2_dfrbp_1 _29292_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net388),
    .D(_02858_),
    .Q_N(_10644_),
    .Q(\atari2600.address_bus_r[5] ));
 sg13g2_dfrbp_1 _29293_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net386),
    .D(_02859_),
    .Q_N(_10643_),
    .Q(\atari2600.address_bus_r[6] ));
 sg13g2_dfrbp_1 _29294_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net384),
    .D(_02860_),
    .Q_N(_10642_),
    .Q(\atari2600.address_bus_r[7] ));
 sg13g2_dfrbp_1 _29295_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net382),
    .D(_02861_),
    .Q_N(_10641_),
    .Q(\atari2600.address_bus_r[8] ));
 sg13g2_dfrbp_1 _29296_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net380),
    .D(_02862_),
    .Q_N(_10640_),
    .Q(\atari2600.address_bus_r[9] ));
 sg13g2_dfrbp_1 _29297_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net378),
    .D(_02863_),
    .Q_N(_10639_),
    .Q(\atari2600.address_bus_r[10] ));
 sg13g2_dfrbp_1 _29298_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net376),
    .D(_02864_),
    .Q_N(_10638_),
    .Q(\atari2600.address_bus_r[11] ));
 sg13g2_dfrbp_1 _29299_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net374),
    .D(_02865_),
    .Q_N(_10637_),
    .Q(\atari2600.address_bus_r[12] ));
 sg13g2_dfrbp_1 _29300_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net372),
    .D(_02866_),
    .Q_N(_10636_),
    .Q(\atari2600.ram[16][0] ));
 sg13g2_dfrbp_1 _29301_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net370),
    .D(_02867_),
    .Q_N(_10635_),
    .Q(\atari2600.ram[16][1] ));
 sg13g2_dfrbp_1 _29302_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net368),
    .D(_02868_),
    .Q_N(_10634_),
    .Q(\atari2600.ram[16][2] ));
 sg13g2_dfrbp_1 _29303_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net366),
    .D(_02869_),
    .Q_N(_10633_),
    .Q(\atari2600.ram[16][3] ));
 sg13g2_dfrbp_1 _29304_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net364),
    .D(_02870_),
    .Q_N(_10632_),
    .Q(\atari2600.ram[16][4] ));
 sg13g2_dfrbp_1 _29305_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net362),
    .D(_02871_),
    .Q_N(_10631_),
    .Q(\atari2600.ram[16][5] ));
 sg13g2_dfrbp_1 _29306_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net360),
    .D(_02872_),
    .Q_N(_10630_),
    .Q(\atari2600.ram[16][6] ));
 sg13g2_dfrbp_1 _29307_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net358),
    .D(_02873_),
    .Q_N(_10629_),
    .Q(\atari2600.ram[16][7] ));
 sg13g2_dfrbp_1 _29308_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net356),
    .D(_02874_),
    .Q_N(_10628_),
    .Q(\atari2600.ram[15][0] ));
 sg13g2_dfrbp_1 _29309_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net354),
    .D(_02875_),
    .Q_N(_10627_),
    .Q(\atari2600.ram[15][1] ));
 sg13g2_dfrbp_1 _29310_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net352),
    .D(_02876_),
    .Q_N(_10626_),
    .Q(\atari2600.ram[15][2] ));
 sg13g2_dfrbp_1 _29311_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net350),
    .D(_02877_),
    .Q_N(_10625_),
    .Q(\atari2600.ram[15][3] ));
 sg13g2_dfrbp_1 _29312_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net348),
    .D(_02878_),
    .Q_N(_10624_),
    .Q(\atari2600.ram[15][4] ));
 sg13g2_dfrbp_1 _29313_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net346),
    .D(_02879_),
    .Q_N(_10623_),
    .Q(\atari2600.ram[15][5] ));
 sg13g2_dfrbp_1 _29314_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net344),
    .D(_02880_),
    .Q_N(_10622_),
    .Q(\atari2600.ram[15][6] ));
 sg13g2_dfrbp_1 _29315_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net342),
    .D(_02881_),
    .Q_N(_10621_),
    .Q(\atari2600.ram[15][7] ));
 sg13g2_dfrbp_1 _29316_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net340),
    .D(_02882_),
    .Q_N(_10620_),
    .Q(\atari2600.ram[126][0] ));
 sg13g2_dfrbp_1 _29317_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net338),
    .D(_02883_),
    .Q_N(_10619_),
    .Q(\atari2600.ram[126][1] ));
 sg13g2_dfrbp_1 _29318_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net336),
    .D(_02884_),
    .Q_N(_10618_),
    .Q(\atari2600.ram[126][2] ));
 sg13g2_dfrbp_1 _29319_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net334),
    .D(_02885_),
    .Q_N(_10617_),
    .Q(\atari2600.ram[126][3] ));
 sg13g2_dfrbp_1 _29320_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net332),
    .D(_02886_),
    .Q_N(_10616_),
    .Q(\atari2600.ram[126][4] ));
 sg13g2_dfrbp_1 _29321_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net330),
    .D(_02887_),
    .Q_N(_10615_),
    .Q(\atari2600.ram[126][5] ));
 sg13g2_dfrbp_1 _29322_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net328),
    .D(_02888_),
    .Q_N(_10614_),
    .Q(\atari2600.ram[126][6] ));
 sg13g2_dfrbp_1 _29323_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net326),
    .D(_02889_),
    .Q_N(_10613_),
    .Q(\atari2600.ram[126][7] ));
 sg13g2_dfrbp_1 _29324_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net324),
    .D(_02890_),
    .Q_N(_10612_),
    .Q(\atari2600.ram[14][0] ));
 sg13g2_dfrbp_1 _29325_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net322),
    .D(_02891_),
    .Q_N(_10611_),
    .Q(\atari2600.ram[14][1] ));
 sg13g2_dfrbp_1 _29326_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net320),
    .D(_02892_),
    .Q_N(_10610_),
    .Q(\atari2600.ram[14][2] ));
 sg13g2_dfrbp_1 _29327_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net318),
    .D(_02893_),
    .Q_N(_10609_),
    .Q(\atari2600.ram[14][3] ));
 sg13g2_dfrbp_1 _29328_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net316),
    .D(_02894_),
    .Q_N(_10608_),
    .Q(\atari2600.ram[14][4] ));
 sg13g2_dfrbp_1 _29329_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net314),
    .D(_02895_),
    .Q_N(_10607_),
    .Q(\atari2600.ram[14][5] ));
 sg13g2_dfrbp_1 _29330_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net312),
    .D(_02896_),
    .Q_N(_10606_),
    .Q(\atari2600.ram[14][6] ));
 sg13g2_dfrbp_1 _29331_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net310),
    .D(_02897_),
    .Q_N(_10605_),
    .Q(\atari2600.ram[14][7] ));
 sg13g2_dfrbp_1 _29332_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net308),
    .D(_02898_),
    .Q_N(_10604_),
    .Q(\atari2600.ram[124][0] ));
 sg13g2_dfrbp_1 _29333_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net306),
    .D(_02899_),
    .Q_N(_10603_),
    .Q(\atari2600.ram[124][1] ));
 sg13g2_dfrbp_1 _29334_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net304),
    .D(_02900_),
    .Q_N(_10602_),
    .Q(\atari2600.ram[124][2] ));
 sg13g2_dfrbp_1 _29335_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net302),
    .D(_02901_),
    .Q_N(_10601_),
    .Q(\atari2600.ram[124][3] ));
 sg13g2_dfrbp_1 _29336_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net300),
    .D(_02902_),
    .Q_N(_10600_),
    .Q(\atari2600.ram[124][4] ));
 sg13g2_dfrbp_1 _29337_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net298),
    .D(_02903_),
    .Q_N(_10599_),
    .Q(\atari2600.ram[124][5] ));
 sg13g2_dfrbp_1 _29338_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net296),
    .D(_02904_),
    .Q_N(_10598_),
    .Q(\atari2600.ram[124][6] ));
 sg13g2_dfrbp_1 _29339_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net294),
    .D(_02905_),
    .Q_N(_10597_),
    .Q(\atari2600.ram[124][7] ));
 sg13g2_dfrbp_1 _29340_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net292),
    .D(_02906_),
    .Q_N(_10596_),
    .Q(\atari2600.ram[125][0] ));
 sg13g2_dfrbp_1 _29341_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net290),
    .D(_02907_),
    .Q_N(_10595_),
    .Q(\atari2600.ram[125][1] ));
 sg13g2_dfrbp_1 _29342_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net288),
    .D(_02908_),
    .Q_N(_10594_),
    .Q(\atari2600.ram[125][2] ));
 sg13g2_dfrbp_1 _29343_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net286),
    .D(_02909_),
    .Q_N(_10593_),
    .Q(\atari2600.ram[125][3] ));
 sg13g2_dfrbp_1 _29344_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net284),
    .D(_02910_),
    .Q_N(_10592_),
    .Q(\atari2600.ram[125][4] ));
 sg13g2_dfrbp_1 _29345_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net282),
    .D(_02911_),
    .Q_N(_10591_),
    .Q(\atari2600.ram[125][5] ));
 sg13g2_dfrbp_1 _29346_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net280),
    .D(_02912_),
    .Q_N(_10590_),
    .Q(\atari2600.ram[125][6] ));
 sg13g2_dfrbp_1 _29347_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net278),
    .D(_02913_),
    .Q_N(_10589_),
    .Q(\atari2600.ram[125][7] ));
 sg13g2_dfrbp_1 _29348_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net276),
    .D(_02914_),
    .Q_N(_10588_),
    .Q(\flash_rom.nibbles_remaining[0] ));
 sg13g2_dfrbp_1 _29349_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net272),
    .D(_02915_),
    .Q_N(_10587_),
    .Q(\flash_rom.nibbles_remaining[1] ));
 sg13g2_dfrbp_1 _29350_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net268),
    .D(_02916_),
    .Q_N(_10586_),
    .Q(\flash_rom.nibbles_remaining[2] ));
 sg13g2_dfrbp_1 _29351_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net264),
    .D(_02917_),
    .Q_N(_00138_),
    .Q(\flash_rom.fsm_state[0] ));
 sg13g2_dfrbp_1 _29352_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net260),
    .D(_02918_),
    .Q_N(_10585_),
    .Q(\flash_rom.fsm_state[1] ));
 sg13g2_dfrbp_1 _29353_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net256),
    .D(_02919_),
    .Q_N(_00102_),
    .Q(\flash_rom.fsm_state[2] ));
 sg13g2_dfrbp_1 _29354_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net252),
    .D(_02920_),
    .Q_N(_10584_),
    .Q(\atari2600.rom_data[0] ));
 sg13g2_dfrbp_1 _29355_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net250),
    .D(_02921_),
    .Q_N(_10583_),
    .Q(\atari2600.rom_data[1] ));
 sg13g2_dfrbp_1 _29356_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net248),
    .D(_02922_),
    .Q_N(_10582_),
    .Q(\atari2600.rom_data[2] ));
 sg13g2_dfrbp_1 _29357_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net246),
    .D(_02923_),
    .Q_N(_10581_),
    .Q(\atari2600.rom_data[3] ));
 sg13g2_dfrbp_1 _29358_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net244),
    .D(net3173),
    .Q_N(_10580_),
    .Q(\atari2600.rom_data[4] ));
 sg13g2_dfrbp_1 _29359_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net242),
    .D(net3002),
    .Q_N(_10579_),
    .Q(\atari2600.rom_data[5] ));
 sg13g2_dfrbp_1 _29360_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net240),
    .D(net3966),
    .Q_N(_10578_),
    .Q(\atari2600.rom_data[6] ));
 sg13g2_dfrbp_1 _29361_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net238),
    .D(net3355),
    .Q_N(_10577_),
    .Q(\atari2600.rom_data[7] ));
 sg13g2_dfrbp_1 _29362_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net236),
    .D(_02928_),
    .Q_N(_00137_),
    .Q(\flash_rom.spi_clk_out ));
 sg13g2_dfrbp_1 _29363_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net232),
    .D(_02929_),
    .Q_N(_10576_),
    .Q(uio_oe[1]));
 sg13g2_dfrbp_1 _29364_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net228),
    .D(net7216),
    .Q_N(_10575_),
    .Q(uio_oe[5]));
 sg13g2_dfrbp_1 _29365_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net224),
    .D(_02931_),
    .Q_N(_10574_),
    .Q(\atari2600.tia.p1_spacing[4] ));
 sg13g2_dfrbp_1 _29366_ (.CLK(clknet_leaf_307_clk),
    .RESET_B(net220),
    .D(_02932_),
    .Q_N(_10573_),
    .Q(\atari2600.tia.p1_spacing[5] ));
 sg13g2_dfrbp_1 _29367_ (.CLK(clknet_leaf_308_clk),
    .RESET_B(net216),
    .D(_02933_),
    .Q_N(_10572_),
    .Q(\atari2600.tia.p1_spacing[6] ));
 sg13g2_dfrbp_1 _29368_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net212),
    .D(_02934_),
    .Q_N(_10571_),
    .Q(\atari2600.ram[40][0] ));
 sg13g2_dfrbp_1 _29369_ (.CLK(clknet_leaf_349_clk),
    .RESET_B(net210),
    .D(_02935_),
    .Q_N(_10570_),
    .Q(\atari2600.ram[40][1] ));
 sg13g2_dfrbp_1 _29370_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net208),
    .D(_02936_),
    .Q_N(_10569_),
    .Q(\atari2600.ram[40][2] ));
 sg13g2_dfrbp_1 _29371_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net206),
    .D(_02937_),
    .Q_N(_10568_),
    .Q(\atari2600.ram[40][3] ));
 sg13g2_dfrbp_1 _29372_ (.CLK(clknet_leaf_350_clk),
    .RESET_B(net204),
    .D(_02938_),
    .Q_N(_10567_),
    .Q(\atari2600.ram[40][4] ));
 sg13g2_dfrbp_1 _29373_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net202),
    .D(_02939_),
    .Q_N(_10566_),
    .Q(\atari2600.ram[40][5] ));
 sg13g2_dfrbp_1 _29374_ (.CLK(clknet_leaf_350_clk),
    .RESET_B(net200),
    .D(_02940_),
    .Q_N(_10565_),
    .Q(\atari2600.ram[40][6] ));
 sg13g2_dfrbp_1 _29375_ (.CLK(clknet_leaf_350_clk),
    .RESET_B(net198),
    .D(_02941_),
    .Q_N(_10564_),
    .Q(\atari2600.ram[40][7] ));
 sg13g2_dfrbp_1 _29376_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net196),
    .D(_02942_),
    .Q_N(_10563_),
    .Q(\atari2600.ram[41][0] ));
 sg13g2_dfrbp_1 _29377_ (.CLK(clknet_leaf_349_clk),
    .RESET_B(net194),
    .D(_02943_),
    .Q_N(_10562_),
    .Q(\atari2600.ram[41][1] ));
 sg13g2_dfrbp_1 _29378_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net192),
    .D(_02944_),
    .Q_N(_10561_),
    .Q(\atari2600.ram[41][2] ));
 sg13g2_dfrbp_1 _29379_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net190),
    .D(_02945_),
    .Q_N(_10560_),
    .Q(\atari2600.ram[41][3] ));
 sg13g2_dfrbp_1 _29380_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net188),
    .D(_02946_),
    .Q_N(_10559_),
    .Q(\atari2600.ram[41][4] ));
 sg13g2_dfrbp_1 _29381_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net186),
    .D(_02947_),
    .Q_N(_10558_),
    .Q(\atari2600.ram[41][5] ));
 sg13g2_dfrbp_1 _29382_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net64),
    .D(_02948_),
    .Q_N(_10557_),
    .Q(\atari2600.ram[41][6] ));
 sg13g2_dfrbp_1 _29383_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net62),
    .D(_02949_),
    .Q_N(_10556_),
    .Q(\atari2600.ram[41][7] ));
 sg13g2_dfrbp_1 _29384_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net60),
    .D(_02950_),
    .Q_N(_10555_),
    .Q(\atari2600.ram[3][0] ));
 sg13g2_dfrbp_1 _29385_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net58),
    .D(_02951_),
    .Q_N(_10554_),
    .Q(\atari2600.ram[3][1] ));
 sg13g2_dfrbp_1 _29386_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net56),
    .D(_02952_),
    .Q_N(_10553_),
    .Q(\atari2600.ram[3][2] ));
 sg13g2_dfrbp_1 _29387_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net54),
    .D(_02953_),
    .Q_N(_10552_),
    .Q(\atari2600.ram[3][3] ));
 sg13g2_dfrbp_1 _29388_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net52),
    .D(_02954_),
    .Q_N(_10551_),
    .Q(\atari2600.ram[3][4] ));
 sg13g2_dfrbp_1 _29389_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net50),
    .D(_02955_),
    .Q_N(_10550_),
    .Q(\atari2600.ram[3][5] ));
 sg13g2_dfrbp_1 _29390_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net48),
    .D(_02956_),
    .Q_N(_10549_),
    .Q(\atari2600.ram[3][6] ));
 sg13g2_dfrbp_1 _29391_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net46),
    .D(_02957_),
    .Q_N(_10548_),
    .Q(\atari2600.ram[3][7] ));
 sg13g2_dfrbp_1 _29392_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net44),
    .D(_02958_),
    .Q_N(_10547_),
    .Q(\atari2600.ram[38][0] ));
 sg13g2_dfrbp_1 _29393_ (.CLK(clknet_leaf_351_clk),
    .RESET_B(net42),
    .D(_02959_),
    .Q_N(_10546_),
    .Q(\atari2600.ram[38][1] ));
 sg13g2_dfrbp_1 _29394_ (.CLK(clknet_leaf_358_clk),
    .RESET_B(net2867),
    .D(_02960_),
    .Q_N(_10545_),
    .Q(\atari2600.ram[38][2] ));
 sg13g2_dfrbp_1 _29395_ (.CLK(clknet_leaf_351_clk),
    .RESET_B(net2858),
    .D(_02961_),
    .Q_N(_10544_),
    .Q(\atari2600.ram[38][3] ));
 sg13g2_dfrbp_1 _29396_ (.CLK(clknet_leaf_351_clk),
    .RESET_B(net2847),
    .D(_02962_),
    .Q_N(_10543_),
    .Q(\atari2600.ram[38][4] ));
 sg13g2_dfrbp_1 _29397_ (.CLK(clknet_leaf_351_clk),
    .RESET_B(net2837),
    .D(_02963_),
    .Q_N(_10542_),
    .Q(\atari2600.ram[38][5] ));
 sg13g2_dfrbp_1 _29398_ (.CLK(clknet_leaf_350_clk),
    .RESET_B(net2835),
    .D(_02964_),
    .Q_N(_10541_),
    .Q(\atari2600.ram[38][6] ));
 sg13g2_dfrbp_1 _29399_ (.CLK(clknet_leaf_358_clk),
    .RESET_B(net2739),
    .D(_02965_),
    .Q_N(_10540_),
    .Q(\atari2600.ram[38][7] ));
 sg13g2_dfrbp_1 _29400_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net2737),
    .D(_02966_),
    .Q_N(_10539_),
    .Q(\atari2600.ram[37][0] ));
 sg13g2_dfrbp_1 _29401_ (.CLK(clknet_leaf_356_clk),
    .RESET_B(net2735),
    .D(_02967_),
    .Q_N(_10538_),
    .Q(\atari2600.ram[37][1] ));
 sg13g2_dfrbp_1 _29402_ (.CLK(clknet_leaf_360_clk),
    .RESET_B(net2733),
    .D(_02968_),
    .Q_N(_10537_),
    .Q(\atari2600.ram[37][2] ));
 sg13g2_dfrbp_1 _29403_ (.CLK(clknet_leaf_360_clk),
    .RESET_B(net2731),
    .D(_02969_),
    .Q_N(_10536_),
    .Q(\atari2600.ram[37][3] ));
 sg13g2_dfrbp_1 _29404_ (.CLK(clknet_leaf_357_clk),
    .RESET_B(net2729),
    .D(_02970_),
    .Q_N(_10535_),
    .Q(\atari2600.ram[37][4] ));
 sg13g2_dfrbp_1 _29405_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net2727),
    .D(_02971_),
    .Q_N(_10534_),
    .Q(\atari2600.ram[37][5] ));
 sg13g2_dfrbp_1 _29406_ (.CLK(clknet_leaf_358_clk),
    .RESET_B(net2725),
    .D(_02972_),
    .Q_N(_10533_),
    .Q(\atari2600.ram[37][6] ));
 sg13g2_dfrbp_1 _29407_ (.CLK(clknet_leaf_358_clk),
    .RESET_B(net2723),
    .D(_02973_),
    .Q_N(_10532_),
    .Q(\atari2600.ram[37][7] ));
 sg13g2_dfrbp_1 _29408_ (.CLK(clknet_leaf_359_clk),
    .RESET_B(net2705),
    .D(_02974_),
    .Q_N(_10531_),
    .Q(\atari2600.ram[36][0] ));
 sg13g2_dfrbp_1 _29409_ (.CLK(clknet_leaf_357_clk),
    .RESET_B(net2703),
    .D(_02975_),
    .Q_N(_10530_),
    .Q(\atari2600.ram[36][1] ));
 sg13g2_dfrbp_1 _29410_ (.CLK(clknet_leaf_357_clk),
    .RESET_B(net2701),
    .D(_02976_),
    .Q_N(_10529_),
    .Q(\atari2600.ram[36][2] ));
 sg13g2_dfrbp_1 _29411_ (.CLK(clknet_leaf_357_clk),
    .RESET_B(net2699),
    .D(_02977_),
    .Q_N(_10528_),
    .Q(\atari2600.ram[36][3] ));
 sg13g2_dfrbp_1 _29412_ (.CLK(clknet_leaf_358_clk),
    .RESET_B(net2697),
    .D(_02978_),
    .Q_N(_10527_),
    .Q(\atari2600.ram[36][4] ));
 sg13g2_dfrbp_1 _29413_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net2695),
    .D(_02979_),
    .Q_N(_10526_),
    .Q(\atari2600.ram[36][5] ));
 sg13g2_dfrbp_1 _29414_ (.CLK(clknet_leaf_356_clk),
    .RESET_B(net2693),
    .D(_02980_),
    .Q_N(_10525_),
    .Q(\atari2600.ram[36][6] ));
 sg13g2_dfrbp_1 _29415_ (.CLK(clknet_leaf_357_clk),
    .RESET_B(net2691),
    .D(_02981_),
    .Q_N(_10524_),
    .Q(\atari2600.ram[36][7] ));
 sg13g2_dfrbp_1 _29416_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net2689),
    .D(net6174),
    .Q_N(_10523_),
    .Q(\atari2600.cpu.ABH[5] ));
 sg13g2_dfrbp_1 _29417_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net2687),
    .D(net7038),
    .Q_N(_10522_),
    .Q(\atari2600.cpu.ABH[6] ));
 sg13g2_dfrbp_1 _29418_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net274),
    .D(net6331),
    .Q_N(_10521_),
    .Q(\atari2600.cpu.ABH[7] ));
 sg13g2_dfrbp_1 _29419_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net270),
    .D(_02985_),
    .Q_N(_10520_),
    .Q(\atari2600.cpu.dst_reg[1] ));
 sg13g2_dfrbp_1 _29420_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net262),
    .D(_02986_),
    .Q_N(_10519_),
    .Q(\atari2600.cpu.dst_reg[0] ));
 sg13g2_dfrbp_1 _29421_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net254),
    .D(_02987_),
    .Q_N(_00081_),
    .Q(\atari2600.cpu.src_reg[1] ));
 sg13g2_dfrbp_1 _29422_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net230),
    .D(_02988_),
    .Q_N(_00080_),
    .Q(\atari2600.cpu.src_reg[0] ));
 sg13g2_dfrbp_1 _29423_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net222),
    .D(_02989_),
    .Q_N(_10518_),
    .Q(\atari2600.cpu.op[3] ));
 sg13g2_dfrbp_1 _29424_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net214),
    .D(_02990_),
    .Q_N(_10517_),
    .Q(\atari2600.cpu.op[2] ));
 sg13g2_dfrbp_1 _29425_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net258),
    .D(_02991_),
    .Q_N(_10516_),
    .Q(\atari2600.cpu.op[1] ));
 sg13g2_dfrbp_1 _29426_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net226),
    .D(_02992_),
    .Q_N(_10515_),
    .Q(\atari2600.cpu.op[0] ));
 sg13g2_dfrbp_1 _29427_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net266),
    .D(_02993_),
    .Q_N(_10514_),
    .Q(\atari2600.tia.dat_o[7] ));
 sg13g2_dfrbp_1 _29428_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net218),
    .D(net2957),
    .Q_N(_10513_),
    .Q(\atari2600.tia.dat_o[6] ));
 sg13g2_tiehi _28842__13 (.L_HI(net13));
 sg13g2_tiehi _28841__14 (.L_HI(net14));
 sg13g2_tiehi _28840__15 (.L_HI(net15));
 sg13g2_tiehi _28839__16 (.L_HI(net16));
 sg13g2_tiehi _28838__17 (.L_HI(net17));
 sg13g2_tiehi _28837__18 (.L_HI(net18));
 sg13g2_tiehi _28836__19 (.L_HI(net19));
 sg13g2_tiehi _28835__20 (.L_HI(net20));
 sg13g2_tiehi _28834__21 (.L_HI(net21));
 sg13g2_tiehi _28833__22 (.L_HI(net22));
 sg13g2_tiehi _28832__23 (.L_HI(net23));
 sg13g2_tiehi _28831__24 (.L_HI(net24));
 sg13g2_tiehi _28830__25 (.L_HI(net25));
 sg13g2_tiehi _28829__26 (.L_HI(net26));
 sg13g2_tiehi _28824__27 (.L_HI(net27));
 sg13g2_tiehi _28823__28 (.L_HI(net28));
 sg13g2_tiehi _28822__29 (.L_HI(net29));
 sg13g2_tiehi _28821__30 (.L_HI(net30));
 sg13g2_tiehi _28820__31 (.L_HI(net31));
 sg13g2_tiehi _28819__32 (.L_HI(net32));
 sg13g2_tiehi _28818__33 (.L_HI(net33));
 sg13g2_tiehi _28817__34 (.L_HI(net34));
 sg13g2_tiehi _28816__35 (.L_HI(net35));
 sg13g2_tiehi _28815__36 (.L_HI(net36));
 sg13g2_tiehi _28814__37 (.L_HI(net37));
 sg13g2_tiehi _28813__38 (.L_HI(net38));
 sg13g2_tiehi _28812__39 (.L_HI(net39));
 sg13g2_tiehi _28811__40 (.L_HI(net40));
 sg13g2_tiehi _28810__41 (.L_HI(net41));
 sg13g2_tiehi _29393__42 (.L_HI(net42));
 sg13g2_tiehi _28809__43 (.L_HI(net43));
 sg13g2_tiehi _29392__44 (.L_HI(net44));
 sg13g2_tiehi _28808__45 (.L_HI(net45));
 sg13g2_tiehi _29391__46 (.L_HI(net46));
 sg13g2_tiehi _28807__47 (.L_HI(net47));
 sg13g2_tiehi _29390__48 (.L_HI(net48));
 sg13g2_tiehi _28806__49 (.L_HI(net49));
 sg13g2_tiehi _29389__50 (.L_HI(net50));
 sg13g2_tiehi _28805__51 (.L_HI(net51));
 sg13g2_tiehi _29388__52 (.L_HI(net52));
 sg13g2_tiehi _28804__53 (.L_HI(net53));
 sg13g2_tiehi _29387__54 (.L_HI(net54));
 sg13g2_tiehi _28803__55 (.L_HI(net55));
 sg13g2_tiehi _29386__56 (.L_HI(net56));
 sg13g2_tiehi _28802__57 (.L_HI(net57));
 sg13g2_tiehi _29385__58 (.L_HI(net58));
 sg13g2_tiehi _28801__59 (.L_HI(net59));
 sg13g2_tiehi _29384__60 (.L_HI(net60));
 sg13g2_tiehi _28800__61 (.L_HI(net61));
 sg13g2_tiehi _29383__62 (.L_HI(net62));
 sg13g2_tiehi _28799__63 (.L_HI(net63));
 sg13g2_tiehi _29382__64 (.L_HI(net64));
 sg13g2_tiehi _28798__65 (.L_HI(net65));
 sg13g2_tiehi _28797__66 (.L_HI(net66));
 sg13g2_tiehi _28796__67 (.L_HI(net67));
 sg13g2_tiehi _28795__68 (.L_HI(net68));
 sg13g2_tiehi _28794__69 (.L_HI(net69));
 sg13g2_tiehi _28793__70 (.L_HI(net70));
 sg13g2_tiehi _28792__71 (.L_HI(net71));
 sg13g2_tiehi _28791__72 (.L_HI(net72));
 sg13g2_tiehi _28790__73 (.L_HI(net73));
 sg13g2_tiehi _28789__74 (.L_HI(net74));
 sg13g2_tiehi _28788__75 (.L_HI(net75));
 sg13g2_tiehi _28787__76 (.L_HI(net76));
 sg13g2_tiehi _28786__77 (.L_HI(net77));
 sg13g2_tiehi _28785__78 (.L_HI(net78));
 sg13g2_tiehi _28784__79 (.L_HI(net79));
 sg13g2_tiehi _28783__80 (.L_HI(net80));
 sg13g2_tiehi _28782__81 (.L_HI(net81));
 sg13g2_tiehi _28781__82 (.L_HI(net82));
 sg13g2_tiehi _28780__83 (.L_HI(net83));
 sg13g2_tiehi _28779__84 (.L_HI(net84));
 sg13g2_tiehi _28778__85 (.L_HI(net85));
 sg13g2_tiehi _28777__86 (.L_HI(net86));
 sg13g2_tiehi _28776__87 (.L_HI(net87));
 sg13g2_tiehi _28775__88 (.L_HI(net88));
 sg13g2_tiehi _28774__89 (.L_HI(net89));
 sg13g2_tiehi _28773__90 (.L_HI(net90));
 sg13g2_tiehi _28772__91 (.L_HI(net91));
 sg13g2_tiehi _28771__92 (.L_HI(net92));
 sg13g2_tiehi _28770__93 (.L_HI(net93));
 sg13g2_tiehi _28769__94 (.L_HI(net94));
 sg13g2_tiehi _28768__95 (.L_HI(net95));
 sg13g2_tiehi _28767__96 (.L_HI(net96));
 sg13g2_tiehi _28766__97 (.L_HI(net97));
 sg13g2_tiehi _28765__98 (.L_HI(net98));
 sg13g2_tiehi _28764__99 (.L_HI(net99));
 sg13g2_tiehi _28763__100 (.L_HI(net100));
 sg13g2_tiehi _28762__101 (.L_HI(net101));
 sg13g2_tiehi _28761__102 (.L_HI(net102));
 sg13g2_tiehi _28760__103 (.L_HI(net103));
 sg13g2_tiehi _28759__104 (.L_HI(net104));
 sg13g2_tiehi _28758__105 (.L_HI(net105));
 sg13g2_tiehi _28757__106 (.L_HI(net106));
 sg13g2_tiehi _28756__107 (.L_HI(net107));
 sg13g2_tiehi _28755__108 (.L_HI(net108));
 sg13g2_tiehi _28754__109 (.L_HI(net109));
 sg13g2_tiehi _28753__110 (.L_HI(net110));
 sg13g2_tiehi _28752__111 (.L_HI(net111));
 sg13g2_tiehi _28751__112 (.L_HI(net112));
 sg13g2_tiehi _28750__113 (.L_HI(net113));
 sg13g2_tiehi _28749__114 (.L_HI(net114));
 sg13g2_tiehi _28748__115 (.L_HI(net115));
 sg13g2_tiehi _28747__116 (.L_HI(net116));
 sg13g2_tiehi _28746__117 (.L_HI(net117));
 sg13g2_tiehi _28745__118 (.L_HI(net118));
 sg13g2_tiehi _28744__119 (.L_HI(net119));
 sg13g2_tiehi _28743__120 (.L_HI(net120));
 sg13g2_tiehi _28742__121 (.L_HI(net121));
 sg13g2_tiehi _28741__122 (.L_HI(net122));
 sg13g2_tiehi _28740__123 (.L_HI(net123));
 sg13g2_tiehi _28739__124 (.L_HI(net124));
 sg13g2_tiehi _28738__125 (.L_HI(net125));
 sg13g2_tiehi _28737__126 (.L_HI(net126));
 sg13g2_tiehi _28736__127 (.L_HI(net127));
 sg13g2_tiehi _28735__128 (.L_HI(net128));
 sg13g2_tiehi _28734__129 (.L_HI(net129));
 sg13g2_tiehi _28733__130 (.L_HI(net130));
 sg13g2_tiehi _28732__131 (.L_HI(net131));
 sg13g2_tiehi _28731__132 (.L_HI(net132));
 sg13g2_tiehi _28730__133 (.L_HI(net133));
 sg13g2_tiehi _28729__134 (.L_HI(net134));
 sg13g2_tiehi _28728__135 (.L_HI(net135));
 sg13g2_tiehi _28727__136 (.L_HI(net136));
 sg13g2_tiehi _28726__137 (.L_HI(net137));
 sg13g2_tiehi _28725__138 (.L_HI(net138));
 sg13g2_tiehi _28724__139 (.L_HI(net139));
 sg13g2_tiehi _28723__140 (.L_HI(net140));
 sg13g2_tiehi _28722__141 (.L_HI(net141));
 sg13g2_tiehi _28721__142 (.L_HI(net142));
 sg13g2_tiehi _28720__143 (.L_HI(net143));
 sg13g2_tiehi _28719__144 (.L_HI(net144));
 sg13g2_tiehi _28718__145 (.L_HI(net145));
 sg13g2_tiehi _28717__146 (.L_HI(net146));
 sg13g2_tiehi _28716__147 (.L_HI(net147));
 sg13g2_tiehi _28715__148 (.L_HI(net148));
 sg13g2_tiehi _28714__149 (.L_HI(net149));
 sg13g2_tiehi _28713__150 (.L_HI(net150));
 sg13g2_tiehi _28712__151 (.L_HI(net151));
 sg13g2_tiehi _28711__152 (.L_HI(net152));
 sg13g2_tiehi _28710__153 (.L_HI(net153));
 sg13g2_tiehi _28709__154 (.L_HI(net154));
 sg13g2_tiehi _28708__155 (.L_HI(net155));
 sg13g2_tiehi _28707__156 (.L_HI(net156));
 sg13g2_tiehi _28706__157 (.L_HI(net157));
 sg13g2_tiehi _28705__158 (.L_HI(net158));
 sg13g2_tiehi _28704__159 (.L_HI(net159));
 sg13g2_tiehi _28703__160 (.L_HI(net160));
 sg13g2_tiehi _28702__161 (.L_HI(net161));
 sg13g2_tiehi _28701__162 (.L_HI(net162));
 sg13g2_tiehi _28700__163 (.L_HI(net163));
 sg13g2_tiehi _28699__164 (.L_HI(net164));
 sg13g2_tiehi _28698__165 (.L_HI(net165));
 sg13g2_tiehi _28697__166 (.L_HI(net166));
 sg13g2_tiehi _28696__167 (.L_HI(net167));
 sg13g2_tiehi _28695__168 (.L_HI(net168));
 sg13g2_tiehi _28694__169 (.L_HI(net169));
 sg13g2_tiehi _28693__170 (.L_HI(net170));
 sg13g2_tiehi _28692__171 (.L_HI(net171));
 sg13g2_tiehi _28691__172 (.L_HI(net172));
 sg13g2_tiehi _28690__173 (.L_HI(net173));
 sg13g2_tiehi _28689__174 (.L_HI(net174));
 sg13g2_tiehi _28688__175 (.L_HI(net175));
 sg13g2_tiehi _28687__176 (.L_HI(net176));
 sg13g2_tiehi _28686__177 (.L_HI(net177));
 sg13g2_tiehi _28685__178 (.L_HI(net178));
 sg13g2_tiehi _28684__179 (.L_HI(net179));
 sg13g2_tiehi _28683__180 (.L_HI(net180));
 sg13g2_tiehi _28682__181 (.L_HI(net181));
 sg13g2_tiehi _28681__182 (.L_HI(net182));
 sg13g2_tiehi _28680__183 (.L_HI(net183));
 sg13g2_tiehi _28679__184 (.L_HI(net184));
 sg13g2_tiehi _28678__185 (.L_HI(net185));
 sg13g2_tiehi _29381__186 (.L_HI(net186));
 sg13g2_tiehi _28677__187 (.L_HI(net187));
 sg13g2_tiehi _29380__188 (.L_HI(net188));
 sg13g2_tiehi _28676__189 (.L_HI(net189));
 sg13g2_tiehi _29379__190 (.L_HI(net190));
 sg13g2_tiehi _28675__191 (.L_HI(net191));
 sg13g2_tiehi _29378__192 (.L_HI(net192));
 sg13g2_tiehi _28674__193 (.L_HI(net193));
 sg13g2_tiehi _29377__194 (.L_HI(net194));
 sg13g2_tiehi _28673__195 (.L_HI(net195));
 sg13g2_tiehi _29376__196 (.L_HI(net196));
 sg13g2_tiehi _28672__197 (.L_HI(net197));
 sg13g2_tiehi _29375__198 (.L_HI(net198));
 sg13g2_tiehi _28671__199 (.L_HI(net199));
 sg13g2_tiehi _29374__200 (.L_HI(net200));
 sg13g2_tiehi _28670__201 (.L_HI(net201));
 sg13g2_tiehi _29373__202 (.L_HI(net202));
 sg13g2_tiehi _28669__203 (.L_HI(net203));
 sg13g2_tiehi _29372__204 (.L_HI(net204));
 sg13g2_tiehi _28668__205 (.L_HI(net205));
 sg13g2_tiehi _29371__206 (.L_HI(net206));
 sg13g2_tiehi _28667__207 (.L_HI(net207));
 sg13g2_tiehi _29370__208 (.L_HI(net208));
 sg13g2_tiehi _28666__209 (.L_HI(net209));
 sg13g2_tiehi _29369__210 (.L_HI(net210));
 sg13g2_tiehi _28665__211 (.L_HI(net211));
 sg13g2_tiehi _29368__212 (.L_HI(net212));
 sg13g2_tiehi _28664__213 (.L_HI(net213));
 sg13g2_tiehi _29424__214 (.L_HI(net214));
 sg13g2_tiehi _28663__215 (.L_HI(net215));
 sg13g2_tiehi _29367__216 (.L_HI(net216));
 sg13g2_tiehi _28662__217 (.L_HI(net217));
 sg13g2_tiehi _29428__218 (.L_HI(net218));
 sg13g2_tiehi _28661__219 (.L_HI(net219));
 sg13g2_tiehi _29366__220 (.L_HI(net220));
 sg13g2_tiehi _28660__221 (.L_HI(net221));
 sg13g2_tiehi _29423__222 (.L_HI(net222));
 sg13g2_tiehi _28659__223 (.L_HI(net223));
 sg13g2_tiehi _29365__224 (.L_HI(net224));
 sg13g2_tiehi _28658__225 (.L_HI(net225));
 sg13g2_tiehi _29426__226 (.L_HI(net226));
 sg13g2_tiehi _28657__227 (.L_HI(net227));
 sg13g2_tiehi _29364__228 (.L_HI(net228));
 sg13g2_tiehi _28656__229 (.L_HI(net229));
 sg13g2_tiehi _29422__230 (.L_HI(net230));
 sg13g2_tiehi _28655__231 (.L_HI(net231));
 sg13g2_tiehi _29363__232 (.L_HI(net232));
 sg13g2_tiehi _28654__233 (.L_HI(net233));
 sg13g2_tiehi _29028__234 (.L_HI(net234));
 sg13g2_tiehi _28653__235 (.L_HI(net235));
 sg13g2_tiehi _29362__236 (.L_HI(net236));
 sg13g2_tiehi _28652__237 (.L_HI(net237));
 sg13g2_tiehi _29361__238 (.L_HI(net238));
 sg13g2_tiehi _28651__239 (.L_HI(net239));
 sg13g2_tiehi _29360__240 (.L_HI(net240));
 sg13g2_tiehi _28650__241 (.L_HI(net241));
 sg13g2_tiehi _29359__242 (.L_HI(net242));
 sg13g2_tiehi _28649__243 (.L_HI(net243));
 sg13g2_tiehi _29358__244 (.L_HI(net244));
 sg13g2_tiehi _28648__245 (.L_HI(net245));
 sg13g2_tiehi _29357__246 (.L_HI(net246));
 sg13g2_tiehi _28647__247 (.L_HI(net247));
 sg13g2_tiehi _29356__248 (.L_HI(net248));
 sg13g2_tiehi _28646__249 (.L_HI(net249));
 sg13g2_tiehi _29355__250 (.L_HI(net250));
 sg13g2_tiehi _28645__251 (.L_HI(net251));
 sg13g2_tiehi _29354__252 (.L_HI(net252));
 sg13g2_tiehi _28644__253 (.L_HI(net253));
 sg13g2_tiehi _29421__254 (.L_HI(net254));
 sg13g2_tiehi _28643__255 (.L_HI(net255));
 sg13g2_tiehi _29353__256 (.L_HI(net256));
 sg13g2_tiehi _28642__257 (.L_HI(net257));
 sg13g2_tiehi _29425__258 (.L_HI(net258));
 sg13g2_tiehi _28641__259 (.L_HI(net259));
 sg13g2_tiehi _29352__260 (.L_HI(net260));
 sg13g2_tiehi _28640__261 (.L_HI(net261));
 sg13g2_tiehi _29420__262 (.L_HI(net262));
 sg13g2_tiehi _28639__263 (.L_HI(net263));
 sg13g2_tiehi _29351__264 (.L_HI(net264));
 sg13g2_tiehi _28638__265 (.L_HI(net265));
 sg13g2_tiehi _29427__266 (.L_HI(net266));
 sg13g2_tiehi _28637__267 (.L_HI(net267));
 sg13g2_tiehi _29350__268 (.L_HI(net268));
 sg13g2_tiehi _28636__269 (.L_HI(net269));
 sg13g2_tiehi _29419__270 (.L_HI(net270));
 sg13g2_tiehi _28635__271 (.L_HI(net271));
 sg13g2_tiehi _29349__272 (.L_HI(net272));
 sg13g2_tiehi _28634__273 (.L_HI(net273));
 sg13g2_tiehi _29418__274 (.L_HI(net274));
 sg13g2_tiehi _28633__275 (.L_HI(net275));
 sg13g2_tiehi _29348__276 (.L_HI(net276));
 sg13g2_tiehi _28632__277 (.L_HI(net277));
 sg13g2_tiehi _29347__278 (.L_HI(net278));
 sg13g2_tiehi _28631__279 (.L_HI(net279));
 sg13g2_tiehi _29346__280 (.L_HI(net280));
 sg13g2_tiehi _28630__281 (.L_HI(net281));
 sg13g2_tiehi _29345__282 (.L_HI(net282));
 sg13g2_tiehi _28629__283 (.L_HI(net283));
 sg13g2_tiehi _29344__284 (.L_HI(net284));
 sg13g2_tiehi _28628__285 (.L_HI(net285));
 sg13g2_tiehi _29343__286 (.L_HI(net286));
 sg13g2_tiehi _28627__287 (.L_HI(net287));
 sg13g2_tiehi _29342__288 (.L_HI(net288));
 sg13g2_tiehi _28626__289 (.L_HI(net289));
 sg13g2_tiehi _29341__290 (.L_HI(net290));
 sg13g2_tiehi _28625__291 (.L_HI(net291));
 sg13g2_tiehi _29340__292 (.L_HI(net292));
 sg13g2_tiehi _28624__293 (.L_HI(net293));
 sg13g2_tiehi _29339__294 (.L_HI(net294));
 sg13g2_tiehi _28623__295 (.L_HI(net295));
 sg13g2_tiehi _29338__296 (.L_HI(net296));
 sg13g2_tiehi _28622__297 (.L_HI(net297));
 sg13g2_tiehi _29337__298 (.L_HI(net298));
 sg13g2_tiehi _28621__299 (.L_HI(net299));
 sg13g2_tiehi _29336__300 (.L_HI(net300));
 sg13g2_tiehi _28620__301 (.L_HI(net301));
 sg13g2_tiehi _29335__302 (.L_HI(net302));
 sg13g2_tiehi _28619__303 (.L_HI(net303));
 sg13g2_tiehi _29334__304 (.L_HI(net304));
 sg13g2_tiehi _28618__305 (.L_HI(net305));
 sg13g2_tiehi _29333__306 (.L_HI(net306));
 sg13g2_tiehi _28617__307 (.L_HI(net307));
 sg13g2_tiehi _29332__308 (.L_HI(net308));
 sg13g2_tiehi _28616__309 (.L_HI(net309));
 sg13g2_tiehi _29331__310 (.L_HI(net310));
 sg13g2_tiehi _28615__311 (.L_HI(net311));
 sg13g2_tiehi _29330__312 (.L_HI(net312));
 sg13g2_tiehi _28614__313 (.L_HI(net313));
 sg13g2_tiehi _29329__314 (.L_HI(net314));
 sg13g2_tiehi _28598__315 (.L_HI(net315));
 sg13g2_tiehi _29328__316 (.L_HI(net316));
 sg13g2_tiehi _28597__317 (.L_HI(net317));
 sg13g2_tiehi _29327__318 (.L_HI(net318));
 sg13g2_tiehi _28596__319 (.L_HI(net319));
 sg13g2_tiehi _29326__320 (.L_HI(net320));
 sg13g2_tiehi _28595__321 (.L_HI(net321));
 sg13g2_tiehi _29325__322 (.L_HI(net322));
 sg13g2_tiehi _28594__323 (.L_HI(net323));
 sg13g2_tiehi _29324__324 (.L_HI(net324));
 sg13g2_tiehi _28593__325 (.L_HI(net325));
 sg13g2_tiehi _29323__326 (.L_HI(net326));
 sg13g2_tiehi _28592__327 (.L_HI(net327));
 sg13g2_tiehi _29322__328 (.L_HI(net328));
 sg13g2_tiehi _28591__329 (.L_HI(net329));
 sg13g2_tiehi _29321__330 (.L_HI(net330));
 sg13g2_tiehi _28590__331 (.L_HI(net331));
 sg13g2_tiehi _29320__332 (.L_HI(net332));
 sg13g2_tiehi _28589__333 (.L_HI(net333));
 sg13g2_tiehi _29319__334 (.L_HI(net334));
 sg13g2_tiehi _28588__335 (.L_HI(net335));
 sg13g2_tiehi _29318__336 (.L_HI(net336));
 sg13g2_tiehi _28587__337 (.L_HI(net337));
 sg13g2_tiehi _29317__338 (.L_HI(net338));
 sg13g2_tiehi _28586__339 (.L_HI(net339));
 sg13g2_tiehi _29316__340 (.L_HI(net340));
 sg13g2_tiehi _28585__341 (.L_HI(net341));
 sg13g2_tiehi _29315__342 (.L_HI(net342));
 sg13g2_tiehi _28584__343 (.L_HI(net343));
 sg13g2_tiehi _29314__344 (.L_HI(net344));
 sg13g2_tiehi _28583__345 (.L_HI(net345));
 sg13g2_tiehi _29313__346 (.L_HI(net346));
 sg13g2_tiehi _28582__347 (.L_HI(net347));
 sg13g2_tiehi _29312__348 (.L_HI(net348));
 sg13g2_tiehi _28581__349 (.L_HI(net349));
 sg13g2_tiehi _29311__350 (.L_HI(net350));
 sg13g2_tiehi _28580__351 (.L_HI(net351));
 sg13g2_tiehi _29310__352 (.L_HI(net352));
 sg13g2_tiehi _28579__353 (.L_HI(net353));
 sg13g2_tiehi _29309__354 (.L_HI(net354));
 sg13g2_tiehi _28578__355 (.L_HI(net355));
 sg13g2_tiehi _29308__356 (.L_HI(net356));
 sg13g2_tiehi _28577__357 (.L_HI(net357));
 sg13g2_tiehi _29307__358 (.L_HI(net358));
 sg13g2_tiehi _28576__359 (.L_HI(net359));
 sg13g2_tiehi _29306__360 (.L_HI(net360));
 sg13g2_tiehi _28575__361 (.L_HI(net361));
 sg13g2_tiehi _29305__362 (.L_HI(net362));
 sg13g2_tiehi _28574__363 (.L_HI(net363));
 sg13g2_tiehi _29304__364 (.L_HI(net364));
 sg13g2_tiehi _28573__365 (.L_HI(net365));
 sg13g2_tiehi _29303__366 (.L_HI(net366));
 sg13g2_tiehi _28572__367 (.L_HI(net367));
 sg13g2_tiehi _29302__368 (.L_HI(net368));
 sg13g2_tiehi _28571__369 (.L_HI(net369));
 sg13g2_tiehi _29301__370 (.L_HI(net370));
 sg13g2_tiehi _28570__371 (.L_HI(net371));
 sg13g2_tiehi _29300__372 (.L_HI(net372));
 sg13g2_tiehi _28569__373 (.L_HI(net373));
 sg13g2_tiehi _29299__374 (.L_HI(net374));
 sg13g2_tiehi _28568__375 (.L_HI(net375));
 sg13g2_tiehi _29298__376 (.L_HI(net376));
 sg13g2_tiehi _28567__377 (.L_HI(net377));
 sg13g2_tiehi _29297__378 (.L_HI(net378));
 sg13g2_tiehi _28566__379 (.L_HI(net379));
 sg13g2_tiehi _29296__380 (.L_HI(net380));
 sg13g2_tiehi _28565__381 (.L_HI(net381));
 sg13g2_tiehi _29295__382 (.L_HI(net382));
 sg13g2_tiehi _28564__383 (.L_HI(net383));
 sg13g2_tiehi _29294__384 (.L_HI(net384));
 sg13g2_tiehi _28563__385 (.L_HI(net385));
 sg13g2_tiehi _29293__386 (.L_HI(net386));
 sg13g2_tiehi _28562__387 (.L_HI(net387));
 sg13g2_tiehi _29292__388 (.L_HI(net388));
 sg13g2_tiehi _28561__389 (.L_HI(net389));
 sg13g2_tiehi _29291__390 (.L_HI(net390));
 sg13g2_tiehi _28560__391 (.L_HI(net391));
 sg13g2_tiehi _29290__392 (.L_HI(net392));
 sg13g2_tiehi _28559__393 (.L_HI(net393));
 sg13g2_tiehi _29289__394 (.L_HI(net394));
 sg13g2_tiehi _28558__395 (.L_HI(net395));
 sg13g2_tiehi _29288__396 (.L_HI(net396));
 sg13g2_tiehi _28557__397 (.L_HI(net397));
 sg13g2_tiehi _29287__398 (.L_HI(net398));
 sg13g2_tiehi _28556__399 (.L_HI(net399));
 sg13g2_tiehi _29286__400 (.L_HI(net400));
 sg13g2_tiehi _28555__401 (.L_HI(net401));
 sg13g2_tiehi _29285__402 (.L_HI(net402));
 sg13g2_tiehi _28554__403 (.L_HI(net403));
 sg13g2_tiehi _29284__404 (.L_HI(net404));
 sg13g2_tiehi _28553__405 (.L_HI(net405));
 sg13g2_tiehi _29283__406 (.L_HI(net406));
 sg13g2_tiehi _28552__407 (.L_HI(net407));
 sg13g2_tiehi _29282__408 (.L_HI(net408));
 sg13g2_tiehi _28551__409 (.L_HI(net409));
 sg13g2_tiehi _29281__410 (.L_HI(net410));
 sg13g2_tiehi _28550__411 (.L_HI(net411));
 sg13g2_tiehi _29280__412 (.L_HI(net412));
 sg13g2_tiehi _28549__413 (.L_HI(net413));
 sg13g2_tiehi _29279__414 (.L_HI(net414));
 sg13g2_tiehi _28548__415 (.L_HI(net415));
 sg13g2_tiehi _29278__416 (.L_HI(net416));
 sg13g2_tiehi _28547__417 (.L_HI(net417));
 sg13g2_tiehi _29277__418 (.L_HI(net418));
 sg13g2_tiehi _28546__419 (.L_HI(net419));
 sg13g2_tiehi _29276__420 (.L_HI(net420));
 sg13g2_tiehi _28545__421 (.L_HI(net421));
 sg13g2_tiehi _29275__422 (.L_HI(net422));
 sg13g2_tiehi _28544__423 (.L_HI(net423));
 sg13g2_tiehi _29274__424 (.L_HI(net424));
 sg13g2_tiehi _28543__425 (.L_HI(net425));
 sg13g2_tiehi _29273__426 (.L_HI(net426));
 sg13g2_tiehi _28542__427 (.L_HI(net427));
 sg13g2_tiehi _29272__428 (.L_HI(net428));
 sg13g2_tiehi _28541__429 (.L_HI(net429));
 sg13g2_tiehi _29271__430 (.L_HI(net430));
 sg13g2_tiehi _28540__431 (.L_HI(net431));
 sg13g2_tiehi _29270__432 (.L_HI(net432));
 sg13g2_tiehi _28539__433 (.L_HI(net433));
 sg13g2_tiehi _29269__434 (.L_HI(net434));
 sg13g2_tiehi _28538__435 (.L_HI(net435));
 sg13g2_tiehi _29268__436 (.L_HI(net436));
 sg13g2_tiehi _28537__437 (.L_HI(net437));
 sg13g2_tiehi _29267__438 (.L_HI(net438));
 sg13g2_tiehi _28536__439 (.L_HI(net439));
 sg13g2_tiehi _29266__440 (.L_HI(net440));
 sg13g2_tiehi _28535__441 (.L_HI(net441));
 sg13g2_tiehi _29265__442 (.L_HI(net442));
 sg13g2_tiehi _28534__443 (.L_HI(net443));
 sg13g2_tiehi _29264__444 (.L_HI(net444));
 sg13g2_tiehi _28533__445 (.L_HI(net445));
 sg13g2_tiehi _29263__446 (.L_HI(net446));
 sg13g2_tiehi _28532__447 (.L_HI(net447));
 sg13g2_tiehi _28531__448 (.L_HI(net448));
 sg13g2_tiehi _28530__449 (.L_HI(net449));
 sg13g2_tiehi _28529__450 (.L_HI(net450));
 sg13g2_tiehi _28528__451 (.L_HI(net451));
 sg13g2_tiehi _28527__452 (.L_HI(net452));
 sg13g2_tiehi _28526__453 (.L_HI(net453));
 sg13g2_tiehi _28525__454 (.L_HI(net454));
 sg13g2_tiehi _28524__455 (.L_HI(net455));
 sg13g2_tiehi _28523__456 (.L_HI(net456));
 sg13g2_tiehi _28522__457 (.L_HI(net457));
 sg13g2_tiehi _28521__458 (.L_HI(net458));
 sg13g2_tiehi _28520__459 (.L_HI(net459));
 sg13g2_tiehi _28519__460 (.L_HI(net460));
 sg13g2_tiehi _28518__461 (.L_HI(net461));
 sg13g2_tiehi _28517__462 (.L_HI(net462));
 sg13g2_tiehi _29262__463 (.L_HI(net463));
 sg13g2_tiehi _28516__464 (.L_HI(net464));
 sg13g2_tiehi _29261__465 (.L_HI(net465));
 sg13g2_tiehi _28515__466 (.L_HI(net466));
 sg13g2_tiehi _29260__467 (.L_HI(net467));
 sg13g2_tiehi _28514__468 (.L_HI(net468));
 sg13g2_tiehi _29259__469 (.L_HI(net469));
 sg13g2_tiehi _28513__470 (.L_HI(net470));
 sg13g2_tiehi _29258__471 (.L_HI(net471));
 sg13g2_tiehi _28512__472 (.L_HI(net472));
 sg13g2_tiehi _29257__473 (.L_HI(net473));
 sg13g2_tiehi _28511__474 (.L_HI(net474));
 sg13g2_tiehi _29256__475 (.L_HI(net475));
 sg13g2_tiehi _28510__476 (.L_HI(net476));
 sg13g2_tiehi _29255__477 (.L_HI(net477));
 sg13g2_tiehi _28509__478 (.L_HI(net478));
 sg13g2_tiehi _29254__479 (.L_HI(net479));
 sg13g2_tiehi _28508__480 (.L_HI(net480));
 sg13g2_tiehi _29253__481 (.L_HI(net481));
 sg13g2_tiehi _28507__482 (.L_HI(net482));
 sg13g2_tiehi _29252__483 (.L_HI(net483));
 sg13g2_tiehi _28506__484 (.L_HI(net484));
 sg13g2_tiehi _29251__485 (.L_HI(net485));
 sg13g2_tiehi _28505__486 (.L_HI(net486));
 sg13g2_tiehi _29250__487 (.L_HI(net487));
 sg13g2_tiehi _28504__488 (.L_HI(net488));
 sg13g2_tiehi _29249__489 (.L_HI(net489));
 sg13g2_tiehi _28503__490 (.L_HI(net490));
 sg13g2_tiehi _29248__491 (.L_HI(net491));
 sg13g2_tiehi _28502__492 (.L_HI(net492));
 sg13g2_tiehi _29247__493 (.L_HI(net493));
 sg13g2_tiehi _28501__494 (.L_HI(net494));
 sg13g2_tiehi _29246__495 (.L_HI(net495));
 sg13g2_tiehi _28500__496 (.L_HI(net496));
 sg13g2_tiehi _29245__497 (.L_HI(net497));
 sg13g2_tiehi _28499__498 (.L_HI(net498));
 sg13g2_tiehi _29244__499 (.L_HI(net499));
 sg13g2_tiehi _28498__500 (.L_HI(net500));
 sg13g2_tiehi _29243__501 (.L_HI(net501));
 sg13g2_tiehi _28497__502 (.L_HI(net502));
 sg13g2_tiehi _29242__503 (.L_HI(net503));
 sg13g2_tiehi _28496__504 (.L_HI(net504));
 sg13g2_tiehi _29241__505 (.L_HI(net505));
 sg13g2_tiehi _28495__506 (.L_HI(net506));
 sg13g2_tiehi _29240__507 (.L_HI(net507));
 sg13g2_tiehi _28494__508 (.L_HI(net508));
 sg13g2_tiehi _28493__509 (.L_HI(net509));
 sg13g2_tiehi _28492__510 (.L_HI(net510));
 sg13g2_tiehi _28491__511 (.L_HI(net511));
 sg13g2_tiehi _28490__512 (.L_HI(net512));
 sg13g2_tiehi _28489__513 (.L_HI(net513));
 sg13g2_tiehi _28488__514 (.L_HI(net514));
 sg13g2_tiehi _28487__515 (.L_HI(net515));
 sg13g2_tiehi _29239__516 (.L_HI(net516));
 sg13g2_tiehi _28486__517 (.L_HI(net517));
 sg13g2_tiehi _29238__518 (.L_HI(net518));
 sg13g2_tiehi _28485__519 (.L_HI(net519));
 sg13g2_tiehi _29237__520 (.L_HI(net520));
 sg13g2_tiehi _28484__521 (.L_HI(net521));
 sg13g2_tiehi _29236__522 (.L_HI(net522));
 sg13g2_tiehi _28483__523 (.L_HI(net523));
 sg13g2_tiehi _29235__524 (.L_HI(net524));
 sg13g2_tiehi _28482__525 (.L_HI(net525));
 sg13g2_tiehi _29234__526 (.L_HI(net526));
 sg13g2_tiehi _28481__527 (.L_HI(net527));
 sg13g2_tiehi _29233__528 (.L_HI(net528));
 sg13g2_tiehi _28480__529 (.L_HI(net529));
 sg13g2_tiehi _29232__530 (.L_HI(net530));
 sg13g2_tiehi _28479__531 (.L_HI(net531));
 sg13g2_tiehi _29231__532 (.L_HI(net532));
 sg13g2_tiehi _28478__533 (.L_HI(net533));
 sg13g2_tiehi _29230__534 (.L_HI(net534));
 sg13g2_tiehi _28477__535 (.L_HI(net535));
 sg13g2_tiehi _29229__536 (.L_HI(net536));
 sg13g2_tiehi _28476__537 (.L_HI(net537));
 sg13g2_tiehi _29228__538 (.L_HI(net538));
 sg13g2_tiehi _28475__539 (.L_HI(net539));
 sg13g2_tiehi _29227__540 (.L_HI(net540));
 sg13g2_tiehi _28474__541 (.L_HI(net541));
 sg13g2_tiehi _29226__542 (.L_HI(net542));
 sg13g2_tiehi _28473__543 (.L_HI(net543));
 sg13g2_tiehi _29225__544 (.L_HI(net544));
 sg13g2_tiehi _28472__545 (.L_HI(net545));
 sg13g2_tiehi _29224__546 (.L_HI(net546));
 sg13g2_tiehi _28471__547 (.L_HI(net547));
 sg13g2_tiehi _29223__548 (.L_HI(net548));
 sg13g2_tiehi _28470__549 (.L_HI(net549));
 sg13g2_tiehi _29222__550 (.L_HI(net550));
 sg13g2_tiehi _28469__551 (.L_HI(net551));
 sg13g2_tiehi _29221__552 (.L_HI(net552));
 sg13g2_tiehi _28468__553 (.L_HI(net553));
 sg13g2_tiehi _29220__554 (.L_HI(net554));
 sg13g2_tiehi _28467__555 (.L_HI(net555));
 sg13g2_tiehi _29219__556 (.L_HI(net556));
 sg13g2_tiehi _28466__557 (.L_HI(net557));
 sg13g2_tiehi _29218__558 (.L_HI(net558));
 sg13g2_tiehi _28465__559 (.L_HI(net559));
 sg13g2_tiehi _29217__560 (.L_HI(net560));
 sg13g2_tiehi _28464__561 (.L_HI(net561));
 sg13g2_tiehi _29216__562 (.L_HI(net562));
 sg13g2_tiehi _28463__563 (.L_HI(net563));
 sg13g2_tiehi _29215__564 (.L_HI(net564));
 sg13g2_tiehi _28462__565 (.L_HI(net565));
 sg13g2_tiehi _29214__566 (.L_HI(net566));
 sg13g2_tiehi _28461__567 (.L_HI(net567));
 sg13g2_tiehi _29213__568 (.L_HI(net568));
 sg13g2_tiehi _28460__569 (.L_HI(net569));
 sg13g2_tiehi _29212__570 (.L_HI(net570));
 sg13g2_tiehi _28459__571 (.L_HI(net571));
 sg13g2_tiehi _29211__572 (.L_HI(net572));
 sg13g2_tiehi _28458__573 (.L_HI(net573));
 sg13g2_tiehi _29210__574 (.L_HI(net574));
 sg13g2_tiehi _28457__575 (.L_HI(net575));
 sg13g2_tiehi _29209__576 (.L_HI(net576));
 sg13g2_tiehi _28456__577 (.L_HI(net577));
 sg13g2_tiehi _28455__578 (.L_HI(net578));
 sg13g2_tiehi _28454__579 (.L_HI(net579));
 sg13g2_tiehi _28453__580 (.L_HI(net580));
 sg13g2_tiehi _29208__581 (.L_HI(net581));
 sg13g2_tiehi _28452__582 (.L_HI(net582));
 sg13g2_tiehi _29207__583 (.L_HI(net583));
 sg13g2_tiehi _28451__584 (.L_HI(net584));
 sg13g2_tiehi _29206__585 (.L_HI(net585));
 sg13g2_tiehi _28450__586 (.L_HI(net586));
 sg13g2_tiehi _29205__587 (.L_HI(net587));
 sg13g2_tiehi _28432__588 (.L_HI(net588));
 sg13g2_tiehi _29204__589 (.L_HI(net589));
 sg13g2_tiehi _28431__590 (.L_HI(net590));
 sg13g2_tiehi _29203__591 (.L_HI(net591));
 sg13g2_tiehi _28430__592 (.L_HI(net592));
 sg13g2_tiehi _29202__593 (.L_HI(net593));
 sg13g2_tiehi _28429__594 (.L_HI(net594));
 sg13g2_tiehi _29201__595 (.L_HI(net595));
 sg13g2_tiehi _28428__596 (.L_HI(net596));
 sg13g2_tiehi _29200__597 (.L_HI(net597));
 sg13g2_tiehi _28427__598 (.L_HI(net598));
 sg13g2_tiehi _29199__599 (.L_HI(net599));
 sg13g2_tiehi _28426__600 (.L_HI(net600));
 sg13g2_tiehi _29198__601 (.L_HI(net601));
 sg13g2_tiehi _28425__602 (.L_HI(net602));
 sg13g2_tiehi _29197__603 (.L_HI(net603));
 sg13g2_tiehi _28424__604 (.L_HI(net604));
 sg13g2_tiehi _29196__605 (.L_HI(net605));
 sg13g2_tiehi _28423__606 (.L_HI(net606));
 sg13g2_tiehi _29195__607 (.L_HI(net607));
 sg13g2_tiehi _28422__608 (.L_HI(net608));
 sg13g2_tiehi _29194__609 (.L_HI(net609));
 sg13g2_tiehi _28421__610 (.L_HI(net610));
 sg13g2_tiehi _29193__611 (.L_HI(net611));
 sg13g2_tiehi _28420__612 (.L_HI(net612));
 sg13g2_tiehi _29192__613 (.L_HI(net613));
 sg13g2_tiehi _28419__614 (.L_HI(net614));
 sg13g2_tiehi _29191__615 (.L_HI(net615));
 sg13g2_tiehi _28418__616 (.L_HI(net616));
 sg13g2_tiehi _29190__617 (.L_HI(net617));
 sg13g2_tiehi _28417__618 (.L_HI(net618));
 sg13g2_tiehi _29189__619 (.L_HI(net619));
 sg13g2_tiehi _28416__620 (.L_HI(net620));
 sg13g2_tiehi _29188__621 (.L_HI(net621));
 sg13g2_tiehi _28415__622 (.L_HI(net622));
 sg13g2_tiehi _29187__623 (.L_HI(net623));
 sg13g2_tiehi _28414__624 (.L_HI(net624));
 sg13g2_tiehi _29186__625 (.L_HI(net625));
 sg13g2_tiehi _28413__626 (.L_HI(net626));
 sg13g2_tiehi _29185__627 (.L_HI(net627));
 sg13g2_tiehi _28412__628 (.L_HI(net628));
 sg13g2_tiehi _29184__629 (.L_HI(net629));
 sg13g2_tiehi _28411__630 (.L_HI(net630));
 sg13g2_tiehi _29183__631 (.L_HI(net631));
 sg13g2_tiehi _28410__632 (.L_HI(net632));
 sg13g2_tiehi _29182__633 (.L_HI(net633));
 sg13g2_tiehi _28409__634 (.L_HI(net634));
 sg13g2_tiehi _29181__635 (.L_HI(net635));
 sg13g2_tiehi _28408__636 (.L_HI(net636));
 sg13g2_tiehi _29180__637 (.L_HI(net637));
 sg13g2_tiehi _28407__638 (.L_HI(net638));
 sg13g2_tiehi _29179__639 (.L_HI(net639));
 sg13g2_tiehi _28406__640 (.L_HI(net640));
 sg13g2_tiehi _29178__641 (.L_HI(net641));
 sg13g2_tiehi _28405__642 (.L_HI(net642));
 sg13g2_tiehi _29177__643 (.L_HI(net643));
 sg13g2_tiehi _28404__644 (.L_HI(net644));
 sg13g2_tiehi _29176__645 (.L_HI(net645));
 sg13g2_tiehi _28403__646 (.L_HI(net646));
 sg13g2_tiehi _29175__647 (.L_HI(net647));
 sg13g2_tiehi _28402__648 (.L_HI(net648));
 sg13g2_tiehi _29174__649 (.L_HI(net649));
 sg13g2_tiehi _28401__650 (.L_HI(net650));
 sg13g2_tiehi _29173__651 (.L_HI(net651));
 sg13g2_tiehi _28400__652 (.L_HI(net652));
 sg13g2_tiehi _29172__653 (.L_HI(net653));
 sg13g2_tiehi _28399__654 (.L_HI(net654));
 sg13g2_tiehi _28398__655 (.L_HI(net655));
 sg13g2_tiehi _28397__656 (.L_HI(net656));
 sg13g2_tiehi _28396__657 (.L_HI(net657));
 sg13g2_tiehi _28395__658 (.L_HI(net658));
 sg13g2_tiehi _28394__659 (.L_HI(net659));
 sg13g2_tiehi _28393__660 (.L_HI(net660));
 sg13g2_tiehi _28392__661 (.L_HI(net661));
 sg13g2_tiehi _28391__662 (.L_HI(net662));
 sg13g2_tiehi _28390__663 (.L_HI(net663));
 sg13g2_tiehi _28389__664 (.L_HI(net664));
 sg13g2_tiehi _28388__665 (.L_HI(net665));
 sg13g2_tiehi _28387__666 (.L_HI(net666));
 sg13g2_tiehi _28386__667 (.L_HI(net667));
 sg13g2_tiehi _28385__668 (.L_HI(net668));
 sg13g2_tiehi _28384__669 (.L_HI(net669));
 sg13g2_tiehi _28383__670 (.L_HI(net670));
 sg13g2_tiehi _28382__671 (.L_HI(net671));
 sg13g2_tiehi _28381__672 (.L_HI(net672));
 sg13g2_tiehi _28380__673 (.L_HI(net673));
 sg13g2_tiehi _28379__674 (.L_HI(net674));
 sg13g2_tiehi _28378__675 (.L_HI(net675));
 sg13g2_tiehi _28377__676 (.L_HI(net676));
 sg13g2_tiehi _28376__677 (.L_HI(net677));
 sg13g2_tiehi _28375__678 (.L_HI(net678));
 sg13g2_tiehi _28374__679 (.L_HI(net679));
 sg13g2_tiehi _28373__680 (.L_HI(net680));
 sg13g2_tiehi _28372__681 (.L_HI(net681));
 sg13g2_tiehi _28371__682 (.L_HI(net682));
 sg13g2_tiehi _28370__683 (.L_HI(net683));
 sg13g2_tiehi _28369__684 (.L_HI(net684));
 sg13g2_tiehi _28368__685 (.L_HI(net685));
 sg13g2_tiehi _28367__686 (.L_HI(net686));
 sg13g2_tiehi _28366__687 (.L_HI(net687));
 sg13g2_tiehi _28365__688 (.L_HI(net688));
 sg13g2_tiehi _28364__689 (.L_HI(net689));
 sg13g2_tiehi _28363__690 (.L_HI(net690));
 sg13g2_tiehi _28362__691 (.L_HI(net691));
 sg13g2_tiehi _28361__692 (.L_HI(net692));
 sg13g2_tiehi _28360__693 (.L_HI(net693));
 sg13g2_tiehi _28359__694 (.L_HI(net694));
 sg13g2_tiehi _28358__695 (.L_HI(net695));
 sg13g2_tiehi _28357__696 (.L_HI(net696));
 sg13g2_tiehi _28356__697 (.L_HI(net697));
 sg13g2_tiehi _28355__698 (.L_HI(net698));
 sg13g2_tiehi _28354__699 (.L_HI(net699));
 sg13g2_tiehi _28353__700 (.L_HI(net700));
 sg13g2_tiehi _28352__701 (.L_HI(net701));
 sg13g2_tiehi _28351__702 (.L_HI(net702));
 sg13g2_tiehi _28350__703 (.L_HI(net703));
 sg13g2_tiehi _28349__704 (.L_HI(net704));
 sg13g2_tiehi _28348__705 (.L_HI(net705));
 sg13g2_tiehi _28347__706 (.L_HI(net706));
 sg13g2_tiehi _28346__707 (.L_HI(net707));
 sg13g2_tiehi _28345__708 (.L_HI(net708));
 sg13g2_tiehi _28344__709 (.L_HI(net709));
 sg13g2_tiehi _28343__710 (.L_HI(net710));
 sg13g2_tiehi _28342__711 (.L_HI(net711));
 sg13g2_tiehi _28341__712 (.L_HI(net712));
 sg13g2_tiehi _28340__713 (.L_HI(net713));
 sg13g2_tiehi _28339__714 (.L_HI(net714));
 sg13g2_tiehi _28338__715 (.L_HI(net715));
 sg13g2_tiehi _28337__716 (.L_HI(net716));
 sg13g2_tiehi _28336__717 (.L_HI(net717));
 sg13g2_tiehi _28335__718 (.L_HI(net718));
 sg13g2_tiehi _28334__719 (.L_HI(net719));
 sg13g2_tiehi _28333__720 (.L_HI(net720));
 sg13g2_tiehi _28332__721 (.L_HI(net721));
 sg13g2_tiehi _28331__722 (.L_HI(net722));
 sg13g2_tiehi _28330__723 (.L_HI(net723));
 sg13g2_tiehi _28329__724 (.L_HI(net724));
 sg13g2_tiehi _28328__725 (.L_HI(net725));
 sg13g2_tiehi _28327__726 (.L_HI(net726));
 sg13g2_tiehi _28326__727 (.L_HI(net727));
 sg13g2_tiehi _28325__728 (.L_HI(net728));
 sg13g2_tiehi _28324__729 (.L_HI(net729));
 sg13g2_tiehi _28323__730 (.L_HI(net730));
 sg13g2_tiehi _28322__731 (.L_HI(net731));
 sg13g2_tiehi _28321__732 (.L_HI(net732));
 sg13g2_tiehi _28320__733 (.L_HI(net733));
 sg13g2_tiehi _28319__734 (.L_HI(net734));
 sg13g2_tiehi _28318__735 (.L_HI(net735));
 sg13g2_tiehi _28317__736 (.L_HI(net736));
 sg13g2_tiehi _28316__737 (.L_HI(net737));
 sg13g2_tiehi _28315__738 (.L_HI(net738));
 sg13g2_tiehi _28314__739 (.L_HI(net739));
 sg13g2_tiehi _28313__740 (.L_HI(net740));
 sg13g2_tiehi _28312__741 (.L_HI(net741));
 sg13g2_tiehi _29171__742 (.L_HI(net742));
 sg13g2_tiehi _28311__743 (.L_HI(net743));
 sg13g2_tiehi _29170__744 (.L_HI(net744));
 sg13g2_tiehi _28310__745 (.L_HI(net745));
 sg13g2_tiehi _29169__746 (.L_HI(net746));
 sg13g2_tiehi _28309__747 (.L_HI(net747));
 sg13g2_tiehi _29168__748 (.L_HI(net748));
 sg13g2_tiehi _28308__749 (.L_HI(net749));
 sg13g2_tiehi _29167__750 (.L_HI(net750));
 sg13g2_tiehi _28307__751 (.L_HI(net751));
 sg13g2_tiehi _28306__752 (.L_HI(net752));
 sg13g2_tiehi _28305__753 (.L_HI(net753));
 sg13g2_tiehi _28304__754 (.L_HI(net754));
 sg13g2_tiehi _28303__755 (.L_HI(net755));
 sg13g2_tiehi _28302__756 (.L_HI(net756));
 sg13g2_tiehi _28301__757 (.L_HI(net757));
 sg13g2_tiehi _28300__758 (.L_HI(net758));
 sg13g2_tiehi _28299__759 (.L_HI(net759));
 sg13g2_tiehi _28298__760 (.L_HI(net760));
 sg13g2_tiehi _28297__761 (.L_HI(net761));
 sg13g2_tiehi _28296__762 (.L_HI(net762));
 sg13g2_tiehi _28295__763 (.L_HI(net763));
 sg13g2_tiehi _28294__764 (.L_HI(net764));
 sg13g2_tiehi _28293__765 (.L_HI(net765));
 sg13g2_tiehi _28292__766 (.L_HI(net766));
 sg13g2_tiehi _28291__767 (.L_HI(net767));
 sg13g2_tiehi _28290__768 (.L_HI(net768));
 sg13g2_tiehi _28289__769 (.L_HI(net769));
 sg13g2_tiehi _28288__770 (.L_HI(net770));
 sg13g2_tiehi _28287__771 (.L_HI(net771));
 sg13g2_tiehi _28286__772 (.L_HI(net772));
 sg13g2_tiehi _28285__773 (.L_HI(net773));
 sg13g2_tiehi _28284__774 (.L_HI(net774));
 sg13g2_tiehi _28283__775 (.L_HI(net775));
 sg13g2_tiehi _28282__776 (.L_HI(net776));
 sg13g2_tiehi _28281__777 (.L_HI(net777));
 sg13g2_tiehi _28280__778 (.L_HI(net778));
 sg13g2_tiehi _28279__779 (.L_HI(net779));
 sg13g2_tiehi _28278__780 (.L_HI(net780));
 sg13g2_tiehi _28277__781 (.L_HI(net781));
 sg13g2_tiehi _28276__782 (.L_HI(net782));
 sg13g2_tiehi _28275__783 (.L_HI(net783));
 sg13g2_tiehi _28274__784 (.L_HI(net784));
 sg13g2_tiehi _28273__785 (.L_HI(net785));
 sg13g2_tiehi _28272__786 (.L_HI(net786));
 sg13g2_tiehi _28271__787 (.L_HI(net787));
 sg13g2_tiehi _28270__788 (.L_HI(net788));
 sg13g2_tiehi _28269__789 (.L_HI(net789));
 sg13g2_tiehi _28268__790 (.L_HI(net790));
 sg13g2_tiehi _28267__791 (.L_HI(net791));
 sg13g2_tiehi _28266__792 (.L_HI(net792));
 sg13g2_tiehi _28265__793 (.L_HI(net793));
 sg13g2_tiehi _28264__794 (.L_HI(net794));
 sg13g2_tiehi _28263__795 (.L_HI(net795));
 sg13g2_tiehi _28262__796 (.L_HI(net796));
 sg13g2_tiehi _28261__797 (.L_HI(net797));
 sg13g2_tiehi _28260__798 (.L_HI(net798));
 sg13g2_tiehi _28259__799 (.L_HI(net799));
 sg13g2_tiehi _28258__800 (.L_HI(net800));
 sg13g2_tiehi _28257__801 (.L_HI(net801));
 sg13g2_tiehi _28256__802 (.L_HI(net802));
 sg13g2_tiehi _28255__803 (.L_HI(net803));
 sg13g2_tiehi _28254__804 (.L_HI(net804));
 sg13g2_tiehi _28253__805 (.L_HI(net805));
 sg13g2_tiehi _28252__806 (.L_HI(net806));
 sg13g2_tiehi _28251__807 (.L_HI(net807));
 sg13g2_tiehi _28250__808 (.L_HI(net808));
 sg13g2_tiehi _29166__809 (.L_HI(net809));
 sg13g2_tiehi _28249__810 (.L_HI(net810));
 sg13g2_tiehi _29165__811 (.L_HI(net811));
 sg13g2_tiehi _28248__812 (.L_HI(net812));
 sg13g2_tiehi _29164__813 (.L_HI(net813));
 sg13g2_tiehi _28247__814 (.L_HI(net814));
 sg13g2_tiehi _29163__815 (.L_HI(net815));
 sg13g2_tiehi _28246__816 (.L_HI(net816));
 sg13g2_tiehi _29162__817 (.L_HI(net817));
 sg13g2_tiehi _28245__818 (.L_HI(net818));
 sg13g2_tiehi _29161__819 (.L_HI(net819));
 sg13g2_tiehi _28244__820 (.L_HI(net820));
 sg13g2_tiehi _29160__821 (.L_HI(net821));
 sg13g2_tiehi _28243__822 (.L_HI(net822));
 sg13g2_tiehi _29159__823 (.L_HI(net823));
 sg13g2_tiehi _28242__824 (.L_HI(net824));
 sg13g2_tiehi _29158__825 (.L_HI(net825));
 sg13g2_tiehi _28241__826 (.L_HI(net826));
 sg13g2_tiehi _29157__827 (.L_HI(net827));
 sg13g2_tiehi _28240__828 (.L_HI(net828));
 sg13g2_tiehi _29156__829 (.L_HI(net829));
 sg13g2_tiehi _28239__830 (.L_HI(net830));
 sg13g2_tiehi _29155__831 (.L_HI(net831));
 sg13g2_tiehi _28238__832 (.L_HI(net832));
 sg13g2_tiehi _29154__833 (.L_HI(net833));
 sg13g2_tiehi _28237__834 (.L_HI(net834));
 sg13g2_tiehi _29153__835 (.L_HI(net835));
 sg13g2_tiehi _28236__836 (.L_HI(net836));
 sg13g2_tiehi _29152__837 (.L_HI(net837));
 sg13g2_tiehi _28235__838 (.L_HI(net838));
 sg13g2_tiehi _29151__839 (.L_HI(net839));
 sg13g2_tiehi _28234__840 (.L_HI(net840));
 sg13g2_tiehi _29150__841 (.L_HI(net841));
 sg13g2_tiehi _28233__842 (.L_HI(net842));
 sg13g2_tiehi _29149__843 (.L_HI(net843));
 sg13g2_tiehi _28232__844 (.L_HI(net844));
 sg13g2_tiehi _29148__845 (.L_HI(net845));
 sg13g2_tiehi _28231__846 (.L_HI(net846));
 sg13g2_tiehi _29147__847 (.L_HI(net847));
 sg13g2_tiehi _28230__848 (.L_HI(net848));
 sg13g2_tiehi _29146__849 (.L_HI(net849));
 sg13g2_tiehi _28229__850 (.L_HI(net850));
 sg13g2_tiehi _29145__851 (.L_HI(net851));
 sg13g2_tiehi _28228__852 (.L_HI(net852));
 sg13g2_tiehi _29144__853 (.L_HI(net853));
 sg13g2_tiehi _28227__854 (.L_HI(net854));
 sg13g2_tiehi _29143__855 (.L_HI(net855));
 sg13g2_tiehi _28226__856 (.L_HI(net856));
 sg13g2_tiehi _29142__857 (.L_HI(net857));
 sg13g2_tiehi _28225__858 (.L_HI(net858));
 sg13g2_tiehi _29141__859 (.L_HI(net859));
 sg13g2_tiehi _28224__860 (.L_HI(net860));
 sg13g2_tiehi _29140__861 (.L_HI(net861));
 sg13g2_tiehi _28223__862 (.L_HI(net862));
 sg13g2_tiehi _29139__863 (.L_HI(net863));
 sg13g2_tiehi _28222__864 (.L_HI(net864));
 sg13g2_tiehi _28221__865 (.L_HI(net865));
 sg13g2_tiehi _28220__866 (.L_HI(net866));
 sg13g2_tiehi _28219__867 (.L_HI(net867));
 sg13g2_tiehi _28218__868 (.L_HI(net868));
 sg13g2_tiehi _28217__869 (.L_HI(net869));
 sg13g2_tiehi _28216__870 (.L_HI(net870));
 sg13g2_tiehi _28215__871 (.L_HI(net871));
 sg13g2_tiehi _28214__872 (.L_HI(net872));
 sg13g2_tiehi _28213__873 (.L_HI(net873));
 sg13g2_tiehi _28212__874 (.L_HI(net874));
 sg13g2_tiehi _28211__875 (.L_HI(net875));
 sg13g2_tiehi _28210__876 (.L_HI(net876));
 sg13g2_tiehi _28209__877 (.L_HI(net877));
 sg13g2_tiehi _28208__878 (.L_HI(net878));
 sg13g2_tiehi _28207__879 (.L_HI(net879));
 sg13g2_tiehi _28206__880 (.L_HI(net880));
 sg13g2_tiehi _28205__881 (.L_HI(net881));
 sg13g2_tiehi _28204__882 (.L_HI(net882));
 sg13g2_tiehi _28203__883 (.L_HI(net883));
 sg13g2_tiehi _28202__884 (.L_HI(net884));
 sg13g2_tiehi _28201__885 (.L_HI(net885));
 sg13g2_tiehi _28200__886 (.L_HI(net886));
 sg13g2_tiehi _28199__887 (.L_HI(net887));
 sg13g2_tiehi _28198__888 (.L_HI(net888));
 sg13g2_tiehi _28197__889 (.L_HI(net889));
 sg13g2_tiehi _28196__890 (.L_HI(net890));
 sg13g2_tiehi _28195__891 (.L_HI(net891));
 sg13g2_tiehi _28194__892 (.L_HI(net892));
 sg13g2_tiehi _28193__893 (.L_HI(net893));
 sg13g2_tiehi _28192__894 (.L_HI(net894));
 sg13g2_tiehi _28191__895 (.L_HI(net895));
 sg13g2_tiehi _28190__896 (.L_HI(net896));
 sg13g2_tiehi _28189__897 (.L_HI(net897));
 sg13g2_tiehi _28188__898 (.L_HI(net898));
 sg13g2_tiehi _28187__899 (.L_HI(net899));
 sg13g2_tiehi _28186__900 (.L_HI(net900));
 sg13g2_tiehi _28185__901 (.L_HI(net901));
 sg13g2_tiehi _28184__902 (.L_HI(net902));
 sg13g2_tiehi _28183__903 (.L_HI(net903));
 sg13g2_tiehi _29138__904 (.L_HI(net904));
 sg13g2_tiehi _28182__905 (.L_HI(net905));
 sg13g2_tiehi _29137__906 (.L_HI(net906));
 sg13g2_tiehi _28181__907 (.L_HI(net907));
 sg13g2_tiehi _29136__908 (.L_HI(net908));
 sg13g2_tiehi _28180__909 (.L_HI(net909));
 sg13g2_tiehi _29135__910 (.L_HI(net910));
 sg13g2_tiehi _28179__911 (.L_HI(net911));
 sg13g2_tiehi _29134__912 (.L_HI(net912));
 sg13g2_tiehi _28178__913 (.L_HI(net913));
 sg13g2_tiehi _29133__914 (.L_HI(net914));
 sg13g2_tiehi _28177__915 (.L_HI(net915));
 sg13g2_tiehi _29132__916 (.L_HI(net916));
 sg13g2_tiehi _28176__917 (.L_HI(net917));
 sg13g2_tiehi _29131__918 (.L_HI(net918));
 sg13g2_tiehi _28175__919 (.L_HI(net919));
 sg13g2_tiehi _29130__920 (.L_HI(net920));
 sg13g2_tiehi _28174__921 (.L_HI(net921));
 sg13g2_tiehi _29129__922 (.L_HI(net922));
 sg13g2_tiehi _28173__923 (.L_HI(net923));
 sg13g2_tiehi _29128__924 (.L_HI(net924));
 sg13g2_tiehi _28172__925 (.L_HI(net925));
 sg13g2_tiehi _29127__926 (.L_HI(net926));
 sg13g2_tiehi _28171__927 (.L_HI(net927));
 sg13g2_tiehi _29126__928 (.L_HI(net928));
 sg13g2_tiehi _28170__929 (.L_HI(net929));
 sg13g2_tiehi _29125__930 (.L_HI(net930));
 sg13g2_tiehi _28169__931 (.L_HI(net931));
 sg13g2_tiehi _29124__932 (.L_HI(net932));
 sg13g2_tiehi _28168__933 (.L_HI(net933));
 sg13g2_tiehi _29123__934 (.L_HI(net934));
 sg13g2_tiehi _28167__935 (.L_HI(net935));
 sg13g2_tiehi _29122__936 (.L_HI(net936));
 sg13g2_tiehi _28166__937 (.L_HI(net937));
 sg13g2_tiehi _29121__938 (.L_HI(net938));
 sg13g2_tiehi _28165__939 (.L_HI(net939));
 sg13g2_tiehi _29120__940 (.L_HI(net940));
 sg13g2_tiehi _28164__941 (.L_HI(net941));
 sg13g2_tiehi _29119__942 (.L_HI(net942));
 sg13g2_tiehi _28163__943 (.L_HI(net943));
 sg13g2_tiehi _29118__944 (.L_HI(net944));
 sg13g2_tiehi _28162__945 (.L_HI(net945));
 sg13g2_tiehi _29117__946 (.L_HI(net946));
 sg13g2_tiehi _28161__947 (.L_HI(net947));
 sg13g2_tiehi _29116__948 (.L_HI(net948));
 sg13g2_tiehi _28160__949 (.L_HI(net949));
 sg13g2_tiehi _29115__950 (.L_HI(net950));
 sg13g2_tiehi _28159__951 (.L_HI(net951));
 sg13g2_tiehi _28158__952 (.L_HI(net952));
 sg13g2_tiehi _28157__953 (.L_HI(net953));
 sg13g2_tiehi _28156__954 (.L_HI(net954));
 sg13g2_tiehi _28155__955 (.L_HI(net955));
 sg13g2_tiehi _28154__956 (.L_HI(net956));
 sg13g2_tiehi _28153__957 (.L_HI(net957));
 sg13g2_tiehi _28152__958 (.L_HI(net958));
 sg13g2_tiehi _28151__959 (.L_HI(net959));
 sg13g2_tiehi _29114__960 (.L_HI(net960));
 sg13g2_tiehi _28150__961 (.L_HI(net961));
 sg13g2_tiehi _29113__962 (.L_HI(net962));
 sg13g2_tiehi _28149__963 (.L_HI(net963));
 sg13g2_tiehi _29112__964 (.L_HI(net964));
 sg13g2_tiehi _28148__965 (.L_HI(net965));
 sg13g2_tiehi _29111__966 (.L_HI(net966));
 sg13g2_tiehi _28147__967 (.L_HI(net967));
 sg13g2_tiehi _29110__968 (.L_HI(net968));
 sg13g2_tiehi _28146__969 (.L_HI(net969));
 sg13g2_tiehi _29109__970 (.L_HI(net970));
 sg13g2_tiehi _28145__971 (.L_HI(net971));
 sg13g2_tiehi _29108__972 (.L_HI(net972));
 sg13g2_tiehi _28144__973 (.L_HI(net973));
 sg13g2_tiehi _29107__974 (.L_HI(net974));
 sg13g2_tiehi _28143__975 (.L_HI(net975));
 sg13g2_tiehi _29106__976 (.L_HI(net976));
 sg13g2_tiehi _28142__977 (.L_HI(net977));
 sg13g2_tiehi _28141__978 (.L_HI(net978));
 sg13g2_tiehi _28140__979 (.L_HI(net979));
 sg13g2_tiehi _28139__980 (.L_HI(net980));
 sg13g2_tiehi _28138__981 (.L_HI(net981));
 sg13g2_tiehi _28137__982 (.L_HI(net982));
 sg13g2_tiehi _28136__983 (.L_HI(net983));
 sg13g2_tiehi _28135__984 (.L_HI(net984));
 sg13g2_tiehi _28134__985 (.L_HI(net985));
 sg13g2_tiehi _28133__986 (.L_HI(net986));
 sg13g2_tiehi _28132__987 (.L_HI(net987));
 sg13g2_tiehi _28131__988 (.L_HI(net988));
 sg13g2_tiehi _28130__989 (.L_HI(net989));
 sg13g2_tiehi _28129__990 (.L_HI(net990));
 sg13g2_tiehi _28128__991 (.L_HI(net991));
 sg13g2_tiehi _28127__992 (.L_HI(net992));
 sg13g2_tiehi _28126__993 (.L_HI(net993));
 sg13g2_tiehi _28125__994 (.L_HI(net994));
 sg13g2_tiehi _28124__995 (.L_HI(net995));
 sg13g2_tiehi _28123__996 (.L_HI(net996));
 sg13g2_tiehi _28122__997 (.L_HI(net997));
 sg13g2_tiehi _28121__998 (.L_HI(net998));
 sg13g2_tiehi _28120__999 (.L_HI(net999));
 sg13g2_tiehi _28119__1000 (.L_HI(net1000));
 sg13g2_tiehi _28118__1001 (.L_HI(net1001));
 sg13g2_tiehi _28117__1002 (.L_HI(net1002));
 sg13g2_tiehi _28116__1003 (.L_HI(net1003));
 sg13g2_tiehi _28115__1004 (.L_HI(net1004));
 sg13g2_tiehi _28114__1005 (.L_HI(net1005));
 sg13g2_tiehi _28113__1006 (.L_HI(net1006));
 sg13g2_tiehi _28112__1007 (.L_HI(net1007));
 sg13g2_tiehi _28111__1008 (.L_HI(net1008));
 sg13g2_tiehi _28110__1009 (.L_HI(net1009));
 sg13g2_tiehi _28109__1010 (.L_HI(net1010));
 sg13g2_tiehi _28108__1011 (.L_HI(net1011));
 sg13g2_tiehi _28107__1012 (.L_HI(net1012));
 sg13g2_tiehi _28106__1013 (.L_HI(net1013));
 sg13g2_tiehi _28105__1014 (.L_HI(net1014));
 sg13g2_tiehi _28104__1015 (.L_HI(net1015));
 sg13g2_tiehi _28103__1016 (.L_HI(net1016));
 sg13g2_tiehi _28102__1017 (.L_HI(net1017));
 sg13g2_tiehi _28101__1018 (.L_HI(net1018));
 sg13g2_tiehi _28100__1019 (.L_HI(net1019));
 sg13g2_tiehi _28099__1020 (.L_HI(net1020));
 sg13g2_tiehi _28098__1021 (.L_HI(net1021));
 sg13g2_tiehi _28097__1022 (.L_HI(net1022));
 sg13g2_tiehi _28096__1023 (.L_HI(net1023));
 sg13g2_tiehi _28095__1024 (.L_HI(net1024));
 sg13g2_tiehi _28094__1025 (.L_HI(net1025));
 sg13g2_tiehi _28093__1026 (.L_HI(net1026));
 sg13g2_tiehi _28092__1027 (.L_HI(net1027));
 sg13g2_tiehi _28091__1028 (.L_HI(net1028));
 sg13g2_tiehi _28090__1029 (.L_HI(net1029));
 sg13g2_tiehi _28089__1030 (.L_HI(net1030));
 sg13g2_tiehi _28088__1031 (.L_HI(net1031));
 sg13g2_tiehi _28087__1032 (.L_HI(net1032));
 sg13g2_tiehi _28086__1033 (.L_HI(net1033));
 sg13g2_tiehi _28085__1034 (.L_HI(net1034));
 sg13g2_tiehi _28084__1035 (.L_HI(net1035));
 sg13g2_tiehi _28083__1036 (.L_HI(net1036));
 sg13g2_tiehi _28082__1037 (.L_HI(net1037));
 sg13g2_tiehi _28081__1038 (.L_HI(net1038));
 sg13g2_tiehi _28080__1039 (.L_HI(net1039));
 sg13g2_tiehi _28079__1040 (.L_HI(net1040));
 sg13g2_tiehi _28078__1041 (.L_HI(net1041));
 sg13g2_tiehi _28077__1042 (.L_HI(net1042));
 sg13g2_tiehi _28076__1043 (.L_HI(net1043));
 sg13g2_tiehi _28075__1044 (.L_HI(net1044));
 sg13g2_tiehi _28074__1045 (.L_HI(net1045));
 sg13g2_tiehi _28073__1046 (.L_HI(net1046));
 sg13g2_tiehi _28072__1047 (.L_HI(net1047));
 sg13g2_tiehi _28071__1048 (.L_HI(net1048));
 sg13g2_tiehi _28070__1049 (.L_HI(net1049));
 sg13g2_tiehi _28069__1050 (.L_HI(net1050));
 sg13g2_tiehi _28068__1051 (.L_HI(net1051));
 sg13g2_tiehi _28067__1052 (.L_HI(net1052));
 sg13g2_tiehi _28066__1053 (.L_HI(net1053));
 sg13g2_tiehi _28065__1054 (.L_HI(net1054));
 sg13g2_tiehi _28064__1055 (.L_HI(net1055));
 sg13g2_tiehi _28063__1056 (.L_HI(net1056));
 sg13g2_tiehi _28062__1057 (.L_HI(net1057));
 sg13g2_tiehi _28061__1058 (.L_HI(net1058));
 sg13g2_tiehi _28060__1059 (.L_HI(net1059));
 sg13g2_tiehi _28059__1060 (.L_HI(net1060));
 sg13g2_tiehi _28058__1061 (.L_HI(net1061));
 sg13g2_tiehi _28057__1062 (.L_HI(net1062));
 sg13g2_tiehi _28056__1063 (.L_HI(net1063));
 sg13g2_tiehi _28055__1064 (.L_HI(net1064));
 sg13g2_tiehi _28054__1065 (.L_HI(net1065));
 sg13g2_tiehi _28053__1066 (.L_HI(net1066));
 sg13g2_tiehi _28052__1067 (.L_HI(net1067));
 sg13g2_tiehi _28051__1068 (.L_HI(net1068));
 sg13g2_tiehi _28050__1069 (.L_HI(net1069));
 sg13g2_tiehi _28049__1070 (.L_HI(net1070));
 sg13g2_tiehi _28048__1071 (.L_HI(net1071));
 sg13g2_tiehi _28047__1072 (.L_HI(net1072));
 sg13g2_tiehi _28046__1073 (.L_HI(net1073));
 sg13g2_tiehi _28045__1074 (.L_HI(net1074));
 sg13g2_tiehi _28044__1075 (.L_HI(net1075));
 sg13g2_tiehi _28043__1076 (.L_HI(net1076));
 sg13g2_tiehi _28042__1077 (.L_HI(net1077));
 sg13g2_tiehi _28041__1078 (.L_HI(net1078));
 sg13g2_tiehi _28040__1079 (.L_HI(net1079));
 sg13g2_tiehi _28039__1080 (.L_HI(net1080));
 sg13g2_tiehi _28038__1081 (.L_HI(net1081));
 sg13g2_tiehi _28037__1082 (.L_HI(net1082));
 sg13g2_tiehi _28036__1083 (.L_HI(net1083));
 sg13g2_tiehi _28035__1084 (.L_HI(net1084));
 sg13g2_tiehi _28034__1085 (.L_HI(net1085));
 sg13g2_tiehi _28033__1086 (.L_HI(net1086));
 sg13g2_tiehi _28032__1087 (.L_HI(net1087));
 sg13g2_tiehi _28031__1088 (.L_HI(net1088));
 sg13g2_tiehi _28030__1089 (.L_HI(net1089));
 sg13g2_tiehi _28029__1090 (.L_HI(net1090));
 sg13g2_tiehi _28028__1091 (.L_HI(net1091));
 sg13g2_tiehi _28027__1092 (.L_HI(net1092));
 sg13g2_tiehi _28026__1093 (.L_HI(net1093));
 sg13g2_tiehi _28025__1094 (.L_HI(net1094));
 sg13g2_tiehi _28024__1095 (.L_HI(net1095));
 sg13g2_tiehi _28023__1096 (.L_HI(net1096));
 sg13g2_tiehi _28022__1097 (.L_HI(net1097));
 sg13g2_tiehi _28021__1098 (.L_HI(net1098));
 sg13g2_tiehi _28020__1099 (.L_HI(net1099));
 sg13g2_tiehi _28019__1100 (.L_HI(net1100));
 sg13g2_tiehi _28018__1101 (.L_HI(net1101));
 sg13g2_tiehi _28017__1102 (.L_HI(net1102));
 sg13g2_tiehi _28016__1103 (.L_HI(net1103));
 sg13g2_tiehi _28015__1104 (.L_HI(net1104));
 sg13g2_tiehi _28014__1105 (.L_HI(net1105));
 sg13g2_tiehi _28013__1106 (.L_HI(net1106));
 sg13g2_tiehi _28012__1107 (.L_HI(net1107));
 sg13g2_tiehi _28011__1108 (.L_HI(net1108));
 sg13g2_tiehi _28010__1109 (.L_HI(net1109));
 sg13g2_tiehi _28009__1110 (.L_HI(net1110));
 sg13g2_tiehi _28008__1111 (.L_HI(net1111));
 sg13g2_tiehi _28007__1112 (.L_HI(net1112));
 sg13g2_tiehi _28006__1113 (.L_HI(net1113));
 sg13g2_tiehi _28005__1114 (.L_HI(net1114));
 sg13g2_tiehi _28004__1115 (.L_HI(net1115));
 sg13g2_tiehi _28003__1116 (.L_HI(net1116));
 sg13g2_tiehi _28002__1117 (.L_HI(net1117));
 sg13g2_tiehi _28001__1118 (.L_HI(net1118));
 sg13g2_tiehi _28000__1119 (.L_HI(net1119));
 sg13g2_tiehi _27999__1120 (.L_HI(net1120));
 sg13g2_tiehi _27998__1121 (.L_HI(net1121));
 sg13g2_tiehi _27997__1122 (.L_HI(net1122));
 sg13g2_tiehi _27996__1123 (.L_HI(net1123));
 sg13g2_tiehi _27995__1124 (.L_HI(net1124));
 sg13g2_tiehi _27994__1125 (.L_HI(net1125));
 sg13g2_tiehi _27993__1126 (.L_HI(net1126));
 sg13g2_tiehi _27992__1127 (.L_HI(net1127));
 sg13g2_tiehi _27991__1128 (.L_HI(net1128));
 sg13g2_tiehi _27990__1129 (.L_HI(net1129));
 sg13g2_tiehi _27989__1130 (.L_HI(net1130));
 sg13g2_tiehi _27988__1131 (.L_HI(net1131));
 sg13g2_tiehi _27987__1132 (.L_HI(net1132));
 sg13g2_tiehi _27986__1133 (.L_HI(net1133));
 sg13g2_tiehi _27985__1134 (.L_HI(net1134));
 sg13g2_tiehi _27984__1135 (.L_HI(net1135));
 sg13g2_tiehi _27983__1136 (.L_HI(net1136));
 sg13g2_tiehi _27982__1137 (.L_HI(net1137));
 sg13g2_tiehi _27981__1138 (.L_HI(net1138));
 sg13g2_tiehi _27980__1139 (.L_HI(net1139));
 sg13g2_tiehi _27979__1140 (.L_HI(net1140));
 sg13g2_tiehi _27978__1141 (.L_HI(net1141));
 sg13g2_tiehi _27977__1142 (.L_HI(net1142));
 sg13g2_tiehi _27976__1143 (.L_HI(net1143));
 sg13g2_tiehi _27975__1144 (.L_HI(net1144));
 sg13g2_tiehi _27974__1145 (.L_HI(net1145));
 sg13g2_tiehi _27973__1146 (.L_HI(net1146));
 sg13g2_tiehi _27972__1147 (.L_HI(net1147));
 sg13g2_tiehi _27971__1148 (.L_HI(net1148));
 sg13g2_tiehi _27970__1149 (.L_HI(net1149));
 sg13g2_tiehi _27969__1150 (.L_HI(net1150));
 sg13g2_tiehi _27968__1151 (.L_HI(net1151));
 sg13g2_tiehi _27967__1152 (.L_HI(net1152));
 sg13g2_tiehi _27966__1153 (.L_HI(net1153));
 sg13g2_tiehi _27965__1154 (.L_HI(net1154));
 sg13g2_tiehi _27964__1155 (.L_HI(net1155));
 sg13g2_tiehi _27963__1156 (.L_HI(net1156));
 sg13g2_tiehi _27962__1157 (.L_HI(net1157));
 sg13g2_tiehi _27961__1158 (.L_HI(net1158));
 sg13g2_tiehi _27960__1159 (.L_HI(net1159));
 sg13g2_tiehi _27959__1160 (.L_HI(net1160));
 sg13g2_tiehi _27958__1161 (.L_HI(net1161));
 sg13g2_tiehi _27957__1162 (.L_HI(net1162));
 sg13g2_tiehi _27956__1163 (.L_HI(net1163));
 sg13g2_tiehi _27955__1164 (.L_HI(net1164));
 sg13g2_tiehi _27954__1165 (.L_HI(net1165));
 sg13g2_tiehi _27953__1166 (.L_HI(net1166));
 sg13g2_tiehi _27952__1167 (.L_HI(net1167));
 sg13g2_tiehi _27951__1168 (.L_HI(net1168));
 sg13g2_tiehi _27950__1169 (.L_HI(net1169));
 sg13g2_tiehi _27949__1170 (.L_HI(net1170));
 sg13g2_tiehi _27948__1171 (.L_HI(net1171));
 sg13g2_tiehi _27947__1172 (.L_HI(net1172));
 sg13g2_tiehi _27946__1173 (.L_HI(net1173));
 sg13g2_tiehi _27945__1174 (.L_HI(net1174));
 sg13g2_tiehi _27944__1175 (.L_HI(net1175));
 sg13g2_tiehi _27943__1176 (.L_HI(net1176));
 sg13g2_tiehi _27942__1177 (.L_HI(net1177));
 sg13g2_tiehi _27941__1178 (.L_HI(net1178));
 sg13g2_tiehi _27940__1179 (.L_HI(net1179));
 sg13g2_tiehi _27939__1180 (.L_HI(net1180));
 sg13g2_tiehi _27938__1181 (.L_HI(net1181));
 sg13g2_tiehi _27937__1182 (.L_HI(net1182));
 sg13g2_tiehi _27936__1183 (.L_HI(net1183));
 sg13g2_tiehi _27935__1184 (.L_HI(net1184));
 sg13g2_tiehi _27934__1185 (.L_HI(net1185));
 sg13g2_tiehi _27933__1186 (.L_HI(net1186));
 sg13g2_tiehi _27932__1187 (.L_HI(net1187));
 sg13g2_tiehi _27931__1188 (.L_HI(net1188));
 sg13g2_tiehi _27930__1189 (.L_HI(net1189));
 sg13g2_tiehi _27929__1190 (.L_HI(net1190));
 sg13g2_tiehi _27928__1191 (.L_HI(net1191));
 sg13g2_tiehi _27927__1192 (.L_HI(net1192));
 sg13g2_tiehi _27926__1193 (.L_HI(net1193));
 sg13g2_tiehi _27925__1194 (.L_HI(net1194));
 sg13g2_tiehi _27924__1195 (.L_HI(net1195));
 sg13g2_tiehi _27923__1196 (.L_HI(net1196));
 sg13g2_tiehi _27922__1197 (.L_HI(net1197));
 sg13g2_tiehi _27921__1198 (.L_HI(net1198));
 sg13g2_tiehi _27920__1199 (.L_HI(net1199));
 sg13g2_tiehi _27919__1200 (.L_HI(net1200));
 sg13g2_tiehi _27918__1201 (.L_HI(net1201));
 sg13g2_tiehi _27917__1202 (.L_HI(net1202));
 sg13g2_tiehi _27916__1203 (.L_HI(net1203));
 sg13g2_tiehi _27915__1204 (.L_HI(net1204));
 sg13g2_tiehi _27914__1205 (.L_HI(net1205));
 sg13g2_tiehi _27913__1206 (.L_HI(net1206));
 sg13g2_tiehi _27912__1207 (.L_HI(net1207));
 sg13g2_tiehi _27911__1208 (.L_HI(net1208));
 sg13g2_tiehi _27910__1209 (.L_HI(net1209));
 sg13g2_tiehi _27909__1210 (.L_HI(net1210));
 sg13g2_tiehi _27908__1211 (.L_HI(net1211));
 sg13g2_tiehi _27907__1212 (.L_HI(net1212));
 sg13g2_tiehi _27906__1213 (.L_HI(net1213));
 sg13g2_tiehi _27905__1214 (.L_HI(net1214));
 sg13g2_tiehi _27904__1215 (.L_HI(net1215));
 sg13g2_tiehi _27903__1216 (.L_HI(net1216));
 sg13g2_tiehi _27902__1217 (.L_HI(net1217));
 sg13g2_tiehi _27901__1218 (.L_HI(net1218));
 sg13g2_tiehi _27900__1219 (.L_HI(net1219));
 sg13g2_tiehi _27899__1220 (.L_HI(net1220));
 sg13g2_tiehi _27898__1221 (.L_HI(net1221));
 sg13g2_tiehi _27897__1222 (.L_HI(net1222));
 sg13g2_tiehi _27896__1223 (.L_HI(net1223));
 sg13g2_tiehi _27895__1224 (.L_HI(net1224));
 sg13g2_tiehi _27894__1225 (.L_HI(net1225));
 sg13g2_tiehi _27893__1226 (.L_HI(net1226));
 sg13g2_tiehi _27892__1227 (.L_HI(net1227));
 sg13g2_tiehi _27891__1228 (.L_HI(net1228));
 sg13g2_tiehi _27890__1229 (.L_HI(net1229));
 sg13g2_tiehi _27889__1230 (.L_HI(net1230));
 sg13g2_tiehi _27888__1231 (.L_HI(net1231));
 sg13g2_tiehi _27887__1232 (.L_HI(net1232));
 sg13g2_tiehi _26549__1233 (.L_HI(net1233));
 sg13g2_tiehi _27097__1234 (.L_HI(net1234));
 sg13g2_tiehi _27098__1235 (.L_HI(net1235));
 sg13g2_tiehi _27099__1236 (.L_HI(net1236));
 sg13g2_tiehi _27100__1237 (.L_HI(net1237));
 sg13g2_tiehi _27101__1238 (.L_HI(net1238));
 sg13g2_tiehi _27102__1239 (.L_HI(net1239));
 sg13g2_tiehi _27103__1240 (.L_HI(net1240));
 sg13g2_tiehi _27886__1241 (.L_HI(net1241));
 sg13g2_tiehi _27885__1242 (.L_HI(net1242));
 sg13g2_tiehi _27884__1243 (.L_HI(net1243));
 sg13g2_tiehi _27883__1244 (.L_HI(net1244));
 sg13g2_tiehi _27882__1245 (.L_HI(net1245));
 sg13g2_tiehi _27881__1246 (.L_HI(net1246));
 sg13g2_tiehi _27880__1247 (.L_HI(net1247));
 sg13g2_tiehi _27879__1248 (.L_HI(net1248));
 sg13g2_tiehi _27878__1249 (.L_HI(net1249));
 sg13g2_tiehi _27877__1250 (.L_HI(net1250));
 sg13g2_tiehi _27876__1251 (.L_HI(net1251));
 sg13g2_tiehi _27875__1252 (.L_HI(net1252));
 sg13g2_tiehi _27874__1253 (.L_HI(net1253));
 sg13g2_tiehi _27873__1254 (.L_HI(net1254));
 sg13g2_tiehi _27872__1255 (.L_HI(net1255));
 sg13g2_tiehi _27871__1256 (.L_HI(net1256));
 sg13g2_tiehi _27870__1257 (.L_HI(net1257));
 sg13g2_tiehi _27869__1258 (.L_HI(net1258));
 sg13g2_tiehi _27868__1259 (.L_HI(net1259));
 sg13g2_tiehi _27867__1260 (.L_HI(net1260));
 sg13g2_tiehi _27866__1261 (.L_HI(net1261));
 sg13g2_tiehi _27865__1262 (.L_HI(net1262));
 sg13g2_tiehi _27864__1263 (.L_HI(net1263));
 sg13g2_tiehi _27863__1264 (.L_HI(net1264));
 sg13g2_tiehi _27862__1265 (.L_HI(net1265));
 sg13g2_tiehi _27861__1266 (.L_HI(net1266));
 sg13g2_tiehi _27860__1267 (.L_HI(net1267));
 sg13g2_tiehi _27859__1268 (.L_HI(net1268));
 sg13g2_tiehi _27858__1269 (.L_HI(net1269));
 sg13g2_tiehi _27857__1270 (.L_HI(net1270));
 sg13g2_tiehi _27856__1271 (.L_HI(net1271));
 sg13g2_tiehi _27855__1272 (.L_HI(net1272));
 sg13g2_tiehi _27854__1273 (.L_HI(net1273));
 sg13g2_tiehi _27853__1274 (.L_HI(net1274));
 sg13g2_tiehi _27852__1275 (.L_HI(net1275));
 sg13g2_tiehi _27851__1276 (.L_HI(net1276));
 sg13g2_tiehi _27850__1277 (.L_HI(net1277));
 sg13g2_tiehi _27849__1278 (.L_HI(net1278));
 sg13g2_tiehi _27848__1279 (.L_HI(net1279));
 sg13g2_tiehi _27847__1280 (.L_HI(net1280));
 sg13g2_tiehi _27846__1281 (.L_HI(net1281));
 sg13g2_tiehi _27845__1282 (.L_HI(net1282));
 sg13g2_tiehi _27844__1283 (.L_HI(net1283));
 sg13g2_tiehi _27843__1284 (.L_HI(net1284));
 sg13g2_tiehi _27842__1285 (.L_HI(net1285));
 sg13g2_tiehi _27841__1286 (.L_HI(net1286));
 sg13g2_tiehi _27840__1287 (.L_HI(net1287));
 sg13g2_tiehi _27839__1288 (.L_HI(net1288));
 sg13g2_tiehi _27838__1289 (.L_HI(net1289));
 sg13g2_tiehi _27837__1290 (.L_HI(net1290));
 sg13g2_tiehi _27836__1291 (.L_HI(net1291));
 sg13g2_tiehi _27835__1292 (.L_HI(net1292));
 sg13g2_tiehi _27834__1293 (.L_HI(net1293));
 sg13g2_tiehi _27833__1294 (.L_HI(net1294));
 sg13g2_tiehi _27832__1295 (.L_HI(net1295));
 sg13g2_tiehi _27831__1296 (.L_HI(net1296));
 sg13g2_tiehi _27830__1297 (.L_HI(net1297));
 sg13g2_tiehi _27829__1298 (.L_HI(net1298));
 sg13g2_tiehi _27828__1299 (.L_HI(net1299));
 sg13g2_tiehi _27827__1300 (.L_HI(net1300));
 sg13g2_tiehi _27826__1301 (.L_HI(net1301));
 sg13g2_tiehi _27825__1302 (.L_HI(net1302));
 sg13g2_tiehi _27824__1303 (.L_HI(net1303));
 sg13g2_tiehi _27823__1304 (.L_HI(net1304));
 sg13g2_tiehi _27822__1305 (.L_HI(net1305));
 sg13g2_tiehi _27821__1306 (.L_HI(net1306));
 sg13g2_tiehi _27820__1307 (.L_HI(net1307));
 sg13g2_tiehi _27819__1308 (.L_HI(net1308));
 sg13g2_tiehi _27818__1309 (.L_HI(net1309));
 sg13g2_tiehi _27817__1310 (.L_HI(net1310));
 sg13g2_tiehi _27816__1311 (.L_HI(net1311));
 sg13g2_tiehi _27815__1312 (.L_HI(net1312));
 sg13g2_tiehi _27814__1313 (.L_HI(net1313));
 sg13g2_tiehi _27813__1314 (.L_HI(net1314));
 sg13g2_tiehi _27812__1315 (.L_HI(net1315));
 sg13g2_tiehi _27811__1316 (.L_HI(net1316));
 sg13g2_tiehi _27810__1317 (.L_HI(net1317));
 sg13g2_tiehi _27809__1318 (.L_HI(net1318));
 sg13g2_tiehi _27808__1319 (.L_HI(net1319));
 sg13g2_tiehi _27807__1320 (.L_HI(net1320));
 sg13g2_tiehi _27806__1321 (.L_HI(net1321));
 sg13g2_tiehi _27805__1322 (.L_HI(net1322));
 sg13g2_tiehi _27804__1323 (.L_HI(net1323));
 sg13g2_tiehi _27803__1324 (.L_HI(net1324));
 sg13g2_tiehi _27802__1325 (.L_HI(net1325));
 sg13g2_tiehi _27801__1326 (.L_HI(net1326));
 sg13g2_tiehi _27800__1327 (.L_HI(net1327));
 sg13g2_tiehi _27799__1328 (.L_HI(net1328));
 sg13g2_tiehi _27798__1329 (.L_HI(net1329));
 sg13g2_tiehi _27797__1330 (.L_HI(net1330));
 sg13g2_tiehi _27796__1331 (.L_HI(net1331));
 sg13g2_tiehi _27795__1332 (.L_HI(net1332));
 sg13g2_tiehi _27794__1333 (.L_HI(net1333));
 sg13g2_tiehi _27793__1334 (.L_HI(net1334));
 sg13g2_tiehi _27792__1335 (.L_HI(net1335));
 sg13g2_tiehi _27791__1336 (.L_HI(net1336));
 sg13g2_tiehi _27790__1337 (.L_HI(net1337));
 sg13g2_tiehi _27789__1338 (.L_HI(net1338));
 sg13g2_tiehi _27788__1339 (.L_HI(net1339));
 sg13g2_tiehi _27787__1340 (.L_HI(net1340));
 sg13g2_tiehi _27786__1341 (.L_HI(net1341));
 sg13g2_tiehi _27785__1342 (.L_HI(net1342));
 sg13g2_tiehi _27784__1343 (.L_HI(net1343));
 sg13g2_tiehi _27783__1344 (.L_HI(net1344));
 sg13g2_tiehi _27782__1345 (.L_HI(net1345));
 sg13g2_tiehi _27781__1346 (.L_HI(net1346));
 sg13g2_tiehi _27780__1347 (.L_HI(net1347));
 sg13g2_tiehi _27779__1348 (.L_HI(net1348));
 sg13g2_tiehi _27778__1349 (.L_HI(net1349));
 sg13g2_tiehi _27777__1350 (.L_HI(net1350));
 sg13g2_tiehi _27776__1351 (.L_HI(net1351));
 sg13g2_tiehi _27775__1352 (.L_HI(net1352));
 sg13g2_tiehi _27774__1353 (.L_HI(net1353));
 sg13g2_tiehi _27773__1354 (.L_HI(net1354));
 sg13g2_tiehi _27772__1355 (.L_HI(net1355));
 sg13g2_tiehi _27771__1356 (.L_HI(net1356));
 sg13g2_tiehi _27770__1357 (.L_HI(net1357));
 sg13g2_tiehi _27769__1358 (.L_HI(net1358));
 sg13g2_tiehi _27768__1359 (.L_HI(net1359));
 sg13g2_tiehi _27767__1360 (.L_HI(net1360));
 sg13g2_tiehi _27766__1361 (.L_HI(net1361));
 sg13g2_tiehi _27765__1362 (.L_HI(net1362));
 sg13g2_tiehi _27764__1363 (.L_HI(net1363));
 sg13g2_tiehi _27763__1364 (.L_HI(net1364));
 sg13g2_tiehi _27762__1365 (.L_HI(net1365));
 sg13g2_tiehi _27761__1366 (.L_HI(net1366));
 sg13g2_tiehi _27760__1367 (.L_HI(net1367));
 sg13g2_tiehi _27759__1368 (.L_HI(net1368));
 sg13g2_tiehi _27758__1369 (.L_HI(net1369));
 sg13g2_tiehi _27757__1370 (.L_HI(net1370));
 sg13g2_tiehi _27756__1371 (.L_HI(net1371));
 sg13g2_tiehi _27755__1372 (.L_HI(net1372));
 sg13g2_tiehi _27754__1373 (.L_HI(net1373));
 sg13g2_tiehi _27753__1374 (.L_HI(net1374));
 sg13g2_tiehi _27752__1375 (.L_HI(net1375));
 sg13g2_tiehi _27751__1376 (.L_HI(net1376));
 sg13g2_tiehi _27750__1377 (.L_HI(net1377));
 sg13g2_tiehi _27749__1378 (.L_HI(net1378));
 sg13g2_tiehi _27748__1379 (.L_HI(net1379));
 sg13g2_tiehi _27747__1380 (.L_HI(net1380));
 sg13g2_tiehi _27746__1381 (.L_HI(net1381));
 sg13g2_tiehi _27745__1382 (.L_HI(net1382));
 sg13g2_tiehi _27744__1383 (.L_HI(net1383));
 sg13g2_tiehi _27743__1384 (.L_HI(net1384));
 sg13g2_tiehi _27742__1385 (.L_HI(net1385));
 sg13g2_tiehi _27741__1386 (.L_HI(net1386));
 sg13g2_tiehi _27740__1387 (.L_HI(net1387));
 sg13g2_tiehi _27739__1388 (.L_HI(net1388));
 sg13g2_tiehi _27738__1389 (.L_HI(net1389));
 sg13g2_tiehi _27737__1390 (.L_HI(net1390));
 sg13g2_tiehi _27736__1391 (.L_HI(net1391));
 sg13g2_tiehi _27735__1392 (.L_HI(net1392));
 sg13g2_tiehi _27734__1393 (.L_HI(net1393));
 sg13g2_tiehi _27733__1394 (.L_HI(net1394));
 sg13g2_tiehi _27732__1395 (.L_HI(net1395));
 sg13g2_tiehi _27731__1396 (.L_HI(net1396));
 sg13g2_tiehi _27730__1397 (.L_HI(net1397));
 sg13g2_tiehi _27729__1398 (.L_HI(net1398));
 sg13g2_tiehi _27728__1399 (.L_HI(net1399));
 sg13g2_tiehi _27727__1400 (.L_HI(net1400));
 sg13g2_tiehi _27726__1401 (.L_HI(net1401));
 sg13g2_tiehi _27725__1402 (.L_HI(net1402));
 sg13g2_tiehi _27724__1403 (.L_HI(net1403));
 sg13g2_tiehi _27723__1404 (.L_HI(net1404));
 sg13g2_tiehi _27722__1405 (.L_HI(net1405));
 sg13g2_tiehi _27721__1406 (.L_HI(net1406));
 sg13g2_tiehi _27720__1407 (.L_HI(net1407));
 sg13g2_tiehi _27719__1408 (.L_HI(net1408));
 sg13g2_tiehi _27718__1409 (.L_HI(net1409));
 sg13g2_tiehi _27717__1410 (.L_HI(net1410));
 sg13g2_tiehi _27716__1411 (.L_HI(net1411));
 sg13g2_tiehi _27715__1412 (.L_HI(net1412));
 sg13g2_tiehi _27714__1413 (.L_HI(net1413));
 sg13g2_tiehi _27713__1414 (.L_HI(net1414));
 sg13g2_tiehi _27712__1415 (.L_HI(net1415));
 sg13g2_tiehi _27711__1416 (.L_HI(net1416));
 sg13g2_tiehi _27710__1417 (.L_HI(net1417));
 sg13g2_tiehi _27709__1418 (.L_HI(net1418));
 sg13g2_tiehi _27708__1419 (.L_HI(net1419));
 sg13g2_tiehi _27707__1420 (.L_HI(net1420));
 sg13g2_tiehi _27706__1421 (.L_HI(net1421));
 sg13g2_tiehi _27705__1422 (.L_HI(net1422));
 sg13g2_tiehi _27704__1423 (.L_HI(net1423));
 sg13g2_tiehi _27703__1424 (.L_HI(net1424));
 sg13g2_tiehi _27702__1425 (.L_HI(net1425));
 sg13g2_tiehi _27701__1426 (.L_HI(net1426));
 sg13g2_tiehi _27700__1427 (.L_HI(net1427));
 sg13g2_tiehi _27699__1428 (.L_HI(net1428));
 sg13g2_tiehi _27698__1429 (.L_HI(net1429));
 sg13g2_tiehi _27697__1430 (.L_HI(net1430));
 sg13g2_tiehi _27696__1431 (.L_HI(net1431));
 sg13g2_tiehi _27695__1432 (.L_HI(net1432));
 sg13g2_tiehi _27694__1433 (.L_HI(net1433));
 sg13g2_tiehi _27693__1434 (.L_HI(net1434));
 sg13g2_tiehi _27692__1435 (.L_HI(net1435));
 sg13g2_tiehi _27691__1436 (.L_HI(net1436));
 sg13g2_tiehi _27690__1437 (.L_HI(net1437));
 sg13g2_tiehi _27689__1438 (.L_HI(net1438));
 sg13g2_tiehi _27688__1439 (.L_HI(net1439));
 sg13g2_tiehi _27687__1440 (.L_HI(net1440));
 sg13g2_tiehi _27686__1441 (.L_HI(net1441));
 sg13g2_tiehi _27685__1442 (.L_HI(net1442));
 sg13g2_tiehi _27684__1443 (.L_HI(net1443));
 sg13g2_tiehi _27683__1444 (.L_HI(net1444));
 sg13g2_tiehi _27682__1445 (.L_HI(net1445));
 sg13g2_tiehi _27681__1446 (.L_HI(net1446));
 sg13g2_tiehi _27680__1447 (.L_HI(net1447));
 sg13g2_tiehi _27679__1448 (.L_HI(net1448));
 sg13g2_tiehi _27678__1449 (.L_HI(net1449));
 sg13g2_tiehi _27677__1450 (.L_HI(net1450));
 sg13g2_tiehi _27676__1451 (.L_HI(net1451));
 sg13g2_tiehi _27675__1452 (.L_HI(net1452));
 sg13g2_tiehi _27674__1453 (.L_HI(net1453));
 sg13g2_tiehi _27673__1454 (.L_HI(net1454));
 sg13g2_tiehi _27672__1455 (.L_HI(net1455));
 sg13g2_tiehi _27671__1456 (.L_HI(net1456));
 sg13g2_tiehi _27670__1457 (.L_HI(net1457));
 sg13g2_tiehi _27669__1458 (.L_HI(net1458));
 sg13g2_tiehi _27668__1459 (.L_HI(net1459));
 sg13g2_tiehi _27667__1460 (.L_HI(net1460));
 sg13g2_tiehi _27666__1461 (.L_HI(net1461));
 sg13g2_tiehi _27665__1462 (.L_HI(net1462));
 sg13g2_tiehi _27664__1463 (.L_HI(net1463));
 sg13g2_tiehi _27663__1464 (.L_HI(net1464));
 sg13g2_tiehi _27662__1465 (.L_HI(net1465));
 sg13g2_tiehi _27661__1466 (.L_HI(net1466));
 sg13g2_tiehi _27660__1467 (.L_HI(net1467));
 sg13g2_tiehi _27659__1468 (.L_HI(net1468));
 sg13g2_tiehi _27658__1469 (.L_HI(net1469));
 sg13g2_tiehi _27657__1470 (.L_HI(net1470));
 sg13g2_tiehi _27656__1471 (.L_HI(net1471));
 sg13g2_tiehi _29105__1472 (.L_HI(net1472));
 sg13g2_tiehi _27648__1473 (.L_HI(net1473));
 sg13g2_tiehi _27647__1474 (.L_HI(net1474));
 sg13g2_tiehi _27646__1475 (.L_HI(net1475));
 sg13g2_tiehi _27645__1476 (.L_HI(net1476));
 sg13g2_tiehi _27644__1477 (.L_HI(net1477));
 sg13g2_tiehi _27643__1478 (.L_HI(net1478));
 sg13g2_tiehi _27642__1479 (.L_HI(net1479));
 sg13g2_tiehi _27641__1480 (.L_HI(net1480));
 sg13g2_tiehi _27640__1481 (.L_HI(net1481));
 sg13g2_tiehi _27639__1482 (.L_HI(net1482));
 sg13g2_tiehi _27638__1483 (.L_HI(net1483));
 sg13g2_tiehi _27637__1484 (.L_HI(net1484));
 sg13g2_tiehi _27636__1485 (.L_HI(net1485));
 sg13g2_tiehi _27635__1486 (.L_HI(net1486));
 sg13g2_tiehi _27634__1487 (.L_HI(net1487));
 sg13g2_tiehi _27633__1488 (.L_HI(net1488));
 sg13g2_tiehi _27632__1489 (.L_HI(net1489));
 sg13g2_tiehi _27631__1490 (.L_HI(net1490));
 sg13g2_tiehi _27630__1491 (.L_HI(net1491));
 sg13g2_tiehi _27629__1492 (.L_HI(net1492));
 sg13g2_tiehi _27628__1493 (.L_HI(net1493));
 sg13g2_tiehi _27627__1494 (.L_HI(net1494));
 sg13g2_tiehi _27626__1495 (.L_HI(net1495));
 sg13g2_tiehi _27625__1496 (.L_HI(net1496));
 sg13g2_tiehi _27624__1497 (.L_HI(net1497));
 sg13g2_tiehi _27623__1498 (.L_HI(net1498));
 sg13g2_tiehi _27622__1499 (.L_HI(net1499));
 sg13g2_tiehi _27621__1500 (.L_HI(net1500));
 sg13g2_tiehi _27620__1501 (.L_HI(net1501));
 sg13g2_tiehi _27619__1502 (.L_HI(net1502));
 sg13g2_tiehi _27618__1503 (.L_HI(net1503));
 sg13g2_tiehi _27617__1504 (.L_HI(net1504));
 sg13g2_tiehi _27616__1505 (.L_HI(net1505));
 sg13g2_tiehi _27615__1506 (.L_HI(net1506));
 sg13g2_tiehi _27614__1507 (.L_HI(net1507));
 sg13g2_tiehi _27613__1508 (.L_HI(net1508));
 sg13g2_tiehi _27612__1509 (.L_HI(net1509));
 sg13g2_tiehi _27611__1510 (.L_HI(net1510));
 sg13g2_tiehi _27610__1511 (.L_HI(net1511));
 sg13g2_tiehi _27609__1512 (.L_HI(net1512));
 sg13g2_tiehi _27608__1513 (.L_HI(net1513));
 sg13g2_tiehi _27607__1514 (.L_HI(net1514));
 sg13g2_tiehi _27606__1515 (.L_HI(net1515));
 sg13g2_tiehi _27605__1516 (.L_HI(net1516));
 sg13g2_tiehi _27604__1517 (.L_HI(net1517));
 sg13g2_tiehi _29104__1518 (.L_HI(net1518));
 sg13g2_tiehi _27603__1519 (.L_HI(net1519));
 sg13g2_tiehi _29103__1520 (.L_HI(net1520));
 sg13g2_tiehi _27602__1521 (.L_HI(net1521));
 sg13g2_tiehi _29102__1522 (.L_HI(net1522));
 sg13g2_tiehi _27601__1523 (.L_HI(net1523));
 sg13g2_tiehi _29101__1524 (.L_HI(net1524));
 sg13g2_tiehi _27600__1525 (.L_HI(net1525));
 sg13g2_tiehi _29100__1526 (.L_HI(net1526));
 sg13g2_tiehi _27599__1527 (.L_HI(net1527));
 sg13g2_tiehi _29099__1528 (.L_HI(net1528));
 sg13g2_tiehi _27598__1529 (.L_HI(net1529));
 sg13g2_tiehi _29098__1530 (.L_HI(net1530));
 sg13g2_tiehi _27597__1531 (.L_HI(net1531));
 sg13g2_tiehi _29097__1532 (.L_HI(net1532));
 sg13g2_tiehi _27596__1533 (.L_HI(net1533));
 sg13g2_tiehi _29096__1534 (.L_HI(net1534));
 sg13g2_tiehi _27595__1535 (.L_HI(net1535));
 sg13g2_tiehi _29095__1536 (.L_HI(net1536));
 sg13g2_tiehi _27594__1537 (.L_HI(net1537));
 sg13g2_tiehi _29094__1538 (.L_HI(net1538));
 sg13g2_tiehi _27593__1539 (.L_HI(net1539));
 sg13g2_tiehi _29093__1540 (.L_HI(net1540));
 sg13g2_tiehi _27592__1541 (.L_HI(net1541));
 sg13g2_tiehi _27591__1542 (.L_HI(net1542));
 sg13g2_tiehi _27590__1543 (.L_HI(net1543));
 sg13g2_tiehi _27589__1544 (.L_HI(net1544));
 sg13g2_tiehi _27588__1545 (.L_HI(net1545));
 sg13g2_tiehi _27587__1546 (.L_HI(net1546));
 sg13g2_tiehi _27586__1547 (.L_HI(net1547));
 sg13g2_tiehi _27585__1548 (.L_HI(net1548));
 sg13g2_tiehi _29092__1549 (.L_HI(net1549));
 sg13g2_tiehi _27584__1550 (.L_HI(net1550));
 sg13g2_tiehi _29091__1551 (.L_HI(net1551));
 sg13g2_tiehi _27582__1552 (.L_HI(net1552));
 sg13g2_tiehi _29090__1553 (.L_HI(net1553));
 sg13g2_tiehi _27581__1554 (.L_HI(net1554));
 sg13g2_tiehi _27580__1555 (.L_HI(net1555));
 sg13g2_tiehi _27579__1556 (.L_HI(net1556));
 sg13g2_tiehi _27578__1557 (.L_HI(net1557));
 sg13g2_tiehi _27577__1558 (.L_HI(net1558));
 sg13g2_tiehi _27576__1559 (.L_HI(net1559));
 sg13g2_tiehi _27575__1560 (.L_HI(net1560));
 sg13g2_tiehi _27574__1561 (.L_HI(net1561));
 sg13g2_tiehi _27573__1562 (.L_HI(net1562));
 sg13g2_tiehi _27572__1563 (.L_HI(net1563));
 sg13g2_tiehi _27571__1564 (.L_HI(net1564));
 sg13g2_tiehi _27570__1565 (.L_HI(net1565));
 sg13g2_tiehi _27569__1566 (.L_HI(net1566));
 sg13g2_tiehi _27568__1567 (.L_HI(net1567));
 sg13g2_tiehi _27567__1568 (.L_HI(net1568));
 sg13g2_tiehi _27566__1569 (.L_HI(net1569));
 sg13g2_tiehi _27565__1570 (.L_HI(net1570));
 sg13g2_tiehi _27564__1571 (.L_HI(net1571));
 sg13g2_tiehi _27563__1572 (.L_HI(net1572));
 sg13g2_tiehi _27562__1573 (.L_HI(net1573));
 sg13g2_tiehi _27561__1574 (.L_HI(net1574));
 sg13g2_tiehi _27560__1575 (.L_HI(net1575));
 sg13g2_tiehi _27559__1576 (.L_HI(net1576));
 sg13g2_tiehi _27558__1577 (.L_HI(net1577));
 sg13g2_tiehi _27557__1578 (.L_HI(net1578));
 sg13g2_tiehi _27556__1579 (.L_HI(net1579));
 sg13g2_tiehi _27555__1580 (.L_HI(net1580));
 sg13g2_tiehi _27554__1581 (.L_HI(net1581));
 sg13g2_tiehi _27553__1582 (.L_HI(net1582));
 sg13g2_tiehi _27552__1583 (.L_HI(net1583));
 sg13g2_tiehi _27551__1584 (.L_HI(net1584));
 sg13g2_tiehi _27550__1585 (.L_HI(net1585));
 sg13g2_tiehi _27549__1586 (.L_HI(net1586));
 sg13g2_tiehi _27548__1587 (.L_HI(net1587));
 sg13g2_tiehi _27547__1588 (.L_HI(net1588));
 sg13g2_tiehi _27546__1589 (.L_HI(net1589));
 sg13g2_tiehi _27545__1590 (.L_HI(net1590));
 sg13g2_tiehi _27544__1591 (.L_HI(net1591));
 sg13g2_tiehi _27543__1592 (.L_HI(net1592));
 sg13g2_tiehi _27542__1593 (.L_HI(net1593));
 sg13g2_tiehi _27541__1594 (.L_HI(net1594));
 sg13g2_tiehi _27540__1595 (.L_HI(net1595));
 sg13g2_tiehi _27539__1596 (.L_HI(net1596));
 sg13g2_tiehi _27538__1597 (.L_HI(net1597));
 sg13g2_tiehi _27537__1598 (.L_HI(net1598));
 sg13g2_tiehi _27536__1599 (.L_HI(net1599));
 sg13g2_tiehi _27535__1600 (.L_HI(net1600));
 sg13g2_tiehi _27534__1601 (.L_HI(net1601));
 sg13g2_tiehi _27533__1602 (.L_HI(net1602));
 sg13g2_tiehi _27532__1603 (.L_HI(net1603));
 sg13g2_tiehi _27531__1604 (.L_HI(net1604));
 sg13g2_tiehi _27530__1605 (.L_HI(net1605));
 sg13g2_tiehi _27529__1606 (.L_HI(net1606));
 sg13g2_tiehi _27528__1607 (.L_HI(net1607));
 sg13g2_tiehi _27527__1608 (.L_HI(net1608));
 sg13g2_tiehi _27526__1609 (.L_HI(net1609));
 sg13g2_tiehi _27525__1610 (.L_HI(net1610));
 sg13g2_tiehi _27524__1611 (.L_HI(net1611));
 sg13g2_tiehi _27523__1612 (.L_HI(net1612));
 sg13g2_tiehi _27522__1613 (.L_HI(net1613));
 sg13g2_tiehi _27521__1614 (.L_HI(net1614));
 sg13g2_tiehi _27520__1615 (.L_HI(net1615));
 sg13g2_tiehi _27519__1616 (.L_HI(net1616));
 sg13g2_tiehi _27518__1617 (.L_HI(net1617));
 sg13g2_tiehi _27517__1618 (.L_HI(net1618));
 sg13g2_tiehi _27516__1619 (.L_HI(net1619));
 sg13g2_tiehi _27515__1620 (.L_HI(net1620));
 sg13g2_tiehi _27514__1621 (.L_HI(net1621));
 sg13g2_tiehi _27513__1622 (.L_HI(net1622));
 sg13g2_tiehi _27512__1623 (.L_HI(net1623));
 sg13g2_tiehi _27511__1624 (.L_HI(net1624));
 sg13g2_tiehi _27510__1625 (.L_HI(net1625));
 sg13g2_tiehi _27509__1626 (.L_HI(net1626));
 sg13g2_tiehi _27508__1627 (.L_HI(net1627));
 sg13g2_tiehi _27507__1628 (.L_HI(net1628));
 sg13g2_tiehi _27506__1629 (.L_HI(net1629));
 sg13g2_tiehi _27505__1630 (.L_HI(net1630));
 sg13g2_tiehi _27504__1631 (.L_HI(net1631));
 sg13g2_tiehi _29089__1632 (.L_HI(net1632));
 sg13g2_tiehi _27503__1633 (.L_HI(net1633));
 sg13g2_tiehi _29088__1634 (.L_HI(net1634));
 sg13g2_tiehi _27104__1635 (.L_HI(net1635));
 sg13g2_tiehi _27501__1636 (.L_HI(net1636));
 sg13g2_tiehi _27500__1637 (.L_HI(net1637));
 sg13g2_tiehi _27499__1638 (.L_HI(net1638));
 sg13g2_tiehi _27498__1639 (.L_HI(net1639));
 sg13g2_tiehi _27497__1640 (.L_HI(net1640));
 sg13g2_tiehi _27496__1641 (.L_HI(net1641));
 sg13g2_tiehi _27495__1642 (.L_HI(net1642));
 sg13g2_tiehi _27494__1643 (.L_HI(net1643));
 sg13g2_tiehi _27493__1644 (.L_HI(net1644));
 sg13g2_tiehi _27492__1645 (.L_HI(net1645));
 sg13g2_tiehi _27491__1646 (.L_HI(net1646));
 sg13g2_tiehi _27490__1647 (.L_HI(net1647));
 sg13g2_tiehi _27489__1648 (.L_HI(net1648));
 sg13g2_tiehi _27488__1649 (.L_HI(net1649));
 sg13g2_tiehi _27487__1650 (.L_HI(net1650));
 sg13g2_tiehi _27486__1651 (.L_HI(net1651));
 sg13g2_tiehi _27485__1652 (.L_HI(net1652));
 sg13g2_tiehi _27484__1653 (.L_HI(net1653));
 sg13g2_tiehi _27483__1654 (.L_HI(net1654));
 sg13g2_tiehi _27482__1655 (.L_HI(net1655));
 sg13g2_tiehi _27481__1656 (.L_HI(net1656));
 sg13g2_tiehi _27480__1657 (.L_HI(net1657));
 sg13g2_tiehi _27479__1658 (.L_HI(net1658));
 sg13g2_tiehi _27478__1659 (.L_HI(net1659));
 sg13g2_tiehi _27477__1660 (.L_HI(net1660));
 sg13g2_tiehi _27476__1661 (.L_HI(net1661));
 sg13g2_tiehi _27475__1662 (.L_HI(net1662));
 sg13g2_tiehi _27474__1663 (.L_HI(net1663));
 sg13g2_tiehi _27473__1664 (.L_HI(net1664));
 sg13g2_tiehi _27472__1665 (.L_HI(net1665));
 sg13g2_tiehi _27471__1666 (.L_HI(net1666));
 sg13g2_tiehi _27470__1667 (.L_HI(net1667));
 sg13g2_tiehi _27469__1668 (.L_HI(net1668));
 sg13g2_tiehi _27468__1669 (.L_HI(net1669));
 sg13g2_tiehi _27467__1670 (.L_HI(net1670));
 sg13g2_tiehi _27466__1671 (.L_HI(net1671));
 sg13g2_tiehi _27465__1672 (.L_HI(net1672));
 sg13g2_tiehi _27464__1673 (.L_HI(net1673));
 sg13g2_tiehi _27463__1674 (.L_HI(net1674));
 sg13g2_tiehi _27462__1675 (.L_HI(net1675));
 sg13g2_tiehi _27461__1676 (.L_HI(net1676));
 sg13g2_tiehi _27460__1677 (.L_HI(net1677));
 sg13g2_tiehi _27459__1678 (.L_HI(net1678));
 sg13g2_tiehi _27458__1679 (.L_HI(net1679));
 sg13g2_tiehi _27457__1680 (.L_HI(net1680));
 sg13g2_tiehi _27456__1681 (.L_HI(net1681));
 sg13g2_tiehi _27455__1682 (.L_HI(net1682));
 sg13g2_tiehi _27454__1683 (.L_HI(net1683));
 sg13g2_tiehi _27453__1684 (.L_HI(net1684));
 sg13g2_tiehi _27452__1685 (.L_HI(net1685));
 sg13g2_tiehi _27451__1686 (.L_HI(net1686));
 sg13g2_tiehi _27450__1687 (.L_HI(net1687));
 sg13g2_tiehi _27449__1688 (.L_HI(net1688));
 sg13g2_tiehi _27448__1689 (.L_HI(net1689));
 sg13g2_tiehi _27447__1690 (.L_HI(net1690));
 sg13g2_tiehi _27446__1691 (.L_HI(net1691));
 sg13g2_tiehi _27445__1692 (.L_HI(net1692));
 sg13g2_tiehi _27444__1693 (.L_HI(net1693));
 sg13g2_tiehi _27443__1694 (.L_HI(net1694));
 sg13g2_tiehi _27442__1695 (.L_HI(net1695));
 sg13g2_tiehi _27441__1696 (.L_HI(net1696));
 sg13g2_tiehi _27440__1697 (.L_HI(net1697));
 sg13g2_tiehi _27439__1698 (.L_HI(net1698));
 sg13g2_tiehi _27438__1699 (.L_HI(net1699));
 sg13g2_tiehi _27437__1700 (.L_HI(net1700));
 sg13g2_tiehi _27436__1701 (.L_HI(net1701));
 sg13g2_tiehi _27435__1702 (.L_HI(net1702));
 sg13g2_tiehi _27434__1703 (.L_HI(net1703));
 sg13g2_tiehi _27433__1704 (.L_HI(net1704));
 sg13g2_tiehi _27432__1705 (.L_HI(net1705));
 sg13g2_tiehi _27431__1706 (.L_HI(net1706));
 sg13g2_tiehi _27430__1707 (.L_HI(net1707));
 sg13g2_tiehi _27429__1708 (.L_HI(net1708));
 sg13g2_tiehi _27428__1709 (.L_HI(net1709));
 sg13g2_tiehi _27427__1710 (.L_HI(net1710));
 sg13g2_tiehi _27426__1711 (.L_HI(net1711));
 sg13g2_tiehi _27425__1712 (.L_HI(net1712));
 sg13g2_tiehi _27424__1713 (.L_HI(net1713));
 sg13g2_tiehi _27423__1714 (.L_HI(net1714));
 sg13g2_tiehi _27422__1715 (.L_HI(net1715));
 sg13g2_tiehi _27421__1716 (.L_HI(net1716));
 sg13g2_tiehi _27502__1717 (.L_HI(net1717));
 sg13g2_tiehi _27420__1718 (.L_HI(net1718));
 sg13g2_tiehi _27419__1719 (.L_HI(net1719));
 sg13g2_tiehi _27418__1720 (.L_HI(net1720));
 sg13g2_tiehi _27417__1721 (.L_HI(net1721));
 sg13g2_tiehi _27416__1722 (.L_HI(net1722));
 sg13g2_tiehi _27415__1723 (.L_HI(net1723));
 sg13g2_tiehi _27414__1724 (.L_HI(net1724));
 sg13g2_tiehi _27413__1725 (.L_HI(net1725));
 sg13g2_tiehi _27412__1726 (.L_HI(net1726));
 sg13g2_tiehi _27411__1727 (.L_HI(net1727));
 sg13g2_tiehi _27410__1728 (.L_HI(net1728));
 sg13g2_tiehi _27409__1729 (.L_HI(net1729));
 sg13g2_tiehi _27408__1730 (.L_HI(net1730));
 sg13g2_tiehi _27407__1731 (.L_HI(net1731));
 sg13g2_tiehi _27406__1732 (.L_HI(net1732));
 sg13g2_tiehi _27405__1733 (.L_HI(net1733));
 sg13g2_tiehi _27404__1734 (.L_HI(net1734));
 sg13g2_tiehi _27403__1735 (.L_HI(net1735));
 sg13g2_tiehi _27402__1736 (.L_HI(net1736));
 sg13g2_tiehi _27401__1737 (.L_HI(net1737));
 sg13g2_tiehi _27400__1738 (.L_HI(net1738));
 sg13g2_tiehi _27399__1739 (.L_HI(net1739));
 sg13g2_tiehi _27398__1740 (.L_HI(net1740));
 sg13g2_tiehi _27397__1741 (.L_HI(net1741));
 sg13g2_tiehi _27396__1742 (.L_HI(net1742));
 sg13g2_tiehi _27395__1743 (.L_HI(net1743));
 sg13g2_tiehi _27394__1744 (.L_HI(net1744));
 sg13g2_tiehi _27393__1745 (.L_HI(net1745));
 sg13g2_tiehi _27392__1746 (.L_HI(net1746));
 sg13g2_tiehi _27391__1747 (.L_HI(net1747));
 sg13g2_tiehi _27390__1748 (.L_HI(net1748));
 sg13g2_tiehi _27389__1749 (.L_HI(net1749));
 sg13g2_tiehi _27388__1750 (.L_HI(net1750));
 sg13g2_tiehi _27387__1751 (.L_HI(net1751));
 sg13g2_tiehi _27386__1752 (.L_HI(net1752));
 sg13g2_tiehi _27385__1753 (.L_HI(net1753));
 sg13g2_tiehi _27384__1754 (.L_HI(net1754));
 sg13g2_tiehi _27383__1755 (.L_HI(net1755));
 sg13g2_tiehi _27382__1756 (.L_HI(net1756));
 sg13g2_tiehi _27381__1757 (.L_HI(net1757));
 sg13g2_tiehi _27380__1758 (.L_HI(net1758));
 sg13g2_tiehi _27379__1759 (.L_HI(net1759));
 sg13g2_tiehi _27378__1760 (.L_HI(net1760));
 sg13g2_tiehi _27377__1761 (.L_HI(net1761));
 sg13g2_tiehi _27376__1762 (.L_HI(net1762));
 sg13g2_tiehi _27375__1763 (.L_HI(net1763));
 sg13g2_tiehi _27374__1764 (.L_HI(net1764));
 sg13g2_tiehi _27373__1765 (.L_HI(net1765));
 sg13g2_tiehi _27372__1766 (.L_HI(net1766));
 sg13g2_tiehi _27371__1767 (.L_HI(net1767));
 sg13g2_tiehi _27370__1768 (.L_HI(net1768));
 sg13g2_tiehi _27369__1769 (.L_HI(net1769));
 sg13g2_tiehi _27368__1770 (.L_HI(net1770));
 sg13g2_tiehi _27367__1771 (.L_HI(net1771));
 sg13g2_tiehi _27366__1772 (.L_HI(net1772));
 sg13g2_tiehi _27365__1773 (.L_HI(net1773));
 sg13g2_tiehi _27364__1774 (.L_HI(net1774));
 sg13g2_tiehi _27363__1775 (.L_HI(net1775));
 sg13g2_tiehi _27362__1776 (.L_HI(net1776));
 sg13g2_tiehi _27361__1777 (.L_HI(net1777));
 sg13g2_tiehi _27360__1778 (.L_HI(net1778));
 sg13g2_tiehi _27359__1779 (.L_HI(net1779));
 sg13g2_tiehi _27358__1780 (.L_HI(net1780));
 sg13g2_tiehi _27357__1781 (.L_HI(net1781));
 sg13g2_tiehi _27356__1782 (.L_HI(net1782));
 sg13g2_tiehi _27583__1783 (.L_HI(net1783));
 sg13g2_tiehi _27649__1784 (.L_HI(net1784));
 sg13g2_tiehi _27355__1785 (.L_HI(net1785));
 sg13g2_tiehi _27354__1786 (.L_HI(net1786));
 sg13g2_tiehi _27353__1787 (.L_HI(net1787));
 sg13g2_tiehi _27352__1788 (.L_HI(net1788));
 sg13g2_tiehi _27351__1789 (.L_HI(net1789));
 sg13g2_tiehi _27350__1790 (.L_HI(net1790));
 sg13g2_tiehi _27349__1791 (.L_HI(net1791));
 sg13g2_tiehi _27348__1792 (.L_HI(net1792));
 sg13g2_tiehi _27347__1793 (.L_HI(net1793));
 sg13g2_tiehi _27346__1794 (.L_HI(net1794));
 sg13g2_tiehi _27345__1795 (.L_HI(net1795));
 sg13g2_tiehi _27344__1796 (.L_HI(net1796));
 sg13g2_tiehi _27343__1797 (.L_HI(net1797));
 sg13g2_tiehi _27342__1798 (.L_HI(net1798));
 sg13g2_tiehi _27341__1799 (.L_HI(net1799));
 sg13g2_tiehi _27340__1800 (.L_HI(net1800));
 sg13g2_tiehi _27339__1801 (.L_HI(net1801));
 sg13g2_tiehi _27338__1802 (.L_HI(net1802));
 sg13g2_tiehi _27337__1803 (.L_HI(net1803));
 sg13g2_tiehi _27336__1804 (.L_HI(net1804));
 sg13g2_tiehi _27335__1805 (.L_HI(net1805));
 sg13g2_tiehi _27334__1806 (.L_HI(net1806));
 sg13g2_tiehi _27333__1807 (.L_HI(net1807));
 sg13g2_tiehi _27332__1808 (.L_HI(net1808));
 sg13g2_tiehi _27331__1809 (.L_HI(net1809));
 sg13g2_tiehi _27330__1810 (.L_HI(net1810));
 sg13g2_tiehi _27329__1811 (.L_HI(net1811));
 sg13g2_tiehi _27328__1812 (.L_HI(net1812));
 sg13g2_tiehi _27327__1813 (.L_HI(net1813));
 sg13g2_tiehi _27326__1814 (.L_HI(net1814));
 sg13g2_tiehi _27325__1815 (.L_HI(net1815));
 sg13g2_tiehi _27324__1816 (.L_HI(net1816));
 sg13g2_tiehi _27323__1817 (.L_HI(net1817));
 sg13g2_tiehi _27322__1818 (.L_HI(net1818));
 sg13g2_tiehi _27321__1819 (.L_HI(net1819));
 sg13g2_tiehi _27320__1820 (.L_HI(net1820));
 sg13g2_tiehi _27319__1821 (.L_HI(net1821));
 sg13g2_tiehi _27318__1822 (.L_HI(net1822));
 sg13g2_tiehi _27317__1823 (.L_HI(net1823));
 sg13g2_tiehi _27316__1824 (.L_HI(net1824));
 sg13g2_tiehi _27315__1825 (.L_HI(net1825));
 sg13g2_tiehi _27314__1826 (.L_HI(net1826));
 sg13g2_tiehi _27313__1827 (.L_HI(net1827));
 sg13g2_tiehi _27312__1828 (.L_HI(net1828));
 sg13g2_tiehi _27311__1829 (.L_HI(net1829));
 sg13g2_tiehi _27310__1830 (.L_HI(net1830));
 sg13g2_tiehi _27309__1831 (.L_HI(net1831));
 sg13g2_tiehi _27308__1832 (.L_HI(net1832));
 sg13g2_tiehi _27307__1833 (.L_HI(net1833));
 sg13g2_tiehi _27306__1834 (.L_HI(net1834));
 sg13g2_tiehi _27305__1835 (.L_HI(net1835));
 sg13g2_tiehi _27304__1836 (.L_HI(net1836));
 sg13g2_tiehi _27303__1837 (.L_HI(net1837));
 sg13g2_tiehi _27302__1838 (.L_HI(net1838));
 sg13g2_tiehi _27301__1839 (.L_HI(net1839));
 sg13g2_tiehi _27300__1840 (.L_HI(net1840));
 sg13g2_tiehi _27299__1841 (.L_HI(net1841));
 sg13g2_tiehi _27298__1842 (.L_HI(net1842));
 sg13g2_tiehi _27297__1843 (.L_HI(net1843));
 sg13g2_tiehi _27296__1844 (.L_HI(net1844));
 sg13g2_tiehi _27295__1845 (.L_HI(net1845));
 sg13g2_tiehi _27294__1846 (.L_HI(net1846));
 sg13g2_tiehi _27293__1847 (.L_HI(net1847));
 sg13g2_tiehi _27292__1848 (.L_HI(net1848));
 sg13g2_tiehi _27291__1849 (.L_HI(net1849));
 sg13g2_tiehi _27290__1850 (.L_HI(net1850));
 sg13g2_tiehi _27289__1851 (.L_HI(net1851));
 sg13g2_tiehi _27288__1852 (.L_HI(net1852));
 sg13g2_tiehi _27287__1853 (.L_HI(net1853));
 sg13g2_tiehi _27286__1854 (.L_HI(net1854));
 sg13g2_tiehi _27285__1855 (.L_HI(net1855));
 sg13g2_tiehi _27284__1856 (.L_HI(net1856));
 sg13g2_tiehi _27283__1857 (.L_HI(net1857));
 sg13g2_tiehi _27282__1858 (.L_HI(net1858));
 sg13g2_tiehi _27281__1859 (.L_HI(net1859));
 sg13g2_tiehi _27280__1860 (.L_HI(net1860));
 sg13g2_tiehi _27279__1861 (.L_HI(net1861));
 sg13g2_tiehi _27278__1862 (.L_HI(net1862));
 sg13g2_tiehi _27277__1863 (.L_HI(net1863));
 sg13g2_tiehi _27276__1864 (.L_HI(net1864));
 sg13g2_tiehi _27275__1865 (.L_HI(net1865));
 sg13g2_tiehi _27274__1866 (.L_HI(net1866));
 sg13g2_tiehi _27273__1867 (.L_HI(net1867));
 sg13g2_tiehi _27272__1868 (.L_HI(net1868));
 sg13g2_tiehi _27271__1869 (.L_HI(net1869));
 sg13g2_tiehi _27270__1870 (.L_HI(net1870));
 sg13g2_tiehi _27269__1871 (.L_HI(net1871));
 sg13g2_tiehi _27268__1872 (.L_HI(net1872));
 sg13g2_tiehi _27267__1873 (.L_HI(net1873));
 sg13g2_tiehi _27266__1874 (.L_HI(net1874));
 sg13g2_tiehi _27265__1875 (.L_HI(net1875));
 sg13g2_tiehi _27264__1876 (.L_HI(net1876));
 sg13g2_tiehi _27263__1877 (.L_HI(net1877));
 sg13g2_tiehi _27262__1878 (.L_HI(net1878));
 sg13g2_tiehi _27261__1879 (.L_HI(net1879));
 sg13g2_tiehi _27260__1880 (.L_HI(net1880));
 sg13g2_tiehi _27259__1881 (.L_HI(net1881));
 sg13g2_tiehi _27258__1882 (.L_HI(net1882));
 sg13g2_tiehi _27257__1883 (.L_HI(net1883));
 sg13g2_tiehi _27256__1884 (.L_HI(net1884));
 sg13g2_tiehi _27255__1885 (.L_HI(net1885));
 sg13g2_tiehi _27254__1886 (.L_HI(net1886));
 sg13g2_tiehi _27253__1887 (.L_HI(net1887));
 sg13g2_tiehi _27252__1888 (.L_HI(net1888));
 sg13g2_tiehi _27251__1889 (.L_HI(net1889));
 sg13g2_tiehi _27250__1890 (.L_HI(net1890));
 sg13g2_tiehi _27249__1891 (.L_HI(net1891));
 sg13g2_tiehi _27248__1892 (.L_HI(net1892));
 sg13g2_tiehi _27247__1893 (.L_HI(net1893));
 sg13g2_tiehi _27246__1894 (.L_HI(net1894));
 sg13g2_tiehi _27245__1895 (.L_HI(net1895));
 sg13g2_tiehi _27244__1896 (.L_HI(net1896));
 sg13g2_tiehi _27243__1897 (.L_HI(net1897));
 sg13g2_tiehi _27242__1898 (.L_HI(net1898));
 sg13g2_tiehi _27241__1899 (.L_HI(net1899));
 sg13g2_tiehi _27240__1900 (.L_HI(net1900));
 sg13g2_tiehi _27239__1901 (.L_HI(net1901));
 sg13g2_tiehi _27238__1902 (.L_HI(net1902));
 sg13g2_tiehi _27237__1903 (.L_HI(net1903));
 sg13g2_tiehi _27236__1904 (.L_HI(net1904));
 sg13g2_tiehi _27235__1905 (.L_HI(net1905));
 sg13g2_tiehi _27234__1906 (.L_HI(net1906));
 sg13g2_tiehi _27233__1907 (.L_HI(net1907));
 sg13g2_tiehi _27232__1908 (.L_HI(net1908));
 sg13g2_tiehi _27231__1909 (.L_HI(net1909));
 sg13g2_tiehi _27230__1910 (.L_HI(net1910));
 sg13g2_tiehi _27229__1911 (.L_HI(net1911));
 sg13g2_tiehi _27228__1912 (.L_HI(net1912));
 sg13g2_tiehi _27227__1913 (.L_HI(net1913));
 sg13g2_tiehi _27226__1914 (.L_HI(net1914));
 sg13g2_tiehi _27225__1915 (.L_HI(net1915));
 sg13g2_tiehi _27224__1916 (.L_HI(net1916));
 sg13g2_tiehi _27223__1917 (.L_HI(net1917));
 sg13g2_tiehi _27222__1918 (.L_HI(net1918));
 sg13g2_tiehi _27221__1919 (.L_HI(net1919));
 sg13g2_tiehi _27220__1920 (.L_HI(net1920));
 sg13g2_tiehi _27219__1921 (.L_HI(net1921));
 sg13g2_tiehi _27218__1922 (.L_HI(net1922));
 sg13g2_tiehi _27217__1923 (.L_HI(net1923));
 sg13g2_tiehi _27216__1924 (.L_HI(net1924));
 sg13g2_tiehi _27215__1925 (.L_HI(net1925));
 sg13g2_tiehi _27214__1926 (.L_HI(net1926));
 sg13g2_tiehi _27213__1927 (.L_HI(net1927));
 sg13g2_tiehi _27212__1928 (.L_HI(net1928));
 sg13g2_tiehi _27211__1929 (.L_HI(net1929));
 sg13g2_tiehi _27210__1930 (.L_HI(net1930));
 sg13g2_tiehi _27209__1931 (.L_HI(net1931));
 sg13g2_tiehi _27208__1932 (.L_HI(net1932));
 sg13g2_tiehi _27207__1933 (.L_HI(net1933));
 sg13g2_tiehi _27206__1934 (.L_HI(net1934));
 sg13g2_tiehi _27205__1935 (.L_HI(net1935));
 sg13g2_tiehi _27204__1936 (.L_HI(net1936));
 sg13g2_tiehi _27203__1937 (.L_HI(net1937));
 sg13g2_tiehi _27202__1938 (.L_HI(net1938));
 sg13g2_tiehi _27201__1939 (.L_HI(net1939));
 sg13g2_tiehi _27200__1940 (.L_HI(net1940));
 sg13g2_tiehi _27199__1941 (.L_HI(net1941));
 sg13g2_tiehi _27198__1942 (.L_HI(net1942));
 sg13g2_tiehi _27197__1943 (.L_HI(net1943));
 sg13g2_tiehi _27196__1944 (.L_HI(net1944));
 sg13g2_tiehi _27195__1945 (.L_HI(net1945));
 sg13g2_tiehi _27194__1946 (.L_HI(net1946));
 sg13g2_tiehi _27193__1947 (.L_HI(net1947));
 sg13g2_tiehi _27192__1948 (.L_HI(net1948));
 sg13g2_tiehi _27191__1949 (.L_HI(net1949));
 sg13g2_tiehi _27190__1950 (.L_HI(net1950));
 sg13g2_tiehi _27189__1951 (.L_HI(net1951));
 sg13g2_tiehi _27188__1952 (.L_HI(net1952));
 sg13g2_tiehi _27187__1953 (.L_HI(net1953));
 sg13g2_tiehi _27186__1954 (.L_HI(net1954));
 sg13g2_tiehi _27185__1955 (.L_HI(net1955));
 sg13g2_tiehi _27184__1956 (.L_HI(net1956));
 sg13g2_tiehi _27183__1957 (.L_HI(net1957));
 sg13g2_tiehi _27182__1958 (.L_HI(net1958));
 sg13g2_tiehi _27181__1959 (.L_HI(net1959));
 sg13g2_tiehi _27180__1960 (.L_HI(net1960));
 sg13g2_tiehi _27179__1961 (.L_HI(net1961));
 sg13g2_tiehi _27178__1962 (.L_HI(net1962));
 sg13g2_tiehi _27177__1963 (.L_HI(net1963));
 sg13g2_tiehi _27176__1964 (.L_HI(net1964));
 sg13g2_tiehi _27175__1965 (.L_HI(net1965));
 sg13g2_tiehi _27174__1966 (.L_HI(net1966));
 sg13g2_tiehi _27173__1967 (.L_HI(net1967));
 sg13g2_tiehi _27172__1968 (.L_HI(net1968));
 sg13g2_tiehi _27171__1969 (.L_HI(net1969));
 sg13g2_tiehi _27170__1970 (.L_HI(net1970));
 sg13g2_tiehi _27169__1971 (.L_HI(net1971));
 sg13g2_tiehi _27168__1972 (.L_HI(net1972));
 sg13g2_tiehi _27167__1973 (.L_HI(net1973));
 sg13g2_tiehi _27166__1974 (.L_HI(net1974));
 sg13g2_tiehi _27165__1975 (.L_HI(net1975));
 sg13g2_tiehi _27164__1976 (.L_HI(net1976));
 sg13g2_tiehi _27163__1977 (.L_HI(net1977));
 sg13g2_tiehi _27162__1978 (.L_HI(net1978));
 sg13g2_tiehi _27161__1979 (.L_HI(net1979));
 sg13g2_tiehi _27160__1980 (.L_HI(net1980));
 sg13g2_tiehi _27159__1981 (.L_HI(net1981));
 sg13g2_tiehi _27158__1982 (.L_HI(net1982));
 sg13g2_tiehi _27157__1983 (.L_HI(net1983));
 sg13g2_tiehi _27156__1984 (.L_HI(net1984));
 sg13g2_tiehi _27155__1985 (.L_HI(net1985));
 sg13g2_tiehi _27154__1986 (.L_HI(net1986));
 sg13g2_tiehi _27153__1987 (.L_HI(net1987));
 sg13g2_tiehi _27152__1988 (.L_HI(net1988));
 sg13g2_tiehi _27151__1989 (.L_HI(net1989));
 sg13g2_tiehi _27150__1990 (.L_HI(net1990));
 sg13g2_tiehi _27149__1991 (.L_HI(net1991));
 sg13g2_tiehi _27148__1992 (.L_HI(net1992));
 sg13g2_tiehi _27147__1993 (.L_HI(net1993));
 sg13g2_tiehi _27146__1994 (.L_HI(net1994));
 sg13g2_tiehi _27145__1995 (.L_HI(net1995));
 sg13g2_tiehi _27144__1996 (.L_HI(net1996));
 sg13g2_tiehi _27143__1997 (.L_HI(net1997));
 sg13g2_tiehi _27142__1998 (.L_HI(net1998));
 sg13g2_tiehi _27141__1999 (.L_HI(net1999));
 sg13g2_tiehi _27140__2000 (.L_HI(net2000));
 sg13g2_tiehi _27139__2001 (.L_HI(net2001));
 sg13g2_tiehi _27138__2002 (.L_HI(net2002));
 sg13g2_tiehi _27137__2003 (.L_HI(net2003));
 sg13g2_tiehi _27136__2004 (.L_HI(net2004));
 sg13g2_tiehi _27135__2005 (.L_HI(net2005));
 sg13g2_tiehi _27134__2006 (.L_HI(net2006));
 sg13g2_tiehi _27133__2007 (.L_HI(net2007));
 sg13g2_tiehi _27132__2008 (.L_HI(net2008));
 sg13g2_tiehi _27131__2009 (.L_HI(net2009));
 sg13g2_tiehi _27130__2010 (.L_HI(net2010));
 sg13g2_tiehi _27129__2011 (.L_HI(net2011));
 sg13g2_tiehi _27128__2012 (.L_HI(net2012));
 sg13g2_tiehi _27127__2013 (.L_HI(net2013));
 sg13g2_tiehi _27126__2014 (.L_HI(net2014));
 sg13g2_tiehi _27125__2015 (.L_HI(net2015));
 sg13g2_tiehi _27124__2016 (.L_HI(net2016));
 sg13g2_tiehi _27123__2017 (.L_HI(net2017));
 sg13g2_tiehi _27122__2018 (.L_HI(net2018));
 sg13g2_tiehi _27121__2019 (.L_HI(net2019));
 sg13g2_tiehi _27120__2020 (.L_HI(net2020));
 sg13g2_tiehi _27119__2021 (.L_HI(net2021));
 sg13g2_tiehi _27118__2022 (.L_HI(net2022));
 sg13g2_tiehi _27117__2023 (.L_HI(net2023));
 sg13g2_tiehi _27116__2024 (.L_HI(net2024));
 sg13g2_tiehi _27115__2025 (.L_HI(net2025));
 sg13g2_tiehi _27114__2026 (.L_HI(net2026));
 sg13g2_tiehi _27113__2027 (.L_HI(net2027));
 sg13g2_tiehi _27112__2028 (.L_HI(net2028));
 sg13g2_tiehi _27111__2029 (.L_HI(net2029));
 sg13g2_tiehi _27110__2030 (.L_HI(net2030));
 sg13g2_tiehi _27109__2031 (.L_HI(net2031));
 sg13g2_tiehi _27108__2032 (.L_HI(net2032));
 sg13g2_tiehi _27107__2033 (.L_HI(net2033));
 sg13g2_tiehi _27106__2034 (.L_HI(net2034));
 sg13g2_tiehi _27105__2035 (.L_HI(net2035));
 sg13g2_tiehi _27096__2036 (.L_HI(net2036));
 sg13g2_tiehi _27095__2037 (.L_HI(net2037));
 sg13g2_tiehi _27094__2038 (.L_HI(net2038));
 sg13g2_tiehi _27093__2039 (.L_HI(net2039));
 sg13g2_tiehi _27092__2040 (.L_HI(net2040));
 sg13g2_tiehi _27091__2041 (.L_HI(net2041));
 sg13g2_tiehi _27090__2042 (.L_HI(net2042));
 sg13g2_tiehi _27089__2043 (.L_HI(net2043));
 sg13g2_tiehi _27088__2044 (.L_HI(net2044));
 sg13g2_tiehi _27087__2045 (.L_HI(net2045));
 sg13g2_tiehi _27086__2046 (.L_HI(net2046));
 sg13g2_tiehi _27085__2047 (.L_HI(net2047));
 sg13g2_tiehi _27084__2048 (.L_HI(net2048));
 sg13g2_tiehi _27083__2049 (.L_HI(net2049));
 sg13g2_tiehi _27082__2050 (.L_HI(net2050));
 sg13g2_tiehi _27081__2051 (.L_HI(net2051));
 sg13g2_tiehi _27080__2052 (.L_HI(net2052));
 sg13g2_tiehi _27079__2053 (.L_HI(net2053));
 sg13g2_tiehi _27078__2054 (.L_HI(net2054));
 sg13g2_tiehi _27077__2055 (.L_HI(net2055));
 sg13g2_tiehi _27076__2056 (.L_HI(net2056));
 sg13g2_tiehi _27075__2057 (.L_HI(net2057));
 sg13g2_tiehi _27074__2058 (.L_HI(net2058));
 sg13g2_tiehi _27073__2059 (.L_HI(net2059));
 sg13g2_tiehi _27072__2060 (.L_HI(net2060));
 sg13g2_tiehi _27071__2061 (.L_HI(net2061));
 sg13g2_tiehi _27070__2062 (.L_HI(net2062));
 sg13g2_tiehi _27069__2063 (.L_HI(net2063));
 sg13g2_tiehi _27068__2064 (.L_HI(net2064));
 sg13g2_tiehi _27067__2065 (.L_HI(net2065));
 sg13g2_tiehi _27066__2066 (.L_HI(net2066));
 sg13g2_tiehi _27065__2067 (.L_HI(net2067));
 sg13g2_tiehi _27064__2068 (.L_HI(net2068));
 sg13g2_tiehi _27063__2069 (.L_HI(net2069));
 sg13g2_tiehi _27062__2070 (.L_HI(net2070));
 sg13g2_tiehi _27061__2071 (.L_HI(net2071));
 sg13g2_tiehi _27060__2072 (.L_HI(net2072));
 sg13g2_tiehi _27059__2073 (.L_HI(net2073));
 sg13g2_tiehi _27058__2074 (.L_HI(net2074));
 sg13g2_tiehi _27057__2075 (.L_HI(net2075));
 sg13g2_tiehi _27056__2076 (.L_HI(net2076));
 sg13g2_tiehi _27055__2077 (.L_HI(net2077));
 sg13g2_tiehi _27054__2078 (.L_HI(net2078));
 sg13g2_tiehi _27053__2079 (.L_HI(net2079));
 sg13g2_tiehi _27052__2080 (.L_HI(net2080));
 sg13g2_tiehi _27051__2081 (.L_HI(net2081));
 sg13g2_tiehi _27050__2082 (.L_HI(net2082));
 sg13g2_tiehi _27049__2083 (.L_HI(net2083));
 sg13g2_tiehi _27048__2084 (.L_HI(net2084));
 sg13g2_tiehi _27047__2085 (.L_HI(net2085));
 sg13g2_tiehi _27046__2086 (.L_HI(net2086));
 sg13g2_tiehi _27045__2087 (.L_HI(net2087));
 sg13g2_tiehi _27044__2088 (.L_HI(net2088));
 sg13g2_tiehi _27043__2089 (.L_HI(net2089));
 sg13g2_tiehi _27042__2090 (.L_HI(net2090));
 sg13g2_tiehi _27041__2091 (.L_HI(net2091));
 sg13g2_tiehi _27040__2092 (.L_HI(net2092));
 sg13g2_tiehi _27039__2093 (.L_HI(net2093));
 sg13g2_tiehi _27038__2094 (.L_HI(net2094));
 sg13g2_tiehi _27037__2095 (.L_HI(net2095));
 sg13g2_tiehi _27036__2096 (.L_HI(net2096));
 sg13g2_tiehi _27035__2097 (.L_HI(net2097));
 sg13g2_tiehi _27034__2098 (.L_HI(net2098));
 sg13g2_tiehi _27033__2099 (.L_HI(net2099));
 sg13g2_tiehi _27032__2100 (.L_HI(net2100));
 sg13g2_tiehi _27031__2101 (.L_HI(net2101));
 sg13g2_tiehi _27030__2102 (.L_HI(net2102));
 sg13g2_tiehi _27029__2103 (.L_HI(net2103));
 sg13g2_tiehi _27028__2104 (.L_HI(net2104));
 sg13g2_tiehi _27027__2105 (.L_HI(net2105));
 sg13g2_tiehi _27026__2106 (.L_HI(net2106));
 sg13g2_tiehi _27025__2107 (.L_HI(net2107));
 sg13g2_tiehi _27024__2108 (.L_HI(net2108));
 sg13g2_tiehi _27023__2109 (.L_HI(net2109));
 sg13g2_tiehi _27022__2110 (.L_HI(net2110));
 sg13g2_tiehi _27021__2111 (.L_HI(net2111));
 sg13g2_tiehi _27020__2112 (.L_HI(net2112));
 sg13g2_tiehi _27019__2113 (.L_HI(net2113));
 sg13g2_tiehi _27018__2114 (.L_HI(net2114));
 sg13g2_tiehi _27017__2115 (.L_HI(net2115));
 sg13g2_tiehi _27016__2116 (.L_HI(net2116));
 sg13g2_tiehi _27015__2117 (.L_HI(net2117));
 sg13g2_tiehi _27014__2118 (.L_HI(net2118));
 sg13g2_tiehi _27013__2119 (.L_HI(net2119));
 sg13g2_tiehi _27012__2120 (.L_HI(net2120));
 sg13g2_tiehi _27011__2121 (.L_HI(net2121));
 sg13g2_tiehi _27010__2122 (.L_HI(net2122));
 sg13g2_tiehi _27009__2123 (.L_HI(net2123));
 sg13g2_tiehi _27008__2124 (.L_HI(net2124));
 sg13g2_tiehi _27007__2125 (.L_HI(net2125));
 sg13g2_tiehi _27006__2126 (.L_HI(net2126));
 sg13g2_tiehi _27005__2127 (.L_HI(net2127));
 sg13g2_tiehi _27004__2128 (.L_HI(net2128));
 sg13g2_tiehi _27003__2129 (.L_HI(net2129));
 sg13g2_tiehi _27002__2130 (.L_HI(net2130));
 sg13g2_tiehi _27001__2131 (.L_HI(net2131));
 sg13g2_tiehi _27000__2132 (.L_HI(net2132));
 sg13g2_tiehi _26999__2133 (.L_HI(net2133));
 sg13g2_tiehi _26998__2134 (.L_HI(net2134));
 sg13g2_tiehi _26997__2135 (.L_HI(net2135));
 sg13g2_tiehi _26996__2136 (.L_HI(net2136));
 sg13g2_tiehi _26995__2137 (.L_HI(net2137));
 sg13g2_tiehi _26994__2138 (.L_HI(net2138));
 sg13g2_tiehi _26993__2139 (.L_HI(net2139));
 sg13g2_tiehi _26992__2140 (.L_HI(net2140));
 sg13g2_tiehi _26991__2141 (.L_HI(net2141));
 sg13g2_tiehi _26990__2142 (.L_HI(net2142));
 sg13g2_tiehi _26989__2143 (.L_HI(net2143));
 sg13g2_tiehi _26988__2144 (.L_HI(net2144));
 sg13g2_tiehi _26987__2145 (.L_HI(net2145));
 sg13g2_tiehi _26986__2146 (.L_HI(net2146));
 sg13g2_tiehi _26985__2147 (.L_HI(net2147));
 sg13g2_tiehi _26984__2148 (.L_HI(net2148));
 sg13g2_tiehi _26983__2149 (.L_HI(net2149));
 sg13g2_tiehi _26982__2150 (.L_HI(net2150));
 sg13g2_tiehi _26981__2151 (.L_HI(net2151));
 sg13g2_tiehi _26980__2152 (.L_HI(net2152));
 sg13g2_tiehi _26979__2153 (.L_HI(net2153));
 sg13g2_tiehi _28433__2154 (.L_HI(net2154));
 sg13g2_tiehi _28434__2155 (.L_HI(net2155));
 sg13g2_tiehi _28435__2156 (.L_HI(net2156));
 sg13g2_tiehi _28436__2157 (.L_HI(net2157));
 sg13g2_tiehi _28437__2158 (.L_HI(net2158));
 sg13g2_tiehi _28438__2159 (.L_HI(net2159));
 sg13g2_tiehi _28439__2160 (.L_HI(net2160));
 sg13g2_tiehi _28440__2161 (.L_HI(net2161));
 sg13g2_tiehi _28441__2162 (.L_HI(net2162));
 sg13g2_tiehi _28442__2163 (.L_HI(net2163));
 sg13g2_tiehi _28443__2164 (.L_HI(net2164));
 sg13g2_tiehi _28444__2165 (.L_HI(net2165));
 sg13g2_tiehi _28445__2166 (.L_HI(net2166));
 sg13g2_tiehi _28446__2167 (.L_HI(net2167));
 sg13g2_tiehi _28447__2168 (.L_HI(net2168));
 sg13g2_tiehi _28448__2169 (.L_HI(net2169));
 sg13g2_tiehi _26978__2170 (.L_HI(net2170));
 sg13g2_tiehi _26977__2171 (.L_HI(net2171));
 sg13g2_tiehi _26976__2172 (.L_HI(net2172));
 sg13g2_tiehi _26975__2173 (.L_HI(net2173));
 sg13g2_tiehi _26974__2174 (.L_HI(net2174));
 sg13g2_tiehi _26973__2175 (.L_HI(net2175));
 sg13g2_tiehi _26972__2176 (.L_HI(net2176));
 sg13g2_tiehi _26971__2177 (.L_HI(net2177));
 sg13g2_tiehi _26970__2178 (.L_HI(net2178));
 sg13g2_tiehi _26969__2179 (.L_HI(net2179));
 sg13g2_tiehi _26968__2180 (.L_HI(net2180));
 sg13g2_tiehi _26967__2181 (.L_HI(net2181));
 sg13g2_tiehi _26966__2182 (.L_HI(net2182));
 sg13g2_tiehi _26965__2183 (.L_HI(net2183));
 sg13g2_tiehi _28449__2184 (.L_HI(net2184));
 sg13g2_tiehi _28599__2185 (.L_HI(net2185));
 sg13g2_tiehi _28600__2186 (.L_HI(net2186));
 sg13g2_tiehi _28601__2187 (.L_HI(net2187));
 sg13g2_tiehi _28602__2188 (.L_HI(net2188));
 sg13g2_tiehi _28603__2189 (.L_HI(net2189));
 sg13g2_tiehi _28604__2190 (.L_HI(net2190));
 sg13g2_tiehi _28605__2191 (.L_HI(net2191));
 sg13g2_tiehi _28606__2192 (.L_HI(net2192));
 sg13g2_tiehi _28607__2193 (.L_HI(net2193));
 sg13g2_tiehi _28608__2194 (.L_HI(net2194));
 sg13g2_tiehi _28609__2195 (.L_HI(net2195));
 sg13g2_tiehi _28610__2196 (.L_HI(net2196));
 sg13g2_tiehi _28611__2197 (.L_HI(net2197));
 sg13g2_tiehi _28612__2198 (.L_HI(net2198));
 sg13g2_tiehi _26964__2199 (.L_HI(net2199));
 sg13g2_tiehi _26963__2200 (.L_HI(net2200));
 sg13g2_tiehi _26962__2201 (.L_HI(net2201));
 sg13g2_tiehi _26961__2202 (.L_HI(net2202));
 sg13g2_tiehi _26960__2203 (.L_HI(net2203));
 sg13g2_tiehi _26959__2204 (.L_HI(net2204));
 sg13g2_tiehi _26958__2205 (.L_HI(net2205));
 sg13g2_tiehi _26957__2206 (.L_HI(net2206));
 sg13g2_tiehi _26956__2207 (.L_HI(net2207));
 sg13g2_tiehi _26955__2208 (.L_HI(net2208));
 sg13g2_tiehi _26954__2209 (.L_HI(net2209));
 sg13g2_tiehi _26953__2210 (.L_HI(net2210));
 sg13g2_tiehi _26952__2211 (.L_HI(net2211));
 sg13g2_tiehi _26951__2212 (.L_HI(net2212));
 sg13g2_tiehi _26950__2213 (.L_HI(net2213));
 sg13g2_tiehi _26949__2214 (.L_HI(net2214));
 sg13g2_tiehi _26948__2215 (.L_HI(net2215));
 sg13g2_tiehi _26947__2216 (.L_HI(net2216));
 sg13g2_tiehi _26946__2217 (.L_HI(net2217));
 sg13g2_tiehi _26945__2218 (.L_HI(net2218));
 sg13g2_tiehi _26944__2219 (.L_HI(net2219));
 sg13g2_tiehi _26943__2220 (.L_HI(net2220));
 sg13g2_tiehi _26942__2221 (.L_HI(net2221));
 sg13g2_tiehi _26941__2222 (.L_HI(net2222));
 sg13g2_tiehi _26940__2223 (.L_HI(net2223));
 sg13g2_tiehi _26939__2224 (.L_HI(net2224));
 sg13g2_tiehi _26938__2225 (.L_HI(net2225));
 sg13g2_tiehi _26937__2226 (.L_HI(net2226));
 sg13g2_tiehi _26936__2227 (.L_HI(net2227));
 sg13g2_tiehi _26935__2228 (.L_HI(net2228));
 sg13g2_tiehi _26934__2229 (.L_HI(net2229));
 sg13g2_tiehi _26933__2230 (.L_HI(net2230));
 sg13g2_tiehi _26932__2231 (.L_HI(net2231));
 sg13g2_tiehi _26931__2232 (.L_HI(net2232));
 sg13g2_tiehi _26930__2233 (.L_HI(net2233));
 sg13g2_tiehi _26929__2234 (.L_HI(net2234));
 sg13g2_tiehi _26928__2235 (.L_HI(net2235));
 sg13g2_tiehi _26927__2236 (.L_HI(net2236));
 sg13g2_tiehi _26926__2237 (.L_HI(net2237));
 sg13g2_tiehi _26925__2238 (.L_HI(net2238));
 sg13g2_tiehi _26924__2239 (.L_HI(net2239));
 sg13g2_tiehi _26923__2240 (.L_HI(net2240));
 sg13g2_tiehi _26922__2241 (.L_HI(net2241));
 sg13g2_tiehi _26921__2242 (.L_HI(net2242));
 sg13g2_tiehi _26920__2243 (.L_HI(net2243));
 sg13g2_tiehi _26919__2244 (.L_HI(net2244));
 sg13g2_tiehi _26918__2245 (.L_HI(net2245));
 sg13g2_tiehi _26917__2246 (.L_HI(net2246));
 sg13g2_tiehi _26916__2247 (.L_HI(net2247));
 sg13g2_tiehi _26915__2248 (.L_HI(net2248));
 sg13g2_tiehi _26914__2249 (.L_HI(net2249));
 sg13g2_tiehi _26913__2250 (.L_HI(net2250));
 sg13g2_tiehi _26912__2251 (.L_HI(net2251));
 sg13g2_tiehi _26911__2252 (.L_HI(net2252));
 sg13g2_tiehi _26910__2253 (.L_HI(net2253));
 sg13g2_tiehi _26909__2254 (.L_HI(net2254));
 sg13g2_tiehi _26908__2255 (.L_HI(net2255));
 sg13g2_tiehi _26907__2256 (.L_HI(net2256));
 sg13g2_tiehi _26906__2257 (.L_HI(net2257));
 sg13g2_tiehi _26905__2258 (.L_HI(net2258));
 sg13g2_tiehi _26904__2259 (.L_HI(net2259));
 sg13g2_tiehi _26903__2260 (.L_HI(net2260));
 sg13g2_tiehi _26902__2261 (.L_HI(net2261));
 sg13g2_tiehi _26901__2262 (.L_HI(net2262));
 sg13g2_tiehi _26900__2263 (.L_HI(net2263));
 sg13g2_tiehi _26899__2264 (.L_HI(net2264));
 sg13g2_tiehi _26898__2265 (.L_HI(net2265));
 sg13g2_tiehi _26897__2266 (.L_HI(net2266));
 sg13g2_tiehi _26896__2267 (.L_HI(net2267));
 sg13g2_tiehi _26895__2268 (.L_HI(net2268));
 sg13g2_tiehi _26894__2269 (.L_HI(net2269));
 sg13g2_tiehi _26893__2270 (.L_HI(net2270));
 sg13g2_tiehi _26892__2271 (.L_HI(net2271));
 sg13g2_tiehi _26891__2272 (.L_HI(net2272));
 sg13g2_tiehi _26890__2273 (.L_HI(net2273));
 sg13g2_tiehi _26889__2274 (.L_HI(net2274));
 sg13g2_tiehi _26888__2275 (.L_HI(net2275));
 sg13g2_tiehi _26887__2276 (.L_HI(net2276));
 sg13g2_tiehi _26886__2277 (.L_HI(net2277));
 sg13g2_tiehi _26885__2278 (.L_HI(net2278));
 sg13g2_tiehi _26884__2279 (.L_HI(net2279));
 sg13g2_tiehi _26883__2280 (.L_HI(net2280));
 sg13g2_tiehi _26882__2281 (.L_HI(net2281));
 sg13g2_tiehi _26881__2282 (.L_HI(net2282));
 sg13g2_tiehi _26880__2283 (.L_HI(net2283));
 sg13g2_tiehi _26879__2284 (.L_HI(net2284));
 sg13g2_tiehi _26878__2285 (.L_HI(net2285));
 sg13g2_tiehi _26877__2286 (.L_HI(net2286));
 sg13g2_tiehi _26876__2287 (.L_HI(net2287));
 sg13g2_tiehi _26875__2288 (.L_HI(net2288));
 sg13g2_tiehi _26874__2289 (.L_HI(net2289));
 sg13g2_tiehi _26873__2290 (.L_HI(net2290));
 sg13g2_tiehi _26872__2291 (.L_HI(net2291));
 sg13g2_tiehi _26871__2292 (.L_HI(net2292));
 sg13g2_tiehi _26870__2293 (.L_HI(net2293));
 sg13g2_tiehi _26869__2294 (.L_HI(net2294));
 sg13g2_tiehi _26868__2295 (.L_HI(net2295));
 sg13g2_tiehi _26867__2296 (.L_HI(net2296));
 sg13g2_tiehi _26866__2297 (.L_HI(net2297));
 sg13g2_tiehi _26865__2298 (.L_HI(net2298));
 sg13g2_tiehi _26864__2299 (.L_HI(net2299));
 sg13g2_tiehi _26863__2300 (.L_HI(net2300));
 sg13g2_tiehi _26862__2301 (.L_HI(net2301));
 sg13g2_tiehi _26861__2302 (.L_HI(net2302));
 sg13g2_tiehi _26860__2303 (.L_HI(net2303));
 sg13g2_tiehi _26859__2304 (.L_HI(net2304));
 sg13g2_tiehi _26858__2305 (.L_HI(net2305));
 sg13g2_tiehi _26857__2306 (.L_HI(net2306));
 sg13g2_tiehi _26856__2307 (.L_HI(net2307));
 sg13g2_tiehi _26855__2308 (.L_HI(net2308));
 sg13g2_tiehi _26854__2309 (.L_HI(net2309));
 sg13g2_tiehi _26853__2310 (.L_HI(net2310));
 sg13g2_tiehi _26852__2311 (.L_HI(net2311));
 sg13g2_tiehi _26851__2312 (.L_HI(net2312));
 sg13g2_tiehi _26850__2313 (.L_HI(net2313));
 sg13g2_tiehi _26849__2314 (.L_HI(net2314));
 sg13g2_tiehi _26848__2315 (.L_HI(net2315));
 sg13g2_tiehi _26847__2316 (.L_HI(net2316));
 sg13g2_tiehi _26846__2317 (.L_HI(net2317));
 sg13g2_tiehi _26845__2318 (.L_HI(net2318));
 sg13g2_tiehi _26844__2319 (.L_HI(net2319));
 sg13g2_tiehi _26843__2320 (.L_HI(net2320));
 sg13g2_tiehi _26842__2321 (.L_HI(net2321));
 sg13g2_tiehi _26841__2322 (.L_HI(net2322));
 sg13g2_tiehi _26840__2323 (.L_HI(net2323));
 sg13g2_tiehi _26839__2324 (.L_HI(net2324));
 sg13g2_tiehi _26838__2325 (.L_HI(net2325));
 sg13g2_tiehi _26837__2326 (.L_HI(net2326));
 sg13g2_tiehi _26836__2327 (.L_HI(net2327));
 sg13g2_tiehi _26835__2328 (.L_HI(net2328));
 sg13g2_tiehi _26834__2329 (.L_HI(net2329));
 sg13g2_tiehi _26833__2330 (.L_HI(net2330));
 sg13g2_tiehi _26832__2331 (.L_HI(net2331));
 sg13g2_tiehi _26831__2332 (.L_HI(net2332));
 sg13g2_tiehi _26830__2333 (.L_HI(net2333));
 sg13g2_tiehi _26829__2334 (.L_HI(net2334));
 sg13g2_tiehi _26828__2335 (.L_HI(net2335));
 sg13g2_tiehi _26827__2336 (.L_HI(net2336));
 sg13g2_tiehi _26826__2337 (.L_HI(net2337));
 sg13g2_tiehi _26825__2338 (.L_HI(net2338));
 sg13g2_tiehi _26824__2339 (.L_HI(net2339));
 sg13g2_tiehi _26823__2340 (.L_HI(net2340));
 sg13g2_tiehi _26822__2341 (.L_HI(net2341));
 sg13g2_tiehi _26821__2342 (.L_HI(net2342));
 sg13g2_tiehi _26820__2343 (.L_HI(net2343));
 sg13g2_tiehi _26819__2344 (.L_HI(net2344));
 sg13g2_tiehi _26818__2345 (.L_HI(net2345));
 sg13g2_tiehi _26817__2346 (.L_HI(net2346));
 sg13g2_tiehi _26816__2347 (.L_HI(net2347));
 sg13g2_tiehi _26815__2348 (.L_HI(net2348));
 sg13g2_tiehi _26814__2349 (.L_HI(net2349));
 sg13g2_tiehi _26813__2350 (.L_HI(net2350));
 sg13g2_tiehi _26812__2351 (.L_HI(net2351));
 sg13g2_tiehi _26811__2352 (.L_HI(net2352));
 sg13g2_tiehi _26810__2353 (.L_HI(net2353));
 sg13g2_tiehi _26809__2354 (.L_HI(net2354));
 sg13g2_tiehi _26808__2355 (.L_HI(net2355));
 sg13g2_tiehi _26807__2356 (.L_HI(net2356));
 sg13g2_tiehi _26806__2357 (.L_HI(net2357));
 sg13g2_tiehi _26805__2358 (.L_HI(net2358));
 sg13g2_tiehi _26804__2359 (.L_HI(net2359));
 sg13g2_tiehi _28613__2360 (.L_HI(net2360));
 sg13g2_tiehi _28825__2361 (.L_HI(net2361));
 sg13g2_tiehi _28826__2362 (.L_HI(net2362));
 sg13g2_tiehi _28827__2363 (.L_HI(net2363));
 sg13g2_tiehi _26803__2364 (.L_HI(net2364));
 sg13g2_tiehi _26802__2365 (.L_HI(net2365));
 sg13g2_tiehi _26801__2366 (.L_HI(net2366));
 sg13g2_tiehi _26800__2367 (.L_HI(net2367));
 sg13g2_tiehi _26799__2368 (.L_HI(net2368));
 sg13g2_tiehi _26798__2369 (.L_HI(net2369));
 sg13g2_tiehi _26797__2370 (.L_HI(net2370));
 sg13g2_tiehi _26796__2371 (.L_HI(net2371));
 sg13g2_tiehi _26795__2372 (.L_HI(net2372));
 sg13g2_tiehi _26794__2373 (.L_HI(net2373));
 sg13g2_tiehi _26793__2374 (.L_HI(net2374));
 sg13g2_tiehi _26792__2375 (.L_HI(net2375));
 sg13g2_tiehi _26791__2376 (.L_HI(net2376));
 sg13g2_tiehi _26790__2377 (.L_HI(net2377));
 sg13g2_tiehi _26789__2378 (.L_HI(net2378));
 sg13g2_tiehi _26788__2379 (.L_HI(net2379));
 sg13g2_tiehi _26787__2380 (.L_HI(net2380));
 sg13g2_tiehi _26786__2381 (.L_HI(net2381));
 sg13g2_tiehi _26785__2382 (.L_HI(net2382));
 sg13g2_tiehi _26784__2383 (.L_HI(net2383));
 sg13g2_tiehi _26783__2384 (.L_HI(net2384));
 sg13g2_tiehi _26782__2385 (.L_HI(net2385));
 sg13g2_tiehi _26781__2386 (.L_HI(net2386));
 sg13g2_tiehi _26780__2387 (.L_HI(net2387));
 sg13g2_tiehi _26779__2388 (.L_HI(net2388));
 sg13g2_tiehi _26778__2389 (.L_HI(net2389));
 sg13g2_tiehi _26777__2390 (.L_HI(net2390));
 sg13g2_tiehi _26776__2391 (.L_HI(net2391));
 sg13g2_tiehi _26775__2392 (.L_HI(net2392));
 sg13g2_tiehi _26774__2393 (.L_HI(net2393));
 sg13g2_tiehi _26773__2394 (.L_HI(net2394));
 sg13g2_tiehi _26772__2395 (.L_HI(net2395));
 sg13g2_tiehi _26771__2396 (.L_HI(net2396));
 sg13g2_tiehi _26770__2397 (.L_HI(net2397));
 sg13g2_tiehi _26769__2398 (.L_HI(net2398));
 sg13g2_tiehi _26768__2399 (.L_HI(net2399));
 sg13g2_tiehi _26767__2400 (.L_HI(net2400));
 sg13g2_tiehi _26766__2401 (.L_HI(net2401));
 sg13g2_tiehi _26765__2402 (.L_HI(net2402));
 sg13g2_tiehi _26764__2403 (.L_HI(net2403));
 sg13g2_tiehi _26763__2404 (.L_HI(net2404));
 sg13g2_tiehi _26762__2405 (.L_HI(net2405));
 sg13g2_tiehi _26761__2406 (.L_HI(net2406));
 sg13g2_tiehi _26760__2407 (.L_HI(net2407));
 sg13g2_tiehi _26759__2408 (.L_HI(net2408));
 sg13g2_tiehi _26758__2409 (.L_HI(net2409));
 sg13g2_tiehi _26757__2410 (.L_HI(net2410));
 sg13g2_tiehi _26756__2411 (.L_HI(net2411));
 sg13g2_tiehi _28828__2412 (.L_HI(net2412));
 sg13g2_tiehi _28877__2413 (.L_HI(net2413));
 sg13g2_tiehi _28878__2414 (.L_HI(net2414));
 sg13g2_tiehi _28879__2415 (.L_HI(net2415));
 sg13g2_tiehi _28880__2416 (.L_HI(net2416));
 sg13g2_tiehi _28881__2417 (.L_HI(net2417));
 sg13g2_tiehi _28882__2418 (.L_HI(net2418));
 sg13g2_tiehi _28883__2419 (.L_HI(net2419));
 sg13g2_tiehi _26755__2420 (.L_HI(net2420));
 sg13g2_tiehi _26754__2421 (.L_HI(net2421));
 sg13g2_tiehi _26753__2422 (.L_HI(net2422));
 sg13g2_tiehi _26752__2423 (.L_HI(net2423));
 sg13g2_tiehi _26751__2424 (.L_HI(net2424));
 sg13g2_tiehi _26750__2425 (.L_HI(net2425));
 sg13g2_tiehi _26749__2426 (.L_HI(net2426));
 sg13g2_tiehi _26748__2427 (.L_HI(net2427));
 sg13g2_tiehi _26747__2428 (.L_HI(net2428));
 sg13g2_tiehi _26746__2429 (.L_HI(net2429));
 sg13g2_tiehi _26745__2430 (.L_HI(net2430));
 sg13g2_tiehi _26744__2431 (.L_HI(net2431));
 sg13g2_tiehi _26743__2432 (.L_HI(net2432));
 sg13g2_tiehi _26742__2433 (.L_HI(net2433));
 sg13g2_tiehi _26741__2434 (.L_HI(net2434));
 sg13g2_tiehi _26740__2435 (.L_HI(net2435));
 sg13g2_tiehi _26739__2436 (.L_HI(net2436));
 sg13g2_tiehi _26738__2437 (.L_HI(net2437));
 sg13g2_tiehi _26737__2438 (.L_HI(net2438));
 sg13g2_tiehi _26736__2439 (.L_HI(net2439));
 sg13g2_tiehi _26735__2440 (.L_HI(net2440));
 sg13g2_tiehi _26734__2441 (.L_HI(net2441));
 sg13g2_tiehi _26733__2442 (.L_HI(net2442));
 sg13g2_tiehi _28884__2443 (.L_HI(net2443));
 sg13g2_tiehi _26732__2444 (.L_HI(net2444));
 sg13g2_tiehi _26731__2445 (.L_HI(net2445));
 sg13g2_tiehi _26730__2446 (.L_HI(net2446));
 sg13g2_tiehi _26729__2447 (.L_HI(net2447));
 sg13g2_tiehi _26728__2448 (.L_HI(net2448));
 sg13g2_tiehi _26727__2449 (.L_HI(net2449));
 sg13g2_tiehi _26726__2450 (.L_HI(net2450));
 sg13g2_tiehi _26725__2451 (.L_HI(net2451));
 sg13g2_tiehi _26724__2452 (.L_HI(net2452));
 sg13g2_tiehi _26723__2453 (.L_HI(net2453));
 sg13g2_tiehi _26722__2454 (.L_HI(net2454));
 sg13g2_tiehi _26721__2455 (.L_HI(net2455));
 sg13g2_tiehi _26720__2456 (.L_HI(net2456));
 sg13g2_tiehi _26719__2457 (.L_HI(net2457));
 sg13g2_tiehi _26718__2458 (.L_HI(net2458));
 sg13g2_tiehi _26717__2459 (.L_HI(net2459));
 sg13g2_tiehi _26716__2460 (.L_HI(net2460));
 sg13g2_tiehi _26715__2461 (.L_HI(net2461));
 sg13g2_tiehi _26714__2462 (.L_HI(net2462));
 sg13g2_tiehi _26713__2463 (.L_HI(net2463));
 sg13g2_tiehi _26712__2464 (.L_HI(net2464));
 sg13g2_tiehi _26711__2465 (.L_HI(net2465));
 sg13g2_tiehi _26710__2466 (.L_HI(net2466));
 sg13g2_tiehi _26709__2467 (.L_HI(net2467));
 sg13g2_tiehi _26708__2468 (.L_HI(net2468));
 sg13g2_tiehi _26707__2469 (.L_HI(net2469));
 sg13g2_tiehi _26706__2470 (.L_HI(net2470));
 sg13g2_tiehi _26705__2471 (.L_HI(net2471));
 sg13g2_tiehi _26704__2472 (.L_HI(net2472));
 sg13g2_tiehi _26703__2473 (.L_HI(net2473));
 sg13g2_tiehi _26702__2474 (.L_HI(net2474));
 sg13g2_tiehi _26701__2475 (.L_HI(net2475));
 sg13g2_tiehi _26700__2476 (.L_HI(net2476));
 sg13g2_tiehi _26699__2477 (.L_HI(net2477));
 sg13g2_tiehi _26698__2478 (.L_HI(net2478));
 sg13g2_tiehi _26697__2479 (.L_HI(net2479));
 sg13g2_tiehi _26696__2480 (.L_HI(net2480));
 sg13g2_tiehi _26695__2481 (.L_HI(net2481));
 sg13g2_tiehi _26694__2482 (.L_HI(net2482));
 sg13g2_tiehi _26693__2483 (.L_HI(net2483));
 sg13g2_tiehi _26692__2484 (.L_HI(net2484));
 sg13g2_tiehi _26691__2485 (.L_HI(net2485));
 sg13g2_tiehi _26690__2486 (.L_HI(net2486));
 sg13g2_tiehi _26689__2487 (.L_HI(net2487));
 sg13g2_tiehi _26688__2488 (.L_HI(net2488));
 sg13g2_tiehi _26687__2489 (.L_HI(net2489));
 sg13g2_tiehi _26686__2490 (.L_HI(net2490));
 sg13g2_tiehi _26685__2491 (.L_HI(net2491));
 sg13g2_tiehi _26684__2492 (.L_HI(net2492));
 sg13g2_tiehi _26683__2493 (.L_HI(net2493));
 sg13g2_tiehi _26682__2494 (.L_HI(net2494));
 sg13g2_tiehi _26681__2495 (.L_HI(net2495));
 sg13g2_tiehi _26680__2496 (.L_HI(net2496));
 sg13g2_tiehi _26679__2497 (.L_HI(net2497));
 sg13g2_tiehi _26678__2498 (.L_HI(net2498));
 sg13g2_tiehi _26677__2499 (.L_HI(net2499));
 sg13g2_tiehi _26676__2500 (.L_HI(net2500));
 sg13g2_tiehi _26675__2501 (.L_HI(net2501));
 sg13g2_tiehi _26674__2502 (.L_HI(net2502));
 sg13g2_tiehi _26673__2503 (.L_HI(net2503));
 sg13g2_tiehi _26672__2504 (.L_HI(net2504));
 sg13g2_tiehi _26671__2505 (.L_HI(net2505));
 sg13g2_tiehi _26670__2506 (.L_HI(net2506));
 sg13g2_tiehi _26669__2507 (.L_HI(net2507));
 sg13g2_tiehi _26668__2508 (.L_HI(net2508));
 sg13g2_tiehi _26667__2509 (.L_HI(net2509));
 sg13g2_tiehi _28908__2510 (.L_HI(net2510));
 sg13g2_tiehi _26666__2511 (.L_HI(net2511));
 sg13g2_tiehi _26665__2512 (.L_HI(net2512));
 sg13g2_tiehi _26664__2513 (.L_HI(net2513));
 sg13g2_tiehi _26663__2514 (.L_HI(net2514));
 sg13g2_tiehi _26662__2515 (.L_HI(net2515));
 sg13g2_tiehi _26661__2516 (.L_HI(net2516));
 sg13g2_tiehi _26660__2517 (.L_HI(net2517));
 sg13g2_tiehi _26659__2518 (.L_HI(net2518));
 sg13g2_tiehi _29017__2519 (.L_HI(net2519));
 sg13g2_tiehi _26658__2520 (.L_HI(net2520));
 sg13g2_tiehi _26657__2521 (.L_HI(net2521));
 sg13g2_tiehi _26656__2522 (.L_HI(net2522));
 sg13g2_tiehi _26655__2523 (.L_HI(net2523));
 sg13g2_tiehi _26654__2524 (.L_HI(net2524));
 sg13g2_tiehi _26653__2525 (.L_HI(net2525));
 sg13g2_tiehi _26652__2526 (.L_HI(net2526));
 sg13g2_tiehi _26651__2527 (.L_HI(net2527));
 sg13g2_tiehi _26650__2528 (.L_HI(net2528));
 sg13g2_tiehi _26649__2529 (.L_HI(net2529));
 sg13g2_tiehi _26648__2530 (.L_HI(net2530));
 sg13g2_tiehi _26647__2531 (.L_HI(net2531));
 sg13g2_tiehi _26646__2532 (.L_HI(net2532));
 sg13g2_tiehi _26645__2533 (.L_HI(net2533));
 sg13g2_tiehi _26644__2534 (.L_HI(net2534));
 sg13g2_tiehi _26643__2535 (.L_HI(net2535));
 sg13g2_tiehi _26642__2536 (.L_HI(net2536));
 sg13g2_tiehi _26641__2537 (.L_HI(net2537));
 sg13g2_tiehi _26640__2538 (.L_HI(net2538));
 sg13g2_tiehi _26639__2539 (.L_HI(net2539));
 sg13g2_tiehi _26638__2540 (.L_HI(net2540));
 sg13g2_tiehi _26637__2541 (.L_HI(net2541));
 sg13g2_tiehi _26636__2542 (.L_HI(net2542));
 sg13g2_tiehi _26635__2543 (.L_HI(net2543));
 sg13g2_tiehi _26634__2544 (.L_HI(net2544));
 sg13g2_tiehi _26633__2545 (.L_HI(net2545));
 sg13g2_tiehi _26632__2546 (.L_HI(net2546));
 sg13g2_tiehi _26631__2547 (.L_HI(net2547));
 sg13g2_tiehi _26630__2548 (.L_HI(net2548));
 sg13g2_tiehi _26629__2549 (.L_HI(net2549));
 sg13g2_tiehi _26628__2550 (.L_HI(net2550));
 sg13g2_tiehi _26627__2551 (.L_HI(net2551));
 sg13g2_tiehi _26626__2552 (.L_HI(net2552));
 sg13g2_tiehi _26625__2553 (.L_HI(net2553));
 sg13g2_tiehi _26624__2554 (.L_HI(net2554));
 sg13g2_tiehi _26623__2555 (.L_HI(net2555));
 sg13g2_tiehi _26622__2556 (.L_HI(net2556));
 sg13g2_tiehi _26621__2557 (.L_HI(net2557));
 sg13g2_tiehi _26620__2558 (.L_HI(net2558));
 sg13g2_tiehi _26619__2559 (.L_HI(net2559));
 sg13g2_tiehi _26618__2560 (.L_HI(net2560));
 sg13g2_tiehi _26617__2561 (.L_HI(net2561));
 sg13g2_tiehi _26616__2562 (.L_HI(net2562));
 sg13g2_tiehi _26615__2563 (.L_HI(net2563));
 sg13g2_tiehi _26614__2564 (.L_HI(net2564));
 sg13g2_tiehi _26613__2565 (.L_HI(net2565));
 sg13g2_tiehi _26612__2566 (.L_HI(net2566));
 sg13g2_tiehi _26611__2567 (.L_HI(net2567));
 sg13g2_tiehi _26610__2568 (.L_HI(net2568));
 sg13g2_tiehi _26609__2569 (.L_HI(net2569));
 sg13g2_tiehi _26608__2570 (.L_HI(net2570));
 sg13g2_tiehi _26607__2571 (.L_HI(net2571));
 sg13g2_tiehi _26606__2572 (.L_HI(net2572));
 sg13g2_tiehi _26605__2573 (.L_HI(net2573));
 sg13g2_tiehi _26604__2574 (.L_HI(net2574));
 sg13g2_tiehi _26603__2575 (.L_HI(net2575));
 sg13g2_tiehi _26602__2576 (.L_HI(net2576));
 sg13g2_tiehi _26601__2577 (.L_HI(net2577));
 sg13g2_tiehi _26600__2578 (.L_HI(net2578));
 sg13g2_tiehi _26599__2579 (.L_HI(net2579));
 sg13g2_tiehi _26598__2580 (.L_HI(net2580));
 sg13g2_tiehi _26597__2581 (.L_HI(net2581));
 sg13g2_tiehi _26596__2582 (.L_HI(net2582));
 sg13g2_tiehi _26595__2583 (.L_HI(net2583));
 sg13g2_tiehi _26594__2584 (.L_HI(net2584));
 sg13g2_tiehi _26593__2585 (.L_HI(net2585));
 sg13g2_tiehi _26592__2586 (.L_HI(net2586));
 sg13g2_tiehi _26591__2587 (.L_HI(net2587));
 sg13g2_tiehi _26590__2588 (.L_HI(net2588));
 sg13g2_tiehi _26589__2589 (.L_HI(net2589));
 sg13g2_tiehi _29087__2590 (.L_HI(net2590));
 sg13g2_tiehi _26588__2591 (.L_HI(net2591));
 sg13g2_tiehi _29086__2592 (.L_HI(net2592));
 sg13g2_tiehi _26587__2593 (.L_HI(net2593));
 sg13g2_tiehi _29085__2594 (.L_HI(net2594));
 sg13g2_tiehi _26586__2595 (.L_HI(net2595));
 sg13g2_tiehi _29084__2596 (.L_HI(net2596));
 sg13g2_tiehi _26585__2597 (.L_HI(net2597));
 sg13g2_tiehi _29083__2598 (.L_HI(net2598));
 sg13g2_tiehi _26584__2599 (.L_HI(net2599));
 sg13g2_tiehi _29082__2600 (.L_HI(net2600));
 sg13g2_tiehi _26583__2601 (.L_HI(net2601));
 sg13g2_tiehi _29081__2602 (.L_HI(net2602));
 sg13g2_tiehi _26582__2603 (.L_HI(net2603));
 sg13g2_tiehi _26581__2604 (.L_HI(net2604));
 sg13g2_tiehi _26580__2605 (.L_HI(net2605));
 sg13g2_tiehi _26579__2606 (.L_HI(net2606));
 sg13g2_tiehi _26578__2607 (.L_HI(net2607));
 sg13g2_tiehi _26577__2608 (.L_HI(net2608));
 sg13g2_tiehi _26576__2609 (.L_HI(net2609));
 sg13g2_tiehi _26575__2610 (.L_HI(net2610));
 sg13g2_tiehi _26574__2611 (.L_HI(net2611));
 sg13g2_tiehi _26573__2612 (.L_HI(net2612));
 sg13g2_tiehi _26572__2613 (.L_HI(net2613));
 sg13g2_tiehi _26571__2614 (.L_HI(net2614));
 sg13g2_tiehi _26570__2615 (.L_HI(net2615));
 sg13g2_tiehi _26569__2616 (.L_HI(net2616));
 sg13g2_tiehi _26568__2617 (.L_HI(net2617));
 sg13g2_tiehi _26567__2618 (.L_HI(net2618));
 sg13g2_tiehi _26566__2619 (.L_HI(net2619));
 sg13g2_tiehi _26565__2620 (.L_HI(net2620));
 sg13g2_tiehi _26564__2621 (.L_HI(net2621));
 sg13g2_tiehi _26563__2622 (.L_HI(net2622));
 sg13g2_tiehi _26562__2623 (.L_HI(net2623));
 sg13g2_tiehi _26561__2624 (.L_HI(net2624));
 sg13g2_tiehi _26560__2625 (.L_HI(net2625));
 sg13g2_tiehi _26559__2626 (.L_HI(net2626));
 sg13g2_tiehi _26558__2627 (.L_HI(net2627));
 sg13g2_tiehi _26557__2628 (.L_HI(net2628));
 sg13g2_tiehi _26556__2629 (.L_HI(net2629));
 sg13g2_tiehi _26555__2630 (.L_HI(net2630));
 sg13g2_tiehi _26554__2631 (.L_HI(net2631));
 sg13g2_tiehi _26553__2632 (.L_HI(net2632));
 sg13g2_tiehi _26552__2633 (.L_HI(net2633));
 sg13g2_tiehi _26551__2634 (.L_HI(net2634));
 sg13g2_tiehi _26550__2635 (.L_HI(net2635));
 sg13g2_tiehi _29080__2636 (.L_HI(net2636));
 sg13g2_tiehi _29079__2637 (.L_HI(net2637));
 sg13g2_tiehi _29078__2638 (.L_HI(net2638));
 sg13g2_tiehi _29077__2639 (.L_HI(net2639));
 sg13g2_tiehi _29076__2640 (.L_HI(net2640));
 sg13g2_tiehi _29075__2641 (.L_HI(net2641));
 sg13g2_tiehi _29074__2642 (.L_HI(net2642));
 sg13g2_tiehi _29073__2643 (.L_HI(net2643));
 sg13g2_tiehi _29072__2644 (.L_HI(net2644));
 sg13g2_tiehi _29071__2645 (.L_HI(net2645));
 sg13g2_tiehi _29070__2646 (.L_HI(net2646));
 sg13g2_tiehi _29069__2647 (.L_HI(net2647));
 sg13g2_tiehi _29068__2648 (.L_HI(net2648));
 sg13g2_tiehi _29067__2649 (.L_HI(net2649));
 sg13g2_tiehi _29066__2650 (.L_HI(net2650));
 sg13g2_tiehi _29065__2651 (.L_HI(net2651));
 sg13g2_tiehi _29064__2652 (.L_HI(net2652));
 sg13g2_tiehi _29063__2653 (.L_HI(net2653));
 sg13g2_tiehi _29062__2654 (.L_HI(net2654));
 sg13g2_tiehi _29061__2655 (.L_HI(net2655));
 sg13g2_tiehi _29060__2656 (.L_HI(net2656));
 sg13g2_tiehi _29059__2657 (.L_HI(net2657));
 sg13g2_tiehi _29058__2658 (.L_HI(net2658));
 sg13g2_tiehi _29057__2659 (.L_HI(net2659));
 sg13g2_tiehi _29056__2660 (.L_HI(net2660));
 sg13g2_tiehi _29055__2661 (.L_HI(net2661));
 sg13g2_tiehi _29054__2662 (.L_HI(net2662));
 sg13g2_tiehi _29053__2663 (.L_HI(net2663));
 sg13g2_tiehi _29052__2664 (.L_HI(net2664));
 sg13g2_tiehi _29051__2665 (.L_HI(net2665));
 sg13g2_tiehi _29050__2666 (.L_HI(net2666));
 sg13g2_tiehi _29049__2667 (.L_HI(net2667));
 sg13g2_tiehi _29048__2668 (.L_HI(net2668));
 sg13g2_tiehi _29047__2669 (.L_HI(net2669));
 sg13g2_tiehi _29046__2670 (.L_HI(net2670));
 sg13g2_tiehi _29045__2671 (.L_HI(net2671));
 sg13g2_tiehi _29044__2672 (.L_HI(net2672));
 sg13g2_tiehi _29043__2673 (.L_HI(net2673));
 sg13g2_tiehi _29042__2674 (.L_HI(net2674));
 sg13g2_tiehi _29041__2675 (.L_HI(net2675));
 sg13g2_tiehi _29040__2676 (.L_HI(net2676));
 sg13g2_tiehi _29039__2677 (.L_HI(net2677));
 sg13g2_tiehi _29038__2678 (.L_HI(net2678));
 sg13g2_tiehi _29037__2679 (.L_HI(net2679));
 sg13g2_tiehi _29036__2680 (.L_HI(net2680));
 sg13g2_tiehi _29035__2681 (.L_HI(net2681));
 sg13g2_tiehi _29034__2682 (.L_HI(net2682));
 sg13g2_tiehi _29033__2683 (.L_HI(net2683));
 sg13g2_tiehi _29032__2684 (.L_HI(net2684));
 sg13g2_tiehi _29031__2685 (.L_HI(net2685));
 sg13g2_tiehi _29030__2686 (.L_HI(net2686));
 sg13g2_tiehi _29417__2687 (.L_HI(net2687));
 sg13g2_tiehi _29029__2688 (.L_HI(net2688));
 sg13g2_tiehi _29416__2689 (.L_HI(net2689));
 sg13g2_tiehi _29027__2690 (.L_HI(net2690));
 sg13g2_tiehi _29415__2691 (.L_HI(net2691));
 sg13g2_tiehi _29026__2692 (.L_HI(net2692));
 sg13g2_tiehi _29414__2693 (.L_HI(net2693));
 sg13g2_tiehi _29025__2694 (.L_HI(net2694));
 sg13g2_tiehi _29413__2695 (.L_HI(net2695));
 sg13g2_tiehi _29024__2696 (.L_HI(net2696));
 sg13g2_tiehi _29412__2697 (.L_HI(net2697));
 sg13g2_tiehi _29023__2698 (.L_HI(net2698));
 sg13g2_tiehi _29411__2699 (.L_HI(net2699));
 sg13g2_tiehi _29022__2700 (.L_HI(net2700));
 sg13g2_tiehi _29410__2701 (.L_HI(net2701));
 sg13g2_tiehi _29021__2702 (.L_HI(net2702));
 sg13g2_tiehi _29409__2703 (.L_HI(net2703));
 sg13g2_tiehi _29020__2704 (.L_HI(net2704));
 sg13g2_tiehi _29408__2705 (.L_HI(net2705));
 sg13g2_tiehi _29019__2706 (.L_HI(net2706));
 sg13g2_tiehi _29018__2707 (.L_HI(net2707));
 sg13g2_tiehi _29016__2708 (.L_HI(net2708));
 sg13g2_tiehi _29015__2709 (.L_HI(net2709));
 sg13g2_tiehi _29014__2710 (.L_HI(net2710));
 sg13g2_tiehi _29013__2711 (.L_HI(net2711));
 sg13g2_tiehi _29012__2712 (.L_HI(net2712));
 sg13g2_tiehi _29011__2713 (.L_HI(net2713));
 sg13g2_tiehi _29010__2714 (.L_HI(net2714));
 sg13g2_tiehi _29009__2715 (.L_HI(net2715));
 sg13g2_tiehi _29008__2716 (.L_HI(net2716));
 sg13g2_tiehi _29007__2717 (.L_HI(net2717));
 sg13g2_tiehi _29006__2718 (.L_HI(net2718));
 sg13g2_tiehi _29005__2719 (.L_HI(net2719));
 sg13g2_tiehi _29004__2720 (.L_HI(net2720));
 sg13g2_tiehi _29003__2721 (.L_HI(net2721));
 sg13g2_tiehi _29002__2722 (.L_HI(net2722));
 sg13g2_tiehi _29407__2723 (.L_HI(net2723));
 sg13g2_tiehi _29001__2724 (.L_HI(net2724));
 sg13g2_tiehi _29406__2725 (.L_HI(net2725));
 sg13g2_tiehi _29000__2726 (.L_HI(net2726));
 sg13g2_tiehi _29405__2727 (.L_HI(net2727));
 sg13g2_tiehi _28999__2728 (.L_HI(net2728));
 sg13g2_tiehi _29404__2729 (.L_HI(net2729));
 sg13g2_tiehi _28998__2730 (.L_HI(net2730));
 sg13g2_tiehi _29403__2731 (.L_HI(net2731));
 sg13g2_tiehi _28997__2732 (.L_HI(net2732));
 sg13g2_tiehi _29402__2733 (.L_HI(net2733));
 sg13g2_tiehi _28996__2734 (.L_HI(net2734));
 sg13g2_tiehi _29401__2735 (.L_HI(net2735));
 sg13g2_tiehi _28995__2736 (.L_HI(net2736));
 sg13g2_tiehi _29400__2737 (.L_HI(net2737));
 sg13g2_tiehi _28994__2738 (.L_HI(net2738));
 sg13g2_tiehi _29399__2739 (.L_HI(net2739));
 sg13g2_tiehi _28993__2740 (.L_HI(net2740));
 sg13g2_tiehi _28992__2741 (.L_HI(net2741));
 sg13g2_tiehi _28991__2742 (.L_HI(net2742));
 sg13g2_tiehi _28990__2743 (.L_HI(net2743));
 sg13g2_tiehi _28989__2744 (.L_HI(net2744));
 sg13g2_tiehi _28988__2745 (.L_HI(net2745));
 sg13g2_tiehi _28987__2746 (.L_HI(net2746));
 sg13g2_tiehi _28986__2747 (.L_HI(net2747));
 sg13g2_tiehi _28985__2748 (.L_HI(net2748));
 sg13g2_tiehi _28984__2749 (.L_HI(net2749));
 sg13g2_tiehi _28983__2750 (.L_HI(net2750));
 sg13g2_tiehi _28982__2751 (.L_HI(net2751));
 sg13g2_tiehi _28981__2752 (.L_HI(net2752));
 sg13g2_tiehi _28980__2753 (.L_HI(net2753));
 sg13g2_tiehi _28979__2754 (.L_HI(net2754));
 sg13g2_tiehi _28978__2755 (.L_HI(net2755));
 sg13g2_tiehi _28977__2756 (.L_HI(net2756));
 sg13g2_tiehi _28976__2757 (.L_HI(net2757));
 sg13g2_tiehi _28975__2758 (.L_HI(net2758));
 sg13g2_tiehi _28974__2759 (.L_HI(net2759));
 sg13g2_tiehi _28973__2760 (.L_HI(net2760));
 sg13g2_tiehi _28972__2761 (.L_HI(net2761));
 sg13g2_tiehi _28971__2762 (.L_HI(net2762));
 sg13g2_tiehi _28970__2763 (.L_HI(net2763));
 sg13g2_tiehi _28969__2764 (.L_HI(net2764));
 sg13g2_tiehi _28968__2765 (.L_HI(net2765));
 sg13g2_tiehi _28967__2766 (.L_HI(net2766));
 sg13g2_tiehi _28966__2767 (.L_HI(net2767));
 sg13g2_tiehi _28965__2768 (.L_HI(net2768));
 sg13g2_tiehi _28964__2769 (.L_HI(net2769));
 sg13g2_tiehi _28963__2770 (.L_HI(net2770));
 sg13g2_tiehi _28962__2771 (.L_HI(net2771));
 sg13g2_tiehi _28961__2772 (.L_HI(net2772));
 sg13g2_tiehi _28960__2773 (.L_HI(net2773));
 sg13g2_tiehi _28959__2774 (.L_HI(net2774));
 sg13g2_tiehi _28958__2775 (.L_HI(net2775));
 sg13g2_tiehi _28957__2776 (.L_HI(net2776));
 sg13g2_tiehi _28956__2777 (.L_HI(net2777));
 sg13g2_tiehi _28955__2778 (.L_HI(net2778));
 sg13g2_tiehi _28954__2779 (.L_HI(net2779));
 sg13g2_tiehi _28953__2780 (.L_HI(net2780));
 sg13g2_tiehi _28952__2781 (.L_HI(net2781));
 sg13g2_tiehi _28951__2782 (.L_HI(net2782));
 sg13g2_tiehi _28950__2783 (.L_HI(net2783));
 sg13g2_tiehi _28949__2784 (.L_HI(net2784));
 sg13g2_tiehi _28948__2785 (.L_HI(net2785));
 sg13g2_tiehi _28947__2786 (.L_HI(net2786));
 sg13g2_tiehi _28946__2787 (.L_HI(net2787));
 sg13g2_tiehi _28945__2788 (.L_HI(net2788));
 sg13g2_tiehi _28944__2789 (.L_HI(net2789));
 sg13g2_tiehi _28943__2790 (.L_HI(net2790));
 sg13g2_tiehi _28942__2791 (.L_HI(net2791));
 sg13g2_tiehi _28941__2792 (.L_HI(net2792));
 sg13g2_tiehi _28940__2793 (.L_HI(net2793));
 sg13g2_tiehi _28939__2794 (.L_HI(net2794));
 sg13g2_tiehi _28938__2795 (.L_HI(net2795));
 sg13g2_tiehi _28937__2796 (.L_HI(net2796));
 sg13g2_tiehi _28936__2797 (.L_HI(net2797));
 sg13g2_tiehi _28935__2798 (.L_HI(net2798));
 sg13g2_tiehi _28934__2799 (.L_HI(net2799));
 sg13g2_tiehi _28933__2800 (.L_HI(net2800));
 sg13g2_tiehi _28932__2801 (.L_HI(net2801));
 sg13g2_tiehi _28931__2802 (.L_HI(net2802));
 sg13g2_tiehi _28930__2803 (.L_HI(net2803));
 sg13g2_tiehi _28929__2804 (.L_HI(net2804));
 sg13g2_tiehi _28928__2805 (.L_HI(net2805));
 sg13g2_tiehi _28927__2806 (.L_HI(net2806));
 sg13g2_tiehi _28926__2807 (.L_HI(net2807));
 sg13g2_tiehi _28925__2808 (.L_HI(net2808));
 sg13g2_tiehi _28924__2809 (.L_HI(net2809));
 sg13g2_tiehi _28923__2810 (.L_HI(net2810));
 sg13g2_tiehi _28922__2811 (.L_HI(net2811));
 sg13g2_tiehi _28921__2812 (.L_HI(net2812));
 sg13g2_tiehi _28920__2813 (.L_HI(net2813));
 sg13g2_tiehi _28919__2814 (.L_HI(net2814));
 sg13g2_tiehi _28918__2815 (.L_HI(net2815));
 sg13g2_tiehi _28917__2816 (.L_HI(net2816));
 sg13g2_tiehi _28916__2817 (.L_HI(net2817));
 sg13g2_tiehi _28915__2818 (.L_HI(net2818));
 sg13g2_tiehi _28914__2819 (.L_HI(net2819));
 sg13g2_tiehi _28913__2820 (.L_HI(net2820));
 sg13g2_tiehi _28912__2821 (.L_HI(net2821));
 sg13g2_tiehi _28911__2822 (.L_HI(net2822));
 sg13g2_tiehi _28910__2823 (.L_HI(net2823));
 sg13g2_tiehi _28909__2824 (.L_HI(net2824));
 sg13g2_tiehi _28907__2825 (.L_HI(net2825));
 sg13g2_tiehi _28906__2826 (.L_HI(net2826));
 sg13g2_tiehi _28905__2827 (.L_HI(net2827));
 sg13g2_tiehi _28904__2828 (.L_HI(net2828));
 sg13g2_tiehi _28903__2829 (.L_HI(net2829));
 sg13g2_tiehi _28902__2830 (.L_HI(net2830));
 sg13g2_tiehi _28901__2831 (.L_HI(net2831));
 sg13g2_tiehi _28900__2832 (.L_HI(net2832));
 sg13g2_tiehi _28899__2833 (.L_HI(net2833));
 sg13g2_tiehi _28898__2834 (.L_HI(net2834));
 sg13g2_tiehi _29398__2835 (.L_HI(net2835));
 sg13g2_tiehi _28897__2836 (.L_HI(net2836));
 sg13g2_tiehi _29397__2837 (.L_HI(net2837));
 sg13g2_tiehi _28896__2838 (.L_HI(net2838));
 sg13g2_tiehi _28895__2839 (.L_HI(net2839));
 sg13g2_tiehi _28894__2840 (.L_HI(net2840));
 sg13g2_tiehi _28893__2841 (.L_HI(net2841));
 sg13g2_tiehi _28892__2842 (.L_HI(net2842));
 sg13g2_tiehi _28891__2843 (.L_HI(net2843));
 sg13g2_tiehi _28890__2844 (.L_HI(net2844));
 sg13g2_tiehi _28889__2845 (.L_HI(net2845));
 sg13g2_tiehi _28888__2846 (.L_HI(net2846));
 sg13g2_tiehi _29396__2847 (.L_HI(net2847));
 sg13g2_tiehi _28887__2848 (.L_HI(net2848));
 sg13g2_tiehi _28886__2849 (.L_HI(net2849));
 sg13g2_tiehi _28885__2850 (.L_HI(net2850));
 sg13g2_tiehi _28876__2851 (.L_HI(net2851));
 sg13g2_tiehi _28875__2852 (.L_HI(net2852));
 sg13g2_tiehi _28874__2853 (.L_HI(net2853));
 sg13g2_tiehi _28873__2854 (.L_HI(net2854));
 sg13g2_tiehi _28872__2855 (.L_HI(net2855));
 sg13g2_tiehi _28871__2856 (.L_HI(net2856));
 sg13g2_tiehi _28870__2857 (.L_HI(net2857));
 sg13g2_tiehi _29395__2858 (.L_HI(net2858));
 sg13g2_tiehi _28869__2859 (.L_HI(net2859));
 sg13g2_tiehi _28868__2860 (.L_HI(net2860));
 sg13g2_tiehi _28867__2861 (.L_HI(net2861));
 sg13g2_tiehi _28866__2862 (.L_HI(net2862));
 sg13g2_tiehi _28865__2863 (.L_HI(net2863));
 sg13g2_tiehi _28864__2864 (.L_HI(net2864));
 sg13g2_tiehi _28863__2865 (.L_HI(net2865));
 sg13g2_tiehi _28862__2866 (.L_HI(net2866));
 sg13g2_tiehi _29394__2867 (.L_HI(net2867));
 sg13g2_tiehi _28861__2868 (.L_HI(net2868));
 sg13g2_tiehi _28860__2869 (.L_HI(net2869));
 sg13g2_tiehi _28859__2870 (.L_HI(net2870));
 sg13g2_tiehi _28858__2871 (.L_HI(net2871));
 sg13g2_tiehi _28857__2872 (.L_HI(net2872));
 sg13g2_tiehi _28856__2873 (.L_HI(net2873));
 sg13g2_tiehi _28855__2874 (.L_HI(net2874));
 sg13g2_tiehi _28854__2875 (.L_HI(net2875));
 sg13g2_tiehi _28853__2876 (.L_HI(net2876));
 sg13g2_tiehi _28852__2877 (.L_HI(net2877));
 sg13g2_tiehi _28851__2878 (.L_HI(net2878));
 sg13g2_tiehi _28850__2879 (.L_HI(net2879));
 sg13g2_tiehi _28849__2880 (.L_HI(net2880));
 sg13g2_tiehi _28848__2881 (.L_HI(net2881));
 sg13g2_tiehi _28847__2882 (.L_HI(net2882));
 sg13g2_tiehi _28846__2883 (.L_HI(net2883));
 sg13g2_tiehi _28845__2884 (.L_HI(net2884));
 sg13g2_tiehi _28844__2885 (.L_HI(net2885));
 sg13g2_tiehi tt_um_rejunity_atari2600_2886 (.L_HI(net2886));
 sg13g2_tiehi tt_um_rejunity_atari2600_2887 (.L_HI(net2887));
 sg13g2_tiehi tt_um_rejunity_atari2600_2888 (.L_HI(net2888));
 sg13g2_tiehi tt_um_rejunity_atari2600_2889 (.L_HI(net2889));
 sg13g2_tiehi tt_um_rejunity_atari2600_2890 (.L_HI(net2890));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _32308_ (.A(uio_oe[5]),
    .X(uio_oe[2]));
 sg13g2_buf_1 _32309_ (.A(uio_oe[5]),
    .X(uio_oe[4]));
 sg13g2_buf_1 _32310_ (.A(net5537),
    .X(uio_out[0]));
 sg13g2_buf_1 _32311_ (.A(\flash_rom.spi_clk_out ),
    .X(uio_out[3]));
 sg13g2_buf_2 _32312_ (.A(audio_pwm),
    .X(uio_out[7]));
 sg13g2_buf_1 _32313_ (.A(\hvsync_gen.vga.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_2 _32314_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout4543 (.A(net4544),
    .X(net4543));
 sg13g2_buf_2 fanout4544 (.A(_07066_),
    .X(net4544));
 sg13g2_buf_2 fanout4545 (.A(net4546),
    .X(net4545));
 sg13g2_buf_2 fanout4546 (.A(_07066_),
    .X(net4546));
 sg13g2_buf_2 fanout4547 (.A(net4549),
    .X(net4547));
 sg13g2_buf_2 fanout4548 (.A(net4549),
    .X(net4548));
 sg13g2_buf_2 fanout4549 (.A(_07017_),
    .X(net4549));
 sg13g2_buf_2 fanout4550 (.A(net4551),
    .X(net4550));
 sg13g2_buf_2 fanout4551 (.A(_07014_),
    .X(net4551));
 sg13g2_buf_4 fanout4552 (.X(net4552),
    .A(_05892_));
 sg13g2_buf_2 fanout4553 (.A(_05892_),
    .X(net4553));
 sg13g2_buf_2 fanout4554 (.A(_06341_),
    .X(net4554));
 sg13g2_buf_2 fanout4555 (.A(_06341_),
    .X(net4555));
 sg13g2_buf_2 fanout4556 (.A(net4557),
    .X(net4556));
 sg13g2_buf_2 fanout4557 (.A(_03237_),
    .X(net4557));
 sg13g2_buf_2 fanout4558 (.A(net4560),
    .X(net4558));
 sg13g2_buf_1 fanout4559 (.A(net4560),
    .X(net4559));
 sg13g2_buf_1 fanout4560 (.A(net4563),
    .X(net4560));
 sg13g2_buf_2 fanout4561 (.A(net4563),
    .X(net4561));
 sg13g2_buf_1 fanout4562 (.A(net4563),
    .X(net4562));
 sg13g2_buf_2 fanout4563 (.A(_03236_),
    .X(net4563));
 sg13g2_buf_2 fanout4564 (.A(net4566),
    .X(net4564));
 sg13g2_buf_1 fanout4565 (.A(net4566),
    .X(net4565));
 sg13g2_buf_2 fanout4566 (.A(net4569),
    .X(net4566));
 sg13g2_buf_2 fanout4567 (.A(net4569),
    .X(net4567));
 sg13g2_buf_2 fanout4568 (.A(net4569),
    .X(net4568));
 sg13g2_buf_2 fanout4569 (.A(_10446_),
    .X(net4569));
 sg13g2_buf_2 fanout4570 (.A(_10446_),
    .X(net4570));
 sg13g2_buf_1 fanout4571 (.A(_10446_),
    .X(net4571));
 sg13g2_buf_2 fanout4572 (.A(_07638_),
    .X(net4572));
 sg13g2_buf_2 fanout4573 (.A(_07840_),
    .X(net4573));
 sg13g2_buf_2 fanout4574 (.A(_07840_),
    .X(net4574));
 sg13g2_buf_4 fanout4575 (.X(net4575),
    .A(_07763_));
 sg13g2_buf_4 fanout4576 (.X(net4576),
    .A(_07709_));
 sg13g2_buf_4 fanout4577 (.X(net4577),
    .A(_07671_));
 sg13g2_buf_2 fanout4578 (.A(_05353_),
    .X(net4578));
 sg13g2_buf_2 fanout4579 (.A(_05353_),
    .X(net4579));
 sg13g2_buf_2 fanout4580 (.A(_05352_),
    .X(net4580));
 sg13g2_buf_1 fanout4581 (.A(_05352_),
    .X(net4581));
 sg13g2_buf_2 fanout4582 (.A(net4584),
    .X(net4582));
 sg13g2_buf_2 fanout4583 (.A(net4584),
    .X(net4583));
 sg13g2_buf_4 fanout4584 (.X(net4584),
    .A(_09986_));
 sg13g2_buf_4 fanout4585 (.X(net4585),
    .A(_07858_));
 sg13g2_buf_4 fanout4586 (.X(net4586),
    .A(_07856_));
 sg13g2_buf_2 fanout4587 (.A(net4588),
    .X(net4587));
 sg13g2_buf_2 fanout4588 (.A(_07848_),
    .X(net4588));
 sg13g2_buf_4 fanout4589 (.X(net4589),
    .A(_07838_));
 sg13g2_buf_4 fanout4590 (.X(net4590),
    .A(_07836_));
 sg13g2_buf_4 fanout4591 (.X(net4591),
    .A(_07783_));
 sg13g2_buf_4 fanout4592 (.X(net4592),
    .A(_07781_));
 sg13g2_buf_2 fanout4593 (.A(net4594),
    .X(net4593));
 sg13g2_buf_2 fanout4594 (.A(_07773_),
    .X(net4594));
 sg13g2_buf_2 fanout4595 (.A(net4596),
    .X(net4595));
 sg13g2_buf_2 fanout4596 (.A(_07765_),
    .X(net4596));
 sg13g2_buf_4 fanout4597 (.X(net4597),
    .A(_07761_));
 sg13g2_buf_4 fanout4598 (.X(net4598),
    .A(_07759_));
 sg13g2_buf_2 fanout4599 (.A(_07751_),
    .X(net4599));
 sg13g2_buf_2 fanout4600 (.A(_07751_),
    .X(net4600));
 sg13g2_buf_2 fanout4601 (.A(net4602),
    .X(net4601));
 sg13g2_buf_2 fanout4602 (.A(_07743_),
    .X(net4602));
 sg13g2_buf_4 fanout4603 (.X(net4603),
    .A(_07741_));
 sg13g2_buf_4 fanout4604 (.X(net4604),
    .A(_07739_));
 sg13g2_buf_4 fanout4605 (.X(net4605),
    .A(_07737_));
 sg13g2_buf_2 fanout4606 (.A(_07729_),
    .X(net4606));
 sg13g2_buf_2 fanout4607 (.A(_07729_),
    .X(net4607));
 sg13g2_buf_4 fanout4608 (.X(net4608),
    .A(_07727_));
 sg13g2_buf_4 fanout4609 (.X(net4609),
    .A(_07725_));
 sg13g2_buf_4 fanout4610 (.X(net4610),
    .A(_07723_));
 sg13g2_buf_2 fanout4611 (.A(_07715_),
    .X(net4611));
 sg13g2_buf_2 fanout4612 (.A(_07715_),
    .X(net4612));
 sg13g2_buf_4 fanout4613 (.X(net4613),
    .A(_07713_));
 sg13g2_buf_4 fanout4614 (.X(net4614),
    .A(_07711_));
 sg13g2_buf_2 fanout4615 (.A(_07701_),
    .X(net4615));
 sg13g2_buf_2 fanout4616 (.A(_07701_),
    .X(net4616));
 sg13g2_buf_4 fanout4617 (.X(net4617),
    .A(_07699_));
 sg13g2_buf_4 fanout4618 (.X(net4618),
    .A(_07697_));
 sg13g2_buf_4 fanout4619 (.X(net4619),
    .A(_07695_));
 sg13g2_buf_2 fanout4620 (.A(_07687_),
    .X(net4620));
 sg13g2_buf_2 fanout4621 (.A(_07687_),
    .X(net4621));
 sg13g2_buf_4 fanout4622 (.X(net4622),
    .A(_07685_));
 sg13g2_buf_4 fanout4623 (.X(net4623),
    .A(_07683_));
 sg13g2_buf_4 fanout4624 (.X(net4624),
    .A(_07681_));
 sg13g2_buf_2 fanout4625 (.A(_07673_),
    .X(net4625));
 sg13g2_buf_2 fanout4626 (.A(_07673_),
    .X(net4626));
 sg13g2_buf_4 fanout4627 (.X(net4627),
    .A(_07668_));
 sg13g2_buf_4 fanout4628 (.X(net4628),
    .A(_07666_));
 sg13g2_buf_4 fanout4629 (.X(net4629),
    .A(_07664_));
 sg13g2_buf_2 fanout4630 (.A(net4631),
    .X(net4630));
 sg13g2_buf_2 fanout4631 (.A(_07655_),
    .X(net4631));
 sg13g2_buf_2 fanout4632 (.A(net4633),
    .X(net4632));
 sg13g2_buf_2 fanout4633 (.A(_07646_),
    .X(net4633));
 sg13g2_buf_2 fanout4634 (.A(net4635),
    .X(net4634));
 sg13g2_buf_2 fanout4635 (.A(_07604_),
    .X(net4635));
 sg13g2_buf_2 fanout4636 (.A(_07595_),
    .X(net4636));
 sg13g2_buf_2 fanout4637 (.A(_07595_),
    .X(net4637));
 sg13g2_buf_2 fanout4638 (.A(_07579_),
    .X(net4638));
 sg13g2_buf_2 fanout4639 (.A(_07579_),
    .X(net4639));
 sg13g2_buf_2 fanout4640 (.A(_07570_),
    .X(net4640));
 sg13g2_buf_2 fanout4641 (.A(_07570_),
    .X(net4641));
 sg13g2_buf_2 fanout4642 (.A(net4643),
    .X(net4642));
 sg13g2_buf_2 fanout4643 (.A(_07559_),
    .X(net4643));
 sg13g2_buf_2 fanout4644 (.A(net4645),
    .X(net4644));
 sg13g2_buf_2 fanout4645 (.A(_07219_),
    .X(net4645));
 sg13g2_buf_2 fanout4646 (.A(net4647),
    .X(net4646));
 sg13g2_buf_2 fanout4647 (.A(_07133_),
    .X(net4647));
 sg13g2_buf_2 fanout4648 (.A(_07117_),
    .X(net4648));
 sg13g2_buf_2 fanout4649 (.A(_07117_),
    .X(net4649));
 sg13g2_buf_2 fanout4650 (.A(_07106_),
    .X(net4650));
 sg13g2_buf_2 fanout4651 (.A(_07106_),
    .X(net4651));
 sg13g2_buf_2 fanout4652 (.A(net4653),
    .X(net4652));
 sg13g2_buf_2 fanout4653 (.A(_06929_),
    .X(net4653));
 sg13g2_buf_2 fanout4654 (.A(net4655),
    .X(net4654));
 sg13g2_buf_2 fanout4655 (.A(_06883_),
    .X(net4655));
 sg13g2_buf_2 fanout4656 (.A(_06811_),
    .X(net4656));
 sg13g2_buf_2 fanout4657 (.A(_06811_),
    .X(net4657));
 sg13g2_buf_2 fanout4658 (.A(_06735_),
    .X(net4658));
 sg13g2_buf_1 fanout4659 (.A(_06735_),
    .X(net4659));
 sg13g2_buf_2 fanout4660 (.A(net4661),
    .X(net4660));
 sg13g2_buf_2 fanout4661 (.A(_06688_),
    .X(net4661));
 sg13g2_buf_4 fanout4662 (.X(net4662),
    .A(_06620_));
 sg13g2_buf_4 fanout4663 (.X(net4663),
    .A(_06611_));
 sg13g2_buf_2 fanout4664 (.A(_06456_),
    .X(net4664));
 sg13g2_buf_2 fanout4665 (.A(_06456_),
    .X(net4665));
 sg13g2_buf_2 fanout4666 (.A(net4667),
    .X(net4666));
 sg13g2_buf_2 fanout4667 (.A(_06422_),
    .X(net4667));
 sg13g2_buf_2 fanout4668 (.A(_05480_),
    .X(net4668));
 sg13g2_buf_2 fanout4669 (.A(_05480_),
    .X(net4669));
 sg13g2_buf_2 fanout4670 (.A(net4671),
    .X(net4670));
 sg13g2_buf_2 fanout4671 (.A(_05400_),
    .X(net4671));
 sg13g2_buf_2 fanout4672 (.A(_05381_),
    .X(net4672));
 sg13g2_buf_2 fanout4673 (.A(_05381_),
    .X(net4673));
 sg13g2_buf_2 fanout4674 (.A(_05256_),
    .X(net4674));
 sg13g2_buf_2 fanout4675 (.A(_05109_),
    .X(net4675));
 sg13g2_buf_2 fanout4676 (.A(_05109_),
    .X(net4676));
 sg13g2_buf_2 fanout4677 (.A(net4678),
    .X(net4677));
 sg13g2_buf_2 fanout4678 (.A(_05099_),
    .X(net4678));
 sg13g2_buf_2 fanout4679 (.A(_05087_),
    .X(net4679));
 sg13g2_buf_2 fanout4680 (.A(_05087_),
    .X(net4680));
 sg13g2_buf_2 fanout4681 (.A(net4682),
    .X(net4681));
 sg13g2_buf_2 fanout4682 (.A(_05078_),
    .X(net4682));
 sg13g2_buf_2 fanout4683 (.A(_05017_),
    .X(net4683));
 sg13g2_buf_2 fanout4684 (.A(_05017_),
    .X(net4684));
 sg13g2_buf_2 fanout4685 (.A(net4686),
    .X(net4685));
 sg13g2_buf_2 fanout4686 (.A(_05004_),
    .X(net4686));
 sg13g2_buf_2 fanout4687 (.A(_04992_),
    .X(net4687));
 sg13g2_buf_2 fanout4688 (.A(_04992_),
    .X(net4688));
 sg13g2_buf_2 fanout4689 (.A(_04979_),
    .X(net4689));
 sg13g2_buf_2 fanout4690 (.A(_04979_),
    .X(net4690));
 sg13g2_buf_2 fanout4691 (.A(_04970_),
    .X(net4691));
 sg13g2_buf_2 fanout4692 (.A(_04970_),
    .X(net4692));
 sg13g2_buf_2 fanout4693 (.A(_04959_),
    .X(net4693));
 sg13g2_buf_2 fanout4694 (.A(_04959_),
    .X(net4694));
 sg13g2_buf_2 fanout4695 (.A(net4696),
    .X(net4695));
 sg13g2_buf_2 fanout4696 (.A(_04946_),
    .X(net4696));
 sg13g2_buf_2 fanout4697 (.A(net4698),
    .X(net4697));
 sg13g2_buf_2 fanout4698 (.A(_04934_),
    .X(net4698));
 sg13g2_buf_2 fanout4699 (.A(_04922_),
    .X(net4699));
 sg13g2_buf_2 fanout4700 (.A(_04922_),
    .X(net4700));
 sg13g2_buf_2 fanout4701 (.A(net4702),
    .X(net4701));
 sg13g2_buf_2 fanout4702 (.A(_04913_),
    .X(net4702));
 sg13g2_buf_2 fanout4703 (.A(net4704),
    .X(net4703));
 sg13g2_buf_2 fanout4704 (.A(_04904_),
    .X(net4704));
 sg13g2_buf_2 fanout4705 (.A(net4706),
    .X(net4705));
 sg13g2_buf_2 fanout4706 (.A(_04894_),
    .X(net4706));
 sg13g2_buf_2 fanout4707 (.A(_04848_),
    .X(net4707));
 sg13g2_buf_2 fanout4708 (.A(_04848_),
    .X(net4708));
 sg13g2_buf_2 fanout4709 (.A(net4710),
    .X(net4709));
 sg13g2_buf_2 fanout4710 (.A(_04837_),
    .X(net4710));
 sg13g2_buf_2 fanout4711 (.A(_04828_),
    .X(net4711));
 sg13g2_buf_2 fanout4712 (.A(_04828_),
    .X(net4712));
 sg13g2_buf_2 fanout4713 (.A(net4714),
    .X(net4713));
 sg13g2_buf_2 fanout4714 (.A(_04818_),
    .X(net4714));
 sg13g2_buf_2 fanout4715 (.A(_04802_),
    .X(net4715));
 sg13g2_buf_2 fanout4716 (.A(_04802_),
    .X(net4716));
 sg13g2_buf_2 fanout4717 (.A(_03091_),
    .X(net4717));
 sg13g2_buf_2 fanout4718 (.A(_03091_),
    .X(net4718));
 sg13g2_buf_2 fanout4719 (.A(_03062_),
    .X(net4719));
 sg13g2_buf_2 fanout4720 (.A(_03062_),
    .X(net4720));
 sg13g2_buf_2 fanout4721 (.A(_03050_),
    .X(net4721));
 sg13g2_buf_2 fanout4722 (.A(_03050_),
    .X(net4722));
 sg13g2_buf_4 fanout4723 (.X(net4723),
    .A(net4724));
 sg13g2_buf_4 fanout4724 (.X(net4724),
    .A(_08633_));
 sg13g2_buf_2 fanout4725 (.A(_06994_),
    .X(net4725));
 sg13g2_buf_4 fanout4726 (.X(net4726),
    .A(_06623_));
 sg13g2_buf_2 fanout4727 (.A(net4728),
    .X(net4727));
 sg13g2_buf_2 fanout4728 (.A(_06495_),
    .X(net4728));
 sg13g2_buf_2 fanout4729 (.A(_06433_),
    .X(net4729));
 sg13g2_buf_4 fanout4730 (.X(net4730),
    .A(_05449_));
 sg13g2_buf_2 fanout4731 (.A(_05398_),
    .X(net4731));
 sg13g2_buf_2 fanout4732 (.A(_05249_),
    .X(net4732));
 sg13g2_buf_8 fanout4733 (.A(_04816_),
    .X(net4733));
 sg13g2_buf_4 fanout4734 (.X(net4734),
    .A(_04816_));
 sg13g2_buf_8 fanout4735 (.A(_03167_),
    .X(net4735));
 sg13g2_buf_4 fanout4736 (.X(net4736),
    .A(_03167_));
 sg13g2_buf_8 fanout4737 (.A(_03159_),
    .X(net4737));
 sg13g2_buf_8 fanout4738 (.A(_03159_),
    .X(net4738));
 sg13g2_buf_8 fanout4739 (.A(_03090_),
    .X(net4739));
 sg13g2_buf_8 fanout4740 (.A(_03090_),
    .X(net4740));
 sg13g2_buf_8 fanout4741 (.A(_03061_),
    .X(net4741));
 sg13g2_buf_8 fanout4742 (.A(_03061_),
    .X(net4742));
 sg13g2_buf_8 fanout4743 (.A(_03049_),
    .X(net4743));
 sg13g2_buf_8 fanout4744 (.A(_03049_),
    .X(net4744));
 sg13g2_buf_8 fanout4745 (.A(_03044_),
    .X(net4745));
 sg13g2_buf_8 fanout4746 (.A(_03044_),
    .X(net4746));
 sg13g2_buf_8 fanout4747 (.A(net4748),
    .X(net4747));
 sg13g2_buf_8 fanout4748 (.A(_03009_),
    .X(net4748));
 sg13g2_buf_4 fanout4749 (.X(net4749),
    .A(_10257_));
 sg13g2_buf_1 fanout4750 (.A(_10257_),
    .X(net4750));
 sg13g2_buf_4 fanout4751 (.X(net4751),
    .A(_08632_));
 sg13g2_buf_2 fanout4752 (.A(_06809_),
    .X(net4752));
 sg13g2_buf_2 fanout4753 (.A(_06738_),
    .X(net4753));
 sg13g2_buf_2 fanout4754 (.A(_06616_),
    .X(net4754));
 sg13g2_buf_2 fanout4755 (.A(_06616_),
    .X(net4755));
 sg13g2_buf_4 fanout4756 (.X(net4756),
    .A(net4759));
 sg13g2_buf_2 fanout4757 (.A(net4759),
    .X(net4757));
 sg13g2_buf_2 fanout4758 (.A(net4759),
    .X(net4758));
 sg13g2_buf_2 fanout4759 (.A(_06616_),
    .X(net4759));
 sg13g2_buf_2 fanout4760 (.A(net4761),
    .X(net4760));
 sg13g2_buf_1 fanout4761 (.A(net4762),
    .X(net4761));
 sg13g2_buf_2 fanout4762 (.A(_05248_),
    .X(net4762));
 sg13g2_buf_4 fanout4763 (.X(net4763),
    .A(_03158_));
 sg13g2_buf_2 fanout4764 (.A(_10180_),
    .X(net4764));
 sg13g2_buf_1 fanout4765 (.A(net4766),
    .X(net4765));
 sg13g2_buf_4 fanout4766 (.X(net4766),
    .A(_10180_));
 sg13g2_buf_2 fanout4767 (.A(net4768),
    .X(net4767));
 sg13g2_buf_4 fanout4768 (.X(net4768),
    .A(_10051_));
 sg13g2_buf_2 fanout4769 (.A(net4770),
    .X(net4769));
 sg13g2_buf_2 fanout4770 (.A(_09820_),
    .X(net4770));
 sg13g2_buf_4 fanout4771 (.X(net4771),
    .A(net4772));
 sg13g2_buf_4 fanout4772 (.X(net4772),
    .A(_08783_));
 sg13g2_buf_2 fanout4773 (.A(net4774),
    .X(net4773));
 sg13g2_buf_4 fanout4774 (.X(net4774),
    .A(net4775));
 sg13g2_buf_8 fanout4775 (.A(_08754_),
    .X(net4775));
 sg13g2_buf_4 fanout4776 (.X(net4776),
    .A(_08729_));
 sg13g2_buf_2 fanout4777 (.A(net4780),
    .X(net4777));
 sg13g2_buf_4 fanout4778 (.X(net4778),
    .A(net4780));
 sg13g2_buf_1 fanout4779 (.A(net4780),
    .X(net4779));
 sg13g2_buf_4 fanout4780 (.X(net4780),
    .A(_08630_));
 sg13g2_buf_2 fanout4781 (.A(_10424_),
    .X(net4781));
 sg13g2_buf_2 fanout4782 (.A(net4784),
    .X(net4782));
 sg13g2_buf_1 fanout4783 (.A(net4784),
    .X(net4783));
 sg13g2_buf_2 fanout4784 (.A(_10115_),
    .X(net4784));
 sg13g2_buf_4 fanout4785 (.X(net4785),
    .A(net4788));
 sg13g2_buf_2 fanout4786 (.A(net4788),
    .X(net4786));
 sg13g2_buf_4 fanout4787 (.X(net4787),
    .A(net4788));
 sg13g2_buf_2 fanout4788 (.A(net4797),
    .X(net4788));
 sg13g2_buf_4 fanout4789 (.X(net4789),
    .A(net4797));
 sg13g2_buf_4 fanout4790 (.X(net4790),
    .A(net4797));
 sg13g2_buf_4 fanout4791 (.X(net4791),
    .A(net4793));
 sg13g2_buf_4 fanout4792 (.X(net4792),
    .A(net4793));
 sg13g2_buf_4 fanout4793 (.X(net4793),
    .A(net4796));
 sg13g2_buf_4 fanout4794 (.X(net4794),
    .A(net4796));
 sg13g2_buf_4 fanout4795 (.X(net4795),
    .A(net4796));
 sg13g2_buf_2 fanout4796 (.A(net4797),
    .X(net4796));
 sg13g2_buf_2 fanout4797 (.A(_08734_),
    .X(net4797));
 sg13g2_buf_4 fanout4798 (.X(net4798),
    .A(net4800));
 sg13g2_buf_4 fanout4799 (.X(net4799),
    .A(net4800));
 sg13g2_buf_4 fanout4800 (.X(net4800),
    .A(net4807));
 sg13g2_buf_4 fanout4801 (.X(net4801),
    .A(net4806));
 sg13g2_buf_4 fanout4802 (.X(net4802),
    .A(net4805));
 sg13g2_buf_4 fanout4803 (.X(net4803),
    .A(net4805));
 sg13g2_buf_2 fanout4804 (.A(net4805),
    .X(net4804));
 sg13g2_buf_2 fanout4805 (.A(net4806),
    .X(net4805));
 sg13g2_buf_2 fanout4806 (.A(net4807),
    .X(net4806));
 sg13g2_buf_2 fanout4807 (.A(_08734_),
    .X(net4807));
 sg13g2_buf_4 fanout4808 (.X(net4808),
    .A(net4810));
 sg13g2_buf_4 fanout4809 (.X(net4809),
    .A(net4810));
 sg13g2_buf_2 fanout4810 (.A(net4817),
    .X(net4810));
 sg13g2_buf_4 fanout4811 (.X(net4811),
    .A(net4812));
 sg13g2_buf_4 fanout4812 (.X(net4812),
    .A(net4817));
 sg13g2_buf_4 fanout4813 (.X(net4813),
    .A(net4815));
 sg13g2_buf_2 fanout4814 (.A(net4815),
    .X(net4814));
 sg13g2_buf_2 fanout4815 (.A(net4817),
    .X(net4815));
 sg13g2_buf_4 fanout4816 (.X(net4816),
    .A(net4817));
 sg13g2_buf_4 fanout4817 (.X(net4817),
    .A(net4829));
 sg13g2_buf_4 fanout4818 (.X(net4818),
    .A(net4824));
 sg13g2_buf_2 fanout4819 (.A(net4824),
    .X(net4819));
 sg13g2_buf_4 fanout4820 (.X(net4820),
    .A(net4821));
 sg13g2_buf_4 fanout4821 (.X(net4821),
    .A(net4824));
 sg13g2_buf_4 fanout4822 (.X(net4822),
    .A(net4823));
 sg13g2_buf_4 fanout4823 (.X(net4823),
    .A(net4824));
 sg13g2_buf_2 fanout4824 (.A(net4829),
    .X(net4824));
 sg13g2_buf_4 fanout4825 (.X(net4825),
    .A(net4826));
 sg13g2_buf_2 fanout4826 (.A(net4829),
    .X(net4826));
 sg13g2_buf_4 fanout4827 (.X(net4827),
    .A(net4828));
 sg13g2_buf_2 fanout4828 (.A(net4829),
    .X(net4828));
 sg13g2_buf_4 fanout4829 (.X(net4829),
    .A(_08734_));
 sg13g2_buf_4 fanout4830 (.X(net4830),
    .A(net4833));
 sg13g2_buf_2 fanout4831 (.A(net4833),
    .X(net4831));
 sg13g2_buf_4 fanout4832 (.X(net4832),
    .A(net4833));
 sg13g2_buf_2 fanout4833 (.A(net4836),
    .X(net4833));
 sg13g2_buf_4 fanout4834 (.X(net4834),
    .A(net4835));
 sg13g2_buf_4 fanout4835 (.X(net4835),
    .A(net4836));
 sg13g2_buf_2 fanout4836 (.A(net4852),
    .X(net4836));
 sg13g2_buf_4 fanout4837 (.X(net4837),
    .A(net4839));
 sg13g2_buf_4 fanout4838 (.X(net4838),
    .A(net4839));
 sg13g2_buf_2 fanout4839 (.A(net4842),
    .X(net4839));
 sg13g2_buf_4 fanout4840 (.X(net4840),
    .A(net4841));
 sg13g2_buf_4 fanout4841 (.X(net4841),
    .A(net4842));
 sg13g2_buf_2 fanout4842 (.A(net4852),
    .X(net4842));
 sg13g2_buf_4 fanout4843 (.X(net4843),
    .A(net4845));
 sg13g2_buf_4 fanout4844 (.X(net4844),
    .A(net4845));
 sg13g2_buf_4 fanout4845 (.X(net4845),
    .A(net4852));
 sg13g2_buf_4 fanout4846 (.X(net4846),
    .A(net4847));
 sg13g2_buf_4 fanout4847 (.X(net4847),
    .A(net4851));
 sg13g2_buf_4 fanout4848 (.X(net4848),
    .A(net4850));
 sg13g2_buf_2 fanout4849 (.A(net4850),
    .X(net4849));
 sg13g2_buf_4 fanout4850 (.X(net4850),
    .A(net4851));
 sg13g2_buf_4 fanout4851 (.X(net4851),
    .A(net4852));
 sg13g2_buf_4 fanout4852 (.X(net4852),
    .A(net4875));
 sg13g2_buf_4 fanout4853 (.X(net4853),
    .A(net4855));
 sg13g2_buf_4 fanout4854 (.X(net4854),
    .A(net4855));
 sg13g2_buf_2 fanout4855 (.A(net4858),
    .X(net4855));
 sg13g2_buf_4 fanout4856 (.X(net4856),
    .A(net4858));
 sg13g2_buf_4 fanout4857 (.X(net4857),
    .A(net4858));
 sg13g2_buf_2 fanout4858 (.A(net4875),
    .X(net4858));
 sg13g2_buf_4 fanout4859 (.X(net4859),
    .A(net4860));
 sg13g2_buf_4 fanout4860 (.X(net4860),
    .A(net4862));
 sg13g2_buf_4 fanout4861 (.X(net4861),
    .A(net4862));
 sg13g2_buf_4 fanout4862 (.X(net4862),
    .A(net4875));
 sg13g2_buf_4 fanout4863 (.X(net4863),
    .A(net4866));
 sg13g2_buf_2 fanout4864 (.A(net4866),
    .X(net4864));
 sg13g2_buf_4 fanout4865 (.X(net4865),
    .A(net4866));
 sg13g2_buf_2 fanout4866 (.A(net4874),
    .X(net4866));
 sg13g2_buf_4 fanout4867 (.X(net4867),
    .A(net4874));
 sg13g2_buf_2 fanout4868 (.A(net4874),
    .X(net4868));
 sg13g2_buf_4 fanout4869 (.X(net4869),
    .A(net4874));
 sg13g2_buf_2 fanout4870 (.A(net4874),
    .X(net4870));
 sg13g2_buf_4 fanout4871 (.X(net4871),
    .A(net4873));
 sg13g2_buf_2 fanout4872 (.A(net4873),
    .X(net4872));
 sg13g2_buf_2 fanout4873 (.A(net4874),
    .X(net4873));
 sg13g2_buf_4 fanout4874 (.X(net4874),
    .A(net4875));
 sg13g2_buf_4 fanout4875 (.X(net4875),
    .A(_08731_));
 sg13g2_buf_4 fanout4876 (.X(net4876),
    .A(net4877));
 sg13g2_buf_4 fanout4877 (.X(net4877),
    .A(net4879));
 sg13g2_buf_4 fanout4878 (.X(net4878),
    .A(net4879));
 sg13g2_buf_4 fanout4879 (.X(net4879),
    .A(_08617_));
 sg13g2_buf_4 fanout4880 (.X(net4880),
    .A(net4882));
 sg13g2_buf_2 fanout4881 (.A(net4882),
    .X(net4881));
 sg13g2_buf_4 fanout4882 (.X(net4882),
    .A(net4891));
 sg13g2_buf_4 fanout4883 (.X(net4883),
    .A(net4891));
 sg13g2_buf_2 fanout4884 (.A(net4891),
    .X(net4884));
 sg13g2_buf_4 fanout4885 (.X(net4885),
    .A(net4887));
 sg13g2_buf_2 fanout4886 (.A(net4887),
    .X(net4886));
 sg13g2_buf_2 fanout4887 (.A(net4890),
    .X(net4887));
 sg13g2_buf_2 fanout4888 (.A(net4890),
    .X(net4888));
 sg13g2_buf_4 fanout4889 (.X(net4889),
    .A(net4890));
 sg13g2_buf_2 fanout4890 (.A(net4891),
    .X(net4890));
 sg13g2_buf_4 fanout4891 (.X(net4891),
    .A(_08564_));
 sg13g2_buf_4 fanout4892 (.X(net4892),
    .A(net4894));
 sg13g2_buf_2 fanout4893 (.A(net4895),
    .X(net4893));
 sg13g2_buf_1 fanout4894 (.A(net4895),
    .X(net4894));
 sg13g2_buf_4 fanout4895 (.X(net4895),
    .A(net4901));
 sg13g2_buf_4 fanout4896 (.X(net4896),
    .A(net4900));
 sg13g2_buf_2 fanout4897 (.A(net4899),
    .X(net4897));
 sg13g2_buf_2 fanout4898 (.A(net4899),
    .X(net4898));
 sg13g2_buf_2 fanout4899 (.A(net4900),
    .X(net4899));
 sg13g2_buf_2 fanout4900 (.A(net4901),
    .X(net4900));
 sg13g2_buf_2 fanout4901 (.A(_08564_),
    .X(net4901));
 sg13g2_buf_4 fanout4902 (.X(net4902),
    .A(net4904));
 sg13g2_buf_4 fanout4903 (.X(net4903),
    .A(net4904));
 sg13g2_buf_2 fanout4904 (.A(net4912),
    .X(net4904));
 sg13g2_buf_4 fanout4905 (.X(net4905),
    .A(net4907));
 sg13g2_buf_2 fanout4906 (.A(net4907),
    .X(net4906));
 sg13g2_buf_4 fanout4907 (.X(net4907),
    .A(net4912));
 sg13g2_buf_4 fanout4908 (.X(net4908),
    .A(net4909));
 sg13g2_buf_2 fanout4909 (.A(net4912),
    .X(net4909));
 sg13g2_buf_4 fanout4910 (.X(net4910),
    .A(net4911));
 sg13g2_buf_2 fanout4911 (.A(net4912),
    .X(net4911));
 sg13g2_buf_2 fanout4912 (.A(net4924),
    .X(net4912));
 sg13g2_buf_2 fanout4913 (.A(net4919),
    .X(net4913));
 sg13g2_buf_2 fanout4914 (.A(net4919),
    .X(net4914));
 sg13g2_buf_4 fanout4915 (.X(net4915),
    .A(net4916));
 sg13g2_buf_4 fanout4916 (.X(net4916),
    .A(net4919));
 sg13g2_buf_2 fanout4917 (.A(net4918),
    .X(net4917));
 sg13g2_buf_2 fanout4918 (.A(net4919),
    .X(net4918));
 sg13g2_buf_2 fanout4919 (.A(net4924),
    .X(net4919));
 sg13g2_buf_2 fanout4920 (.A(net4921),
    .X(net4920));
 sg13g2_buf_2 fanout4921 (.A(net4924),
    .X(net4921));
 sg13g2_buf_4 fanout4922 (.X(net4922),
    .A(net4923));
 sg13g2_buf_2 fanout4923 (.A(net4924),
    .X(net4923));
 sg13g2_buf_4 fanout4924 (.X(net4924),
    .A(_08564_));
 sg13g2_buf_2 fanout4925 (.A(net4926),
    .X(net4925));
 sg13g2_buf_4 fanout4926 (.X(net4926),
    .A(net4936));
 sg13g2_buf_2 fanout4927 (.A(net4929),
    .X(net4927));
 sg13g2_buf_4 fanout4928 (.X(net4928),
    .A(net4929));
 sg13g2_buf_4 fanout4929 (.X(net4929),
    .A(net4936));
 sg13g2_buf_4 fanout4930 (.X(net4930),
    .A(net4931));
 sg13g2_buf_2 fanout4931 (.A(net4932),
    .X(net4931));
 sg13g2_buf_4 fanout4932 (.X(net4932),
    .A(net4935));
 sg13g2_buf_2 fanout4933 (.A(net4934),
    .X(net4933));
 sg13g2_buf_4 fanout4934 (.X(net4934),
    .A(net4935));
 sg13g2_buf_4 fanout4935 (.X(net4935),
    .A(net4936));
 sg13g2_buf_2 fanout4936 (.A(_08747_),
    .X(net4936));
 sg13g2_buf_4 fanout4937 (.X(net4937),
    .A(net4939));
 sg13g2_buf_4 fanout4938 (.X(net4938),
    .A(net4939));
 sg13g2_buf_4 fanout4939 (.X(net4939),
    .A(net4940));
 sg13g2_buf_4 fanout4940 (.X(net4940),
    .A(net4947));
 sg13g2_buf_4 fanout4941 (.X(net4941),
    .A(net4947));
 sg13g2_buf_4 fanout4942 (.X(net4942),
    .A(net4947));
 sg13g2_buf_4 fanout4943 (.X(net4943),
    .A(net4944));
 sg13g2_buf_4 fanout4944 (.X(net4944),
    .A(net4946));
 sg13g2_buf_4 fanout4945 (.X(net4945),
    .A(net4946));
 sg13g2_buf_4 fanout4946 (.X(net4946),
    .A(net4947));
 sg13g2_buf_2 fanout4947 (.A(_08742_),
    .X(net4947));
 sg13g2_buf_8 fanout4948 (.A(_08732_),
    .X(net4948));
 sg13g2_buf_4 fanout4949 (.X(net4949),
    .A(net4951));
 sg13g2_buf_4 fanout4950 (.X(net4950),
    .A(net4951));
 sg13g2_buf_4 fanout4951 (.X(net4951),
    .A(net4953));
 sg13g2_buf_4 fanout4952 (.X(net4952),
    .A(net4953));
 sg13g2_buf_4 fanout4953 (.X(net4953),
    .A(_08730_));
 sg13g2_buf_4 fanout4954 (.X(net4954),
    .A(net4955));
 sg13g2_buf_2 fanout4955 (.A(net4956),
    .X(net4955));
 sg13g2_buf_4 fanout4956 (.X(net4956),
    .A(_08730_));
 sg13g2_buf_4 fanout4957 (.X(net4957),
    .A(net4958));
 sg13g2_buf_4 fanout4958 (.X(net4958),
    .A(net4959));
 sg13g2_buf_4 fanout4959 (.X(net4959),
    .A(_08730_));
 sg13g2_buf_4 fanout4960 (.X(net4960),
    .A(net4963));
 sg13g2_buf_1 fanout4961 (.A(net4963),
    .X(net4961));
 sg13g2_buf_4 fanout4962 (.X(net4962),
    .A(net4963));
 sg13g2_buf_2 fanout4963 (.A(net4966),
    .X(net4963));
 sg13g2_buf_2 fanout4964 (.A(net4965),
    .X(net4964));
 sg13g2_buf_2 fanout4965 (.A(net4966),
    .X(net4965));
 sg13g2_buf_2 fanout4966 (.A(net4982),
    .X(net4966));
 sg13g2_buf_4 fanout4967 (.X(net4967),
    .A(net4969));
 sg13g2_buf_4 fanout4968 (.X(net4968),
    .A(net4969));
 sg13g2_buf_4 fanout4969 (.X(net4969),
    .A(net4982));
 sg13g2_buf_4 fanout4970 (.X(net4970),
    .A(net4972));
 sg13g2_buf_1 fanout4971 (.A(net4972),
    .X(net4971));
 sg13g2_buf_4 fanout4972 (.X(net4972),
    .A(net4982));
 sg13g2_buf_2 fanout4973 (.A(net4975),
    .X(net4973));
 sg13g2_buf_2 fanout4974 (.A(net4975),
    .X(net4974));
 sg13g2_buf_4 fanout4975 (.X(net4975),
    .A(net4982));
 sg13g2_buf_2 fanout4976 (.A(net4978),
    .X(net4976));
 sg13g2_buf_4 fanout4977 (.X(net4977),
    .A(net4978));
 sg13g2_buf_2 fanout4978 (.A(net4981),
    .X(net4978));
 sg13g2_buf_4 fanout4979 (.X(net4979),
    .A(net4980));
 sg13g2_buf_2 fanout4980 (.A(net4981),
    .X(net4980));
 sg13g2_buf_2 fanout4981 (.A(net4982),
    .X(net4981));
 sg13g2_buf_4 fanout4982 (.X(net4982),
    .A(net5005));
 sg13g2_buf_4 fanout4983 (.X(net4983),
    .A(net4985));
 sg13g2_buf_2 fanout4984 (.A(net4985),
    .X(net4984));
 sg13g2_buf_2 fanout4985 (.A(net4993),
    .X(net4985));
 sg13g2_buf_4 fanout4986 (.X(net4986),
    .A(net4987));
 sg13g2_buf_4 fanout4987 (.X(net4987),
    .A(net4993));
 sg13g2_buf_2 fanout4988 (.A(net4993),
    .X(net4988));
 sg13g2_buf_4 fanout4989 (.X(net4989),
    .A(net4990));
 sg13g2_buf_2 fanout4990 (.A(net4992),
    .X(net4990));
 sg13g2_buf_2 fanout4991 (.A(net4992),
    .X(net4991));
 sg13g2_buf_2 fanout4992 (.A(net4993),
    .X(net4992));
 sg13g2_buf_2 fanout4993 (.A(net5005),
    .X(net4993));
 sg13g2_buf_4 fanout4994 (.X(net4994),
    .A(net4996));
 sg13g2_buf_1 fanout4995 (.A(net4996),
    .X(net4995));
 sg13g2_buf_4 fanout4996 (.X(net4996),
    .A(net4999));
 sg13g2_buf_4 fanout4997 (.X(net4997),
    .A(net4998));
 sg13g2_buf_4 fanout4998 (.X(net4998),
    .A(net4999));
 sg13g2_buf_2 fanout4999 (.A(net5005),
    .X(net4999));
 sg13g2_buf_4 fanout5000 (.X(net5000),
    .A(net5001));
 sg13g2_buf_2 fanout5001 (.A(net5004),
    .X(net5001));
 sg13g2_buf_4 fanout5002 (.X(net5002),
    .A(net5004));
 sg13g2_buf_1 fanout5003 (.A(net5004),
    .X(net5003));
 sg13g2_buf_2 fanout5004 (.A(net5005),
    .X(net5004));
 sg13g2_buf_4 fanout5005 (.X(net5005),
    .A(_08675_));
 sg13g2_buf_4 fanout5006 (.X(net5006),
    .A(net5011));
 sg13g2_buf_2 fanout5007 (.A(net5010),
    .X(net5007));
 sg13g2_buf_4 fanout5008 (.X(net5008),
    .A(net5009));
 sg13g2_buf_4 fanout5009 (.X(net5009),
    .A(net5010));
 sg13g2_buf_4 fanout5010 (.X(net5010),
    .A(net5011));
 sg13g2_buf_4 fanout5011 (.X(net5011),
    .A(net5017));
 sg13g2_buf_4 fanout5012 (.X(net5012),
    .A(net5014));
 sg13g2_buf_2 fanout5013 (.A(net5014),
    .X(net5013));
 sg13g2_buf_2 fanout5014 (.A(net5017),
    .X(net5014));
 sg13g2_buf_4 fanout5015 (.X(net5015),
    .A(net5017));
 sg13g2_buf_4 fanout5016 (.X(net5016),
    .A(net5017));
 sg13g2_buf_4 fanout5017 (.X(net5017),
    .A(_08582_));
 sg13g2_buf_2 fanout5018 (.A(_06510_),
    .X(net5018));
 sg13g2_buf_2 fanout5019 (.A(_06510_),
    .X(net5019));
 sg13g2_buf_4 fanout5020 (.X(net5020),
    .A(net5021));
 sg13g2_buf_8 fanout5021 (.A(net5022),
    .X(net5021));
 sg13g2_buf_8 fanout5022 (.A(_08728_),
    .X(net5022));
 sg13g2_buf_2 fanout5023 (.A(net5024),
    .X(net5023));
 sg13g2_buf_8 fanout5024 (.A(_08727_),
    .X(net5024));
 sg13g2_buf_4 fanout5025 (.X(net5025),
    .A(net5026));
 sg13g2_buf_8 fanout5026 (.A(_08629_),
    .X(net5026));
 sg13g2_buf_8 fanout5027 (.A(_08628_),
    .X(net5027));
 sg13g2_buf_8 fanout5028 (.A(_08628_),
    .X(net5028));
 sg13g2_buf_4 fanout5029 (.X(net5029),
    .A(net5031));
 sg13g2_buf_2 fanout5030 (.A(net5031),
    .X(net5030));
 sg13g2_buf_8 fanout5031 (.A(_08578_),
    .X(net5031));
 sg13g2_buf_8 fanout5032 (.A(_08577_),
    .X(net5032));
 sg13g2_buf_4 fanout5033 (.X(net5033),
    .A(_08577_));
 sg13g2_buf_4 fanout5034 (.X(net5034),
    .A(_08562_));
 sg13g2_buf_4 fanout5035 (.X(net5035),
    .A(_08553_));
 sg13g2_buf_8 fanout5036 (.A(_08545_),
    .X(net5036));
 sg13g2_buf_8 fanout5037 (.A(net5039),
    .X(net5037));
 sg13g2_buf_2 fanout5038 (.A(net5039),
    .X(net5038));
 sg13g2_buf_8 fanout5039 (.A(_08544_),
    .X(net5039));
 sg13g2_buf_4 fanout5040 (.X(net5040),
    .A(net5042));
 sg13g2_buf_2 fanout5041 (.A(net5042),
    .X(net5041));
 sg13g2_buf_4 fanout5042 (.X(net5042),
    .A(net5048));
 sg13g2_buf_4 fanout5043 (.X(net5043),
    .A(net5048));
 sg13g2_buf_2 fanout5044 (.A(net5048),
    .X(net5044));
 sg13g2_buf_4 fanout5045 (.X(net5045),
    .A(net5047));
 sg13g2_buf_2 fanout5046 (.A(net5047),
    .X(net5046));
 sg13g2_buf_8 fanout5047 (.A(net5048),
    .X(net5047));
 sg13g2_buf_2 fanout5048 (.A(_03040_),
    .X(net5048));
 sg13g2_buf_4 fanout5049 (.X(net5049),
    .A(net5052));
 sg13g2_buf_4 fanout5050 (.X(net5050),
    .A(net5051));
 sg13g2_buf_4 fanout5051 (.X(net5051),
    .A(net5052));
 sg13g2_buf_2 fanout5052 (.A(_03040_),
    .X(net5052));
 sg13g2_buf_4 fanout5053 (.X(net5053),
    .A(net5054));
 sg13g2_buf_8 fanout5054 (.A(_03040_),
    .X(net5054));
 sg13g2_buf_8 fanout5055 (.A(net5058),
    .X(net5055));
 sg13g2_buf_8 fanout5056 (.A(net5058),
    .X(net5056));
 sg13g2_buf_4 fanout5057 (.X(net5057),
    .A(net5058));
 sg13g2_buf_8 fanout5058 (.A(_03039_),
    .X(net5058));
 sg13g2_buf_8 fanout5059 (.A(net5063),
    .X(net5059));
 sg13g2_buf_4 fanout5060 (.X(net5060),
    .A(net5061));
 sg13g2_buf_2 fanout5061 (.A(net5062),
    .X(net5061));
 sg13g2_buf_4 fanout5062 (.X(net5062),
    .A(net5063));
 sg13g2_buf_4 fanout5063 (.X(net5063),
    .A(_03039_));
 sg13g2_buf_4 fanout5064 (.X(net5064),
    .A(net5065));
 sg13g2_buf_4 fanout5065 (.X(net5065),
    .A(net5068));
 sg13g2_buf_4 fanout5066 (.X(net5066),
    .A(net5067));
 sg13g2_buf_4 fanout5067 (.X(net5067),
    .A(net5068));
 sg13g2_buf_4 fanout5068 (.X(net5068),
    .A(_03034_));
 sg13g2_buf_4 fanout5069 (.X(net5069),
    .A(net5070));
 sg13g2_buf_4 fanout5070 (.X(net5070),
    .A(net5071));
 sg13g2_buf_4 fanout5071 (.X(net5071),
    .A(_03034_));
 sg13g2_buf_4 fanout5072 (.X(net5072),
    .A(net5077));
 sg13g2_buf_4 fanout5073 (.X(net5073),
    .A(net5077));
 sg13g2_buf_4 fanout5074 (.X(net5074),
    .A(net5077));
 sg13g2_buf_4 fanout5075 (.X(net5075),
    .A(net5077));
 sg13g2_buf_2 fanout5076 (.A(net5077),
    .X(net5076));
 sg13g2_buf_4 fanout5077 (.X(net5077),
    .A(_03034_));
 sg13g2_buf_8 fanout5078 (.A(net5082),
    .X(net5078));
 sg13g2_buf_2 fanout5079 (.A(net5082),
    .X(net5079));
 sg13g2_buf_4 fanout5080 (.X(net5080),
    .A(net5082));
 sg13g2_buf_1 fanout5081 (.A(net5082),
    .X(net5081));
 sg13g2_buf_8 fanout5082 (.A(_03033_),
    .X(net5082));
 sg13g2_buf_8 fanout5083 (.A(net5087),
    .X(net5083));
 sg13g2_buf_4 fanout5084 (.X(net5084),
    .A(net5085));
 sg13g2_buf_4 fanout5085 (.X(net5085),
    .A(net5086));
 sg13g2_buf_4 fanout5086 (.X(net5086),
    .A(net5087));
 sg13g2_buf_4 fanout5087 (.X(net5087),
    .A(_03033_));
 sg13g2_buf_4 fanout5088 (.X(net5088),
    .A(net5089));
 sg13g2_buf_4 fanout5089 (.X(net5089),
    .A(net5090));
 sg13g2_buf_4 fanout5090 (.X(net5090),
    .A(net5097));
 sg13g2_buf_4 fanout5091 (.X(net5091),
    .A(net5092));
 sg13g2_buf_4 fanout5092 (.X(net5092),
    .A(net5097));
 sg13g2_buf_4 fanout5093 (.X(net5093),
    .A(net5096));
 sg13g2_buf_4 fanout5094 (.X(net5094),
    .A(net5095));
 sg13g2_buf_4 fanout5095 (.X(net5095),
    .A(net5096));
 sg13g2_buf_4 fanout5096 (.X(net5096),
    .A(net5097));
 sg13g2_buf_2 fanout5097 (.A(_03016_),
    .X(net5097));
 sg13g2_buf_4 fanout5098 (.X(net5098),
    .A(net5102));
 sg13g2_buf_2 fanout5099 (.A(net5102),
    .X(net5099));
 sg13g2_buf_4 fanout5100 (.X(net5100),
    .A(net5101));
 sg13g2_buf_8 fanout5101 (.A(net5102),
    .X(net5101));
 sg13g2_buf_8 fanout5102 (.A(_03016_),
    .X(net5102));
 sg13g2_buf_8 fanout5103 (.A(net5106),
    .X(net5103));
 sg13g2_buf_4 fanout5104 (.X(net5104),
    .A(net5106));
 sg13g2_buf_2 fanout5105 (.A(net5106),
    .X(net5105));
 sg13g2_buf_8 fanout5106 (.A(_03015_),
    .X(net5106));
 sg13g2_buf_4 fanout5107 (.X(net5107),
    .A(net5112));
 sg13g2_buf_2 fanout5108 (.A(net5109),
    .X(net5108));
 sg13g2_buf_4 fanout5109 (.X(net5109),
    .A(net5110));
 sg13g2_buf_2 fanout5110 (.A(net5111),
    .X(net5110));
 sg13g2_buf_4 fanout5111 (.X(net5111),
    .A(net5112));
 sg13g2_buf_4 fanout5112 (.X(net5112),
    .A(_03015_));
 sg13g2_buf_4 fanout5113 (.X(net5113),
    .A(_10265_));
 sg13g2_buf_4 fanout5114 (.X(net5114),
    .A(_10233_));
 sg13g2_buf_4 fanout5115 (.X(net5115),
    .A(net5116));
 sg13g2_buf_4 fanout5116 (.X(net5116),
    .A(net5125));
 sg13g2_buf_2 fanout5117 (.A(net5125),
    .X(net5117));
 sg13g2_buf_4 fanout5118 (.X(net5118),
    .A(net5119));
 sg13g2_buf_4 fanout5119 (.X(net5119),
    .A(net5125));
 sg13g2_buf_4 fanout5120 (.X(net5120),
    .A(net5125));
 sg13g2_buf_4 fanout5121 (.X(net5121),
    .A(net5125));
 sg13g2_buf_4 fanout5122 (.X(net5122),
    .A(net5124));
 sg13g2_buf_2 fanout5123 (.A(net5124),
    .X(net5123));
 sg13g2_buf_4 fanout5124 (.X(net5124),
    .A(net5125));
 sg13g2_buf_4 fanout5125 (.X(net5125),
    .A(_08656_));
 sg13g2_buf_4 fanout5126 (.X(net5126),
    .A(net5127));
 sg13g2_buf_4 fanout5127 (.X(net5127),
    .A(net5128));
 sg13g2_buf_4 fanout5128 (.X(net5128),
    .A(net5130));
 sg13g2_buf_8 fanout5129 (.A(net5130),
    .X(net5129));
 sg13g2_buf_4 fanout5130 (.X(net5130),
    .A(_08656_));
 sg13g2_buf_8 fanout5131 (.A(net5134),
    .X(net5131));
 sg13g2_buf_4 fanout5132 (.X(net5132),
    .A(net5133));
 sg13g2_buf_4 fanout5133 (.X(net5133),
    .A(net5134));
 sg13g2_buf_8 fanout5134 (.A(net5140),
    .X(net5134));
 sg13g2_buf_8 fanout5135 (.A(net5140),
    .X(net5135));
 sg13g2_buf_4 fanout5136 (.X(net5136),
    .A(net5140));
 sg13g2_buf_4 fanout5137 (.X(net5137),
    .A(net5138));
 sg13g2_buf_2 fanout5138 (.A(net5139),
    .X(net5138));
 sg13g2_buf_4 fanout5139 (.X(net5139),
    .A(net5140));
 sg13g2_buf_8 fanout5140 (.A(_08655_),
    .X(net5140));
 sg13g2_buf_2 fanout5141 (.A(_05207_),
    .X(net5141));
 sg13g2_buf_2 fanout5142 (.A(net5143),
    .X(net5142));
 sg13g2_buf_2 fanout5143 (.A(_04063_),
    .X(net5143));
 sg13g2_buf_4 fanout5144 (.X(net5144),
    .A(_04061_));
 sg13g2_buf_2 fanout5145 (.A(_04061_),
    .X(net5145));
 sg13g2_buf_8 fanout5146 (.A(net5149),
    .X(net5146));
 sg13g2_buf_4 fanout5147 (.X(net5147),
    .A(net5149));
 sg13g2_buf_4 fanout5148 (.X(net5148),
    .A(net5149));
 sg13g2_buf_4 fanout5149 (.X(net5149),
    .A(net5156));
 sg13g2_buf_4 fanout5150 (.X(net5150),
    .A(net5156));
 sg13g2_buf_4 fanout5151 (.X(net5151),
    .A(net5156));
 sg13g2_buf_2 fanout5152 (.A(net5154),
    .X(net5152));
 sg13g2_buf_2 fanout5153 (.A(net5154),
    .X(net5153));
 sg13g2_buf_4 fanout5154 (.X(net5154),
    .A(net5155));
 sg13g2_buf_2 fanout5155 (.A(net5156),
    .X(net5155));
 sg13g2_buf_4 fanout5156 (.X(net5156),
    .A(_03028_));
 sg13g2_buf_4 fanout5157 (.X(net5157),
    .A(net5158));
 sg13g2_buf_4 fanout5158 (.X(net5158),
    .A(net5161));
 sg13g2_buf_4 fanout5159 (.X(net5159),
    .A(net5160));
 sg13g2_buf_4 fanout5160 (.X(net5160),
    .A(net5161));
 sg13g2_buf_2 fanout5161 (.A(net5172),
    .X(net5161));
 sg13g2_buf_4 fanout5162 (.X(net5162),
    .A(net5164));
 sg13g2_buf_4 fanout5163 (.X(net5163),
    .A(net5164));
 sg13g2_buf_4 fanout5164 (.X(net5164),
    .A(net5172));
 sg13g2_buf_4 fanout5165 (.X(net5165),
    .A(net5168));
 sg13g2_buf_4 fanout5166 (.X(net5166),
    .A(net5168));
 sg13g2_buf_1 fanout5167 (.A(net5168),
    .X(net5167));
 sg13g2_buf_2 fanout5168 (.A(net5169),
    .X(net5168));
 sg13g2_buf_2 fanout5169 (.A(net5172),
    .X(net5169));
 sg13g2_buf_4 fanout5170 (.X(net5170),
    .A(net5171));
 sg13g2_buf_2 fanout5171 (.A(net5172),
    .X(net5171));
 sg13g2_buf_8 fanout5172 (.A(_03027_),
    .X(net5172));
 sg13g2_buf_4 fanout5173 (.X(net5173),
    .A(net5175));
 sg13g2_buf_4 fanout5174 (.X(net5174),
    .A(net5175));
 sg13g2_buf_4 fanout5175 (.X(net5175),
    .A(_03022_));
 sg13g2_buf_4 fanout5176 (.X(net5176),
    .A(net5178));
 sg13g2_buf_4 fanout5177 (.X(net5177),
    .A(net5178));
 sg13g2_buf_4 fanout5178 (.X(net5178),
    .A(_03022_));
 sg13g2_buf_4 fanout5179 (.X(net5179),
    .A(net5180));
 sg13g2_buf_8 fanout5180 (.A(net5184),
    .X(net5180));
 sg13g2_buf_4 fanout5181 (.X(net5181),
    .A(net5183));
 sg13g2_buf_2 fanout5182 (.A(net5183),
    .X(net5182));
 sg13g2_buf_4 fanout5183 (.X(net5183),
    .A(net5184));
 sg13g2_buf_4 fanout5184 (.X(net5184),
    .A(_03022_));
 sg13g2_buf_4 fanout5185 (.X(net5185),
    .A(net5187));
 sg13g2_buf_4 fanout5186 (.X(net5186),
    .A(net5187));
 sg13g2_buf_4 fanout5187 (.X(net5187),
    .A(net5191));
 sg13g2_buf_4 fanout5188 (.X(net5188),
    .A(net5190));
 sg13g2_buf_4 fanout5189 (.X(net5189),
    .A(net5190));
 sg13g2_buf_8 fanout5190 (.A(net5191),
    .X(net5190));
 sg13g2_buf_2 fanout5191 (.A(net5196),
    .X(net5191));
 sg13g2_buf_4 fanout5192 (.X(net5192),
    .A(net5194));
 sg13g2_buf_4 fanout5193 (.X(net5193),
    .A(net5194));
 sg13g2_buf_2 fanout5194 (.A(net5196),
    .X(net5194));
 sg13g2_buf_4 fanout5195 (.X(net5195),
    .A(net5196));
 sg13g2_buf_8 fanout5196 (.A(_03021_),
    .X(net5196));
 sg13g2_buf_2 fanout5197 (.A(net5198),
    .X(net5197));
 sg13g2_buf_2 fanout5198 (.A(_09660_),
    .X(net5198));
 sg13g2_buf_4 fanout5199 (.X(net5199),
    .A(_08247_));
 sg13g2_buf_2 fanout5200 (.A(net5201),
    .X(net5200));
 sg13g2_buf_2 fanout5201 (.A(_08222_),
    .X(net5201));
 sg13g2_buf_4 fanout5202 (.X(net5202),
    .A(_08203_));
 sg13g2_buf_2 fanout5203 (.A(_08184_),
    .X(net5203));
 sg13g2_buf_2 fanout5204 (.A(net5206),
    .X(net5204));
 sg13g2_buf_2 fanout5205 (.A(net5206),
    .X(net5205));
 sg13g2_buf_2 fanout5206 (.A(_08179_),
    .X(net5206));
 sg13g2_buf_2 fanout5207 (.A(net5209),
    .X(net5207));
 sg13g2_buf_2 fanout5208 (.A(net5209),
    .X(net5208));
 sg13g2_buf_2 fanout5209 (.A(_05242_),
    .X(net5209));
 sg13g2_buf_4 fanout5210 (.X(net5210),
    .A(net5211));
 sg13g2_buf_4 fanout5211 (.X(net5211),
    .A(_04891_));
 sg13g2_buf_4 fanout5212 (.X(net5212),
    .A(_04054_));
 sg13g2_buf_2 fanout5213 (.A(net5214),
    .X(net5213));
 sg13g2_buf_4 fanout5214 (.X(net5214),
    .A(_04040_));
 sg13g2_buf_2 fanout5215 (.A(_03446_),
    .X(net5215));
 sg13g2_buf_4 fanout5216 (.X(net5216),
    .A(_09826_));
 sg13g2_buf_4 fanout5217 (.X(net5217),
    .A(net5218));
 sg13g2_buf_4 fanout5218 (.X(net5218),
    .A(net5219));
 sg13g2_buf_2 fanout5219 (.A(net5227),
    .X(net5219));
 sg13g2_buf_4 fanout5220 (.X(net5220),
    .A(net5227));
 sg13g2_buf_4 fanout5221 (.X(net5221),
    .A(net5227));
 sg13g2_buf_4 fanout5222 (.X(net5222),
    .A(net5226));
 sg13g2_buf_4 fanout5223 (.X(net5223),
    .A(net5226));
 sg13g2_buf_4 fanout5224 (.X(net5224),
    .A(net5226));
 sg13g2_buf_2 fanout5225 (.A(net5226),
    .X(net5225));
 sg13g2_buf_4 fanout5226 (.X(net5226),
    .A(net5227));
 sg13g2_buf_2 fanout5227 (.A(net5233),
    .X(net5227));
 sg13g2_buf_4 fanout5228 (.X(net5228),
    .A(net5229));
 sg13g2_buf_4 fanout5229 (.X(net5229),
    .A(net5230));
 sg13g2_buf_4 fanout5230 (.X(net5230),
    .A(net5233));
 sg13g2_buf_4 fanout5231 (.X(net5231),
    .A(net5232));
 sg13g2_buf_8 fanout5232 (.A(net5233),
    .X(net5232));
 sg13g2_buf_8 fanout5233 (.A(_08665_),
    .X(net5233));
 sg13g2_buf_8 fanout5234 (.A(net5237),
    .X(net5234));
 sg13g2_buf_4 fanout5235 (.X(net5235),
    .A(net5237));
 sg13g2_buf_2 fanout5236 (.A(net5237),
    .X(net5236));
 sg13g2_buf_8 fanout5237 (.A(_08664_),
    .X(net5237));
 sg13g2_buf_4 fanout5238 (.X(net5238),
    .A(net5239));
 sg13g2_buf_4 fanout5239 (.X(net5239),
    .A(net5243));
 sg13g2_buf_4 fanout5240 (.X(net5240),
    .A(net5242));
 sg13g2_buf_1 fanout5241 (.A(net5242),
    .X(net5241));
 sg13g2_buf_4 fanout5242 (.X(net5242),
    .A(net5243));
 sg13g2_buf_4 fanout5243 (.X(net5243),
    .A(_08664_));
 sg13g2_buf_4 fanout5244 (.X(net5244),
    .A(net5245));
 sg13g2_buf_4 fanout5245 (.X(net5245),
    .A(net5250));
 sg13g2_buf_4 fanout5246 (.X(net5246),
    .A(net5249));
 sg13g2_buf_2 fanout5247 (.A(net5249),
    .X(net5247));
 sg13g2_buf_4 fanout5248 (.X(net5248),
    .A(net5249));
 sg13g2_buf_2 fanout5249 (.A(net5250),
    .X(net5249));
 sg13g2_buf_2 fanout5250 (.A(net5259),
    .X(net5250));
 sg13g2_buf_4 fanout5251 (.X(net5251),
    .A(net5253));
 sg13g2_buf_2 fanout5252 (.A(net5253),
    .X(net5252));
 sg13g2_buf_4 fanout5253 (.X(net5253),
    .A(net5254));
 sg13g2_buf_8 fanout5254 (.A(net5259),
    .X(net5254));
 sg13g2_buf_4 fanout5255 (.X(net5255),
    .A(net5256));
 sg13g2_buf_4 fanout5256 (.X(net5256),
    .A(net5257));
 sg13g2_buf_4 fanout5257 (.X(net5257),
    .A(net5259));
 sg13g2_buf_4 fanout5258 (.X(net5258),
    .A(net5259));
 sg13g2_buf_8 fanout5259 (.A(_08649_),
    .X(net5259));
 sg13g2_buf_8 fanout5260 (.A(net5263),
    .X(net5260));
 sg13g2_buf_4 fanout5261 (.X(net5261),
    .A(net5262));
 sg13g2_buf_8 fanout5262 (.A(net5263),
    .X(net5262));
 sg13g2_buf_8 fanout5263 (.A(net5269),
    .X(net5263));
 sg13g2_buf_8 fanout5264 (.A(net5269),
    .X(net5264));
 sg13g2_buf_4 fanout5265 (.X(net5265),
    .A(net5269));
 sg13g2_buf_4 fanout5266 (.X(net5266),
    .A(net5267));
 sg13g2_buf_2 fanout5267 (.A(net5268),
    .X(net5267));
 sg13g2_buf_4 fanout5268 (.X(net5268),
    .A(net5269));
 sg13g2_buf_8 fanout5269 (.A(_08648_),
    .X(net5269));
 sg13g2_buf_2 fanout5270 (.A(net5271),
    .X(net5270));
 sg13g2_buf_4 fanout5271 (.X(net5271),
    .A(_08213_));
 sg13g2_buf_2 fanout5272 (.A(_08213_),
    .X(net5272));
 sg13g2_buf_4 fanout5273 (.X(net5273),
    .A(\atari2600.cpu.DIMUX[7] ));
 sg13g2_buf_4 fanout5274 (.X(net5274),
    .A(_08176_));
 sg13g2_buf_2 fanout5275 (.A(_08176_),
    .X(net5275));
 sg13g2_buf_2 fanout5276 (.A(net5277),
    .X(net5276));
 sg13g2_buf_2 fanout5277 (.A(net5278),
    .X(net5277));
 sg13g2_buf_4 fanout5278 (.X(net5278),
    .A(net5279));
 sg13g2_buf_2 fanout5279 (.A(net5280),
    .X(net5279));
 sg13g2_buf_4 fanout5280 (.X(net5280),
    .A(_05495_));
 sg13g2_buf_2 fanout5281 (.A(_04088_),
    .X(net5281));
 sg13g2_buf_4 fanout5282 (.X(net5282),
    .A(_04067_));
 sg13g2_buf_2 fanout5283 (.A(_04049_),
    .X(net5283));
 sg13g2_buf_4 fanout5284 (.X(net5284),
    .A(_04043_));
 sg13g2_buf_2 fanout5285 (.A(_03941_),
    .X(net5285));
 sg13g2_buf_1 fanout5286 (.A(_03941_),
    .X(net5286));
 sg13g2_buf_2 fanout5287 (.A(net5288),
    .X(net5287));
 sg13g2_buf_2 fanout5288 (.A(_03540_),
    .X(net5288));
 sg13g2_buf_2 fanout5289 (.A(_03540_),
    .X(net5289));
 sg13g2_buf_2 fanout5290 (.A(_03540_),
    .X(net5290));
 sg13g2_buf_2 fanout5291 (.A(net5293),
    .X(net5291));
 sg13g2_buf_4 fanout5292 (.X(net5292),
    .A(net5298));
 sg13g2_buf_1 fanout5293 (.A(net5298),
    .X(net5293));
 sg13g2_buf_2 fanout5294 (.A(net5295),
    .X(net5294));
 sg13g2_buf_2 fanout5295 (.A(net5298),
    .X(net5295));
 sg13g2_buf_2 fanout5296 (.A(net5298),
    .X(net5296));
 sg13g2_buf_2 fanout5297 (.A(net5298),
    .X(net5297));
 sg13g2_buf_2 fanout5298 (.A(_03539_),
    .X(net5298));
 sg13g2_buf_4 fanout5299 (.X(net5299),
    .A(net5300));
 sg13g2_buf_2 fanout5300 (.A(_03445_),
    .X(net5300));
 sg13g2_buf_2 fanout5301 (.A(_03445_),
    .X(net5301));
 sg13g2_buf_2 fanout5302 (.A(_03445_),
    .X(net5302));
 sg13g2_buf_2 fanout5303 (.A(net5305),
    .X(net5303));
 sg13g2_buf_2 fanout5304 (.A(net5305),
    .X(net5304));
 sg13g2_buf_2 fanout5305 (.A(_08671_),
    .X(net5305));
 sg13g2_buf_2 fanout5306 (.A(_08671_),
    .X(net5306));
 sg13g2_buf_4 fanout5307 (.X(net5307),
    .A(net5309));
 sg13g2_buf_2 fanout5308 (.A(net5309),
    .X(net5308));
 sg13g2_buf_2 fanout5309 (.A(_08534_),
    .X(net5309));
 sg13g2_buf_2 fanout5310 (.A(net5311),
    .X(net5310));
 sg13g2_buf_2 fanout5311 (.A(net5312),
    .X(net5311));
 sg13g2_buf_4 fanout5312 (.X(net5312),
    .A(net5315));
 sg13g2_buf_4 fanout5313 (.X(net5313),
    .A(net5315));
 sg13g2_buf_2 fanout5314 (.A(net5315),
    .X(net5314));
 sg13g2_buf_4 fanout5315 (.X(net5315),
    .A(_08165_));
 sg13g2_buf_4 fanout5316 (.X(net5316),
    .A(_08163_));
 sg13g2_buf_4 fanout5317 (.X(net5317),
    .A(_07461_));
 sg13g2_buf_2 fanout5318 (.A(_07240_),
    .X(net5318));
 sg13g2_buf_2 fanout5319 (.A(_07240_),
    .X(net5319));
 sg13g2_buf_2 fanout5320 (.A(_06016_),
    .X(net5320));
 sg13g2_buf_2 fanout5321 (.A(_05642_),
    .X(net5321));
 sg13g2_buf_4 fanout5322 (.X(net5322),
    .A(_05204_));
 sg13g2_buf_2 fanout5323 (.A(_05130_),
    .X(net5323));
 sg13g2_buf_2 fanout5324 (.A(_05130_),
    .X(net5324));
 sg13g2_buf_4 fanout5325 (.X(net5325),
    .A(_04085_));
 sg13g2_buf_4 fanout5326 (.X(net5326),
    .A(_03934_));
 sg13g2_buf_2 fanout5327 (.A(_03934_),
    .X(net5327));
 sg13g2_buf_4 fanout5328 (.X(net5328),
    .A(_03930_));
 sg13g2_buf_1 fanout5329 (.A(_03930_),
    .X(net5329));
 sg13g2_buf_4 fanout5330 (.X(net5330),
    .A(_03928_));
 sg13g2_buf_2 fanout5331 (.A(_03733_),
    .X(net5331));
 sg13g2_buf_4 fanout5332 (.X(net5332),
    .A(net5336));
 sg13g2_buf_2 fanout5333 (.A(net5335),
    .X(net5333));
 sg13g2_buf_1 fanout5334 (.A(net5335),
    .X(net5334));
 sg13g2_buf_2 fanout5335 (.A(net5336),
    .X(net5335));
 sg13g2_buf_2 fanout5336 (.A(_03636_),
    .X(net5336));
 sg13g2_buf_2 fanout5337 (.A(net5339),
    .X(net5337));
 sg13g2_buf_2 fanout5338 (.A(net5339),
    .X(net5338));
 sg13g2_buf_2 fanout5339 (.A(_03635_),
    .X(net5339));
 sg13g2_buf_2 fanout5340 (.A(_03635_),
    .X(net5340));
 sg13g2_buf_1 fanout5341 (.A(net5342),
    .X(net5341));
 sg13g2_buf_2 fanout5342 (.A(_03635_),
    .X(net5342));
 sg13g2_buf_4 fanout5343 (.X(net5343),
    .A(net5344));
 sg13g2_buf_4 fanout5344 (.X(net5344),
    .A(_08670_));
 sg13g2_buf_2 fanout5345 (.A(_08529_),
    .X(net5345));
 sg13g2_buf_2 fanout5346 (.A(net5348),
    .X(net5346));
 sg13g2_buf_2 fanout5347 (.A(net5348),
    .X(net5347));
 sg13g2_buf_2 fanout5348 (.A(_08214_),
    .X(net5348));
 sg13g2_buf_4 fanout5349 (.X(net5349),
    .A(_08214_));
 sg13g2_buf_2 fanout5350 (.A(_08214_),
    .X(net5350));
 sg13g2_buf_4 fanout5351 (.X(net5351),
    .A(net7363));
 sg13g2_buf_4 fanout5352 (.X(net5352),
    .A(net5354));
 sg13g2_buf_4 fanout5353 (.X(net5353),
    .A(net5354));
 sg13g2_buf_8 fanout5354 (.A(_08162_),
    .X(net5354));
 sg13g2_buf_2 fanout5355 (.A(net5357),
    .X(net5355));
 sg13g2_buf_2 fanout5356 (.A(net5357),
    .X(net5356));
 sg13g2_buf_1 fanout5357 (.A(_05133_),
    .X(net5357));
 sg13g2_buf_2 fanout5358 (.A(_05131_),
    .X(net5358));
 sg13g2_buf_1 fanout5359 (.A(_05131_),
    .X(net5359));
 sg13g2_buf_4 fanout5360 (.X(net5360),
    .A(_03731_));
 sg13g2_buf_4 fanout5361 (.X(net5361),
    .A(_08522_));
 sg13g2_buf_2 fanout5362 (.A(net5363),
    .X(net5362));
 sg13g2_buf_4 fanout5363 (.X(net5363),
    .A(net5384));
 sg13g2_buf_2 fanout5364 (.A(net5367),
    .X(net5364));
 sg13g2_buf_2 fanout5365 (.A(net5367),
    .X(net5365));
 sg13g2_buf_1 fanout5366 (.A(net5367),
    .X(net5366));
 sg13g2_buf_2 fanout5367 (.A(net5384),
    .X(net5367));
 sg13g2_buf_2 fanout5368 (.A(net5369),
    .X(net5368));
 sg13g2_buf_1 fanout5369 (.A(net5373),
    .X(net5369));
 sg13g2_buf_2 fanout5370 (.A(net5373),
    .X(net5370));
 sg13g2_buf_1 fanout5371 (.A(net5373),
    .X(net5371));
 sg13g2_buf_2 fanout5372 (.A(net5373),
    .X(net5372));
 sg13g2_buf_1 fanout5373 (.A(net5379),
    .X(net5373));
 sg13g2_buf_2 fanout5374 (.A(net5375),
    .X(net5374));
 sg13g2_buf_2 fanout5375 (.A(net5378),
    .X(net5375));
 sg13g2_buf_2 fanout5376 (.A(net5377),
    .X(net5376));
 sg13g2_buf_1 fanout5377 (.A(net5378),
    .X(net5377));
 sg13g2_buf_2 fanout5378 (.A(net5379),
    .X(net5378));
 sg13g2_buf_2 fanout5379 (.A(net5380),
    .X(net5379));
 sg13g2_buf_2 fanout5380 (.A(net5383),
    .X(net5380));
 sg13g2_buf_2 fanout5381 (.A(net5382),
    .X(net5381));
 sg13g2_buf_4 fanout5382 (.X(net5382),
    .A(net5383));
 sg13g2_buf_2 fanout5383 (.A(net5384),
    .X(net5383));
 sg13g2_buf_4 fanout5384 (.X(net5384),
    .A(_08164_));
 sg13g2_buf_2 fanout5385 (.A(_08160_),
    .X(net5385));
 sg13g2_buf_2 fanout5386 (.A(_08160_),
    .X(net5386));
 sg13g2_buf_2 fanout5387 (.A(net5388),
    .X(net5387));
 sg13g2_buf_2 fanout5388 (.A(_04874_),
    .X(net5388));
 sg13g2_buf_2 fanout5389 (.A(_10196_),
    .X(net5389));
 sg13g2_buf_4 fanout5390 (.X(net5390),
    .A(_10190_));
 sg13g2_buf_1 fanout5391 (.A(_10190_),
    .X(net5391));
 sg13g2_buf_2 fanout5392 (.A(_08532_),
    .X(net5392));
 sg13g2_buf_2 fanout5393 (.A(net5395),
    .X(net5393));
 sg13g2_buf_2 fanout5394 (.A(net5395),
    .X(net5394));
 sg13g2_buf_2 fanout5395 (.A(_10448_),
    .X(net5395));
 sg13g2_buf_2 fanout5396 (.A(_08531_),
    .X(net5396));
 sg13g2_buf_2 fanout5397 (.A(_08519_),
    .X(net5397));
 sg13g2_buf_2 fanout5398 (.A(_08500_),
    .X(net5398));
 sg13g2_buf_4 fanout5399 (.X(net5399),
    .A(_07819_));
 sg13g2_buf_2 fanout5400 (.A(_06054_),
    .X(net5400));
 sg13g2_buf_2 fanout5401 (.A(_05570_),
    .X(net5401));
 sg13g2_buf_4 fanout5402 (.X(net5402),
    .A(_04881_));
 sg13g2_buf_2 fanout5403 (.A(net5405),
    .X(net5403));
 sg13g2_buf_2 fanout5404 (.A(net5405),
    .X(net5404));
 sg13g2_buf_2 fanout5405 (.A(_03350_),
    .X(net5405));
 sg13g2_buf_4 fanout5406 (.X(net5406),
    .A(_03350_));
 sg13g2_buf_4 fanout5407 (.X(net5407),
    .A(_03349_));
 sg13g2_buf_2 fanout5408 (.A(_03349_),
    .X(net5408));
 sg13g2_buf_4 fanout5409 (.X(net5409),
    .A(net5410));
 sg13g2_buf_2 fanout5410 (.A(_03349_),
    .X(net5410));
 sg13g2_buf_8 fanout5411 (.A(_03124_),
    .X(net5411));
 sg13g2_buf_8 fanout5412 (.A(_03113_),
    .X(net5412));
 sg13g2_buf_4 fanout5413 (.X(net5413),
    .A(_03105_));
 sg13g2_buf_4 fanout5414 (.X(net5414),
    .A(_03082_));
 sg13g2_buf_4 fanout5415 (.X(net5415),
    .A(_03079_));
 sg13g2_buf_8 fanout5416 (.A(_03074_),
    .X(net5416));
 sg13g2_buf_4 fanout5417 (.X(net5417),
    .A(net5418));
 sg13g2_buf_4 fanout5418 (.X(net5418),
    .A(_03072_));
 sg13g2_buf_8 fanout5419 (.A(_10507_),
    .X(net5419));
 sg13g2_buf_4 fanout5420 (.X(net5420),
    .A(net5421));
 sg13g2_buf_4 fanout5421 (.X(net5421),
    .A(_10501_));
 sg13g2_buf_4 fanout5422 (.X(net5422),
    .A(_10498_));
 sg13g2_buf_2 fanout5423 (.A(_10498_),
    .X(net5423));
 sg13g2_buf_8 fanout5424 (.A(_10497_),
    .X(net5424));
 sg13g2_buf_4 fanout5425 (.X(net5425),
    .A(_10481_));
 sg13g2_buf_2 fanout5426 (.A(net5429),
    .X(net5426));
 sg13g2_buf_1 fanout5427 (.A(net5429),
    .X(net5427));
 sg13g2_buf_2 fanout5428 (.A(net5429),
    .X(net5428));
 sg13g2_buf_2 fanout5429 (.A(_10447_),
    .X(net5429));
 sg13g2_buf_4 fanout5430 (.X(net5430),
    .A(_10384_));
 sg13g2_buf_4 fanout5431 (.X(net5431),
    .A(_10376_));
 sg13g2_buf_2 fanout5432 (.A(_10376_),
    .X(net5432));
 sg13g2_buf_2 fanout5433 (.A(_08497_),
    .X(net5433));
 sg13g2_buf_2 fanout5434 (.A(_08496_),
    .X(net5434));
 sg13g2_buf_4 fanout5435 (.X(net5435),
    .A(_08413_));
 sg13g2_buf_4 fanout5436 (.X(net5436),
    .A(_08389_));
 sg13g2_buf_4 fanout5437 (.X(net5437),
    .A(_08363_));
 sg13g2_buf_2 fanout5438 (.A(_08363_),
    .X(net5438));
 sg13g2_buf_2 fanout5439 (.A(net5440),
    .X(net5439));
 sg13g2_buf_2 fanout5440 (.A(_08362_),
    .X(net5440));
 sg13g2_buf_2 fanout5441 (.A(net5443),
    .X(net5441));
 sg13g2_buf_1 fanout5442 (.A(net5443),
    .X(net5442));
 sg13g2_buf_2 fanout5443 (.A(net5444),
    .X(net5443));
 sg13g2_buf_2 fanout5444 (.A(_08361_),
    .X(net5444));
 sg13g2_buf_2 fanout5445 (.A(_08335_),
    .X(net5445));
 sg13g2_buf_2 fanout5446 (.A(_06076_),
    .X(net5446));
 sg13g2_buf_2 fanout5447 (.A(_06005_),
    .X(net5447));
 sg13g2_buf_1 fanout5448 (.A(_06005_),
    .X(net5448));
 sg13g2_buf_2 fanout5449 (.A(_05957_),
    .X(net5449));
 sg13g2_buf_2 fanout5450 (.A(_05957_),
    .X(net5450));
 sg13g2_buf_2 fanout5451 (.A(net5452),
    .X(net5451));
 sg13g2_buf_1 fanout5452 (.A(_05956_),
    .X(net5452));
 sg13g2_buf_4 fanout5453 (.X(net5453),
    .A(_05553_));
 sg13g2_buf_4 fanout5454 (.X(net5454),
    .A(_05552_));
 sg13g2_buf_4 fanout5455 (.X(net5455),
    .A(_03393_));
 sg13g2_buf_4 fanout5456 (.X(net5456),
    .A(net5458));
 sg13g2_buf_2 fanout5457 (.A(net5458),
    .X(net5457));
 sg13g2_buf_4 fanout5458 (.X(net5458),
    .A(net5462));
 sg13g2_buf_2 fanout5459 (.A(net5462),
    .X(net5459));
 sg13g2_buf_2 fanout5460 (.A(net5461),
    .X(net5460));
 sg13g2_buf_4 fanout5461 (.X(net5461),
    .A(net5462));
 sg13g2_buf_2 fanout5462 (.A(_03347_),
    .X(net5462));
 sg13g2_buf_2 fanout5463 (.A(net5466),
    .X(net5463));
 sg13g2_buf_2 fanout5464 (.A(net5465),
    .X(net5464));
 sg13g2_buf_2 fanout5465 (.A(net5466),
    .X(net5465));
 sg13g2_buf_2 fanout5466 (.A(_03233_),
    .X(net5466));
 sg13g2_buf_8 fanout5467 (.A(_02998_),
    .X(net5467));
 sg13g2_buf_8 fanout5468 (.A(_10509_),
    .X(net5468));
 sg13g2_buf_4 fanout5469 (.X(net5469),
    .A(net5470));
 sg13g2_buf_4 fanout5470 (.X(net5470),
    .A(_10506_));
 sg13g2_buf_8 fanout5471 (.A(_10504_),
    .X(net5471));
 sg13g2_buf_8 fanout5472 (.A(_10334_),
    .X(net5472));
 sg13g2_buf_8 fanout5473 (.A(_10334_),
    .X(net5473));
 sg13g2_buf_4 fanout5474 (.X(net5474),
    .A(_10211_));
 sg13g2_buf_4 fanout5475 (.X(net5475),
    .A(_08314_));
 sg13g2_buf_2 fanout5476 (.A(_08257_),
    .X(net5476));
 sg13g2_buf_2 fanout5477 (.A(_08257_),
    .X(net5477));
 sg13g2_buf_4 fanout5478 (.X(net5478),
    .A(_08256_));
 sg13g2_buf_4 fanout5479 (.X(net5479),
    .A(_08231_));
 sg13g2_buf_4 fanout5480 (.X(net5480),
    .A(_08211_));
 sg13g2_buf_2 fanout5481 (.A(net5482),
    .X(net5481));
 sg13g2_buf_2 fanout5482 (.A(_05564_),
    .X(net5482));
 sg13g2_buf_2 fanout5483 (.A(net5484),
    .X(net5483));
 sg13g2_buf_4 fanout5484 (.X(net5484),
    .A(net5485));
 sg13g2_buf_8 fanout5485 (.A(_03357_),
    .X(net5485));
 sg13g2_buf_4 fanout5486 (.X(net5486),
    .A(net5488));
 sg13g2_buf_2 fanout5487 (.A(net5488),
    .X(net5487));
 sg13g2_buf_2 fanout5488 (.A(_03356_),
    .X(net5488));
 sg13g2_buf_4 fanout5489 (.X(net5489),
    .A(net5490));
 sg13g2_buf_4 fanout5490 (.X(net5490),
    .A(net5494));
 sg13g2_buf_4 fanout5491 (.X(net5491),
    .A(net5492));
 sg13g2_buf_4 fanout5492 (.X(net5492),
    .A(net5493));
 sg13g2_buf_4 fanout5493 (.X(net5493),
    .A(net5494));
 sg13g2_buf_4 fanout5494 (.X(net5494),
    .A(_03356_));
 sg13g2_buf_2 fanout5495 (.A(_03234_),
    .X(net5495));
 sg13g2_buf_2 fanout5496 (.A(_03234_),
    .X(net5496));
 sg13g2_buf_4 fanout5497 (.X(net5497),
    .A(net5499));
 sg13g2_buf_2 fanout5498 (.A(net5499),
    .X(net5498));
 sg13g2_buf_8 fanout5499 (.A(_03228_),
    .X(net5499));
 sg13g2_buf_4 fanout5500 (.X(net5500),
    .A(net5503));
 sg13g2_buf_2 fanout5501 (.A(net5503),
    .X(net5501));
 sg13g2_buf_4 fanout5502 (.X(net5502),
    .A(net5503));
 sg13g2_buf_2 fanout5503 (.A(_03227_),
    .X(net5503));
 sg13g2_buf_4 fanout5504 (.X(net5504),
    .A(net5508));
 sg13g2_buf_4 fanout5505 (.X(net5505),
    .A(net5508));
 sg13g2_buf_4 fanout5506 (.X(net5506),
    .A(net5507));
 sg13g2_buf_4 fanout5507 (.X(net5507),
    .A(net5508));
 sg13g2_buf_4 fanout5508 (.X(net5508),
    .A(_03227_));
 sg13g2_buf_8 fanout5509 (.A(_03225_),
    .X(net5509));
 sg13g2_buf_2 fanout5510 (.A(_03225_),
    .X(net5510));
 sg13g2_buf_4 fanout5511 (.X(net5511),
    .A(_10210_));
 sg13g2_buf_4 fanout5512 (.X(net5512),
    .A(net5513));
 sg13g2_buf_2 fanout5513 (.A(_08698_),
    .X(net5513));
 sg13g2_buf_4 fanout5514 (.X(net5514),
    .A(net5516));
 sg13g2_buf_2 fanout5515 (.A(net5516),
    .X(net5515));
 sg13g2_buf_4 fanout5516 (.X(net5516),
    .A(_08693_));
 sg13g2_buf_4 fanout5517 (.X(net5517),
    .A(net5519));
 sg13g2_buf_2 fanout5518 (.A(net5519),
    .X(net5518));
 sg13g2_buf_4 fanout5519 (.X(net5519),
    .A(_08692_));
 sg13g2_buf_4 fanout5520 (.X(net5520),
    .A(net5521));
 sg13g2_buf_4 fanout5521 (.X(net5521),
    .A(net5524));
 sg13g2_buf_4 fanout5522 (.X(net5522),
    .A(net5523));
 sg13g2_buf_4 fanout5523 (.X(net5523),
    .A(net5524));
 sg13g2_buf_4 fanout5524 (.X(net5524),
    .A(_08692_));
 sg13g2_buf_2 fanout5525 (.A(net5526),
    .X(net5525));
 sg13g2_buf_2 fanout5526 (.A(net5527),
    .X(net5526));
 sg13g2_buf_2 fanout5527 (.A(net5528),
    .X(net5527));
 sg13g2_buf_4 fanout5528 (.X(net5528),
    .A(_08689_));
 sg13g2_buf_4 fanout5529 (.X(net5529),
    .A(net5530));
 sg13g2_buf_4 fanout5530 (.X(net5530),
    .A(net5531));
 sg13g2_buf_4 fanout5531 (.X(net5531),
    .A(_08688_));
 sg13g2_buf_4 fanout5532 (.X(net5532),
    .A(net5536));
 sg13g2_buf_2 fanout5533 (.A(net5536),
    .X(net5533));
 sg13g2_buf_4 fanout5534 (.X(net5534),
    .A(net5535));
 sg13g2_buf_4 fanout5535 (.X(net5535),
    .A(net5536));
 sg13g2_buf_4 fanout5536 (.X(net5536),
    .A(_08688_));
 sg13g2_buf_2 fanout5537 (.A(\flash_rom.spi_select ),
    .X(net5537));
 sg13g2_buf_2 fanout5538 (.A(_08277_),
    .X(net5538));
 sg13g2_buf_2 fanout5539 (.A(_08228_),
    .X(net5539));
 sg13g2_buf_2 fanout5540 (.A(_08227_),
    .X(net5540));
 sg13g2_buf_4 fanout5541 (.X(net5541),
    .A(_08226_));
 sg13g2_buf_2 fanout5542 (.A(_08225_),
    .X(net5542));
 sg13g2_buf_1 fanout5543 (.A(_08225_),
    .X(net5543));
 sg13g2_buf_2 fanout5544 (.A(_08209_),
    .X(net5544));
 sg13g2_buf_4 fanout5545 (.X(net5545),
    .A(_08208_));
 sg13g2_buf_2 fanout5546 (.A(_08208_),
    .X(net5546));
 sg13g2_buf_2 fanout5547 (.A(_08207_),
    .X(net5547));
 sg13g2_buf_2 fanout5548 (.A(_08170_),
    .X(net5548));
 sg13g2_buf_2 fanout5549 (.A(_08168_),
    .X(net5549));
 sg13g2_buf_4 fanout5550 (.X(net5550),
    .A(_08167_));
 sg13g2_buf_2 fanout5551 (.A(_08166_),
    .X(net5551));
 sg13g2_buf_4 fanout5552 (.X(net5552),
    .A(_08119_));
 sg13g2_buf_4 fanout5553 (.X(net5553),
    .A(net5556));
 sg13g2_buf_4 fanout5554 (.X(net5554),
    .A(net5556));
 sg13g2_buf_4 fanout5555 (.X(net5555),
    .A(net5556));
 sg13g2_buf_2 fanout5556 (.A(_08118_),
    .X(net5556));
 sg13g2_buf_4 fanout5557 (.X(net5557),
    .A(_08114_));
 sg13g2_buf_4 fanout5558 (.X(net5558),
    .A(_08113_));
 sg13g2_buf_4 fanout5559 (.X(net5559),
    .A(_08112_));
 sg13g2_buf_4 fanout5560 (.X(net5560),
    .A(_08111_));
 sg13g2_buf_4 fanout5561 (.X(net5561),
    .A(net5562));
 sg13g2_buf_4 fanout5562 (.X(net5562),
    .A(_08110_));
 sg13g2_buf_4 fanout5563 (.X(net5563),
    .A(_08109_));
 sg13g2_buf_4 fanout5564 (.X(net5564),
    .A(_08109_));
 sg13g2_buf_2 fanout5565 (.A(_08009_),
    .X(net5565));
 sg13g2_buf_2 fanout5566 (.A(_08009_),
    .X(net5566));
 sg13g2_buf_2 fanout5567 (.A(net7357),
    .X(net5567));
 sg13g2_buf_4 fanout5568 (.X(net5568),
    .A(net7344));
 sg13g2_buf_4 fanout5569 (.X(net5569),
    .A(net7322));
 sg13g2_buf_4 fanout5570 (.X(net5570),
    .A(net7325));
 sg13g2_buf_4 fanout5571 (.X(net5571),
    .A(net7361));
 sg13g2_buf_4 fanout5572 (.X(net5572),
    .A(net7374));
 sg13g2_buf_2 fanout5573 (.A(net5575),
    .X(net5573));
 sg13g2_buf_1 fanout5574 (.A(net5575),
    .X(net5574));
 sg13g2_buf_2 fanout5575 (.A(net5576),
    .X(net5575));
 sg13g2_buf_2 fanout5576 (.A(\atari2600.cpu.IRHOLD_valid ),
    .X(net5576));
 sg13g2_buf_2 fanout5577 (.A(net7367),
    .X(net5577));
 sg13g2_buf_2 fanout5578 (.A(net7354),
    .X(net5578));
 sg13g2_buf_2 fanout5579 (.A(net7343),
    .X(net5579));
 sg13g2_buf_2 fanout5580 (.A(net5581),
    .X(net5580));
 sg13g2_buf_1 fanout5581 (.A(net7262),
    .X(net5581));
 sg13g2_buf_2 fanout5582 (.A(\atari2600.tia.audf0[0] ),
    .X(net5582));
 sg13g2_buf_2 fanout5583 (.A(net7351),
    .X(net5583));
 sg13g2_buf_2 fanout5584 (.A(\atari2600.tia.hmbl[3] ),
    .X(net5584));
 sg13g2_buf_4 fanout5585 (.X(net5585),
    .A(net7341));
 sg13g2_buf_4 fanout5586 (.X(net5586),
    .A(\atari2600.tia.hmm0[3] ));
 sg13g2_buf_4 fanout5587 (.X(net5587),
    .A(\atari2600.tia.hmp1[3] ));
 sg13g2_buf_4 fanout5588 (.X(net5588),
    .A(\atari2600.tia.hmp0[3] ));
 sg13g2_buf_4 fanout5589 (.X(net5589),
    .A(net7334));
 sg13g2_buf_2 fanout5590 (.A(net7353),
    .X(net5590));
 sg13g2_buf_1 fanout5591 (.A(\atari2600.tia.diag[60] ),
    .X(net5591));
 sg13g2_buf_4 fanout5592 (.X(net5592),
    .A(net7340));
 sg13g2_buf_4 fanout5593 (.X(net5593),
    .A(net7352));
 sg13g2_buf_2 fanout5594 (.A(\atari2600.tia.diag[68] ),
    .X(net5594));
 sg13g2_buf_4 fanout5595 (.X(net5595),
    .A(net7345));
 sg13g2_buf_4 fanout5596 (.X(net5596),
    .A(net7358));
 sg13g2_buf_2 fanout5597 (.A(net5598),
    .X(net5597));
 sg13g2_buf_2 fanout5598 (.A(net5599),
    .X(net5598));
 sg13g2_buf_2 fanout5599 (.A(\atari2600.tia.vid_out[6] ),
    .X(net5599));
 sg13g2_buf_4 fanout5600 (.X(net5600),
    .A(net5606));
 sg13g2_buf_4 fanout5601 (.X(net5601),
    .A(net5603));
 sg13g2_buf_1 fanout5602 (.A(net5603),
    .X(net5602));
 sg13g2_buf_4 fanout5603 (.X(net5603),
    .A(net5606));
 sg13g2_buf_2 fanout5604 (.A(net5605),
    .X(net5604));
 sg13g2_buf_4 fanout5605 (.X(net5605),
    .A(net5606));
 sg13g2_buf_2 fanout5606 (.A(\atari2600.tia.vid_out[6] ),
    .X(net5606));
 sg13g2_buf_4 fanout5607 (.X(net5607),
    .A(net5611));
 sg13g2_buf_2 fanout5608 (.A(net5611),
    .X(net5608));
 sg13g2_buf_4 fanout5609 (.X(net5609),
    .A(net5611));
 sg13g2_buf_1 fanout5610 (.A(net5611),
    .X(net5610));
 sg13g2_buf_1 fanout5611 (.A(net5625),
    .X(net5611));
 sg13g2_buf_2 fanout5612 (.A(net5615),
    .X(net5612));
 sg13g2_buf_2 fanout5613 (.A(net5615),
    .X(net5613));
 sg13g2_buf_4 fanout5614 (.X(net5614),
    .A(net5625));
 sg13g2_buf_2 fanout5615 (.A(net5625),
    .X(net5615));
 sg13g2_buf_4 fanout5616 (.X(net5616),
    .A(net5620));
 sg13g2_buf_2 fanout5617 (.A(net5620),
    .X(net5617));
 sg13g2_buf_4 fanout5618 (.X(net5618),
    .A(net5620));
 sg13g2_buf_1 fanout5619 (.A(net5620),
    .X(net5619));
 sg13g2_buf_2 fanout5620 (.A(net5625),
    .X(net5620));
 sg13g2_buf_2 fanout5621 (.A(net5623),
    .X(net5621));
 sg13g2_buf_4 fanout5622 (.X(net5622),
    .A(net5623));
 sg13g2_buf_4 fanout5623 (.X(net5623),
    .A(net5625));
 sg13g2_buf_1 fanout5624 (.A(net5625),
    .X(net5624));
 sg13g2_buf_4 fanout5625 (.X(net5625),
    .A(\atari2600.tia.vid_out[6] ));
 sg13g2_buf_2 fanout5626 (.A(net5633),
    .X(net5626));
 sg13g2_buf_1 fanout5627 (.A(net5633),
    .X(net5627));
 sg13g2_buf_4 fanout5628 (.X(net5628),
    .A(net5630));
 sg13g2_buf_1 fanout5629 (.A(net5630),
    .X(net5629));
 sg13g2_buf_2 fanout5630 (.A(net5633),
    .X(net5630));
 sg13g2_buf_2 fanout5631 (.A(net5633),
    .X(net5631));
 sg13g2_buf_1 fanout5632 (.A(net5633),
    .X(net5632));
 sg13g2_buf_4 fanout5633 (.X(net5633),
    .A(net5654));
 sg13g2_buf_4 fanout5634 (.X(net5634),
    .A(net5637));
 sg13g2_buf_1 fanout5635 (.A(net5637),
    .X(net5635));
 sg13g2_buf_4 fanout5636 (.X(net5636),
    .A(net5637));
 sg13g2_buf_2 fanout5637 (.A(net5654),
    .X(net5637));
 sg13g2_buf_4 fanout5638 (.X(net5638),
    .A(net5645));
 sg13g2_buf_2 fanout5639 (.A(net5645),
    .X(net5639));
 sg13g2_buf_2 fanout5640 (.A(net5641),
    .X(net5640));
 sg13g2_buf_4 fanout5641 (.X(net5641),
    .A(net5645));
 sg13g2_buf_2 fanout5642 (.A(net5644),
    .X(net5642));
 sg13g2_buf_4 fanout5643 (.X(net5643),
    .A(net5644));
 sg13g2_buf_4 fanout5644 (.X(net5644),
    .A(net5645));
 sg13g2_buf_4 fanout5645 (.X(net5645),
    .A(net5654));
 sg13g2_buf_2 fanout5646 (.A(net5647),
    .X(net5646));
 sg13g2_buf_1 fanout5647 (.A(net5653),
    .X(net5647));
 sg13g2_buf_2 fanout5648 (.A(net5653),
    .X(net5648));
 sg13g2_buf_1 fanout5649 (.A(net5653),
    .X(net5649));
 sg13g2_buf_2 fanout5650 (.A(net5651),
    .X(net5650));
 sg13g2_buf_2 fanout5651 (.A(net5652),
    .X(net5651));
 sg13g2_buf_4 fanout5652 (.X(net5652),
    .A(net5653));
 sg13g2_buf_4 fanout5653 (.X(net5653),
    .A(net5654));
 sg13g2_buf_8 fanout5654 (.A(\atari2600.tia.vid_out[5] ),
    .X(net5654));
 sg13g2_buf_2 fanout5655 (.A(net5656),
    .X(net5655));
 sg13g2_buf_4 fanout5656 (.X(net5656),
    .A(net5657));
 sg13g2_buf_2 fanout5657 (.A(net5683),
    .X(net5657));
 sg13g2_buf_4 fanout5658 (.X(net5658),
    .A(net5659));
 sg13g2_buf_4 fanout5659 (.X(net5659),
    .A(net5660));
 sg13g2_buf_2 fanout5660 (.A(net5664),
    .X(net5660));
 sg13g2_buf_4 fanout5661 (.X(net5661),
    .A(net5664));
 sg13g2_buf_2 fanout5662 (.A(net5664),
    .X(net5662));
 sg13g2_buf_1 fanout5663 (.A(net5664),
    .X(net5663));
 sg13g2_buf_2 fanout5664 (.A(net5683),
    .X(net5664));
 sg13g2_buf_4 fanout5665 (.X(net5665),
    .A(net5674));
 sg13g2_buf_2 fanout5666 (.A(net5674),
    .X(net5666));
 sg13g2_buf_2 fanout5667 (.A(net5668),
    .X(net5667));
 sg13g2_buf_2 fanout5668 (.A(net5669),
    .X(net5668));
 sg13g2_buf_2 fanout5669 (.A(net5674),
    .X(net5669));
 sg13g2_buf_2 fanout5670 (.A(net5671),
    .X(net5670));
 sg13g2_buf_2 fanout5671 (.A(net5672),
    .X(net5671));
 sg13g2_buf_4 fanout5672 (.X(net5672),
    .A(net5673));
 sg13g2_buf_2 fanout5673 (.A(net5674),
    .X(net5673));
 sg13g2_buf_2 fanout5674 (.A(net5682),
    .X(net5674));
 sg13g2_buf_2 fanout5675 (.A(net5679),
    .X(net5675));
 sg13g2_buf_2 fanout5676 (.A(net5679),
    .X(net5676));
 sg13g2_buf_4 fanout5677 (.X(net5677),
    .A(net5679));
 sg13g2_buf_2 fanout5678 (.A(net5679),
    .X(net5678));
 sg13g2_buf_4 fanout5679 (.X(net5679),
    .A(net5682));
 sg13g2_buf_4 fanout5680 (.X(net5680),
    .A(net5682));
 sg13g2_buf_4 fanout5681 (.X(net5681),
    .A(net5682));
 sg13g2_buf_4 fanout5682 (.X(net5682),
    .A(net5683));
 sg13g2_buf_2 fanout5683 (.A(\atari2600.tia.vid_out[4] ),
    .X(net5683));
 sg13g2_buf_2 fanout5684 (.A(net5685),
    .X(net5684));
 sg13g2_buf_2 fanout5685 (.A(net5712),
    .X(net5685));
 sg13g2_buf_4 fanout5686 (.X(net5686),
    .A(net5687));
 sg13g2_buf_2 fanout5687 (.A(net5712),
    .X(net5687));
 sg13g2_buf_4 fanout5688 (.X(net5688),
    .A(net5690));
 sg13g2_buf_4 fanout5689 (.X(net5689),
    .A(net5690));
 sg13g2_buf_4 fanout5690 (.X(net5690),
    .A(net5692));
 sg13g2_buf_2 fanout5691 (.A(net5692),
    .X(net5691));
 sg13g2_buf_2 fanout5692 (.A(net5712),
    .X(net5692));
 sg13g2_buf_4 fanout5693 (.X(net5693),
    .A(net5697));
 sg13g2_buf_2 fanout5694 (.A(net5697),
    .X(net5694));
 sg13g2_buf_2 fanout5695 (.A(net5697),
    .X(net5695));
 sg13g2_buf_1 fanout5696 (.A(net5697),
    .X(net5696));
 sg13g2_buf_4 fanout5697 (.X(net5697),
    .A(net5701));
 sg13g2_buf_4 fanout5698 (.X(net5698),
    .A(net5700));
 sg13g2_buf_1 fanout5699 (.A(net5700),
    .X(net5699));
 sg13g2_buf_2 fanout5700 (.A(net5701),
    .X(net5700));
 sg13g2_buf_2 fanout5701 (.A(net5712),
    .X(net5701));
 sg13g2_buf_2 fanout5702 (.A(net5704),
    .X(net5702));
 sg13g2_buf_2 fanout5703 (.A(net5704),
    .X(net5703));
 sg13g2_buf_4 fanout5704 (.X(net5704),
    .A(net5705));
 sg13g2_buf_4 fanout5705 (.X(net5705),
    .A(net5711));
 sg13g2_buf_2 fanout5706 (.A(net5711),
    .X(net5706));
 sg13g2_buf_2 fanout5707 (.A(net5711),
    .X(net5707));
 sg13g2_buf_2 fanout5708 (.A(net5709),
    .X(net5708));
 sg13g2_buf_2 fanout5709 (.A(net5710),
    .X(net5709));
 sg13g2_buf_2 fanout5710 (.A(net5711),
    .X(net5710));
 sg13g2_buf_2 fanout5711 (.A(net5712),
    .X(net5711));
 sg13g2_buf_8 fanout5712 (.A(\atari2600.tia.vid_out[3] ),
    .X(net5712));
 sg13g2_buf_2 fanout5713 (.A(net5741),
    .X(net5713));
 sg13g2_buf_2 fanout5714 (.A(net5741),
    .X(net5714));
 sg13g2_buf_4 fanout5715 (.X(net5715),
    .A(net5716));
 sg13g2_buf_4 fanout5716 (.X(net5716),
    .A(net5721));
 sg13g2_buf_4 fanout5717 (.X(net5717),
    .A(net5718));
 sg13g2_buf_4 fanout5718 (.X(net5718),
    .A(net5721));
 sg13g2_buf_4 fanout5719 (.X(net5719),
    .A(net5721));
 sg13g2_buf_2 fanout5720 (.A(net5721),
    .X(net5720));
 sg13g2_buf_2 fanout5721 (.A(net5741),
    .X(net5721));
 sg13g2_buf_4 fanout5722 (.X(net5722),
    .A(net5726));
 sg13g2_buf_2 fanout5723 (.A(net5726),
    .X(net5723));
 sg13g2_buf_4 fanout5724 (.X(net5724),
    .A(net5726));
 sg13g2_buf_2 fanout5725 (.A(net5726),
    .X(net5725));
 sg13g2_buf_2 fanout5726 (.A(net5729),
    .X(net5726));
 sg13g2_buf_2 fanout5727 (.A(net5728),
    .X(net5727));
 sg13g2_buf_2 fanout5728 (.A(net5729),
    .X(net5728));
 sg13g2_buf_4 fanout5729 (.X(net5729),
    .A(net5741));
 sg13g2_buf_2 fanout5730 (.A(net5734),
    .X(net5730));
 sg13g2_buf_1 fanout5731 (.A(net5734),
    .X(net5731));
 sg13g2_buf_4 fanout5732 (.X(net5732),
    .A(net5734));
 sg13g2_buf_1 fanout5733 (.A(net5734),
    .X(net5733));
 sg13g2_buf_2 fanout5734 (.A(net5740),
    .X(net5734));
 sg13g2_buf_2 fanout5735 (.A(net5737),
    .X(net5735));
 sg13g2_buf_4 fanout5736 (.X(net5736),
    .A(net5737));
 sg13g2_buf_2 fanout5737 (.A(net5740),
    .X(net5737));
 sg13g2_buf_4 fanout5738 (.X(net5738),
    .A(net5740));
 sg13g2_buf_1 fanout5739 (.A(net5740),
    .X(net5739));
 sg13g2_buf_4 fanout5740 (.X(net5740),
    .A(net5741));
 sg13g2_buf_8 fanout5741 (.A(\atari2600.tia.vid_out[2] ),
    .X(net5741));
 sg13g2_buf_2 fanout5742 (.A(net5744),
    .X(net5742));
 sg13g2_buf_2 fanout5743 (.A(net5744),
    .X(net5743));
 sg13g2_buf_4 fanout5744 (.X(net5744),
    .A(net5770));
 sg13g2_buf_4 fanout5745 (.X(net5745),
    .A(net5748));
 sg13g2_buf_2 fanout5746 (.A(net5748),
    .X(net5746));
 sg13g2_buf_4 fanout5747 (.X(net5747),
    .A(net5748));
 sg13g2_buf_2 fanout5748 (.A(net5770),
    .X(net5748));
 sg13g2_buf_2 fanout5749 (.A(net5750),
    .X(net5749));
 sg13g2_buf_4 fanout5750 (.X(net5750),
    .A(net5751));
 sg13g2_buf_2 fanout5751 (.A(net5770),
    .X(net5751));
 sg13g2_buf_4 fanout5752 (.X(net5752),
    .A(net5755));
 sg13g2_buf_4 fanout5753 (.X(net5753),
    .A(net5755));
 sg13g2_buf_2 fanout5754 (.A(net5755),
    .X(net5754));
 sg13g2_buf_4 fanout5755 (.X(net5755),
    .A(net5770));
 sg13g2_buf_2 fanout5756 (.A(net5760),
    .X(net5756));
 sg13g2_buf_2 fanout5757 (.A(net5760),
    .X(net5757));
 sg13g2_buf_4 fanout5758 (.X(net5758),
    .A(net5759));
 sg13g2_buf_2 fanout5759 (.A(net5760),
    .X(net5759));
 sg13g2_buf_2 fanout5760 (.A(net5770),
    .X(net5760));
 sg13g2_buf_2 fanout5761 (.A(net5765),
    .X(net5761));
 sg13g2_buf_1 fanout5762 (.A(net5765),
    .X(net5762));
 sg13g2_buf_2 fanout5763 (.A(net5765),
    .X(net5763));
 sg13g2_buf_1 fanout5764 (.A(net5765),
    .X(net5764));
 sg13g2_buf_4 fanout5765 (.X(net5765),
    .A(net5769));
 sg13g2_buf_4 fanout5766 (.X(net5766),
    .A(net5768));
 sg13g2_buf_2 fanout5767 (.A(net5768),
    .X(net5767));
 sg13g2_buf_4 fanout5768 (.X(net5768),
    .A(net5769));
 sg13g2_buf_4 fanout5769 (.X(net5769),
    .A(net5770));
 sg13g2_buf_8 fanout5770 (.A(\atari2600.tia.vid_out[1] ),
    .X(net5770));
 sg13g2_buf_2 fanout5771 (.A(net5780),
    .X(net5771));
 sg13g2_buf_2 fanout5772 (.A(net5780),
    .X(net5772));
 sg13g2_buf_4 fanout5773 (.X(net5773),
    .A(net5774));
 sg13g2_buf_2 fanout5774 (.A(net5775),
    .X(net5774));
 sg13g2_buf_4 fanout5775 (.X(net5775),
    .A(net5780));
 sg13g2_buf_2 fanout5776 (.A(net5778),
    .X(net5776));
 sg13g2_buf_1 fanout5777 (.A(net5778),
    .X(net5777));
 sg13g2_buf_4 fanout5778 (.X(net5778),
    .A(net5779));
 sg13g2_buf_2 fanout5779 (.A(net5780),
    .X(net5779));
 sg13g2_buf_2 fanout5780 (.A(\atari2600.tia.vid_out[0] ),
    .X(net5780));
 sg13g2_buf_2 fanout5781 (.A(net5783),
    .X(net5781));
 sg13g2_buf_1 fanout5782 (.A(net5783),
    .X(net5782));
 sg13g2_buf_4 fanout5783 (.X(net5783),
    .A(net5789));
 sg13g2_buf_4 fanout5784 (.X(net5784),
    .A(net5785));
 sg13g2_buf_4 fanout5785 (.X(net5785),
    .A(net5788));
 sg13g2_buf_2 fanout5786 (.A(net5788),
    .X(net5786));
 sg13g2_buf_2 fanout5787 (.A(net5788),
    .X(net5787));
 sg13g2_buf_2 fanout5788 (.A(net5789),
    .X(net5788));
 sg13g2_buf_2 fanout5789 (.A(\atari2600.tia.vid_out[0] ),
    .X(net5789));
 sg13g2_buf_2 fanout5790 (.A(net5791),
    .X(net5790));
 sg13g2_buf_4 fanout5791 (.X(net5791),
    .A(net5799));
 sg13g2_buf_4 fanout5792 (.X(net5792),
    .A(net5799));
 sg13g2_buf_2 fanout5793 (.A(net5799),
    .X(net5793));
 sg13g2_buf_4 fanout5794 (.X(net5794),
    .A(net5796));
 sg13g2_buf_2 fanout5795 (.A(net5796),
    .X(net5795));
 sg13g2_buf_2 fanout5796 (.A(net5799),
    .X(net5796));
 sg13g2_buf_4 fanout5797 (.X(net5797),
    .A(net5799));
 sg13g2_buf_1 fanout5798 (.A(net5799),
    .X(net5798));
 sg13g2_buf_4 fanout5799 (.X(net5799),
    .A(\atari2600.tia.vid_out[0] ));
 sg13g2_buf_4 fanout5800 (.X(net5800),
    .A(net5802));
 sg13g2_buf_4 fanout5801 (.X(net5801),
    .A(net5802));
 sg13g2_buf_4 fanout5802 (.X(net5802),
    .A(\atari2600.tia.vid_xpos[7] ));
 sg13g2_buf_4 fanout5803 (.X(net5803),
    .A(_00154_));
 sg13g2_buf_4 fanout5804 (.X(net5804),
    .A(\atari2600.tia.vid_xpos[6] ));
 sg13g2_buf_2 fanout5805 (.A(\atari2600.tia.vid_xpos[6] ),
    .X(net5805));
 sg13g2_buf_4 fanout5806 (.X(net5806),
    .A(net5808));
 sg13g2_buf_2 fanout5807 (.A(net5808),
    .X(net5807));
 sg13g2_buf_2 fanout5808 (.A(\atari2600.tia.vid_xpos[6] ),
    .X(net5808));
 sg13g2_buf_4 fanout5809 (.X(net5809),
    .A(_00153_));
 sg13g2_buf_4 fanout5810 (.X(net5810),
    .A(net5813));
 sg13g2_buf_4 fanout5811 (.X(net5811),
    .A(net5812));
 sg13g2_buf_4 fanout5812 (.X(net5812),
    .A(net5813));
 sg13g2_buf_4 fanout5813 (.X(net5813),
    .A(\atari2600.tia.vid_xpos[5] ));
 sg13g2_buf_4 fanout5814 (.X(net5814),
    .A(_00156_));
 sg13g2_buf_2 fanout5815 (.A(net7356),
    .X(net5815));
 sg13g2_buf_4 fanout5816 (.X(net5816),
    .A(net5817));
 sg13g2_buf_2 fanout5817 (.A(net5818),
    .X(net5817));
 sg13g2_buf_4 fanout5818 (.X(net5818),
    .A(\atari2600.tia.vid_xpos[4] ));
 sg13g2_buf_4 fanout5819 (.X(net5819),
    .A(_00152_));
 sg13g2_buf_4 fanout5820 (.X(net5820),
    .A(net5822));
 sg13g2_buf_2 fanout5821 (.A(net5822),
    .X(net5821));
 sg13g2_buf_4 fanout5822 (.X(net5822),
    .A(\atari2600.tia.vid_xpos[3] ));
 sg13g2_buf_8 fanout5823 (.A(\atari2600.tia.vid_xpos[2] ),
    .X(net5823));
 sg13g2_buf_2 fanout5824 (.A(\atari2600.tia.vid_xpos[2] ),
    .X(net5824));
 sg13g2_buf_2 fanout5825 (.A(net5828),
    .X(net5825));
 sg13g2_buf_4 fanout5826 (.X(net5826),
    .A(net5828));
 sg13g2_buf_2 fanout5827 (.A(net5828),
    .X(net5827));
 sg13g2_buf_2 fanout5828 (.A(\atari2600.tia.vid_xpos[1] ),
    .X(net5828));
 sg13g2_buf_4 fanout5829 (.X(net5829),
    .A(net5831));
 sg13g2_buf_4 fanout5830 (.X(net5830),
    .A(net5831));
 sg13g2_buf_4 fanout5831 (.X(net5831),
    .A(\atari2600.tia.vid_xpos[0] ));
 sg13g2_buf_2 fanout5832 (.A(net5833),
    .X(net5832));
 sg13g2_buf_2 fanout5833 (.A(net7306),
    .X(net5833));
 sg13g2_buf_2 fanout5834 (.A(net7266),
    .X(net5834));
 sg13g2_buf_2 fanout5835 (.A(net7313),
    .X(net5835));
 sg13g2_buf_2 fanout5836 (.A(\atari2600.tia.p1_scale[1] ),
    .X(net5836));
 sg13g2_buf_2 fanout5837 (.A(net7267),
    .X(net5837));
 sg13g2_buf_1 fanout5838 (.A(\atari2600.tia.p1_scale[0] ),
    .X(net5838));
 sg13g2_buf_4 fanout5839 (.X(net5839),
    .A(\hvsync_gen.hpos[9] ));
 sg13g2_buf_4 fanout5840 (.X(net5840),
    .A(net7323));
 sg13g2_buf_4 fanout5841 (.X(net5841),
    .A(\hvsync_gen.hpos[8] ));
 sg13g2_buf_4 fanout5842 (.X(net5842),
    .A(net5843));
 sg13g2_buf_4 fanout5843 (.X(net5843),
    .A(\hvsync_gen.hpos[7] ));
 sg13g2_buf_2 fanout5844 (.A(net5846),
    .X(net5844));
 sg13g2_buf_4 fanout5845 (.X(net5845),
    .A(net5846));
 sg13g2_buf_1 fanout5846 (.A(\hvsync_gen.hpos[6] ),
    .X(net5846));
 sg13g2_buf_4 fanout5847 (.X(net5847),
    .A(\hvsync_gen.hpos[6] ));
 sg13g2_buf_2 fanout5848 (.A(\hvsync_gen.hpos[6] ),
    .X(net5848));
 sg13g2_buf_4 fanout5849 (.X(net5849),
    .A(\hvsync_gen.hpos[5] ));
 sg13g2_buf_4 fanout5850 (.X(net5850),
    .A(net7326));
 sg13g2_buf_4 fanout5851 (.X(net5851),
    .A(net5852));
 sg13g2_buf_4 fanout5852 (.X(net5852),
    .A(net5856));
 sg13g2_buf_4 fanout5853 (.X(net5853),
    .A(net5855));
 sg13g2_buf_4 fanout5854 (.X(net5854),
    .A(net5855));
 sg13g2_buf_4 fanout5855 (.X(net5855),
    .A(net5856));
 sg13g2_buf_2 fanout5856 (.A(net5874),
    .X(net5856));
 sg13g2_buf_4 fanout5857 (.X(net5857),
    .A(net5861));
 sg13g2_buf_2 fanout5858 (.A(net5861),
    .X(net5858));
 sg13g2_buf_4 fanout5859 (.X(net5859),
    .A(net5861));
 sg13g2_buf_2 fanout5860 (.A(net5861),
    .X(net5860));
 sg13g2_buf_2 fanout5861 (.A(net5865),
    .X(net5861));
 sg13g2_buf_4 fanout5862 (.X(net5862),
    .A(net5865));
 sg13g2_buf_2 fanout5863 (.A(net5865),
    .X(net5863));
 sg13g2_buf_4 fanout5864 (.X(net5864),
    .A(net5865));
 sg13g2_buf_2 fanout5865 (.A(net5874),
    .X(net5865));
 sg13g2_buf_4 fanout5866 (.X(net5866),
    .A(net5868));
 sg13g2_buf_2 fanout5867 (.A(net5868),
    .X(net5867));
 sg13g2_buf_4 fanout5868 (.X(net5868),
    .A(net5869));
 sg13g2_buf_2 fanout5869 (.A(net5874),
    .X(net5869));
 sg13g2_buf_4 fanout5870 (.X(net5870),
    .A(net5872));
 sg13g2_buf_4 fanout5871 (.X(net5871),
    .A(net5873));
 sg13g2_buf_2 fanout5872 (.A(net5873),
    .X(net5872));
 sg13g2_buf_4 fanout5873 (.X(net5873),
    .A(net5874));
 sg13g2_buf_4 fanout5874 (.X(net5874),
    .A(\hvsync_gen.hpos[3] ));
 sg13g2_buf_4 fanout5875 (.X(net5875),
    .A(net5877));
 sg13g2_buf_4 fanout5876 (.X(net5876),
    .A(net5877));
 sg13g2_buf_2 fanout5877 (.A(net5881),
    .X(net5877));
 sg13g2_buf_4 fanout5878 (.X(net5878),
    .A(net5881));
 sg13g2_buf_2 fanout5879 (.A(net5881),
    .X(net5879));
 sg13g2_buf_4 fanout5880 (.X(net5880),
    .A(net5881));
 sg13g2_buf_1 fanout5881 (.A(net5906),
    .X(net5881));
 sg13g2_buf_4 fanout5882 (.X(net5882),
    .A(net5885));
 sg13g2_buf_4 fanout5883 (.X(net5883),
    .A(net5885));
 sg13g2_buf_2 fanout5884 (.A(net5885),
    .X(net5884));
 sg13g2_buf_2 fanout5885 (.A(net5906),
    .X(net5885));
 sg13g2_buf_4 fanout5886 (.X(net5886),
    .A(net5889));
 sg13g2_buf_4 fanout5887 (.X(net5887),
    .A(net5889));
 sg13g2_buf_2 fanout5888 (.A(net5889),
    .X(net5888));
 sg13g2_buf_2 fanout5889 (.A(net5906),
    .X(net5889));
 sg13g2_buf_4 fanout5890 (.X(net5890),
    .A(net5894));
 sg13g2_buf_2 fanout5891 (.A(net5894),
    .X(net5891));
 sg13g2_buf_4 fanout5892 (.X(net5892),
    .A(net5894));
 sg13g2_buf_2 fanout5893 (.A(net5894),
    .X(net5893));
 sg13g2_buf_2 fanout5894 (.A(net5905),
    .X(net5894));
 sg13g2_buf_4 fanout5895 (.X(net5895),
    .A(net5898));
 sg13g2_buf_4 fanout5896 (.X(net5896),
    .A(net5897));
 sg13g2_buf_4 fanout5897 (.X(net5897),
    .A(net5898));
 sg13g2_buf_2 fanout5898 (.A(net5905),
    .X(net5898));
 sg13g2_buf_4 fanout5899 (.X(net5899),
    .A(net5902));
 sg13g2_buf_4 fanout5900 (.X(net5900),
    .A(net5901));
 sg13g2_buf_4 fanout5901 (.X(net5901),
    .A(net5902));
 sg13g2_buf_2 fanout5902 (.A(net5905),
    .X(net5902));
 sg13g2_buf_4 fanout5903 (.X(net5903),
    .A(net5904));
 sg13g2_buf_4 fanout5904 (.X(net5904),
    .A(net5905));
 sg13g2_buf_4 fanout5905 (.X(net5905),
    .A(net5906));
 sg13g2_buf_4 fanout5906 (.X(net5906),
    .A(\hvsync_gen.hpos[3] ));
 sg13g2_buf_8 fanout5907 (.A(net5908),
    .X(net5907));
 sg13g2_buf_8 fanout5908 (.A(net5912),
    .X(net5908));
 sg13g2_buf_8 fanout5909 (.A(net5911),
    .X(net5909));
 sg13g2_buf_8 fanout5910 (.A(net5911),
    .X(net5910));
 sg13g2_buf_4 fanout5911 (.X(net5911),
    .A(net5912));
 sg13g2_buf_2 fanout5912 (.A(net5930),
    .X(net5912));
 sg13g2_buf_8 fanout5913 (.A(net5917),
    .X(net5913));
 sg13g2_buf_4 fanout5914 (.X(net5914),
    .A(net5917));
 sg13g2_buf_4 fanout5915 (.X(net5915),
    .A(net5917));
 sg13g2_buf_2 fanout5916 (.A(net5917),
    .X(net5916));
 sg13g2_buf_2 fanout5917 (.A(net5930),
    .X(net5917));
 sg13g2_buf_4 fanout5918 (.X(net5918),
    .A(net5921));
 sg13g2_buf_4 fanout5919 (.X(net5919),
    .A(net5921));
 sg13g2_buf_4 fanout5920 (.X(net5920),
    .A(net5921));
 sg13g2_buf_2 fanout5921 (.A(net5930),
    .X(net5921));
 sg13g2_buf_8 fanout5922 (.A(net5923),
    .X(net5922));
 sg13g2_buf_8 fanout5923 (.A(net5924),
    .X(net5923));
 sg13g2_buf_4 fanout5924 (.X(net5924),
    .A(net5930));
 sg13g2_buf_4 fanout5925 (.X(net5925),
    .A(net5928));
 sg13g2_buf_4 fanout5926 (.X(net5926),
    .A(net5927));
 sg13g2_buf_4 fanout5927 (.X(net5927),
    .A(net5928));
 sg13g2_buf_4 fanout5928 (.X(net5928),
    .A(net5929));
 sg13g2_buf_4 fanout5929 (.X(net5929),
    .A(net5930));
 sg13g2_buf_4 fanout5930 (.X(net5930),
    .A(net5968));
 sg13g2_buf_8 fanout5931 (.A(net5934),
    .X(net5931));
 sg13g2_buf_2 fanout5932 (.A(net5934),
    .X(net5932));
 sg13g2_buf_8 fanout5933 (.A(net5934),
    .X(net5933));
 sg13g2_buf_2 fanout5934 (.A(net5947),
    .X(net5934));
 sg13g2_buf_8 fanout5935 (.A(net5937),
    .X(net5935));
 sg13g2_buf_8 fanout5936 (.A(net5947),
    .X(net5936));
 sg13g2_buf_4 fanout5937 (.X(net5937),
    .A(net5947));
 sg13g2_buf_8 fanout5938 (.A(net5941),
    .X(net5938));
 sg13g2_buf_8 fanout5939 (.A(net5941),
    .X(net5939));
 sg13g2_buf_4 fanout5940 (.X(net5940),
    .A(net5941));
 sg13g2_buf_4 fanout5941 (.X(net5941),
    .A(net5947));
 sg13g2_buf_4 fanout5942 (.X(net5942),
    .A(net5946));
 sg13g2_buf_4 fanout5943 (.X(net5943),
    .A(net5946));
 sg13g2_buf_8 fanout5944 (.A(net5946),
    .X(net5944));
 sg13g2_buf_4 fanout5945 (.X(net5945),
    .A(net5946));
 sg13g2_buf_2 fanout5946 (.A(net5947),
    .X(net5946));
 sg13g2_buf_4 fanout5947 (.X(net5947),
    .A(net5968));
 sg13g2_buf_2 fanout5948 (.A(net5949),
    .X(net5948));
 sg13g2_buf_4 fanout5949 (.X(net5949),
    .A(net5950));
 sg13g2_buf_4 fanout5950 (.X(net5950),
    .A(net5958));
 sg13g2_buf_4 fanout5951 (.X(net5951),
    .A(net5958));
 sg13g2_buf_4 fanout5952 (.X(net5952),
    .A(net5958));
 sg13g2_buf_4 fanout5953 (.X(net5953),
    .A(net5958));
 sg13g2_buf_4 fanout5954 (.X(net5954),
    .A(net5958));
 sg13g2_buf_4 fanout5955 (.X(net5955),
    .A(net5957));
 sg13g2_buf_2 fanout5956 (.A(net5957),
    .X(net5956));
 sg13g2_buf_4 fanout5957 (.X(net5957),
    .A(net5958));
 sg13g2_buf_4 fanout5958 (.X(net5958),
    .A(net5968));
 sg13g2_buf_4 fanout5959 (.X(net5959),
    .A(net5960));
 sg13g2_buf_4 fanout5960 (.X(net5960),
    .A(net5967));
 sg13g2_buf_4 fanout5961 (.X(net5961),
    .A(net5967));
 sg13g2_buf_2 fanout5962 (.A(net5963),
    .X(net5962));
 sg13g2_buf_4 fanout5963 (.X(net5963),
    .A(net5967));
 sg13g2_buf_8 fanout5964 (.A(net5966),
    .X(net5964));
 sg13g2_buf_2 fanout5965 (.A(net5966),
    .X(net5965));
 sg13g2_buf_8 fanout5966 (.A(net5967),
    .X(net5966));
 sg13g2_buf_2 fanout5967 (.A(net5968),
    .X(net5967));
 sg13g2_buf_4 fanout5968 (.X(net5968),
    .A(\hvsync_gen.hpos[2] ));
 sg13g2_buf_2 fanout5969 (.A(net5970),
    .X(net5969));
 sg13g2_buf_4 fanout5970 (.X(net5970),
    .A(\atari2600.cpu.state[5] ));
 sg13g2_buf_2 fanout5971 (.A(\atari2600.cpu.state[4] ),
    .X(net5971));
 sg13g2_buf_1 fanout5972 (.A(\atari2600.cpu.state[4] ),
    .X(net5972));
 sg13g2_buf_4 fanout5973 (.X(net5973),
    .A(\atari2600.cpu.state[3] ));
 sg13g2_buf_2 fanout5974 (.A(\atari2600.cpu.state[1] ),
    .X(net5974));
 sg13g2_buf_2 fanout5975 (.A(\atari2600.cpu.state[0] ),
    .X(net5975));
 sg13g2_buf_2 fanout5976 (.A(net5977),
    .X(net5976));
 sg13g2_buf_2 fanout5977 (.A(net5978),
    .X(net5977));
 sg13g2_buf_2 fanout5978 (.A(net5979),
    .X(net5978));
 sg13g2_buf_2 fanout5979 (.A(net5981),
    .X(net5979));
 sg13g2_buf_4 fanout5980 (.X(net5980),
    .A(net5981));
 sg13g2_buf_2 fanout5981 (.A(net5982),
    .X(net5981));
 sg13g2_buf_4 fanout5982 (.X(net5982),
    .A(net5993));
 sg13g2_buf_4 fanout5983 (.X(net5983),
    .A(net5984));
 sg13g2_buf_4 fanout5984 (.X(net5984),
    .A(net5993));
 sg13g2_buf_2 fanout5985 (.A(net5986),
    .X(net5985));
 sg13g2_buf_2 fanout5986 (.A(net5987),
    .X(net5986));
 sg13g2_buf_2 fanout5987 (.A(net5988),
    .X(net5987));
 sg13g2_buf_2 fanout5988 (.A(net5989),
    .X(net5988));
 sg13g2_buf_2 fanout5989 (.A(net5993),
    .X(net5989));
 sg13g2_buf_2 fanout5990 (.A(net5992),
    .X(net5990));
 sg13g2_buf_4 fanout5991 (.X(net5991),
    .A(net5992));
 sg13g2_buf_4 fanout5992 (.X(net5992),
    .A(net5993));
 sg13g2_buf_8 fanout5993 (.A(_08097_),
    .X(net5993));
 sg13g2_buf_2 fanout5994 (.A(net6),
    .X(net5994));
 sg13g2_buf_2 fanout5995 (.A(ui_in[5]),
    .X(net5995));
 sg13g2_buf_2 fanout5996 (.A(ui_in[5]),
    .X(net5996));
 sg13g2_buf_4 fanout5997 (.X(net5997),
    .A(net5998));
 sg13g2_buf_2 fanout5998 (.A(net5999),
    .X(net5998));
 sg13g2_buf_4 fanout5999 (.X(net5999),
    .A(net6002));
 sg13g2_buf_4 fanout6000 (.X(net6000),
    .A(net6002));
 sg13g2_buf_2 fanout6001 (.A(net6002),
    .X(net6001));
 sg13g2_buf_2 fanout6002 (.A(net6039),
    .X(net6002));
 sg13g2_buf_2 fanout6003 (.A(net6005),
    .X(net6003));
 sg13g2_buf_2 fanout6004 (.A(net6005),
    .X(net6004));
 sg13g2_buf_2 fanout6005 (.A(net6015),
    .X(net6005));
 sg13g2_buf_2 fanout6006 (.A(net6008),
    .X(net6006));
 sg13g2_buf_2 fanout6007 (.A(net6008),
    .X(net6007));
 sg13g2_buf_4 fanout6008 (.X(net6008),
    .A(net6015));
 sg13g2_buf_4 fanout6009 (.X(net6009),
    .A(net6011));
 sg13g2_buf_2 fanout6010 (.A(net6015),
    .X(net6010));
 sg13g2_buf_1 fanout6011 (.A(net6015),
    .X(net6011));
 sg13g2_buf_2 fanout6012 (.A(net6014),
    .X(net6012));
 sg13g2_buf_2 fanout6013 (.A(net6014),
    .X(net6013));
 sg13g2_buf_2 fanout6014 (.A(net6015),
    .X(net6014));
 sg13g2_buf_4 fanout6015 (.X(net6015),
    .A(net6016));
 sg13g2_buf_4 fanout6016 (.X(net6016),
    .A(net6039));
 sg13g2_buf_4 fanout6017 (.X(net6017),
    .A(net6018));
 sg13g2_buf_2 fanout6018 (.A(net6026),
    .X(net6018));
 sg13g2_buf_2 fanout6019 (.A(net6021),
    .X(net6019));
 sg13g2_buf_1 fanout6020 (.A(net6021),
    .X(net6020));
 sg13g2_buf_2 fanout6021 (.A(net6026),
    .X(net6021));
 sg13g2_buf_2 fanout6022 (.A(net6023),
    .X(net6022));
 sg13g2_buf_2 fanout6023 (.A(net6025),
    .X(net6023));
 sg13g2_buf_2 fanout6024 (.A(net6025),
    .X(net6024));
 sg13g2_buf_1 fanout6025 (.A(net6026),
    .X(net6025));
 sg13g2_buf_2 fanout6026 (.A(net6039),
    .X(net6026));
 sg13g2_buf_2 fanout6027 (.A(net6028),
    .X(net6027));
 sg13g2_buf_2 fanout6028 (.A(net6029),
    .X(net6028));
 sg13g2_buf_2 fanout6029 (.A(net6031),
    .X(net6029));
 sg13g2_buf_2 fanout6030 (.A(net6031),
    .X(net6030));
 sg13g2_buf_2 fanout6031 (.A(net6038),
    .X(net6031));
 sg13g2_buf_4 fanout6032 (.X(net6032),
    .A(net6033));
 sg13g2_buf_2 fanout6033 (.A(net6038),
    .X(net6033));
 sg13g2_buf_2 fanout6034 (.A(net6035),
    .X(net6034));
 sg13g2_buf_2 fanout6035 (.A(net6038),
    .X(net6035));
 sg13g2_buf_4 fanout6036 (.X(net6036),
    .A(net6037));
 sg13g2_buf_4 fanout6037 (.X(net6037),
    .A(net6038));
 sg13g2_buf_4 fanout6038 (.X(net6038),
    .A(net6039));
 sg13g2_buf_8 fanout6039 (.A(rst_n),
    .X(net6039));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[6]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[1]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[4]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[5]),
    .X(net11));
 sg13g2_tiehi _28843__12 (.L_HI(net12));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_72_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_74_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_2 clkbuf_leaf_75_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_2 clkbuf_leaf_76_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_2 clkbuf_leaf_77_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_2 clkbuf_leaf_78_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_2 clkbuf_leaf_79_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_2 clkbuf_leaf_80_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_2 clkbuf_leaf_81_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_2 clkbuf_leaf_82_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_2 clkbuf_leaf_83_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_2 clkbuf_leaf_84_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_2 clkbuf_leaf_85_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_2 clkbuf_leaf_86_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_2 clkbuf_leaf_87_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_2 clkbuf_leaf_88_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_2 clkbuf_leaf_89_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_2 clkbuf_leaf_90_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_2 clkbuf_leaf_91_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_2 clkbuf_leaf_92_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_2 clkbuf_leaf_93_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_2 clkbuf_leaf_94_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_2 clkbuf_leaf_95_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_2 clkbuf_leaf_96_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_2 clkbuf_leaf_97_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_2 clkbuf_leaf_98_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_2 clkbuf_leaf_99_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_2 clkbuf_leaf_100_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_2 clkbuf_leaf_101_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_2 clkbuf_leaf_102_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_2 clkbuf_leaf_103_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_2 clkbuf_leaf_104_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_2 clkbuf_leaf_105_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_2 clkbuf_leaf_106_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_2 clkbuf_leaf_107_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_2 clkbuf_leaf_108_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_2 clkbuf_leaf_109_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_2 clkbuf_leaf_110_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_2 clkbuf_leaf_111_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_2 clkbuf_leaf_112_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_2 clkbuf_leaf_113_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_2 clkbuf_leaf_114_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_2 clkbuf_leaf_115_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_2 clkbuf_leaf_116_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_2 clkbuf_leaf_117_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_2 clkbuf_leaf_118_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_2 clkbuf_leaf_119_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_2 clkbuf_leaf_120_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_2 clkbuf_leaf_121_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_2 clkbuf_leaf_122_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_2 clkbuf_leaf_123_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_2 clkbuf_leaf_124_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_2 clkbuf_leaf_125_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_2 clkbuf_leaf_126_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_2 clkbuf_leaf_127_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_2 clkbuf_leaf_128_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_2 clkbuf_leaf_129_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_2 clkbuf_leaf_130_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_2 clkbuf_leaf_131_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_2 clkbuf_leaf_132_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_2 clkbuf_leaf_133_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_2 clkbuf_leaf_134_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_2 clkbuf_leaf_135_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_2 clkbuf_leaf_136_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_2 clkbuf_leaf_137_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_2 clkbuf_leaf_138_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_2 clkbuf_leaf_139_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_2 clkbuf_leaf_140_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_2 clkbuf_leaf_141_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_2 clkbuf_leaf_142_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_2 clkbuf_leaf_143_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_2 clkbuf_leaf_144_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_2 clkbuf_leaf_145_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_2 clkbuf_leaf_146_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_2 clkbuf_leaf_147_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_2 clkbuf_leaf_148_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_2 clkbuf_leaf_149_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_2 clkbuf_leaf_150_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_2 clkbuf_leaf_151_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_2 clkbuf_leaf_152_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_2 clkbuf_leaf_153_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_2 clkbuf_leaf_154_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_2 clkbuf_leaf_155_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_2 clkbuf_leaf_156_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_2 clkbuf_leaf_158_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_2 clkbuf_leaf_159_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_2 clkbuf_leaf_160_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_2 clkbuf_leaf_161_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_2 clkbuf_leaf_162_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_2 clkbuf_leaf_163_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_2 clkbuf_leaf_164_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_2 clkbuf_leaf_165_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_2 clkbuf_leaf_166_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_2 clkbuf_leaf_167_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_2 clkbuf_leaf_168_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_2 clkbuf_leaf_169_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_2 clkbuf_leaf_170_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_2 clkbuf_leaf_171_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_2 clkbuf_leaf_172_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_2 clkbuf_leaf_173_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_2 clkbuf_leaf_174_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_2 clkbuf_leaf_175_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_2 clkbuf_leaf_176_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_2 clkbuf_leaf_177_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_2 clkbuf_leaf_178_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_2 clkbuf_leaf_179_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_2 clkbuf_leaf_180_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_2 clkbuf_leaf_181_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_2 clkbuf_leaf_182_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_2 clkbuf_leaf_183_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_2 clkbuf_leaf_184_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_2 clkbuf_leaf_185_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_2 clkbuf_leaf_186_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_2 clkbuf_leaf_187_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_2 clkbuf_leaf_188_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_2 clkbuf_leaf_189_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_2 clkbuf_leaf_190_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_2 clkbuf_leaf_191_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_2 clkbuf_leaf_192_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_2 clkbuf_leaf_193_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_2 clkbuf_leaf_194_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_2 clkbuf_leaf_195_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_2 clkbuf_leaf_196_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_2 clkbuf_leaf_197_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_2 clkbuf_leaf_198_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_2 clkbuf_leaf_199_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_2 clkbuf_leaf_200_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_2 clkbuf_leaf_201_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_2 clkbuf_leaf_202_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_2 clkbuf_leaf_203_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_2 clkbuf_leaf_204_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_2 clkbuf_leaf_205_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_2 clkbuf_leaf_206_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_2 clkbuf_leaf_207_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_2 clkbuf_leaf_208_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_2 clkbuf_leaf_209_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_2 clkbuf_leaf_210_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_2 clkbuf_leaf_211_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_2 clkbuf_leaf_212_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_2 clkbuf_leaf_213_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_2 clkbuf_leaf_214_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_2 clkbuf_leaf_215_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_2 clkbuf_leaf_216_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_2 clkbuf_leaf_217_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_2 clkbuf_leaf_218_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_2 clkbuf_leaf_219_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_2 clkbuf_leaf_220_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_2 clkbuf_leaf_221_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_2 clkbuf_leaf_222_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_2 clkbuf_leaf_223_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_2 clkbuf_leaf_224_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_2 clkbuf_leaf_225_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_2 clkbuf_leaf_226_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_2 clkbuf_leaf_227_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_2 clkbuf_leaf_228_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_2 clkbuf_leaf_229_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_2 clkbuf_leaf_230_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_2 clkbuf_leaf_231_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_2 clkbuf_leaf_232_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_2 clkbuf_leaf_233_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_2 clkbuf_leaf_234_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_2 clkbuf_leaf_235_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_2 clkbuf_leaf_236_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_2 clkbuf_leaf_237_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_2 clkbuf_leaf_238_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_2 clkbuf_leaf_239_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_2 clkbuf_leaf_240_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_2 clkbuf_leaf_241_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_2 clkbuf_leaf_242_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_2 clkbuf_leaf_243_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_2 clkbuf_leaf_244_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_2 clkbuf_leaf_245_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_2 clkbuf_leaf_246_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_2 clkbuf_leaf_247_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_2 clkbuf_leaf_248_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_2 clkbuf_leaf_249_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_2 clkbuf_leaf_250_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_2 clkbuf_leaf_251_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_2 clkbuf_leaf_252_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_2 clkbuf_leaf_253_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_2 clkbuf_leaf_254_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_2 clkbuf_leaf_255_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_2 clkbuf_leaf_256_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_2 clkbuf_leaf_257_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_2 clkbuf_leaf_258_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_2 clkbuf_leaf_259_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_2 clkbuf_leaf_260_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_2 clkbuf_leaf_261_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_2 clkbuf_leaf_262_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_2 clkbuf_leaf_263_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_2 clkbuf_leaf_264_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_2 clkbuf_leaf_265_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_2 clkbuf_leaf_266_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_2 clkbuf_leaf_267_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_2 clkbuf_leaf_268_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_2 clkbuf_leaf_269_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_2 clkbuf_leaf_270_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_2 clkbuf_leaf_271_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_2 clkbuf_leaf_272_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_2 clkbuf_leaf_273_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_2 clkbuf_leaf_274_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_2 clkbuf_leaf_275_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_2 clkbuf_leaf_276_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_2 clkbuf_leaf_277_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_2 clkbuf_leaf_278_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_2 clkbuf_leaf_279_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_2 clkbuf_leaf_280_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_2 clkbuf_leaf_281_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_2 clkbuf_leaf_282_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_2 clkbuf_leaf_283_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_2 clkbuf_leaf_284_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_2 clkbuf_leaf_285_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_2 clkbuf_leaf_286_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_2 clkbuf_leaf_287_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_2 clkbuf_leaf_288_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_2 clkbuf_leaf_289_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_2 clkbuf_leaf_290_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_2 clkbuf_leaf_291_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_2 clkbuf_leaf_292_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_2 clkbuf_leaf_293_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_2 clkbuf_leaf_294_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_2 clkbuf_leaf_295_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_2 clkbuf_leaf_296_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_2 clkbuf_leaf_297_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_2 clkbuf_leaf_298_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_2 clkbuf_leaf_299_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_2 clkbuf_leaf_300_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_2 clkbuf_leaf_301_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_2 clkbuf_leaf_302_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_2 clkbuf_leaf_303_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_2 clkbuf_leaf_304_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_2 clkbuf_leaf_305_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_2 clkbuf_leaf_306_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_2 clkbuf_leaf_307_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_2 clkbuf_leaf_308_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_2 clkbuf_leaf_309_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_2 clkbuf_leaf_310_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_2 clkbuf_leaf_311_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_311_clk));
 sg13g2_buf_2 clkbuf_leaf_312_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_312_clk));
 sg13g2_buf_2 clkbuf_leaf_313_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_313_clk));
 sg13g2_buf_2 clkbuf_leaf_314_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_314_clk));
 sg13g2_buf_2 clkbuf_leaf_315_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_315_clk));
 sg13g2_buf_2 clkbuf_leaf_316_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_316_clk));
 sg13g2_buf_2 clkbuf_leaf_317_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_317_clk));
 sg13g2_buf_2 clkbuf_leaf_318_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_318_clk));
 sg13g2_buf_2 clkbuf_leaf_319_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_319_clk));
 sg13g2_buf_2 clkbuf_leaf_320_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_320_clk));
 sg13g2_buf_2 clkbuf_leaf_321_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_321_clk));
 sg13g2_buf_2 clkbuf_leaf_322_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_322_clk));
 sg13g2_buf_2 clkbuf_leaf_323_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_323_clk));
 sg13g2_buf_2 clkbuf_leaf_324_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_324_clk));
 sg13g2_buf_2 clkbuf_leaf_325_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_325_clk));
 sg13g2_buf_2 clkbuf_leaf_326_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_326_clk));
 sg13g2_buf_2 clkbuf_leaf_327_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_327_clk));
 sg13g2_buf_2 clkbuf_leaf_328_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_328_clk));
 sg13g2_buf_2 clkbuf_leaf_329_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_329_clk));
 sg13g2_buf_2 clkbuf_leaf_330_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_330_clk));
 sg13g2_buf_2 clkbuf_leaf_331_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_331_clk));
 sg13g2_buf_2 clkbuf_leaf_332_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_332_clk));
 sg13g2_buf_2 clkbuf_leaf_333_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_333_clk));
 sg13g2_buf_2 clkbuf_leaf_334_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_334_clk));
 sg13g2_buf_2 clkbuf_leaf_335_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_335_clk));
 sg13g2_buf_2 clkbuf_leaf_336_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_336_clk));
 sg13g2_buf_2 clkbuf_leaf_337_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_337_clk));
 sg13g2_buf_2 clkbuf_leaf_338_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_338_clk));
 sg13g2_buf_2 clkbuf_leaf_339_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_339_clk));
 sg13g2_buf_2 clkbuf_leaf_340_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_340_clk));
 sg13g2_buf_2 clkbuf_leaf_341_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_341_clk));
 sg13g2_buf_2 clkbuf_leaf_342_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_342_clk));
 sg13g2_buf_2 clkbuf_leaf_343_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_343_clk));
 sg13g2_buf_2 clkbuf_leaf_344_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_344_clk));
 sg13g2_buf_2 clkbuf_leaf_345_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_345_clk));
 sg13g2_buf_2 clkbuf_leaf_346_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_346_clk));
 sg13g2_buf_2 clkbuf_leaf_347_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_347_clk));
 sg13g2_buf_2 clkbuf_leaf_348_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_348_clk));
 sg13g2_buf_2 clkbuf_leaf_349_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_349_clk));
 sg13g2_buf_2 clkbuf_leaf_350_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_350_clk));
 sg13g2_buf_2 clkbuf_leaf_351_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_351_clk));
 sg13g2_buf_2 clkbuf_leaf_352_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_352_clk));
 sg13g2_buf_2 clkbuf_leaf_353_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_353_clk));
 sg13g2_buf_2 clkbuf_leaf_354_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_354_clk));
 sg13g2_buf_2 clkbuf_leaf_355_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_355_clk));
 sg13g2_buf_2 clkbuf_leaf_356_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_356_clk));
 sg13g2_buf_2 clkbuf_leaf_357_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_357_clk));
 sg13g2_buf_2 clkbuf_leaf_358_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_358_clk));
 sg13g2_buf_2 clkbuf_leaf_359_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_359_clk));
 sg13g2_buf_2 clkbuf_leaf_360_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_360_clk));
 sg13g2_buf_2 clkbuf_leaf_361_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_361_clk));
 sg13g2_buf_2 clkbuf_leaf_362_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_362_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_2 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_2 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_2 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_2 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_2 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_2 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_2 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_2 clkbuf_6_0__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_0__leaf_clk));
 sg13g2_buf_2 clkbuf_6_1__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_1__leaf_clk));
 sg13g2_buf_2 clkbuf_6_2__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_2__leaf_clk));
 sg13g2_buf_2 clkbuf_6_3__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_3__leaf_clk));
 sg13g2_buf_2 clkbuf_6_4__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_4__leaf_clk));
 sg13g2_buf_2 clkbuf_6_5__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_5__leaf_clk));
 sg13g2_buf_2 clkbuf_6_6__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_6__leaf_clk));
 sg13g2_buf_2 clkbuf_6_7__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_7__leaf_clk));
 sg13g2_buf_2 clkbuf_6_8__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_8__leaf_clk));
 sg13g2_buf_2 clkbuf_6_9__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_9__leaf_clk));
 sg13g2_buf_2 clkbuf_6_10__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_10__leaf_clk));
 sg13g2_buf_2 clkbuf_6_11__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_11__leaf_clk));
 sg13g2_buf_2 clkbuf_6_12__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_12__leaf_clk));
 sg13g2_buf_2 clkbuf_6_13__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_13__leaf_clk));
 sg13g2_buf_2 clkbuf_6_14__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_14__leaf_clk));
 sg13g2_buf_2 clkbuf_6_15__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_15__leaf_clk));
 sg13g2_buf_2 clkbuf_6_16__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_16__leaf_clk));
 sg13g2_buf_2 clkbuf_6_17__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_17__leaf_clk));
 sg13g2_buf_2 clkbuf_6_18__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_18__leaf_clk));
 sg13g2_buf_2 clkbuf_6_19__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_19__leaf_clk));
 sg13g2_buf_2 clkbuf_6_20__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_20__leaf_clk));
 sg13g2_buf_2 clkbuf_6_21__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_21__leaf_clk));
 sg13g2_buf_2 clkbuf_6_22__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_22__leaf_clk));
 sg13g2_buf_2 clkbuf_6_23__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_23__leaf_clk));
 sg13g2_buf_2 clkbuf_6_24__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_24__leaf_clk));
 sg13g2_buf_2 clkbuf_6_25__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_25__leaf_clk));
 sg13g2_buf_2 clkbuf_6_26__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_26__leaf_clk));
 sg13g2_buf_2 clkbuf_6_27__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_27__leaf_clk));
 sg13g2_buf_2 clkbuf_6_28__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_28__leaf_clk));
 sg13g2_buf_2 clkbuf_6_29__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_29__leaf_clk));
 sg13g2_buf_2 clkbuf_6_30__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_30__leaf_clk));
 sg13g2_buf_2 clkbuf_6_31__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_31__leaf_clk));
 sg13g2_buf_2 clkbuf_6_32__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_32__leaf_clk));
 sg13g2_buf_2 clkbuf_6_33__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_33__leaf_clk));
 sg13g2_buf_2 clkbuf_6_34__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_34__leaf_clk));
 sg13g2_buf_2 clkbuf_6_35__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_35__leaf_clk));
 sg13g2_buf_2 clkbuf_6_36__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_36__leaf_clk));
 sg13g2_buf_2 clkbuf_6_37__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_37__leaf_clk));
 sg13g2_buf_2 clkbuf_6_38__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_38__leaf_clk));
 sg13g2_buf_2 clkbuf_6_39__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_39__leaf_clk));
 sg13g2_buf_2 clkbuf_6_40__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_40__leaf_clk));
 sg13g2_buf_2 clkbuf_6_41__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_41__leaf_clk));
 sg13g2_buf_2 clkbuf_6_42__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_42__leaf_clk));
 sg13g2_buf_2 clkbuf_6_43__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_43__leaf_clk));
 sg13g2_buf_2 clkbuf_6_44__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_44__leaf_clk));
 sg13g2_buf_2 clkbuf_6_45__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_45__leaf_clk));
 sg13g2_buf_2 clkbuf_6_46__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_46__leaf_clk));
 sg13g2_buf_2 clkbuf_6_47__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_47__leaf_clk));
 sg13g2_buf_2 clkbuf_6_48__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_48__leaf_clk));
 sg13g2_buf_2 clkbuf_6_49__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_49__leaf_clk));
 sg13g2_buf_2 clkbuf_6_50__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_50__leaf_clk));
 sg13g2_buf_2 clkbuf_6_51__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_51__leaf_clk));
 sg13g2_buf_2 clkbuf_6_52__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_52__leaf_clk));
 sg13g2_buf_2 clkbuf_6_53__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_53__leaf_clk));
 sg13g2_buf_2 clkbuf_6_54__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_54__leaf_clk));
 sg13g2_buf_2 clkbuf_6_55__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_55__leaf_clk));
 sg13g2_buf_2 clkbuf_6_56__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_56__leaf_clk));
 sg13g2_buf_2 clkbuf_6_57__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_57__leaf_clk));
 sg13g2_buf_2 clkbuf_6_58__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_58__leaf_clk));
 sg13g2_buf_2 clkbuf_6_59__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_59__leaf_clk));
 sg13g2_buf_2 clkbuf_6_60__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_60__leaf_clk));
 sg13g2_buf_2 clkbuf_6_61__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_61__leaf_clk));
 sg13g2_buf_2 clkbuf_6_62__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_62__leaf_clk));
 sg13g2_buf_2 clkbuf_6_63__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_63__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_6_3__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_6_7__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_6_11__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_6_13__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_6_19__leaf_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_2 clkload7 (.A(clknet_6_27__leaf_clk));
 sg13g2_buf_2 clkload8 (.A(clknet_6_29__leaf_clk));
 sg13g2_buf_2 clkload9 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_2 clkload10 (.A(clknet_6_35__leaf_clk));
 sg13g2_buf_2 clkload11 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_2 clkload12 (.A(clknet_6_43__leaf_clk));
 sg13g2_buf_2 clkload13 (.A(clknet_6_45__leaf_clk));
 sg13g2_buf_2 clkload14 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_2 clkload15 (.A(clknet_6_51__leaf_clk));
 sg13g2_buf_2 clkload16 (.A(clknet_6_53__leaf_clk));
 sg13g2_buf_1 clkload17 (.A(clknet_6_55__leaf_clk));
 sg13g2_buf_2 clkload18 (.A(clknet_6_59__leaf_clk));
 sg13g2_buf_2 clkload19 (.A(clknet_6_61__leaf_clk));
 sg13g2_buf_2 clkload20 (.A(clknet_6_63__leaf_clk));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_362_clk));
 sg13g2_inv_8 clkload22 (.A(clknet_leaf_15_clk));
 sg13g2_inv_4 clkload23 (.A(clknet_leaf_16_clk));
 sg13g2_inv_4 clkload24 (.A(clknet_leaf_149_clk));
 sg13g2_inv_1 clkload25 (.A(clknet_leaf_150_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_00171_),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold2 (.A(\flash_rom.data_ready ),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold3 (.A(_00170_),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold4 (.A(_07619_),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold5 (.A(_00169_),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold6 (.A(_01201_),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold7 (.A(_00048_),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold8 (.A(\atari2600.clk_counter[6] ),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold9 (.A(\flash_rom.fsm_state[0] ),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold10 (.A(\flash_rom.spi_select ),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold11 (.A(\r_pwm_odd[2] ),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold12 (.A(\atari2600.clk_counter[7] ),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold13 (.A(_00168_),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold14 (.A(_06340_),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold15 (.A(_02028_),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold16 (.A(\atari2600.ram[37][4] ),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold17 (.A(\atari2600.clk_counter[3] ),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold18 (.A(_00049_),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold19 (.A(\atari2600.ram[53][4] ),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold20 (.A(\g_pwm_odd[2] ),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold21 (.A(\flash_rom.addr[1] ),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold22 (.A(\atari2600.ram[51][4] ),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold23 (.A(\atari2600.clk_counter[2] ),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold24 (.A(\atari2600.ram[4][4] ),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold25 (.A(\atari2600.ram[60][4] ),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold26 (.A(\atari2600.ram[124][4] ),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold27 (.A(\atari2600.ram[41][4] ),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold28 (.A(\atari2600.tia.cx[2] ),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold29 (.A(\atari2600.ram[57][4] ),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold30 (.A(\flash_rom.addr[3] ),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold31 (.A(\atari2600.ram[52][4] ),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold32 (.A(\atari2600.ram[64][4] ),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold33 (.A(\atari2600.cpu.cld ),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold34 (.A(\atari2600.tia.p1_scale[1] ),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold35 (.A(\flash_rom.addr[2] ),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold36 (.A(\atari2600.ram[68][4] ),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold37 (.A(\atari2600.clk_counter[4] ),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold38 (.A(\atari2600.ram[35][4] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold39 (.A(\atari2600.tia.cx[7] ),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold40 (.A(_00053_),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold41 (.A(_00045_),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold42 (.A(\atari2600.ram[125][4] ),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold43 (.A(\atari2600.tia.cx[6] ),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold44 (.A(\atari2600.tia.old_grp1[7] ),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold45 (.A(_01827_),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold46 (.A(\atari2600.tia.audv0[0] ),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold47 (.A(\atari2600.ram[16][4] ),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold48 (.A(\atari2600.clk_counter[5] ),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold49 (.A(\atari2600.ram[5][4] ),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold50 (.A(\atari2600.tia.old_grp1[2] ),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold51 (.A(_01822_),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold52 (.A(\atari2600.ram[25][4] ),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold53 (.A(\atari2600.ram[65][4] ),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold54 (.A(\atari2600.ram[61][4] ),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold55 (.A(\atari2600.ram[36][4] ),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold56 (.A(\atari2600.ram[40][4] ),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold57 (.A(\atari2600.tia.old_grp1[0] ),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold58 (.A(_01820_),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold59 (.A(\atari2600.ram[20][4] ),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold60 (.A(\atari2600.tia.audf0[4] ),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold61 (.A(\atari2600.ram[33][4] ),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold62 (.A(\atari2600.ram[67][4] ),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold63 (.A(\atari2600.tia.cx[14] ),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold64 (.A(_10250_),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold65 (.A(\atari2600.ram[55][4] ),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold66 (.A(\atari2600.tia.dat_o[6] ),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold67 (.A(_02994_),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold68 (.A(\atari2600.tia.p1_copies[2] ),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold69 (.A(\atari2600.ram[17][4] ),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold70 (.A(\atari2600.ram[63][4] ),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold71 (.A(\atari2600.ram[56][4] ),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold72 (.A(\atari2600.tia.cx[5] ),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold73 (.A(\atari2600.tia.cx_clr ),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold74 (.A(\atari2600.tia.old_grp1[6] ),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold75 (.A(_01826_),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold76 (.A(\atari2600.cpu.sed ),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold77 (.A(\flash_rom.addr[0] ),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold78 (.A(\atari2600.ram[76][7] ),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold79 (.A(\scanline[124][1] ),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold80 (.A(\atari2600.tia.audio_left_counter[15] ),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold81 (.A(_05954_),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold82 (.A(\atari2600.tia.dat_o[7] ),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold83 (.A(\atari2600.ram[73][1] ),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold84 (.A(\atari2600.tia.audio_left_counter[14] ),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold85 (.A(_02026_),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold86 (.A(\atari2600.tia.cx[8] ),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold87 (.A(\atari2600.ram[73][0] ),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold88 (.A(\atari2600.tia.diag[77] ),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold89 (.A(\atari2600.ram[15][4] ),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold90 (.A(\atari2600.ram[89][4] ),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold91 (.A(\atari2600.tia.p0_copies[2] ),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold92 (.A(\atari2600.ram[92][7] ),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold93 (.A(\atari2600.cpu.cli ),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold94 (.A(\atari2600.ram[93][4] ),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold95 (.A(\atari2600.tia.cx[4] ),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold96 (.A(\atari2600.ram[72][2] ),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold97 (.A(\atari2600.ram[1][1] ),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold98 (.A(\atari2600.tia.audv0[2] ),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold99 (.A(\atari2600.tia.old_grp1[1] ),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold100 (.A(_01821_),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold101 (.A(\atari2600.tia.cx[13] ),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold102 (.A(\atari2600.tia.audv0[1] ),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold103 (.A(\atari2600.tia.diag[79] ),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold104 (.A(\atari2600.ram[30][5] ),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold105 (.A(\atari2600.input_joystick_0[2] ),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold106 (.A(_01213_),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold107 (.A(\atari2600.ram[78][6] ),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold108 (.A(\atari2600.ram[89][2] ),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold109 (.A(\atari2600.ram[88][1] ),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold110 (.A(\atari2600.tia.audio_right_counter[15] ),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold111 (.A(\atari2600.rom_data[5] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold112 (.A(_02925_),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold113 (.A(\atari2600.ram[74][0] ),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold114 (.A(\atari2600.ram[94][1] ),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold115 (.A(\atari2600.ram[72][1] ),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold116 (.A(\atari2600.ram[3][2] ),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold117 (.A(\atari2600.ram[38][1] ),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold118 (.A(\atari2600.ram[78][4] ),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold119 (.A(\atari2600.ram[93][0] ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold120 (.A(\atari2600.ram[72][7] ),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold121 (.A(\atari2600.ram[54][2] ),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold122 (.A(\atari2600.ram[93][3] ),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold123 (.A(\atari2600.ram[89][5] ),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold124 (.A(\atari2600.tia.cx[1] ),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold125 (.A(\atari2600.ram[1][7] ),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold126 (.A(\atari2600.ram[106][3] ),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold127 (.A(\atari2600.ram[102][0] ),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold128 (.A(\atari2600.ram[92][6] ),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold129 (.A(\atari2600.ram[92][2] ),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold130 (.A(\atari2600.ram[90][3] ),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold131 (.A(\flash_rom.addr[9] ),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold132 (.A(_01921_),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold133 (.A(\atari2600.ram[91][0] ),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold134 (.A(\atari2600.ram[79][0] ),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold135 (.A(\atari2600.tia.cx[9] ),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold136 (.A(\atari2600.ram[92][3] ),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold137 (.A(\atari2600.ram[66][7] ),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold138 (.A(\atari2600.cpu.sei ),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold139 (.A(\atari2600.ram[10][3] ),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold140 (.A(\atari2600.ram[58][7] ),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold141 (.A(\atari2600.ram[73][4] ),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold142 (.A(\atari2600.ram[122][3] ),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold143 (.A(\atari2600.ram[62][1] ),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold144 (.A(\scanline[112][0] ),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold145 (.A(\atari2600.ram[77][6] ),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold146 (.A(\atari2600.ram[98][2] ),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold147 (.A(\atari2600.tia.cx[10] ),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold148 (.A(\atari2600.ram[3][6] ),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold149 (.A(\atari2600.ram[78][5] ),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold150 (.A(\atari2600.ram[58][2] ),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold151 (.A(\atari2600.ram[122][7] ),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold152 (.A(\atari2600.ram[93][6] ),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold153 (.A(\atari2600.ram[34][4] ),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold154 (.A(\atari2600.pia.swa_dir[5] ),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold155 (.A(\atari2600.ram[14][2] ),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold156 (.A(\atari2600.ram[66][3] ),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold157 (.A(\atari2600.ram[91][7] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold158 (.A(\atari2600.ram[77][0] ),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold159 (.A(\atari2600.ram[98][1] ),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold160 (.A(\atari2600.ram[106][0] ),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold161 (.A(\atari2600.ram[46][0] ),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold162 (.A(\atari2600.ram[58][0] ),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold163 (.A(\atari2600.ram[58][1] ),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold164 (.A(\atari2600.tia.old_grp1[3] ),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold165 (.A(_01823_),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold166 (.A(\atari2600.tia.poly5_r.x[2] ),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold167 (.A(_02246_),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold168 (.A(\atari2600.ram[93][5] ),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold169 (.A(\atari2600.ram[94][7] ),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold170 (.A(\atari2600.ram[77][4] ),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold171 (.A(\atari2600.ram[88][7] ),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold172 (.A(\atari2600.ram[73][6] ),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold173 (.A(\atari2600.ram[62][6] ),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold174 (.A(\atari2600.ram[6][7] ),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold175 (.A(\atari2600.pia.dat_o[6] ),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold176 (.A(_01770_),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold177 (.A(\scanline[110][4] ),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold178 (.A(\atari2600.ram[18][1] ),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold179 (.A(\atari2600.tia.audio_left_counter[7] ),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold180 (.A(_05919_),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold181 (.A(\atari2600.cpu.IRHOLD[7] ),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold182 (.A(_02464_),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold183 (.A(\atari2600.ram[38][7] ),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold184 (.A(\atari2600.ram[70][5] ),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold185 (.A(\atari2600.ram[30][1] ),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold186 (.A(\atari2600.ram[30][2] ),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold187 (.A(\atari2600.ram[14][3] ),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold188 (.A(\atari2600.ram[74][4] ),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold189 (.A(\atari2600.ram[78][2] ),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold190 (.A(\atari2600.ram[77][3] ),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold191 (.A(\atari2600.ram[1][5] ),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold192 (.A(\atari2600.ram[26][2] ),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold193 (.A(\atari2600.tia.vblank ),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold194 (.A(\atari2600.ram[106][6] ),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold195 (.A(\atari2600.ram[95][7] ),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold196 (.A(\atari2600.pia.swb_dir[4] ),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold197 (.A(\atari2600.ram[90][4] ),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold198 (.A(\atari2600.ram[78][0] ),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold199 (.A(\atari2600.ram[70][0] ),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold200 (.A(\atari2600.ram[126][5] ),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold201 (.A(\atari2600.ram[75][6] ),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold202 (.A(\atari2600.ram[75][0] ),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold203 (.A(\atari2600.ram[14][6] ),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold204 (.A(\atari2600.ram[14][0] ),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold205 (.A(\atari2600.ram[74][3] ),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold206 (.A(\atari2600.ram[10][1] ),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold207 (.A(\atari2600.ram[72][3] ),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold208 (.A(\atari2600.ram[92][4] ),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold209 (.A(\atari2600.ram[70][4] ),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold210 (.A(\atari2600.ram[79][7] ),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold211 (.A(\atari2600.ram[1][6] ),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold212 (.A(\atari2600.ram[34][5] ),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold213 (.A(\atari2600.ram[77][5] ),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold214 (.A(\atari2600.ram[95][4] ),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold215 (.A(\atari2600.ram[72][4] ),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold216 (.A(\atari2600.ram[54][3] ),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold217 (.A(\scanline[45][2] ),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold218 (.A(\atari2600.ram[6][0] ),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold219 (.A(\atari2600.ram[95][3] ),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold220 (.A(\atari2600.ram[38][6] ),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold221 (.A(\atari2600.ram[66][1] ),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold222 (.A(\atari2600.ram[82][6] ),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold223 (.A(\atari2600.ram[95][2] ),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold224 (.A(\atari2600.ram[102][1] ),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold225 (.A(\atari2600.ram[62][0] ),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold226 (.A(\scanline[124][6] ),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold227 (.A(\atari2600.cpu.ALU.BI7 ),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold228 (.A(\atari2600.tia.audio_left_counter[12] ),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold229 (.A(_02024_),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold230 (.A(\atari2600.ram[70][7] ),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold231 (.A(\scanline[90][1] ),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold232 (.A(spi_restart),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold233 (.A(\atari2600.ram[118][0] ),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold234 (.A(\atari2600.ram[50][6] ),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold235 (.A(\atari2600.ram[86][4] ),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold236 (.A(\atari2600.ram[122][2] ),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold237 (.A(\scanline[121][0] ),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold238 (.A(\atari2600.ram[98][0] ),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold239 (.A(\atari2600.ram[110][4] ),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold240 (.A(\atari2600.tia.p0_copies[1] ),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold241 (.A(\scanline[119][6] ),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold242 (.A(\atari2600.ram[91][3] ),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold243 (.A(\atari2600.tia.audio_left_counter[4] ),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold244 (.A(_02016_),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold245 (.A(\scanline[29][2] ),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold246 (.A(\atari2600.ram[118][5] ),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold247 (.A(\atari2600.ram[34][3] ),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold248 (.A(\scanline[62][6] ),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold249 (.A(\atari2600.ram[77][7] ),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold250 (.A(\scanline[158][2] ),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold251 (.A(\scanline[117][4] ),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold252 (.A(\scanline[53][6] ),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold253 (.A(\atari2600.ram[110][1] ),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold254 (.A(\atari2600.ram[88][3] ),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold255 (.A(\atari2600.tia.audio_left_counter[8] ),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold256 (.A(_02020_),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold257 (.A(\atari2600.ram[2][7] ),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold258 (.A(\scanline[78][3] ),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold259 (.A(\atari2600.ram[54][6] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold260 (.A(\scanline[95][4] ),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold261 (.A(\atari2600.ram[46][4] ),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold262 (.A(\scanline[45][5] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold263 (.A(\atari2600.ram[95][1] ),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold264 (.A(\scanline[95][1] ),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold265 (.A(\atari2600.pia.instat[0] ),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold266 (.A(_02309_),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold267 (.A(\scanline[109][0] ),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold268 (.A(\atari2600.ram[76][5] ),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold269 (.A(_00142_),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold270 (.A(_07594_),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold271 (.A(\atari2600.ram[90][7] ),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold272 (.A(\atari2600.ram[94][0] ),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold273 (.A(\scanline[126][6] ),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold274 (.A(\scanline[54][6] ),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold275 (.A(\atari2600.ram[76][6] ),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold276 (.A(\atari2600.ram[110][5] ),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold277 (.A(\scanline[53][0] ),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold278 (.A(\atari2600.pia.time_counter[5] ),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold279 (.A(_05307_),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold280 (.A(\scanline[89][4] ),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold281 (.A(\atari2600.ram[93][7] ),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold282 (.A(\atari2600.rom_data[4] ),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold283 (.A(_02924_),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold284 (.A(\atari2600.ram[22][2] ),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold285 (.A(\atari2600.ram[42][4] ),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold286 (.A(\atari2600.ram[86][7] ),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold287 (.A(\scanline[119][3] ),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold288 (.A(\scanline[101][3] ),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold289 (.A(\atari2600.ram[58][4] ),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold290 (.A(\scanline[123][6] ),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold291 (.A(\scanline[85][2] ),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold292 (.A(\scanline[45][1] ),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold293 (.A(\scanline[89][3] ),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold294 (.A(\scanline[105][5] ),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold295 (.A(\atari2600.ram[106][5] ),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold296 (.A(\atari2600.ram[46][2] ),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold297 (.A(\scanline[30][4] ),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold298 (.A(\atari2600.ram[26][7] ),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold299 (.A(\scanline[102][5] ),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold300 (.A(\scanline[57][6] ),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold301 (.A(\atari2600.ram[93][2] ),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold302 (.A(\scanline[15][1] ),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold303 (.A(\atari2600.ram[58][6] ),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold304 (.A(\scanline[29][5] ),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold305 (.A(\atari2600.ram[73][3] ),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold306 (.A(\scanline[90][5] ),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold307 (.A(\atari2600.ram[54][4] ),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold308 (.A(\scanline[91][3] ),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold309 (.A(\atari2600.ram[79][1] ),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold310 (.A(\scanline[110][3] ),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold311 (.A(\atari2600.tia.old_grp0[3] ),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold312 (.A(_02123_),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold313 (.A(\atari2600.ram[88][0] ),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold314 (.A(\scanline[159][4] ),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold315 (.A(\scanline[151][4] ),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold316 (.A(\scanline[121][1] ),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold317 (.A(\atari2600.ram[88][5] ),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold318 (.A(\atari2600.ram[34][1] ),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold319 (.A(\scanline[86][5] ),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold320 (.A(\atari2600.ram[78][7] ),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold321 (.A(\scanline[101][4] ),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold322 (.A(\scanline[118][0] ),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold323 (.A(\scanline[87][2] ),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold324 (.A(\scanline[158][4] ),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold325 (.A(\scanline[118][6] ),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold326 (.A(\scanline[125][4] ),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold327 (.A(\atari2600.ram[76][1] ),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold328 (.A(\atari2600.tia.old_grp0[5] ),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold329 (.A(_02125_),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold330 (.A(\scanline[143][6] ),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold331 (.A(\scanline[62][3] ),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold332 (.A(\atari2600.tia.cx[12] ),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold333 (.A(\scanline[149][2] ),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold334 (.A(\scanline[141][2] ),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold335 (.A(\scanline[86][1] ),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold336 (.A(\atari2600.ram[42][2] ),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold337 (.A(\scanline[111][1] ),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold338 (.A(\scanline[55][2] ),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold339 (.A(\scanline[119][5] ),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold340 (.A(\atari2600.ram[30][0] ),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold341 (.A(\atari2600.ram[10][6] ),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold342 (.A(\atari2600.tia.poly5_l.x[1] ),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold343 (.A(_02227_),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold344 (.A(\scanline[114][2] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold345 (.A(\scanline[109][2] ),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold346 (.A(\scanline[111][2] ),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold347 (.A(\atari2600.ram[30][6] ),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold348 (.A(\scanline[51][6] ),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold349 (.A(\atari2600.tia.old_grp0[6] ),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold350 (.A(_02126_),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold351 (.A(\atari2600.tia.poly9_l.x[2] ),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold352 (.A(_02233_),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold353 (.A(\atari2600.ram[18][4] ),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold354 (.A(\atari2600.pia.swb_dir[2] ),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold355 (.A(\atari2600.ram[114][6] ),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold356 (.A(\scanline[125][3] ),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold357 (.A(\atari2600.ram[76][3] ),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold358 (.A(\scanline[147][0] ),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold359 (.A(\atari2600.ram[88][4] ),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold360 (.A(\scanline[105][1] ),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold361 (.A(\scanline[54][4] ),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold362 (.A(\atari2600.ram[22][4] ),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold363 (.A(\atari2600.ram[22][5] ),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold364 (.A(\scanline[118][1] ),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold365 (.A(\scanline[126][3] ),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold366 (.A(\atari2600.ram[88][2] ),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold367 (.A(\atari2600.ram[34][2] ),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold368 (.A(\scanline[114][5] ),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold369 (.A(\scanline[46][3] ),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold370 (.A(\scanline[107][2] ),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold371 (.A(\scanline[14][2] ),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold372 (.A(\atari2600.ram[54][5] ),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold373 (.A(\scanline[106][3] ),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold374 (.A(\scanline[46][1] ),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold375 (.A(\scanline[15][0] ),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold376 (.A(\scanline[83][2] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold377 (.A(\atari2600.ram[74][1] ),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold378 (.A(\atari2600.ram[79][4] ),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold379 (.A(\atari2600.ram[2][1] ),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold380 (.A(\scanline[123][0] ),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold381 (.A(\atari2600.tia.old_grp0[7] ),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold382 (.A(_02127_),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold383 (.A(\scanline[121][3] ),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold384 (.A(\scanline[77][6] ),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold385 (.A(\atari2600.ram[86][0] ),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold386 (.A(\scanline[89][2] ),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold387 (.A(\atari2600.tia.audv1[1] ),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold388 (.A(\scanline[15][5] ),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold389 (.A(\atari2600.ram[46][3] ),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold390 (.A(_00050_),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold391 (.A(\atari2600.ram[110][6] ),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold392 (.A(\scanline[53][2] ),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold393 (.A(\scanline[110][1] ),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold394 (.A(\scanline[95][3] ),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold395 (.A(\scanline[113][2] ),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold396 (.A(\atari2600.ram[79][3] ),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold397 (.A(\scanline[93][1] ),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold398 (.A(\atari2600.ram[79][2] ),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold399 (.A(\atari2600.ram[3][1] ),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold400 (.A(\scanline[61][6] ),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold401 (.A(\scanline[45][4] ),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold402 (.A(\atari2600.ram[92][0] ),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold403 (.A(\scanline[154][2] ),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold404 (.A(\scanline[127][2] ),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold405 (.A(\atari2600.ram[10][4] ),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold406 (.A(\scanline[61][1] ),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold407 (.A(\scanline[102][3] ),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold408 (.A(\atari2600.ram[118][3] ),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold409 (.A(\scanline[126][0] ),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold410 (.A(\atari2600.ram[73][7] ),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold411 (.A(\scanline[155][0] ),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold412 (.A(\scanline[157][5] ),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold413 (.A(\scanline[30][3] ),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold414 (.A(\atari2600.ram[2][3] ),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold415 (.A(\atari2600.cpu.src_reg[1] ),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold416 (.A(\scanline[77][2] ),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold417 (.A(\scanline[101][6] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold418 (.A(\scanline[154][0] ),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold419 (.A(\atari2600.ram[70][1] ),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold420 (.A(\scanline[58][0] ),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold421 (.A(\scanline[59][6] ),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold422 (.A(\scanline[15][2] ),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold423 (.A(\atari2600.pia.dat_o[2] ),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold424 (.A(_01766_),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold425 (.A(\scanline[119][1] ),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold426 (.A(\scanline[93][0] ),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold427 (.A(\scanline[55][3] ),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold428 (.A(\atari2600.ram[74][6] ),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold429 (.A(\atari2600.ram[3][4] ),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold430 (.A(\atari2600.ram[89][6] ),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold431 (.A(\scanline[141][5] ),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold432 (.A(\atari2600.ram[1][4] ),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold433 (.A(\scanline[110][5] ),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold434 (.A(\scanline[55][4] ),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold435 (.A(\atari2600.ram[10][7] ),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold436 (.A(\atari2600.ram[93][1] ),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold437 (.A(\scanline[117][5] ),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold438 (.A(\atari2600.tia.audio_left_counter[11] ),
    .X(net3328));
 sg13g2_dlygate4sd3_1 hold439 (.A(_05937_),
    .X(net3329));
 sg13g2_dlygate4sd3_1 hold440 (.A(\atari2600.ram[62][4] ),
    .X(net3330));
 sg13g2_dlygate4sd3_1 hold441 (.A(\atari2600.ram[14][4] ),
    .X(net3331));
 sg13g2_dlygate4sd3_1 hold442 (.A(\scanline[127][5] ),
    .X(net3332));
 sg13g2_dlygate4sd3_1 hold443 (.A(\scanline[105][2] ),
    .X(net3333));
 sg13g2_dlygate4sd3_1 hold444 (.A(\scanline[119][0] ),
    .X(net3334));
 sg13g2_dlygate4sd3_1 hold445 (.A(\scanline[109][4] ),
    .X(net3335));
 sg13g2_dlygate4sd3_1 hold446 (.A(\atari2600.ram[82][2] ),
    .X(net3336));
 sg13g2_dlygate4sd3_1 hold447 (.A(\scanline[155][2] ),
    .X(net3337));
 sg13g2_dlygate4sd3_1 hold448 (.A(\scanline[29][6] ),
    .X(net3338));
 sg13g2_dlygate4sd3_1 hold449 (.A(\atari2600.ram[110][2] ),
    .X(net3339));
 sg13g2_dlygate4sd3_1 hold450 (.A(\atari2600.ram[18][2] ),
    .X(net3340));
 sg13g2_dlygate4sd3_1 hold451 (.A(\scanline[94][4] ),
    .X(net3341));
 sg13g2_dlygate4sd3_1 hold452 (.A(\scanline[95][0] ),
    .X(net3342));
 sg13g2_dlygate4sd3_1 hold453 (.A(\scanline[54][0] ),
    .X(net3343));
 sg13g2_dlygate4sd3_1 hold454 (.A(\atari2600.ram[102][2] ),
    .X(net3344));
 sg13g2_dlygate4sd3_1 hold455 (.A(\scanline[122][6] ),
    .X(net3345));
 sg13g2_dlygate4sd3_1 hold456 (.A(\scanline[105][3] ),
    .X(net3346));
 sg13g2_dlygate4sd3_1 hold457 (.A(\scanline[29][1] ),
    .X(net3347));
 sg13g2_dlygate4sd3_1 hold458 (.A(\atari2600.ram[42][5] ),
    .X(net3348));
 sg13g2_dlygate4sd3_1 hold459 (.A(\scanline[107][3] ),
    .X(net3349));
 sg13g2_dlygate4sd3_1 hold460 (.A(\scanline[151][6] ),
    .X(net3350));
 sg13g2_dlygate4sd3_1 hold461 (.A(\atari2600.pia.swa_dir[3] ),
    .X(net3351));
 sg13g2_dlygate4sd3_1 hold462 (.A(\scanline[106][6] ),
    .X(net3352));
 sg13g2_dlygate4sd3_1 hold463 (.A(\atari2600.ram[82][4] ),
    .X(net3353));
 sg13g2_dlygate4sd3_1 hold464 (.A(\atari2600.rom_data[7] ),
    .X(net3354));
 sg13g2_dlygate4sd3_1 hold465 (.A(_02927_),
    .X(net3355));
 sg13g2_dlygate4sd3_1 hold466 (.A(\scanline[29][3] ),
    .X(net3356));
 sg13g2_dlygate4sd3_1 hold467 (.A(\scanline[122][2] ),
    .X(net3357));
 sg13g2_dlygate4sd3_1 hold468 (.A(\scanline[85][5] ),
    .X(net3358));
 sg13g2_dlygate4sd3_1 hold469 (.A(\atari2600.ram[6][5] ),
    .X(net3359));
 sg13g2_dlygate4sd3_1 hold470 (.A(\scanline[86][0] ),
    .X(net3360));
 sg13g2_dlygate4sd3_1 hold471 (.A(\scanline[54][1] ),
    .X(net3361));
 sg13g2_dlygate4sd3_1 hold472 (.A(\scanline[78][1] ),
    .X(net3362));
 sg13g2_dlygate4sd3_1 hold473 (.A(\scanline[114][0] ),
    .X(net3363));
 sg13g2_dlygate4sd3_1 hold474 (.A(\atari2600.tia.old_grp0[4] ),
    .X(net3364));
 sg13g2_dlygate4sd3_1 hold475 (.A(_02124_),
    .X(net3365));
 sg13g2_dlygate4sd3_1 hold476 (.A(\atari2600.ram[26][6] ),
    .X(net3366));
 sg13g2_dlygate4sd3_1 hold477 (.A(\scanline[142][1] ),
    .X(net3367));
 sg13g2_dlygate4sd3_1 hold478 (.A(\scanline[147][4] ),
    .X(net3368));
 sg13g2_dlygate4sd3_1 hold479 (.A(\atari2600.tia.diag[105] ),
    .X(net3369));
 sg13g2_dlygate4sd3_1 hold480 (.A(_02121_),
    .X(net3370));
 sg13g2_dlygate4sd3_1 hold481 (.A(\atari2600.cpu.ABL[6] ),
    .X(net3371));
 sg13g2_dlygate4sd3_1 hold482 (.A(\atari2600.ram[91][4] ),
    .X(net3372));
 sg13g2_dlygate4sd3_1 hold483 (.A(\scanline[141][4] ),
    .X(net3373));
 sg13g2_dlygate4sd3_1 hold484 (.A(\scanline[13][4] ),
    .X(net3374));
 sg13g2_dlygate4sd3_1 hold485 (.A(\scanline[90][4] ),
    .X(net3375));
 sg13g2_dlygate4sd3_1 hold486 (.A(\scanline[57][0] ),
    .X(net3376));
 sg13g2_dlygate4sd3_1 hold487 (.A(\atari2600.ram[98][7] ),
    .X(net3377));
 sg13g2_dlygate4sd3_1 hold488 (.A(\atari2600.tia.audv0[3] ),
    .X(net3378));
 sg13g2_dlygate4sd3_1 hold489 (.A(\atari2600.tia.audv1[0] ),
    .X(net3379));
 sg13g2_dlygate4sd3_1 hold490 (.A(\atari2600.ram[89][3] ),
    .X(net3380));
 sg13g2_dlygate4sd3_1 hold491 (.A(\scanline[126][5] ),
    .X(net3381));
 sg13g2_dlygate4sd3_1 hold492 (.A(\atari2600.ram[86][2] ),
    .X(net3382));
 sg13g2_dlygate4sd3_1 hold493 (.A(\atari2600.ram[76][2] ),
    .X(net3383));
 sg13g2_dlygate4sd3_1 hold494 (.A(\scanline[14][3] ),
    .X(net3384));
 sg13g2_dlygate4sd3_1 hold495 (.A(\scanline[55][6] ),
    .X(net3385));
 sg13g2_dlygate4sd3_1 hold496 (.A(\scanline[29][0] ),
    .X(net3386));
 sg13g2_dlygate4sd3_1 hold497 (.A(\scanline[125][5] ),
    .X(net3387));
 sg13g2_dlygate4sd3_1 hold498 (.A(\scanline[89][1] ),
    .X(net3388));
 sg13g2_dlygate4sd3_1 hold499 (.A(\scanline[155][6] ),
    .X(net3389));
 sg13g2_dlygate4sd3_1 hold500 (.A(\scanline[159][3] ),
    .X(net3390));
 sg13g2_dlygate4sd3_1 hold501 (.A(\scanline[115][6] ),
    .X(net3391));
 sg13g2_dlygate4sd3_1 hold502 (.A(\scanline[61][3] ),
    .X(net3392));
 sg13g2_dlygate4sd3_1 hold503 (.A(\scanline[158][0] ),
    .X(net3393));
 sg13g2_dlygate4sd3_1 hold504 (.A(\scanline[91][1] ),
    .X(net3394));
 sg13g2_dlygate4sd3_1 hold505 (.A(\scanline[93][4] ),
    .X(net3395));
 sg13g2_dlygate4sd3_1 hold506 (.A(\scanline[77][5] ),
    .X(net3396));
 sg13g2_dlygate4sd3_1 hold507 (.A(\atari2600.ram[66][5] ),
    .X(net3397));
 sg13g2_dlygate4sd3_1 hold508 (.A(\scanline[149][1] ),
    .X(net3398));
 sg13g2_dlygate4sd3_1 hold509 (.A(\scanline[29][4] ),
    .X(net3399));
 sg13g2_dlygate4sd3_1 hold510 (.A(\scanline[109][1] ),
    .X(net3400));
 sg13g2_dlygate4sd3_1 hold511 (.A(\scanline[59][1] ),
    .X(net3401));
 sg13g2_dlygate4sd3_1 hold512 (.A(\scanline[119][2] ),
    .X(net3402));
 sg13g2_dlygate4sd3_1 hold513 (.A(\scanline[153][6] ),
    .X(net3403));
 sg13g2_dlygate4sd3_1 hold514 (.A(\atari2600.ram[38][3] ),
    .X(net3404));
 sg13g2_dlygate4sd3_1 hold515 (.A(\scanline[118][3] ),
    .X(net3405));
 sg13g2_dlygate4sd3_1 hold516 (.A(\atari2600.ram[14][1] ),
    .X(net3406));
 sg13g2_dlygate4sd3_1 hold517 (.A(\atari2600.ram[30][7] ),
    .X(net3407));
 sg13g2_dlygate4sd3_1 hold518 (.A(\scanline[62][1] ),
    .X(net3408));
 sg13g2_dlygate4sd3_1 hold519 (.A(\atari2600.pia.dat_o[7] ),
    .X(net3409));
 sg13g2_dlygate4sd3_1 hold520 (.A(_01771_),
    .X(net3410));
 sg13g2_dlygate4sd3_1 hold521 (.A(\atari2600.tia.audio_left_counter[3] ),
    .X(net3411));
 sg13g2_dlygate4sd3_1 hold522 (.A(_05902_),
    .X(net3412));
 sg13g2_dlygate4sd3_1 hold523 (.A(\scanline[83][3] ),
    .X(net3413));
 sg13g2_dlygate4sd3_1 hold524 (.A(\atari2600.pia.time_counter[18] ),
    .X(net3414));
 sg13g2_dlygate4sd3_1 hold525 (.A(_05339_),
    .X(net3415));
 sg13g2_dlygate4sd3_1 hold526 (.A(_01790_),
    .X(net3416));
 sg13g2_dlygate4sd3_1 hold527 (.A(\scanline[61][2] ),
    .X(net3417));
 sg13g2_dlygate4sd3_1 hold528 (.A(\scanline[89][6] ),
    .X(net3418));
 sg13g2_dlygate4sd3_1 hold529 (.A(\scanline[142][0] ),
    .X(net3419));
 sg13g2_dlygate4sd3_1 hold530 (.A(\scanline[94][2] ),
    .X(net3420));
 sg13g2_dlygate4sd3_1 hold531 (.A(\atari2600.ram[1][2] ),
    .X(net3421));
 sg13g2_dlygate4sd3_1 hold532 (.A(\scanline[57][3] ),
    .X(net3422));
 sg13g2_dlygate4sd3_1 hold533 (.A(\scanline[46][2] ),
    .X(net3423));
 sg13g2_dlygate4sd3_1 hold534 (.A(\scanline[111][3] ),
    .X(net3424));
 sg13g2_dlygate4sd3_1 hold535 (.A(\atari2600.ram[91][2] ),
    .X(net3425));
 sg13g2_dlygate4sd3_1 hold536 (.A(\atari2600.ram[114][2] ),
    .X(net3426));
 sg13g2_dlygate4sd3_1 hold537 (.A(\scanline[115][4] ),
    .X(net3427));
 sg13g2_dlygate4sd3_1 hold538 (.A(\scanline[53][3] ),
    .X(net3428));
 sg13g2_dlygate4sd3_1 hold539 (.A(\scanline[123][3] ),
    .X(net3429));
 sg13g2_dlygate4sd3_1 hold540 (.A(\atari2600.cpu.ABL[3] ),
    .X(net3430));
 sg13g2_dlygate4sd3_1 hold541 (.A(_02482_),
    .X(net3431));
 sg13g2_dlygate4sd3_1 hold542 (.A(\scanline[111][5] ),
    .X(net3432));
 sg13g2_dlygate4sd3_1 hold543 (.A(\scanline[95][5] ),
    .X(net3433));
 sg13g2_dlygate4sd3_1 hold544 (.A(\scanline[124][5] ),
    .X(net3434));
 sg13g2_dlygate4sd3_1 hold545 (.A(\scanline[102][1] ),
    .X(net3435));
 sg13g2_dlygate4sd3_1 hold546 (.A(\scanline[118][5] ),
    .X(net3436));
 sg13g2_dlygate4sd3_1 hold547 (.A(\scanline[14][5] ),
    .X(net3437));
 sg13g2_dlygate4sd3_1 hold548 (.A(\scanline[77][1] ),
    .X(net3438));
 sg13g2_dlygate4sd3_1 hold549 (.A(\atari2600.ram[106][2] ),
    .X(net3439));
 sg13g2_dlygate4sd3_1 hold550 (.A(\scanline[143][4] ),
    .X(net3440));
 sg13g2_dlygate4sd3_1 hold551 (.A(\scanline[79][1] ),
    .X(net3441));
 sg13g2_dlygate4sd3_1 hold552 (.A(\scanline[110][2] ),
    .X(net3442));
 sg13g2_dlygate4sd3_1 hold553 (.A(\scanline[91][6] ),
    .X(net3443));
 sg13g2_dlygate4sd3_1 hold554 (.A(\scanline[86][6] ),
    .X(net3444));
 sg13g2_dlygate4sd3_1 hold555 (.A(\scanline[85][4] ),
    .X(net3445));
 sg13g2_dlygate4sd3_1 hold556 (.A(\scanline[122][3] ),
    .X(net3446));
 sg13g2_dlygate4sd3_1 hold557 (.A(\atari2600.ram[62][5] ),
    .X(net3447));
 sg13g2_dlygate4sd3_1 hold558 (.A(\scanline[127][4] ),
    .X(net3448));
 sg13g2_dlygate4sd3_1 hold559 (.A(\scanline[159][0] ),
    .X(net3449));
 sg13g2_dlygate4sd3_1 hold560 (.A(\scanline[31][5] ),
    .X(net3450));
 sg13g2_dlygate4sd3_1 hold561 (.A(\scanline[157][2] ),
    .X(net3451));
 sg13g2_dlygate4sd3_1 hold562 (.A(\atari2600.ram[46][6] ),
    .X(net3452));
 sg13g2_dlygate4sd3_1 hold563 (.A(\scanline[158][1] ),
    .X(net3453));
 sg13g2_dlygate4sd3_1 hold564 (.A(\atari2600.ram[6][6] ),
    .X(net3454));
 sg13g2_dlygate4sd3_1 hold565 (.A(\atari2600.ram[94][2] ),
    .X(net3455));
 sg13g2_dlygate4sd3_1 hold566 (.A(\atari2600.ram[18][6] ),
    .X(net3456));
 sg13g2_dlygate4sd3_1 hold567 (.A(\scanline[87][6] ),
    .X(net3457));
 sg13g2_dlygate4sd3_1 hold568 (.A(\scanline[124][2] ),
    .X(net3458));
 sg13g2_dlygate4sd3_1 hold569 (.A(\scanline[90][2] ),
    .X(net3459));
 sg13g2_dlygate4sd3_1 hold570 (.A(\scanline[30][1] ),
    .X(net3460));
 sg13g2_dlygate4sd3_1 hold571 (.A(\atari2600.tia.old_grp0[0] ),
    .X(net3461));
 sg13g2_dlygate4sd3_1 hold572 (.A(_02120_),
    .X(net3462));
 sg13g2_dlygate4sd3_1 hold573 (.A(\scanline[91][4] ),
    .X(net3463));
 sg13g2_dlygate4sd3_1 hold574 (.A(_00106_),
    .X(net3464));
 sg13g2_dlygate4sd3_1 hold575 (.A(_05890_),
    .X(net3465));
 sg13g2_dlygate4sd3_1 hold576 (.A(_02012_),
    .X(net3466));
 sg13g2_dlygate4sd3_1 hold577 (.A(\scanline[63][4] ),
    .X(net3467));
 sg13g2_dlygate4sd3_1 hold578 (.A(\scanline[79][3] ),
    .X(net3468));
 sg13g2_dlygate4sd3_1 hold579 (.A(\scanline[78][4] ),
    .X(net3469));
 sg13g2_dlygate4sd3_1 hold580 (.A(\scanline[123][1] ),
    .X(net3470));
 sg13g2_dlygate4sd3_1 hold581 (.A(\atari2600.ram[70][2] ),
    .X(net3471));
 sg13g2_dlygate4sd3_1 hold582 (.A(\atari2600.ram[22][7] ),
    .X(net3472));
 sg13g2_dlygate4sd3_1 hold583 (.A(\atari2600.tia.audio_left_counter[5] ),
    .X(net3473));
 sg13g2_dlygate4sd3_1 hold584 (.A(_05910_),
    .X(net3474));
 sg13g2_dlygate4sd3_1 hold585 (.A(\scanline[78][0] ),
    .X(net3475));
 sg13g2_dlygate4sd3_1 hold586 (.A(\scanline[153][4] ),
    .X(net3476));
 sg13g2_dlygate4sd3_1 hold587 (.A(\atari2600.ram[90][5] ),
    .X(net3477));
 sg13g2_dlygate4sd3_1 hold588 (.A(\scanline[115][5] ),
    .X(net3478));
 sg13g2_dlygate4sd3_1 hold589 (.A(_00060_),
    .X(net3479));
 sg13g2_dlygate4sd3_1 hold590 (.A(_04867_),
    .X(net3480));
 sg13g2_dlygate4sd3_1 hold591 (.A(\scanline[113][0] ),
    .X(net3481));
 sg13g2_dlygate4sd3_1 hold592 (.A(\scanline[78][2] ),
    .X(net3482));
 sg13g2_dlygate4sd3_1 hold593 (.A(\scanline[126][2] ),
    .X(net3483));
 sg13g2_dlygate4sd3_1 hold594 (.A(\scanline[115][0] ),
    .X(net3484));
 sg13g2_dlygate4sd3_1 hold595 (.A(\atari2600.ram[2][6] ),
    .X(net3485));
 sg13g2_dlygate4sd3_1 hold596 (.A(\scanline[13][2] ),
    .X(net3486));
 sg13g2_dlygate4sd3_1 hold597 (.A(\atari2600.cpu.ABL[4] ),
    .X(net3487));
 sg13g2_dlygate4sd3_1 hold598 (.A(\atari2600.ram[91][5] ),
    .X(net3488));
 sg13g2_dlygate4sd3_1 hold599 (.A(\atari2600.ram[92][5] ),
    .X(net3489));
 sg13g2_dlygate4sd3_1 hold600 (.A(\scanline[118][4] ),
    .X(net3490));
 sg13g2_dlygate4sd3_1 hold601 (.A(\atari2600.cpu.AXYS[1][1] ),
    .X(net3491));
 sg13g2_dlygate4sd3_1 hold602 (.A(\atari2600.cpu.AXYS[3][1] ),
    .X(net3492));
 sg13g2_dlygate4sd3_1 hold603 (.A(\scanline[58][2] ),
    .X(net3493));
 sg13g2_dlygate4sd3_1 hold604 (.A(\scanline[153][0] ),
    .X(net3494));
 sg13g2_dlygate4sd3_1 hold605 (.A(\scanline[153][2] ),
    .X(net3495));
 sg13g2_dlygate4sd3_1 hold606 (.A(\atari2600.ram[66][4] ),
    .X(net3496));
 sg13g2_dlygate4sd3_1 hold607 (.A(\atari2600.ram[88][6] ),
    .X(net3497));
 sg13g2_dlygate4sd3_1 hold608 (.A(\scanline[87][3] ),
    .X(net3498));
 sg13g2_dlygate4sd3_1 hold609 (.A(\scanline[58][1] ),
    .X(net3499));
 sg13g2_dlygate4sd3_1 hold610 (.A(\atari2600.ram[114][1] ),
    .X(net3500));
 sg13g2_dlygate4sd3_1 hold611 (.A(\atari2600.cpu.AXYS[0][0] ),
    .X(net3501));
 sg13g2_dlygate4sd3_1 hold612 (.A(\scanline[105][0] ),
    .X(net3502));
 sg13g2_dlygate4sd3_1 hold613 (.A(\scanline[87][5] ),
    .X(net3503));
 sg13g2_dlygate4sd3_1 hold614 (.A(\scanline[102][0] ),
    .X(net3504));
 sg13g2_dlygate4sd3_1 hold615 (.A(\atari2600.tia.poly4_l.x[2] ),
    .X(net3505));
 sg13g2_dlygate4sd3_1 hold616 (.A(_02225_),
    .X(net3506));
 sg13g2_dlygate4sd3_1 hold617 (.A(\scanline[115][3] ),
    .X(net3507));
 sg13g2_dlygate4sd3_1 hold618 (.A(\atari2600.ram[74][7] ),
    .X(net3508));
 sg13g2_dlygate4sd3_1 hold619 (.A(\scanline[141][6] ),
    .X(net3509));
 sg13g2_dlygate4sd3_1 hold620 (.A(\scanline[117][6] ),
    .X(net3510));
 sg13g2_dlygate4sd3_1 hold621 (.A(\scanline[63][6] ),
    .X(net3511));
 sg13g2_dlygate4sd3_1 hold622 (.A(\scanline[99][0] ),
    .X(net3512));
 sg13g2_dlygate4sd3_1 hold623 (.A(\scanline[53][1] ),
    .X(net3513));
 sg13g2_dlygate4sd3_1 hold624 (.A(\scanline[155][3] ),
    .X(net3514));
 sg13g2_dlygate4sd3_1 hold625 (.A(\scanline[57][2] ),
    .X(net3515));
 sg13g2_dlygate4sd3_1 hold626 (.A(\scanline[58][4] ),
    .X(net3516));
 sg13g2_dlygate4sd3_1 hold627 (.A(\scanline[103][6] ),
    .X(net3517));
 sg13g2_dlygate4sd3_1 hold628 (.A(\scanline[90][0] ),
    .X(net3518));
 sg13g2_dlygate4sd3_1 hold629 (.A(\scanline[83][4] ),
    .X(net3519));
 sg13g2_dlygate4sd3_1 hold630 (.A(\scanline[86][4] ),
    .X(net3520));
 sg13g2_dlygate4sd3_1 hold631 (.A(\scanline[61][0] ),
    .X(net3521));
 sg13g2_dlygate4sd3_1 hold632 (.A(\scanline[107][4] ),
    .X(net3522));
 sg13g2_dlygate4sd3_1 hold633 (.A(\scanline[157][0] ),
    .X(net3523));
 sg13g2_dlygate4sd3_1 hold634 (.A(\scanline[78][5] ),
    .X(net3524));
 sg13g2_dlygate4sd3_1 hold635 (.A(\atari2600.ram[38][2] ),
    .X(net3525));
 sg13g2_dlygate4sd3_1 hold636 (.A(\scanline[79][0] ),
    .X(net3526));
 sg13g2_dlygate4sd3_1 hold637 (.A(\scanline[93][3] ),
    .X(net3527));
 sg13g2_dlygate4sd3_1 hold638 (.A(\frame_counter[2] ),
    .X(net3528));
 sg13g2_dlygate4sd3_1 hold639 (.A(_01202_),
    .X(net3529));
 sg13g2_dlygate4sd3_1 hold640 (.A(\atari2600.ram[50][3] ),
    .X(net3530));
 sg13g2_dlygate4sd3_1 hold641 (.A(\scanline[61][5] ),
    .X(net3531));
 sg13g2_dlygate4sd3_1 hold642 (.A(\atari2600.ram[6][2] ),
    .X(net3532));
 sg13g2_dlygate4sd3_1 hold643 (.A(\atari2600.ram[50][4] ),
    .X(net3533));
 sg13g2_dlygate4sd3_1 hold644 (.A(\scanline[141][3] ),
    .X(net3534));
 sg13g2_dlygate4sd3_1 hold645 (.A(\scanline[141][1] ),
    .X(net3535));
 sg13g2_dlygate4sd3_1 hold646 (.A(\scanline[59][3] ),
    .X(net3536));
 sg13g2_dlygate4sd3_1 hold647 (.A(\scanline[77][3] ),
    .X(net3537));
 sg13g2_dlygate4sd3_1 hold648 (.A(\scanline[147][6] ),
    .X(net3538));
 sg13g2_dlygate4sd3_1 hold649 (.A(\scanline[127][6] ),
    .X(net3539));
 sg13g2_dlygate4sd3_1 hold650 (.A(\scanline[99][2] ),
    .X(net3540));
 sg13g2_dlygate4sd3_1 hold651 (.A(\scanline[150][3] ),
    .X(net3541));
 sg13g2_dlygate4sd3_1 hold652 (.A(\scanline[87][4] ),
    .X(net3542));
 sg13g2_dlygate4sd3_1 hold653 (.A(\scanline[117][3] ),
    .X(net3543));
 sg13g2_dlygate4sd3_1 hold654 (.A(\scanline[79][5] ),
    .X(net3544));
 sg13g2_dlygate4sd3_1 hold655 (.A(\scanline[79][4] ),
    .X(net3545));
 sg13g2_dlygate4sd3_1 hold656 (.A(\scanline[107][5] ),
    .X(net3546));
 sg13g2_dlygate4sd3_1 hold657 (.A(\scanline[13][5] ),
    .X(net3547));
 sg13g2_dlygate4sd3_1 hold658 (.A(\scanline[99][5] ),
    .X(net3548));
 sg13g2_dlygate4sd3_1 hold659 (.A(\scanline[151][3] ),
    .X(net3549));
 sg13g2_dlygate4sd3_1 hold660 (.A(\scanline[122][0] ),
    .X(net3550));
 sg13g2_dlygate4sd3_1 hold661 (.A(\scanline[51][0] ),
    .X(net3551));
 sg13g2_dlygate4sd3_1 hold662 (.A(\scanline[86][2] ),
    .X(net3552));
 sg13g2_dlygate4sd3_1 hold663 (.A(\atari2600.ram[72][5] ),
    .X(net3553));
 sg13g2_dlygate4sd3_1 hold664 (.A(\atari2600.ram[42][0] ),
    .X(net3554));
 sg13g2_dlygate4sd3_1 hold665 (.A(\scanline[31][0] ),
    .X(net3555));
 sg13g2_dlygate4sd3_1 hold666 (.A(\scanline[63][0] ),
    .X(net3556));
 sg13g2_dlygate4sd3_1 hold667 (.A(\atari2600.cpu.AXYS[1][0] ),
    .X(net3557));
 sg13g2_dlygate4sd3_1 hold668 (.A(\scanline[151][5] ),
    .X(net3558));
 sg13g2_dlygate4sd3_1 hold669 (.A(\scanline[13][3] ),
    .X(net3559));
 sg13g2_dlygate4sd3_1 hold670 (.A(\scanline[154][3] ),
    .X(net3560));
 sg13g2_dlygate4sd3_1 hold671 (.A(\scanline[31][1] ),
    .X(net3561));
 sg13g2_dlygate4sd3_1 hold672 (.A(\scanline[91][2] ),
    .X(net3562));
 sg13g2_dlygate4sd3_1 hold673 (.A(\scanline[121][6] ),
    .X(net3563));
 sg13g2_dlygate4sd3_1 hold674 (.A(\scanline[105][6] ),
    .X(net3564));
 sg13g2_dlygate4sd3_1 hold675 (.A(\scanline[62][2] ),
    .X(net3565));
 sg13g2_dlygate4sd3_1 hold676 (.A(\atari2600.ram[122][6] ),
    .X(net3566));
 sg13g2_dlygate4sd3_1 hold677 (.A(\scanline[113][5] ),
    .X(net3567));
 sg13g2_dlygate4sd3_1 hold678 (.A(\atari2600.ram[126][4] ),
    .X(net3568));
 sg13g2_dlygate4sd3_1 hold679 (.A(\scanline[101][5] ),
    .X(net3569));
 sg13g2_dlygate4sd3_1 hold680 (.A(\scanline[13][6] ),
    .X(net3570));
 sg13g2_dlygate4sd3_1 hold681 (.A(\scanline[63][1] ),
    .X(net3571));
 sg13g2_dlygate4sd3_1 hold682 (.A(\atari2600.ram[62][2] ),
    .X(net3572));
 sg13g2_dlygate4sd3_1 hold683 (.A(\scanline[127][1] ),
    .X(net3573));
 sg13g2_dlygate4sd3_1 hold684 (.A(\scanline[111][4] ),
    .X(net3574));
 sg13g2_dlygate4sd3_1 hold685 (.A(\scanline[109][5] ),
    .X(net3575));
 sg13g2_dlygate4sd3_1 hold686 (.A(\atari2600.ram[26][0] ),
    .X(net3576));
 sg13g2_dlygate4sd3_1 hold687 (.A(\scanline[94][0] ),
    .X(net3577));
 sg13g2_dlygate4sd3_1 hold688 (.A(\scanline[31][3] ),
    .X(net3578));
 sg13g2_dlygate4sd3_1 hold689 (.A(\atari2600.ram[14][7] ),
    .X(net3579));
 sg13g2_dlygate4sd3_1 hold690 (.A(\atari2600.pia.time_counter[20] ),
    .X(net3580));
 sg13g2_dlygate4sd3_1 hold691 (.A(_05342_),
    .X(net3581));
 sg13g2_dlygate4sd3_1 hold692 (.A(_01792_),
    .X(net3582));
 sg13g2_dlygate4sd3_1 hold693 (.A(\scanline[123][4] ),
    .X(net3583));
 sg13g2_dlygate4sd3_1 hold694 (.A(\scanline[103][4] ),
    .X(net3584));
 sg13g2_dlygate4sd3_1 hold695 (.A(\scanline[101][1] ),
    .X(net3585));
 sg13g2_dlygate4sd3_1 hold696 (.A(\scanline[159][2] ),
    .X(net3586));
 sg13g2_dlygate4sd3_1 hold697 (.A(\scanline[86][3] ),
    .X(net3587));
 sg13g2_dlygate4sd3_1 hold698 (.A(\atari2600.ram[77][2] ),
    .X(net3588));
 sg13g2_dlygate4sd3_1 hold699 (.A(\scanline[105][4] ),
    .X(net3589));
 sg13g2_dlygate4sd3_1 hold700 (.A(\scanline[90][6] ),
    .X(net3590));
 sg13g2_dlygate4sd3_1 hold701 (.A(\scanline[143][0] ),
    .X(net3591));
 sg13g2_dlygate4sd3_1 hold702 (.A(\scanline[113][4] ),
    .X(net3592));
 sg13g2_dlygate4sd3_1 hold703 (.A(\scanline[51][5] ),
    .X(net3593));
 sg13g2_dlygate4sd3_1 hold704 (.A(\scanline[115][2] ),
    .X(net3594));
 sg13g2_dlygate4sd3_1 hold705 (.A(\scanline[147][5] ),
    .X(net3595));
 sg13g2_dlygate4sd3_1 hold706 (.A(\atari2600.ram[50][7] ),
    .X(net3596));
 sg13g2_dlygate4sd3_1 hold707 (.A(\scanline[63][2] ),
    .X(net3597));
 sg13g2_dlygate4sd3_1 hold708 (.A(\scanline[114][1] ),
    .X(net3598));
 sg13g2_dlygate4sd3_1 hold709 (.A(\scanline[101][0] ),
    .X(net3599));
 sg13g2_dlygate4sd3_1 hold710 (.A(\scanline[113][1] ),
    .X(net3600));
 sg13g2_dlygate4sd3_1 hold711 (.A(\scanline[119][4] ),
    .X(net3601));
 sg13g2_dlygate4sd3_1 hold712 (.A(\atari2600.pia.swa_dir[2] ),
    .X(net3602));
 sg13g2_dlygate4sd3_1 hold713 (.A(\scanline[117][0] ),
    .X(net3603));
 sg13g2_dlygate4sd3_1 hold714 (.A(\atari2600.ram[114][3] ),
    .X(net3604));
 sg13g2_dlygate4sd3_1 hold715 (.A(\scanline[45][0] ),
    .X(net3605));
 sg13g2_dlygate4sd3_1 hold716 (.A(\scanline[95][2] ),
    .X(net3606));
 sg13g2_dlygate4sd3_1 hold717 (.A(\scanline[109][6] ),
    .X(net3607));
 sg13g2_dlygate4sd3_1 hold718 (.A(\scanline[150][6] ),
    .X(net3608));
 sg13g2_dlygate4sd3_1 hold719 (.A(\scanline[159][6] ),
    .X(net3609));
 sg13g2_dlygate4sd3_1 hold720 (.A(\atari2600.ram[94][5] ),
    .X(net3610));
 sg13g2_dlygate4sd3_1 hold721 (.A(\atari2600.ram[90][1] ),
    .X(net3611));
 sg13g2_dlygate4sd3_1 hold722 (.A(\scanline[59][0] ),
    .X(net3612));
 sg13g2_dlygate4sd3_1 hold723 (.A(\scanline[114][4] ),
    .X(net3613));
 sg13g2_dlygate4sd3_1 hold724 (.A(\scanline[159][5] ),
    .X(net3614));
 sg13g2_dlygate4sd3_1 hold725 (.A(\scanline[55][1] ),
    .X(net3615));
 sg13g2_dlygate4sd3_1 hold726 (.A(\scanline[15][6] ),
    .X(net3616));
 sg13g2_dlygate4sd3_1 hold727 (.A(\scanline[151][1] ),
    .X(net3617));
 sg13g2_dlygate4sd3_1 hold728 (.A(\scanline[94][5] ),
    .X(net3618));
 sg13g2_dlygate4sd3_1 hold729 (.A(\scanline[59][2] ),
    .X(net3619));
 sg13g2_dlygate4sd3_1 hold730 (.A(\scanline[113][6] ),
    .X(net3620));
 sg13g2_dlygate4sd3_1 hold731 (.A(\atari2600.ram[118][1] ),
    .X(net3621));
 sg13g2_dlygate4sd3_1 hold732 (.A(\scanline[13][1] ),
    .X(net3622));
 sg13g2_dlygate4sd3_1 hold733 (.A(\atari2600.ram[75][1] ),
    .X(net3623));
 sg13g2_dlygate4sd3_1 hold734 (.A(\scanline[99][1] ),
    .X(net3624));
 sg13g2_dlygate4sd3_1 hold735 (.A(\scanline[114][6] ),
    .X(net3625));
 sg13g2_dlygate4sd3_1 hold736 (.A(\scanline[47][5] ),
    .X(net3626));
 sg13g2_dlygate4sd3_1 hold737 (.A(\atari2600.tia.old_grp0[2] ),
    .X(net3627));
 sg13g2_dlygate4sd3_1 hold738 (.A(_02122_),
    .X(net3628));
 sg13g2_dlygate4sd3_1 hold739 (.A(\scanline[124][4] ),
    .X(net3629));
 sg13g2_dlygate4sd3_1 hold740 (.A(\scanline[127][3] ),
    .X(net3630));
 sg13g2_dlygate4sd3_1 hold741 (.A(\scanline[153][1] ),
    .X(net3631));
 sg13g2_dlygate4sd3_1 hold742 (.A(\atari2600.ram[54][7] ),
    .X(net3632));
 sg13g2_dlygate4sd3_1 hold743 (.A(\atari2600.ram[126][2] ),
    .X(net3633));
 sg13g2_dlygate4sd3_1 hold744 (.A(\scanline[114][3] ),
    .X(net3634));
 sg13g2_dlygate4sd3_1 hold745 (.A(\atari2600.ram[102][5] ),
    .X(net3635));
 sg13g2_dlygate4sd3_1 hold746 (.A(\scanline[15][4] ),
    .X(net3636));
 sg13g2_dlygate4sd3_1 hold747 (.A(\atari2600.ram[90][2] ),
    .X(net3637));
 sg13g2_dlygate4sd3_1 hold748 (.A(\scanline[142][6] ),
    .X(net3638));
 sg13g2_dlygate4sd3_1 hold749 (.A(\atari2600.ram[89][0] ),
    .X(net3639));
 sg13g2_dlygate4sd3_1 hold750 (.A(\scanline[46][6] ),
    .X(net3640));
 sg13g2_dlygate4sd3_1 hold751 (.A(\scanline[30][6] ),
    .X(net3641));
 sg13g2_dlygate4sd3_1 hold752 (.A(\atari2600.ram[70][6] ),
    .X(net3642));
 sg13g2_dlygate4sd3_1 hold753 (.A(\scanline[103][5] ),
    .X(net3643));
 sg13g2_dlygate4sd3_1 hold754 (.A(\atari2600.pia.instat[1] ),
    .X(net3644));
 sg13g2_dlygate4sd3_1 hold755 (.A(\scanline[155][4] ),
    .X(net3645));
 sg13g2_dlygate4sd3_1 hold756 (.A(\flash_rom.addr[14] ),
    .X(net3646));
 sg13g2_dlygate4sd3_1 hold757 (.A(_00214_),
    .X(net3647));
 sg13g2_dlygate4sd3_1 hold758 (.A(\scanline[63][3] ),
    .X(net3648));
 sg13g2_dlygate4sd3_1 hold759 (.A(\scanline[55][0] ),
    .X(net3649));
 sg13g2_dlygate4sd3_1 hold760 (.A(\atari2600.ram[95][6] ),
    .X(net3650));
 sg13g2_dlygate4sd3_1 hold761 (.A(\scanline[85][0] ),
    .X(net3651));
 sg13g2_dlygate4sd3_1 hold762 (.A(\atari2600.ram[50][1] ),
    .X(net3652));
 sg13g2_dlygate4sd3_1 hold763 (.A(\atari2600.ram[126][1] ),
    .X(net3653));
 sg13g2_dlygate4sd3_1 hold764 (.A(\scanline[45][6] ),
    .X(net3654));
 sg13g2_dlygate4sd3_1 hold765 (.A(\scanline[46][0] ),
    .X(net3655));
 sg13g2_dlygate4sd3_1 hold766 (.A(\scanline[151][2] ),
    .X(net3656));
 sg13g2_dlygate4sd3_1 hold767 (.A(\atari2600.ram[38][0] ),
    .X(net3657));
 sg13g2_dlygate4sd3_1 hold768 (.A(\scanline[59][5] ),
    .X(net3658));
 sg13g2_dlygate4sd3_1 hold769 (.A(\atari2600.tia.diag[78] ),
    .X(net3659));
 sg13g2_dlygate4sd3_1 hold770 (.A(\atari2600.ram[2][5] ),
    .X(net3660));
 sg13g2_dlygate4sd3_1 hold771 (.A(\scanline[150][4] ),
    .X(net3661));
 sg13g2_dlygate4sd3_1 hold772 (.A(\atari2600.ram[110][3] ),
    .X(net3662));
 sg13g2_dlygate4sd3_1 hold773 (.A(\atari2600.ram[50][5] ),
    .X(net3663));
 sg13g2_dlygate4sd3_1 hold774 (.A(\scanline[30][5] ),
    .X(net3664));
 sg13g2_dlygate4sd3_1 hold775 (.A(\scanline[124][3] ),
    .X(net3665));
 sg13g2_dlygate4sd3_1 hold776 (.A(\atari2600.ram[78][3] ),
    .X(net3666));
 sg13g2_dlygate4sd3_1 hold777 (.A(\scanline[14][1] ),
    .X(net3667));
 sg13g2_dlygate4sd3_1 hold778 (.A(\atari2600.ram[54][1] ),
    .X(net3668));
 sg13g2_dlygate4sd3_1 hold779 (.A(\atari2600.ram[110][0] ),
    .X(net3669));
 sg13g2_dlygate4sd3_1 hold780 (.A(\scanline[94][1] ),
    .X(net3670));
 sg13g2_dlygate4sd3_1 hold781 (.A(\atari2600.ram[14][5] ),
    .X(net3671));
 sg13g2_dlygate4sd3_1 hold782 (.A(\scanline[121][2] ),
    .X(net3672));
 sg13g2_dlygate4sd3_1 hold783 (.A(\scanline[89][0] ),
    .X(net3673));
 sg13g2_dlygate4sd3_1 hold784 (.A(\scanline[90][3] ),
    .X(net3674));
 sg13g2_dlygate4sd3_1 hold785 (.A(\scanline[87][1] ),
    .X(net3675));
 sg13g2_dlygate4sd3_1 hold786 (.A(\atari2600.tia.audio_left_counter[13] ),
    .X(net3676));
 sg13g2_dlygate4sd3_1 hold787 (.A(_05946_),
    .X(net3677));
 sg13g2_dlygate4sd3_1 hold788 (.A(\scanline[142][4] ),
    .X(net3678));
 sg13g2_dlygate4sd3_1 hold789 (.A(_00077_),
    .X(net3679));
 sg13g2_dlygate4sd3_1 hold790 (.A(_00043_),
    .X(net3680));
 sg13g2_dlygate4sd3_1 hold791 (.A(\scanline[58][3] ),
    .X(net3681));
 sg13g2_dlygate4sd3_1 hold792 (.A(\scanline[115][1] ),
    .X(net3682));
 sg13g2_dlygate4sd3_1 hold793 (.A(\scanline[117][1] ),
    .X(net3683));
 sg13g2_dlygate4sd3_1 hold794 (.A(\atari2600.cpu.V ),
    .X(net3684));
 sg13g2_dlygate4sd3_1 hold795 (.A(_02467_),
    .X(net3685));
 sg13g2_dlygate4sd3_1 hold796 (.A(\scanline[93][6] ),
    .X(net3686));
 sg13g2_dlygate4sd3_1 hold797 (.A(\atari2600.ram[42][1] ),
    .X(net3687));
 sg13g2_dlygate4sd3_1 hold798 (.A(\scanline[127][0] ),
    .X(net3688));
 sg13g2_dlygate4sd3_1 hold799 (.A(\scanline[126][4] ),
    .X(net3689));
 sg13g2_dlygate4sd3_1 hold800 (.A(\scanline[30][2] ),
    .X(net3690));
 sg13g2_dlygate4sd3_1 hold801 (.A(\scanline[15][3] ),
    .X(net3691));
 sg13g2_dlygate4sd3_1 hold802 (.A(\atari2600.ram[22][1] ),
    .X(net3692));
 sg13g2_dlygate4sd3_1 hold803 (.A(\scanline[57][1] ),
    .X(net3693));
 sg13g2_dlygate4sd3_1 hold804 (.A(\atari2600.ram[72][6] ),
    .X(net3694));
 sg13g2_dlygate4sd3_1 hold805 (.A(\scanline[102][6] ),
    .X(net3695));
 sg13g2_dlygate4sd3_1 hold806 (.A(\scanline[14][6] ),
    .X(net3696));
 sg13g2_dlygate4sd3_1 hold807 (.A(\atari2600.ram[86][1] ),
    .X(net3697));
 sg13g2_dlygate4sd3_1 hold808 (.A(\atari2600.ram[106][7] ),
    .X(net3698));
 sg13g2_dlygate4sd3_1 hold809 (.A(\scanline[125][0] ),
    .X(net3699));
 sg13g2_dlygate4sd3_1 hold810 (.A(\atari2600.ram[34][6] ),
    .X(net3700));
 sg13g2_dlygate4sd3_1 hold811 (.A(\atari2600.pia.swa_dir[6] ),
    .X(net3701));
 sg13g2_dlygate4sd3_1 hold812 (.A(\scanline[107][6] ),
    .X(net3702));
 sg13g2_dlygate4sd3_1 hold813 (.A(\atari2600.ram[114][0] ),
    .X(net3703));
 sg13g2_dlygate4sd3_1 hold814 (.A(\atari2600.tia.cx[11] ),
    .X(net3704));
 sg13g2_dlygate4sd3_1 hold815 (.A(\scanline[151][0] ),
    .X(net3705));
 sg13g2_dlygate4sd3_1 hold816 (.A(\atari2600.ram[75][4] ),
    .X(net3706));
 sg13g2_dlygate4sd3_1 hold817 (.A(\flash_rom.addr[19] ),
    .X(net3707));
 sg13g2_dlygate4sd3_1 hold818 (.A(_00218_),
    .X(net3708));
 sg13g2_dlygate4sd3_1 hold819 (.A(\scanline[79][2] ),
    .X(net3709));
 sg13g2_dlygate4sd3_1 hold820 (.A(\flash_rom.addr[22] ),
    .X(net3710));
 sg13g2_dlygate4sd3_1 hold821 (.A(_00217_),
    .X(net3711));
 sg13g2_dlygate4sd3_1 hold822 (.A(\scanline[102][2] ),
    .X(net3712));
 sg13g2_dlygate4sd3_1 hold823 (.A(\atari2600.ram[1][0] ),
    .X(net3713));
 sg13g2_dlygate4sd3_1 hold824 (.A(\scanline[110][0] ),
    .X(net3714));
 sg13g2_dlygate4sd3_1 hold825 (.A(\scanline[55][5] ),
    .X(net3715));
 sg13g2_dlygate4sd3_1 hold826 (.A(\scanline[149][5] ),
    .X(net3716));
 sg13g2_dlygate4sd3_1 hold827 (.A(\scanline[57][4] ),
    .X(net3717));
 sg13g2_dlygate4sd3_1 hold828 (.A(\scanline[83][0] ),
    .X(net3718));
 sg13g2_dlygate4sd3_1 hold829 (.A(\scanline[155][5] ),
    .X(net3719));
 sg13g2_dlygate4sd3_1 hold830 (.A(\atari2600.ram[122][0] ),
    .X(net3720));
 sg13g2_dlygate4sd3_1 hold831 (.A(\scanline[142][3] ),
    .X(net3721));
 sg13g2_dlygate4sd3_1 hold832 (.A(\atari2600.ram[72][0] ),
    .X(net3722));
 sg13g2_dlygate4sd3_1 hold833 (.A(\atari2600.tia.p1_copies[1] ),
    .X(net3723));
 sg13g2_dlygate4sd3_1 hold834 (.A(\atari2600.ram[114][5] ),
    .X(net3724));
 sg13g2_dlygate4sd3_1 hold835 (.A(\scanline[125][2] ),
    .X(net3725));
 sg13g2_dlygate4sd3_1 hold836 (.A(\scanline[143][1] ),
    .X(net3726));
 sg13g2_dlygate4sd3_1 hold837 (.A(\scanline[106][0] ),
    .X(net3727));
 sg13g2_dlygate4sd3_1 hold838 (.A(\scanline[124][0] ),
    .X(net3728));
 sg13g2_dlygate4sd3_1 hold839 (.A(\atari2600.ram[82][1] ),
    .X(net3729));
 sg13g2_dlygate4sd3_1 hold840 (.A(\atari2600.ram[75][7] ),
    .X(net3730));
 sg13g2_dlygate4sd3_1 hold841 (.A(\scanline[157][6] ),
    .X(net3731));
 sg13g2_dlygate4sd3_1 hold842 (.A(\scanline[63][5] ),
    .X(net3732));
 sg13g2_dlygate4sd3_1 hold843 (.A(\r_pwm_even[1] ),
    .X(net3733));
 sg13g2_dlygate4sd3_1 hold844 (.A(_04572_),
    .X(net3734));
 sg13g2_dlygate4sd3_1 hold845 (.A(_01183_),
    .X(net3735));
 sg13g2_dlygate4sd3_1 hold846 (.A(\scanline[125][6] ),
    .X(net3736));
 sg13g2_dlygate4sd3_1 hold847 (.A(\scanline[153][3] ),
    .X(net3737));
 sg13g2_dlygate4sd3_1 hold848 (.A(\atari2600.ram[75][2] ),
    .X(net3738));
 sg13g2_dlygate4sd3_1 hold849 (.A(\scanline[142][2] ),
    .X(net3739));
 sg13g2_dlygate4sd3_1 hold850 (.A(\scanline[58][6] ),
    .X(net3740));
 sg13g2_dlygate4sd3_1 hold851 (.A(\scanline[158][5] ),
    .X(net3741));
 sg13g2_dlygate4sd3_1 hold852 (.A(\scanline[47][1] ),
    .X(net3742));
 sg13g2_dlygate4sd3_1 hold853 (.A(\atari2600.ram[3][0] ),
    .X(net3743));
 sg13g2_dlygate4sd3_1 hold854 (.A(\atari2600.ram[66][6] ),
    .X(net3744));
 sg13g2_dlygate4sd3_1 hold855 (.A(\scanline[14][4] ),
    .X(net3745));
 sg13g2_dlygate4sd3_1 hold856 (.A(\scanline[109][3] ),
    .X(net3746));
 sg13g2_dlygate4sd3_1 hold857 (.A(\atari2600.ram[92][1] ),
    .X(net3747));
 sg13g2_dlygate4sd3_1 hold858 (.A(\scanline[99][4] ),
    .X(net3748));
 sg13g2_dlygate4sd3_1 hold859 (.A(\atari2600.cpu.AXYS[0][1] ),
    .X(net3749));
 sg13g2_dlygate4sd3_1 hold860 (.A(\scanline[106][2] ),
    .X(net3750));
 sg13g2_dlygate4sd3_1 hold861 (.A(\scanline[154][4] ),
    .X(net3751));
 sg13g2_dlygate4sd3_1 hold862 (.A(\scanline[53][5] ),
    .X(net3752));
 sg13g2_dlygate4sd3_1 hold863 (.A(\atari2600.tia.poly9_l.x[3] ),
    .X(net3753));
 sg13g2_dlygate4sd3_1 hold864 (.A(\atari2600.tia.audio_right_counter[11] ),
    .X(net3754));
 sg13g2_dlygate4sd3_1 hold865 (.A(_02039_),
    .X(net3755));
 sg13g2_dlygate4sd3_1 hold866 (.A(\scanline[47][3] ),
    .X(net3756));
 sg13g2_dlygate4sd3_1 hold867 (.A(\atari2600.ram[91][1] ),
    .X(net3757));
 sg13g2_dlygate4sd3_1 hold868 (.A(\scanline[150][0] ),
    .X(net3758));
 sg13g2_dlygate4sd3_1 hold869 (.A(\atari2600.ram[58][3] ),
    .X(net3759));
 sg13g2_dlygate4sd3_1 hold870 (.A(\atari2600.ram[3][7] ),
    .X(net3760));
 sg13g2_dlygate4sd3_1 hold871 (.A(\g_pwm_even[1] ),
    .X(net3761));
 sg13g2_dlygate4sd3_1 hold872 (.A(_04641_),
    .X(net3762));
 sg13g2_dlygate4sd3_1 hold873 (.A(_01192_),
    .X(net3763));
 sg13g2_dlygate4sd3_1 hold874 (.A(\atari2600.ram[94][4] ),
    .X(net3764));
 sg13g2_dlygate4sd3_1 hold875 (.A(\scanline[53][4] ),
    .X(net3765));
 sg13g2_dlygate4sd3_1 hold876 (.A(\atari2600.ram[89][1] ),
    .X(net3766));
 sg13g2_dlygate4sd3_1 hold877 (.A(\scanline[99][6] ),
    .X(net3767));
 sg13g2_dlygate4sd3_1 hold878 (.A(\scanline[121][4] ),
    .X(net3768));
 sg13g2_dlygate4sd3_1 hold879 (.A(\scanline[83][1] ),
    .X(net3769));
 sg13g2_dlygate4sd3_1 hold880 (.A(\scanline[157][4] ),
    .X(net3770));
 sg13g2_dlygate4sd3_1 hold881 (.A(_00669_),
    .X(net3771));
 sg13g2_dlygate4sd3_1 hold882 (.A(\atari2600.ram[30][3] ),
    .X(net3772));
 sg13g2_dlygate4sd3_1 hold883 (.A(\atari2600.ram[22][3] ),
    .X(net3773));
 sg13g2_dlygate4sd3_1 hold884 (.A(\scanline[94][3] ),
    .X(net3774));
 sg13g2_dlygate4sd3_1 hold885 (.A(\atari2600.ram[42][6] ),
    .X(net3775));
 sg13g2_dlygate4sd3_1 hold886 (.A(\scanline[143][5] ),
    .X(net3776));
 sg13g2_dlygate4sd3_1 hold887 (.A(\atari2600.cpu.AXYS[3][0] ),
    .X(net3777));
 sg13g2_dlygate4sd3_1 hold888 (.A(\atari2600.ram[114][4] ),
    .X(net3778));
 sg13g2_dlygate4sd3_1 hold889 (.A(\scanline[155][1] ),
    .X(net3779));
 sg13g2_dlygate4sd3_1 hold890 (.A(\atari2600.ram[42][3] ),
    .X(net3780));
 sg13g2_dlygate4sd3_1 hold891 (.A(\atari2600.ram[126][6] ),
    .X(net3781));
 sg13g2_dlygate4sd3_1 hold892 (.A(\scanline[47][4] ),
    .X(net3782));
 sg13g2_dlygate4sd3_1 hold893 (.A(\scanline[103][1] ),
    .X(net3783));
 sg13g2_dlygate4sd3_1 hold894 (.A(\scanline[83][5] ),
    .X(net3784));
 sg13g2_dlygate4sd3_1 hold895 (.A(\scanline[45][3] ),
    .X(net3785));
 sg13g2_dlygate4sd3_1 hold896 (.A(\atari2600.ram[76][0] ),
    .X(net3786));
 sg13g2_dlygate4sd3_1 hold897 (.A(\scanline[54][3] ),
    .X(net3787));
 sg13g2_dlygate4sd3_1 hold898 (.A(\atari2600.tia.pf_priority ),
    .X(net3788));
 sg13g2_dlygate4sd3_1 hold899 (.A(\scanline[93][5] ),
    .X(net3789));
 sg13g2_dlygate4sd3_1 hold900 (.A(\scanline[118][2] ),
    .X(net3790));
 sg13g2_dlygate4sd3_1 hold901 (.A(\scanline[85][6] ),
    .X(net3791));
 sg13g2_dlygate4sd3_1 hold902 (.A(\scanline[87][0] ),
    .X(net3792));
 sg13g2_dlygate4sd3_1 hold903 (.A(\atari2600.ram[38][4] ),
    .X(net3793));
 sg13g2_dlygate4sd3_1 hold904 (.A(\atari2600.pia.time_counter[14] ),
    .X(net3794));
 sg13g2_dlygate4sd3_1 hold905 (.A(_05329_),
    .X(net3795));
 sg13g2_dlygate4sd3_1 hold906 (.A(_01786_),
    .X(net3796));
 sg13g2_dlygate4sd3_1 hold907 (.A(\atari2600.ram[2][4] ),
    .X(net3797));
 sg13g2_dlygate4sd3_1 hold908 (.A(\atari2600.ram[46][1] ),
    .X(net3798));
 sg13g2_dlygate4sd3_1 hold909 (.A(\scanline[141][0] ),
    .X(net3799));
 sg13g2_dlygate4sd3_1 hold910 (.A(\atari2600.ram[22][0] ),
    .X(net3800));
 sg13g2_dlygate4sd3_1 hold911 (.A(\atari2600.tia.poly9_l.x[1] ),
    .X(net3801));
 sg13g2_dlygate4sd3_1 hold912 (.A(_02232_),
    .X(net3802));
 sg13g2_dlygate4sd3_1 hold913 (.A(\scanline[77][0] ),
    .X(net3803));
 sg13g2_dlygate4sd3_1 hold914 (.A(\atari2600.cpu.AXYS[2][0] ),
    .X(net3804));
 sg13g2_dlygate4sd3_1 hold915 (.A(\atari2600.tia.audio_left_counter[10] ),
    .X(net3805));
 sg13g2_dlygate4sd3_1 hold916 (.A(_02022_),
    .X(net3806));
 sg13g2_dlygate4sd3_1 hold917 (.A(\atari2600.ram[10][0] ),
    .X(net3807));
 sg13g2_dlygate4sd3_1 hold918 (.A(\atari2600.tia.cx[3] ),
    .X(net3808));
 sg13g2_dlygate4sd3_1 hold919 (.A(\scanline[79][6] ),
    .X(net3809));
 sg13g2_dlygate4sd3_1 hold920 (.A(\atari2600.ram[42][7] ),
    .X(net3810));
 sg13g2_dlygate4sd3_1 hold921 (.A(\atari2600.ram[82][5] ),
    .X(net3811));
 sg13g2_dlygate4sd3_1 hold922 (.A(\atari2600.ram[118][7] ),
    .X(net3812));
 sg13g2_dlygate4sd3_1 hold923 (.A(\scanline[89][5] ),
    .X(net3813));
 sg13g2_dlygate4sd3_1 hold924 (.A(\scanline[149][6] ),
    .X(net3814));
 sg13g2_dlygate4sd3_1 hold925 (.A(\atari2600.ram[94][6] ),
    .X(net3815));
 sg13g2_dlygate4sd3_1 hold926 (.A(\scanline[149][4] ),
    .X(net3816));
 sg13g2_dlygate4sd3_1 hold927 (.A(\atari2600.ram[82][7] ),
    .X(net3817));
 sg13g2_dlygate4sd3_1 hold928 (.A(\scanline[110][6] ),
    .X(net3818));
 sg13g2_dlygate4sd3_1 hold929 (.A(\scanline[46][5] ),
    .X(net3819));
 sg13g2_dlygate4sd3_1 hold930 (.A(\scanline[51][2] ),
    .X(net3820));
 sg13g2_dlygate4sd3_1 hold931 (.A(\scanline[61][4] ),
    .X(net3821));
 sg13g2_dlygate4sd3_1 hold932 (.A(_00059_),
    .X(net3822));
 sg13g2_dlygate4sd3_1 hold933 (.A(_04871_),
    .X(net3823));
 sg13g2_dlygate4sd3_1 hold934 (.A(\atari2600.ram[18][0] ),
    .X(net3824));
 sg13g2_dlygate4sd3_1 hold935 (.A(\atari2600.ram[73][5] ),
    .X(net3825));
 sg13g2_dlygate4sd3_1 hold936 (.A(\scanline[107][1] ),
    .X(net3826));
 sg13g2_dlygate4sd3_1 hold937 (.A(\scanline[147][1] ),
    .X(net3827));
 sg13g2_dlygate4sd3_1 hold938 (.A(\scanline[111][0] ),
    .X(net3828));
 sg13g2_dlygate4sd3_1 hold939 (.A(\atari2600.pia.diag[4] ),
    .X(net3829));
 sg13g2_dlygate4sd3_1 hold940 (.A(_01759_),
    .X(net3830));
 sg13g2_dlygate4sd3_1 hold941 (.A(\scanline[59][4] ),
    .X(net3831));
 sg13g2_dlygate4sd3_1 hold942 (.A(\scanline[122][4] ),
    .X(net3832));
 sg13g2_dlygate4sd3_1 hold943 (.A(\atari2600.ram[78][1] ),
    .X(net3833));
 sg13g2_dlygate4sd3_1 hold944 (.A(\scanline[150][2] ),
    .X(net3834));
 sg13g2_dlygate4sd3_1 hold945 (.A(\atari2600.ram[6][4] ),
    .X(net3835));
 sg13g2_dlygate4sd3_1 hold946 (.A(\scanline[93][2] ),
    .X(net3836));
 sg13g2_dlygate4sd3_1 hold947 (.A(\atari2600.ram[74][2] ),
    .X(net3837));
 sg13g2_dlygate4sd3_1 hold948 (.A(\atari2600.tia.audio_right_counter[3] ),
    .X(net3838));
 sg13g2_dlygate4sd3_1 hold949 (.A(_02031_),
    .X(net3839));
 sg13g2_dlygate4sd3_1 hold950 (.A(\atari2600.ram[118][2] ),
    .X(net3840));
 sg13g2_dlygate4sd3_1 hold951 (.A(\scanline[150][5] ),
    .X(net3841));
 sg13g2_dlygate4sd3_1 hold952 (.A(\scanline[31][2] ),
    .X(net3842));
 sg13g2_dlygate4sd3_1 hold953 (.A(\scanline[31][6] ),
    .X(net3843));
 sg13g2_dlygate4sd3_1 hold954 (.A(\atari2600.ram[82][3] ),
    .X(net3844));
 sg13g2_dlygate4sd3_1 hold955 (.A(\atari2600.pia.swb_dir[5] ),
    .X(net3845));
 sg13g2_dlygate4sd3_1 hold956 (.A(\flash_rom.addr[11] ),
    .X(net3846));
 sg13g2_dlygate4sd3_1 hold957 (.A(_01923_),
    .X(net3847));
 sg13g2_dlygate4sd3_1 hold958 (.A(\scanline[47][6] ),
    .X(net3848));
 sg13g2_dlygate4sd3_1 hold959 (.A(\atari2600.ram[6][3] ),
    .X(net3849));
 sg13g2_dlygate4sd3_1 hold960 (.A(\scanline[154][1] ),
    .X(net3850));
 sg13g2_dlygate4sd3_1 hold961 (.A(\atari2600.ram[90][0] ),
    .X(net3851));
 sg13g2_dlygate4sd3_1 hold962 (.A(\scanline[103][3] ),
    .X(net3852));
 sg13g2_dlygate4sd3_1 hold963 (.A(\atari2600.ram[79][6] ),
    .X(net3853));
 sg13g2_dlygate4sd3_1 hold964 (.A(\atari2600.ram[122][1] ),
    .X(net3854));
 sg13g2_dlygate4sd3_1 hold965 (.A(\atari2600.ram[74][5] ),
    .X(net3855));
 sg13g2_dlygate4sd3_1 hold966 (.A(\atari2600.tia.audio_right_counter[13] ),
    .X(net3856));
 sg13g2_dlygate4sd3_1 hold967 (.A(_02041_),
    .X(net3857));
 sg13g2_dlygate4sd3_1 hold968 (.A(\atari2600.cpu.src_reg[0] ),
    .X(net3858));
 sg13g2_dlygate4sd3_1 hold969 (.A(\atari2600.ram[126][7] ),
    .X(net3859));
 sg13g2_dlygate4sd3_1 hold970 (.A(\scanline[94][6] ),
    .X(net3860));
 sg13g2_dlygate4sd3_1 hold971 (.A(\atari2600.ram[76][4] ),
    .X(net3861));
 sg13g2_dlygate4sd3_1 hold972 (.A(\scanline[85][3] ),
    .X(net3862));
 sg13g2_dlygate4sd3_1 hold973 (.A(\atari2600.ram[26][4] ),
    .X(net3863));
 sg13g2_dlygate4sd3_1 hold974 (.A(\scanline[157][1] ),
    .X(net3864));
 sg13g2_dlygate4sd3_1 hold975 (.A(\atari2600.tia.poly4_l.x[1] ),
    .X(net3865));
 sg13g2_dlygate4sd3_1 hold976 (.A(\scanline[143][2] ),
    .X(net3866));
 sg13g2_dlygate4sd3_1 hold977 (.A(\scanline[154][6] ),
    .X(net3867));
 sg13g2_dlygate4sd3_1 hold978 (.A(\atari2600.ram[75][3] ),
    .X(net3868));
 sg13g2_dlygate4sd3_1 hold979 (.A(\atari2600.ram[3][5] ),
    .X(net3869));
 sg13g2_dlygate4sd3_1 hold980 (.A(\atari2600.pia.time_counter[9] ),
    .X(net3870));
 sg13g2_dlygate4sd3_1 hold981 (.A(_05316_),
    .X(net3871));
 sg13g2_dlygate4sd3_1 hold982 (.A(_01781_),
    .X(net3872));
 sg13g2_dlygate4sd3_1 hold983 (.A(\scanline[154][5] ),
    .X(net3873));
 sg13g2_dlygate4sd3_1 hold984 (.A(\scanline[62][0] ),
    .X(net3874));
 sg13g2_dlygate4sd3_1 hold985 (.A(\atari2600.ram[46][7] ),
    .X(net3875));
 sg13g2_dlygate4sd3_1 hold986 (.A(\atari2600.ram[98][6] ),
    .X(net3876));
 sg13g2_dlygate4sd3_1 hold987 (.A(\scanline[95][6] ),
    .X(net3877));
 sg13g2_dlygate4sd3_1 hold988 (.A(\atari2600.ram[82][0] ),
    .X(net3878));
 sg13g2_dlygate4sd3_1 hold989 (.A(\atari2600.ram[75][5] ),
    .X(net3879));
 sg13g2_dlygate4sd3_1 hold990 (.A(\atari2600.ram[86][6] ),
    .X(net3880));
 sg13g2_dlygate4sd3_1 hold991 (.A(\scanline[101][2] ),
    .X(net3881));
 sg13g2_dlygate4sd3_1 hold992 (.A(\scanline[62][4] ),
    .X(net3882));
 sg13g2_dlygate4sd3_1 hold993 (.A(\atari2600.pia.time_counter[6] ),
    .X(net3883));
 sg13g2_dlygate4sd3_1 hold994 (.A(_05311_),
    .X(net3884));
 sg13g2_dlygate4sd3_1 hold995 (.A(\scanline[122][1] ),
    .X(net3885));
 sg13g2_dlygate4sd3_1 hold996 (.A(\scanline[46][4] ),
    .X(net3886));
 sg13g2_dlygate4sd3_1 hold997 (.A(_00061_),
    .X(net3887));
 sg13g2_dlygate4sd3_1 hold998 (.A(_04863_),
    .X(net3888));
 sg13g2_dlygate4sd3_1 hold999 (.A(\atari2600.ram[106][4] ),
    .X(net3889));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\atari2600.ram[26][3] ),
    .X(net3890));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\scanline[51][3] ),
    .X(net3891));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\scanline[54][5] ),
    .X(net3892));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\atari2600.tia.audv1[2] ),
    .X(net3893));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\scanline[102][4] ),
    .X(net3894));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\atari2600.ram[122][5] ),
    .X(net3895));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\scanline[85][1] ),
    .X(net3896));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\atari2600.ram[89][7] ),
    .X(net3897));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\atari2600.ram[26][1] ),
    .X(net3898));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\atari2600.ram[2][0] ),
    .X(net3899));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\atari2600.ram[90][6] ),
    .X(net3900));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\atari2600.ram[10][2] ),
    .X(net3901));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\scanline[123][2] ),
    .X(net3902));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\scanline[57][5] ),
    .X(net3903));
 sg13g2_dlygate4sd3_1 hold1014 (.A(\scanline[142][5] ),
    .X(net3904));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\atari2600.tia.audio_left_counter[9] ),
    .X(net3905));
 sg13g2_dlygate4sd3_1 hold1016 (.A(_05928_),
    .X(net3906));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\scanline[47][2] ),
    .X(net3907));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\atari2600.cpu.ABL[5] ),
    .X(net3908));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\atari2600.ram[118][4] ),
    .X(net3909));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\scanline[91][5] ),
    .X(net3910));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\scanline[149][3] ),
    .X(net3911));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\atari2600.ram[77][1] ),
    .X(net3912));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\atari2600.tia.poly5_l.x[3] ),
    .X(net3913));
 sg13g2_dlygate4sd3_1 hold1024 (.A(_02230_),
    .X(net3914));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\atari2600.ram[3][3] ),
    .X(net3915));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\atari2600.pia.swa_dir[4] ),
    .X(net3916));
 sg13g2_dlygate4sd3_1 hold1027 (.A(\scanline[14][0] ),
    .X(net3917));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\atari2600.ram[79][5] ),
    .X(net3918));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\scanline[30][0] ),
    .X(net3919));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\atari2600.pia.swa_dir[1] ),
    .X(net3920));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\atari2600.ram[46][5] ),
    .X(net3921));
 sg13g2_dlygate4sd3_1 hold1032 (.A(\scanline[123][5] ),
    .X(net3922));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\atari2600.cpu.AXYS[2][1] ),
    .X(net3923));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\scanline[147][3] ),
    .X(net3924));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\scanline[150][1] ),
    .X(net3925));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\atari2600.tia.audio_right_counter[7] ),
    .X(net3926));
 sg13g2_dlygate4sd3_1 hold1037 (.A(_02035_),
    .X(net3927));
 sg13g2_dlygate4sd3_1 hold1038 (.A(\atari2600.ram[18][3] ),
    .X(net3928));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\scanline[107][0] ),
    .X(net3929));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\atari2600.tia.poly5_l.x[2] ),
    .X(net3930));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\atari2600.cpu.Z ),
    .X(net3931));
 sg13g2_dlygate4sd3_1 hold1042 (.A(_07288_),
    .X(net3932));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\atari2600.tia.audio_left_counter[2] ),
    .X(net3933));
 sg13g2_dlygate4sd3_1 hold1044 (.A(_02014_),
    .X(net3934));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\scanline[158][3] ),
    .X(net3935));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\scanline[106][1] ),
    .X(net3936));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\scanline[31][4] ),
    .X(net3937));
 sg13g2_dlygate4sd3_1 hold1048 (.A(\scanline[153][5] ),
    .X(net3938));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\scanline[62][5] ),
    .X(net3939));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\scanline[122][5] ),
    .X(net3940));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\atari2600.pia.swa_dir[0] ),
    .X(net3941));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\atari2600.tia.poly9_l.x[8] ),
    .X(net3942));
 sg13g2_dlygate4sd3_1 hold1053 (.A(_02239_),
    .X(net3943));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\scanline[121][5] ),
    .X(net3944));
 sg13g2_dlygate4sd3_1 hold1055 (.A(\scanline[103][0] ),
    .X(net3945));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\atari2600.ram[6][1] ),
    .X(net3946));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\atari2600.ram[91][6] ),
    .X(net3947));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\scanline[158][6] ),
    .X(net3948));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\scanline[77][4] ),
    .X(net3949));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\scanline[99][3] ),
    .X(net3950));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\atari2600.ram[102][3] ),
    .X(net3951));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\flash_rom.addr[15] ),
    .X(net3952));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\atari2600.ram[86][3] ),
    .X(net3953));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\scanline[78][6] ),
    .X(net3954));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\atari2600.tia.cx[0] ),
    .X(net3955));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\scanline[83][6] ),
    .X(net3956));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\atari2600.ram[73][2] ),
    .X(net3957));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\atari2600.rom_data[3] ),
    .X(net3958));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\atari2600.tia.diag[103] ),
    .X(net3959));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\atari2600.ram[58][5] ),
    .X(net3960));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\scanline[130][3] ),
    .X(net3961));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\scanline[106][5] ),
    .X(net3962));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\atari2600.ram[62][3] ),
    .X(net3963));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\scanline[143][3] ),
    .X(net3964));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\atari2600.rom_data[6] ),
    .X(net3965));
 sg13g2_dlygate4sd3_1 hold1076 (.A(_02926_),
    .X(net3966));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\atari2600.ram[95][5] ),
    .X(net3967));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\atari2600.ram[94][3] ),
    .X(net3968));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\atari2600.ram[2][2] ),
    .X(net3969));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\atari2600.cpu.clc ),
    .X(net3970));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\atari2600.ram[30][4] ),
    .X(net3971));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\atari2600.cpu.load_reg ),
    .X(net3972));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\scanline[126][1] ),
    .X(net3973));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\rom_last_read_addr[4] ),
    .X(net3974));
 sg13g2_dlygate4sd3_1 hold1085 (.A(_01130_),
    .X(net3975));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\atari2600.ram[98][3] ),
    .X(net3976));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\rom_last_read_addr[5] ),
    .X(net3977));
 sg13g2_dlygate4sd3_1 hold1088 (.A(_01131_),
    .X(net3978));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\atari2600.ram[126][0] ),
    .X(net3979));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\scanline[13][0] ),
    .X(net3980));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\atari2600.cpu.op[3] ),
    .X(net3981));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\atari2600.tia.audio_right_counter[9] ),
    .X(net3982));
 sg13g2_dlygate4sd3_1 hold1093 (.A(_02037_),
    .X(net3983));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\atari2600.ram[38][5] ),
    .X(net3984));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\atari2600.ram[53][1] ),
    .X(net3985));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\atari2600.ram[70][3] ),
    .X(net3986));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\atari2600.pia.dat_o[1] ),
    .X(net3987));
 sg13g2_dlygate4sd3_1 hold1098 (.A(_01765_),
    .X(net3988));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\atari2600.cpu.op[2] ),
    .X(net3989));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\atari2600.pia.swa_dir[7] ),
    .X(net3990));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\scanline[159][1] ),
    .X(net3991));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\atari2600.tia.audio_left_counter[6] ),
    .X(net3992));
 sg13g2_dlygate4sd3_1 hold1103 (.A(_02018_),
    .X(net3993));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\atari2600.ram[62][7] ),
    .X(net3994));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\scanline[47][0] ),
    .X(net3995));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\atari2600.ram[29][3] ),
    .X(net3996));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\scanline[117][2] ),
    .X(net3997));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\atari2600.ram[106][1] ),
    .X(net3998));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\scanline[106][4] ),
    .X(net3999));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\atari2600.ram[113][1] ),
    .X(net4000));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\atari2600.ram[10][5] ),
    .X(net4001));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\scanline[111][6] ),
    .X(net4002));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\atari2600.ram[110][7] ),
    .X(net4003));
 sg13g2_dlygate4sd3_1 hold1114 (.A(\scanline[54][2] ),
    .X(net4004));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\atari2600.ram[18][7] ),
    .X(net4005));
 sg13g2_dlygate4sd3_1 hold1116 (.A(\atari2600.ram[101][0] ),
    .X(net4006));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\atari2600.tia.audio_right_counter[14] ),
    .X(net4007));
 sg13g2_dlygate4sd3_1 hold1118 (.A(_02042_),
    .X(net4008));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\flash_rom.addr[17] ),
    .X(net4009));
 sg13g2_dlygate4sd3_1 hold1120 (.A(_00213_),
    .X(net4010));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\atari2600.ram[61][5] ),
    .X(net4011));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\atari2600.ram[24][5] ),
    .X(net4012));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\atari2600.ram[125][1] ),
    .X(net4013));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\atari2600.tia.diag[110] ),
    .X(net4014));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\scanline[58][5] ),
    .X(net4015));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\atari2600.ram[55][1] ),
    .X(net4016));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\atari2600.ram[8][6] ),
    .X(net4017));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\atari2600.ram[41][1] ),
    .X(net4018));
 sg13g2_dlygate4sd3_1 hold1129 (.A(\atari2600.pia.dat_o[0] ),
    .X(net4019));
 sg13g2_dlygate4sd3_1 hold1130 (.A(_01764_),
    .X(net4020));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\atari2600.ram[45][0] ),
    .X(net4021));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\atari2600.pia.time_counter[11] ),
    .X(net4022));
 sg13g2_dlygate4sd3_1 hold1133 (.A(_05322_),
    .X(net4023));
 sg13g2_dlygate4sd3_1 hold1134 (.A(_01783_),
    .X(net4024));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\atari2600.ram[55][3] ),
    .X(net4025));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\atari2600.ram[1][3] ),
    .X(net4026));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\atari2600.ram[25][5] ),
    .X(net4027));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\atari2600.ram[45][4] ),
    .X(net4028));
 sg13g2_dlygate4sd3_1 hold1139 (.A(\scanline[113][3] ),
    .X(net4029));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\atari2600.ram[49][4] ),
    .X(net4030));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\atari2600.ram[12][2] ),
    .X(net4031));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\scanline[91][0] ),
    .X(net4032));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\atari2600.ram[44][3] ),
    .X(net4033));
 sg13g2_dlygate4sd3_1 hold1144 (.A(\atari2600.ram[5][0] ),
    .X(net4034));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\atari2600.ram[49][3] ),
    .X(net4035));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\scanline[157][3] ),
    .X(net4036));
 sg13g2_dlygate4sd3_1 hold1147 (.A(\atari2600.ram[21][6] ),
    .X(net4037));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\atari2600.ram[29][5] ),
    .X(net4038));
 sg13g2_dlygate4sd3_1 hold1149 (.A(\atari2600.ram[0][5] ),
    .X(net4039));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\atari2600.ram[84][4] ),
    .X(net4040));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\atari2600.ram[97][7] ),
    .X(net4041));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\atari2600.ram[49][7] ),
    .X(net4042));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\atari2600.ram[60][0] ),
    .X(net4043));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\atari2600.ram[121][5] ),
    .X(net4044));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\atari2600.ram[61][1] ),
    .X(net4045));
 sg13g2_dlygate4sd3_1 hold1156 (.A(\atari2600.ram[95][0] ),
    .X(net4046));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\atari2600.ram[109][7] ),
    .X(net4047));
 sg13g2_dlygate4sd3_1 hold1158 (.A(\atari2600.ram[34][0] ),
    .X(net4048));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\atari2600.ram[126][3] ),
    .X(net4049));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\atari2600.ram[121][7] ),
    .X(net4050));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\atari2600.ram[24][7] ),
    .X(net4051));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\atari2600.ram[69][2] ),
    .X(net4052));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\atari2600.ram[26][5] ),
    .X(net4053));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\atari2600.ram[69][7] ),
    .X(net4054));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\atari2600.ram[81][7] ),
    .X(net4055));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\atari2600.ram[53][3] ),
    .X(net4056));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\atari2600.ram[114][7] ),
    .X(net4057));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\atari2600.cpu.PC[9] ),
    .X(net4058));
 sg13g2_dlygate4sd3_1 hold1169 (.A(_02507_),
    .X(net4059));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\atari2600.ram[119][1] ),
    .X(net4060));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\scanline[147][2] ),
    .X(net4061));
 sg13g2_dlygate4sd3_1 hold1172 (.A(\atari2600.ram[100][6] ),
    .X(net4062));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\atari2600.ram[105][7] ),
    .X(net4063));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\atari2600.ram[50][2] ),
    .X(net4064));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\atari2600.ram[32][4] ),
    .X(net4065));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\flash_rom.addr[10] ),
    .X(net4066));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\atari2600.ram[68][5] ),
    .X(net4067));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\atari2600.ram[45][3] ),
    .X(net4068));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\atari2600.ram[45][5] ),
    .X(net4069));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\atari2600.ram[125][3] ),
    .X(net4070));
 sg13g2_dlygate4sd3_1 hold1181 (.A(\atari2600.ram[108][7] ),
    .X(net4071));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\atari2600.ram[41][0] ),
    .X(net4072));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\atari2600.tia.diag[99] ),
    .X(net4073));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\atari2600.ram[108][0] ),
    .X(net4074));
 sg13g2_dlygate4sd3_1 hold1185 (.A(\scanline[51][4] ),
    .X(net4075));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\atari2600.ram[20][1] ),
    .X(net4076));
 sg13g2_dlygate4sd3_1 hold1187 (.A(\atari2600.ram[113][4] ),
    .X(net4077));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\atari2600.ram[121][6] ),
    .X(net4078));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\atari2600.ram[28][3] ),
    .X(net4079));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\atari2600.ram[21][5] ),
    .X(net4080));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\atari2600.ram[17][2] ),
    .X(net4081));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\atari2600.ram[48][7] ),
    .X(net4082));
 sg13g2_dlygate4sd3_1 hold1193 (.A(\atari2600.ram[49][0] ),
    .X(net4083));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\atari2600.ram[117][0] ),
    .X(net4084));
 sg13g2_dlygate4sd3_1 hold1195 (.A(\atari2600.ram[21][2] ),
    .X(net4085));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\atari2600.ram[64][0] ),
    .X(net4086));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\atari2600.ram[96][4] ),
    .X(net4087));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\atari2600.tia.diag[102] ),
    .X(net4088));
 sg13g2_dlygate4sd3_1 hold1199 (.A(\atari2600.cpu.N ),
    .X(net4089));
 sg13g2_dlygate4sd3_1 hold1200 (.A(_02468_),
    .X(net4090));
 sg13g2_dlygate4sd3_1 hold1201 (.A(\atari2600.ram[0][2] ),
    .X(net4091));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\atari2600.ram[104][2] ),
    .X(net4092));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\atari2600.ram[109][2] ),
    .X(net4093));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\scanline[149][0] ),
    .X(net4094));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\atari2600.ram[28][0] ),
    .X(net4095));
 sg13g2_dlygate4sd3_1 hold1206 (.A(\atari2600.ram[50][0] ),
    .X(net4096));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\atari2600.ram[64][1] ),
    .X(net4097));
 sg13g2_dlygate4sd3_1 hold1208 (.A(\atari2600.tia.poly9_l.x[4] ),
    .X(net4098));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\atari2600.ram[84][3] ),
    .X(net4099));
 sg13g2_dlygate4sd3_1 hold1210 (.A(\atari2600.ram[25][2] ),
    .X(net4100));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\atari2600.ram[48][4] ),
    .X(net4101));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\atari2600.cpu.sec ),
    .X(net4102));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\atari2600.ram[100][4] ),
    .X(net4103));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\scanline[125][1] ),
    .X(net4104));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\atari2600.tia.refp1 ),
    .X(net4105));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\atari2600.ram[61][7] ),
    .X(net4106));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\atari2600.ram[45][7] ),
    .X(net4107));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\atari2600.ram[44][7] ),
    .X(net4108));
 sg13g2_dlygate4sd3_1 hold1219 (.A(\atari2600.cpu.AXYS[3][5] ),
    .X(net4109));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\atari2600.ram[104][6] ),
    .X(net4110));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\atari2600.ram[100][3] ),
    .X(net4111));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\atari2600.cpu.AXYS[0][3] ),
    .X(net4112));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\atari2600.ram[52][0] ),
    .X(net4113));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\atari2600.ram[85][2] ),
    .X(net4114));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\atari2600.ram[9][1] ),
    .X(net4115));
 sg13g2_dlygate4sd3_1 hold1226 (.A(\atari2600.ram[69][0] ),
    .X(net4116));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\atari2600.ram[96][7] ),
    .X(net4117));
 sg13g2_dlygate4sd3_1 hold1228 (.A(\atari2600.ram[65][0] ),
    .X(net4118));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\atari2600.tia.poly9_l.x[5] ),
    .X(net4119));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\atari2600.ram[113][6] ),
    .X(net4120));
 sg13g2_dlygate4sd3_1 hold1231 (.A(\atari2600.ram[28][6] ),
    .X(net4121));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\atari2600.ram[56][7] ),
    .X(net4122));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\atari2600.ram[124][3] ),
    .X(net4123));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\atari2600.ram[20][6] ),
    .X(net4124));
 sg13g2_dlygate4sd3_1 hold1235 (.A(\atari2600.ram[44][1] ),
    .X(net4125));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\atari2600.cpu.ABL[7] ),
    .X(net4126));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\atari2600.ram[8][4] ),
    .X(net4127));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\atari2600.ram[57][3] ),
    .X(net4128));
 sg13g2_dlygate4sd3_1 hold1239 (.A(\atari2600.ram[20][2] ),
    .X(net4129));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\atari2600.ram[49][2] ),
    .X(net4130));
 sg13g2_dlygate4sd3_1 hold1241 (.A(\atari2600.ram[41][2] ),
    .X(net4131));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\atari2600.ram[116][1] ),
    .X(net4132));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\atari2600.ram[120][6] ),
    .X(net4133));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\scanline[120][0] ),
    .X(net4134));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\atari2600.tia.audio_right_counter[5] ),
    .X(net4135));
 sg13g2_dlygate4sd3_1 hold1246 (.A(_02033_),
    .X(net4136));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\atari2600.ram[109][5] ),
    .X(net4137));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\atari2600.ram[105][3] ),
    .X(net4138));
 sg13g2_dlygate4sd3_1 hold1249 (.A(\atari2600.ram[68][3] ),
    .X(net4139));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\atari2600.ram[48][2] ),
    .X(net4140));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\atari2600.ram[98][5] ),
    .X(net4141));
 sg13g2_dlygate4sd3_1 hold1252 (.A(\atari2600.ram[85][0] ),
    .X(net4142));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\atari2600.tia.colup0[1] ),
    .X(net4143));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\atari2600.ram[0][3] ),
    .X(net4144));
 sg13g2_dlygate4sd3_1 hold1255 (.A(\atari2600.ram[20][0] ),
    .X(net4145));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\atari2600.cpu.I ),
    .X(net4146));
 sg13g2_dlygate4sd3_1 hold1257 (.A(_07261_),
    .X(net4147));
 sg13g2_dlygate4sd3_1 hold1258 (.A(_02466_),
    .X(net4148));
 sg13g2_dlygate4sd3_1 hold1259 (.A(\atari2600.ram[48][6] ),
    .X(net4149));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\atari2600.ram[9][6] ),
    .X(net4150));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\atari2600.ram[61][2] ),
    .X(net4151));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\atari2600.ram[5][2] ),
    .X(net4152));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\atari2600.ram[108][1] ),
    .X(net4153));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\atari2600.ram[29][2] ),
    .X(net4154));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\atari2600.ram[81][3] ),
    .X(net4155));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\atari2600.ram[40][6] ),
    .X(net4156));
 sg13g2_dlygate4sd3_1 hold1267 (.A(\atari2600.ram[32][7] ),
    .X(net4157));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\atari2600.ram[9][3] ),
    .X(net4158));
 sg13g2_dlygate4sd3_1 hold1269 (.A(\atari2600.ram[54][0] ),
    .X(net4159));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\atari2600.ram[103][5] ),
    .X(net4160));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\atari2600.ram[24][6] ),
    .X(net4161));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\atari2600.ram[16][7] ),
    .X(net4162));
 sg13g2_dlygate4sd3_1 hold1273 (.A(\atari2600.tia.diag[96] ),
    .X(net4163));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\scanline[76][1] ),
    .X(net4164));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\flash_rom.addr[12] ),
    .X(net4165));
 sg13g2_dlygate4sd3_1 hold1276 (.A(_01920_),
    .X(net4166));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\atari2600.ram[125][5] ),
    .X(net4167));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\atari2600.ram[117][3] ),
    .X(net4168));
 sg13g2_dlygate4sd3_1 hold1279 (.A(\scanline[68][6] ),
    .X(net4169));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\atari2600.ram[0][6] ),
    .X(net4170));
 sg13g2_dlygate4sd3_1 hold1281 (.A(\atari2600.ram[8][1] ),
    .X(net4171));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\scanline[70][6] ),
    .X(net4172));
 sg13g2_dlygate4sd3_1 hold1283 (.A(\atari2600.ram[112][3] ),
    .X(net4173));
 sg13g2_dlygate4sd3_1 hold1284 (.A(\atari2600.ram[5][1] ),
    .X(net4174));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\atari2600.ram[7][7] ),
    .X(net4175));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\atari2600.ram[113][2] ),
    .X(net4176));
 sg13g2_dlygate4sd3_1 hold1287 (.A(\atari2600.ram[4][5] ),
    .X(net4177));
 sg13g2_dlygate4sd3_1 hold1288 (.A(\atari2600.ram[120][0] ),
    .X(net4178));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\atari2600.pia.reset_timer[1] ),
    .X(net4179));
 sg13g2_dlygate4sd3_1 hold1290 (.A(\atari2600.pia.time_counter[17] ),
    .X(net4180));
 sg13g2_dlygate4sd3_1 hold1291 (.A(_05338_),
    .X(net4181));
 sg13g2_dlygate4sd3_1 hold1292 (.A(\atari2600.ram[11][7] ),
    .X(net4182));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\atari2600.ram[0][1] ),
    .X(net4183));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\atari2600.ram[24][0] ),
    .X(net4184));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\atari2600.ram[108][2] ),
    .X(net4185));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\atari2600.ram[108][4] ),
    .X(net4186));
 sg13g2_dlygate4sd3_1 hold1297 (.A(\atari2600.tia.poly9_l.x[6] ),
    .X(net4187));
 sg13g2_dlygate4sd3_1 hold1298 (.A(\atari2600.ram[45][2] ),
    .X(net4188));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\scanline[116][4] ),
    .X(net4189));
 sg13g2_dlygate4sd3_1 hold1300 (.A(\atari2600.ram[65][2] ),
    .X(net4190));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\atari2600.cpu.dst_reg[0] ),
    .X(net4191));
 sg13g2_dlygate4sd3_1 hold1302 (.A(\atari2600.ram[9][4] ),
    .X(net4192));
 sg13g2_dlygate4sd3_1 hold1303 (.A(\atari2600.ram[56][6] ),
    .X(net4193));
 sg13g2_dlygate4sd3_1 hold1304 (.A(\atari2600.ram[24][2] ),
    .X(net4194));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\atari2600.ram[8][5] ),
    .X(net4195));
 sg13g2_dlygate4sd3_1 hold1306 (.A(\atari2600.ram[24][4] ),
    .X(net4196));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\atari2600.ram[125][6] ),
    .X(net4197));
 sg13g2_dlygate4sd3_1 hold1308 (.A(\atari2600.ram[40][3] ),
    .X(net4198));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\scanline[120][4] ),
    .X(net4199));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\atari2600.ram[16][0] ),
    .X(net4200));
 sg13g2_dlygate4sd3_1 hold1311 (.A(\atari2600.ram[80][7] ),
    .X(net4201));
 sg13g2_dlygate4sd3_1 hold1312 (.A(\atari2600.ram[84][6] ),
    .X(net4202));
 sg13g2_dlygate4sd3_1 hold1313 (.A(\atari2600.ram[108][3] ),
    .X(net4203));
 sg13g2_dlygate4sd3_1 hold1314 (.A(\atari2600.ram[59][6] ),
    .X(net4204));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\atari2600.ram[97][3] ),
    .X(net4205));
 sg13g2_dlygate4sd3_1 hold1316 (.A(\scanline[4][2] ),
    .X(net4206));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\atari2600.ram[17][1] ),
    .X(net4207));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\atari2600.ram[53][5] ),
    .X(net4208));
 sg13g2_dlygate4sd3_1 hold1319 (.A(\atari2600.ram[112][6] ),
    .X(net4209));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\atari2600.ram[122][4] ),
    .X(net4210));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\atari2600.ram[86][5] ),
    .X(net4211));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\atari2600.ram[109][1] ),
    .X(net4212));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\atari2600.ram[109][3] ),
    .X(net4213));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\atari2600.ram[43][1] ),
    .X(net4214));
 sg13g2_dlygate4sd3_1 hold1325 (.A(\flash_rom.addr[21] ),
    .X(net4215));
 sg13g2_dlygate4sd3_1 hold1326 (.A(_10492_),
    .X(net4216));
 sg13g2_dlygate4sd3_1 hold1327 (.A(\atari2600.ram[80][5] ),
    .X(net4217));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\atari2600.ram[18][5] ),
    .X(net4218));
 sg13g2_dlygate4sd3_1 hold1329 (.A(\atari2600.ram[125][0] ),
    .X(net4219));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\atari2600.ram[85][3] ),
    .X(net4220));
 sg13g2_dlygate4sd3_1 hold1331 (.A(\flash_rom.addr[16] ),
    .X(net4221));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\scanline[80][4] ),
    .X(net4222));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\scanline[103][2] ),
    .X(net4223));
 sg13g2_dlygate4sd3_1 hold1334 (.A(\atari2600.tia.audv1[3] ),
    .X(net4224));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\atari2600.ram[101][5] ),
    .X(net4225));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\atari2600.ram[121][3] ),
    .X(net4226));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\atari2600.ram[127][2] ),
    .X(net4227));
 sg13g2_dlygate4sd3_1 hold1338 (.A(\atari2600.ram[39][3] ),
    .X(net4228));
 sg13g2_dlygate4sd3_1 hold1339 (.A(\atari2600.rom_data[1] ),
    .X(net4229));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\scanline[51][1] ),
    .X(net4230));
 sg13g2_dlygate4sd3_1 hold1341 (.A(\atari2600.cpu.AXYS[1][3] ),
    .X(net4231));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\scanline[137][3] ),
    .X(net4232));
 sg13g2_dlygate4sd3_1 hold1343 (.A(\atari2600.ram[5][7] ),
    .X(net4233));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\atari2600.ram[12][1] ),
    .X(net4234));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\atari2600.ram[25][1] ),
    .X(net4235));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\atari2600.ram[29][4] ),
    .X(net4236));
 sg13g2_dlygate4sd3_1 hold1347 (.A(\atari2600.ram[55][5] ),
    .X(net4237));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\atari2600.ram[39][4] ),
    .X(net4238));
 sg13g2_dlygate4sd3_1 hold1349 (.A(\atari2600.ram[32][2] ),
    .X(net4239));
 sg13g2_dlygate4sd3_1 hold1350 (.A(\atari2600.ram[64][6] ),
    .X(net4240));
 sg13g2_dlygate4sd3_1 hold1351 (.A(\atari2600.ram[45][6] ),
    .X(net4241));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\atari2600.ram[125][7] ),
    .X(net4242));
 sg13g2_dlygate4sd3_1 hold1353 (.A(\scanline[34][1] ),
    .X(net4243));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\scanline[17][1] ),
    .X(net4244));
 sg13g2_dlygate4sd3_1 hold1355 (.A(\atari2600.ram[119][5] ),
    .X(net4245));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\scanline[28][0] ),
    .X(net4246));
 sg13g2_dlygate4sd3_1 hold1357 (.A(\atari2600.ram[112][1] ),
    .X(net4247));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\atari2600.ram[120][1] ),
    .X(net4248));
 sg13g2_dlygate4sd3_1 hold1359 (.A(\atari2600.ram[107][3] ),
    .X(net4249));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\atari2600.ram[44][6] ),
    .X(net4250));
 sg13g2_dlygate4sd3_1 hold1361 (.A(\atari2600.ram[48][0] ),
    .X(net4251));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\atari2600.ram[123][1] ),
    .X(net4252));
 sg13g2_dlygate4sd3_1 hold1363 (.A(\atari2600.cpu.AXYS[1][6] ),
    .X(net4253));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\atari2600.ram[63][1] ),
    .X(net4254));
 sg13g2_dlygate4sd3_1 hold1365 (.A(\atari2600.ram[7][1] ),
    .X(net4255));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\atari2600.ram[120][2] ),
    .X(net4256));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\scanline[18][5] ),
    .X(net4257));
 sg13g2_dlygate4sd3_1 hold1368 (.A(\atari2600.ram[13][7] ),
    .X(net4258));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\atari2600.ram[84][7] ),
    .X(net4259));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\atari2600.ram[65][7] ),
    .X(net4260));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\atari2600.ram[120][7] ),
    .X(net4261));
 sg13g2_dlygate4sd3_1 hold1372 (.A(\scanline[137][0] ),
    .X(net4262));
 sg13g2_dlygate4sd3_1 hold1373 (.A(\atari2600.ram[39][7] ),
    .X(net4263));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\atari2600.ram[84][5] ),
    .X(net4264));
 sg13g2_dlygate4sd3_1 hold1375 (.A(\atari2600.ram[80][6] ),
    .X(net4265));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\atari2600.ram[71][5] ),
    .X(net4266));
 sg13g2_dlygate4sd3_1 hold1377 (.A(\scanline[76][4] ),
    .X(net4267));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\atari2600.ram[16][1] ),
    .X(net4268));
 sg13g2_dlygate4sd3_1 hold1379 (.A(\atari2600.ram[39][1] ),
    .X(net4269));
 sg13g2_dlygate4sd3_1 hold1380 (.A(\atari2600.ram[52][2] ),
    .X(net4270));
 sg13g2_dlygate4sd3_1 hold1381 (.A(\atari2600.ram[9][0] ),
    .X(net4271));
 sg13g2_dlygate4sd3_1 hold1382 (.A(\atari2600.ram[68][2] ),
    .X(net4272));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\atari2600.ram[96][1] ),
    .X(net4273));
 sg13g2_dlygate4sd3_1 hold1384 (.A(\atari2600.ram[69][1] ),
    .X(net4274));
 sg13g2_dlygate4sd3_1 hold1385 (.A(\atari2600.ram[27][2] ),
    .X(net4275));
 sg13g2_dlygate4sd3_1 hold1386 (.A(\atari2600.cpu.AXYS[1][7] ),
    .X(net4276));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\atari2600.ram[32][3] ),
    .X(net4277));
 sg13g2_dlygate4sd3_1 hold1388 (.A(\atari2600.tia.diag[98] ),
    .X(net4278));
 sg13g2_dlygate4sd3_1 hold1389 (.A(\atari2600.cpu.ABL[0] ),
    .X(net4279));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\scanline[136][0] ),
    .X(net4280));
 sg13g2_dlygate4sd3_1 hold1391 (.A(\atari2600.ram[44][5] ),
    .X(net4281));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\scanline[25][5] ),
    .X(net4282));
 sg13g2_dlygate4sd3_1 hold1393 (.A(\atari2600.cpu.AXYS[0][4] ),
    .X(net4283));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\scanline[34][0] ),
    .X(net4284));
 sg13g2_dlygate4sd3_1 hold1395 (.A(\atari2600.ram[35][2] ),
    .X(net4285));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\scanline[36][2] ),
    .X(net4286));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\atari2600.ram[34][7] ),
    .X(net4287));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\scanline[97][0] ),
    .X(net4288));
 sg13g2_dlygate4sd3_1 hold1399 (.A(\scanline[25][1] ),
    .X(net4289));
 sg13g2_dlygate4sd3_1 hold1400 (.A(\atari2600.ram[21][4] ),
    .X(net4290));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\atari2600.cpu.ABL[2] ),
    .X(net4291));
 sg13g2_dlygate4sd3_1 hold1402 (.A(_02481_),
    .X(net4292));
 sg13g2_dlygate4sd3_1 hold1403 (.A(\scanline[76][0] ),
    .X(net4293));
 sg13g2_dlygate4sd3_1 hold1404 (.A(\atari2600.ram[104][0] ),
    .X(net4294));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\atari2600.ram[35][1] ),
    .X(net4295));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\atari2600.ram[104][1] ),
    .X(net4296));
 sg13g2_dlygate4sd3_1 hold1407 (.A(\atari2600.ram[61][3] ),
    .X(net4297));
 sg13g2_dlygate4sd3_1 hold1408 (.A(\atari2600.ram[37][7] ),
    .X(net4298));
 sg13g2_dlygate4sd3_1 hold1409 (.A(\atari2600.ram[115][5] ),
    .X(net4299));
 sg13g2_dlygate4sd3_1 hold1410 (.A(\atari2600.ram[104][4] ),
    .X(net4300));
 sg13g2_dlygate4sd3_1 hold1411 (.A(\scanline[81][5] ),
    .X(net4301));
 sg13g2_dlygate4sd3_1 hold1412 (.A(\scanline[138][0] ),
    .X(net4302));
 sg13g2_dlygate4sd3_1 hold1413 (.A(\scanline[7][4] ),
    .X(net4303));
 sg13g2_dlygate4sd3_1 hold1414 (.A(\atari2600.ram[56][2] ),
    .X(net4304));
 sg13g2_dlygate4sd3_1 hold1415 (.A(\scanline[74][3] ),
    .X(net4305));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\atari2600.ram[55][7] ),
    .X(net4306));
 sg13g2_dlygate4sd3_1 hold1417 (.A(\scanline[144][4] ),
    .X(net4307));
 sg13g2_dlygate4sd3_1 hold1418 (.A(\scanline[81][6] ),
    .X(net4308));
 sg13g2_dlygate4sd3_1 hold1419 (.A(\atari2600.ram[56][5] ),
    .X(net4309));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\atari2600.ram[112][4] ),
    .X(net4310));
 sg13g2_dlygate4sd3_1 hold1421 (.A(\scanline[129][3] ),
    .X(net4311));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\atari2600.ram[57][1] ),
    .X(net4312));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\atari2600.cpu.AXYS[3][4] ),
    .X(net4313));
 sg13g2_dlygate4sd3_1 hold1424 (.A(\atari2600.ram[35][0] ),
    .X(net4314));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\atari2600.ram[49][1] ),
    .X(net4315));
 sg13g2_dlygate4sd3_1 hold1426 (.A(\atari2600.ram[120][4] ),
    .X(net4316));
 sg13g2_dlygate4sd3_1 hold1427 (.A(\atari2600.tia.diag[100] ),
    .X(net4317));
 sg13g2_dlygate4sd3_1 hold1428 (.A(_01824_),
    .X(net4318));
 sg13g2_dlygate4sd3_1 hold1429 (.A(\scanline[100][4] ),
    .X(net4319));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\atari2600.ram[52][3] ),
    .X(net4320));
 sg13g2_dlygate4sd3_1 hold1431 (.A(\atari2600.ram[12][7] ),
    .X(net4321));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\scanline[6][1] ),
    .X(net4322));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\scanline[116][2] ),
    .X(net4323));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\atari2600.ram[12][4] ),
    .X(net4324));
 sg13g2_dlygate4sd3_1 hold1435 (.A(\atari2600.ram[24][3] ),
    .X(net4325));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\atari2600.ram[56][0] ),
    .X(net4326));
 sg13g2_dlygate4sd3_1 hold1437 (.A(\atari2600.ram[101][6] ),
    .X(net4327));
 sg13g2_dlygate4sd3_1 hold1438 (.A(\scanline[56][0] ),
    .X(net4328));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\scanline[21][0] ),
    .X(net4329));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\scanline[21][2] ),
    .X(net4330));
 sg13g2_dlygate4sd3_1 hold1441 (.A(\atari2600.ram[102][4] ),
    .X(net4331));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\atari2600.ram[87][0] ),
    .X(net4332));
 sg13g2_dlygate4sd3_1 hold1443 (.A(\atari2600.ram[102][6] ),
    .X(net4333));
 sg13g2_dlygate4sd3_1 hold1444 (.A(\atari2600.ram[59][4] ),
    .X(net4334));
 sg13g2_dlygate4sd3_1 hold1445 (.A(\atari2600.ram[12][3] ),
    .X(net4335));
 sg13g2_dlygate4sd3_1 hold1446 (.A(\atari2600.ram[23][7] ),
    .X(net4336));
 sg13g2_dlygate4sd3_1 hold1447 (.A(\scanline[84][2] ),
    .X(net4337));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\atari2600.ram[31][5] ),
    .X(net4338));
 sg13g2_dlygate4sd3_1 hold1449 (.A(\scanline[8][2] ),
    .X(net4339));
 sg13g2_dlygate4sd3_1 hold1450 (.A(\atari2600.ram[101][3] ),
    .X(net4340));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\atari2600.ram[31][6] ),
    .X(net4341));
 sg13g2_dlygate4sd3_1 hold1452 (.A(\atari2600.ram[125][2] ),
    .X(net4342));
 sg13g2_dlygate4sd3_1 hold1453 (.A(\atari2600.ram[63][2] ),
    .X(net4343));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\scanline[12][4] ),
    .X(net4344));
 sg13g2_dlygate4sd3_1 hold1455 (.A(\atari2600.ram[111][3] ),
    .X(net4345));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\atari2600.ram[43][0] ),
    .X(net4346));
 sg13g2_dlygate4sd3_1 hold1457 (.A(\atari2600.ram[57][5] ),
    .X(net4347));
 sg13g2_dlygate4sd3_1 hold1458 (.A(\scanline[108][6] ),
    .X(net4348));
 sg13g2_dlygate4sd3_1 hold1459 (.A(\atari2600.ram[111][2] ),
    .X(net4349));
 sg13g2_dlygate4sd3_1 hold1460 (.A(\scanline[38][5] ),
    .X(net4350));
 sg13g2_dlygate4sd3_1 hold1461 (.A(\atari2600.ram[116][4] ),
    .X(net4351));
 sg13g2_dlygate4sd3_1 hold1462 (.A(\scanline[20][3] ),
    .X(net4352));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\atari2600.ram[124][5] ),
    .X(net4353));
 sg13g2_dlygate4sd3_1 hold1464 (.A(\atari2600.ram[4][3] ),
    .X(net4354));
 sg13g2_dlygate4sd3_1 hold1465 (.A(\scanline[10][4] ),
    .X(net4355));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\atari2600.ram[59][7] ),
    .X(net4356));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\atari2600.tia.poly9_r.x[8] ),
    .X(net4357));
 sg13g2_dlygate4sd3_1 hold1468 (.A(_02258_),
    .X(net4358));
 sg13g2_dlygate4sd3_1 hold1469 (.A(\scanline[120][3] ),
    .X(net4359));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\scanline[70][1] ),
    .X(net4360));
 sg13g2_dlygate4sd3_1 hold1471 (.A(\atari2600.ram[39][0] ),
    .X(net4361));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\atari2600.ram[20][5] ),
    .X(net4362));
 sg13g2_dlygate4sd3_1 hold1473 (.A(\atari2600.ram[21][3] ),
    .X(net4363));
 sg13g2_dlygate4sd3_1 hold1474 (.A(\atari2600.ram[103][3] ),
    .X(net4364));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\atari2600.ram[117][4] ),
    .X(net4365));
 sg13g2_dlygate4sd3_1 hold1476 (.A(\scanline[140][1] ),
    .X(net4366));
 sg13g2_dlygate4sd3_1 hold1477 (.A(\atari2600.ram[40][1] ),
    .X(net4367));
 sg13g2_dlygate4sd3_1 hold1478 (.A(\scanline[140][4] ),
    .X(net4368));
 sg13g2_dlygate4sd3_1 hold1479 (.A(\scanline[50][6] ),
    .X(net4369));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\atari2600.ram[0][0] ),
    .X(net4370));
 sg13g2_dlygate4sd3_1 hold1481 (.A(\atari2600.ram[112][5] ),
    .X(net4371));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\scanline[60][6] ),
    .X(net4372));
 sg13g2_dlygate4sd3_1 hold1483 (.A(\scanline[129][1] ),
    .X(net4373));
 sg13g2_dlygate4sd3_1 hold1484 (.A(\scanline[144][0] ),
    .X(net4374));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\atari2600.ram[55][2] ),
    .X(net4375));
 sg13g2_dlygate4sd3_1 hold1486 (.A(\atari2600.ram[97][5] ),
    .X(net4376));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\scanline[36][6] ),
    .X(net4377));
 sg13g2_dlygate4sd3_1 hold1488 (.A(\atari2600.ram[4][0] ),
    .X(net4378));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\atari2600.ram[51][6] ),
    .X(net4379));
 sg13g2_dlygate4sd3_1 hold1490 (.A(\scanline[100][3] ),
    .X(net4380));
 sg13g2_dlygate4sd3_1 hold1491 (.A(\atari2600.ram[29][1] ),
    .X(net4381));
 sg13g2_dlygate4sd3_1 hold1492 (.A(\scanline[130][6] ),
    .X(net4382));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\atari2600.ram[87][5] ),
    .X(net4383));
 sg13g2_dlygate4sd3_1 hold1494 (.A(\atari2600.ram[84][0] ),
    .X(net4384));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\atari2600.ram[20][7] ),
    .X(net4385));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\atari2600.ram[48][1] ),
    .X(net4386));
 sg13g2_dlygate4sd3_1 hold1497 (.A(\atari2600.cpu.AXYS[1][4] ),
    .X(net4387));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\atari2600.ram[39][2] ),
    .X(net4388));
 sg13g2_dlygate4sd3_1 hold1499 (.A(\scanline[35][6] ),
    .X(net4389));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\atari2600.ram[28][1] ),
    .X(net4390));
 sg13g2_dlygate4sd3_1 hold1501 (.A(\atari2600.ram[47][1] ),
    .X(net4391));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\atari2600.cpu.AXYS[3][2] ),
    .X(net4392));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\atari2600.ram[101][1] ),
    .X(net4393));
 sg13g2_dlygate4sd3_1 hold1504 (.A(\scanline[56][2] ),
    .X(net4394));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\atari2600.ram[15][3] ),
    .X(net4395));
 sg13g2_dlygate4sd3_1 hold1506 (.A(\atari2600.ram[8][0] ),
    .X(net4396));
 sg13g2_dlygate4sd3_1 hold1507 (.A(\scanline[137][4] ),
    .X(net4397));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\atari2600.ram[11][0] ),
    .X(net4398));
 sg13g2_dlygate4sd3_1 hold1509 (.A(\scanline[28][5] ),
    .X(net4399));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\atari2600.tia.ball_w[2] ),
    .X(net4400));
 sg13g2_dlygate4sd3_1 hold1511 (.A(\atari2600.ram[108][5] ),
    .X(net4401));
 sg13g2_dlygate4sd3_1 hold1512 (.A(\atari2600.ram[40][2] ),
    .X(net4402));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\atari2600.ram[80][1] ),
    .X(net4403));
 sg13g2_dlygate4sd3_1 hold1514 (.A(\scanline[98][6] ),
    .X(net4404));
 sg13g2_dlygate4sd3_1 hold1515 (.A(\atari2600.ram[28][4] ),
    .X(net4405));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\scanline[133][5] ),
    .X(net4406));
 sg13g2_dlygate4sd3_1 hold1517 (.A(\scanline[28][6] ),
    .X(net4407));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\atari2600.ram[49][5] ),
    .X(net4408));
 sg13g2_dlygate4sd3_1 hold1519 (.A(\atari2600.ram[64][2] ),
    .X(net4409));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\atari2600.cpu.write_back ),
    .X(net4410));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\atari2600.ram[127][1] ),
    .X(net4411));
 sg13g2_dlygate4sd3_1 hold1522 (.A(\atari2600.ram[59][2] ),
    .X(net4412));
 sg13g2_dlygate4sd3_1 hold1523 (.A(\scanline[37][3] ),
    .X(net4413));
 sg13g2_dlygate4sd3_1 hold1524 (.A(\atari2600.tia.poly9_r.x[3] ),
    .X(net4414));
 sg13g2_dlygate4sd3_1 hold1525 (.A(_02253_),
    .X(net4415));
 sg13g2_dlygate4sd3_1 hold1526 (.A(\scanline[144][1] ),
    .X(net4416));
 sg13g2_dlygate4sd3_1 hold1527 (.A(\scanline[36][5] ),
    .X(net4417));
 sg13g2_dlygate4sd3_1 hold1528 (.A(\atari2600.ram[15][6] ),
    .X(net4418));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\atari2600.ram[41][5] ),
    .X(net4419));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\atari2600.ram[117][2] ),
    .X(net4420));
 sg13g2_dlygate4sd3_1 hold1531 (.A(\atari2600.ram[47][7] ),
    .X(net4421));
 sg13g2_dlygate4sd3_1 hold1532 (.A(\atari2600.ram[101][2] ),
    .X(net4422));
 sg13g2_dlygate4sd3_1 hold1533 (.A(\atari2600.ram[111][5] ),
    .X(net4423));
 sg13g2_dlygate4sd3_1 hold1534 (.A(\atari2600.ram[57][0] ),
    .X(net4424));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\atari2600.cpu.AXYS[2][4] ),
    .X(net4425));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\scanline[40][2] ),
    .X(net4426));
 sg13g2_dlygate4sd3_1 hold1537 (.A(\atari2600.ram[7][2] ),
    .X(net4427));
 sg13g2_dlygate4sd3_1 hold1538 (.A(\scanline[33][1] ),
    .X(net4428));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\atari2600.ram[99][4] ),
    .X(net4429));
 sg13g2_dlygate4sd3_1 hold1540 (.A(\scanline[148][6] ),
    .X(net4430));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\atari2600.ram[60][5] ),
    .X(net4431));
 sg13g2_dlygate4sd3_1 hold1542 (.A(\atari2600.ram[5][6] ),
    .X(net4432));
 sg13g2_dlygate4sd3_1 hold1543 (.A(\scanline[148][2] ),
    .X(net4433));
 sg13g2_dlygate4sd3_1 hold1544 (.A(\scanline[144][3] ),
    .X(net4434));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\scanline[116][0] ),
    .X(net4435));
 sg13g2_dlygate4sd3_1 hold1546 (.A(\atari2600.ram[71][0] ),
    .X(net4436));
 sg13g2_dlygate4sd3_1 hold1547 (.A(\atari2600.ram[81][6] ),
    .X(net4437));
 sg13g2_dlygate4sd3_1 hold1548 (.A(\atari2600.ram[69][4] ),
    .X(net4438));
 sg13g2_dlygate4sd3_1 hold1549 (.A(\scanline[137][1] ),
    .X(net4439));
 sg13g2_dlygate4sd3_1 hold1550 (.A(\atari2600.ram[12][5] ),
    .X(net4440));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\atari2600.ram[27][4] ),
    .X(net4441));
 sg13g2_dlygate4sd3_1 hold1552 (.A(\scanline[65][6] ),
    .X(net4442));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\atari2600.ram[60][2] ),
    .X(net4443));
 sg13g2_dlygate4sd3_1 hold1554 (.A(\atari2600.ram[87][4] ),
    .X(net4444));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\atari2600.ram[19][4] ),
    .X(net4445));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\atari2600.ram[19][3] ),
    .X(net4446));
 sg13g2_dlygate4sd3_1 hold1557 (.A(\scanline[41][0] ),
    .X(net4447));
 sg13g2_dlygate4sd3_1 hold1558 (.A(\atari2600.ram[117][1] ),
    .X(net4448));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\atari2600.ram[7][4] ),
    .X(net4449));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\atari2600.ram[60][7] ),
    .X(net4450));
 sg13g2_dlygate4sd3_1 hold1561 (.A(\atari2600.ram[108][6] ),
    .X(net4451));
 sg13g2_dlygate4sd3_1 hold1562 (.A(\atari2600.ram[68][7] ),
    .X(net4452));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\atari2600.ram[29][7] ),
    .X(net4453));
 sg13g2_dlygate4sd3_1 hold1564 (.A(\atari2600.cpu.AXYS[0][2] ),
    .X(net4454));
 sg13g2_dlygate4sd3_1 hold1565 (.A(\scanline[40][6] ),
    .X(net4455));
 sg13g2_dlygate4sd3_1 hold1566 (.A(\atari2600.ram[105][5] ),
    .X(net4456));
 sg13g2_dlygate4sd3_1 hold1567 (.A(\atari2600.ram[47][4] ),
    .X(net4457));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\scanline[24][3] ),
    .X(net4458));
 sg13g2_dlygate4sd3_1 hold1569 (.A(\atari2600.ram[119][2] ),
    .X(net4459));
 sg13g2_dlygate4sd3_1 hold1570 (.A(\atari2600.ram[27][0] ),
    .X(net4460));
 sg13g2_dlygate4sd3_1 hold1571 (.A(\atari2600.ram[116][7] ),
    .X(net4461));
 sg13g2_dlygate4sd3_1 hold1572 (.A(\atari2600.ram[48][3] ),
    .X(net4462));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\atari2600.ram[44][0] ),
    .X(net4463));
 sg13g2_dlygate4sd3_1 hold1574 (.A(\atari2600.ram[23][1] ),
    .X(net4464));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\atari2600.ram[56][1] ),
    .X(net4465));
 sg13g2_dlygate4sd3_1 hold1576 (.A(\scanline[16][5] ),
    .X(net4466));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\scanline[11][3] ),
    .X(net4467));
 sg13g2_dlygate4sd3_1 hold1578 (.A(\atari2600.ram[19][0] ),
    .X(net4468));
 sg13g2_dlygate4sd3_1 hold1579 (.A(\scanline[21][5] ),
    .X(net4469));
 sg13g2_dlygate4sd3_1 hold1580 (.A(\atari2600.ram[39][6] ),
    .X(net4470));
 sg13g2_dlygate4sd3_1 hold1581 (.A(\scanline[145][3] ),
    .X(net4471));
 sg13g2_dlygate4sd3_1 hold1582 (.A(\atari2600.ram[103][1] ),
    .X(net4472));
 sg13g2_dlygate4sd3_1 hold1583 (.A(\atari2600.ram[99][1] ),
    .X(net4473));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\atari2600.ram[31][2] ),
    .X(net4474));
 sg13g2_dlygate4sd3_1 hold1585 (.A(\atari2600.ram[97][6] ),
    .X(net4475));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\scanline[69][1] ),
    .X(net4476));
 sg13g2_dlygate4sd3_1 hold1587 (.A(\atari2600.ram[101][7] ),
    .X(net4477));
 sg13g2_dlygate4sd3_1 hold1588 (.A(\scanline[96][0] ),
    .X(net4478));
 sg13g2_dlygate4sd3_1 hold1589 (.A(\atari2600.ram[96][3] ),
    .X(net4479));
 sg13g2_dlygate4sd3_1 hold1590 (.A(\atari2600.ram[103][0] ),
    .X(net4480));
 sg13g2_dlygate4sd3_1 hold1591 (.A(\scanline[17][3] ),
    .X(net4481));
 sg13g2_dlygate4sd3_1 hold1592 (.A(\atari2600.ram[61][6] ),
    .X(net4482));
 sg13g2_dlygate4sd3_1 hold1593 (.A(\scanline[43][6] ),
    .X(net4483));
 sg13g2_dlygate4sd3_1 hold1594 (.A(\atari2600.ram[9][7] ),
    .X(net4484));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\scanline[108][4] ),
    .X(net4485));
 sg13g2_dlygate4sd3_1 hold1596 (.A(\scanline[128][0] ),
    .X(net4486));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\scanline[19][3] ),
    .X(net4487));
 sg13g2_dlygate4sd3_1 hold1598 (.A(\atari2600.ram[116][2] ),
    .X(net4488));
 sg13g2_dlygate4sd3_1 hold1599 (.A(\atari2600.ram[44][4] ),
    .X(net4489));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\scanline[70][0] ),
    .X(net4490));
 sg13g2_dlygate4sd3_1 hold1601 (.A(\scanline[35][1] ),
    .X(net4491));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\atari2600.ram[85][7] ),
    .X(net4492));
 sg13g2_dlygate4sd3_1 hold1603 (.A(\scanline[37][5] ),
    .X(net4493));
 sg13g2_dlygate4sd3_1 hold1604 (.A(\atari2600.ram[69][6] ),
    .X(net4494));
 sg13g2_dlygate4sd3_1 hold1605 (.A(\atari2600.ram[61][0] ),
    .X(net4495));
 sg13g2_dlygate4sd3_1 hold1606 (.A(\atari2600.ram[4][1] ),
    .X(net4496));
 sg13g2_dlygate4sd3_1 hold1607 (.A(\atari2600.ram[105][1] ),
    .X(net4497));
 sg13g2_dlygate4sd3_1 hold1608 (.A(\atari2600.ram[52][5] ),
    .X(net4498));
 sg13g2_dlygate4sd3_1 hold1609 (.A(\atari2600.ram[22][6] ),
    .X(net4499));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\atari2600.ram[31][1] ),
    .X(net4500));
 sg13g2_dlygate4sd3_1 hold1611 (.A(\scanline[9][1] ),
    .X(net4501));
 sg13g2_dlygate4sd3_1 hold1612 (.A(\scanline[2][6] ),
    .X(net4502));
 sg13g2_dlygate4sd3_1 hold1613 (.A(\scanline[48][2] ),
    .X(net4503));
 sg13g2_dlygate4sd3_1 hold1614 (.A(\atari2600.ram[127][0] ),
    .X(net4504));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\scanline[82][0] ),
    .X(net4505));
 sg13g2_dlygate4sd3_1 hold1616 (.A(\scanline[25][0] ),
    .X(net4506));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\atari2600.ram[36][1] ),
    .X(net4507));
 sg13g2_dlygate4sd3_1 hold1618 (.A(\atari2600.ram[59][3] ),
    .X(net4508));
 sg13g2_dlygate4sd3_1 hold1619 (.A(\atari2600.ram[99][6] ),
    .X(net4509));
 sg13g2_dlygate4sd3_1 hold1620 (.A(\scanline[25][2] ),
    .X(net4510));
 sg13g2_dlygate4sd3_1 hold1621 (.A(\scanline[96][2] ),
    .X(net4511));
 sg13g2_dlygate4sd3_1 hold1622 (.A(\scanline[145][1] ),
    .X(net4512));
 sg13g2_dlygate4sd3_1 hold1623 (.A(\atari2600.ram[100][5] ),
    .X(net4513));
 sg13g2_dlygate4sd3_1 hold1624 (.A(\atari2600.ram[120][3] ),
    .X(net4514));
 sg13g2_dlygate4sd3_1 hold1625 (.A(\scanline[64][1] ),
    .X(net4515));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\scanline[24][1] ),
    .X(net4516));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\atari2600.ram[51][5] ),
    .X(net4517));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\atari2600.ram[17][0] ),
    .X(net4518));
 sg13g2_dlygate4sd3_1 hold1629 (.A(\scanline[152][2] ),
    .X(net4519));
 sg13g2_dlygate4sd3_1 hold1630 (.A(\scanline[8][5] ),
    .X(net4520));
 sg13g2_dlygate4sd3_1 hold1631 (.A(\atari2600.ram[116][3] ),
    .X(net4521));
 sg13g2_dlygate4sd3_1 hold1632 (.A(\atari2600.ram[71][6] ),
    .X(net4522));
 sg13g2_dlygate4sd3_1 hold1633 (.A(\atari2600.ram[85][5] ),
    .X(net4523));
 sg13g2_dlygate4sd3_1 hold1634 (.A(\atari2600.ram[28][7] ),
    .X(net4524));
 sg13g2_dlygate4sd3_1 hold1635 (.A(\atari2600.ram[31][4] ),
    .X(net4525));
 sg13g2_dlygate4sd3_1 hold1636 (.A(\atari2600.ram[17][3] ),
    .X(net4526));
 sg13g2_dlygate4sd3_1 hold1637 (.A(\scanline[74][1] ),
    .X(net4527));
 sg13g2_dlygate4sd3_1 hold1638 (.A(\scanline[131][5] ),
    .X(net4528));
 sg13g2_dlygate4sd3_1 hold1639 (.A(\atari2600.ram[121][0] ),
    .X(net4529));
 sg13g2_dlygate4sd3_1 hold1640 (.A(\scanline[39][5] ),
    .X(net4530));
 sg13g2_dlygate4sd3_1 hold1641 (.A(\atari2600.ram[104][7] ),
    .X(net4531));
 sg13g2_dlygate4sd3_1 hold1642 (.A(\atari2600.pia.dat_o[5] ),
    .X(net4532));
 sg13g2_dlygate4sd3_1 hold1643 (.A(_07159_),
    .X(net4533));
 sg13g2_dlygate4sd3_1 hold1644 (.A(\atari2600.ram[113][5] ),
    .X(net4534));
 sg13g2_dlygate4sd3_1 hold1645 (.A(\scanline[10][3] ),
    .X(net4535));
 sg13g2_dlygate4sd3_1 hold1646 (.A(\atari2600.ram[63][6] ),
    .X(net4536));
 sg13g2_dlygate4sd3_1 hold1647 (.A(\atari2600.ram[4][6] ),
    .X(net4537));
 sg13g2_dlygate4sd3_1 hold1648 (.A(\scanline[69][5] ),
    .X(net4538));
 sg13g2_dlygate4sd3_1 hold1649 (.A(\atari2600.ram[85][1] ),
    .X(net4539));
 sg13g2_dlygate4sd3_1 hold1650 (.A(\atari2600.ram[67][5] ),
    .X(net4540));
 sg13g2_dlygate4sd3_1 hold1651 (.A(\atari2600.ram[81][0] ),
    .X(net4541));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\atari2600.ram[120][5] ),
    .X(net4542));
 sg13g2_dlygate4sd3_1 hold1653 (.A(\atari2600.ram[32][6] ),
    .X(net6040));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\scanline[133][3] ),
    .X(net6041));
 sg13g2_dlygate4sd3_1 hold1655 (.A(\scanline[133][0] ),
    .X(net6042));
 sg13g2_dlygate4sd3_1 hold1656 (.A(\scanline[20][1] ),
    .X(net6043));
 sg13g2_dlygate4sd3_1 hold1657 (.A(\atari2600.ram[12][0] ),
    .X(net6044));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\atari2600.cpu.AXYS[2][2] ),
    .X(net6045));
 sg13g2_dlygate4sd3_1 hold1659 (.A(\atari2600.ram[87][3] ),
    .X(net6046));
 sg13g2_dlygate4sd3_1 hold1660 (.A(\scanline[133][4] ),
    .X(net6047));
 sg13g2_dlygate4sd3_1 hold1661 (.A(\atari2600.ram[33][2] ),
    .X(net6048));
 sg13g2_dlygate4sd3_1 hold1662 (.A(\atari2600.ram[85][4] ),
    .X(net6049));
 sg13g2_dlygate4sd3_1 hold1663 (.A(\atari2600.ram[41][7] ),
    .X(net6050));
 sg13g2_dlygate4sd3_1 hold1664 (.A(\atari2600.ram[112][7] ),
    .X(net6051));
 sg13g2_dlygate4sd3_1 hold1665 (.A(\scanline[5][5] ),
    .X(net6052));
 sg13g2_dlygate4sd3_1 hold1666 (.A(\scanline[92][1] ),
    .X(net6053));
 sg13g2_dlygate4sd3_1 hold1667 (.A(\atari2600.ram[53][7] ),
    .X(net6054));
 sg13g2_dlygate4sd3_1 hold1668 (.A(\atari2600.ram[23][0] ),
    .X(net6055));
 sg13g2_dlygate4sd3_1 hold1669 (.A(\scanline[65][5] ),
    .X(net6056));
 sg13g2_dlygate4sd3_1 hold1670 (.A(\atari2600.ram[109][6] ),
    .X(net6057));
 sg13g2_dlygate4sd3_1 hold1671 (.A(\scanline[39][1] ),
    .X(net6058));
 sg13g2_dlygate4sd3_1 hold1672 (.A(\atari2600.ram[107][6] ),
    .X(net6059));
 sg13g2_dlygate4sd3_1 hold1673 (.A(\atari2600.ram[83][4] ),
    .X(net6060));
 sg13g2_dlygate4sd3_1 hold1674 (.A(\atari2600.ram[111][0] ),
    .X(net6061));
 sg13g2_dlygate4sd3_1 hold1675 (.A(\atari2600.ram[36][7] ),
    .X(net6062));
 sg13g2_dlygate4sd3_1 hold1676 (.A(\atari2600.ram[68][1] ),
    .X(net6063));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\scanline[69][6] ),
    .X(net6064));
 sg13g2_dlygate4sd3_1 hold1678 (.A(\atari2600.ram[8][2] ),
    .X(net6065));
 sg13g2_dlygate4sd3_1 hold1679 (.A(\atari2600.ram_data[2] ),
    .X(net6066));
 sg13g2_dlygate4sd3_1 hold1680 (.A(_07152_),
    .X(net6067));
 sg13g2_dlygate4sd3_1 hold1681 (.A(\scanline[12][6] ),
    .X(net6068));
 sg13g2_dlygate4sd3_1 hold1682 (.A(\atari2600.ram[63][0] ),
    .X(net6069));
 sg13g2_dlygate4sd3_1 hold1683 (.A(\scanline[38][4] ),
    .X(net6070));
 sg13g2_dlygate4sd3_1 hold1684 (.A(\scanline[120][6] ),
    .X(net6071));
 sg13g2_dlygate4sd3_1 hold1685 (.A(\atari2600.ram[81][4] ),
    .X(net6072));
 sg13g2_dlygate4sd3_1 hold1686 (.A(\atari2600.ram[109][4] ),
    .X(net6073));
 sg13g2_dlygate4sd3_1 hold1687 (.A(\scanline[96][1] ),
    .X(net6074));
 sg13g2_dlygate4sd3_1 hold1688 (.A(\atari2600.ram[16][6] ),
    .X(net6075));
 sg13g2_dlygate4sd3_1 hold1689 (.A(\atari2600.ram[56][3] ),
    .X(net6076));
 sg13g2_dlygate4sd3_1 hold1690 (.A(\scanline[16][6] ),
    .X(net6077));
 sg13g2_dlygate4sd3_1 hold1691 (.A(\atari2600.ram[48][5] ),
    .X(net6078));
 sg13g2_dlygate4sd3_1 hold1692 (.A(\scanline[139][4] ),
    .X(net6079));
 sg13g2_dlygate4sd3_1 hold1693 (.A(\scanline[134][0] ),
    .X(net6080));
 sg13g2_dlygate4sd3_1 hold1694 (.A(\scanline[24][0] ),
    .X(net6081));
 sg13g2_dlygate4sd3_1 hold1695 (.A(\atari2600.ram[29][6] ),
    .X(net6082));
 sg13g2_dlygate4sd3_1 hold1696 (.A(\atari2600.ram[16][2] ),
    .X(net6083));
 sg13g2_dlygate4sd3_1 hold1697 (.A(\scanline[17][5] ),
    .X(net6084));
 sg13g2_dlygate4sd3_1 hold1698 (.A(\atari2600.ram[84][1] ),
    .X(net6085));
 sg13g2_dlygate4sd3_1 hold1699 (.A(\atari2600.ram[65][3] ),
    .X(net6086));
 sg13g2_dlygate4sd3_1 hold1700 (.A(\scanline[131][0] ),
    .X(net6087));
 sg13g2_dlygate4sd3_1 hold1701 (.A(\scanline[75][5] ),
    .X(net6088));
 sg13g2_dlygate4sd3_1 hold1702 (.A(\atari2600.ram[100][2] ),
    .X(net6089));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\atari2600.ram[37][1] ),
    .X(net6090));
 sg13g2_dlygate4sd3_1 hold1704 (.A(\atari2600.cpu.ALU.AI7 ),
    .X(net6091));
 sg13g2_dlygate4sd3_1 hold1705 (.A(_02487_),
    .X(net6092));
 sg13g2_dlygate4sd3_1 hold1706 (.A(\scanline[26][3] ),
    .X(net6093));
 sg13g2_dlygate4sd3_1 hold1707 (.A(\atari2600.ram[97][2] ),
    .X(net6094));
 sg13g2_dlygate4sd3_1 hold1708 (.A(\atari2600.ram[68][0] ),
    .X(net6095));
 sg13g2_dlygate4sd3_1 hold1709 (.A(\scanline[42][4] ),
    .X(net6096));
 sg13g2_dlygate4sd3_1 hold1710 (.A(\scanline[44][5] ),
    .X(net6097));
 sg13g2_dlygate4sd3_1 hold1711 (.A(\atari2600.ram[19][1] ),
    .X(net6098));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\scanline[132][1] ),
    .X(net6099));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\scanline[35][3] ),
    .X(net6100));
 sg13g2_dlygate4sd3_1 hold1714 (.A(\scanline[60][5] ),
    .X(net6101));
 sg13g2_dlygate4sd3_1 hold1715 (.A(\atari2600.ram[121][1] ),
    .X(net6102));
 sg13g2_dlygate4sd3_1 hold1716 (.A(\atari2600.ram[25][7] ),
    .X(net6103));
 sg13g2_dlygate4sd3_1 hold1717 (.A(\atari2600.ram[117][6] ),
    .X(net6104));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\atari2600.ram[17][6] ),
    .X(net6105));
 sg13g2_dlygate4sd3_1 hold1719 (.A(\atari2600.ram[27][7] ),
    .X(net6106));
 sg13g2_dlygate4sd3_1 hold1720 (.A(\scanline[0][0] ),
    .X(net6107));
 sg13g2_dlygate4sd3_1 hold1721 (.A(\atari2600.ram[15][7] ),
    .X(net6108));
 sg13g2_dlygate4sd3_1 hold1722 (.A(\atari2600.ram[60][6] ),
    .X(net6109));
 sg13g2_dlygate4sd3_1 hold1723 (.A(\atari2600.ram[127][7] ),
    .X(net6110));
 sg13g2_dlygate4sd3_1 hold1724 (.A(\scanline[5][3] ),
    .X(net6111));
 sg13g2_dlygate4sd3_1 hold1725 (.A(\scanline[43][2] ),
    .X(net6112));
 sg13g2_dlygate4sd3_1 hold1726 (.A(\scanline[68][0] ),
    .X(net6113));
 sg13g2_dlygate4sd3_1 hold1727 (.A(\atari2600.ram[101][4] ),
    .X(net6114));
 sg13g2_dlygate4sd3_1 hold1728 (.A(\scanline[38][3] ),
    .X(net6115));
 sg13g2_dlygate4sd3_1 hold1729 (.A(\scanline[135][2] ),
    .X(net6116));
 sg13g2_dlygate4sd3_1 hold1730 (.A(\atari2600.ram[119][6] ),
    .X(net6117));
 sg13g2_dlygate4sd3_1 hold1731 (.A(\atari2600.ram[29][0] ),
    .X(net6118));
 sg13g2_dlygate4sd3_1 hold1732 (.A(\atari2600.ram[5][5] ),
    .X(net6119));
 sg13g2_dlygate4sd3_1 hold1733 (.A(\atari2600.ram[67][0] ),
    .X(net6120));
 sg13g2_dlygate4sd3_1 hold1734 (.A(\atari2600.ram[123][3] ),
    .X(net6121));
 sg13g2_dlygate4sd3_1 hold1735 (.A(\atari2600.cpu.AXYS[2][5] ),
    .X(net6122));
 sg13g2_dlygate4sd3_1 hold1736 (.A(\scanline[71][2] ),
    .X(net6123));
 sg13g2_dlygate4sd3_1 hold1737 (.A(\atari2600.ram[113][3] ),
    .X(net6124));
 sg13g2_dlygate4sd3_1 hold1738 (.A(\atari2600.ram[83][1] ),
    .X(net6125));
 sg13g2_dlygate4sd3_1 hold1739 (.A(\atari2600.ram[124][6] ),
    .X(net6126));
 sg13g2_dlygate4sd3_1 hold1740 (.A(\atari2600.ram[103][6] ),
    .X(net6127));
 sg13g2_dlygate4sd3_1 hold1741 (.A(\atari2600.ram[63][7] ),
    .X(net6128));
 sg13g2_dlygate4sd3_1 hold1742 (.A(\atari2600.ram[87][7] ),
    .X(net6129));
 sg13g2_dlygate4sd3_1 hold1743 (.A(\atari2600.ram[4][7] ),
    .X(net6130));
 sg13g2_dlygate4sd3_1 hold1744 (.A(\scanline[23][0] ),
    .X(net6131));
 sg13g2_dlygate4sd3_1 hold1745 (.A(\atari2600.ram[35][5] ),
    .X(net6132));
 sg13g2_dlygate4sd3_1 hold1746 (.A(\scanline[40][1] ),
    .X(net6133));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\scanline[132][0] ),
    .X(net6134));
 sg13g2_dlygate4sd3_1 hold1748 (.A(\atari2600.ram[104][3] ),
    .X(net6135));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\scanline[152][4] ),
    .X(net6136));
 sg13g2_dlygate4sd3_1 hold1750 (.A(\scanline[82][3] ),
    .X(net6137));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\atari2600.tia.refp0 ),
    .X(net6138));
 sg13g2_dlygate4sd3_1 hold1752 (.A(\atari2600.ram[45][1] ),
    .X(net6139));
 sg13g2_dlygate4sd3_1 hold1753 (.A(\scanline[32][3] ),
    .X(net6140));
 sg13g2_dlygate4sd3_1 hold1754 (.A(\atari2600.ram[83][0] ),
    .X(net6141));
 sg13g2_dlygate4sd3_1 hold1755 (.A(\atari2600.ram[111][6] ),
    .X(net6142));
 sg13g2_dlygate4sd3_1 hold1756 (.A(\scanline[36][4] ),
    .X(net6143));
 sg13g2_dlygate4sd3_1 hold1757 (.A(\atari2600.ram[13][2] ),
    .X(net6144));
 sg13g2_dlygate4sd3_1 hold1758 (.A(\atari2600.ram[96][2] ),
    .X(net6145));
 sg13g2_dlygate4sd3_1 hold1759 (.A(\atari2600.ram[99][3] ),
    .X(net6146));
 sg13g2_dlygate4sd3_1 hold1760 (.A(\scanline[81][2] ),
    .X(net6147));
 sg13g2_dlygate4sd3_1 hold1761 (.A(\atari2600.ram[64][5] ),
    .X(net6148));
 sg13g2_dlygate4sd3_1 hold1762 (.A(\scanline[44][0] ),
    .X(net6149));
 sg13g2_dlygate4sd3_1 hold1763 (.A(\atari2600.pia.time_counter[8] ),
    .X(net6150));
 sg13g2_dlygate4sd3_1 hold1764 (.A(_01780_),
    .X(net6151));
 sg13g2_dlygate4sd3_1 hold1765 (.A(\scanline[20][2] ),
    .X(net6152));
 sg13g2_dlygate4sd3_1 hold1766 (.A(\atari2600.ram[81][2] ),
    .X(net6153));
 sg13g2_dlygate4sd3_1 hold1767 (.A(\atari2600.ram[66][2] ),
    .X(net6154));
 sg13g2_dlygate4sd3_1 hold1768 (.A(\scanline[128][4] ),
    .X(net6155));
 sg13g2_dlygate4sd3_1 hold1769 (.A(\scanline[39][3] ),
    .X(net6156));
 sg13g2_dlygate4sd3_1 hold1770 (.A(\scanline[60][1] ),
    .X(net6157));
 sg13g2_dlygate4sd3_1 hold1771 (.A(\atari2600.ram[127][5] ),
    .X(net6158));
 sg13g2_dlygate4sd3_1 hold1772 (.A(\scanline[12][5] ),
    .X(net6159));
 sg13g2_dlygate4sd3_1 hold1773 (.A(\atari2600.ram[67][2] ),
    .X(net6160));
 sg13g2_dlygate4sd3_1 hold1774 (.A(\scanline[12][1] ),
    .X(net6161));
 sg13g2_dlygate4sd3_1 hold1775 (.A(\scanline[66][2] ),
    .X(net6162));
 sg13g2_dlygate4sd3_1 hold1776 (.A(\scanline[144][5] ),
    .X(net6163));
 sg13g2_dlygate4sd3_1 hold1777 (.A(\atari2600.tia.colup0[2] ),
    .X(net6164));
 sg13g2_dlygate4sd3_1 hold1778 (.A(\scanline[152][6] ),
    .X(net6165));
 sg13g2_dlygate4sd3_1 hold1779 (.A(\atari2600.ram[19][5] ),
    .X(net6166));
 sg13g2_dlygate4sd3_1 hold1780 (.A(\atari2600.ram[80][4] ),
    .X(net6167));
 sg13g2_dlygate4sd3_1 hold1781 (.A(\scanline[116][3] ),
    .X(net6168));
 sg13g2_dlygate4sd3_1 hold1782 (.A(\atari2600.ram[13][0] ),
    .X(net6169));
 sg13g2_dlygate4sd3_1 hold1783 (.A(\atari2600.tia.diag[85] ),
    .X(net6170));
 sg13g2_dlygate4sd3_1 hold1784 (.A(\atari2600.ram[51][2] ),
    .X(net6171));
 sg13g2_dlygate4sd3_1 hold1785 (.A(\atari2600.ram[43][3] ),
    .X(net6172));
 sg13g2_dlygate4sd3_1 hold1786 (.A(\atari2600.cpu.ABH[5] ),
    .X(net6173));
 sg13g2_dlygate4sd3_1 hold1787 (.A(_02982_),
    .X(net6174));
 sg13g2_dlygate4sd3_1 hold1788 (.A(\atari2600.ram[99][2] ),
    .X(net6175));
 sg13g2_dlygate4sd3_1 hold1789 (.A(\atari2600.ram[117][7] ),
    .X(net6176));
 sg13g2_dlygate4sd3_1 hold1790 (.A(\scanline[92][3] ),
    .X(net6177));
 sg13g2_dlygate4sd3_1 hold1791 (.A(\atari2600.ram[53][6] ),
    .X(net6178));
 sg13g2_dlygate4sd3_1 hold1792 (.A(\atari2600.ram[66][0] ),
    .X(net6179));
 sg13g2_dlygate4sd3_1 hold1793 (.A(\atari2600.ram[116][6] ),
    .X(net6180));
 sg13g2_dlygate4sd3_1 hold1794 (.A(\atari2600.ram[124][7] ),
    .X(net6181));
 sg13g2_dlygate4sd3_1 hold1795 (.A(\scanline[81][0] ),
    .X(net6182));
 sg13g2_dlygate4sd3_1 hold1796 (.A(\scanline[26][1] ),
    .X(net6183));
 sg13g2_dlygate4sd3_1 hold1797 (.A(\scanline[71][4] ),
    .X(net6184));
 sg13g2_dlygate4sd3_1 hold1798 (.A(\atari2600.ram[33][6] ),
    .X(net6185));
 sg13g2_dlygate4sd3_1 hold1799 (.A(\scanline[12][0] ),
    .X(net6186));
 sg13g2_dlygate4sd3_1 hold1800 (.A(\scanline[16][0] ),
    .X(net6187));
 sg13g2_dlygate4sd3_1 hold1801 (.A(\scanline[136][3] ),
    .X(net6188));
 sg13g2_dlygate4sd3_1 hold1802 (.A(\atari2600.ram[40][7] ),
    .X(net6189));
 sg13g2_dlygate4sd3_1 hold1803 (.A(\scanline[72][6] ),
    .X(net6190));
 sg13g2_dlygate4sd3_1 hold1804 (.A(\scanline[135][6] ),
    .X(net6191));
 sg13g2_dlygate4sd3_1 hold1805 (.A(\scanline[69][2] ),
    .X(net6192));
 sg13g2_dlygate4sd3_1 hold1806 (.A(\scanline[80][1] ),
    .X(net6193));
 sg13g2_dlygate4sd3_1 hold1807 (.A(\scanline[22][6] ),
    .X(net6194));
 sg13g2_dlygate4sd3_1 hold1808 (.A(\scanline[120][1] ),
    .X(net6195));
 sg13g2_dlygate4sd3_1 hold1809 (.A(\atari2600.ram[37][3] ),
    .X(net6196));
 sg13g2_dlygate4sd3_1 hold1810 (.A(\scanline[138][6] ),
    .X(net6197));
 sg13g2_dlygate4sd3_1 hold1811 (.A(\atari2600.ram[112][0] ),
    .X(net6198));
 sg13g2_dlygate4sd3_1 hold1812 (.A(\scanline[73][2] ),
    .X(net6199));
 sg13g2_dlygate4sd3_1 hold1813 (.A(\scanline[8][6] ),
    .X(net6200));
 sg13g2_dlygate4sd3_1 hold1814 (.A(\scanline[120][2] ),
    .X(net6201));
 sg13g2_dlygate4sd3_1 hold1815 (.A(\scanline[129][5] ),
    .X(net6202));
 sg13g2_dlygate4sd3_1 hold1816 (.A(\atari2600.tia.audio_right_counter[10] ),
    .X(net6203));
 sg13g2_dlygate4sd3_1 hold1817 (.A(_02038_),
    .X(net6204));
 sg13g2_dlygate4sd3_1 hold1818 (.A(\atari2600.ram[65][1] ),
    .X(net6205));
 sg13g2_dlygate4sd3_1 hold1819 (.A(\atari2600.ram[32][1] ),
    .X(net6206));
 sg13g2_dlygate4sd3_1 hold1820 (.A(\atari2600.ram[55][0] ),
    .X(net6207));
 sg13g2_dlygate4sd3_1 hold1821 (.A(\scanline[88][3] ),
    .X(net6208));
 sg13g2_dlygate4sd3_1 hold1822 (.A(\atari2600.pia.reset_timer[3] ),
    .X(net6209));
 sg13g2_dlygate4sd3_1 hold1823 (.A(\atari2600.ram[109][0] ),
    .X(net6210));
 sg13g2_dlygate4sd3_1 hold1824 (.A(\scanline[28][3] ),
    .X(net6211));
 sg13g2_dlygate4sd3_1 hold1825 (.A(\scanline[18][4] ),
    .X(net6212));
 sg13g2_dlygate4sd3_1 hold1826 (.A(\atari2600.ram[57][7] ),
    .X(net6213));
 sg13g2_dlygate4sd3_1 hold1827 (.A(\atari2600.ram[23][2] ),
    .X(net6214));
 sg13g2_dlygate4sd3_1 hold1828 (.A(\scanline[104][6] ),
    .X(net6215));
 sg13g2_dlygate4sd3_1 hold1829 (.A(\scanline[22][3] ),
    .X(net6216));
 sg13g2_dlygate4sd3_1 hold1830 (.A(\atari2600.ram[87][1] ),
    .X(net6217));
 sg13g2_dlygate4sd3_1 hold1831 (.A(\atari2600.ram[115][2] ),
    .X(net6218));
 sg13g2_dlygate4sd3_1 hold1832 (.A(\scanline[34][3] ),
    .X(net6219));
 sg13g2_dlygate4sd3_1 hold1833 (.A(\atari2600.ram[105][2] ),
    .X(net6220));
 sg13g2_dlygate4sd3_1 hold1834 (.A(\atari2600.ram[115][7] ),
    .X(net6221));
 sg13g2_dlygate4sd3_1 hold1835 (.A(\atari2600.ram[64][3] ),
    .X(net6222));
 sg13g2_dlygate4sd3_1 hold1836 (.A(\atari2600.pia.dat_o[3] ),
    .X(net6223));
 sg13g2_dlygate4sd3_1 hold1837 (.A(_01767_),
    .X(net6224));
 sg13g2_dlygate4sd3_1 hold1838 (.A(\scanline[67][3] ),
    .X(net6225));
 sg13g2_dlygate4sd3_1 hold1839 (.A(\scanline[137][2] ),
    .X(net6226));
 sg13g2_dlygate4sd3_1 hold1840 (.A(\atari2600.ram[15][0] ),
    .X(net6227));
 sg13g2_dlygate4sd3_1 hold1841 (.A(\atari2600.ram[33][7] ),
    .X(net6228));
 sg13g2_dlygate4sd3_1 hold1842 (.A(\atari2600.ram[40][0] ),
    .X(net6229));
 sg13g2_dlygate4sd3_1 hold1843 (.A(\scanline[156][1] ),
    .X(net6230));
 sg13g2_dlygate4sd3_1 hold1844 (.A(\scanline[18][1] ),
    .X(net6231));
 sg13g2_dlygate4sd3_1 hold1845 (.A(\scanline[96][3] ),
    .X(net6232));
 sg13g2_dlygate4sd3_1 hold1846 (.A(\scanline[140][0] ),
    .X(net6233));
 sg13g2_dlygate4sd3_1 hold1847 (.A(\scanline[92][5] ),
    .X(net6234));
 sg13g2_dlygate4sd3_1 hold1848 (.A(\atari2600.ram[63][5] ),
    .X(net6235));
 sg13g2_dlygate4sd3_1 hold1849 (.A(\scanline[134][6] ),
    .X(net6236));
 sg13g2_dlygate4sd3_1 hold1850 (.A(\atari2600.ram[31][7] ),
    .X(net6237));
 sg13g2_dlygate4sd3_1 hold1851 (.A(\scanline[130][2] ),
    .X(net6238));
 sg13g2_dlygate4sd3_1 hold1852 (.A(\atari2600.ram[27][3] ),
    .X(net6239));
 sg13g2_dlygate4sd3_1 hold1853 (.A(\atari2600.cpu.AXYS[3][7] ),
    .X(net6240));
 sg13g2_dlygate4sd3_1 hold1854 (.A(\scanline[52][6] ),
    .X(net6241));
 sg13g2_dlygate4sd3_1 hold1855 (.A(\scanline[0][5] ),
    .X(net6242));
 sg13g2_dlygate4sd3_1 hold1856 (.A(\scanline[3][5] ),
    .X(net6243));
 sg13g2_dlygate4sd3_1 hold1857 (.A(\atari2600.ram[53][0] ),
    .X(net6244));
 sg13g2_dlygate4sd3_1 hold1858 (.A(\scanline[24][5] ),
    .X(net6245));
 sg13g2_dlygate4sd3_1 hold1859 (.A(\scanline[21][3] ),
    .X(net6246));
 sg13g2_dlygate4sd3_1 hold1860 (.A(\scanline[104][3] ),
    .X(net6247));
 sg13g2_dlygate4sd3_1 hold1861 (.A(\scanline[16][1] ),
    .X(net6248));
 sg13g2_dlygate4sd3_1 hold1862 (.A(\scanline[82][5] ),
    .X(net6249));
 sg13g2_dlygate4sd3_1 hold1863 (.A(\scanline[80][0] ),
    .X(net6250));
 sg13g2_dlygate4sd3_1 hold1864 (.A(\atari2600.ram[11][6] ),
    .X(net6251));
 sg13g2_dlygate4sd3_1 hold1865 (.A(\scanline[80][5] ),
    .X(net6252));
 sg13g2_dlygate4sd3_1 hold1866 (.A(\atari2600.ram[8][7] ),
    .X(net6253));
 sg13g2_dlygate4sd3_1 hold1867 (.A(\scanline[49][0] ),
    .X(net6254));
 sg13g2_dlygate4sd3_1 hold1868 (.A(\scanline[84][5] ),
    .X(net6255));
 sg13g2_dlygate4sd3_1 hold1869 (.A(\scanline[66][3] ),
    .X(net6256));
 sg13g2_dlygate4sd3_1 hold1870 (.A(\atari2600.ram[28][5] ),
    .X(net6257));
 sg13g2_dlygate4sd3_1 hold1871 (.A(\scanline[70][2] ),
    .X(net6258));
 sg13g2_dlygate4sd3_1 hold1872 (.A(\scanline[38][1] ),
    .X(net6259));
 sg13g2_dlygate4sd3_1 hold1873 (.A(\atari2600.ram[119][7] ),
    .X(net6260));
 sg13g2_dlygate4sd3_1 hold1874 (.A(\scanline[88][4] ),
    .X(net6261));
 sg13g2_dlygate4sd3_1 hold1875 (.A(\scanline[100][6] ),
    .X(net6262));
 sg13g2_dlygate4sd3_1 hold1876 (.A(\scanline[10][6] ),
    .X(net6263));
 sg13g2_dlygate4sd3_1 hold1877 (.A(\scanline[32][0] ),
    .X(net6264));
 sg13g2_dlygate4sd3_1 hold1878 (.A(\scanline[37][1] ),
    .X(net6265));
 sg13g2_dlygate4sd3_1 hold1879 (.A(\atari2600.ram[67][6] ),
    .X(net6266));
 sg13g2_dlygate4sd3_1 hold1880 (.A(\scanline[148][4] ),
    .X(net6267));
 sg13g2_dlygate4sd3_1 hold1881 (.A(\scanline[9][5] ),
    .X(net6268));
 sg13g2_dlygate4sd3_1 hold1882 (.A(\atari2600.ram[0][4] ),
    .X(net6269));
 sg13g2_dlygate4sd3_1 hold1883 (.A(\scanline[9][3] ),
    .X(net6270));
 sg13g2_dlygate4sd3_1 hold1884 (.A(\scanline[88][6] ),
    .X(net6271));
 sg13g2_dlygate4sd3_1 hold1885 (.A(\scanline[74][6] ),
    .X(net6272));
 sg13g2_dlygate4sd3_1 hold1886 (.A(\atari2600.ram[35][3] ),
    .X(net6273));
 sg13g2_dlygate4sd3_1 hold1887 (.A(\scanline[67][6] ),
    .X(net6274));
 sg13g2_dlygate4sd3_1 hold1888 (.A(\atari2600.ram[96][6] ),
    .X(net6275));
 sg13g2_dlygate4sd3_1 hold1889 (.A(\atari2600.ram[111][7] ),
    .X(net6276));
 sg13g2_dlygate4sd3_1 hold1890 (.A(\scanline[20][5] ),
    .X(net6277));
 sg13g2_dlygate4sd3_1 hold1891 (.A(\scanline[97][6] ),
    .X(net6278));
 sg13g2_dlygate4sd3_1 hold1892 (.A(\atari2600.ram[123][0] ),
    .X(net6279));
 sg13g2_dlygate4sd3_1 hold1893 (.A(\scanline[5][0] ),
    .X(net6280));
 sg13g2_dlygate4sd3_1 hold1894 (.A(\atari2600.ram[96][5] ),
    .X(net6281));
 sg13g2_dlygate4sd3_1 hold1895 (.A(\scanline[80][3] ),
    .X(net6282));
 sg13g2_dlygate4sd3_1 hold1896 (.A(\atari2600.ram[59][0] ),
    .X(net6283));
 sg13g2_dlygate4sd3_1 hold1897 (.A(\atari2600.tia.audio_right_counter[4] ),
    .X(net6284));
 sg13g2_dlygate4sd3_1 hold1898 (.A(_02032_),
    .X(net6285));
 sg13g2_dlygate4sd3_1 hold1899 (.A(\scanline[131][1] ),
    .X(net6286));
 sg13g2_dlygate4sd3_1 hold1900 (.A(\scanline[156][5] ),
    .X(net6287));
 sg13g2_dlygate4sd3_1 hold1901 (.A(\scanline[34][2] ),
    .X(net6288));
 sg13g2_dlygate4sd3_1 hold1902 (.A(\atari2600.ram[71][2] ),
    .X(net6289));
 sg13g2_dlygate4sd3_1 hold1903 (.A(\scanline[88][1] ),
    .X(net6290));
 sg13g2_dlygate4sd3_1 hold1904 (.A(\scanline[12][3] ),
    .X(net6291));
 sg13g2_dlygate4sd3_1 hold1905 (.A(\scanline[20][0] ),
    .X(net6292));
 sg13g2_dlygate4sd3_1 hold1906 (.A(\scanline[148][0] ),
    .X(net6293));
 sg13g2_dlygate4sd3_1 hold1907 (.A(\scanline[146][3] ),
    .X(net6294));
 sg13g2_dlygate4sd3_1 hold1908 (.A(\scanline[52][2] ),
    .X(net6295));
 sg13g2_dlygate4sd3_1 hold1909 (.A(\atari2600.ram[11][3] ),
    .X(net6296));
 sg13g2_dlygate4sd3_1 hold1910 (.A(\atari2600.ram[36][6] ),
    .X(net6297));
 sg13g2_dlygate4sd3_1 hold1911 (.A(\frame_counter[1] ),
    .X(net6298));
 sg13g2_dlygate4sd3_1 hold1912 (.A(_01203_),
    .X(net6299));
 sg13g2_dlygate4sd3_1 hold1913 (.A(\scanline[25][6] ),
    .X(net6300));
 sg13g2_dlygate4sd3_1 hold1914 (.A(\scanline[74][0] ),
    .X(net6301));
 sg13g2_dlygate4sd3_1 hold1915 (.A(\atari2600.ram[43][6] ),
    .X(net6302));
 sg13g2_dlygate4sd3_1 hold1916 (.A(\scanline[8][4] ),
    .X(net6303));
 sg13g2_dlygate4sd3_1 hold1917 (.A(\scanline[5][4] ),
    .X(net6304));
 sg13g2_dlygate4sd3_1 hold1918 (.A(\scanline[24][2] ),
    .X(net6305));
 sg13g2_dlygate4sd3_1 hold1919 (.A(\scanline[6][2] ),
    .X(net6306));
 sg13g2_dlygate4sd3_1 hold1920 (.A(\scanline[135][1] ),
    .X(net6307));
 sg13g2_dlygate4sd3_1 hold1921 (.A(\atari2600.ram[23][4] ),
    .X(net6308));
 sg13g2_dlygate4sd3_1 hold1922 (.A(\atari2600.ram[57][2] ),
    .X(net6309));
 sg13g2_dlygate4sd3_1 hold1923 (.A(\atari2600.ram[49][6] ),
    .X(net6310));
 sg13g2_dlygate4sd3_1 hold1924 (.A(\scanline[56][1] ),
    .X(net6311));
 sg13g2_dlygate4sd3_1 hold1925 (.A(\scanline[152][1] ),
    .X(net6312));
 sg13g2_dlygate4sd3_1 hold1926 (.A(\scanline[129][6] ),
    .X(net6313));
 sg13g2_dlygate4sd3_1 hold1927 (.A(\atari2600.ram[71][4] ),
    .X(net6314));
 sg13g2_dlygate4sd3_1 hold1928 (.A(\scanline[84][6] ),
    .X(net6315));
 sg13g2_dlygate4sd3_1 hold1929 (.A(\scanline[71][5] ),
    .X(net6316));
 sg13g2_dlygate4sd3_1 hold1930 (.A(\scanline[1][1] ),
    .X(net6317));
 sg13g2_dlygate4sd3_1 hold1931 (.A(\atari2600.ram[99][0] ),
    .X(net6318));
 sg13g2_dlygate4sd3_1 hold1932 (.A(\scanline[40][5] ),
    .X(net6319));
 sg13g2_dlygate4sd3_1 hold1933 (.A(\scanline[3][3] ),
    .X(net6320));
 sg13g2_dlygate4sd3_1 hold1934 (.A(\scanline[68][4] ),
    .X(net6321));
 sg13g2_dlygate4sd3_1 hold1935 (.A(\scanline[42][6] ),
    .X(net6322));
 sg13g2_dlygate4sd3_1 hold1936 (.A(\atari2600.input_switches[3] ),
    .X(net6323));
 sg13g2_dlygate4sd3_1 hold1937 (.A(_02301_),
    .X(net6324));
 sg13g2_dlygate4sd3_1 hold1938 (.A(\atari2600.ram[33][1] ),
    .X(net6325));
 sg13g2_dlygate4sd3_1 hold1939 (.A(\scanline[131][2] ),
    .X(net6326));
 sg13g2_dlygate4sd3_1 hold1940 (.A(\scanline[84][1] ),
    .X(net6327));
 sg13g2_dlygate4sd3_1 hold1941 (.A(\scanline[8][1] ),
    .X(net6328));
 sg13g2_dlygate4sd3_1 hold1942 (.A(\scanline[4][6] ),
    .X(net6329));
 sg13g2_dlygate4sd3_1 hold1943 (.A(\atari2600.cpu.ABH[7] ),
    .X(net6330));
 sg13g2_dlygate4sd3_1 hold1944 (.A(_02984_),
    .X(net6331));
 sg13g2_dlygate4sd3_1 hold1945 (.A(\atari2600.ram[68][6] ),
    .X(net6332));
 sg13g2_dlygate4sd3_1 hold1946 (.A(\atari2600.ram[83][3] ),
    .X(net6333));
 sg13g2_dlygate4sd3_1 hold1947 (.A(\scanline[145][2] ),
    .X(net6334));
 sg13g2_dlygate4sd3_1 hold1948 (.A(\atari2600.ram[104][5] ),
    .X(net6335));
 sg13g2_dlygate4sd3_1 hold1949 (.A(\atari2600.ram[51][0] ),
    .X(net6336));
 sg13g2_dlygate4sd3_1 hold1950 (.A(\scanline[33][5] ),
    .X(net6337));
 sg13g2_dlygate4sd3_1 hold1951 (.A(\scanline[132][2] ),
    .X(net6338));
 sg13g2_dlygate4sd3_1 hold1952 (.A(\atari2600.ram[60][1] ),
    .X(net6339));
 sg13g2_dlygate4sd3_1 hold1953 (.A(\atari2600.ram[124][2] ),
    .X(net6340));
 sg13g2_dlygate4sd3_1 hold1954 (.A(\scanline[80][6] ),
    .X(net6341));
 sg13g2_dlygate4sd3_1 hold1955 (.A(\scanline[68][3] ),
    .X(net6342));
 sg13g2_dlygate4sd3_1 hold1956 (.A(\atari2600.ram[67][1] ),
    .X(net6343));
 sg13g2_dlygate4sd3_1 hold1957 (.A(\atari2600.ram[13][5] ),
    .X(net6344));
 sg13g2_dlygate4sd3_1 hold1958 (.A(\atari2600.pia.reset_timer[4] ),
    .X(net6345));
 sg13g2_dlygate4sd3_1 hold1959 (.A(\atari2600.ram[105][4] ),
    .X(net6346));
 sg13g2_dlygate4sd3_1 hold1960 (.A(\atari2600.ram[17][5] ),
    .X(net6347));
 sg13g2_dlygate4sd3_1 hold1961 (.A(\atari2600.ram[51][1] ),
    .X(net6348));
 sg13g2_dlygate4sd3_1 hold1962 (.A(\scanline[1][4] ),
    .X(net6349));
 sg13g2_dlygate4sd3_1 hold1963 (.A(\scanline[16][2] ),
    .X(net6350));
 sg13g2_dlygate4sd3_1 hold1964 (.A(\atari2600.ram[20][3] ),
    .X(net6351));
 sg13g2_dlygate4sd3_1 hold1965 (.A(\scanline[8][0] ),
    .X(net6352));
 sg13g2_dlygate4sd3_1 hold1966 (.A(\scanline[19][6] ),
    .X(net6353));
 sg13g2_dlygate4sd3_1 hold1967 (.A(\atari2600.ram[15][2] ),
    .X(net6354));
 sg13g2_dlygate4sd3_1 hold1968 (.A(\atari2600.ram[7][0] ),
    .X(net6355));
 sg13g2_dlygate4sd3_1 hold1969 (.A(\scanline[50][2] ),
    .X(net6356));
 sg13g2_dlygate4sd3_1 hold1970 (.A(\scanline[100][2] ),
    .X(net6357));
 sg13g2_dlygate4sd3_1 hold1971 (.A(\atari2600.ram[32][0] ),
    .X(net6358));
 sg13g2_dlygate4sd3_1 hold1972 (.A(\scanline[108][1] ),
    .X(net6359));
 sg13g2_dlygate4sd3_1 hold1973 (.A(\atari2600.ram[60][3] ),
    .X(net6360));
 sg13g2_dlygate4sd3_1 hold1974 (.A(\scanline[116][1] ),
    .X(net6361));
 sg13g2_dlygate4sd3_1 hold1975 (.A(\scanline[74][2] ),
    .X(net6362));
 sg13g2_dlygate4sd3_1 hold1976 (.A(\scanline[128][2] ),
    .X(net6363));
 sg13g2_dlygate4sd3_1 hold1977 (.A(\scanline[100][0] ),
    .X(net6364));
 sg13g2_dlygate4sd3_1 hold1978 (.A(\atari2600.ram[115][3] ),
    .X(net6365));
 sg13g2_dlygate4sd3_1 hold1979 (.A(\scanline[134][2] ),
    .X(net6366));
 sg13g2_dlygate4sd3_1 hold1980 (.A(\scanline[104][2] ),
    .X(net6367));
 sg13g2_dlygate4sd3_1 hold1981 (.A(\atari2600.ram[53][2] ),
    .X(net6368));
 sg13g2_dlygate4sd3_1 hold1982 (.A(\atari2600.ram[41][6] ),
    .X(net6369));
 sg13g2_dlygate4sd3_1 hold1983 (.A(\atari2600.ram[43][4] ),
    .X(net6370));
 sg13g2_dlygate4sd3_1 hold1984 (.A(\scanline[32][4] ),
    .X(net6371));
 sg13g2_dlygate4sd3_1 hold1985 (.A(\atari2600.cpu.AXYS[0][5] ),
    .X(net6372));
 sg13g2_dlygate4sd3_1 hold1986 (.A(\scanline[133][2] ),
    .X(net6373));
 sg13g2_dlygate4sd3_1 hold1987 (.A(\scanline[40][0] ),
    .X(net6374));
 sg13g2_dlygate4sd3_1 hold1988 (.A(\scanline[17][4] ),
    .X(net6375));
 sg13g2_dlygate4sd3_1 hold1989 (.A(\scanline[70][4] ),
    .X(net6376));
 sg13g2_dlygate4sd3_1 hold1990 (.A(\scanline[65][1] ),
    .X(net6377));
 sg13g2_dlygate4sd3_1 hold1991 (.A(\atari2600.ram[31][0] ),
    .X(net6378));
 sg13g2_dlygate4sd3_1 hold1992 (.A(\scanline[71][1] ),
    .X(net6379));
 sg13g2_dlygate4sd3_1 hold1993 (.A(\scanline[72][2] ),
    .X(net6380));
 sg13g2_dlygate4sd3_1 hold1994 (.A(\scanline[41][3] ),
    .X(net6381));
 sg13g2_dlygate4sd3_1 hold1995 (.A(\scanline[0][2] ),
    .X(net6382));
 sg13g2_dlygate4sd3_1 hold1996 (.A(\scanline[10][1] ),
    .X(net6383));
 sg13g2_dlygate4sd3_1 hold1997 (.A(\scanline[72][5] ),
    .X(net6384));
 sg13g2_dlygate4sd3_1 hold1998 (.A(\scanline[40][4] ),
    .X(net6385));
 sg13g2_dlygate4sd3_1 hold1999 (.A(\scanline[28][2] ),
    .X(net6386));
 sg13g2_dlygate4sd3_1 hold2000 (.A(\scanline[132][3] ),
    .X(net6387));
 sg13g2_dlygate4sd3_1 hold2001 (.A(\atari2600.ram[43][5] ),
    .X(net6388));
 sg13g2_dlygate4sd3_1 hold2002 (.A(\scanline[42][5] ),
    .X(net6389));
 sg13g2_dlygate4sd3_1 hold2003 (.A(\scanline[60][4] ),
    .X(net6390));
 sg13g2_dlygate4sd3_1 hold2004 (.A(\atari2600.ram[118][6] ),
    .X(net6391));
 sg13g2_dlygate4sd3_1 hold2005 (.A(\atari2600.ram[47][6] ),
    .X(net6392));
 sg13g2_dlygate4sd3_1 hold2006 (.A(\atari2600.ram[25][3] ),
    .X(net6393));
 sg13g2_dlygate4sd3_1 hold2007 (.A(\scanline[66][5] ),
    .X(net6394));
 sg13g2_dlygate4sd3_1 hold2008 (.A(\atari2600.ram[99][5] ),
    .X(net6395));
 sg13g2_dlygate4sd3_1 hold2009 (.A(\scanline[145][5] ),
    .X(net6396));
 sg13g2_dlygate4sd3_1 hold2010 (.A(\scanline[75][2] ),
    .X(net6397));
 sg13g2_dlygate4sd3_1 hold2011 (.A(_00144_),
    .X(net6398));
 sg13g2_dlygate4sd3_1 hold2012 (.A(\atari2600.ram[37][5] ),
    .X(net6399));
 sg13g2_dlygate4sd3_1 hold2013 (.A(\atari2600.ram[52][6] ),
    .X(net6400));
 sg13g2_dlygate4sd3_1 hold2014 (.A(\scanline[34][6] ),
    .X(net6401));
 sg13g2_dlygate4sd3_1 hold2015 (.A(\scanline[18][2] ),
    .X(net6402));
 sg13g2_dlygate4sd3_1 hold2016 (.A(\atari2600.ram[51][7] ),
    .X(net6403));
 sg13g2_dlygate4sd3_1 hold2017 (.A(\atari2600.cpu.IRHOLD[5] ),
    .X(net6404));
 sg13g2_dlygate4sd3_1 hold2018 (.A(\scanline[49][6] ),
    .X(net6405));
 sg13g2_dlygate4sd3_1 hold2019 (.A(\scanline[73][4] ),
    .X(net6406));
 sg13g2_dlygate4sd3_1 hold2020 (.A(\scanline[136][1] ),
    .X(net6407));
 sg13g2_dlygate4sd3_1 hold2021 (.A(\atari2600.ram[98][4] ),
    .X(net6408));
 sg13g2_dlygate4sd3_1 hold2022 (.A(\atari2600.ram[12][6] ),
    .X(net6409));
 sg13g2_dlygate4sd3_1 hold2023 (.A(\atari2600.ram[41][3] ),
    .X(net6410));
 sg13g2_dlygate4sd3_1 hold2024 (.A(\scanline[132][5] ),
    .X(net6411));
 sg13g2_dlygate4sd3_1 hold2025 (.A(\scanline[133][6] ),
    .X(net6412));
 sg13g2_dlygate4sd3_1 hold2026 (.A(\scanline[104][1] ),
    .X(net6413));
 sg13g2_dlygate4sd3_1 hold2027 (.A(\atari2600.ram[27][1] ),
    .X(net6414));
 sg13g2_dlygate4sd3_1 hold2028 (.A(\scanline[16][3] ),
    .X(net6415));
 sg13g2_dlygate4sd3_1 hold2029 (.A(\scanline[49][5] ),
    .X(net6416));
 sg13g2_dlygate4sd3_1 hold2030 (.A(\scanline[138][1] ),
    .X(net6417));
 sg13g2_dlygate4sd3_1 hold2031 (.A(\atari2600.pia.reset_timer[6] ),
    .X(net6418));
 sg13g2_dlygate4sd3_1 hold2032 (.A(\atari2600.ram[35][7] ),
    .X(net6419));
 sg13g2_dlygate4sd3_1 hold2033 (.A(\atari2600.ram[33][0] ),
    .X(net6420));
 sg13g2_dlygate4sd3_1 hold2034 (.A(\atari2600.ram[5][3] ),
    .X(net6421));
 sg13g2_dlygate4sd3_1 hold2035 (.A(\atari2600.ram[115][4] ),
    .X(net6422));
 sg13g2_dlygate4sd3_1 hold2036 (.A(\atari2600.ram[69][3] ),
    .X(net6423));
 sg13g2_dlygate4sd3_1 hold2037 (.A(\atari2600.ram[103][7] ),
    .X(net6424));
 sg13g2_dlygate4sd3_1 hold2038 (.A(\scanline[139][6] ),
    .X(net6425));
 sg13g2_dlygate4sd3_1 hold2039 (.A(\atari2600.ram[63][3] ),
    .X(net6426));
 sg13g2_dlygate4sd3_1 hold2040 (.A(\atari2600.ram[65][5] ),
    .X(net6427));
 sg13g2_dlygate4sd3_1 hold2041 (.A(\scanline[0][3] ),
    .X(net6428));
 sg13g2_dlygate4sd3_1 hold2042 (.A(\atari2600.ram[13][6] ),
    .X(net6429));
 sg13g2_dlygate4sd3_1 hold2043 (.A(\scanline[48][3] ),
    .X(net6430));
 sg13g2_dlygate4sd3_1 hold2044 (.A(\atari2600.ram[19][6] ),
    .X(net6431));
 sg13g2_dlygate4sd3_1 hold2045 (.A(\scanline[120][5] ),
    .X(net6432));
 sg13g2_dlygate4sd3_1 hold2046 (.A(\scanline[42][3] ),
    .X(net6433));
 sg13g2_dlygate4sd3_1 hold2047 (.A(\atari2600.ram[119][4] ),
    .X(net6434));
 sg13g2_dlygate4sd3_1 hold2048 (.A(\scanline[108][2] ),
    .X(net6435));
 sg13g2_dlygate4sd3_1 hold2049 (.A(\scanline[2][1] ),
    .X(net6436));
 sg13g2_dlygate4sd3_1 hold2050 (.A(\atari2600.ram[123][7] ),
    .X(net6437));
 sg13g2_dlygate4sd3_1 hold2051 (.A(\scanline[4][5] ),
    .X(net6438));
 sg13g2_dlygate4sd3_1 hold2052 (.A(\atari2600.ram[13][4] ),
    .X(net6439));
 sg13g2_dlygate4sd3_1 hold2053 (.A(\scanline[28][4] ),
    .X(net6440));
 sg13g2_dlygate4sd3_1 hold2054 (.A(\scanline[52][4] ),
    .X(net6441));
 sg13g2_dlygate4sd3_1 hold2055 (.A(\atari2600.ram[37][0] ),
    .X(net6442));
 sg13g2_dlygate4sd3_1 hold2056 (.A(\scanline[20][6] ),
    .X(net6443));
 sg13g2_dlygate4sd3_1 hold2057 (.A(\scanline[112][4] ),
    .X(net6444));
 sg13g2_dlygate4sd3_1 hold2058 (.A(\atari2600.ram[57][6] ),
    .X(net6445));
 sg13g2_dlygate4sd3_1 hold2059 (.A(\atari2600.ram[15][5] ),
    .X(net6446));
 sg13g2_dlygate4sd3_1 hold2060 (.A(\scanline[128][5] ),
    .X(net6447));
 sg13g2_dlygate4sd3_1 hold2061 (.A(\scanline[82][1] ),
    .X(net6448));
 sg13g2_dlygate4sd3_1 hold2062 (.A(\scanline[137][6] ),
    .X(net6449));
 sg13g2_dlygate4sd3_1 hold2063 (.A(\scanline[25][3] ),
    .X(net6450));
 sg13g2_dlygate4sd3_1 hold2064 (.A(\scanline[32][6] ),
    .X(net6451));
 sg13g2_dlygate4sd3_1 hold2065 (.A(\scanline[72][1] ),
    .X(net6452));
 sg13g2_dlygate4sd3_1 hold2066 (.A(\scanline[9][2] ),
    .X(net6453));
 sg13g2_dlygate4sd3_1 hold2067 (.A(\atari2600.ram[21][0] ),
    .X(net6454));
 sg13g2_dlygate4sd3_1 hold2068 (.A(\atari2600.cpu.AXYS[3][6] ),
    .X(net6455));
 sg13g2_dlygate4sd3_1 hold2069 (.A(\atari2600.ram[71][1] ),
    .X(net6456));
 sg13g2_dlygate4sd3_1 hold2070 (.A(\atari2600.ram[55][6] ),
    .X(net6457));
 sg13g2_dlygate4sd3_1 hold2071 (.A(\atari2600.ram[33][3] ),
    .X(net6458));
 sg13g2_dlygate4sd3_1 hold2072 (.A(\scanline[48][4] ),
    .X(net6459));
 sg13g2_dlygate4sd3_1 hold2073 (.A(\scanline[19][1] ),
    .X(net6460));
 sg13g2_dlygate4sd3_1 hold2074 (.A(\scanline[132][6] ),
    .X(net6461));
 sg13g2_dlygate4sd3_1 hold2075 (.A(\scanline[146][5] ),
    .X(net6462));
 sg13g2_dlygate4sd3_1 hold2076 (.A(\scanline[146][6] ),
    .X(net6463));
 sg13g2_dlygate4sd3_1 hold2077 (.A(\atari2600.ram[0][7] ),
    .X(net6464));
 sg13g2_dlygate4sd3_1 hold2078 (.A(\scanline[38][2] ),
    .X(net6465));
 sg13g2_dlygate4sd3_1 hold2079 (.A(\scanline[52][3] ),
    .X(net6466));
 sg13g2_dlygate4sd3_1 hold2080 (.A(\atari2600.ram[121][4] ),
    .X(net6467));
 sg13g2_dlygate4sd3_1 hold2081 (.A(\atari2600.ram[11][2] ),
    .X(net6468));
 sg13g2_dlygate4sd3_1 hold2082 (.A(\scanline[108][0] ),
    .X(net6469));
 sg13g2_dlygate4sd3_1 hold2083 (.A(\atari2600.ram[67][3] ),
    .X(net6470));
 sg13g2_dlygate4sd3_1 hold2084 (.A(\atari2600.ram[23][5] ),
    .X(net6471));
 sg13g2_dlygate4sd3_1 hold2085 (.A(\atari2600.ram[9][2] ),
    .X(net6472));
 sg13g2_dlygate4sd3_1 hold2086 (.A(\atari2600.ram[87][2] ),
    .X(net6473));
 sg13g2_dlygate4sd3_1 hold2087 (.A(\atari2600.ram[47][5] ),
    .X(net6474));
 sg13g2_dlygate4sd3_1 hold2088 (.A(\scanline[64][4] ),
    .X(net6475));
 sg13g2_dlygate4sd3_1 hold2089 (.A(\scanline[82][4] ),
    .X(net6476));
 sg13g2_dlygate4sd3_1 hold2090 (.A(\scanline[48][1] ),
    .X(net6477));
 sg13g2_dlygate4sd3_1 hold2091 (.A(\atari2600.ram[96][0] ),
    .X(net6478));
 sg13g2_dlygate4sd3_1 hold2092 (.A(\atari2600.ram[116][0] ),
    .X(net6479));
 sg13g2_dlygate4sd3_1 hold2093 (.A(\scanline[27][3] ),
    .X(net6480));
 sg13g2_dlygate4sd3_1 hold2094 (.A(\scanline[73][5] ),
    .X(net6481));
 sg13g2_dlygate4sd3_1 hold2095 (.A(\atari2600.cpu.AXYS[2][7] ),
    .X(net6482));
 sg13g2_dlygate4sd3_1 hold2096 (.A(\scanline[92][2] ),
    .X(net6483));
 sg13g2_dlygate4sd3_1 hold2097 (.A(\atari2600.ram[7][6] ),
    .X(net6484));
 sg13g2_dlygate4sd3_1 hold2098 (.A(\scanline[146][1] ),
    .X(net6485));
 sg13g2_dlygate4sd3_1 hold2099 (.A(\scanline[23][3] ),
    .X(net6486));
 sg13g2_dlygate4sd3_1 hold2100 (.A(\atari2600.ram[117][5] ),
    .X(net6487));
 sg13g2_dlygate4sd3_1 hold2101 (.A(\scanline[97][2] ),
    .X(net6488));
 sg13g2_dlygate4sd3_1 hold2102 (.A(\scanline[74][4] ),
    .X(net6489));
 sg13g2_dlygate4sd3_1 hold2103 (.A(\scanline[50][3] ),
    .X(net6490));
 sg13g2_dlygate4sd3_1 hold2104 (.A(\scanline[108][3] ),
    .X(net6491));
 sg13g2_dlygate4sd3_1 hold2105 (.A(\atari2600.ram[69][5] ),
    .X(net6492));
 sg13g2_dlygate4sd3_1 hold2106 (.A(\scanline[39][4] ),
    .X(net6493));
 sg13g2_dlygate4sd3_1 hold2107 (.A(\atari2600.ram[119][3] ),
    .X(net6494));
 sg13g2_dlygate4sd3_1 hold2108 (.A(\atari2600.ram[107][1] ),
    .X(net6495));
 sg13g2_dlygate4sd3_1 hold2109 (.A(\scanline[36][3] ),
    .X(net6496));
 sg13g2_dlygate4sd3_1 hold2110 (.A(\scanline[7][0] ),
    .X(net6497));
 sg13g2_dlygate4sd3_1 hold2111 (.A(\scanline[81][1] ),
    .X(net6498));
 sg13g2_dlygate4sd3_1 hold2112 (.A(\scanline[64][5] ),
    .X(net6499));
 sg13g2_dlygate4sd3_1 hold2113 (.A(\scanline[139][3] ),
    .X(net6500));
 sg13g2_dlygate4sd3_1 hold2114 (.A(\atari2600.ram[19][2] ),
    .X(net6501));
 sg13g2_dlygate4sd3_1 hold2115 (.A(\scanline[44][6] ),
    .X(net6502));
 sg13g2_dlygate4sd3_1 hold2116 (.A(\scanline[50][0] ),
    .X(net6503));
 sg13g2_dlygate4sd3_1 hold2117 (.A(\atari2600.ram[119][0] ),
    .X(net6504));
 sg13g2_dlygate4sd3_1 hold2118 (.A(\scanline[6][4] ),
    .X(net6505));
 sg13g2_dlygate4sd3_1 hold2119 (.A(\scanline[27][0] ),
    .X(net6506));
 sg13g2_dlygate4sd3_1 hold2120 (.A(\scanline[32][2] ),
    .X(net6507));
 sg13g2_dlygate4sd3_1 hold2121 (.A(\atari2600.ram[107][4] ),
    .X(net6508));
 sg13g2_dlygate4sd3_1 hold2122 (.A(\atari2600.ram[52][1] ),
    .X(net6509));
 sg13g2_dlygate4sd3_1 hold2123 (.A(\scanline[10][5] ),
    .X(net6510));
 sg13g2_dlygate4sd3_1 hold2124 (.A(\scanline[73][1] ),
    .X(net6511));
 sg13g2_dlygate4sd3_1 hold2125 (.A(\atari2600.ram[107][0] ),
    .X(net6512));
 sg13g2_dlygate4sd3_1 hold2126 (.A(\atari2600.ram[115][6] ),
    .X(net6513));
 sg13g2_dlygate4sd3_1 hold2127 (.A(\scanline[138][5] ),
    .X(net6514));
 sg13g2_dlygate4sd3_1 hold2128 (.A(\scanline[34][4] ),
    .X(net6515));
 sg13g2_dlygate4sd3_1 hold2129 (.A(\atari2600.ram[113][0] ),
    .X(net6516));
 sg13g2_dlygate4sd3_1 hold2130 (.A(\scanline[68][5] ),
    .X(net6517));
 sg13g2_dlygate4sd3_1 hold2131 (.A(\scanline[104][5] ),
    .X(net6518));
 sg13g2_dlygate4sd3_1 hold2132 (.A(\atari2600.ram[67][7] ),
    .X(net6519));
 sg13g2_dlygate4sd3_1 hold2133 (.A(\scanline[75][0] ),
    .X(net6520));
 sg13g2_dlygate4sd3_1 hold2134 (.A(\atari2600.ram[123][6] ),
    .X(net6521));
 sg13g2_dlygate4sd3_1 hold2135 (.A(\scanline[41][2] ),
    .X(net6522));
 sg13g2_dlygate4sd3_1 hold2136 (.A(\atari2600.ram[81][5] ),
    .X(net6523));
 sg13g2_dlygate4sd3_1 hold2137 (.A(\scanline[129][4] ),
    .X(net6524));
 sg13g2_dlygate4sd3_1 hold2138 (.A(\scanline[16][4] ),
    .X(net6525));
 sg13g2_dlygate4sd3_1 hold2139 (.A(\atari2600.ram[83][6] ),
    .X(net6526));
 sg13g2_dlygate4sd3_1 hold2140 (.A(\atari2600.ram[107][7] ),
    .X(net6527));
 sg13g2_dlygate4sd3_1 hold2141 (.A(\scanline[116][5] ),
    .X(net6528));
 sg13g2_dlygate4sd3_1 hold2142 (.A(\scanline[2][0] ),
    .X(net6529));
 sg13g2_dlygate4sd3_1 hold2143 (.A(\scanline[0][6] ),
    .X(net6530));
 sg13g2_dlygate4sd3_1 hold2144 (.A(\scanline[76][2] ),
    .X(net6531));
 sg13g2_dlygate4sd3_1 hold2145 (.A(\scanline[23][1] ),
    .X(net6532));
 sg13g2_dlygate4sd3_1 hold2146 (.A(\scanline[7][3] ),
    .X(net6533));
 sg13g2_dlygate4sd3_1 hold2147 (.A(\atari2600.pia.time_counter[19] ),
    .X(net6534));
 sg13g2_dlygate4sd3_1 hold2148 (.A(_01791_),
    .X(net6535));
 sg13g2_dlygate4sd3_1 hold2149 (.A(\scanline[52][1] ),
    .X(net6536));
 sg13g2_dlygate4sd3_1 hold2150 (.A(\scanline[128][6] ),
    .X(net6537));
 sg13g2_dlygate4sd3_1 hold2151 (.A(\atari2600.pia.reset_timer[0] ),
    .X(net6538));
 sg13g2_dlygate4sd3_1 hold2152 (.A(\scanline[140][3] ),
    .X(net6539));
 sg13g2_dlygate4sd3_1 hold2153 (.A(\scanline[37][2] ),
    .X(net6540));
 sg13g2_dlygate4sd3_1 hold2154 (.A(\scanline[23][2] ),
    .X(net6541));
 sg13g2_dlygate4sd3_1 hold2155 (.A(\scanline[140][2] ),
    .X(net6542));
 sg13g2_dlygate4sd3_1 hold2156 (.A(\scanline[70][5] ),
    .X(net6543));
 sg13g2_dlygate4sd3_1 hold2157 (.A(\scanline[50][1] ),
    .X(net6544));
 sg13g2_dlygate4sd3_1 hold2158 (.A(\scanline[23][5] ),
    .X(net6545));
 sg13g2_dlygate4sd3_1 hold2159 (.A(\atari2600.ram[43][2] ),
    .X(net6546));
 sg13g2_dlygate4sd3_1 hold2160 (.A(\scanline[67][1] ),
    .X(net6547));
 sg13g2_dlygate4sd3_1 hold2161 (.A(\scanline[152][3] ),
    .X(net6548));
 sg13g2_dlygate4sd3_1 hold2162 (.A(\scanline[66][1] ),
    .X(net6549));
 sg13g2_dlygate4sd3_1 hold2163 (.A(\atari2600.cpu.AXYS[0][6] ),
    .X(net6550));
 sg13g2_dlygate4sd3_1 hold2164 (.A(\scanline[146][2] ),
    .X(net6551));
 sg13g2_dlygate4sd3_1 hold2165 (.A(\atari2600.ram[23][6] ),
    .X(net6552));
 sg13g2_dlygate4sd3_1 hold2166 (.A(\atari2600.ram[127][4] ),
    .X(net6553));
 sg13g2_dlygate4sd3_1 hold2167 (.A(\scanline[68][1] ),
    .X(net6554));
 sg13g2_dlygate4sd3_1 hold2168 (.A(\atari2600.ram[19][7] ),
    .X(net6555));
 sg13g2_dlygate4sd3_1 hold2169 (.A(\atari2600.ram[105][0] ),
    .X(net6556));
 sg13g2_dlygate4sd3_1 hold2170 (.A(\scanline[74][5] ),
    .X(net6557));
 sg13g2_dlygate4sd3_1 hold2171 (.A(\scanline[43][0] ),
    .X(net6558));
 sg13g2_dlygate4sd3_1 hold2172 (.A(\scanline[28][1] ),
    .X(net6559));
 sg13g2_dlygate4sd3_1 hold2173 (.A(\atari2600.ram[112][2] ),
    .X(net6560));
 sg13g2_dlygate4sd3_1 hold2174 (.A(\scanline[73][6] ),
    .X(net6561));
 sg13g2_dlygate4sd3_1 hold2175 (.A(\scanline[97][3] ),
    .X(net6562));
 sg13g2_dlygate4sd3_1 hold2176 (.A(\atari2600.ram[97][1] ),
    .X(net6563));
 sg13g2_dlygate4sd3_1 hold2177 (.A(\atari2600.ram[27][5] ),
    .X(net6564));
 sg13g2_dlygate4sd3_1 hold2178 (.A(\scanline[2][5] ),
    .X(net6565));
 sg13g2_dlygate4sd3_1 hold2179 (.A(\atari2600.ram[13][3] ),
    .X(net6566));
 sg13g2_dlygate4sd3_1 hold2180 (.A(\scanline[82][2] ),
    .X(net6567));
 sg13g2_dlygate4sd3_1 hold2181 (.A(\atari2600.ram[85][6] ),
    .X(net6568));
 sg13g2_dlygate4sd3_1 hold2182 (.A(\atari2600.ram[7][3] ),
    .X(net6569));
 sg13g2_dlygate4sd3_1 hold2183 (.A(\scanline[133][1] ),
    .X(net6570));
 sg13g2_dlygate4sd3_1 hold2184 (.A(\atari2600.ram[43][7] ),
    .X(net6571));
 sg13g2_dlygate4sd3_1 hold2185 (.A(\atari2600.ram[64][7] ),
    .X(net6572));
 sg13g2_dlygate4sd3_1 hold2186 (.A(\scanline[27][2] ),
    .X(net6573));
 sg13g2_dlygate4sd3_1 hold2187 (.A(\scanline[42][2] ),
    .X(net6574));
 sg13g2_dlygate4sd3_1 hold2188 (.A(\atari2600.ram[100][1] ),
    .X(net6575));
 sg13g2_dlygate4sd3_1 hold2189 (.A(\scanline[43][3] ),
    .X(net6576));
 sg13g2_dlygate4sd3_1 hold2190 (.A(\scanline[26][4] ),
    .X(net6577));
 sg13g2_dlygate4sd3_1 hold2191 (.A(\atari2600.ram[121][2] ),
    .X(net6578));
 sg13g2_dlygate4sd3_1 hold2192 (.A(\scanline[72][0] ),
    .X(net6579));
 sg13g2_dlygate4sd3_1 hold2193 (.A(\atari2600.ram[33][5] ),
    .X(net6580));
 sg13g2_dlygate4sd3_1 hold2194 (.A(\atari2600.cpu.PC[13] ),
    .X(net6581));
 sg13g2_dlygate4sd3_1 hold2195 (.A(_02511_),
    .X(net6582));
 sg13g2_dlygate4sd3_1 hold2196 (.A(\scanline[66][6] ),
    .X(net6583));
 sg13g2_dlygate4sd3_1 hold2197 (.A(\scanline[33][0] ),
    .X(net6584));
 sg13g2_dlygate4sd3_1 hold2198 (.A(\scanline[152][5] ),
    .X(net6585));
 sg13g2_dlygate4sd3_1 hold2199 (.A(\scanline[6][5] ),
    .X(net6586));
 sg13g2_dlygate4sd3_1 hold2200 (.A(\scanline[1][3] ),
    .X(net6587));
 sg13g2_dlygate4sd3_1 hold2201 (.A(\atari2600.ram[16][3] ),
    .X(net6588));
 sg13g2_dlygate4sd3_1 hold2202 (.A(\scanline[73][0] ),
    .X(net6589));
 sg13g2_dlygate4sd3_1 hold2203 (.A(\scanline[69][0] ),
    .X(net6590));
 sg13g2_dlygate4sd3_1 hold2204 (.A(\scanline[139][1] ),
    .X(net6591));
 sg13g2_dlygate4sd3_1 hold2205 (.A(\scanline[26][0] ),
    .X(net6592));
 sg13g2_dlygate4sd3_1 hold2206 (.A(\atari2600.ram[102][7] ),
    .X(net6593));
 sg13g2_dlygate4sd3_1 hold2207 (.A(\scanline[88][2] ),
    .X(net6594));
 sg13g2_dlygate4sd3_1 hold2208 (.A(\scanline[70][3] ),
    .X(net6595));
 sg13g2_dlygate4sd3_1 hold2209 (.A(\scanline[37][6] ),
    .X(net6596));
 sg13g2_dlygate4sd3_1 hold2210 (.A(\scanline[68][2] ),
    .X(net6597));
 sg13g2_dlygate4sd3_1 hold2211 (.A(\atari2600.ram[37][6] ),
    .X(net6598));
 sg13g2_dlygate4sd3_1 hold2212 (.A(\atari2600.pia.dat_o[4] ),
    .X(net6599));
 sg13g2_dlygate4sd3_1 hold2213 (.A(_07157_),
    .X(net6600));
 sg13g2_dlygate4sd3_1 hold2214 (.A(\atari2600.ram[51][3] ),
    .X(net6601));
 sg13g2_dlygate4sd3_1 hold2215 (.A(\scanline[10][0] ),
    .X(net6602));
 sg13g2_dlygate4sd3_1 hold2216 (.A(\scanline[49][4] ),
    .X(net6603));
 sg13g2_dlygate4sd3_1 hold2217 (.A(\scanline[18][0] ),
    .X(net6604));
 sg13g2_dlygate4sd3_1 hold2218 (.A(\scanline[69][3] ),
    .X(net6605));
 sg13g2_dlygate4sd3_1 hold2219 (.A(\scanline[64][3] ),
    .X(net6606));
 sg13g2_dlygate4sd3_1 hold2220 (.A(\atari2600.ram[123][5] ),
    .X(net6607));
 sg13g2_dlygate4sd3_1 hold2221 (.A(\scanline[145][4] ),
    .X(net6608));
 sg13g2_dlygate4sd3_1 hold2222 (.A(\scanline[23][4] ),
    .X(net6609));
 sg13g2_dlygate4sd3_1 hold2223 (.A(\atari2600.ram[40][5] ),
    .X(net6610));
 sg13g2_dlygate4sd3_1 hold2224 (.A(\scanline[35][2] ),
    .X(net6611));
 sg13g2_dlygate4sd3_1 hold2225 (.A(\scanline[116][6] ),
    .X(net6612));
 sg13g2_dlygate4sd3_1 hold2226 (.A(\scanline[138][4] ),
    .X(net6613));
 sg13g2_dlygate4sd3_1 hold2227 (.A(\scanline[44][2] ),
    .X(net6614));
 sg13g2_dlygate4sd3_1 hold2228 (.A(\atari2600.ram[36][3] ),
    .X(net6615));
 sg13g2_dlygate4sd3_1 hold2229 (.A(\scanline[156][0] ),
    .X(net6616));
 sg13g2_dlygate4sd3_1 hold2230 (.A(\scanline[5][1] ),
    .X(net6617));
 sg13g2_dlygate4sd3_1 hold2231 (.A(\rom_last_read_addr[3] ),
    .X(net6618));
 sg13g2_dlygate4sd3_1 hold2232 (.A(_01129_),
    .X(net6619));
 sg13g2_dlygate4sd3_1 hold2233 (.A(\atari2600.ram[47][0] ),
    .X(net6620));
 sg13g2_dlygate4sd3_1 hold2234 (.A(\scanline[11][0] ),
    .X(net6621));
 sg13g2_dlygate4sd3_1 hold2235 (.A(\scanline[43][5] ),
    .X(net6622));
 sg13g2_dlygate4sd3_1 hold2236 (.A(\scanline[76][5] ),
    .X(net6623));
 sg13g2_dlygate4sd3_1 hold2237 (.A(\scanline[97][5] ),
    .X(net6624));
 sg13g2_dlygate4sd3_1 hold2238 (.A(\scanline[64][6] ),
    .X(net6625));
 sg13g2_dlygate4sd3_1 hold2239 (.A(\atari2600.ram[32][5] ),
    .X(net6626));
 sg13g2_dlygate4sd3_1 hold2240 (.A(\scanline[75][1] ),
    .X(net6627));
 sg13g2_dlygate4sd3_1 hold2241 (.A(\atari2600.ram[107][2] ),
    .X(net6628));
 sg13g2_dlygate4sd3_1 hold2242 (.A(\scanline[17][6] ),
    .X(net6629));
 sg13g2_dlygate4sd3_1 hold2243 (.A(\scanline[69][4] ),
    .X(net6630));
 sg13g2_dlygate4sd3_1 hold2244 (.A(\atari2600.ram[13][1] ),
    .X(net6631));
 sg13g2_dlygate4sd3_1 hold2245 (.A(\scanline[156][4] ),
    .X(net6632));
 sg13g2_dlygate4sd3_1 hold2246 (.A(\atari2600.ram[107][5] ),
    .X(net6633));
 sg13g2_dlygate4sd3_1 hold2247 (.A(\atari2600.cpu.IRHOLD[6] ),
    .X(net6634));
 sg13g2_dlygate4sd3_1 hold2248 (.A(\scanline[50][5] ),
    .X(net6635));
 sg13g2_dlygate4sd3_1 hold2249 (.A(\atari2600.ram[15][1] ),
    .X(net6636));
 sg13g2_dlygate4sd3_1 hold2250 (.A(\scanline[136][2] ),
    .X(net6637));
 sg13g2_dlygate4sd3_1 hold2251 (.A(\atari2600.ram[100][7] ),
    .X(net6638));
 sg13g2_dlygate4sd3_1 hold2252 (.A(\scanline[21][6] ),
    .X(net6639));
 sg13g2_dlygate4sd3_1 hold2253 (.A(\atari2600.ram[115][1] ),
    .X(net6640));
 sg13g2_dlygate4sd3_1 hold2254 (.A(\scanline[67][5] ),
    .X(net6641));
 sg13g2_dlygate4sd3_1 hold2255 (.A(\scanline[92][6] ),
    .X(net6642));
 sg13g2_dlygate4sd3_1 hold2256 (.A(\scanline[3][4] ),
    .X(net6643));
 sg13g2_dlygate4sd3_1 hold2257 (.A(\scanline[76][3] ),
    .X(net6644));
 sg13g2_dlygate4sd3_1 hold2258 (.A(\scanline[7][1] ),
    .X(net6645));
 sg13g2_dlygate4sd3_1 hold2259 (.A(\scanline[131][3] ),
    .X(net6646));
 sg13g2_dlygate4sd3_1 hold2260 (.A(\scanline[112][3] ),
    .X(net6647));
 sg13g2_dlygate4sd3_1 hold2261 (.A(\scanline[144][6] ),
    .X(net6648));
 sg13g2_dlygate4sd3_1 hold2262 (.A(\atari2600.ram[84][2] ),
    .X(net6649));
 sg13g2_dlygate4sd3_1 hold2263 (.A(\scanline[75][3] ),
    .X(net6650));
 sg13g2_dlygate4sd3_1 hold2264 (.A(\atari2600.ram[80][0] ),
    .X(net6651));
 sg13g2_dlygate4sd3_1 hold2265 (.A(\scanline[152][0] ),
    .X(net6652));
 sg13g2_dlygate4sd3_1 hold2266 (.A(\scanline[84][4] ),
    .X(net6653));
 sg13g2_dlygate4sd3_1 hold2267 (.A(\scanline[17][0] ),
    .X(net6654));
 sg13g2_dlygate4sd3_1 hold2268 (.A(\atari2600.ram[123][2] ),
    .X(net6655));
 sg13g2_dlygate4sd3_1 hold2269 (.A(\scanline[135][4] ),
    .X(net6656));
 sg13g2_dlygate4sd3_1 hold2270 (.A(\atari2600.ram[7][5] ),
    .X(net6657));
 sg13g2_dlygate4sd3_1 hold2271 (.A(\atari2600.ram[127][3] ),
    .X(net6658));
 sg13g2_dlygate4sd3_1 hold2272 (.A(\atari2600.tia.old_grp1[5] ),
    .X(net6659));
 sg13g2_dlygate4sd3_1 hold2273 (.A(_01825_),
    .X(net6660));
 sg13g2_dlygate4sd3_1 hold2274 (.A(\scanline[98][4] ),
    .X(net6661));
 sg13g2_dlygate4sd3_1 hold2275 (.A(\scanline[130][1] ),
    .X(net6662));
 sg13g2_dlygate4sd3_1 hold2276 (.A(\scanline[136][4] ),
    .X(net6663));
 sg13g2_dlygate4sd3_1 hold2277 (.A(\scanline[66][4] ),
    .X(net6664));
 sg13g2_dlygate4sd3_1 hold2278 (.A(\atari2600.ram[65][6] ),
    .X(net6665));
 sg13g2_dlygate4sd3_1 hold2279 (.A(\scanline[64][0] ),
    .X(net6666));
 sg13g2_dlygate4sd3_1 hold2280 (.A(\scanline[48][5] ),
    .X(net6667));
 sg13g2_dlygate4sd3_1 hold2281 (.A(\scanline[24][4] ),
    .X(net6668));
 sg13g2_dlygate4sd3_1 hold2282 (.A(\scanline[43][4] ),
    .X(net6669));
 sg13g2_dlygate4sd3_1 hold2283 (.A(\atari2600.ram[71][3] ),
    .X(net6670));
 sg13g2_dlygate4sd3_1 hold2284 (.A(\scanline[33][2] ),
    .X(net6671));
 sg13g2_dlygate4sd3_1 hold2285 (.A(\scanline[42][1] ),
    .X(net6672));
 sg13g2_dlygate4sd3_1 hold2286 (.A(\atari2600.cpu.AXYS[2][3] ),
    .X(net6673));
 sg13g2_dlygate4sd3_1 hold2287 (.A(\scanline[22][0] ),
    .X(net6674));
 sg13g2_dlygate4sd3_1 hold2288 (.A(\scanline[26][5] ),
    .X(net6675));
 sg13g2_dlygate4sd3_1 hold2289 (.A(\atari2600.ram[123][4] ),
    .X(net6676));
 sg13g2_dlygate4sd3_1 hold2290 (.A(\scanline[6][6] ),
    .X(net6677));
 sg13g2_dlygate4sd3_1 hold2291 (.A(\atari2600.ram[87][6] ),
    .X(net6678));
 sg13g2_dlygate4sd3_1 hold2292 (.A(\atari2600.ram[59][5] ),
    .X(net6679));
 sg13g2_dlygate4sd3_1 hold2293 (.A(\scanline[65][0] ),
    .X(net6680));
 sg13g2_dlygate4sd3_1 hold2294 (.A(\scanline[3][0] ),
    .X(net6681));
 sg13g2_dlygate4sd3_1 hold2295 (.A(\scanline[41][5] ),
    .X(net6682));
 sg13g2_dlygate4sd3_1 hold2296 (.A(\scanline[144][2] ),
    .X(net6683));
 sg13g2_dlygate4sd3_1 hold2297 (.A(\scanline[8][3] ),
    .X(net6684));
 sg13g2_dlygate4sd3_1 hold2298 (.A(\atari2600.ram[4][2] ),
    .X(net6685));
 sg13g2_dlygate4sd3_1 hold2299 (.A(\atari2600.ram[36][0] ),
    .X(net6686));
 sg13g2_dlygate4sd3_1 hold2300 (.A(\scanline[67][0] ),
    .X(net6687));
 sg13g2_dlygate4sd3_1 hold2301 (.A(\scanline[97][1] ),
    .X(net6688));
 sg13g2_dlygate4sd3_1 hold2302 (.A(\scanline[98][1] ),
    .X(net6689));
 sg13g2_dlygate4sd3_1 hold2303 (.A(\scanline[128][1] ),
    .X(net6690));
 sg13g2_dlygate4sd3_1 hold2304 (.A(\atari2600.ram_data[0] ),
    .X(net6691));
 sg13g2_dlygate4sd3_1 hold2305 (.A(_07148_),
    .X(net6692));
 sg13g2_dlygate4sd3_1 hold2306 (.A(\scanline[22][5] ),
    .X(net6693));
 sg13g2_dlygate4sd3_1 hold2307 (.A(\atari2600.ram[16][5] ),
    .X(net6694));
 sg13g2_dlygate4sd3_1 hold2308 (.A(\scanline[26][2] ),
    .X(net6695));
 sg13g2_dlygate4sd3_1 hold2309 (.A(\atari2600.ram[71][7] ),
    .X(net6696));
 sg13g2_dlygate4sd3_1 hold2310 (.A(\atari2600.ram[124][1] ),
    .X(net6697));
 sg13g2_dlygate4sd3_1 hold2311 (.A(\scanline[5][2] ),
    .X(net6698));
 sg13g2_dlygate4sd3_1 hold2312 (.A(\scanline[112][6] ),
    .X(net6699));
 sg13g2_dlygate4sd3_1 hold2313 (.A(\atari2600.pia.reset_timer[5] ),
    .X(net6700));
 sg13g2_dlygate4sd3_1 hold2314 (.A(\scanline[39][6] ),
    .X(net6701));
 sg13g2_dlygate4sd3_1 hold2315 (.A(\atari2600.ram[113][7] ),
    .X(net6702));
 sg13g2_dlygate4sd3_1 hold2316 (.A(\atari2600.ram[97][0] ),
    .X(net6703));
 sg13g2_dlygate4sd3_1 hold2317 (.A(\scanline[0][1] ),
    .X(net6704));
 sg13g2_dlygate4sd3_1 hold2318 (.A(\scanline[81][4] ),
    .X(net6705));
 sg13g2_dlygate4sd3_1 hold2319 (.A(\scanline[130][0] ),
    .X(net6706));
 sg13g2_dlygate4sd3_1 hold2320 (.A(\atari2600.cpu.AXYS[0][7] ),
    .X(net6707));
 sg13g2_dlygate4sd3_1 hold2321 (.A(\scanline[36][1] ),
    .X(net6708));
 sg13g2_dlygate4sd3_1 hold2322 (.A(\scanline[41][1] ),
    .X(net6709));
 sg13g2_dlygate4sd3_1 hold2323 (.A(\scanline[108][5] ),
    .X(net6710));
 sg13g2_dlygate4sd3_1 hold2324 (.A(\scanline[71][6] ),
    .X(net6711));
 sg13g2_dlygate4sd3_1 hold2325 (.A(\atari2600.ram[24][1] ),
    .X(net6712));
 sg13g2_dlygate4sd3_1 hold2326 (.A(\scanline[60][0] ),
    .X(net6713));
 sg13g2_dlygate4sd3_1 hold2327 (.A(\atari2600.ram[100][0] ),
    .X(net6714));
 sg13g2_dlygate4sd3_1 hold2328 (.A(\scanline[44][4] ),
    .X(net6715));
 sg13g2_dlygate4sd3_1 hold2329 (.A(\atari2600.ram[28][2] ),
    .X(net6716));
 sg13g2_dlygate4sd3_1 hold2330 (.A(\scanline[35][4] ),
    .X(net6717));
 sg13g2_dlygate4sd3_1 hold2331 (.A(\scanline[98][2] ),
    .X(net6718));
 sg13g2_dlygate4sd3_1 hold2332 (.A(\scanline[9][4] ),
    .X(net6719));
 sg13g2_dlygate4sd3_1 hold2333 (.A(\scanline[98][3] ),
    .X(net6720));
 sg13g2_dlygate4sd3_1 hold2334 (.A(\atari2600.ram[11][4] ),
    .X(net6721));
 sg13g2_dlygate4sd3_1 hold2335 (.A(\scanline[37][0] ),
    .X(net6722));
 sg13g2_dlygate4sd3_1 hold2336 (.A(\rom_last_read_addr[6] ),
    .X(net6723));
 sg13g2_dlygate4sd3_1 hold2337 (.A(_01132_),
    .X(net6724));
 sg13g2_dlygate4sd3_1 hold2338 (.A(\scanline[72][3] ),
    .X(net6725));
 sg13g2_dlygate4sd3_1 hold2339 (.A(\scanline[39][0] ),
    .X(net6726));
 sg13g2_dlygate4sd3_1 hold2340 (.A(\scanline[60][2] ),
    .X(net6727));
 sg13g2_dlygate4sd3_1 hold2341 (.A(\scanline[2][2] ),
    .X(net6728));
 sg13g2_dlygate4sd3_1 hold2342 (.A(\scanline[36][0] ),
    .X(net6729));
 sg13g2_dlygate4sd3_1 hold2343 (.A(\scanline[92][4] ),
    .X(net6730));
 sg13g2_dlygate4sd3_1 hold2344 (.A(\scanline[21][1] ),
    .X(net6731));
 sg13g2_dlygate4sd3_1 hold2345 (.A(\scanline[81][3] ),
    .X(net6732));
 sg13g2_dlygate4sd3_1 hold2346 (.A(\atari2600.cpu.D ),
    .X(net6733));
 sg13g2_dlygate4sd3_1 hold2347 (.A(_00014_),
    .X(net6734));
 sg13g2_dlygate4sd3_1 hold2348 (.A(\scanline[4][1] ),
    .X(net6735));
 sg13g2_dlygate4sd3_1 hold2349 (.A(\atari2600.ram[11][5] ),
    .X(net6736));
 sg13g2_dlygate4sd3_1 hold2350 (.A(\atari2600.ram[81][1] ),
    .X(net6737));
 sg13g2_dlygate4sd3_1 hold2351 (.A(\scanline[49][1] ),
    .X(net6738));
 sg13g2_dlygate4sd3_1 hold2352 (.A(\scanline[17][2] ),
    .X(net6739));
 sg13g2_dlygate4sd3_1 hold2353 (.A(\scanline[32][5] ),
    .X(net6740));
 sg13g2_dlygate4sd3_1 hold2354 (.A(\atari2600.ram[23][3] ),
    .X(net6741));
 sg13g2_dlygate4sd3_1 hold2355 (.A(\scanline[71][3] ),
    .X(net6742));
 sg13g2_dlygate4sd3_1 hold2356 (.A(\atari2600.ram[31][3] ),
    .X(net6743));
 sg13g2_dlygate4sd3_1 hold2357 (.A(\scanline[130][5] ),
    .X(net6744));
 sg13g2_dlygate4sd3_1 hold2358 (.A(\atari2600.ram[80][2] ),
    .X(net6745));
 sg13g2_dlygate4sd3_1 hold2359 (.A(\scanline[98][5] ),
    .X(net6746));
 sg13g2_dlygate4sd3_1 hold2360 (.A(\scanline[4][0] ),
    .X(net6747));
 sg13g2_dlygate4sd3_1 hold2361 (.A(\atari2600.tia.poly4_r.x[3] ),
    .X(net6748));
 sg13g2_dlygate4sd3_1 hold2362 (.A(_02244_),
    .X(net6749));
 sg13g2_dlygate4sd3_1 hold2363 (.A(\scanline[2][3] ),
    .X(net6750));
 sg13g2_dlygate4sd3_1 hold2364 (.A(\scanline[148][1] ),
    .X(net6751));
 sg13g2_dlygate4sd3_1 hold2365 (.A(\atari2600.ram[27][6] ),
    .X(net6752));
 sg13g2_dlygate4sd3_1 hold2366 (.A(\scanline[139][5] ),
    .X(net6753));
 sg13g2_dlygate4sd3_1 hold2367 (.A(\scanline[75][6] ),
    .X(net6754));
 sg13g2_dlygate4sd3_1 hold2368 (.A(\scanline[19][4] ),
    .X(net6755));
 sg13g2_dlygate4sd3_1 hold2369 (.A(_00051_),
    .X(net6756));
 sg13g2_dlygate4sd3_1 hold2370 (.A(_00042_),
    .X(net6757));
 sg13g2_dlygate4sd3_1 hold2371 (.A(\scanline[132][4] ),
    .X(net6758));
 sg13g2_dlygate4sd3_1 hold2372 (.A(\scanline[12][2] ),
    .X(net6759));
 sg13g2_dlygate4sd3_1 hold2373 (.A(\scanline[7][2] ),
    .X(net6760));
 sg13g2_dlygate4sd3_1 hold2374 (.A(\atari2600.ram[59][1] ),
    .X(net6761));
 sg13g2_dlygate4sd3_1 hold2375 (.A(\scanline[2][4] ),
    .X(net6762));
 sg13g2_dlygate4sd3_1 hold2376 (.A(\scanline[20][4] ),
    .X(net6763));
 sg13g2_dlygate4sd3_1 hold2377 (.A(\scanline[34][5] ),
    .X(net6764));
 sg13g2_dlygate4sd3_1 hold2378 (.A(\atari2600.ram[124][0] ),
    .X(net6765));
 sg13g2_dlygate4sd3_1 hold2379 (.A(\scanline[100][5] ),
    .X(net6766));
 sg13g2_dlygate4sd3_1 hold2380 (.A(\rom_last_read_addr[11] ),
    .X(net6767));
 sg13g2_dlygate4sd3_1 hold2381 (.A(_01137_),
    .X(net6768));
 sg13g2_dlygate4sd3_1 hold2382 (.A(\atari2600.ram[83][5] ),
    .X(net6769));
 sg13g2_dlygate4sd3_1 hold2383 (.A(\scanline[84][3] ),
    .X(net6770));
 sg13g2_dlygate4sd3_1 hold2384 (.A(\atari2600.ram[83][7] ),
    .X(net6771));
 sg13g2_dlygate4sd3_1 hold2385 (.A(\scanline[22][2] ),
    .X(net6772));
 sg13g2_dlygate4sd3_1 hold2386 (.A(\scanline[67][2] ),
    .X(net6773));
 sg13g2_dlygate4sd3_1 hold2387 (.A(\scanline[134][5] ),
    .X(net6774));
 sg13g2_dlygate4sd3_1 hold2388 (.A(\scanline[98][0] ),
    .X(net6775));
 sg13g2_dlygate4sd3_1 hold2389 (.A(\scanline[64][2] ),
    .X(net6776));
 sg13g2_dlygate4sd3_1 hold2390 (.A(\scanline[11][6] ),
    .X(net6777));
 sg13g2_dlygate4sd3_1 hold2391 (.A(\atari2600.ram[97][4] ),
    .X(net6778));
 sg13g2_dlygate4sd3_1 hold2392 (.A(\scanline[88][0] ),
    .X(net6779));
 sg13g2_dlygate4sd3_1 hold2393 (.A(\scanline[24][6] ),
    .X(net6780));
 sg13g2_dlygate4sd3_1 hold2394 (.A(\scanline[130][4] ),
    .X(net6781));
 sg13g2_dlygate4sd3_1 hold2395 (.A(\scanline[37][4] ),
    .X(net6782));
 sg13g2_dlygate4sd3_1 hold2396 (.A(\scanline[96][5] ),
    .X(net6783));
 sg13g2_dlygate4sd3_1 hold2397 (.A(\scanline[156][3] ),
    .X(net6784));
 sg13g2_dlygate4sd3_1 hold2398 (.A(\atari2600.cpu.AXYS[2][6] ),
    .X(net6785));
 sg13g2_dlygate4sd3_1 hold2399 (.A(\scanline[11][2] ),
    .X(net6786));
 sg13g2_dlygate4sd3_1 hold2400 (.A(\atari2600.cpu.dst_reg[1] ),
    .X(net6787));
 sg13g2_dlygate4sd3_1 hold2401 (.A(\scanline[49][3] ),
    .X(net6788));
 sg13g2_dlygate4sd3_1 hold2402 (.A(\scanline[97][4] ),
    .X(net6789));
 sg13g2_dlygate4sd3_1 hold2403 (.A(\scanline[56][4] ),
    .X(net6790));
 sg13g2_dlygate4sd3_1 hold2404 (.A(\atari2600.tia.audio_right_counter[8] ),
    .X(net6791));
 sg13g2_dlygate4sd3_1 hold2405 (.A(_02036_),
    .X(net6792));
 sg13g2_dlygate4sd3_1 hold2406 (.A(\scanline[41][4] ),
    .X(net6793));
 sg13g2_dlygate4sd3_1 hold2407 (.A(\scanline[138][3] ),
    .X(net6794));
 sg13g2_dlygate4sd3_1 hold2408 (.A(\atari2600.ram[52][7] ),
    .X(net6795));
 sg13g2_dlygate4sd3_1 hold2409 (.A(\scanline[112][5] ),
    .X(net6796));
 sg13g2_dlygate4sd3_1 hold2410 (.A(\scanline[131][4] ),
    .X(net6797));
 sg13g2_dlygate4sd3_1 hold2411 (.A(\scanline[18][6] ),
    .X(net6798));
 sg13g2_dlygate4sd3_1 hold2412 (.A(\scanline[11][5] ),
    .X(net6799));
 sg13g2_dlygate4sd3_1 hold2413 (.A(\scanline[138][2] ),
    .X(net6800));
 sg13g2_dlygate4sd3_1 hold2414 (.A(\scanline[134][1] ),
    .X(net6801));
 sg13g2_dlygate4sd3_1 hold2415 (.A(\scanline[92][0] ),
    .X(net6802));
 sg13g2_dlygate4sd3_1 hold2416 (.A(\scanline[129][0] ),
    .X(net6803));
 sg13g2_dlygate4sd3_1 hold2417 (.A(\atari2600.cpu.AXYS[1][2] ),
    .X(net6804));
 sg13g2_dlygate4sd3_1 hold2418 (.A(\scanline[135][0] ),
    .X(net6805));
 sg13g2_dlygate4sd3_1 hold2419 (.A(\scanline[72][4] ),
    .X(net6806));
 sg13g2_dlygate4sd3_1 hold2420 (.A(\atari2600.ram[39][5] ),
    .X(net6807));
 sg13g2_dlygate4sd3_1 hold2421 (.A(\scanline[139][0] ),
    .X(net6808));
 sg13g2_dlygate4sd3_1 hold2422 (.A(\scanline[40][3] ),
    .X(net6809));
 sg13g2_dlygate4sd3_1 hold2423 (.A(\scanline[19][5] ),
    .X(net6810));
 sg13g2_dlygate4sd3_1 hold2424 (.A(\scanline[11][1] ),
    .X(net6811));
 sg13g2_dlygate4sd3_1 hold2425 (.A(\scanline[43][1] ),
    .X(net6812));
 sg13g2_dlygate4sd3_1 hold2426 (.A(\scanline[65][3] ),
    .X(net6813));
 sg13g2_dlygate4sd3_1 hold2427 (.A(\atari2600.ram[111][4] ),
    .X(net6814));
 sg13g2_dlygate4sd3_1 hold2428 (.A(\scanline[33][4] ),
    .X(net6815));
 sg13g2_dlygate4sd3_1 hold2429 (.A(\atari2600.ram[127][6] ),
    .X(net6816));
 sg13g2_dlygate4sd3_1 hold2430 (.A(\atari2600.ram[47][3] ),
    .X(net6817));
 sg13g2_dlygate4sd3_1 hold2431 (.A(\atari2600.tia.poly9_l.x[7] ),
    .X(net6818));
 sg13g2_dlygate4sd3_1 hold2432 (.A(\scanline[33][6] ),
    .X(net6819));
 sg13g2_dlygate4sd3_1 hold2433 (.A(\atari2600.ram[11][1] ),
    .X(net6820));
 sg13g2_dlygate4sd3_1 hold2434 (.A(\scanline[9][0] ),
    .X(net6821));
 sg13g2_dlygate4sd3_1 hold2435 (.A(\atari2600.tia.diag[89] ),
    .X(net6822));
 sg13g2_dlygate4sd3_1 hold2436 (.A(\scanline[42][0] ),
    .X(net6823));
 sg13g2_dlygate4sd3_1 hold2437 (.A(\scanline[7][5] ),
    .X(net6824));
 sg13g2_dlygate4sd3_1 hold2438 (.A(\atari2600.ram[35][6] ),
    .X(net6825));
 sg13g2_dlygate4sd3_1 hold2439 (.A(\scanline[134][4] ),
    .X(net6826));
 sg13g2_dlygate4sd3_1 hold2440 (.A(\atari2600.ram[105][6] ),
    .X(net6827));
 sg13g2_dlygate4sd3_1 hold2441 (.A(\atari2600.ram[36][2] ),
    .X(net6828));
 sg13g2_dlygate4sd3_1 hold2442 (.A(\scanline[39][2] ),
    .X(net6829));
 sg13g2_dlygate4sd3_1 hold2443 (.A(\scanline[96][6] ),
    .X(net6830));
 sg13g2_dlygate4sd3_1 hold2444 (.A(\scanline[0][4] ),
    .X(net6831));
 sg13g2_dlygate4sd3_1 hold2445 (.A(\atari2600.tia.audio_right_counter[6] ),
    .X(net6832));
 sg13g2_dlygate4sd3_1 hold2446 (.A(\scanline[75][4] ),
    .X(net6833));
 sg13g2_dlygate4sd3_1 hold2447 (.A(\scanline[1][2] ),
    .X(net6834));
 sg13g2_dlygate4sd3_1 hold2448 (.A(\atari2600.ram[83][2] ),
    .X(net6835));
 sg13g2_dlygate4sd3_1 hold2449 (.A(\atari2600.ram[80][3] ),
    .X(net6836));
 sg13g2_dlygate4sd3_1 hold2450 (.A(\scanline[67][4] ),
    .X(net6837));
 sg13g2_dlygate4sd3_1 hold2451 (.A(\scanline[65][2] ),
    .X(net6838));
 sg13g2_dlygate4sd3_1 hold2452 (.A(\scanline[18][3] ),
    .X(net6839));
 sg13g2_dlygate4sd3_1 hold2453 (.A(\scanline[156][6] ),
    .X(net6840));
 sg13g2_dlygate4sd3_1 hold2454 (.A(\atari2600.cpu.rotate ),
    .X(net6841));
 sg13g2_dlygate4sd3_1 hold2455 (.A(\scanline[4][3] ),
    .X(net6842));
 sg13g2_dlygate4sd3_1 hold2456 (.A(\atari2600.cpu.AXYS[1][5] ),
    .X(net6843));
 sg13g2_dlygate4sd3_1 hold2457 (.A(\atari2600.ram[21][1] ),
    .X(net6844));
 sg13g2_dlygate4sd3_1 hold2458 (.A(\scanline[27][6] ),
    .X(net6845));
 sg13g2_dlygate4sd3_1 hold2459 (.A(\scanline[9][6] ),
    .X(net6846));
 sg13g2_dlygate4sd3_1 hold2460 (.A(\scanline[1][0] ),
    .X(net6847));
 sg13g2_dlygate4sd3_1 hold2461 (.A(\scanline[19][0] ),
    .X(net6848));
 sg13g2_dlygate4sd3_1 hold2462 (.A(\atari2600.cpu.AXYS[3][3] ),
    .X(net6849));
 sg13g2_dlygate4sd3_1 hold2463 (.A(\scanline[19][2] ),
    .X(net6850));
 sg13g2_dlygate4sd3_1 hold2464 (.A(\scanline[41][6] ),
    .X(net6851));
 sg13g2_dlygate4sd3_1 hold2465 (.A(\rom_last_read_addr[7] ),
    .X(net6852));
 sg13g2_dlygate4sd3_1 hold2466 (.A(_01133_),
    .X(net6853));
 sg13g2_dlygate4sd3_1 hold2467 (.A(\atari2600.tia.poly5_l.x[4] ),
    .X(net6854));
 sg13g2_dlygate4sd3_1 hold2468 (.A(_02231_),
    .X(net6855));
 sg13g2_dlygate4sd3_1 hold2469 (.A(\scanline[26][6] ),
    .X(net6856));
 sg13g2_dlygate4sd3_1 hold2470 (.A(\scanline[71][0] ),
    .X(net6857));
 sg13g2_dlygate4sd3_1 hold2471 (.A(\scanline[52][0] ),
    .X(net6858));
 sg13g2_dlygate4sd3_1 hold2472 (.A(\atari2600.ram[116][5] ),
    .X(net6859));
 sg13g2_dlygate4sd3_1 hold2473 (.A(\scanline[33][3] ),
    .X(net6860));
 sg13g2_dlygate4sd3_1 hold2474 (.A(\scanline[145][6] ),
    .X(net6861));
 sg13g2_dlygate4sd3_1 hold2475 (.A(\atari2600.ram[25][6] ),
    .X(net6862));
 sg13g2_dlygate4sd3_1 hold2476 (.A(\scanline[66][0] ),
    .X(net6863));
 sg13g2_dlygate4sd3_1 hold2477 (.A(\scanline[104][4] ),
    .X(net6864));
 sg13g2_dlygate4sd3_1 hold2478 (.A(\scanline[56][5] ),
    .X(net6865));
 sg13g2_dlygate4sd3_1 hold2479 (.A(\scanline[60][3] ),
    .X(net6866));
 sg13g2_dlygate4sd3_1 hold2480 (.A(\scanline[100][1] ),
    .X(net6867));
 sg13g2_dlygate4sd3_1 hold2481 (.A(\scanline[6][0] ),
    .X(net6868));
 sg13g2_dlygate4sd3_1 hold2482 (.A(\scanline[135][5] ),
    .X(net6869));
 sg13g2_dlygate4sd3_1 hold2483 (.A(\scanline[27][1] ),
    .X(net6870));
 sg13g2_dlygate4sd3_1 hold2484 (.A(\scanline[131][6] ),
    .X(net6871));
 sg13g2_dlygate4sd3_1 hold2485 (.A(\atari2600.tia.poly5_r.x[4] ),
    .X(net6872));
 sg13g2_dlygate4sd3_1 hold2486 (.A(\scanline[112][2] ),
    .X(net6873));
 sg13g2_dlygate4sd3_1 hold2487 (.A(\scanline[35][0] ),
    .X(net6874));
 sg13g2_dlygate4sd3_1 hold2488 (.A(\scanline[38][0] ),
    .X(net6875));
 sg13g2_dlygate4sd3_1 hold2489 (.A(\atari2600.pia.interval[10] ),
    .X(net6876));
 sg13g2_dlygate4sd3_1 hold2490 (.A(\atari2600.tia.poly4_r.x[1] ),
    .X(net6877));
 sg13g2_dlygate4sd3_1 hold2491 (.A(_02241_),
    .X(net6878));
 sg13g2_dlygate4sd3_1 hold2492 (.A(\scanline[140][6] ),
    .X(net6879));
 sg13g2_dlygate4sd3_1 hold2493 (.A(\scanline[22][1] ),
    .X(net6880));
 sg13g2_dlygate4sd3_1 hold2494 (.A(\atari2600.ram[25][0] ),
    .X(net6881));
 sg13g2_dlygate4sd3_1 hold2495 (.A(_00052_),
    .X(net6882));
 sg13g2_dlygate4sd3_1 hold2496 (.A(_00044_),
    .X(net6883));
 sg13g2_dlygate4sd3_1 hold2497 (.A(\scanline[44][3] ),
    .X(net6884));
 sg13g2_dlygate4sd3_1 hold2498 (.A(\atari2600.ram[99][7] ),
    .X(net6885));
 sg13g2_dlygate4sd3_1 hold2499 (.A(\scanline[104][0] ),
    .X(net6886));
 sg13g2_dlygate4sd3_1 hold2500 (.A(\scanline[27][5] ),
    .X(net6887));
 sg13g2_dlygate4sd3_1 hold2501 (.A(\scanline[3][2] ),
    .X(net6888));
 sg13g2_dlygate4sd3_1 hold2502 (.A(\atari2600.tia.audio_right_counter[2] ),
    .X(net6889));
 sg13g2_dlygate4sd3_1 hold2503 (.A(_02030_),
    .X(net6890));
 sg13g2_dlygate4sd3_1 hold2504 (.A(\atari2600.tia.p4_l ),
    .X(net6891));
 sg13g2_dlygate4sd3_1 hold2505 (.A(\scanline[136][6] ),
    .X(net6892));
 sg13g2_dlygate4sd3_1 hold2506 (.A(\scanline[48][6] ),
    .X(net6893));
 sg13g2_dlygate4sd3_1 hold2507 (.A(\scanline[146][4] ),
    .X(net6894));
 sg13g2_dlygate4sd3_1 hold2508 (.A(\scanline[146][0] ),
    .X(net6895));
 sg13g2_dlygate4sd3_1 hold2509 (.A(\scanline[5][6] ),
    .X(net6896));
 sg13g2_dlygate4sd3_1 hold2510 (.A(\scanline[35][5] ),
    .X(net6897));
 sg13g2_dlygate4sd3_1 hold2511 (.A(\scanline[82][6] ),
    .X(net6898));
 sg13g2_dlygate4sd3_1 hold2512 (.A(\scanline[48][0] ),
    .X(net6899));
 sg13g2_dlygate4sd3_1 hold2513 (.A(\scanline[84][0] ),
    .X(net6900));
 sg13g2_dlygate4sd3_1 hold2514 (.A(\atari2600.ram[115][0] ),
    .X(net6901));
 sg13g2_dlygate4sd3_1 hold2515 (.A(\scanline[88][5] ),
    .X(net6902));
 sg13g2_dlygate4sd3_1 hold2516 (.A(\atari2600.ram[103][4] ),
    .X(net6903));
 sg13g2_dlygate4sd3_1 hold2517 (.A(\scanline[3][1] ),
    .X(net6904));
 sg13g2_dlygate4sd3_1 hold2518 (.A(\atari2600.tia.colup0[0] ),
    .X(net6905));
 sg13g2_dlygate4sd3_1 hold2519 (.A(\atari2600.ram[36][5] ),
    .X(net6906));
 sg13g2_dlygate4sd3_1 hold2520 (.A(\scanline[134][3] ),
    .X(net6907));
 sg13g2_dlygate4sd3_1 hold2521 (.A(\scanline[1][5] ),
    .X(net6908));
 sg13g2_dlygate4sd3_1 hold2522 (.A(\scanline[21][4] ),
    .X(net6909));
 sg13g2_dlygate4sd3_1 hold2523 (.A(\scanline[137][5] ),
    .X(net6910));
 sg13g2_dlygate4sd3_1 hold2524 (.A(\scanline[96][4] ),
    .X(net6911));
 sg13g2_dlygate4sd3_1 hold2525 (.A(\scanline[112][1] ),
    .X(net6912));
 sg13g2_dlygate4sd3_1 hold2526 (.A(\scanline[4][4] ),
    .X(net6913));
 sg13g2_dlygate4sd3_1 hold2527 (.A(\scanline[52][5] ),
    .X(net6914));
 sg13g2_dlygate4sd3_1 hold2528 (.A(\scanline[140][5] ),
    .X(net6915));
 sg13g2_dlygate4sd3_1 hold2529 (.A(\scanline[80][2] ),
    .X(net6916));
 sg13g2_dlygate4sd3_1 hold2530 (.A(\atari2600.cpu.IRHOLD[2] ),
    .X(net6917));
 sg13g2_dlygate4sd3_1 hold2531 (.A(\atari2600.ram[9][5] ),
    .X(net6918));
 sg13g2_dlygate4sd3_1 hold2532 (.A(\atari2600.cpu.PC[12] ),
    .X(net6919));
 sg13g2_dlygate4sd3_1 hold2533 (.A(_02510_),
    .X(net6920));
 sg13g2_dlygate4sd3_1 hold2534 (.A(\scanline[56][3] ),
    .X(net6921));
 sg13g2_dlygate4sd3_1 hold2535 (.A(\atari2600.ram[103][2] ),
    .X(net6922));
 sg13g2_dlygate4sd3_1 hold2536 (.A(\scanline[25][4] ),
    .X(net6923));
 sg13g2_dlygate4sd3_1 hold2537 (.A(\scanline[3][6] ),
    .X(net6924));
 sg13g2_dlygate4sd3_1 hold2538 (.A(\scanline[27][4] ),
    .X(net6925));
 sg13g2_dlygate4sd3_1 hold2539 (.A(\scanline[128][3] ),
    .X(net6926));
 sg13g2_dlygate4sd3_1 hold2540 (.A(\scanline[7][6] ),
    .X(net6927));
 sg13g2_dlygate4sd3_1 hold2541 (.A(\atari2600.cpu.IRHOLD[3] ),
    .X(net6928));
 sg13g2_dlygate4sd3_1 hold2542 (.A(\scanline[50][4] ),
    .X(net6929));
 sg13g2_dlygate4sd3_1 hold2543 (.A(\scanline[76][6] ),
    .X(net6930));
 sg13g2_dlygate4sd3_1 hold2544 (.A(\atari2600.tia.vid_vsync ),
    .X(net6931));
 sg13g2_dlygate4sd3_1 hold2545 (.A(\scanline[23][6] ),
    .X(net6932));
 sg13g2_dlygate4sd3_1 hold2546 (.A(\rom_last_read_addr[2] ),
    .X(net6933));
 sg13g2_dlygate4sd3_1 hold2547 (.A(_01128_),
    .X(net6934));
 sg13g2_dlygate4sd3_1 hold2548 (.A(\atari2600.ram[21][7] ),
    .X(net6935));
 sg13g2_dlygate4sd3_1 hold2549 (.A(\scanline[11][4] ),
    .X(net6936));
 sg13g2_dlygate4sd3_1 hold2550 (.A(\atari2600.cpu.index_y ),
    .X(net6937));
 sg13g2_dlygate4sd3_1 hold2551 (.A(\scanline[10][2] ),
    .X(net6938));
 sg13g2_dlygate4sd3_1 hold2552 (.A(\atari2600.tia.poly9_r.x[4] ),
    .X(net6939));
 sg13g2_dlygate4sd3_1 hold2553 (.A(_02254_),
    .X(net6940));
 sg13g2_dlygate4sd3_1 hold2554 (.A(\atari2600.ram[37][2] ),
    .X(net6941));
 sg13g2_dlygate4sd3_1 hold2555 (.A(\atari2600.tia.diag[82] ),
    .X(net6942));
 sg13g2_dlygate4sd3_1 hold2556 (.A(\atari2600.tia.diag[97] ),
    .X(net6943));
 sg13g2_dlygate4sd3_1 hold2557 (.A(\scanline[148][5] ),
    .X(net6944));
 sg13g2_dlygate4sd3_1 hold2558 (.A(\atari2600.ram[17][7] ),
    .X(net6945));
 sg13g2_dlygate4sd3_1 hold2559 (.A(\atari2600.ram_data[3] ),
    .X(net6946));
 sg13g2_dlygate4sd3_1 hold2560 (.A(\scanline[44][1] ),
    .X(net6947));
 sg13g2_dlygate4sd3_1 hold2561 (.A(\atari2600.ram[8][3] ),
    .X(net6948));
 sg13g2_dlygate4sd3_1 hold2562 (.A(\scanline[139][2] ),
    .X(net6949));
 sg13g2_dlygate4sd3_1 hold2563 (.A(\scanline[49][2] ),
    .X(net6950));
 sg13g2_dlygate4sd3_1 hold2564 (.A(\atari2600.pia.diag[7] ),
    .X(net6951));
 sg13g2_dlygate4sd3_1 hold2565 (.A(_01762_),
    .X(net6952));
 sg13g2_dlygate4sd3_1 hold2566 (.A(\rom_last_read_addr[10] ),
    .X(net6953));
 sg13g2_dlygate4sd3_1 hold2567 (.A(_01136_),
    .X(net6954));
 sg13g2_dlygate4sd3_1 hold2568 (.A(\scanline[22][4] ),
    .X(net6955));
 sg13g2_dlygate4sd3_1 hold2569 (.A(\scanline[148][3] ),
    .X(net6956));
 sg13g2_dlygate4sd3_1 hold2570 (.A(\atari2600.tia.diag[93] ),
    .X(net6957));
 sg13g2_dlygate4sd3_1 hold2571 (.A(\atari2600.tia.colup0[6] ),
    .X(net6958));
 sg13g2_dlygate4sd3_1 hold2572 (.A(\scanline[156][2] ),
    .X(net6959));
 sg13g2_dlygate4sd3_1 hold2573 (.A(\atari2600.pia.time_counter[10] ),
    .X(net6960));
 sg13g2_dlygate4sd3_1 hold2574 (.A(_05321_),
    .X(net6961));
 sg13g2_dlygate4sd3_1 hold2575 (.A(\atari2600.cpu.cond_code[2] ),
    .X(net6962));
 sg13g2_dlygate4sd3_1 hold2576 (.A(\scanline[129][2] ),
    .X(net6963));
 sg13g2_dlygate4sd3_1 hold2577 (.A(\scanline[145][0] ),
    .X(net6964));
 sg13g2_dlygate4sd3_1 hold2578 (.A(\scanline[32][1] ),
    .X(net6965));
 sg13g2_dlygate4sd3_1 hold2579 (.A(\atari2600.ram[111][1] ),
    .X(net6966));
 sg13g2_dlygate4sd3_1 hold2580 (.A(\scanline[65][4] ),
    .X(net6967));
 sg13g2_dlygate4sd3_1 hold2581 (.A(\scanline[73][3] ),
    .X(net6968));
 sg13g2_dlygate4sd3_1 hold2582 (.A(\joypmod[2] ),
    .X(net6969));
 sg13g2_dlygate4sd3_1 hold2583 (.A(\atari2600.pia.time_counter[12] ),
    .X(net6970));
 sg13g2_dlygate4sd3_1 hold2584 (.A(\atari2600.cpu.IRHOLD[0] ),
    .X(net6971));
 sg13g2_dlygate4sd3_1 hold2585 (.A(_02457_),
    .X(net6972));
 sg13g2_dlygate4sd3_1 hold2586 (.A(\atari2600.cpu.inc ),
    .X(net6973));
 sg13g2_dlygate4sd3_1 hold2587 (.A(\scanline[6][3] ),
    .X(net6974));
 sg13g2_dlygate4sd3_1 hold2588 (.A(\atari2600.cpu.IRHOLD[4] ),
    .X(net6975));
 sg13g2_dlygate4sd3_1 hold2589 (.A(\atari2600.ram[47][2] ),
    .X(net6976));
 sg13g2_dlygate4sd3_1 hold2590 (.A(\scanline[135][3] ),
    .X(net6977));
 sg13g2_dlygate4sd3_1 hold2591 (.A(\atari2600.tia.colubk[2] ),
    .X(net6978));
 sg13g2_dlygate4sd3_1 hold2592 (.A(\atari2600.tia.audf0[0] ),
    .X(net6979));
 sg13g2_dlygate4sd3_1 hold2593 (.A(\atari2600.cpu.PC[2] ),
    .X(net6980));
 sg13g2_dlygate4sd3_1 hold2594 (.A(_02500_),
    .X(net6981));
 sg13g2_dlygate4sd3_1 hold2595 (.A(\atari2600.tia.colubk[3] ),
    .X(net6982));
 sg13g2_dlygate4sd3_1 hold2596 (.A(\rom_last_read_addr[1] ),
    .X(net6983));
 sg13g2_dlygate4sd3_1 hold2597 (.A(\rom_last_read_addr[8] ),
    .X(net6984));
 sg13g2_dlygate4sd3_1 hold2598 (.A(_01134_),
    .X(net6985));
 sg13g2_dlygate4sd3_1 hold2599 (.A(\atari2600.input_joystick_0[6] ),
    .X(net6986));
 sg13g2_dlygate4sd3_1 hold2600 (.A(\atari2600.tia.colubk[1] ),
    .X(net6987));
 sg13g2_dlygate4sd3_1 hold2601 (.A(\scanline[38][6] ),
    .X(net6988));
 sg13g2_dlygate4sd3_1 hold2602 (.A(\atari2600.pia.time_counter[2] ),
    .X(net6989));
 sg13g2_dlygate4sd3_1 hold2603 (.A(_05300_),
    .X(net6990));
 sg13g2_dlygate4sd3_1 hold2604 (.A(_01774_),
    .X(net6991));
 sg13g2_dlygate4sd3_1 hold2605 (.A(\atari2600.cpu.bit_ins ),
    .X(net6992));
 sg13g2_dlygate4sd3_1 hold2606 (.A(\atari2600.pia.time_counter[13] ),
    .X(net6993));
 sg13g2_dlygate4sd3_1 hold2607 (.A(_05328_),
    .X(net6994));
 sg13g2_dlygate4sd3_1 hold2608 (.A(\scanline[136][5] ),
    .X(net6995));
 sg13g2_dlygate4sd3_1 hold2609 (.A(\atari2600.cpu.adc_sbc ),
    .X(net6996));
 sg13g2_dlygate4sd3_1 hold2610 (.A(\atari2600.input_switches[0] ),
    .X(net6997));
 sg13g2_dlygate4sd3_1 hold2611 (.A(\atari2600.tia.audio_right_counter[12] ),
    .X(net6998));
 sg13g2_dlygate4sd3_1 hold2612 (.A(\atari2600.cpu.PC[10] ),
    .X(net6999));
 sg13g2_dlygate4sd3_1 hold2613 (.A(_02508_),
    .X(net7000));
 sg13g2_dlygate4sd3_1 hold2614 (.A(\atari2600.tia.poly4_r.x[2] ),
    .X(net7001));
 sg13g2_dlygate4sd3_1 hold2615 (.A(\atari2600.cpu.cond_code[0] ),
    .X(net7002));
 sg13g2_dlygate4sd3_1 hold2616 (.A(\atari2600.cpu.load_only ),
    .X(net7003));
 sg13g2_dlygate4sd3_1 hold2617 (.A(\atari2600.cpu.clv ),
    .X(net7004));
 sg13g2_dlygate4sd3_1 hold2618 (.A(\atari2600.tia.colup1[6] ),
    .X(net7005));
 sg13g2_dlygate4sd3_1 hold2619 (.A(\atari2600.tia.p9_l ),
    .X(net7006));
 sg13g2_dlygate4sd3_1 hold2620 (.A(\atari2600.tia.diag[81] ),
    .X(net7007));
 sg13g2_dlygate4sd3_1 hold2621 (.A(\atari2600.cpu.ABL[1] ),
    .X(net7008));
 sg13g2_dlygate4sd3_1 hold2622 (.A(\atari2600.pia.interval[3] ),
    .X(net7009));
 sg13g2_dlygate4sd3_1 hold2623 (.A(\atari2600.tia.diag[83] ),
    .X(net7010));
 sg13g2_dlygate4sd3_1 hold2624 (.A(\atari2600.cpu.ABH[4] ),
    .X(net7011));
 sg13g2_dlygate4sd3_1 hold2625 (.A(\atari2600.tia.audio_l ),
    .X(net7012));
 sg13g2_dlygate4sd3_1 hold2626 (.A(_01150_),
    .X(net7013));
 sg13g2_dlygate4sd3_1 hold2627 (.A(\atari2600.tia.colubk[4] ),
    .X(net7014));
 sg13g2_dlygate4sd3_1 hold2628 (.A(\atari2600.tia.diag[94] ),
    .X(net7015));
 sg13g2_dlygate4sd3_1 hold2629 (.A(\atari2600.tia.poly5_r.x[3] ),
    .X(net7016));
 sg13g2_dlygate4sd3_1 hold2630 (.A(\atari2600.tia.poly4_l.x[3] ),
    .X(net7017));
 sg13g2_dlygate4sd3_1 hold2631 (.A(_00105_),
    .X(net7018));
 sg13g2_dlygate4sd3_1 hold2632 (.A(_01138_),
    .X(net7019));
 sg13g2_dlygate4sd3_1 hold2633 (.A(\atari2600.input_joystick_0[3] ),
    .X(net7020));
 sg13g2_dlygate4sd3_1 hold2634 (.A(\atari2600.tia.audio_left_counter[1] ),
    .X(net7021));
 sg13g2_dlygate4sd3_1 hold2635 (.A(_02013_),
    .X(net7022));
 sg13g2_dlygate4sd3_1 hold2636 (.A(\atari2600.input_joystick_0[4] ),
    .X(net7023));
 sg13g2_dlygate4sd3_1 hold2637 (.A(\atari2600.tia.colup1[2] ),
    .X(net7024));
 sg13g2_dlygate4sd3_1 hold2638 (.A(\atari2600.tia.diag[91] ),
    .X(net7025));
 sg13g2_dlygate4sd3_1 hold2639 (.A(\atari2600.pia.diag[0] ),
    .X(net7026));
 sg13g2_dlygate4sd3_1 hold2640 (.A(\flash_rom.stall_read ),
    .X(net7027));
 sg13g2_dlygate4sd3_1 hold2641 (.A(_03221_),
    .X(net7028));
 sg13g2_dlygate4sd3_1 hold2642 (.A(\scanline[56][6] ),
    .X(net7029));
 sg13g2_dlygate4sd3_1 hold2643 (.A(\atari2600.tia.diag[90] ),
    .X(net7030));
 sg13g2_dlygate4sd3_1 hold2644 (.A(\atari2600.ram_data[6] ),
    .X(net7031));
 sg13g2_dlygate4sd3_1 hold2645 (.A(\atari2600.cpu.IRHOLD[1] ),
    .X(net7032));
 sg13g2_dlygate4sd3_1 hold2646 (.A(_02458_),
    .X(net7033));
 sg13g2_dlygate4sd3_1 hold2647 (.A(\atari2600.pia.reset_timer[7] ),
    .X(net7034));
 sg13g2_dlygate4sd3_1 hold2648 (.A(_00143_),
    .X(net7035));
 sg13g2_dlygate4sd3_1 hold2649 (.A(\atari2600.tia.colup0[5] ),
    .X(net7036));
 sg13g2_dlygate4sd3_1 hold2650 (.A(\atari2600.cpu.ABH[6] ),
    .X(net7037));
 sg13g2_dlygate4sd3_1 hold2651 (.A(_02983_),
    .X(net7038));
 sg13g2_dlygate4sd3_1 hold2652 (.A(\hvsync_gen.vga.vpos[7] ),
    .X(net7039));
 sg13g2_dlygate4sd3_1 hold2653 (.A(_07634_),
    .X(net7040));
 sg13g2_dlygate4sd3_1 hold2654 (.A(\atari2600.tia.audf1[4] ),
    .X(net7041));
 sg13g2_dlygate4sd3_1 hold2655 (.A(\atari2600.cpu.ALU.HC ),
    .X(net7042));
 sg13g2_dlygate4sd3_1 hold2656 (.A(\atari2600.tia.colubk[6] ),
    .X(net7043));
 sg13g2_dlygate4sd3_1 hold2657 (.A(\atari2600.input_switches[2] ),
    .X(net7044));
 sg13g2_dlygate4sd3_1 hold2658 (.A(\atari2600.rom_data[2] ),
    .X(net7045));
 sg13g2_dlygate4sd3_1 hold2659 (.A(\atari2600.tia.diag[88] ),
    .X(net7046));
 sg13g2_dlygate4sd3_1 hold2660 (.A(\atari2600.tia.diag[95] ),
    .X(net7047));
 sg13g2_dlygate4sd3_1 hold2661 (.A(\atari2600.tia.diag[92] ),
    .X(net7048));
 sg13g2_dlygate4sd3_1 hold2662 (.A(\atari2600.tia.diag[76] ),
    .X(net7049));
 sg13g2_dlygate4sd3_1 hold2663 (.A(\atari2600.tia.diag[87] ),
    .X(net7050));
 sg13g2_dlygate4sd3_1 hold2664 (.A(\scanline[1][6] ),
    .X(net7051));
 sg13g2_dlygate4sd3_1 hold2665 (.A(\atari2600.cpu.PC[14] ),
    .X(net7052));
 sg13g2_dlygate4sd3_1 hold2666 (.A(\rom_last_read_addr[9] ),
    .X(net7053));
 sg13g2_dlygate4sd3_1 hold2667 (.A(_01135_),
    .X(net7054));
 sg13g2_dlygate4sd3_1 hold2668 (.A(\atari2600.cpu.PC[1] ),
    .X(net7055));
 sg13g2_dlygate4sd3_1 hold2669 (.A(_02499_),
    .X(net7056));
 sg13g2_dlygate4sd3_1 hold2670 (.A(\atari2600.rom_data[0] ),
    .X(net7057));
 sg13g2_dlygate4sd3_1 hold2671 (.A(\atari2600.tia.colup1[0] ),
    .X(net7058));
 sg13g2_dlygate4sd3_1 hold2672 (.A(\atari2600.tia.colubk[0] ),
    .X(net7059));
 sg13g2_dlygate4sd3_1 hold2673 (.A(\atari2600.pia.diag[6] ),
    .X(net7060));
 sg13g2_dlygate4sd3_1 hold2674 (.A(_01761_),
    .X(net7061));
 sg13g2_dlygate4sd3_1 hold2675 (.A(\atari2600.pia.time_counter[16] ),
    .X(net7062));
 sg13g2_dlygate4sd3_1 hold2676 (.A(_05334_),
    .X(net7063));
 sg13g2_dlygate4sd3_1 hold2677 (.A(\atari2600.cpu.PC[8] ),
    .X(net7064));
 sg13g2_dlygate4sd3_1 hold2678 (.A(\atari2600.ram_data[1] ),
    .X(net7065));
 sg13g2_dlygate4sd3_1 hold2679 (.A(_00153_),
    .X(net7066));
 sg13g2_dlygate4sd3_1 hold2680 (.A(\atari2600.tia.diag[86] ),
    .X(net7067));
 sg13g2_dlygate4sd3_1 hold2681 (.A(\atari2600.cpu.PC[7] ),
    .X(net7068));
 sg13g2_dlygate4sd3_1 hold2682 (.A(_02505_),
    .X(net7069));
 sg13g2_dlygate4sd3_1 hold2683 (.A(\atari2600.tia.diag[80] ),
    .X(net7070));
 sg13g2_dlygate4sd3_1 hold2684 (.A(\atari2600.pia.time_counter[3] ),
    .X(net7071));
 sg13g2_dlygate4sd3_1 hold2685 (.A(_05302_),
    .X(net7072));
 sg13g2_dlygate4sd3_1 hold2686 (.A(_01775_),
    .X(net7073));
 sg13g2_dlygate4sd3_1 hold2687 (.A(\atari2600.pia.diag[3] ),
    .X(net7074));
 sg13g2_dlygate4sd3_1 hold2688 (.A(\atari2600.pia.diag[5] ),
    .X(net7075));
 sg13g2_dlygate4sd3_1 hold2689 (.A(\atari2600.tia.colubk[5] ),
    .X(net7076));
 sg13g2_dlygate4sd3_1 hold2690 (.A(\atari2600.ram[44][2] ),
    .X(net7077));
 sg13g2_dlygate4sd3_1 hold2691 (.A(\atari2600.cpu.ABH[0] ),
    .X(net7078));
 sg13g2_dlygate4sd3_1 hold2692 (.A(\atari2600.cpu.PC[6] ),
    .X(net7079));
 sg13g2_dlygate4sd3_1 hold2693 (.A(_02504_),
    .X(net7080));
 sg13g2_dlygate4sd3_1 hold2694 (.A(uio_oe[1]),
    .X(net7081));
 sg13g2_dlygate4sd3_1 hold2695 (.A(\atari2600.pia.interval[6] ),
    .X(net7082));
 sg13g2_dlygate4sd3_1 hold2696 (.A(\atari2600.cpu.PC[15] ),
    .X(net7083));
 sg13g2_dlygate4sd3_1 hold2697 (.A(_02513_),
    .X(net7084));
 sg13g2_dlygate4sd3_1 hold2698 (.A(\atari2600.cpu.ABH[3] ),
    .X(net7085));
 sg13g2_dlygate4sd3_1 hold2699 (.A(\rom_next_addr_in_queue[5] ),
    .X(net7086));
 sg13g2_dlygate4sd3_1 hold2700 (.A(\atari2600.pia.diag[1] ),
    .X(net7087));
 sg13g2_dlygate4sd3_1 hold2701 (.A(_01756_),
    .X(net7088));
 sg13g2_dlygate4sd3_1 hold2702 (.A(\atari2600.cpu.PC[11] ),
    .X(net7089));
 sg13g2_dlygate4sd3_1 hold2703 (.A(_02509_),
    .X(net7090));
 sg13g2_dlygate4sd3_1 hold2704 (.A(\atari2600.input_joystick_0[0] ),
    .X(net7091));
 sg13g2_dlygate4sd3_1 hold2705 (.A(\atari2600.tia.colupf[1] ),
    .X(net7092));
 sg13g2_dlygate4sd3_1 hold2706 (.A(\atari2600.tia.diag[104] ),
    .X(net7093));
 sg13g2_dlygate4sd3_1 hold2707 (.A(\atari2600.input_switches[1] ),
    .X(net7094));
 sg13g2_dlygate4sd3_1 hold2708 (.A(\atari2600.pia.time_counter[21] ),
    .X(net7095));
 sg13g2_dlygate4sd3_1 hold2709 (.A(\atari2600.pia.reset_timer[2] ),
    .X(net7096));
 sg13g2_dlygate4sd3_1 hold2710 (.A(\atari2600.tia.colupf[3] ),
    .X(net7097));
 sg13g2_dlygate4sd3_1 hold2711 (.A(\atari2600.tia.diag[108] ),
    .X(net7098));
 sg13g2_dlygate4sd3_1 hold2712 (.A(\atari2600.tia.diag[84] ),
    .X(net7099));
 sg13g2_dlygate4sd3_1 hold2713 (.A(\atari2600.cpu.ABH[2] ),
    .X(net7100));
 sg13g2_dlygate4sd3_1 hold2714 (.A(\atari2600.input_joystick_0[3] ),
    .X(net7101));
 sg13g2_dlygate4sd3_1 hold2715 (.A(\atari2600.input_joystick_0[5] ),
    .X(net7102));
 sg13g2_dlygate4sd3_1 hold2716 (.A(\atari2600.cpu.shift_right ),
    .X(net7103));
 sg13g2_dlygate4sd3_1 hold2717 (.A(\atari2600.tia.p1_spacing[6] ),
    .X(net7104));
 sg13g2_dlygate4sd3_1 hold2718 (.A(\rom_next_addr_in_queue[4] ),
    .X(net7105));
 sg13g2_dlygate4sd3_1 hold2719 (.A(\atari2600.tia.diag[101] ),
    .X(net7106));
 sg13g2_dlygate4sd3_1 hold2720 (.A(\atari2600.cpu.ABH[1] ),
    .X(net7107));
 sg13g2_dlygate4sd3_1 hold2721 (.A(\atari2600.tia.diag[111] ),
    .X(net7108));
 sg13g2_dlygate4sd3_1 hold2722 (.A(\atari2600.pia.time_counter[15] ),
    .X(net7109));
 sg13g2_dlygate4sd3_1 hold2723 (.A(\flash_rom.addr[4] ),
    .X(net7110));
 sg13g2_dlygate4sd3_1 hold2724 (.A(_10468_),
    .X(net7111));
 sg13g2_dlygate4sd3_1 hold2725 (.A(_00201_),
    .X(net7112));
 sg13g2_dlygate4sd3_1 hold2726 (.A(\atari2600.cpu.cond_code[1] ),
    .X(net7113));
 sg13g2_dlygate4sd3_1 hold2727 (.A(\atari2600.tia.hmm0[2] ),
    .X(net7114));
 sg13g2_dlygate4sd3_1 hold2728 (.A(\atari2600.pia.diag[2] ),
    .X(net7115));
 sg13g2_dlygate4sd3_1 hold2729 (.A(\atari2600.tia.colupf[0] ),
    .X(net7116));
 sg13g2_dlygate4sd3_1 hold2730 (.A(\atari2600.pia.time_counter[0] ),
    .X(net7117));
 sg13g2_dlygate4sd3_1 hold2731 (.A(\atari2600.tia.hmm0[3] ),
    .X(net7118));
 sg13g2_dlygate4sd3_1 hold2732 (.A(\rom_next_addr_in_queue[6] ),
    .X(net7119));
 sg13g2_dlygate4sd3_1 hold2733 (.A(\rom_next_addr_in_queue[10] ),
    .X(net7120));
 sg13g2_dlygate4sd3_1 hold2734 (.A(\atari2600.pia.time_counter[22] ),
    .X(net7121));
 sg13g2_dlygate4sd3_1 hold2735 (.A(\atari2600.clk_counter[0] ),
    .X(net7122));
 sg13g2_dlygate4sd3_1 hold2736 (.A(\atari2600.cpu.PC[0] ),
    .X(net7123));
 sg13g2_dlygate4sd3_1 hold2737 (.A(_02498_),
    .X(net7124));
 sg13g2_dlygate4sd3_1 hold2738 (.A(\atari2600.tia.hmp1[2] ),
    .X(net7125));
 sg13g2_dlygate4sd3_1 hold2739 (.A(\atari2600.tia.hmm0[0] ),
    .X(net7126));
 sg13g2_dlygate4sd3_1 hold2740 (.A(\atari2600.tia.m1_w[1] ),
    .X(net7127));
 sg13g2_dlygate4sd3_1 hold2741 (.A(\rom_next_addr_in_queue[7] ),
    .X(net7128));
 sg13g2_dlygate4sd3_1 hold2742 (.A(\atari2600.tia.m1_w[0] ),
    .X(net7129));
 sg13g2_dlygate4sd3_1 hold2743 (.A(\atari2600.tia.m0_w[2] ),
    .X(net7130));
 sg13g2_dlygate4sd3_1 hold2744 (.A(\atari2600.tia.diag[109] ),
    .X(net7131));
 sg13g2_dlygate4sd3_1 hold2745 (.A(\atari2600.cpu.PC[5] ),
    .X(net7132));
 sg13g2_dlygate4sd3_1 hold2746 (.A(_02503_),
    .X(net7133));
 sg13g2_dlygate4sd3_1 hold2747 (.A(\atari2600.tia.hmm0[1] ),
    .X(net7134));
 sg13g2_dlygate4sd3_1 hold2748 (.A(\atari2600.tia.colup1[5] ),
    .X(net7135));
 sg13g2_dlygate4sd3_1 hold2749 (.A(\rom_next_addr_in_queue[3] ),
    .X(net7136));
 sg13g2_dlygate4sd3_1 hold2750 (.A(\atari2600.cpu.php ),
    .X(net7137));
 sg13g2_dlygate4sd3_1 hold2751 (.A(\hvsync_gen.vga.vpos[1] ),
    .X(net7138));
 sg13g2_dlygate4sd3_1 hold2752 (.A(\atari2600.cpu.adc_bcd ),
    .X(net7139));
 sg13g2_dlygate4sd3_1 hold2753 (.A(\flash_rom.addr[7] ),
    .X(net7140));
 sg13g2_dlygate4sd3_1 hold2754 (.A(_00200_),
    .X(net7141));
 sg13g2_dlygate4sd3_1 hold2755 (.A(\hvsync_gen.vga.vpos[9] ),
    .X(net7142));
 sg13g2_dlygate4sd3_1 hold2756 (.A(_02595_),
    .X(net7143));
 sg13g2_dlygate4sd3_1 hold2757 (.A(\atari2600.tia.hmp1[1] ),
    .X(net7144));
 sg13g2_dlygate4sd3_1 hold2758 (.A(\atari2600.tia.p0_w[5] ),
    .X(net7145));
 sg13g2_dlygate4sd3_1 hold2759 (.A(\atari2600.cpu.shift ),
    .X(net7146));
 sg13g2_dlygate4sd3_1 hold2760 (.A(\hvsync_gen.vga.vpos[4] ),
    .X(net7147));
 sg13g2_dlygate4sd3_1 hold2761 (.A(_07627_),
    .X(net7148));
 sg13g2_dlygate4sd3_1 hold2762 (.A(\atari2600.tia.m0_w[1] ),
    .X(net7149));
 sg13g2_dlygate4sd3_1 hold2763 (.A(\atari2600.tia.hmp1[0] ),
    .X(net7150));
 sg13g2_dlygate4sd3_1 hold2764 (.A(\rom_next_addr_in_queue[8] ),
    .X(net7151));
 sg13g2_dlygate4sd3_1 hold2765 (.A(\atari2600.tia.m0_w[0] ),
    .X(net7152));
 sg13g2_dlygate4sd3_1 hold2766 (.A(\flash_rom.addr[20] ),
    .X(net7153));
 sg13g2_dlygate4sd3_1 hold2767 (.A(\atari2600.tia.p0_w[4] ),
    .X(net7154));
 sg13g2_dlygate4sd3_1 hold2768 (.A(\atari2600.cpu.PC[3] ),
    .X(net7155));
 sg13g2_dlygate4sd3_1 hold2769 (.A(_02501_),
    .X(net7156));
 sg13g2_dlygate4sd3_1 hold2770 (.A(\atari2600.tia.colupf[4] ),
    .X(net7157));
 sg13g2_dlygate4sd3_1 hold2771 (.A(\atari2600.tia.colup1[4] ),
    .X(net7158));
 sg13g2_dlygate4sd3_1 hold2772 (.A(\atari2600.pia.time_counter[7] ),
    .X(net7159));
 sg13g2_dlygate4sd3_1 hold2773 (.A(\atari2600.tia.hmp0[2] ),
    .X(net7160));
 sg13g2_dlygate4sd3_1 hold2774 (.A(\atari2600.tia.hmm1[0] ),
    .X(net7161));
 sg13g2_dlygate4sd3_1 hold2775 (.A(\atari2600.tia.hmp0[0] ),
    .X(net7162));
 sg13g2_dlygate4sd3_1 hold2776 (.A(\hvsync_gen.vga.vpos[2] ),
    .X(net7163));
 sg13g2_dlygate4sd3_1 hold2777 (.A(\atari2600.tia.colupf[2] ),
    .X(net7164));
 sg13g2_dlygate4sd3_1 hold2778 (.A(\atari2600.tia.hmm1[2] ),
    .X(net7165));
 sg13g2_dlygate4sd3_1 hold2779 (.A(\atari2600.tia.diag[55] ),
    .X(net7166));
 sg13g2_dlygate4sd3_1 hold2780 (.A(\atari2600.tia.p5_r ),
    .X(net7167));
 sg13g2_dlygate4sd3_1 hold2781 (.A(_02245_),
    .X(net7168));
 sg13g2_dlygate4sd3_1 hold2782 (.A(\atari2600.tia.enam0 ),
    .X(net7169));
 sg13g2_dlygate4sd3_1 hold2783 (.A(\atari2600.tia.m1_w[3] ),
    .X(net7170));
 sg13g2_dlygate4sd3_1 hold2784 (.A(\atari2600.tia.diag[106] ),
    .X(net7171));
 sg13g2_dlygate4sd3_1 hold2785 (.A(\atari2600.pia.time_counter[4] ),
    .X(net7172));
 sg13g2_dlygate4sd3_1 hold2786 (.A(_05306_),
    .X(net7173));
 sg13g2_dlygate4sd3_1 hold2787 (.A(\flash_rom.nibbles_remaining[0] ),
    .X(net7174));
 sg13g2_dlygate4sd3_1 hold2788 (.A(\flash_rom.addr[6] ),
    .X(net7175));
 sg13g2_dlygate4sd3_1 hold2789 (.A(\hvsync_gen.vga.vpos[8] ),
    .X(net7176));
 sg13g2_dlygate4sd3_1 hold2790 (.A(\atari2600.tia.m1_w[2] ),
    .X(net7177));
 sg13g2_dlygate4sd3_1 hold2791 (.A(\atari2600.tia.p1_spacing[4] ),
    .X(net7178));
 sg13g2_dlygate4sd3_1 hold2792 (.A(\hvsync_gen.hpos[1] ),
    .X(net7179));
 sg13g2_dlygate4sd3_1 hold2793 (.A(_03223_),
    .X(net7180));
 sg13g2_dlygate4sd3_1 hold2794 (.A(_01349_),
    .X(net7181));
 sg13g2_dlygate4sd3_1 hold2795 (.A(\atari2600.tia.hmm1[1] ),
    .X(net7182));
 sg13g2_dlygate4sd3_1 hold2796 (.A(\atari2600.tia.diag[107] ),
    .X(net7183));
 sg13g2_dlygate4sd3_1 hold2797 (.A(\atari2600.tia.p1_w[5] ),
    .X(net7184));
 sg13g2_dlygate4sd3_1 hold2798 (.A(\atari2600.address_bus_r[11] ),
    .X(net7185));
 sg13g2_dlygate4sd3_1 hold2799 (.A(\atari2600.tia.colup1[3] ),
    .X(net7186));
 sg13g2_dlygate4sd3_1 hold2800 (.A(\hvsync_gen.vga.vpos[5] ),
    .X(net7187));
 sg13g2_dlygate4sd3_1 hold2801 (.A(_07631_),
    .X(net7188));
 sg13g2_dlygate4sd3_1 hold2802 (.A(\atari2600.cpu.PC[4] ),
    .X(net7189));
 sg13g2_dlygate4sd3_1 hold2803 (.A(\atari2600.tia.colupf[6] ),
    .X(net7190));
 sg13g2_dlygate4sd3_1 hold2804 (.A(\atari2600.tia.hmp0[1] ),
    .X(net7191));
 sg13g2_dlygate4sd3_1 hold2805 (.A(\atari2600.tia.colup0[3] ),
    .X(net7192));
 sg13g2_dlygate4sd3_1 hold2806 (.A(_00137_),
    .X(net7193));
 sg13g2_dlygate4sd3_1 hold2807 (.A(_07820_),
    .X(net7194));
 sg13g2_dlygate4sd3_1 hold2808 (.A(\atari2600.address_bus_r[10] ),
    .X(net7195));
 sg13g2_dlygate4sd3_1 hold2809 (.A(\atari2600.tia.p0_spacing[4] ),
    .X(net7196));
 sg13g2_dlygate4sd3_1 hold2810 (.A(\atari2600.cpu.op[1] ),
    .X(net7197));
 sg13g2_dlygate4sd3_1 hold2811 (.A(\atari2600.tia.p1_w[4] ),
    .X(net7198));
 sg13g2_dlygate4sd3_1 hold2812 (.A(\flash_rom.nibbles_remaining[2] ),
    .X(net7199));
 sg13g2_dlygate4sd3_1 hold2813 (.A(_07804_),
    .X(net7200));
 sg13g2_dlygate4sd3_1 hold2814 (.A(\atari2600.tia.hmbl[0] ),
    .X(net7201));
 sg13g2_dlygate4sd3_1 hold2815 (.A(\atari2600.cpu.DI[7] ),
    .X(net7202));
 sg13g2_dlygate4sd3_1 hold2816 (.A(_02478_),
    .X(net7203));
 sg13g2_dlygate4sd3_1 hold2817 (.A(\atari2600.cpu.op[0] ),
    .X(net7204));
 sg13g2_dlygate4sd3_1 hold2818 (.A(\atari2600.tia.colup1[1] ),
    .X(net7205));
 sg13g2_dlygate4sd3_1 hold2819 (.A(\flash_rom.nibbles_remaining[1] ),
    .X(net7206));
 sg13g2_dlygate4sd3_1 hold2820 (.A(\atari2600.tia.m0_w[3] ),
    .X(net7207));
 sg13g2_dlygate4sd3_1 hold2821 (.A(\atari2600.pia.time_counter[1] ),
    .X(net7208));
 sg13g2_dlygate4sd3_1 hold2822 (.A(\rom_next_addr_in_queue[1] ),
    .X(net7209));
 sg13g2_dlygate4sd3_1 hold2823 (.A(_03267_),
    .X(net7210));
 sg13g2_dlygate4sd3_1 hold2824 (.A(_03268_),
    .X(net7211));
 sg13g2_dlygate4sd3_1 hold2825 (.A(\atari2600.tia.hmp1[3] ),
    .X(net7212));
 sg13g2_dlygate4sd3_1 hold2826 (.A(\rom_last_read_addr[0] ),
    .X(net7213));
 sg13g2_dlygate4sd3_1 hold2827 (.A(_03240_),
    .X(net7214));
 sg13g2_dlygate4sd3_1 hold2828 (.A(uio_oe[5]),
    .X(net7215));
 sg13g2_dlygate4sd3_1 hold2829 (.A(_02930_),
    .X(net7216));
 sg13g2_dlygate4sd3_1 hold2830 (.A(\atari2600.tia.colup0[4] ),
    .X(net7217));
 sg13g2_dlygate4sd3_1 hold2831 (.A(\hvsync_gen.vga.vpos[6] ),
    .X(net7218));
 sg13g2_dlygate4sd3_1 hold2832 (.A(\atari2600.tia.hmbl[1] ),
    .X(net7219));
 sg13g2_dlygate4sd3_1 hold2833 (.A(\flash_rom.addr[5] ),
    .X(net7220));
 sg13g2_dlygate4sd3_1 hold2834 (.A(\atari2600.cpu.compare ),
    .X(net7221));
 sg13g2_dlygate4sd3_1 hold2835 (.A(\atari2600.tia.diag[36] ),
    .X(net7222));
 sg13g2_dlygate4sd3_1 hold2836 (.A(\rom_next_addr_in_queue[11] ),
    .X(net7223));
 sg13g2_dlygate4sd3_1 hold2837 (.A(\atari2600.ram_data[7] ),
    .X(net7224));
 sg13g2_dlygate4sd3_1 hold2838 (.A(\atari2600.cpu.store ),
    .X(net7225));
 sg13g2_dlygate4sd3_1 hold2839 (.A(\atari2600.address_bus_r[4] ),
    .X(net7226));
 sg13g2_dlygate4sd3_1 hold2840 (.A(\atari2600.tia.ball_w[1] ),
    .X(net7227));
 sg13g2_dlygate4sd3_1 hold2841 (.A(\atari2600.cpu.res ),
    .X(net7228));
 sg13g2_dlygate4sd3_1 hold2842 (.A(\flash_rom.spi_clk_out ),
    .X(net7229));
 sg13g2_dlygate4sd3_1 hold2843 (.A(_07643_),
    .X(net7230));
 sg13g2_dlygate4sd3_1 hold2844 (.A(_02596_),
    .X(net7231));
 sg13g2_dlygate4sd3_1 hold2845 (.A(\atari2600.tia.enam1 ),
    .X(net7232));
 sg13g2_dlygate4sd3_1 hold2846 (.A(\atari2600.tia.colupf[5] ),
    .X(net7233));
 sg13g2_dlygate4sd3_1 hold2847 (.A(_00138_),
    .X(net7234));
 sg13g2_dlygate4sd3_1 hold2848 (.A(\atari2600.tia.diag[46] ),
    .X(net7235));
 sg13g2_dlygate4sd3_1 hold2849 (.A(\hvsync_gen.vga.vpos[3] ),
    .X(net7236));
 sg13g2_dlygate4sd3_1 hold2850 (.A(\atari2600.pia.time_counter[23] ),
    .X(net7237));
 sg13g2_dlygate4sd3_1 hold2851 (.A(\atari2600.tia.ball_w[0] ),
    .X(net7238));
 sg13g2_dlygate4sd3_1 hold2852 (.A(\atari2600.tia.enabl ),
    .X(net7239));
 sg13g2_dlygate4sd3_1 hold2853 (.A(\atari2600.tia.p9_r ),
    .X(net7240));
 sg13g2_dlygate4sd3_1 hold2854 (.A(_02250_),
    .X(net7241));
 sg13g2_dlygate4sd3_1 hold2855 (.A(\rom_next_addr_in_queue[2] ),
    .X(net7242));
 sg13g2_dlygate4sd3_1 hold2856 (.A(_01140_),
    .X(net7243));
 sg13g2_dlygate4sd3_1 hold2857 (.A(\atari2600.tia.audio_right_counter[1] ),
    .X(net7244));
 sg13g2_dlygate4sd3_1 hold2858 (.A(_02029_),
    .X(net7245));
 sg13g2_dlygate4sd3_1 hold2859 (.A(\flash_rom.fsm_state[1] ),
    .X(net7246));
 sg13g2_dlygate4sd3_1 hold2860 (.A(\atari2600.tia.diag[56] ),
    .X(net7247));
 sg13g2_dlygate4sd3_1 hold2861 (.A(_02136_),
    .X(net7248));
 sg13g2_dlygate4sd3_1 hold2862 (.A(\atari2600.tia.diag[39] ),
    .X(net7249));
 sg13g2_dlygate4sd3_1 hold2863 (.A(\atari2600.tia.p1_spacing[5] ),
    .X(net7250));
 sg13g2_dlygate4sd3_1 hold2864 (.A(\atari2600.tia.diag[38] ),
    .X(net7251));
 sg13g2_dlygate4sd3_1 hold2865 (.A(\atari2600.tia.hmbl[2] ),
    .X(net7252));
 sg13g2_dlygate4sd3_1 hold2866 (.A(\atari2600.tia.ball_w[3] ),
    .X(net7253));
 sg13g2_dlygate4sd3_1 hold2867 (.A(\atari2600.tia.diag[44] ),
    .X(net7254));
 sg13g2_dlygate4sd3_1 hold2868 (.A(\atari2600.tia.p0_spacing[5] ),
    .X(net7255));
 sg13g2_dlygate4sd3_1 hold2869 (.A(\atari2600.tia.p0_spacing[6] ),
    .X(net7256));
 sg13g2_dlygate4sd3_1 hold2870 (.A(\atari2600.tia.poly9_r.x[2] ),
    .X(net7257));
 sg13g2_dlygate4sd3_1 hold2871 (.A(_07081_),
    .X(net7258));
 sg13g2_dlygate4sd3_1 hold2872 (.A(\atari2600.tia.poly9_r.x[7] ),
    .X(net7259));
 sg13g2_dlygate4sd3_1 hold2873 (.A(\atari2600.tia.diag[52] ),
    .X(net7260));
 sg13g2_dlygate4sd3_1 hold2874 (.A(\atari2600.tia.audc1[1] ),
    .X(net7261));
 sg13g2_dlygate4sd3_1 hold2875 (.A(\atari2600.tia.audf1[0] ),
    .X(net7262));
 sg13g2_dlygate4sd3_1 hold2876 (.A(\atari2600.tia.audf0[2] ),
    .X(net7263));
 sg13g2_dlygate4sd3_1 hold2877 (.A(\atari2600.tia.poly9_r.x[5] ),
    .X(net7264));
 sg13g2_dlygate4sd3_1 hold2878 (.A(_07085_),
    .X(net7265));
 sg13g2_dlygate4sd3_1 hold2879 (.A(\atari2600.tia.p0_scale[1] ),
    .X(net7266));
 sg13g2_dlygate4sd3_1 hold2880 (.A(\atari2600.tia.p1_scale[0] ),
    .X(net7267));
 sg13g2_dlygate4sd3_1 hold2881 (.A(\atari2600.tia.audc1[0] ),
    .X(net7268));
 sg13g2_dlygate4sd3_1 hold2882 (.A(_00062_),
    .X(net7269));
 sg13g2_dlygate4sd3_1 hold2883 (.A(_04646_),
    .X(net7270));
 sg13g2_dlygate4sd3_1 hold2884 (.A(_04649_),
    .X(net7271));
 sg13g2_dlygate4sd3_1 hold2885 (.A(\atari2600.tia.audf0[1] ),
    .X(net7272));
 sg13g2_dlygate4sd3_1 hold2886 (.A(\atari2600.tia.diag[41] ),
    .X(net7273));
 sg13g2_dlygate4sd3_1 hold2887 (.A(_02153_),
    .X(net7274));
 sg13g2_dlygate4sd3_1 hold2888 (.A(\atari2600.tia.audc0[1] ),
    .X(net7275));
 sg13g2_dlygate4sd3_1 hold2889 (.A(\atari2600.tia.poly9_r.x[6] ),
    .X(net7276));
 sg13g2_dlygate4sd3_1 hold2890 (.A(\atari2600.tia.audc0[0] ),
    .X(net7277));
 sg13g2_dlygate4sd3_1 hold2891 (.A(\atari2600.tia.diag[40] ),
    .X(net7278));
 sg13g2_dlygate4sd3_1 hold2892 (.A(\atari2600.cpu.ADD[7] ),
    .X(net7279));
 sg13g2_dlygate4sd3_1 hold2893 (.A(_00141_),
    .X(net7280));
 sg13g2_dlygate4sd3_1 hold2894 (.A(_07297_),
    .X(net7281));
 sg13g2_dlygate4sd3_1 hold2895 (.A(_02470_),
    .X(net7282));
 sg13g2_dlygate4sd3_1 hold2896 (.A(\atari2600.tia.audc0[3] ),
    .X(net7283));
 sg13g2_dlygate4sd3_1 hold2897 (.A(\atari2600.tia.diag[43] ),
    .X(net7284));
 sg13g2_dlygate4sd3_1 hold2898 (.A(\atari2600.tia.diag[64] ),
    .X(net7285));
 sg13g2_dlygate4sd3_1 hold2899 (.A(_02128_),
    .X(net7286));
 sg13g2_dlygate4sd3_1 hold2900 (.A(\atari2600.tia.diag[47] ),
    .X(net7287));
 sg13g2_dlygate4sd3_1 hold2901 (.A(\atari2600.tia.vdelp1 ),
    .X(net7288));
 sg13g2_dlygate4sd3_1 hold2902 (.A(\atari2600.tia.diag[57] ),
    .X(net7289));
 sg13g2_dlygate4sd3_1 hold2903 (.A(_02137_),
    .X(net7290));
 sg13g2_dlygate4sd3_1 hold2904 (.A(\atari2600.tia.audc1[3] ),
    .X(net7291));
 sg13g2_dlygate4sd3_1 hold2905 (.A(\atari2600.tia.vdelp0 ),
    .X(net7292));
 sg13g2_dlygate4sd3_1 hold2906 (.A(\atari2600.tia.audc0[2] ),
    .X(net7293));
 sg13g2_dlygate4sd3_1 hold2907 (.A(\rom_next_addr_in_queue[9] ),
    .X(net7294));
 sg13g2_dlygate4sd3_1 hold2908 (.A(_00063_),
    .X(net7295));
 sg13g2_dlygate4sd3_1 hold2909 (.A(\atari2600.tia.diag[65] ),
    .X(net7296));
 sg13g2_dlygate4sd3_1 hold2910 (.A(_02129_),
    .X(net7297));
 sg13g2_dlygate4sd3_1 hold2911 (.A(\atari2600.tia.diag[33] ),
    .X(net7298));
 sg13g2_dlygate4sd3_1 hold2912 (.A(_02161_),
    .X(net7299));
 sg13g2_dlygate4sd3_1 hold2913 (.A(\atari2600.tia.refpf ),
    .X(net7300));
 sg13g2_dlygate4sd3_1 hold2914 (.A(\atari2600.tia.diag[50] ),
    .X(net7301));
 sg13g2_dlygate4sd3_1 hold2915 (.A(\atari2600.tia.hmbl[3] ),
    .X(net7302));
 sg13g2_dlygate4sd3_1 hold2916 (.A(\atari2600.tia.diag[32] ),
    .X(net7303));
 sg13g2_dlygate4sd3_1 hold2917 (.A(\atari2600.tia.diag[37] ),
    .X(net7304));
 sg13g2_dlygate4sd3_1 hold2918 (.A(\atari2600.tia.diag[48] ),
    .X(net7305));
 sg13g2_dlygate4sd3_1 hold2919 (.A(\atari2600.tia.audio_r ),
    .X(net7306));
 sg13g2_dlygate4sd3_1 hold2920 (.A(_02045_),
    .X(net7307));
 sg13g2_dlygate4sd3_1 hold2921 (.A(\atari2600.cpu.ADD[1] ),
    .X(net7308));
 sg13g2_dlygate4sd3_1 hold2922 (.A(\atari2600.tia.diag[51] ),
    .X(net7309));
 sg13g2_dlygate4sd3_1 hold2923 (.A(_02147_),
    .X(net7310));
 sg13g2_dlygate4sd3_1 hold2924 (.A(\atari2600.tia.audf1[3] ),
    .X(net7311));
 sg13g2_dlygate4sd3_1 hold2925 (.A(\atari2600.tia.diag[42] ),
    .X(net7312));
 sg13g2_dlygate4sd3_1 hold2926 (.A(\atari2600.tia.p0_scale[0] ),
    .X(net7313));
 sg13g2_dlygate4sd3_1 hold2927 (.A(\b_pwm_odd[2] ),
    .X(net7314));
 sg13g2_dlygate4sd3_1 hold2928 (.A(_04410_),
    .X(net7315));
 sg13g2_dlygate4sd3_1 hold2929 (.A(\atari2600.tia.diag[34] ),
    .X(net7316));
 sg13g2_dlygate4sd3_1 hold2930 (.A(\atari2600.tia.diag[35] ),
    .X(net7317));
 sg13g2_dlygate4sd3_1 hold2931 (.A(\atari2600.tia.diag[45] ),
    .X(net7318));
 sg13g2_dlygate4sd3_1 hold2932 (.A(\atari2600.tia.p0_w[3] ),
    .X(net7319));
 sg13g2_dlygate4sd3_1 hold2933 (.A(_00154_),
    .X(net7320));
 sg13g2_dlygate4sd3_1 hold2934 (.A(\atari2600.tia.scorepf ),
    .X(net7321));
 sg13g2_dlygate4sd3_1 hold2935 (.A(\atari2600.cpu.ADD[5] ),
    .X(net7322));
 sg13g2_dlygate4sd3_1 hold2936 (.A(\hvsync_gen.hpos[8] ),
    .X(net7323));
 sg13g2_dlygate4sd3_1 hold2937 (.A(\atari2600.tia.p1_w[3] ),
    .X(net7324));
 sg13g2_dlygate4sd3_1 hold2938 (.A(\atari2600.cpu.ADD[4] ),
    .X(net7325));
 sg13g2_dlygate4sd3_1 hold2939 (.A(\hvsync_gen.hpos[4] ),
    .X(net7326));
 sg13g2_dlygate4sd3_1 hold2940 (.A(\atari2600.tia.diag[61] ),
    .X(net7327));
 sg13g2_dlygate4sd3_1 hold2941 (.A(\atari2600.tia.diag[54] ),
    .X(net7328));
 sg13g2_dlygate4sd3_1 hold2942 (.A(\atari2600.tia.diag[49] ),
    .X(net7329));
 sg13g2_dlygate4sd3_1 hold2943 (.A(\atari2600.tia.diag[58] ),
    .X(net7330));
 sg13g2_dlygate4sd3_1 hold2944 (.A(\atari2600.pia.underflow ),
    .X(net7331));
 sg13g2_dlygate4sd3_1 hold2945 (.A(_01796_),
    .X(net7332));
 sg13g2_dlygate4sd3_1 hold2946 (.A(\atari2600.tia.audf0[3] ),
    .X(net7333));
 sg13g2_dlygate4sd3_1 hold2947 (.A(\atari2600.tia.diag[62] ),
    .X(net7334));
 sg13g2_dlygate4sd3_1 hold2948 (.A(\atari2600.address_bus_r[8] ),
    .X(net7335));
 sg13g2_dlygate4sd3_1 hold2949 (.A(\atari2600.address_bus_r[0] ),
    .X(net7336));
 sg13g2_dlygate4sd3_1 hold2950 (.A(\atari2600.tia.diag[71] ),
    .X(net7337));
 sg13g2_dlygate4sd3_1 hold2951 (.A(\r_pwm_even[3] ),
    .X(net7338));
 sg13g2_dlygate4sd3_1 hold2952 (.A(_04580_),
    .X(net7339));
 sg13g2_dlygate4sd3_1 hold2953 (.A(\atari2600.tia.diag[59] ),
    .X(net7340));
 sg13g2_dlygate4sd3_1 hold2954 (.A(\atari2600.tia.hmm1[3] ),
    .X(net7341));
 sg13g2_dlygate4sd3_1 hold2955 (.A(\atari2600.cpu.DIHOLD[7] ),
    .X(net7342));
 sg13g2_dlygate4sd3_1 hold2956 (.A(\atari2600.tia.audf1[1] ),
    .X(net7343));
 sg13g2_dlygate4sd3_1 hold2957 (.A(\atari2600.cpu.ADD[6] ),
    .X(net7344));
 sg13g2_dlygate4sd3_1 hold2958 (.A(\atari2600.tia.diag[67] ),
    .X(net7345));
 sg13g2_dlygate4sd3_1 hold2959 (.A(\atari2600.tia.diag[63] ),
    .X(net7346));
 sg13g2_dlygate4sd3_1 hold2960 (.A(_00094_),
    .X(net7347));
 sg13g2_dlygate4sd3_1 hold2961 (.A(_08191_),
    .X(net7348));
 sg13g2_dlygate4sd3_1 hold2962 (.A(\atari2600.cpu.ADD[3] ),
    .X(net7349));
 sg13g2_dlygate4sd3_1 hold2963 (.A(\atari2600.tia.diag[53] ),
    .X(net7350));
 sg13g2_dlygate4sd3_1 hold2964 (.A(\atari2600.tia.audc1[2] ),
    .X(net7351));
 sg13g2_dlygate4sd3_1 hold2965 (.A(\atari2600.tia.diag[69] ),
    .X(net7352));
 sg13g2_dlygate4sd3_1 hold2966 (.A(\atari2600.tia.diag[60] ),
    .X(net7353));
 sg13g2_dlygate4sd3_1 hold2967 (.A(\atari2600.tia.audf1[2] ),
    .X(net7354));
 sg13g2_dlygate4sd3_1 hold2968 (.A(\atari2600.tia.diag[70] ),
    .X(net7355));
 sg13g2_dlygate4sd3_1 hold2969 (.A(_00156_),
    .X(net7356));
 sg13g2_dlygate4sd3_1 hold2970 (.A(\flash_rom.fsm_state[2] ),
    .X(net7357));
 sg13g2_dlygate4sd3_1 hold2971 (.A(\atari2600.tia.diag[66] ),
    .X(net7358));
 sg13g2_dlygate4sd3_1 hold2972 (.A(_00164_),
    .X(net7359));
 sg13g2_dlygate4sd3_1 hold2973 (.A(\audio_pwm_accumulator[4] ),
    .X(net7360));
 sg13g2_dlygate4sd3_1 hold2974 (.A(\atari2600.cpu.ADD[2] ),
    .X(net7361));
 sg13g2_dlygate4sd3_1 hold2975 (.A(\atari2600.cpu.DIHOLD[5] ),
    .X(net7362));
 sg13g2_dlygate4sd3_1 hold2976 (.A(\atari2600.cpu.DIMUX[5] ),
    .X(net7363));
 sg13g2_dlygate4sd3_1 hold2977 (.A(\atari2600.stall_cpu ),
    .X(net7364));
 sg13g2_dlygate4sd3_1 hold2978 (.A(_00088_),
    .X(net7365));
 sg13g2_dlygate4sd3_1 hold2979 (.A(_00146_),
    .X(net7366));
 sg13g2_dlygate4sd3_1 hold2980 (.A(\atari2600.cpu.plp ),
    .X(net7367));
 sg13g2_dlygate4sd3_1 hold2981 (.A(_00165_),
    .X(net7368));
 sg13g2_dlygate4sd3_1 hold2982 (.A(\hvsync_gen.vga.vpos[8] ),
    .X(net7369));
 sg13g2_dlygate4sd3_1 hold2983 (.A(_08493_),
    .X(net7370));
 sg13g2_dlygate4sd3_1 hold2984 (.A(_08495_),
    .X(net7371));
 sg13g2_dlygate4sd3_1 hold2985 (.A(\atari2600.address_bus_r[9] ),
    .X(net7372));
 sg13g2_dlygate4sd3_1 hold2986 (.A(_00150_),
    .X(net7373));
 sg13g2_dlygate4sd3_1 hold2987 (.A(\atari2600.cpu.ADD[0] ),
    .X(net7374));
 sg13g2_dlygate4sd3_1 hold2988 (.A(\b_pwm_odd[1] ),
    .X(net7375));
 sg13g2_dlygate4sd3_1 hold2989 (.A(\hvsync_gen.vga.vpos[6] ),
    .X(net7376));
 sg13g2_dlygate4sd3_1 hold2990 (.A(\atari2600.pia.diag[0] ),
    .X(net7377));
 sg13g2_dlygate4sd3_1 hold2991 (.A(_05246_),
    .X(net7378));
 sg13g2_dlygate4sd3_1 hold2992 (.A(\atari2600.tia.cx_clr ),
    .X(net7379));
 sg13g2_dlygate4sd3_1 hold2993 (.A(\atari2600.tia.enam0 ),
    .X(net7380));
 sg13g2_antennanp ANTENNA_1 (.A(_00001_));
 sg13g2_antennanp ANTENNA_2 (.A(_00008_));
 sg13g2_antennanp ANTENNA_3 (.A(_00013_));
 sg13g2_antennanp ANTENNA_4 (.A(_01155_));
 sg13g2_antennanp ANTENNA_5 (.A(_01163_));
 sg13g2_antennanp ANTENNA_6 (.A(_01778_));
 sg13g2_antennanp ANTENNA_7 (.A(_01782_));
 sg13g2_antennanp ANTENNA_8 (.A(_03601_));
 sg13g2_antennanp ANTENNA_9 (.A(_05302_));
 sg13g2_antennanp ANTENNA_10 (.A(_05334_));
 sg13g2_antennanp ANTENNA_11 (.A(_05334_));
 sg13g2_antennanp ANTENNA_12 (.A(_07899_));
 sg13g2_antennanp ANTENNA_13 (.A(_07910_));
 sg13g2_antennanp ANTENNA_14 (.A(_07918_));
 sg13g2_antennanp ANTENNA_15 (.A(_08164_));
 sg13g2_antennanp ANTENNA_16 (.A(_10257_));
 sg13g2_antennanp ANTENNA_17 (.A(_10257_));
 sg13g2_antennanp ANTENNA_18 (.A(\atari2600.input_joystick_0[1] ));
 sg13g2_antennanp ANTENNA_19 (.A(\atari2600.input_joystick_0[1] ));
 sg13g2_antennanp ANTENNA_20 (.A(\atari2600.input_joystick_0[1] ));
 sg13g2_antennanp ANTENNA_21 (.A(\atari2600.input_joystick_0[1] ));
 sg13g2_antennanp ANTENNA_22 (.A(clk));
 sg13g2_antennanp ANTENNA_23 (.A(clk));
 sg13g2_antennanp ANTENNA_24 (.A(rom_data_pending));
 sg13g2_antennanp ANTENNA_25 (.A(rom_data_pending));
 sg13g2_antennanp ANTENNA_26 (.A(rom_data_pending));
 sg13g2_antennanp ANTENNA_27 (.A(rom_data_pending));
 sg13g2_antennanp ANTENNA_28 (.A(net4875));
 sg13g2_antennanp ANTENNA_29 (.A(net4875));
 sg13g2_antennanp ANTENNA_30 (.A(net4875));
 sg13g2_antennanp ANTENNA_31 (.A(net4875));
 sg13g2_antennanp ANTENNA_32 (.A(net4875));
 sg13g2_antennanp ANTENNA_33 (.A(net4875));
 sg13g2_antennanp ANTENNA_34 (.A(net4875));
 sg13g2_antennanp ANTENNA_35 (.A(net4875));
 sg13g2_antennanp ANTENNA_36 (.A(net4875));
 sg13g2_antennanp ANTENNA_37 (.A(net4875));
 sg13g2_antennanp ANTENNA_38 (.A(net4875));
 sg13g2_antennanp ANTENNA_39 (.A(net4875));
 sg13g2_antennanp ANTENNA_40 (.A(net5682));
 sg13g2_antennanp ANTENNA_41 (.A(net5682));
 sg13g2_antennanp ANTENNA_42 (.A(net5682));
 sg13g2_antennanp ANTENNA_43 (.A(net5682));
 sg13g2_antennanp ANTENNA_44 (.A(_00001_));
 sg13g2_antennanp ANTENNA_45 (.A(_00002_));
 sg13g2_antennanp ANTENNA_46 (.A(_00005_));
 sg13g2_antennanp ANTENNA_47 (.A(_00006_));
 sg13g2_antennanp ANTENNA_48 (.A(_00007_));
 sg13g2_antennanp ANTENNA_49 (.A(_00013_));
 sg13g2_antennanp ANTENNA_50 (.A(_01155_));
 sg13g2_antennanp ANTENNA_51 (.A(_01199_));
 sg13g2_antennanp ANTENNA_52 (.A(_01773_));
 sg13g2_antennanp ANTENNA_53 (.A(_01778_));
 sg13g2_antennanp ANTENNA_54 (.A(_01784_));
 sg13g2_antennanp ANTENNA_55 (.A(_01784_));
 sg13g2_antennanp ANTENNA_56 (.A(_01787_));
 sg13g2_antennanp ANTENNA_57 (.A(_01788_));
 sg13g2_antennanp ANTENNA_58 (.A(_01788_));
 sg13g2_antennanp ANTENNA_59 (.A(_01793_));
 sg13g2_antennanp ANTENNA_60 (.A(_01793_));
 sg13g2_antennanp ANTENNA_61 (.A(_01793_));
 sg13g2_antennanp ANTENNA_62 (.A(_03601_));
 sg13g2_antennanp ANTENNA_63 (.A(_05302_));
 sg13g2_antennanp ANTENNA_64 (.A(_07899_));
 sg13g2_antennanp ANTENNA_65 (.A(_07910_));
 sg13g2_antennanp ANTENNA_66 (.A(_07918_));
 sg13g2_antennanp ANTENNA_67 (.A(_08164_));
 sg13g2_antennanp ANTENNA_68 (.A(_10257_));
 sg13g2_antennanp ANTENNA_69 (.A(_10257_));
 sg13g2_antennanp ANTENNA_70 (.A(\atari2600.input_joystick_0[1] ));
 sg13g2_antennanp ANTENNA_71 (.A(\atari2600.input_joystick_0[1] ));
 sg13g2_antennanp ANTENNA_72 (.A(\atari2600.tia.hmbl[3] ));
 sg13g2_antennanp ANTENNA_73 (.A(\atari2600.tia.hmbl[3] ));
 sg13g2_antennanp ANTENNA_74 (.A(\atari2600.tia.hmbl[3] ));
 sg13g2_antennanp ANTENNA_75 (.A(\atari2600.tia.hmbl[3] ));
 sg13g2_antennanp ANTENNA_76 (.A(\atari2600.tia.hmbl[3] ));
 sg13g2_antennanp ANTENNA_77 (.A(clk));
 sg13g2_antennanp ANTENNA_78 (.A(clk));
 sg13g2_antennanp ANTENNA_79 (.A(rom_data_pending));
 sg13g2_antennanp ANTENNA_80 (.A(rom_data_pending));
 sg13g2_antennanp ANTENNA_81 (.A(rom_data_pending));
 sg13g2_antennanp ANTENNA_82 (.A(rom_data_pending));
 sg13g2_antennanp ANTENNA_83 (.A(net5682));
 sg13g2_antennanp ANTENNA_84 (.A(net5682));
 sg13g2_antennanp ANTENNA_85 (.A(net5682));
 sg13g2_antennanp ANTENNA_86 (.A(net5682));
 sg13g2_antennanp ANTENNA_87 (.A(_00001_));
 sg13g2_antennanp ANTENNA_88 (.A(_00002_));
 sg13g2_antennanp ANTENNA_89 (.A(_00006_));
 sg13g2_antennanp ANTENNA_90 (.A(_00008_));
 sg13g2_antennanp ANTENNA_91 (.A(_00013_));
 sg13g2_antennanp ANTENNA_92 (.A(_01155_));
 sg13g2_antennanp ANTENNA_93 (.A(_01199_));
 sg13g2_antennanp ANTENNA_94 (.A(_01773_));
 sg13g2_antennanp ANTENNA_95 (.A(_01778_));
 sg13g2_antennanp ANTENNA_96 (.A(_01782_));
 sg13g2_antennanp ANTENNA_97 (.A(_01784_));
 sg13g2_antennanp ANTENNA_98 (.A(_01787_));
 sg13g2_antennanp ANTENNA_99 (.A(_01788_));
 sg13g2_antennanp ANTENNA_100 (.A(_03601_));
 sg13g2_antennanp ANTENNA_101 (.A(_05302_));
 sg13g2_antennanp ANTENNA_102 (.A(_05334_));
 sg13g2_antennanp ANTENNA_103 (.A(_07756_));
 sg13g2_antennanp ANTENNA_104 (.A(_07910_));
 sg13g2_antennanp ANTENNA_105 (.A(_07918_));
 sg13g2_antennanp ANTENNA_106 (.A(_08164_));
 sg13g2_antennanp ANTENNA_107 (.A(_10257_));
 sg13g2_antennanp ANTENNA_108 (.A(_10257_));
 sg13g2_antennanp ANTENNA_109 (.A(\atari2600.input_joystick_0[1] ));
 sg13g2_antennanp ANTENNA_110 (.A(\atari2600.input_joystick_0[1] ));
 sg13g2_antennanp ANTENNA_111 (.A(clk));
 sg13g2_antennanp ANTENNA_112 (.A(clk));
 sg13g2_antennanp ANTENNA_113 (.A(rom_data_pending));
 sg13g2_antennanp ANTENNA_114 (.A(rom_data_pending));
 sg13g2_antennanp ANTENNA_115 (.A(rom_data_pending));
 sg13g2_antennanp ANTENNA_116 (.A(rom_data_pending));
 sg13g2_antennanp ANTENNA_117 (.A(net5682));
 sg13g2_antennanp ANTENNA_118 (.A(net5682));
 sg13g2_antennanp ANTENNA_119 (.A(net5682));
 sg13g2_antennanp ANTENNA_120 (.A(net5682));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_fill_1 FILLER_0_161 ();
 sg13g2_fill_1 FILLER_0_350 ();
 sg13g2_fill_2 FILLER_0_364 ();
 sg13g2_fill_2 FILLER_0_416 ();
 sg13g2_fill_1 FILLER_0_432 ();
 sg13g2_fill_2 FILLER_0_472 ();
 sg13g2_fill_1 FILLER_0_474 ();
 sg13g2_fill_2 FILLER_0_518 ();
 sg13g2_fill_1 FILLER_0_564 ();
 sg13g2_fill_2 FILLER_0_610 ();
 sg13g2_fill_1 FILLER_0_612 ();
 sg13g2_fill_1 FILLER_0_682 ();
 sg13g2_fill_1 FILLER_0_687 ();
 sg13g2_fill_2 FILLER_0_777 ();
 sg13g2_fill_1 FILLER_0_889 ();
 sg13g2_fill_2 FILLER_0_995 ();
 sg13g2_fill_1 FILLER_0_1023 ();
 sg13g2_fill_2 FILLER_0_1050 ();
 sg13g2_fill_1 FILLER_0_1052 ();
 sg13g2_fill_2 FILLER_0_1092 ();
 sg13g2_fill_2 FILLER_0_1112 ();
 sg13g2_fill_1 FILLER_0_1124 ();
 sg13g2_fill_1 FILLER_0_1133 ();
 sg13g2_fill_1 FILLER_0_1169 ();
 sg13g2_fill_1 FILLER_0_1212 ();
 sg13g2_fill_2 FILLER_0_1297 ();
 sg13g2_fill_2 FILLER_0_1343 ();
 sg13g2_fill_1 FILLER_0_1345 ();
 sg13g2_decap_4 FILLER_0_1381 ();
 sg13g2_fill_2 FILLER_0_1459 ();
 sg13g2_fill_1 FILLER_0_1461 ();
 sg13g2_fill_2 FILLER_0_1516 ();
 sg13g2_fill_2 FILLER_0_1590 ();
 sg13g2_fill_2 FILLER_0_1605 ();
 sg13g2_fill_1 FILLER_0_1617 ();
 sg13g2_fill_2 FILLER_0_1662 ();
 sg13g2_fill_1 FILLER_0_1664 ();
 sg13g2_fill_2 FILLER_0_1704 ();
 sg13g2_fill_1 FILLER_0_1706 ();
 sg13g2_fill_2 FILLER_0_1749 ();
 sg13g2_fill_1 FILLER_0_1751 ();
 sg13g2_fill_1 FILLER_0_1776 ();
 sg13g2_fill_2 FILLER_0_1787 ();
 sg13g2_fill_2 FILLER_0_1830 ();
 sg13g2_fill_1 FILLER_0_1832 ();
 sg13g2_fill_1 FILLER_0_1903 ();
 sg13g2_fill_2 FILLER_0_1928 ();
 sg13g2_fill_1 FILLER_0_1930 ();
 sg13g2_fill_2 FILLER_0_1987 ();
 sg13g2_fill_1 FILLER_0_1989 ();
 sg13g2_fill_2 FILLER_0_2068 ();
 sg13g2_fill_1 FILLER_0_2070 ();
 sg13g2_fill_2 FILLER_0_2092 ();
 sg13g2_fill_1 FILLER_0_2094 ();
 sg13g2_fill_2 FILLER_0_2113 ();
 sg13g2_fill_2 FILLER_0_2198 ();
 sg13g2_fill_1 FILLER_0_2200 ();
 sg13g2_fill_2 FILLER_0_2246 ();
 sg13g2_fill_1 FILLER_0_2248 ();
 sg13g2_fill_2 FILLER_0_2288 ();
 sg13g2_fill_2 FILLER_0_2313 ();
 sg13g2_fill_1 FILLER_0_2315 ();
 sg13g2_fill_2 FILLER_0_2342 ();
 sg13g2_fill_1 FILLER_0_2344 ();
 sg13g2_fill_1 FILLER_0_2355 ();
 sg13g2_fill_2 FILLER_0_2408 ();
 sg13g2_fill_2 FILLER_0_2465 ();
 sg13g2_fill_1 FILLER_0_2467 ();
 sg13g2_fill_2 FILLER_0_2486 ();
 sg13g2_decap_8 FILLER_0_2545 ();
 sg13g2_decap_8 FILLER_0_2552 ();
 sg13g2_decap_8 FILLER_0_2559 ();
 sg13g2_decap_8 FILLER_0_2566 ();
 sg13g2_decap_8 FILLER_0_2573 ();
 sg13g2_decap_8 FILLER_0_2580 ();
 sg13g2_decap_8 FILLER_0_2587 ();
 sg13g2_decap_8 FILLER_0_2594 ();
 sg13g2_decap_8 FILLER_0_2601 ();
 sg13g2_decap_8 FILLER_0_2608 ();
 sg13g2_decap_8 FILLER_0_2615 ();
 sg13g2_decap_8 FILLER_0_2622 ();
 sg13g2_decap_8 FILLER_0_2629 ();
 sg13g2_decap_8 FILLER_0_2636 ();
 sg13g2_decap_8 FILLER_0_2643 ();
 sg13g2_decap_8 FILLER_0_2650 ();
 sg13g2_decap_8 FILLER_0_2657 ();
 sg13g2_decap_8 FILLER_0_2664 ();
 sg13g2_fill_2 FILLER_0_2671 ();
 sg13g2_fill_1 FILLER_0_2673 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_4 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_153 ();
 sg13g2_decap_8 FILLER_1_160 ();
 sg13g2_decap_4 FILLER_1_167 ();
 sg13g2_fill_2 FILLER_1_171 ();
 sg13g2_fill_1 FILLER_1_220 ();
 sg13g2_fill_2 FILLER_1_248 ();
 sg13g2_fill_2 FILLER_1_284 ();
 sg13g2_fill_1 FILLER_1_491 ();
 sg13g2_fill_2 FILLER_1_574 ();
 sg13g2_fill_1 FILLER_1_576 ();
 sg13g2_fill_1 FILLER_1_707 ();
 sg13g2_fill_2 FILLER_1_762 ();
 sg13g2_fill_1 FILLER_1_764 ();
 sg13g2_fill_2 FILLER_1_810 ();
 sg13g2_fill_1 FILLER_1_812 ();
 sg13g2_fill_2 FILLER_1_903 ();
 sg13g2_fill_1 FILLER_1_940 ();
 sg13g2_fill_2 FILLER_1_990 ();
 sg13g2_fill_1 FILLER_1_1002 ();
 sg13g2_fill_2 FILLER_1_1051 ();
 sg13g2_fill_1 FILLER_1_1063 ();
 sg13g2_fill_2 FILLER_1_1146 ();
 sg13g2_fill_1 FILLER_1_1148 ();
 sg13g2_fill_1 FILLER_1_1278 ();
 sg13g2_fill_2 FILLER_1_1348 ();
 sg13g2_fill_2 FILLER_1_1433 ();
 sg13g2_fill_2 FILLER_1_1581 ();
 sg13g2_fill_2 FILLER_1_1613 ();
 sg13g2_fill_2 FILLER_1_1668 ();
 sg13g2_fill_1 FILLER_1_1670 ();
 sg13g2_fill_2 FILLER_1_1715 ();
 sg13g2_fill_1 FILLER_1_1717 ();
 sg13g2_fill_2 FILLER_1_1881 ();
 sg13g2_fill_1 FILLER_1_1935 ();
 sg13g2_fill_2 FILLER_1_1960 ();
 sg13g2_fill_1 FILLER_1_1962 ();
 sg13g2_fill_1 FILLER_1_2050 ();
 sg13g2_fill_2 FILLER_1_2087 ();
 sg13g2_fill_1 FILLER_1_2089 ();
 sg13g2_fill_1 FILLER_1_2116 ();
 sg13g2_fill_2 FILLER_1_2157 ();
 sg13g2_fill_1 FILLER_1_2159 ();
 sg13g2_fill_2 FILLER_1_2199 ();
 sg13g2_fill_2 FILLER_1_2220 ();
 sg13g2_fill_1 FILLER_1_2222 ();
 sg13g2_fill_2 FILLER_1_2263 ();
 sg13g2_fill_1 FILLER_1_2265 ();
 sg13g2_fill_2 FILLER_1_2302 ();
 sg13g2_fill_2 FILLER_1_2330 ();
 sg13g2_fill_2 FILLER_1_2509 ();
 sg13g2_fill_1 FILLER_1_2511 ();
 sg13g2_fill_1 FILLER_1_2550 ();
 sg13g2_decap_8 FILLER_1_2555 ();
 sg13g2_decap_8 FILLER_1_2562 ();
 sg13g2_decap_4 FILLER_1_2569 ();
 sg13g2_decap_8 FILLER_1_2582 ();
 sg13g2_decap_8 FILLER_1_2589 ();
 sg13g2_decap_8 FILLER_1_2596 ();
 sg13g2_decap_8 FILLER_1_2603 ();
 sg13g2_decap_8 FILLER_1_2610 ();
 sg13g2_decap_8 FILLER_1_2617 ();
 sg13g2_decap_8 FILLER_1_2624 ();
 sg13g2_decap_8 FILLER_1_2631 ();
 sg13g2_decap_8 FILLER_1_2638 ();
 sg13g2_decap_8 FILLER_1_2645 ();
 sg13g2_decap_8 FILLER_1_2652 ();
 sg13g2_decap_8 FILLER_1_2659 ();
 sg13g2_decap_8 FILLER_1_2666 ();
 sg13g2_fill_1 FILLER_1_2673 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_fill_1 FILLER_2_133 ();
 sg13g2_decap_4 FILLER_2_138 ();
 sg13g2_fill_2 FILLER_2_152 ();
 sg13g2_fill_1 FILLER_2_154 ();
 sg13g2_fill_1 FILLER_2_159 ();
 sg13g2_fill_2 FILLER_2_179 ();
 sg13g2_fill_1 FILLER_2_181 ();
 sg13g2_fill_2 FILLER_2_192 ();
 sg13g2_fill_1 FILLER_2_194 ();
 sg13g2_fill_1 FILLER_2_205 ();
 sg13g2_fill_2 FILLER_2_219 ();
 sg13g2_fill_2 FILLER_2_304 ();
 sg13g2_fill_1 FILLER_2_318 ();
 sg13g2_fill_2 FILLER_2_350 ();
 sg13g2_fill_1 FILLER_2_352 ();
 sg13g2_fill_1 FILLER_2_393 ();
 sg13g2_fill_2 FILLER_2_403 ();
 sg13g2_fill_1 FILLER_2_405 ();
 sg13g2_fill_1 FILLER_2_484 ();
 sg13g2_fill_2 FILLER_2_495 ();
 sg13g2_fill_1 FILLER_2_497 ();
 sg13g2_fill_1 FILLER_2_511 ();
 sg13g2_fill_1 FILLER_2_525 ();
 sg13g2_fill_1 FILLER_2_578 ();
 sg13g2_fill_2 FILLER_2_647 ();
 sg13g2_fill_1 FILLER_2_649 ();
 sg13g2_fill_2 FILLER_2_669 ();
 sg13g2_fill_1 FILLER_2_671 ();
 sg13g2_fill_1 FILLER_2_682 ();
 sg13g2_fill_1 FILLER_2_696 ();
 sg13g2_fill_1 FILLER_2_733 ();
 sg13g2_fill_2 FILLER_2_800 ();
 sg13g2_fill_1 FILLER_2_828 ();
 sg13g2_fill_2 FILLER_2_852 ();
 sg13g2_fill_1 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_898 ();
 sg13g2_fill_1 FILLER_2_914 ();
 sg13g2_fill_1 FILLER_2_960 ();
 sg13g2_fill_1 FILLER_2_1031 ();
 sg13g2_fill_1 FILLER_2_1067 ();
 sg13g2_fill_2 FILLER_2_1131 ();
 sg13g2_fill_2 FILLER_2_1147 ();
 sg13g2_fill_2 FILLER_2_1250 ();
 sg13g2_fill_1 FILLER_2_1282 ();
 sg13g2_fill_1 FILLER_2_1292 ();
 sg13g2_fill_1 FILLER_2_1303 ();
 sg13g2_fill_2 FILLER_2_1309 ();
 sg13g2_fill_1 FILLER_2_1311 ();
 sg13g2_fill_1 FILLER_2_1342 ();
 sg13g2_fill_1 FILLER_2_1353 ();
 sg13g2_fill_1 FILLER_2_1420 ();
 sg13g2_fill_1 FILLER_2_1488 ();
 sg13g2_fill_2 FILLER_2_1550 ();
 sg13g2_fill_2 FILLER_2_1619 ();
 sg13g2_fill_2 FILLER_2_1700 ();
 sg13g2_fill_2 FILLER_2_1737 ();
 sg13g2_fill_1 FILLER_2_1739 ();
 sg13g2_fill_2 FILLER_2_1827 ();
 sg13g2_fill_2 FILLER_2_1843 ();
 sg13g2_fill_1 FILLER_2_1845 ();
 sg13g2_fill_2 FILLER_2_1876 ();
 sg13g2_fill_1 FILLER_2_1878 ();
 sg13g2_fill_2 FILLER_2_1909 ();
 sg13g2_fill_1 FILLER_2_1911 ();
 sg13g2_fill_1 FILLER_2_1922 ();
 sg13g2_fill_1 FILLER_2_1974 ();
 sg13g2_fill_2 FILLER_2_2053 ();
 sg13g2_fill_2 FILLER_2_2095 ();
 sg13g2_fill_1 FILLER_2_2097 ();
 sg13g2_fill_2 FILLER_2_2184 ();
 sg13g2_fill_1 FILLER_2_2186 ();
 sg13g2_fill_1 FILLER_2_2227 ();
 sg13g2_fill_2 FILLER_2_2297 ();
 sg13g2_fill_2 FILLER_2_2337 ();
 sg13g2_fill_1 FILLER_2_2360 ();
 sg13g2_fill_2 FILLER_2_2413 ();
 sg13g2_fill_1 FILLER_2_2442 ();
 sg13g2_fill_2 FILLER_2_2457 ();
 sg13g2_fill_2 FILLER_2_2507 ();
 sg13g2_fill_2 FILLER_2_2523 ();
 sg13g2_fill_1 FILLER_2_2525 ();
 sg13g2_fill_2 FILLER_2_2551 ();
 sg13g2_fill_2 FILLER_2_2558 ();
 sg13g2_fill_2 FILLER_2_2574 ();
 sg13g2_fill_1 FILLER_2_2576 ();
 sg13g2_decap_8 FILLER_2_2587 ();
 sg13g2_fill_2 FILLER_2_2594 ();
 sg13g2_decap_8 FILLER_2_2609 ();
 sg13g2_decap_8 FILLER_2_2616 ();
 sg13g2_decap_8 FILLER_2_2623 ();
 sg13g2_decap_8 FILLER_2_2630 ();
 sg13g2_decap_8 FILLER_2_2637 ();
 sg13g2_decap_8 FILLER_2_2644 ();
 sg13g2_decap_8 FILLER_2_2651 ();
 sg13g2_decap_8 FILLER_2_2658 ();
 sg13g2_decap_8 FILLER_2_2665 ();
 sg13g2_fill_2 FILLER_2_2672 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_4 FILLER_3_112 ();
 sg13g2_fill_2 FILLER_3_194 ();
 sg13g2_fill_1 FILLER_3_206 ();
 sg13g2_fill_1 FILLER_3_252 ();
 sg13g2_fill_2 FILLER_3_287 ();
 sg13g2_fill_1 FILLER_3_289 ();
 sg13g2_fill_1 FILLER_3_374 ();
 sg13g2_fill_1 FILLER_3_546 ();
 sg13g2_fill_1 FILLER_3_572 ();
 sg13g2_fill_1 FILLER_3_708 ();
 sg13g2_fill_1 FILLER_3_761 ();
 sg13g2_fill_2 FILLER_3_776 ();
 sg13g2_fill_1 FILLER_3_778 ();
 sg13g2_fill_2 FILLER_3_807 ();
 sg13g2_fill_1 FILLER_3_809 ();
 sg13g2_fill_2 FILLER_3_859 ();
 sg13g2_fill_2 FILLER_3_918 ();
 sg13g2_fill_1 FILLER_3_920 ();
 sg13g2_fill_2 FILLER_3_956 ();
 sg13g2_fill_1 FILLER_3_1000 ();
 sg13g2_fill_2 FILLER_3_1016 ();
 sg13g2_fill_1 FILLER_3_1018 ();
 sg13g2_fill_2 FILLER_3_1028 ();
 sg13g2_fill_2 FILLER_3_1093 ();
 sg13g2_fill_1 FILLER_3_1149 ();
 sg13g2_fill_1 FILLER_3_1160 ();
 sg13g2_fill_2 FILLER_3_1273 ();
 sg13g2_fill_2 FILLER_3_1345 ();
 sg13g2_fill_1 FILLER_3_1439 ();
 sg13g2_fill_1 FILLER_3_1458 ();
 sg13g2_fill_2 FILLER_3_1490 ();
 sg13g2_fill_1 FILLER_3_1513 ();
 sg13g2_fill_2 FILLER_3_1543 ();
 sg13g2_fill_1 FILLER_3_1545 ();
 sg13g2_fill_1 FILLER_3_1560 ();
 sg13g2_fill_2 FILLER_3_1600 ();
 sg13g2_fill_1 FILLER_3_1630 ();
 sg13g2_fill_1 FILLER_3_1666 ();
 sg13g2_fill_2 FILLER_3_1689 ();
 sg13g2_fill_1 FILLER_3_1691 ();
 sg13g2_fill_2 FILLER_3_1728 ();
 sg13g2_fill_1 FILLER_3_1730 ();
 sg13g2_fill_1 FILLER_3_1777 ();
 sg13g2_fill_1 FILLER_3_1797 ();
 sg13g2_fill_2 FILLER_3_1970 ();
 sg13g2_fill_1 FILLER_3_1972 ();
 sg13g2_fill_2 FILLER_3_2017 ();
 sg13g2_fill_1 FILLER_3_2019 ();
 sg13g2_fill_1 FILLER_3_2079 ();
 sg13g2_fill_2 FILLER_3_2131 ();
 sg13g2_fill_1 FILLER_3_2133 ();
 sg13g2_fill_2 FILLER_3_2206 ();
 sg13g2_fill_1 FILLER_3_2208 ();
 sg13g2_fill_2 FILLER_3_2219 ();
 sg13g2_fill_1 FILLER_3_2221 ();
 sg13g2_fill_1 FILLER_3_2271 ();
 sg13g2_fill_2 FILLER_3_2293 ();
 sg13g2_fill_1 FILLER_3_2295 ();
 sg13g2_fill_1 FILLER_3_2343 ();
 sg13g2_fill_2 FILLER_3_2398 ();
 sg13g2_fill_1 FILLER_3_2400 ();
 sg13g2_fill_2 FILLER_3_2474 ();
 sg13g2_fill_1 FILLER_3_2476 ();
 sg13g2_fill_2 FILLER_3_2517 ();
 sg13g2_fill_1 FILLER_3_2519 ();
 sg13g2_fill_2 FILLER_3_2582 ();
 sg13g2_fill_1 FILLER_3_2584 ();
 sg13g2_decap_8 FILLER_3_2611 ();
 sg13g2_decap_8 FILLER_3_2618 ();
 sg13g2_decap_8 FILLER_3_2625 ();
 sg13g2_decap_8 FILLER_3_2632 ();
 sg13g2_decap_8 FILLER_3_2639 ();
 sg13g2_decap_8 FILLER_3_2646 ();
 sg13g2_decap_8 FILLER_3_2653 ();
 sg13g2_decap_8 FILLER_3_2660 ();
 sg13g2_decap_8 FILLER_3_2667 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_fill_2 FILLER_4_164 ();
 sg13g2_fill_1 FILLER_4_166 ();
 sg13g2_fill_2 FILLER_4_281 ();
 sg13g2_fill_1 FILLER_4_283 ();
 sg13g2_fill_2 FILLER_4_308 ();
 sg13g2_fill_1 FILLER_4_351 ();
 sg13g2_fill_2 FILLER_4_390 ();
 sg13g2_fill_1 FILLER_4_392 ();
 sg13g2_fill_1 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_444 ();
 sg13g2_fill_1 FILLER_4_465 ();
 sg13g2_fill_1 FILLER_4_551 ();
 sg13g2_fill_2 FILLER_4_607 ();
 sg13g2_fill_2 FILLER_4_635 ();
 sg13g2_fill_1 FILLER_4_669 ();
 sg13g2_fill_1 FILLER_4_729 ();
 sg13g2_fill_1 FILLER_4_740 ();
 sg13g2_fill_2 FILLER_4_756 ();
 sg13g2_fill_1 FILLER_4_758 ();
 sg13g2_fill_2 FILLER_4_795 ();
 sg13g2_fill_2 FILLER_4_861 ();
 sg13g2_fill_2 FILLER_4_887 ();
 sg13g2_fill_1 FILLER_4_889 ();
 sg13g2_fill_1 FILLER_4_947 ();
 sg13g2_fill_2 FILLER_4_966 ();
 sg13g2_fill_1 FILLER_4_1020 ();
 sg13g2_fill_1 FILLER_4_1051 ();
 sg13g2_fill_2 FILLER_4_1068 ();
 sg13g2_fill_1 FILLER_4_1114 ();
 sg13g2_fill_2 FILLER_4_1124 ();
 sg13g2_fill_1 FILLER_4_1126 ();
 sg13g2_fill_2 FILLER_4_1206 ();
 sg13g2_fill_2 FILLER_4_1239 ();
 sg13g2_fill_1 FILLER_4_1297 ();
 sg13g2_fill_2 FILLER_4_1304 ();
 sg13g2_fill_1 FILLER_4_1306 ();
 sg13g2_fill_2 FILLER_4_1329 ();
 sg13g2_fill_2 FILLER_4_1335 ();
 sg13g2_fill_1 FILLER_4_1337 ();
 sg13g2_fill_1 FILLER_4_1343 ();
 sg13g2_fill_2 FILLER_4_1367 ();
 sg13g2_fill_2 FILLER_4_1377 ();
 sg13g2_fill_1 FILLER_4_1379 ();
 sg13g2_fill_2 FILLER_4_1390 ();
 sg13g2_fill_2 FILLER_4_1400 ();
 sg13g2_fill_1 FILLER_4_1402 ();
 sg13g2_fill_2 FILLER_4_1408 ();
 sg13g2_fill_1 FILLER_4_1419 ();
 sg13g2_fill_2 FILLER_4_1477 ();
 sg13g2_fill_1 FILLER_4_1479 ();
 sg13g2_fill_1 FILLER_4_1499 ();
 sg13g2_fill_2 FILLER_4_1534 ();
 sg13g2_fill_2 FILLER_4_1577 ();
 sg13g2_fill_2 FILLER_4_1605 ();
 sg13g2_fill_1 FILLER_4_1625 ();
 sg13g2_fill_1 FILLER_4_1636 ();
 sg13g2_fill_1 FILLER_4_1703 ();
 sg13g2_fill_2 FILLER_4_1811 ();
 sg13g2_fill_2 FILLER_4_1823 ();
 sg13g2_fill_1 FILLER_4_1825 ();
 sg13g2_fill_2 FILLER_4_1990 ();
 sg13g2_fill_2 FILLER_4_2050 ();
 sg13g2_fill_1 FILLER_4_2052 ();
 sg13g2_fill_2 FILLER_4_2068 ();
 sg13g2_fill_1 FILLER_4_2100 ();
 sg13g2_fill_2 FILLER_4_2111 ();
 sg13g2_fill_2 FILLER_4_2123 ();
 sg13g2_fill_2 FILLER_4_2139 ();
 sg13g2_fill_1 FILLER_4_2164 ();
 sg13g2_fill_2 FILLER_4_2190 ();
 sg13g2_fill_2 FILLER_4_2248 ();
 sg13g2_fill_1 FILLER_4_2286 ();
 sg13g2_fill_2 FILLER_4_2382 ();
 sg13g2_fill_2 FILLER_4_2429 ();
 sg13g2_fill_2 FILLER_4_2457 ();
 sg13g2_fill_1 FILLER_4_2459 ();
 sg13g2_fill_2 FILLER_4_2469 ();
 sg13g2_fill_1 FILLER_4_2471 ();
 sg13g2_fill_2 FILLER_4_2487 ();
 sg13g2_fill_1 FILLER_4_2489 ();
 sg13g2_fill_2 FILLER_4_2503 ();
 sg13g2_fill_1 FILLER_4_2505 ();
 sg13g2_fill_2 FILLER_4_2562 ();
 sg13g2_decap_8 FILLER_4_2611 ();
 sg13g2_decap_8 FILLER_4_2618 ();
 sg13g2_decap_8 FILLER_4_2625 ();
 sg13g2_decap_8 FILLER_4_2632 ();
 sg13g2_decap_8 FILLER_4_2639 ();
 sg13g2_decap_8 FILLER_4_2646 ();
 sg13g2_decap_8 FILLER_4_2653 ();
 sg13g2_decap_8 FILLER_4_2660 ();
 sg13g2_decap_8 FILLER_4_2667 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_fill_2 FILLER_5_240 ();
 sg13g2_fill_1 FILLER_5_242 ();
 sg13g2_fill_1 FILLER_5_249 ();
 sg13g2_fill_2 FILLER_5_279 ();
 sg13g2_fill_1 FILLER_5_281 ();
 sg13g2_fill_1 FILLER_5_317 ();
 sg13g2_fill_2 FILLER_5_363 ();
 sg13g2_fill_1 FILLER_5_365 ();
 sg13g2_fill_2 FILLER_5_418 ();
 sg13g2_fill_2 FILLER_5_457 ();
 sg13g2_fill_2 FILLER_5_475 ();
 sg13g2_fill_2 FILLER_5_518 ();
 sg13g2_fill_1 FILLER_5_520 ();
 sg13g2_fill_2 FILLER_5_556 ();
 sg13g2_fill_2 FILLER_5_608 ();
 sg13g2_fill_1 FILLER_5_654 ();
 sg13g2_fill_2 FILLER_5_696 ();
 sg13g2_fill_2 FILLER_5_812 ();
 sg13g2_fill_1 FILLER_5_814 ();
 sg13g2_fill_2 FILLER_5_891 ();
 sg13g2_fill_2 FILLER_5_903 ();
 sg13g2_fill_1 FILLER_5_905 ();
 sg13g2_fill_1 FILLER_5_934 ();
 sg13g2_fill_2 FILLER_5_980 ();
 sg13g2_fill_1 FILLER_5_982 ();
 sg13g2_fill_1 FILLER_5_992 ();
 sg13g2_fill_2 FILLER_5_997 ();
 sg13g2_fill_1 FILLER_5_999 ();
 sg13g2_fill_2 FILLER_5_1012 ();
 sg13g2_fill_1 FILLER_5_1058 ();
 sg13g2_fill_1 FILLER_5_1152 ();
 sg13g2_fill_1 FILLER_5_1197 ();
 sg13g2_fill_2 FILLER_5_1236 ();
 sg13g2_fill_1 FILLER_5_1275 ();
 sg13g2_fill_1 FILLER_5_1293 ();
 sg13g2_fill_2 FILLER_5_1306 ();
 sg13g2_fill_1 FILLER_5_1308 ();
 sg13g2_fill_1 FILLER_5_1317 ();
 sg13g2_fill_2 FILLER_5_1374 ();
 sg13g2_decap_4 FILLER_5_1385 ();
 sg13g2_fill_2 FILLER_5_1401 ();
 sg13g2_fill_2 FILLER_5_1434 ();
 sg13g2_fill_2 FILLER_5_1515 ();
 sg13g2_fill_1 FILLER_5_1546 ();
 sg13g2_fill_2 FILLER_5_1663 ();
 sg13g2_fill_1 FILLER_5_1705 ();
 sg13g2_fill_2 FILLER_5_1740 ();
 sg13g2_fill_1 FILLER_5_1742 ();
 sg13g2_fill_2 FILLER_5_1785 ();
 sg13g2_fill_1 FILLER_5_1787 ();
 sg13g2_fill_2 FILLER_5_1890 ();
 sg13g2_fill_1 FILLER_5_1892 ();
 sg13g2_fill_1 FILLER_5_1944 ();
 sg13g2_fill_1 FILLER_5_2010 ();
 sg13g2_fill_1 FILLER_5_2087 ();
 sg13g2_fill_2 FILLER_5_2114 ();
 sg13g2_fill_1 FILLER_5_2116 ();
 sg13g2_fill_2 FILLER_5_2212 ();
 sg13g2_fill_2 FILLER_5_2294 ();
 sg13g2_fill_1 FILLER_5_2296 ();
 sg13g2_fill_1 FILLER_5_2307 ();
 sg13g2_fill_1 FILLER_5_2351 ();
 sg13g2_fill_2 FILLER_5_2378 ();
 sg13g2_fill_1 FILLER_5_2380 ();
 sg13g2_fill_1 FILLER_5_2422 ();
 sg13g2_fill_2 FILLER_5_2596 ();
 sg13g2_decap_8 FILLER_5_2611 ();
 sg13g2_decap_8 FILLER_5_2618 ();
 sg13g2_decap_8 FILLER_5_2625 ();
 sg13g2_decap_8 FILLER_5_2632 ();
 sg13g2_decap_8 FILLER_5_2639 ();
 sg13g2_decap_8 FILLER_5_2646 ();
 sg13g2_decap_8 FILLER_5_2653 ();
 sg13g2_decap_8 FILLER_5_2660 ();
 sg13g2_decap_8 FILLER_5_2667 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_fill_2 FILLER_6_112 ();
 sg13g2_fill_1 FILLER_6_114 ();
 sg13g2_fill_1 FILLER_6_174 ();
 sg13g2_fill_1 FILLER_6_191 ();
 sg13g2_fill_1 FILLER_6_198 ();
 sg13g2_fill_1 FILLER_6_273 ();
 sg13g2_fill_1 FILLER_6_290 ();
 sg13g2_fill_2 FILLER_6_329 ();
 sg13g2_fill_2 FILLER_6_394 ();
 sg13g2_fill_2 FILLER_6_482 ();
 sg13g2_fill_2 FILLER_6_545 ();
 sg13g2_fill_1 FILLER_6_547 ();
 sg13g2_fill_2 FILLER_6_567 ();
 sg13g2_fill_1 FILLER_6_569 ();
 sg13g2_fill_2 FILLER_6_584 ();
 sg13g2_fill_1 FILLER_6_604 ();
 sg13g2_fill_1 FILLER_6_610 ();
 sg13g2_fill_2 FILLER_6_635 ();
 sg13g2_fill_2 FILLER_6_673 ();
 sg13g2_fill_1 FILLER_6_675 ();
 sg13g2_fill_2 FILLER_6_712 ();
 sg13g2_fill_1 FILLER_6_749 ();
 sg13g2_fill_2 FILLER_6_789 ();
 sg13g2_fill_1 FILLER_6_898 ();
 sg13g2_fill_1 FILLER_6_924 ();
 sg13g2_fill_2 FILLER_6_964 ();
 sg13g2_fill_2 FILLER_6_1051 ();
 sg13g2_fill_1 FILLER_6_1053 ();
 sg13g2_fill_1 FILLER_6_1113 ();
 sg13g2_fill_1 FILLER_6_1127 ();
 sg13g2_fill_1 FILLER_6_1147 ();
 sg13g2_fill_2 FILLER_6_1296 ();
 sg13g2_fill_1 FILLER_6_1304 ();
 sg13g2_fill_2 FILLER_6_1314 ();
 sg13g2_fill_1 FILLER_6_1383 ();
 sg13g2_decap_4 FILLER_6_1388 ();
 sg13g2_decap_4 FILLER_6_1395 ();
 sg13g2_fill_1 FILLER_6_1399 ();
 sg13g2_fill_2 FILLER_6_1413 ();
 sg13g2_fill_2 FILLER_6_1444 ();
 sg13g2_fill_1 FILLER_6_1446 ();
 sg13g2_fill_1 FILLER_6_1452 ();
 sg13g2_fill_2 FILLER_6_1500 ();
 sg13g2_fill_2 FILLER_6_1531 ();
 sg13g2_fill_2 FILLER_6_1570 ();
 sg13g2_fill_2 FILLER_6_1599 ();
 sg13g2_fill_1 FILLER_6_1608 ();
 sg13g2_fill_1 FILLER_6_1677 ();
 sg13g2_fill_2 FILLER_6_1713 ();
 sg13g2_fill_2 FILLER_6_1802 ();
 sg13g2_fill_1 FILLER_6_1804 ();
 sg13g2_fill_2 FILLER_6_1818 ();
 sg13g2_fill_2 FILLER_6_2038 ();
 sg13g2_fill_2 FILLER_6_2085 ();
 sg13g2_fill_1 FILLER_6_2087 ();
 sg13g2_fill_2 FILLER_6_2143 ();
 sg13g2_fill_2 FILLER_6_2154 ();
 sg13g2_fill_1 FILLER_6_2176 ();
 sg13g2_fill_2 FILLER_6_2285 ();
 sg13g2_fill_2 FILLER_6_2327 ();
 sg13g2_fill_2 FILLER_6_2350 ();
 sg13g2_fill_1 FILLER_6_2378 ();
 sg13g2_fill_1 FILLER_6_2409 ();
 sg13g2_fill_1 FILLER_6_2443 ();
 sg13g2_fill_2 FILLER_6_2458 ();
 sg13g2_fill_1 FILLER_6_2460 ();
 sg13g2_fill_2 FILLER_6_2521 ();
 sg13g2_fill_1 FILLER_6_2523 ();
 sg13g2_fill_1 FILLER_6_2554 ();
 sg13g2_fill_2 FILLER_6_2575 ();
 sg13g2_fill_1 FILLER_6_2577 ();
 sg13g2_decap_8 FILLER_6_2606 ();
 sg13g2_decap_8 FILLER_6_2613 ();
 sg13g2_decap_8 FILLER_6_2620 ();
 sg13g2_decap_8 FILLER_6_2627 ();
 sg13g2_decap_8 FILLER_6_2634 ();
 sg13g2_decap_8 FILLER_6_2641 ();
 sg13g2_decap_8 FILLER_6_2648 ();
 sg13g2_decap_8 FILLER_6_2655 ();
 sg13g2_decap_8 FILLER_6_2662 ();
 sg13g2_decap_4 FILLER_6_2669 ();
 sg13g2_fill_1 FILLER_6_2673 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_fill_2 FILLER_7_119 ();
 sg13g2_fill_1 FILLER_7_121 ();
 sg13g2_fill_1 FILLER_7_148 ();
 sg13g2_fill_1 FILLER_7_231 ();
 sg13g2_fill_1 FILLER_7_273 ();
 sg13g2_fill_1 FILLER_7_284 ();
 sg13g2_fill_1 FILLER_7_316 ();
 sg13g2_fill_1 FILLER_7_406 ();
 sg13g2_fill_2 FILLER_7_451 ();
 sg13g2_fill_1 FILLER_7_517 ();
 sg13g2_fill_1 FILLER_7_541 ();
 sg13g2_fill_1 FILLER_7_548 ();
 sg13g2_fill_1 FILLER_7_651 ();
 sg13g2_fill_1 FILLER_7_672 ();
 sg13g2_fill_2 FILLER_7_729 ();
 sg13g2_fill_1 FILLER_7_750 ();
 sg13g2_fill_1 FILLER_7_761 ();
 sg13g2_fill_1 FILLER_7_779 ();
 sg13g2_fill_2 FILLER_7_936 ();
 sg13g2_fill_2 FILLER_7_953 ();
 sg13g2_fill_2 FILLER_7_966 ();
 sg13g2_fill_1 FILLER_7_979 ();
 sg13g2_fill_2 FILLER_7_989 ();
 sg13g2_fill_1 FILLER_7_991 ();
 sg13g2_fill_2 FILLER_7_1057 ();
 sg13g2_fill_2 FILLER_7_1160 ();
 sg13g2_fill_2 FILLER_7_1190 ();
 sg13g2_fill_1 FILLER_7_1201 ();
 sg13g2_fill_2 FILLER_7_1266 ();
 sg13g2_fill_2 FILLER_7_1286 ();
 sg13g2_fill_1 FILLER_7_1328 ();
 sg13g2_fill_2 FILLER_7_1353 ();
 sg13g2_fill_1 FILLER_7_1355 ();
 sg13g2_fill_2 FILLER_7_1369 ();
 sg13g2_fill_1 FILLER_7_1371 ();
 sg13g2_fill_2 FILLER_7_1423 ();
 sg13g2_fill_1 FILLER_7_1425 ();
 sg13g2_decap_8 FILLER_7_1441 ();
 sg13g2_fill_1 FILLER_7_1513 ();
 sg13g2_fill_1 FILLER_7_1570 ();
 sg13g2_fill_2 FILLER_7_1703 ();
 sg13g2_fill_2 FILLER_7_1748 ();
 sg13g2_fill_1 FILLER_7_1750 ();
 sg13g2_fill_2 FILLER_7_1764 ();
 sg13g2_fill_2 FILLER_7_1806 ();
 sg13g2_fill_1 FILLER_7_1808 ();
 sg13g2_fill_2 FILLER_7_1853 ();
 sg13g2_fill_1 FILLER_7_1868 ();
 sg13g2_fill_2 FILLER_7_1890 ();
 sg13g2_fill_2 FILLER_7_1917 ();
 sg13g2_fill_2 FILLER_7_1934 ();
 sg13g2_fill_1 FILLER_7_1936 ();
 sg13g2_fill_2 FILLER_7_1947 ();
 sg13g2_fill_2 FILLER_7_2011 ();
 sg13g2_fill_1 FILLER_7_2062 ();
 sg13g2_fill_2 FILLER_7_2116 ();
 sg13g2_fill_1 FILLER_7_2313 ();
 sg13g2_fill_1 FILLER_7_2379 ();
 sg13g2_fill_2 FILLER_7_2480 ();
 sg13g2_fill_1 FILLER_7_2482 ();
 sg13g2_fill_1 FILLER_7_2508 ();
 sg13g2_fill_1 FILLER_7_2539 ();
 sg13g2_fill_2 FILLER_7_2570 ();
 sg13g2_fill_1 FILLER_7_2572 ();
 sg13g2_decap_8 FILLER_7_2625 ();
 sg13g2_decap_8 FILLER_7_2632 ();
 sg13g2_decap_8 FILLER_7_2639 ();
 sg13g2_decap_8 FILLER_7_2646 ();
 sg13g2_decap_8 FILLER_7_2653 ();
 sg13g2_decap_8 FILLER_7_2660 ();
 sg13g2_decap_8 FILLER_7_2667 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_fill_2 FILLER_8_177 ();
 sg13g2_fill_2 FILLER_8_189 ();
 sg13g2_fill_2 FILLER_8_322 ();
 sg13g2_fill_1 FILLER_8_324 ();
 sg13g2_fill_1 FILLER_8_342 ();
 sg13g2_fill_1 FILLER_8_491 ();
 sg13g2_fill_2 FILLER_8_509 ();
 sg13g2_fill_1 FILLER_8_534 ();
 sg13g2_fill_1 FILLER_8_541 ();
 sg13g2_fill_2 FILLER_8_562 ();
 sg13g2_fill_2 FILLER_8_582 ();
 sg13g2_fill_1 FILLER_8_584 ();
 sg13g2_fill_1 FILLER_8_648 ();
 sg13g2_fill_2 FILLER_8_675 ();
 sg13g2_fill_2 FILLER_8_703 ();
 sg13g2_fill_1 FILLER_8_705 ();
 sg13g2_fill_1 FILLER_8_715 ();
 sg13g2_fill_2 FILLER_8_778 ();
 sg13g2_fill_1 FILLER_8_780 ();
 sg13g2_fill_2 FILLER_8_794 ();
 sg13g2_fill_2 FILLER_8_812 ();
 sg13g2_fill_1 FILLER_8_814 ();
 sg13g2_fill_2 FILLER_8_847 ();
 sg13g2_fill_1 FILLER_8_849 ();
 sg13g2_fill_2 FILLER_8_976 ();
 sg13g2_fill_1 FILLER_8_1040 ();
 sg13g2_fill_2 FILLER_8_1050 ();
 sg13g2_fill_1 FILLER_8_1052 ();
 sg13g2_fill_2 FILLER_8_1100 ();
 sg13g2_fill_1 FILLER_8_1102 ();
 sg13g2_fill_1 FILLER_8_1119 ();
 sg13g2_fill_1 FILLER_8_1156 ();
 sg13g2_fill_2 FILLER_8_1248 ();
 sg13g2_fill_2 FILLER_8_1260 ();
 sg13g2_fill_1 FILLER_8_1262 ();
 sg13g2_fill_2 FILLER_8_1303 ();
 sg13g2_fill_1 FILLER_8_1305 ();
 sg13g2_fill_2 FILLER_8_1315 ();
 sg13g2_fill_1 FILLER_8_1317 ();
 sg13g2_fill_1 FILLER_8_1344 ();
 sg13g2_fill_1 FILLER_8_1383 ();
 sg13g2_fill_2 FILLER_8_1401 ();
 sg13g2_fill_1 FILLER_8_1403 ();
 sg13g2_fill_1 FILLER_8_1457 ();
 sg13g2_fill_2 FILLER_8_1462 ();
 sg13g2_fill_1 FILLER_8_1464 ();
 sg13g2_fill_2 FILLER_8_1479 ();
 sg13g2_decap_8 FILLER_8_1485 ();
 sg13g2_decap_4 FILLER_8_1492 ();
 sg13g2_fill_2 FILLER_8_1509 ();
 sg13g2_fill_1 FILLER_8_1511 ();
 sg13g2_fill_1 FILLER_8_1533 ();
 sg13g2_fill_2 FILLER_8_1591 ();
 sg13g2_fill_1 FILLER_8_1593 ();
 sg13g2_decap_4 FILLER_8_1614 ();
 sg13g2_fill_2 FILLER_8_1618 ();
 sg13g2_fill_2 FILLER_8_1628 ();
 sg13g2_fill_2 FILLER_8_1657 ();
 sg13g2_fill_1 FILLER_8_1659 ();
 sg13g2_fill_2 FILLER_8_1728 ();
 sg13g2_fill_1 FILLER_8_1730 ();
 sg13g2_fill_2 FILLER_8_1803 ();
 sg13g2_fill_1 FILLER_8_1805 ();
 sg13g2_fill_1 FILLER_8_1834 ();
 sg13g2_fill_1 FILLER_8_1871 ();
 sg13g2_fill_2 FILLER_8_1948 ();
 sg13g2_fill_1 FILLER_8_1950 ();
 sg13g2_fill_2 FILLER_8_2005 ();
 sg13g2_fill_2 FILLER_8_2037 ();
 sg13g2_fill_1 FILLER_8_2105 ();
 sg13g2_fill_2 FILLER_8_2200 ();
 sg13g2_fill_2 FILLER_8_2382 ();
 sg13g2_fill_1 FILLER_8_2384 ();
 sg13g2_fill_2 FILLER_8_2429 ();
 sg13g2_fill_1 FILLER_8_2431 ();
 sg13g2_decap_8 FILLER_8_2624 ();
 sg13g2_decap_8 FILLER_8_2631 ();
 sg13g2_decap_8 FILLER_8_2638 ();
 sg13g2_decap_8 FILLER_8_2645 ();
 sg13g2_decap_8 FILLER_8_2652 ();
 sg13g2_decap_8 FILLER_8_2659 ();
 sg13g2_decap_8 FILLER_8_2666 ();
 sg13g2_fill_1 FILLER_8_2673 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_fill_2 FILLER_9_161 ();
 sg13g2_fill_2 FILLER_9_178 ();
 sg13g2_fill_2 FILLER_9_215 ();
 sg13g2_fill_1 FILLER_9_217 ();
 sg13g2_fill_2 FILLER_9_243 ();
 sg13g2_fill_1 FILLER_9_245 ();
 sg13g2_fill_2 FILLER_9_315 ();
 sg13g2_fill_1 FILLER_9_317 ();
 sg13g2_fill_1 FILLER_9_354 ();
 sg13g2_fill_2 FILLER_9_385 ();
 sg13g2_fill_1 FILLER_9_397 ();
 sg13g2_fill_1 FILLER_9_417 ();
 sg13g2_fill_1 FILLER_9_438 ();
 sg13g2_fill_1 FILLER_9_448 ();
 sg13g2_fill_1 FILLER_9_486 ();
 sg13g2_fill_2 FILLER_9_653 ();
 sg13g2_fill_2 FILLER_9_660 ();
 sg13g2_fill_1 FILLER_9_704 ();
 sg13g2_fill_2 FILLER_9_733 ();
 sg13g2_fill_1 FILLER_9_735 ();
 sg13g2_fill_1 FILLER_9_755 ();
 sg13g2_fill_1 FILLER_9_790 ();
 sg13g2_fill_1 FILLER_9_825 ();
 sg13g2_fill_1 FILLER_9_924 ();
 sg13g2_fill_1 FILLER_9_1028 ();
 sg13g2_fill_2 FILLER_9_1084 ();
 sg13g2_fill_1 FILLER_9_1086 ();
 sg13g2_fill_1 FILLER_9_1146 ();
 sg13g2_fill_1 FILLER_9_1219 ();
 sg13g2_fill_2 FILLER_9_1272 ();
 sg13g2_fill_1 FILLER_9_1287 ();
 sg13g2_fill_1 FILLER_9_1318 ();
 sg13g2_fill_2 FILLER_9_1324 ();
 sg13g2_fill_1 FILLER_9_1326 ();
 sg13g2_fill_2 FILLER_9_1337 ();
 sg13g2_fill_2 FILLER_9_1352 ();
 sg13g2_fill_1 FILLER_9_1354 ();
 sg13g2_fill_2 FILLER_9_1364 ();
 sg13g2_fill_1 FILLER_9_1366 ();
 sg13g2_fill_1 FILLER_9_1406 ();
 sg13g2_fill_1 FILLER_9_1439 ();
 sg13g2_decap_8 FILLER_9_1453 ();
 sg13g2_decap_4 FILLER_9_1460 ();
 sg13g2_decap_4 FILLER_9_1479 ();
 sg13g2_fill_1 FILLER_9_1483 ();
 sg13g2_fill_2 FILLER_9_1500 ();
 sg13g2_fill_2 FILLER_9_1507 ();
 sg13g2_fill_2 FILLER_9_1526 ();
 sg13g2_fill_2 FILLER_9_1540 ();
 sg13g2_fill_1 FILLER_9_1542 ();
 sg13g2_fill_2 FILLER_9_1571 ();
 sg13g2_fill_1 FILLER_9_1573 ();
 sg13g2_fill_1 FILLER_9_1604 ();
 sg13g2_fill_1 FILLER_9_1643 ();
 sg13g2_fill_1 FILLER_9_1652 ();
 sg13g2_fill_2 FILLER_9_1674 ();
 sg13g2_fill_1 FILLER_9_1676 ();
 sg13g2_fill_2 FILLER_9_1775 ();
 sg13g2_fill_1 FILLER_9_1777 ();
 sg13g2_fill_1 FILLER_9_1800 ();
 sg13g2_fill_2 FILLER_9_1814 ();
 sg13g2_fill_1 FILLER_9_1922 ();
 sg13g2_fill_2 FILLER_9_1932 ();
 sg13g2_fill_2 FILLER_9_2019 ();
 sg13g2_fill_1 FILLER_9_2021 ();
 sg13g2_fill_2 FILLER_9_2048 ();
 sg13g2_fill_2 FILLER_9_2064 ();
 sg13g2_fill_2 FILLER_9_2080 ();
 sg13g2_fill_1 FILLER_9_2108 ();
 sg13g2_fill_2 FILLER_9_2133 ();
 sg13g2_fill_2 FILLER_9_2171 ();
 sg13g2_fill_1 FILLER_9_2173 ();
 sg13g2_fill_2 FILLER_9_2218 ();
 sg13g2_fill_1 FILLER_9_2220 ();
 sg13g2_fill_2 FILLER_9_2292 ();
 sg13g2_fill_1 FILLER_9_2319 ();
 sg13g2_fill_2 FILLER_9_2346 ();
 sg13g2_fill_2 FILLER_9_2386 ();
 sg13g2_fill_2 FILLER_9_2402 ();
 sg13g2_fill_2 FILLER_9_2413 ();
 sg13g2_fill_1 FILLER_9_2415 ();
 sg13g2_fill_2 FILLER_9_2491 ();
 sg13g2_fill_1 FILLER_9_2493 ();
 sg13g2_fill_2 FILLER_9_2580 ();
 sg13g2_fill_1 FILLER_9_2592 ();
 sg13g2_decap_8 FILLER_9_2619 ();
 sg13g2_decap_8 FILLER_9_2626 ();
 sg13g2_decap_8 FILLER_9_2633 ();
 sg13g2_decap_8 FILLER_9_2640 ();
 sg13g2_decap_8 FILLER_9_2647 ();
 sg13g2_decap_8 FILLER_9_2654 ();
 sg13g2_decap_8 FILLER_9_2661 ();
 sg13g2_decap_4 FILLER_9_2668 ();
 sg13g2_fill_2 FILLER_9_2672 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_fill_1 FILLER_10_98 ();
 sg13g2_fill_2 FILLER_10_165 ();
 sg13g2_fill_2 FILLER_10_191 ();
 sg13g2_fill_1 FILLER_10_193 ();
 sg13g2_fill_2 FILLER_10_211 ();
 sg13g2_fill_2 FILLER_10_257 ();
 sg13g2_fill_2 FILLER_10_445 ();
 sg13g2_fill_1 FILLER_10_447 ();
 sg13g2_fill_2 FILLER_10_508 ();
 sg13g2_fill_1 FILLER_10_510 ();
 sg13g2_fill_1 FILLER_10_552 ();
 sg13g2_fill_1 FILLER_10_564 ();
 sg13g2_fill_1 FILLER_10_586 ();
 sg13g2_fill_1 FILLER_10_600 ();
 sg13g2_fill_1 FILLER_10_606 ();
 sg13g2_fill_1 FILLER_10_660 ();
 sg13g2_fill_1 FILLER_10_722 ();
 sg13g2_fill_2 FILLER_10_728 ();
 sg13g2_fill_2 FILLER_10_898 ();
 sg13g2_fill_2 FILLER_10_946 ();
 sg13g2_fill_1 FILLER_10_948 ();
 sg13g2_fill_1 FILLER_10_1014 ();
 sg13g2_fill_2 FILLER_10_1095 ();
 sg13g2_fill_2 FILLER_10_1105 ();
 sg13g2_fill_2 FILLER_10_1136 ();
 sg13g2_fill_1 FILLER_10_1138 ();
 sg13g2_fill_2 FILLER_10_1184 ();
 sg13g2_fill_2 FILLER_10_1248 ();
 sg13g2_fill_1 FILLER_10_1278 ();
 sg13g2_fill_2 FILLER_10_1287 ();
 sg13g2_fill_1 FILLER_10_1289 ();
 sg13g2_fill_2 FILLER_10_1300 ();
 sg13g2_fill_1 FILLER_10_1302 ();
 sg13g2_fill_2 FILLER_10_1308 ();
 sg13g2_fill_1 FILLER_10_1310 ();
 sg13g2_fill_2 FILLER_10_1323 ();
 sg13g2_fill_1 FILLER_10_1346 ();
 sg13g2_fill_2 FILLER_10_1357 ();
 sg13g2_fill_2 FILLER_10_1377 ();
 sg13g2_fill_1 FILLER_10_1379 ();
 sg13g2_fill_2 FILLER_10_1393 ();
 sg13g2_fill_1 FILLER_10_1395 ();
 sg13g2_fill_2 FILLER_10_1404 ();
 sg13g2_fill_1 FILLER_10_1406 ();
 sg13g2_decap_4 FILLER_10_1427 ();
 sg13g2_fill_2 FILLER_10_1431 ();
 sg13g2_fill_1 FILLER_10_1442 ();
 sg13g2_fill_1 FILLER_10_1486 ();
 sg13g2_fill_2 FILLER_10_1546 ();
 sg13g2_fill_1 FILLER_10_1574 ();
 sg13g2_fill_2 FILLER_10_1583 ();
 sg13g2_fill_2 FILLER_10_1601 ();
 sg13g2_fill_1 FILLER_10_1603 ();
 sg13g2_fill_2 FILLER_10_1654 ();
 sg13g2_fill_2 FILLER_10_1666 ();
 sg13g2_fill_1 FILLER_10_1702 ();
 sg13g2_fill_2 FILLER_10_1724 ();
 sg13g2_fill_1 FILLER_10_1780 ();
 sg13g2_fill_1 FILLER_10_1816 ();
 sg13g2_fill_1 FILLER_10_1878 ();
 sg13g2_fill_1 FILLER_10_1898 ();
 sg13g2_fill_1 FILLER_10_1939 ();
 sg13g2_fill_2 FILLER_10_2010 ();
 sg13g2_fill_1 FILLER_10_2026 ();
 sg13g2_fill_2 FILLER_10_2053 ();
 sg13g2_fill_1 FILLER_10_2237 ();
 sg13g2_fill_1 FILLER_10_2266 ();
 sg13g2_fill_1 FILLER_10_2276 ();
 sg13g2_fill_1 FILLER_10_2303 ();
 sg13g2_fill_1 FILLER_10_2336 ();
 sg13g2_fill_2 FILLER_10_2424 ();
 sg13g2_fill_1 FILLER_10_2426 ();
 sg13g2_fill_2 FILLER_10_2462 ();
 sg13g2_fill_1 FILLER_10_2464 ();
 sg13g2_fill_2 FILLER_10_2496 ();
 sg13g2_fill_1 FILLER_10_2498 ();
 sg13g2_fill_1 FILLER_10_2554 ();
 sg13g2_fill_2 FILLER_10_2565 ();
 sg13g2_decap_8 FILLER_10_2623 ();
 sg13g2_decap_8 FILLER_10_2630 ();
 sg13g2_decap_8 FILLER_10_2637 ();
 sg13g2_decap_8 FILLER_10_2644 ();
 sg13g2_decap_8 FILLER_10_2651 ();
 sg13g2_decap_8 FILLER_10_2658 ();
 sg13g2_decap_8 FILLER_10_2665 ();
 sg13g2_fill_2 FILLER_10_2672 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_fill_2 FILLER_11_84 ();
 sg13g2_fill_1 FILLER_11_158 ();
 sg13g2_fill_1 FILLER_11_175 ();
 sg13g2_fill_1 FILLER_11_239 ();
 sg13g2_fill_2 FILLER_11_270 ();
 sg13g2_fill_1 FILLER_11_272 ();
 sg13g2_fill_2 FILLER_11_313 ();
 sg13g2_fill_1 FILLER_11_315 ();
 sg13g2_fill_1 FILLER_11_365 ();
 sg13g2_fill_2 FILLER_11_398 ();
 sg13g2_fill_2 FILLER_11_458 ();
 sg13g2_fill_1 FILLER_11_460 ();
 sg13g2_fill_2 FILLER_11_487 ();
 sg13g2_fill_1 FILLER_11_511 ();
 sg13g2_fill_1 FILLER_11_527 ();
 sg13g2_fill_1 FILLER_11_577 ();
 sg13g2_fill_2 FILLER_11_622 ();
 sg13g2_fill_1 FILLER_11_624 ();
 sg13g2_fill_2 FILLER_11_634 ();
 sg13g2_fill_2 FILLER_11_677 ();
 sg13g2_fill_2 FILLER_11_703 ();
 sg13g2_fill_1 FILLER_11_705 ();
 sg13g2_fill_2 FILLER_11_730 ();
 sg13g2_fill_1 FILLER_11_732 ();
 sg13g2_fill_1 FILLER_11_812 ();
 sg13g2_fill_1 FILLER_11_830 ();
 sg13g2_fill_2 FILLER_11_871 ();
 sg13g2_fill_1 FILLER_11_919 ();
 sg13g2_fill_2 FILLER_11_934 ();
 sg13g2_fill_1 FILLER_11_962 ();
 sg13g2_fill_2 FILLER_11_1062 ();
 sg13g2_fill_2 FILLER_11_1073 ();
 sg13g2_fill_2 FILLER_11_1101 ();
 sg13g2_fill_1 FILLER_11_1103 ();
 sg13g2_fill_2 FILLER_11_1140 ();
 sg13g2_fill_2 FILLER_11_1269 ();
 sg13g2_fill_1 FILLER_11_1271 ();
 sg13g2_fill_2 FILLER_11_1293 ();
 sg13g2_fill_1 FILLER_11_1295 ();
 sg13g2_fill_2 FILLER_11_1345 ();
 sg13g2_fill_2 FILLER_11_1412 ();
 sg13g2_fill_2 FILLER_11_1419 ();
 sg13g2_fill_2 FILLER_11_1439 ();
 sg13g2_decap_8 FILLER_11_1476 ();
 sg13g2_decap_4 FILLER_11_1483 ();
 sg13g2_decap_4 FILLER_11_1516 ();
 sg13g2_fill_2 FILLER_11_1520 ();
 sg13g2_decap_4 FILLER_11_1535 ();
 sg13g2_fill_1 FILLER_11_1544 ();
 sg13g2_fill_2 FILLER_11_1553 ();
 sg13g2_fill_1 FILLER_11_1555 ();
 sg13g2_fill_2 FILLER_11_1586 ();
 sg13g2_fill_2 FILLER_11_1606 ();
 sg13g2_fill_1 FILLER_11_1608 ();
 sg13g2_fill_2 FILLER_11_1619 ();
 sg13g2_fill_1 FILLER_11_1621 ();
 sg13g2_fill_1 FILLER_11_1650 ();
 sg13g2_decap_4 FILLER_11_1677 ();
 sg13g2_fill_1 FILLER_11_1685 ();
 sg13g2_fill_1 FILLER_11_1699 ();
 sg13g2_fill_2 FILLER_11_1794 ();
 sg13g2_fill_2 FILLER_11_1830 ();
 sg13g2_fill_1 FILLER_11_1832 ();
 sg13g2_fill_2 FILLER_11_1907 ();
 sg13g2_fill_2 FILLER_11_1925 ();
 sg13g2_fill_1 FILLER_11_1927 ();
 sg13g2_fill_2 FILLER_11_1959 ();
 sg13g2_fill_1 FILLER_11_1974 ();
 sg13g2_fill_2 FILLER_11_2004 ();
 sg13g2_fill_1 FILLER_11_2006 ();
 sg13g2_fill_2 FILLER_11_2060 ();
 sg13g2_fill_1 FILLER_11_2062 ();
 sg13g2_fill_1 FILLER_11_2100 ();
 sg13g2_fill_2 FILLER_11_2155 ();
 sg13g2_fill_1 FILLER_11_2281 ();
 sg13g2_fill_1 FILLER_11_2292 ();
 sg13g2_fill_1 FILLER_11_2303 ();
 sg13g2_fill_1 FILLER_11_2336 ();
 sg13g2_fill_2 FILLER_11_2373 ();
 sg13g2_fill_1 FILLER_11_2375 ();
 sg13g2_fill_2 FILLER_11_2418 ();
 sg13g2_fill_2 FILLER_11_2439 ();
 sg13g2_fill_1 FILLER_11_2538 ();
 sg13g2_fill_2 FILLER_11_2565 ();
 sg13g2_fill_1 FILLER_11_2567 ();
 sg13g2_fill_1 FILLER_11_2591 ();
 sg13g2_decap_8 FILLER_11_2626 ();
 sg13g2_decap_8 FILLER_11_2633 ();
 sg13g2_decap_8 FILLER_11_2640 ();
 sg13g2_decap_8 FILLER_11_2647 ();
 sg13g2_decap_8 FILLER_11_2654 ();
 sg13g2_decap_8 FILLER_11_2661 ();
 sg13g2_decap_4 FILLER_11_2668 ();
 sg13g2_fill_2 FILLER_11_2672 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_4 FILLER_12_70 ();
 sg13g2_fill_1 FILLER_12_128 ();
 sg13g2_fill_1 FILLER_12_167 ();
 sg13g2_fill_2 FILLER_12_207 ();
 sg13g2_fill_2 FILLER_12_219 ();
 sg13g2_fill_1 FILLER_12_221 ();
 sg13g2_fill_1 FILLER_12_253 ();
 sg13g2_fill_1 FILLER_12_301 ();
 sg13g2_fill_2 FILLER_12_340 ();
 sg13g2_fill_2 FILLER_12_397 ();
 sg13g2_fill_1 FILLER_12_399 ();
 sg13g2_fill_1 FILLER_12_415 ();
 sg13g2_fill_2 FILLER_12_425 ();
 sg13g2_fill_1 FILLER_12_435 ();
 sg13g2_fill_2 FILLER_12_481 ();
 sg13g2_fill_1 FILLER_12_513 ();
 sg13g2_fill_2 FILLER_12_540 ();
 sg13g2_fill_1 FILLER_12_542 ();
 sg13g2_fill_2 FILLER_12_571 ();
 sg13g2_fill_1 FILLER_12_573 ();
 sg13g2_fill_1 FILLER_12_584 ();
 sg13g2_fill_1 FILLER_12_639 ();
 sg13g2_fill_2 FILLER_12_665 ();
 sg13g2_fill_1 FILLER_12_667 ();
 sg13g2_fill_2 FILLER_12_694 ();
 sg13g2_fill_2 FILLER_12_770 ();
 sg13g2_fill_2 FILLER_12_814 ();
 sg13g2_fill_1 FILLER_12_816 ();
 sg13g2_fill_2 FILLER_12_833 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_fill_2 FILLER_12_888 ();
 sg13g2_fill_1 FILLER_12_934 ();
 sg13g2_fill_1 FILLER_12_970 ();
 sg13g2_fill_1 FILLER_12_993 ();
 sg13g2_fill_2 FILLER_12_1013 ();
 sg13g2_fill_1 FILLER_12_1015 ();
 sg13g2_fill_1 FILLER_12_1067 ();
 sg13g2_fill_2 FILLER_12_1101 ();
 sg13g2_fill_1 FILLER_12_1103 ();
 sg13g2_fill_1 FILLER_12_1123 ();
 sg13g2_fill_2 FILLER_12_1152 ();
 sg13g2_fill_1 FILLER_12_1173 ();
 sg13g2_fill_1 FILLER_12_1226 ();
 sg13g2_fill_1 FILLER_12_1241 ();
 sg13g2_fill_1 FILLER_12_1304 ();
 sg13g2_fill_1 FILLER_12_1317 ();
 sg13g2_decap_4 FILLER_12_1322 ();
 sg13g2_fill_2 FILLER_12_1362 ();
 sg13g2_fill_1 FILLER_12_1375 ();
 sg13g2_fill_2 FILLER_12_1408 ();
 sg13g2_fill_2 FILLER_12_1429 ();
 sg13g2_fill_2 FILLER_12_1457 ();
 sg13g2_fill_2 FILLER_12_1510 ();
 sg13g2_fill_2 FILLER_12_1541 ();
 sg13g2_fill_1 FILLER_12_1543 ();
 sg13g2_fill_1 FILLER_12_1565 ();
 sg13g2_fill_1 FILLER_12_1592 ();
 sg13g2_fill_1 FILLER_12_1639 ();
 sg13g2_fill_1 FILLER_12_1647 ();
 sg13g2_fill_1 FILLER_12_1669 ();
 sg13g2_fill_2 FILLER_12_1706 ();
 sg13g2_fill_2 FILLER_12_1760 ();
 sg13g2_fill_1 FILLER_12_1762 ();
 sg13g2_fill_1 FILLER_12_1869 ();
 sg13g2_fill_1 FILLER_12_1880 ();
 sg13g2_fill_2 FILLER_12_1943 ();
 sg13g2_fill_2 FILLER_12_2003 ();
 sg13g2_fill_1 FILLER_12_2005 ();
 sg13g2_fill_1 FILLER_12_2016 ();
 sg13g2_fill_2 FILLER_12_2043 ();
 sg13g2_fill_1 FILLER_12_2045 ();
 sg13g2_fill_2 FILLER_12_2072 ();
 sg13g2_fill_1 FILLER_12_2136 ();
 sg13g2_fill_2 FILLER_12_2257 ();
 sg13g2_fill_1 FILLER_12_2259 ();
 sg13g2_fill_2 FILLER_12_2312 ();
 sg13g2_fill_2 FILLER_12_2323 ();
 sg13g2_fill_1 FILLER_12_2325 ();
 sg13g2_fill_2 FILLER_12_2377 ();
 sg13g2_fill_1 FILLER_12_2477 ();
 sg13g2_fill_2 FILLER_12_2511 ();
 sg13g2_decap_8 FILLER_12_2637 ();
 sg13g2_decap_8 FILLER_12_2644 ();
 sg13g2_decap_8 FILLER_12_2651 ();
 sg13g2_decap_8 FILLER_12_2658 ();
 sg13g2_decap_8 FILLER_12_2665 ();
 sg13g2_fill_2 FILLER_12_2672 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_4 FILLER_13_63 ();
 sg13g2_fill_2 FILLER_13_75 ();
 sg13g2_fill_1 FILLER_13_77 ();
 sg13g2_fill_1 FILLER_13_86 ();
 sg13g2_fill_2 FILLER_13_117 ();
 sg13g2_fill_2 FILLER_13_232 ();
 sg13g2_fill_1 FILLER_13_262 ();
 sg13g2_fill_2 FILLER_13_293 ();
 sg13g2_fill_1 FILLER_13_295 ();
 sg13g2_fill_2 FILLER_13_322 ();
 sg13g2_fill_2 FILLER_13_360 ();
 sg13g2_fill_2 FILLER_13_372 ();
 sg13g2_fill_1 FILLER_13_389 ();
 sg13g2_fill_2 FILLER_13_428 ();
 sg13g2_fill_2 FILLER_13_497 ();
 sg13g2_fill_2 FILLER_13_514 ();
 sg13g2_fill_1 FILLER_13_530 ();
 sg13g2_fill_2 FILLER_13_548 ();
 sg13g2_fill_1 FILLER_13_576 ();
 sg13g2_fill_2 FILLER_13_650 ();
 sg13g2_fill_1 FILLER_13_652 ();
 sg13g2_fill_1 FILLER_13_739 ();
 sg13g2_fill_1 FILLER_13_780 ();
 sg13g2_fill_1 FILLER_13_791 ();
 sg13g2_fill_1 FILLER_13_852 ();
 sg13g2_fill_1 FILLER_13_867 ();
 sg13g2_fill_2 FILLER_13_873 ();
 sg13g2_fill_1 FILLER_13_875 ();
 sg13g2_fill_2 FILLER_13_894 ();
 sg13g2_fill_2 FILLER_13_932 ();
 sg13g2_fill_1 FILLER_13_934 ();
 sg13g2_fill_1 FILLER_13_949 ();
 sg13g2_fill_1 FILLER_13_1009 ();
 sg13g2_fill_2 FILLER_13_1130 ();
 sg13g2_fill_2 FILLER_13_1145 ();
 sg13g2_fill_2 FILLER_13_1189 ();
 sg13g2_fill_1 FILLER_13_1240 ();
 sg13g2_fill_2 FILLER_13_1269 ();
 sg13g2_fill_1 FILLER_13_1271 ();
 sg13g2_fill_2 FILLER_13_1281 ();
 sg13g2_fill_2 FILLER_13_1326 ();
 sg13g2_fill_1 FILLER_13_1349 ();
 sg13g2_fill_2 FILLER_13_1354 ();
 sg13g2_fill_2 FILLER_13_1364 ();
 sg13g2_fill_1 FILLER_13_1366 ();
 sg13g2_fill_2 FILLER_13_1373 ();
 sg13g2_fill_2 FILLER_13_1389 ();
 sg13g2_fill_1 FILLER_13_1396 ();
 sg13g2_fill_1 FILLER_13_1441 ();
 sg13g2_decap_4 FILLER_13_1447 ();
 sg13g2_fill_1 FILLER_13_1451 ();
 sg13g2_fill_2 FILLER_13_1474 ();
 sg13g2_decap_4 FILLER_13_1501 ();
 sg13g2_decap_8 FILLER_13_1515 ();
 sg13g2_decap_4 FILLER_13_1522 ();
 sg13g2_fill_2 FILLER_13_1526 ();
 sg13g2_decap_4 FILLER_13_1532 ();
 sg13g2_fill_2 FILLER_13_1536 ();
 sg13g2_fill_1 FILLER_13_1547 ();
 sg13g2_fill_1 FILLER_13_1558 ();
 sg13g2_fill_2 FILLER_13_1574 ();
 sg13g2_decap_4 FILLER_13_1604 ();
 sg13g2_decap_8 FILLER_13_1623 ();
 sg13g2_fill_2 FILLER_13_1635 ();
 sg13g2_fill_1 FILLER_13_1663 ();
 sg13g2_decap_4 FILLER_13_1672 ();
 sg13g2_fill_2 FILLER_13_1676 ();
 sg13g2_fill_2 FILLER_13_1723 ();
 sg13g2_fill_2 FILLER_13_1744 ();
 sg13g2_fill_1 FILLER_13_1746 ();
 sg13g2_fill_1 FILLER_13_1841 ();
 sg13g2_fill_2 FILLER_13_1906 ();
 sg13g2_fill_1 FILLER_13_1908 ();
 sg13g2_fill_2 FILLER_13_1923 ();
 sg13g2_fill_2 FILLER_13_1952 ();
 sg13g2_fill_1 FILLER_13_1962 ();
 sg13g2_fill_2 FILLER_13_1985 ();
 sg13g2_fill_2 FILLER_13_2018 ();
 sg13g2_fill_1 FILLER_13_2020 ();
 sg13g2_fill_2 FILLER_13_2053 ();
 sg13g2_fill_1 FILLER_13_2055 ();
 sg13g2_fill_2 FILLER_13_2065 ();
 sg13g2_fill_1 FILLER_13_2067 ();
 sg13g2_fill_1 FILLER_13_2099 ();
 sg13g2_fill_2 FILLER_13_2214 ();
 sg13g2_fill_1 FILLER_13_2216 ();
 sg13g2_fill_2 FILLER_13_2246 ();
 sg13g2_fill_1 FILLER_13_2318 ();
 sg13g2_fill_2 FILLER_13_2349 ();
 sg13g2_fill_1 FILLER_13_2351 ();
 sg13g2_fill_2 FILLER_13_2403 ();
 sg13g2_fill_2 FILLER_13_2443 ();
 sg13g2_fill_1 FILLER_13_2445 ();
 sg13g2_fill_2 FILLER_13_2520 ();
 sg13g2_fill_1 FILLER_13_2522 ();
 sg13g2_fill_1 FILLER_13_2558 ();
 sg13g2_fill_2 FILLER_13_2580 ();
 sg13g2_fill_1 FILLER_13_2582 ();
 sg13g2_decap_8 FILLER_13_2641 ();
 sg13g2_decap_8 FILLER_13_2648 ();
 sg13g2_decap_8 FILLER_13_2655 ();
 sg13g2_decap_8 FILLER_13_2662 ();
 sg13g2_decap_4 FILLER_13_2669 ();
 sg13g2_fill_1 FILLER_13_2673 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_fill_2 FILLER_14_49 ();
 sg13g2_fill_1 FILLER_14_51 ();
 sg13g2_decap_4 FILLER_14_55 ();
 sg13g2_fill_2 FILLER_14_59 ();
 sg13g2_fill_1 FILLER_14_78 ();
 sg13g2_fill_1 FILLER_14_191 ();
 sg13g2_fill_2 FILLER_14_201 ();
 sg13g2_fill_2 FILLER_14_212 ();
 sg13g2_fill_2 FILLER_14_226 ();
 sg13g2_fill_1 FILLER_14_236 ();
 sg13g2_fill_1 FILLER_14_270 ();
 sg13g2_fill_1 FILLER_14_285 ();
 sg13g2_fill_1 FILLER_14_295 ();
 sg13g2_fill_2 FILLER_14_301 ();
 sg13g2_fill_1 FILLER_14_303 ();
 sg13g2_fill_2 FILLER_14_326 ();
 sg13g2_fill_2 FILLER_14_347 ();
 sg13g2_fill_1 FILLER_14_384 ();
 sg13g2_fill_2 FILLER_14_408 ();
 sg13g2_fill_2 FILLER_14_469 ();
 sg13g2_fill_1 FILLER_14_471 ();
 sg13g2_fill_1 FILLER_14_482 ();
 sg13g2_fill_2 FILLER_14_513 ();
 sg13g2_fill_1 FILLER_14_515 ();
 sg13g2_fill_2 FILLER_14_602 ();
 sg13g2_fill_1 FILLER_14_604 ();
 sg13g2_fill_2 FILLER_14_656 ();
 sg13g2_fill_1 FILLER_14_773 ();
 sg13g2_fill_1 FILLER_14_804 ();
 sg13g2_fill_2 FILLER_14_860 ();
 sg13g2_fill_2 FILLER_14_981 ();
 sg13g2_fill_1 FILLER_14_983 ();
 sg13g2_fill_2 FILLER_14_1004 ();
 sg13g2_fill_1 FILLER_14_1006 ();
 sg13g2_fill_1 FILLER_14_1029 ();
 sg13g2_fill_1 FILLER_14_1035 ();
 sg13g2_fill_2 FILLER_14_1041 ();
 sg13g2_fill_1 FILLER_14_1043 ();
 sg13g2_fill_1 FILLER_14_1067 ();
 sg13g2_fill_2 FILLER_14_1078 ();
 sg13g2_fill_1 FILLER_14_1101 ();
 sg13g2_fill_2 FILLER_14_1117 ();
 sg13g2_fill_2 FILLER_14_1154 ();
 sg13g2_fill_1 FILLER_14_1170 ();
 sg13g2_fill_1 FILLER_14_1180 ();
 sg13g2_fill_2 FILLER_14_1293 ();
 sg13g2_fill_1 FILLER_14_1295 ();
 sg13g2_fill_2 FILLER_14_1324 ();
 sg13g2_fill_1 FILLER_14_1326 ();
 sg13g2_fill_1 FILLER_14_1345 ();
 sg13g2_fill_1 FILLER_14_1372 ();
 sg13g2_fill_2 FILLER_14_1429 ();
 sg13g2_decap_4 FILLER_14_1447 ();
 sg13g2_decap_4 FILLER_14_1486 ();
 sg13g2_fill_2 FILLER_14_1506 ();
 sg13g2_fill_1 FILLER_14_1508 ();
 sg13g2_decap_4 FILLER_14_1601 ();
 sg13g2_fill_1 FILLER_14_1605 ();
 sg13g2_fill_2 FILLER_14_1616 ();
 sg13g2_decap_4 FILLER_14_1644 ();
 sg13g2_fill_1 FILLER_14_1668 ();
 sg13g2_fill_2 FILLER_14_1772 ();
 sg13g2_fill_2 FILLER_14_1801 ();
 sg13g2_decap_4 FILLER_14_1813 ();
 sg13g2_fill_2 FILLER_14_1817 ();
 sg13g2_fill_2 FILLER_14_1870 ();
 sg13g2_fill_2 FILLER_14_1882 ();
 sg13g2_fill_2 FILLER_14_1946 ();
 sg13g2_fill_1 FILLER_14_1948 ();
 sg13g2_fill_1 FILLER_14_1972 ();
 sg13g2_fill_2 FILLER_14_2009 ();
 sg13g2_fill_1 FILLER_14_2011 ();
 sg13g2_fill_2 FILLER_14_2022 ();
 sg13g2_fill_1 FILLER_14_2024 ();
 sg13g2_fill_2 FILLER_14_2089 ();
 sg13g2_fill_1 FILLER_14_2091 ();
 sg13g2_fill_2 FILLER_14_2123 ();
 sg13g2_fill_1 FILLER_14_2125 ();
 sg13g2_fill_1 FILLER_14_2143 ();
 sg13g2_fill_2 FILLER_14_2199 ();
 sg13g2_fill_1 FILLER_14_2224 ();
 sg13g2_fill_2 FILLER_14_2260 ();
 sg13g2_fill_2 FILLER_14_2284 ();
 sg13g2_fill_2 FILLER_14_2294 ();
 sg13g2_fill_1 FILLER_14_2347 ();
 sg13g2_fill_2 FILLER_14_2367 ();
 sg13g2_fill_1 FILLER_14_2369 ();
 sg13g2_fill_2 FILLER_14_2375 ();
 sg13g2_fill_2 FILLER_14_2413 ();
 sg13g2_fill_2 FILLER_14_2429 ();
 sg13g2_fill_2 FILLER_14_2444 ();
 sg13g2_fill_1 FILLER_14_2446 ();
 sg13g2_fill_2 FILLER_14_2502 ();
 sg13g2_fill_2 FILLER_14_2530 ();
 sg13g2_fill_1 FILLER_14_2532 ();
 sg13g2_fill_2 FILLER_14_2569 ();
 sg13g2_fill_1 FILLER_14_2601 ();
 sg13g2_fill_1 FILLER_14_2612 ();
 sg13g2_decap_8 FILLER_14_2648 ();
 sg13g2_decap_8 FILLER_14_2655 ();
 sg13g2_decap_8 FILLER_14_2662 ();
 sg13g2_decap_4 FILLER_14_2669 ();
 sg13g2_fill_1 FILLER_14_2673 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_fill_1 FILLER_15_42 ();
 sg13g2_fill_1 FILLER_15_143 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_fill_2 FILLER_15_263 ();
 sg13g2_fill_1 FILLER_15_270 ();
 sg13g2_fill_2 FILLER_15_281 ();
 sg13g2_fill_1 FILLER_15_283 ();
 sg13g2_fill_2 FILLER_15_292 ();
 sg13g2_fill_2 FILLER_15_325 ();
 sg13g2_fill_2 FILLER_15_350 ();
 sg13g2_fill_2 FILLER_15_361 ();
 sg13g2_fill_1 FILLER_15_363 ();
 sg13g2_fill_1 FILLER_15_443 ();
 sg13g2_fill_1 FILLER_15_463 ();
 sg13g2_fill_1 FILLER_15_507 ();
 sg13g2_fill_2 FILLER_15_514 ();
 sg13g2_fill_2 FILLER_15_565 ();
 sg13g2_fill_2 FILLER_15_617 ();
 sg13g2_fill_2 FILLER_15_691 ();
 sg13g2_fill_2 FILLER_15_701 ();
 sg13g2_fill_1 FILLER_15_703 ();
 sg13g2_fill_2 FILLER_15_722 ();
 sg13g2_fill_1 FILLER_15_724 ();
 sg13g2_fill_2 FILLER_15_735 ();
 sg13g2_fill_1 FILLER_15_737 ();
 sg13g2_fill_2 FILLER_15_780 ();
 sg13g2_fill_1 FILLER_15_782 ();
 sg13g2_fill_2 FILLER_15_842 ();
 sg13g2_fill_1 FILLER_15_853 ();
 sg13g2_fill_2 FILLER_15_952 ();
 sg13g2_fill_1 FILLER_15_968 ();
 sg13g2_fill_2 FILLER_15_1025 ();
 sg13g2_fill_1 FILLER_15_1069 ();
 sg13g2_fill_2 FILLER_15_1126 ();
 sg13g2_fill_1 FILLER_15_1128 ();
 sg13g2_fill_1 FILLER_15_1274 ();
 sg13g2_fill_2 FILLER_15_1284 ();
 sg13g2_fill_2 FILLER_15_1312 ();
 sg13g2_fill_1 FILLER_15_1335 ();
 sg13g2_decap_8 FILLER_15_1361 ();
 sg13g2_fill_2 FILLER_15_1368 ();
 sg13g2_fill_1 FILLER_15_1370 ();
 sg13g2_fill_2 FILLER_15_1403 ();
 sg13g2_fill_1 FILLER_15_1405 ();
 sg13g2_fill_1 FILLER_15_1433 ();
 sg13g2_decap_8 FILLER_15_1454 ();
 sg13g2_fill_1 FILLER_15_1461 ();
 sg13g2_fill_2 FILLER_15_1466 ();
 sg13g2_fill_1 FILLER_15_1468 ();
 sg13g2_decap_4 FILLER_15_1515 ();
 sg13g2_fill_1 FILLER_15_1519 ();
 sg13g2_fill_2 FILLER_15_1524 ();
 sg13g2_decap_4 FILLER_15_1530 ();
 sg13g2_fill_1 FILLER_15_1534 ();
 sg13g2_fill_1 FILLER_15_1545 ();
 sg13g2_fill_2 FILLER_15_1554 ();
 sg13g2_fill_2 FILLER_15_1582 ();
 sg13g2_fill_1 FILLER_15_1584 ();
 sg13g2_fill_2 FILLER_15_1604 ();
 sg13g2_decap_4 FILLER_15_1624 ();
 sg13g2_fill_1 FILLER_15_1628 ();
 sg13g2_decap_4 FILLER_15_1672 ();
 sg13g2_fill_2 FILLER_15_1676 ();
 sg13g2_fill_2 FILLER_15_1691 ();
 sg13g2_fill_1 FILLER_15_1733 ();
 sg13g2_fill_1 FILLER_15_1748 ();
 sg13g2_fill_2 FILLER_15_1783 ();
 sg13g2_fill_1 FILLER_15_1808 ();
 sg13g2_fill_1 FILLER_15_1857 ();
 sg13g2_fill_2 FILLER_15_1920 ();
 sg13g2_fill_1 FILLER_15_1922 ();
 sg13g2_fill_1 FILLER_15_1962 ();
 sg13g2_fill_2 FILLER_15_1989 ();
 sg13g2_fill_1 FILLER_15_1991 ();
 sg13g2_fill_1 FILLER_15_2103 ();
 sg13g2_fill_1 FILLER_15_2123 ();
 sg13g2_fill_1 FILLER_15_2178 ();
 sg13g2_fill_2 FILLER_15_2239 ();
 sg13g2_fill_1 FILLER_15_2241 ();
 sg13g2_fill_1 FILLER_15_2334 ();
 sg13g2_fill_1 FILLER_15_2382 ();
 sg13g2_fill_2 FILLER_15_2529 ();
 sg13g2_fill_1 FILLER_15_2531 ();
 sg13g2_fill_2 FILLER_15_2561 ();
 sg13g2_fill_1 FILLER_15_2563 ();
 sg13g2_fill_2 FILLER_15_2589 ();
 sg13g2_fill_1 FILLER_15_2591 ();
 sg13g2_fill_1 FILLER_15_2613 ();
 sg13g2_decap_8 FILLER_15_2653 ();
 sg13g2_decap_8 FILLER_15_2660 ();
 sg13g2_decap_8 FILLER_15_2667 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_4 FILLER_16_21 ();
 sg13g2_fill_1 FILLER_16_25 ();
 sg13g2_fill_1 FILLER_16_117 ();
 sg13g2_fill_1 FILLER_16_133 ();
 sg13g2_fill_1 FILLER_16_139 ();
 sg13g2_fill_1 FILLER_16_194 ();
 sg13g2_fill_1 FILLER_16_216 ();
 sg13g2_fill_1 FILLER_16_224 ();
 sg13g2_fill_2 FILLER_16_236 ();
 sg13g2_fill_1 FILLER_16_238 ();
 sg13g2_fill_1 FILLER_16_268 ();
 sg13g2_fill_1 FILLER_16_289 ();
 sg13g2_fill_2 FILLER_16_295 ();
 sg13g2_fill_2 FILLER_16_392 ();
 sg13g2_fill_1 FILLER_16_394 ();
 sg13g2_fill_2 FILLER_16_425 ();
 sg13g2_fill_1 FILLER_16_427 ();
 sg13g2_fill_1 FILLER_16_433 ();
 sg13g2_fill_2 FILLER_16_477 ();
 sg13g2_fill_2 FILLER_16_520 ();
 sg13g2_fill_1 FILLER_16_522 ();
 sg13g2_fill_2 FILLER_16_593 ();
 sg13g2_fill_2 FILLER_16_642 ();
 sg13g2_fill_1 FILLER_16_673 ();
 sg13g2_fill_1 FILLER_16_770 ();
 sg13g2_fill_2 FILLER_16_797 ();
 sg13g2_fill_2 FILLER_16_812 ();
 sg13g2_fill_1 FILLER_16_814 ();
 sg13g2_fill_2 FILLER_16_888 ();
 sg13g2_fill_1 FILLER_16_890 ();
 sg13g2_fill_2 FILLER_16_936 ();
 sg13g2_fill_1 FILLER_16_983 ();
 sg13g2_fill_1 FILLER_16_1008 ();
 sg13g2_fill_2 FILLER_16_1023 ();
 sg13g2_fill_2 FILLER_16_1039 ();
 sg13g2_fill_2 FILLER_16_1067 ();
 sg13g2_fill_1 FILLER_16_1074 ();
 sg13g2_fill_2 FILLER_16_1134 ();
 sg13g2_fill_2 FILLER_16_1165 ();
 sg13g2_fill_1 FILLER_16_1208 ();
 sg13g2_fill_2 FILLER_16_1277 ();
 sg13g2_fill_1 FILLER_16_1279 ();
 sg13g2_fill_2 FILLER_16_1300 ();
 sg13g2_fill_1 FILLER_16_1302 ();
 sg13g2_fill_2 FILLER_16_1322 ();
 sg13g2_fill_2 FILLER_16_1329 ();
 sg13g2_fill_2 FILLER_16_1352 ();
 sg13g2_fill_2 FILLER_16_1375 ();
 sg13g2_fill_2 FILLER_16_1382 ();
 sg13g2_fill_1 FILLER_16_1389 ();
 sg13g2_fill_1 FILLER_16_1425 ();
 sg13g2_fill_1 FILLER_16_1451 ();
 sg13g2_fill_1 FILLER_16_1460 ();
 sg13g2_fill_2 FILLER_16_1466 ();
 sg13g2_fill_1 FILLER_16_1468 ();
 sg13g2_fill_1 FILLER_16_1474 ();
 sg13g2_fill_1 FILLER_16_1487 ();
 sg13g2_fill_1 FILLER_16_1514 ();
 sg13g2_decap_4 FILLER_16_1519 ();
 sg13g2_fill_2 FILLER_16_1523 ();
 sg13g2_fill_2 FILLER_16_1542 ();
 sg13g2_fill_1 FILLER_16_1544 ();
 sg13g2_fill_2 FILLER_16_1571 ();
 sg13g2_fill_1 FILLER_16_1573 ();
 sg13g2_fill_1 FILLER_16_1596 ();
 sg13g2_decap_4 FILLER_16_1600 ();
 sg13g2_fill_1 FILLER_16_1604 ();
 sg13g2_fill_2 FILLER_16_1644 ();
 sg13g2_fill_1 FILLER_16_1646 ();
 sg13g2_fill_2 FILLER_16_1664 ();
 sg13g2_fill_2 FILLER_16_1702 ();
 sg13g2_fill_2 FILLER_16_1765 ();
 sg13g2_fill_1 FILLER_16_1767 ();
 sg13g2_fill_2 FILLER_16_1847 ();
 sg13g2_fill_1 FILLER_16_1849 ();
 sg13g2_fill_2 FILLER_16_1866 ();
 sg13g2_fill_2 FILLER_16_1893 ();
 sg13g2_fill_1 FILLER_16_1895 ();
 sg13g2_fill_1 FILLER_16_1942 ();
 sg13g2_fill_1 FILLER_16_1953 ();
 sg13g2_fill_2 FILLER_16_1975 ();
 sg13g2_fill_2 FILLER_16_1987 ();
 sg13g2_fill_1 FILLER_16_1989 ();
 sg13g2_fill_2 FILLER_16_2046 ();
 sg13g2_fill_1 FILLER_16_2048 ();
 sg13g2_fill_2 FILLER_16_2068 ();
 sg13g2_fill_1 FILLER_16_2070 ();
 sg13g2_fill_2 FILLER_16_2081 ();
 sg13g2_fill_2 FILLER_16_2129 ();
 sg13g2_fill_1 FILLER_16_2131 ();
 sg13g2_fill_2 FILLER_16_2147 ();
 sg13g2_fill_1 FILLER_16_2149 ();
 sg13g2_fill_2 FILLER_16_2206 ();
 sg13g2_fill_1 FILLER_16_2208 ();
 sg13g2_fill_2 FILLER_16_2241 ();
 sg13g2_fill_1 FILLER_16_2243 ();
 sg13g2_fill_2 FILLER_16_2299 ();
 sg13g2_fill_2 FILLER_16_2370 ();
 sg13g2_fill_1 FILLER_16_2384 ();
 sg13g2_fill_1 FILLER_16_2391 ();
 sg13g2_fill_2 FILLER_16_2438 ();
 sg13g2_fill_1 FILLER_16_2524 ();
 sg13g2_fill_2 FILLER_16_2538 ();
 sg13g2_fill_1 FILLER_16_2540 ();
 sg13g2_fill_2 FILLER_16_2567 ();
 sg13g2_fill_1 FILLER_16_2569 ();
 sg13g2_fill_1 FILLER_16_2605 ();
 sg13g2_fill_2 FILLER_16_2625 ();
 sg13g2_decap_8 FILLER_16_2656 ();
 sg13g2_decap_8 FILLER_16_2663 ();
 sg13g2_decap_4 FILLER_16_2670 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_fill_2 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_51 ();
 sg13g2_fill_2 FILLER_17_85 ();
 sg13g2_fill_2 FILLER_17_110 ();
 sg13g2_fill_2 FILLER_17_247 ();
 sg13g2_fill_1 FILLER_17_249 ();
 sg13g2_fill_2 FILLER_17_265 ();
 sg13g2_fill_2 FILLER_17_272 ();
 sg13g2_fill_2 FILLER_17_292 ();
 sg13g2_fill_1 FILLER_17_333 ();
 sg13g2_fill_2 FILLER_17_348 ();
 sg13g2_fill_2 FILLER_17_398 ();
 sg13g2_fill_2 FILLER_17_442 ();
 sg13g2_fill_1 FILLER_17_470 ();
 sg13g2_fill_2 FILLER_17_484 ();
 sg13g2_fill_1 FILLER_17_486 ();
 sg13g2_fill_2 FILLER_17_513 ();
 sg13g2_fill_1 FILLER_17_515 ();
 sg13g2_fill_1 FILLER_17_521 ();
 sg13g2_fill_1 FILLER_17_543 ();
 sg13g2_fill_2 FILLER_17_579 ();
 sg13g2_fill_1 FILLER_17_581 ();
 sg13g2_fill_2 FILLER_17_638 ();
 sg13g2_fill_1 FILLER_17_640 ();
 sg13g2_fill_2 FILLER_17_649 ();
 sg13g2_fill_1 FILLER_17_651 ();
 sg13g2_fill_2 FILLER_17_720 ();
 sg13g2_fill_1 FILLER_17_722 ();
 sg13g2_fill_2 FILLER_17_733 ();
 sg13g2_fill_2 FILLER_17_741 ();
 sg13g2_fill_1 FILLER_17_743 ();
 sg13g2_fill_2 FILLER_17_758 ();
 sg13g2_fill_1 FILLER_17_760 ();
 sg13g2_fill_1 FILLER_17_785 ();
 sg13g2_fill_1 FILLER_17_822 ();
 sg13g2_fill_1 FILLER_17_890 ();
 sg13g2_fill_1 FILLER_17_902 ();
 sg13g2_fill_1 FILLER_17_912 ();
 sg13g2_fill_2 FILLER_17_947 ();
 sg13g2_fill_2 FILLER_17_1014 ();
 sg13g2_fill_2 FILLER_17_1047 ();
 sg13g2_fill_2 FILLER_17_1059 ();
 sg13g2_fill_1 FILLER_17_1100 ();
 sg13g2_fill_2 FILLER_17_1111 ();
 sg13g2_fill_2 FILLER_17_1169 ();
 sg13g2_fill_1 FILLER_17_1240 ();
 sg13g2_decap_8 FILLER_17_1296 ();
 sg13g2_fill_1 FILLER_17_1341 ();
 sg13g2_fill_2 FILLER_17_1378 ();
 sg13g2_fill_2 FILLER_17_1385 ();
 sg13g2_fill_1 FILLER_17_1392 ();
 sg13g2_fill_2 FILLER_17_1423 ();
 sg13g2_fill_2 FILLER_17_1440 ();
 sg13g2_fill_1 FILLER_17_1498 ();
 sg13g2_fill_1 FILLER_17_1555 ();
 sg13g2_fill_2 FILLER_17_1595 ();
 sg13g2_fill_1 FILLER_17_1623 ();
 sg13g2_fill_2 FILLER_17_1632 ();
 sg13g2_fill_1 FILLER_17_1634 ();
 sg13g2_fill_2 FILLER_17_1661 ();
 sg13g2_fill_1 FILLER_17_1735 ();
 sg13g2_fill_2 FILLER_17_1758 ();
 sg13g2_fill_1 FILLER_17_1760 ();
 sg13g2_fill_2 FILLER_17_1794 ();
 sg13g2_fill_1 FILLER_17_1796 ();
 sg13g2_fill_1 FILLER_17_1837 ();
 sg13g2_fill_1 FILLER_17_1880 ();
 sg13g2_fill_1 FILLER_17_2009 ();
 sg13g2_fill_2 FILLER_17_2080 ();
 sg13g2_fill_2 FILLER_17_2090 ();
 sg13g2_fill_1 FILLER_17_2092 ();
 sg13g2_fill_1 FILLER_17_2145 ();
 sg13g2_fill_2 FILLER_17_2161 ();
 sg13g2_fill_1 FILLER_17_2172 ();
 sg13g2_fill_2 FILLER_17_2182 ();
 sg13g2_fill_1 FILLER_17_2219 ();
 sg13g2_fill_2 FILLER_17_2246 ();
 sg13g2_fill_2 FILLER_17_2274 ();
 sg13g2_fill_1 FILLER_17_2276 ();
 sg13g2_fill_2 FILLER_17_2324 ();
 sg13g2_fill_1 FILLER_17_2326 ();
 sg13g2_fill_2 FILLER_17_2342 ();
 sg13g2_fill_1 FILLER_17_2344 ();
 sg13g2_fill_2 FILLER_17_2472 ();
 sg13g2_fill_1 FILLER_17_2474 ();
 sg13g2_fill_1 FILLER_17_2489 ();
 sg13g2_fill_1 FILLER_17_2570 ();
 sg13g2_fill_1 FILLER_17_2617 ();
 sg13g2_decap_8 FILLER_17_2648 ();
 sg13g2_decap_8 FILLER_17_2655 ();
 sg13g2_decap_8 FILLER_17_2662 ();
 sg13g2_decap_4 FILLER_17_2669 ();
 sg13g2_fill_1 FILLER_17_2673 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_51 ();
 sg13g2_fill_2 FILLER_18_59 ();
 sg13g2_fill_1 FILLER_18_71 ();
 sg13g2_fill_1 FILLER_18_133 ();
 sg13g2_fill_2 FILLER_18_154 ();
 sg13g2_fill_1 FILLER_18_205 ();
 sg13g2_fill_2 FILLER_18_219 ();
 sg13g2_fill_1 FILLER_18_221 ();
 sg13g2_fill_2 FILLER_18_275 ();
 sg13g2_fill_1 FILLER_18_277 ();
 sg13g2_fill_1 FILLER_18_291 ();
 sg13g2_fill_2 FILLER_18_324 ();
 sg13g2_fill_2 FILLER_18_370 ();
 sg13g2_fill_2 FILLER_18_438 ();
 sg13g2_fill_2 FILLER_18_464 ();
 sg13g2_fill_1 FILLER_18_484 ();
 sg13g2_fill_2 FILLER_18_511 ();
 sg13g2_fill_1 FILLER_18_513 ();
 sg13g2_fill_1 FILLER_18_682 ();
 sg13g2_fill_2 FILLER_18_691 ();
 sg13g2_fill_2 FILLER_18_735 ();
 sg13g2_fill_1 FILLER_18_737 ();
 sg13g2_fill_1 FILLER_18_774 ();
 sg13g2_fill_1 FILLER_18_784 ();
 sg13g2_fill_2 FILLER_18_795 ();
 sg13g2_fill_2 FILLER_18_802 ();
 sg13g2_fill_1 FILLER_18_822 ();
 sg13g2_fill_2 FILLER_18_872 ();
 sg13g2_fill_1 FILLER_18_925 ();
 sg13g2_fill_2 FILLER_18_943 ();
 sg13g2_fill_2 FILLER_18_980 ();
 sg13g2_fill_1 FILLER_18_1013 ();
 sg13g2_fill_1 FILLER_18_1085 ();
 sg13g2_fill_1 FILLER_18_1117 ();
 sg13g2_fill_2 FILLER_18_1174 ();
 sg13g2_fill_1 FILLER_18_1257 ();
 sg13g2_fill_1 FILLER_18_1267 ();
 sg13g2_fill_2 FILLER_18_1282 ();
 sg13g2_fill_1 FILLER_18_1284 ();
 sg13g2_fill_1 FILLER_18_1361 ();
 sg13g2_decap_4 FILLER_18_1420 ();
 sg13g2_fill_2 FILLER_18_1424 ();
 sg13g2_fill_2 FILLER_18_1450 ();
 sg13g2_fill_1 FILLER_18_1452 ();
 sg13g2_fill_2 FILLER_18_1484 ();
 sg13g2_fill_1 FILLER_18_1486 ();
 sg13g2_fill_1 FILLER_18_1491 ();
 sg13g2_decap_4 FILLER_18_1519 ();
 sg13g2_fill_2 FILLER_18_1523 ();
 sg13g2_fill_1 FILLER_18_1542 ();
 sg13g2_decap_4 FILLER_18_1555 ();
 sg13g2_fill_2 FILLER_18_1564 ();
 sg13g2_fill_1 FILLER_18_1566 ();
 sg13g2_decap_8 FILLER_18_1575 ();
 sg13g2_fill_1 FILLER_18_1582 ();
 sg13g2_fill_2 FILLER_18_1596 ();
 sg13g2_fill_1 FILLER_18_1598 ();
 sg13g2_fill_2 FILLER_18_1626 ();
 sg13g2_fill_2 FILLER_18_1641 ();
 sg13g2_fill_1 FILLER_18_1653 ();
 sg13g2_fill_2 FILLER_18_1719 ();
 sg13g2_fill_1 FILLER_18_1721 ();
 sg13g2_fill_1 FILLER_18_1743 ();
 sg13g2_fill_2 FILLER_18_1748 ();
 sg13g2_fill_1 FILLER_18_1826 ();
 sg13g2_fill_2 FILLER_18_1833 ();
 sg13g2_fill_1 FILLER_18_1835 ();
 sg13g2_fill_1 FILLER_18_1846 ();
 sg13g2_fill_1 FILLER_18_1902 ();
 sg13g2_fill_2 FILLER_18_1939 ();
 sg13g2_fill_1 FILLER_18_1941 ();
 sg13g2_fill_2 FILLER_18_1968 ();
 sg13g2_fill_1 FILLER_18_2056 ();
 sg13g2_fill_2 FILLER_18_2107 ();
 sg13g2_fill_2 FILLER_18_2118 ();
 sg13g2_fill_2 FILLER_18_2193 ();
 sg13g2_fill_2 FILLER_18_2212 ();
 sg13g2_fill_1 FILLER_18_2262 ();
 sg13g2_fill_1 FILLER_18_2287 ();
 sg13g2_fill_2 FILLER_18_2343 ();
 sg13g2_fill_1 FILLER_18_2345 ();
 sg13g2_fill_1 FILLER_18_2494 ();
 sg13g2_fill_2 FILLER_18_2539 ();
 sg13g2_fill_1 FILLER_18_2541 ();
 sg13g2_decap_8 FILLER_18_2651 ();
 sg13g2_decap_8 FILLER_18_2658 ();
 sg13g2_decap_8 FILLER_18_2665 ();
 sg13g2_fill_2 FILLER_18_2672 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_7 ();
 sg13g2_fill_1 FILLER_19_13 ();
 sg13g2_fill_2 FILLER_19_49 ();
 sg13g2_fill_2 FILLER_19_59 ();
 sg13g2_fill_1 FILLER_19_147 ();
 sg13g2_fill_1 FILLER_19_195 ();
 sg13g2_fill_2 FILLER_19_201 ();
 sg13g2_fill_1 FILLER_19_203 ();
 sg13g2_fill_1 FILLER_19_209 ();
 sg13g2_fill_1 FILLER_19_264 ();
 sg13g2_fill_1 FILLER_19_316 ();
 sg13g2_fill_1 FILLER_19_335 ();
 sg13g2_fill_2 FILLER_19_396 ();
 sg13g2_fill_2 FILLER_19_418 ();
 sg13g2_fill_2 FILLER_19_429 ();
 sg13g2_fill_1 FILLER_19_431 ();
 sg13g2_fill_2 FILLER_19_446 ();
 sg13g2_fill_1 FILLER_19_474 ();
 sg13g2_fill_1 FILLER_19_489 ();
 sg13g2_fill_2 FILLER_19_511 ();
 sg13g2_fill_1 FILLER_19_513 ();
 sg13g2_fill_1 FILLER_19_560 ();
 sg13g2_fill_2 FILLER_19_584 ();
 sg13g2_fill_1 FILLER_19_613 ();
 sg13g2_fill_2 FILLER_19_630 ();
 sg13g2_fill_1 FILLER_19_632 ();
 sg13g2_fill_2 FILLER_19_713 ();
 sg13g2_fill_2 FILLER_19_738 ();
 sg13g2_fill_1 FILLER_19_855 ();
 sg13g2_fill_1 FILLER_19_887 ();
 sg13g2_fill_2 FILLER_19_897 ();
 sg13g2_fill_1 FILLER_19_899 ();
 sg13g2_fill_1 FILLER_19_936 ();
 sg13g2_fill_2 FILLER_19_942 ();
 sg13g2_fill_1 FILLER_19_944 ();
 sg13g2_fill_1 FILLER_19_993 ();
 sg13g2_fill_1 FILLER_19_1024 ();
 sg13g2_fill_2 FILLER_19_1080 ();
 sg13g2_fill_1 FILLER_19_1082 ();
 sg13g2_fill_2 FILLER_19_1248 ();
 sg13g2_decap_4 FILLER_19_1286 ();
 sg13g2_decap_4 FILLER_19_1305 ();
 sg13g2_fill_2 FILLER_19_1314 ();
 sg13g2_decap_4 FILLER_19_1343 ();
 sg13g2_decap_4 FILLER_19_1361 ();
 sg13g2_fill_2 FILLER_19_1365 ();
 sg13g2_decap_8 FILLER_19_1371 ();
 sg13g2_decap_4 FILLER_19_1382 ();
 sg13g2_fill_2 FILLER_19_1396 ();
 sg13g2_fill_1 FILLER_19_1398 ();
 sg13g2_fill_2 FILLER_19_1437 ();
 sg13g2_fill_1 FILLER_19_1546 ();
 sg13g2_decap_4 FILLER_19_1570 ();
 sg13g2_fill_2 FILLER_19_1574 ();
 sg13g2_fill_1 FILLER_19_1588 ();
 sg13g2_fill_1 FILLER_19_1594 ();
 sg13g2_fill_1 FILLER_19_1620 ();
 sg13g2_fill_1 FILLER_19_1647 ();
 sg13g2_fill_2 FILLER_19_1660 ();
 sg13g2_fill_1 FILLER_19_1662 ();
 sg13g2_fill_1 FILLER_19_1676 ();
 sg13g2_fill_2 FILLER_19_1703 ();
 sg13g2_fill_1 FILLER_19_1736 ();
 sg13g2_fill_1 FILLER_19_1763 ();
 sg13g2_fill_1 FILLER_19_1774 ();
 sg13g2_fill_2 FILLER_19_1789 ();
 sg13g2_fill_1 FILLER_19_1791 ();
 sg13g2_fill_1 FILLER_19_1870 ();
 sg13g2_fill_2 FILLER_19_1886 ();
 sg13g2_fill_2 FILLER_19_1919 ();
 sg13g2_fill_1 FILLER_19_1921 ();
 sg13g2_fill_2 FILLER_19_1969 ();
 sg13g2_fill_1 FILLER_19_2005 ();
 sg13g2_fill_2 FILLER_19_2045 ();
 sg13g2_fill_1 FILLER_19_2047 ();
 sg13g2_fill_2 FILLER_19_2173 ();
 sg13g2_fill_1 FILLER_19_2175 ();
 sg13g2_fill_2 FILLER_19_2284 ();
 sg13g2_fill_1 FILLER_19_2312 ();
 sg13g2_fill_2 FILLER_19_2331 ();
 sg13g2_fill_1 FILLER_19_2333 ();
 sg13g2_fill_1 FILLER_19_2353 ();
 sg13g2_fill_1 FILLER_19_2397 ();
 sg13g2_fill_1 FILLER_19_2441 ();
 sg13g2_fill_1 FILLER_19_2491 ();
 sg13g2_fill_1 FILLER_19_2522 ();
 sg13g2_fill_2 FILLER_19_2600 ();
 sg13g2_decap_8 FILLER_19_2650 ();
 sg13g2_decap_8 FILLER_19_2657 ();
 sg13g2_decap_8 FILLER_19_2664 ();
 sg13g2_fill_2 FILLER_19_2671 ();
 sg13g2_fill_1 FILLER_19_2673 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_25 ();
 sg13g2_fill_1 FILLER_20_54 ();
 sg13g2_fill_1 FILLER_20_80 ();
 sg13g2_fill_1 FILLER_20_86 ();
 sg13g2_fill_2 FILLER_20_140 ();
 sg13g2_fill_2 FILLER_20_187 ();
 sg13g2_fill_2 FILLER_20_211 ();
 sg13g2_fill_1 FILLER_20_231 ();
 sg13g2_fill_2 FILLER_20_237 ();
 sg13g2_fill_1 FILLER_20_249 ();
 sg13g2_fill_2 FILLER_20_296 ();
 sg13g2_fill_1 FILLER_20_343 ();
 sg13g2_fill_2 FILLER_20_458 ();
 sg13g2_fill_1 FILLER_20_491 ();
 sg13g2_fill_1 FILLER_20_535 ();
 sg13g2_fill_2 FILLER_20_541 ();
 sg13g2_fill_2 FILLER_20_579 ();
 sg13g2_fill_1 FILLER_20_581 ();
 sg13g2_fill_2 FILLER_20_648 ();
 sg13g2_fill_2 FILLER_20_690 ();
 sg13g2_fill_1 FILLER_20_711 ();
 sg13g2_fill_1 FILLER_20_741 ();
 sg13g2_fill_2 FILLER_20_763 ();
 sg13g2_fill_2 FILLER_20_800 ();
 sg13g2_fill_2 FILLER_20_843 ();
 sg13g2_fill_1 FILLER_20_870 ();
 sg13g2_fill_1 FILLER_20_877 ();
 sg13g2_fill_2 FILLER_20_908 ();
 sg13g2_fill_2 FILLER_20_915 ();
 sg13g2_fill_1 FILLER_20_917 ();
 sg13g2_fill_1 FILLER_20_969 ();
 sg13g2_fill_1 FILLER_20_1018 ();
 sg13g2_fill_2 FILLER_20_1094 ();
 sg13g2_fill_2 FILLER_20_1120 ();
 sg13g2_fill_2 FILLER_20_1153 ();
 sg13g2_fill_1 FILLER_20_1155 ();
 sg13g2_fill_2 FILLER_20_1173 ();
 sg13g2_fill_1 FILLER_20_1175 ();
 sg13g2_fill_2 FILLER_20_1223 ();
 sg13g2_fill_1 FILLER_20_1225 ();
 sg13g2_fill_2 FILLER_20_1245 ();
 sg13g2_fill_1 FILLER_20_1247 ();
 sg13g2_fill_2 FILLER_20_1269 ();
 sg13g2_fill_1 FILLER_20_1271 ();
 sg13g2_fill_1 FILLER_20_1281 ();
 sg13g2_decap_8 FILLER_20_1298 ();
 sg13g2_fill_1 FILLER_20_1328 ();
 sg13g2_fill_1 FILLER_20_1334 ();
 sg13g2_fill_1 FILLER_20_1347 ();
 sg13g2_decap_4 FILLER_20_1398 ();
 sg13g2_fill_2 FILLER_20_1402 ();
 sg13g2_decap_8 FILLER_20_1418 ();
 sg13g2_fill_2 FILLER_20_1425 ();
 sg13g2_fill_2 FILLER_20_1432 ();
 sg13g2_decap_8 FILLER_20_1443 ();
 sg13g2_decap_8 FILLER_20_1454 ();
 sg13g2_fill_1 FILLER_20_1461 ();
 sg13g2_fill_1 FILLER_20_1488 ();
 sg13g2_decap_4 FILLER_20_1503 ();
 sg13g2_fill_1 FILLER_20_1507 ();
 sg13g2_fill_1 FILLER_20_1535 ();
 sg13g2_fill_2 FILLER_20_1573 ();
 sg13g2_fill_1 FILLER_20_1575 ();
 sg13g2_fill_1 FILLER_20_1594 ();
 sg13g2_fill_2 FILLER_20_1603 ();
 sg13g2_fill_1 FILLER_20_1605 ();
 sg13g2_fill_2 FILLER_20_1616 ();
 sg13g2_fill_1 FILLER_20_1632 ();
 sg13g2_fill_2 FILLER_20_1642 ();
 sg13g2_fill_1 FILLER_20_1676 ();
 sg13g2_fill_1 FILLER_20_1689 ();
 sg13g2_fill_1 FILLER_20_1709 ();
 sg13g2_fill_1 FILLER_20_1753 ();
 sg13g2_fill_2 FILLER_20_1768 ();
 sg13g2_fill_1 FILLER_20_1770 ();
 sg13g2_fill_1 FILLER_20_1829 ();
 sg13g2_decap_4 FILLER_20_1866 ();
 sg13g2_fill_1 FILLER_20_1870 ();
 sg13g2_fill_2 FILLER_20_1883 ();
 sg13g2_fill_1 FILLER_20_1885 ();
 sg13g2_fill_2 FILLER_20_1907 ();
 sg13g2_fill_2 FILLER_20_1963 ();
 sg13g2_fill_2 FILLER_20_1984 ();
 sg13g2_fill_2 FILLER_20_2034 ();
 sg13g2_fill_1 FILLER_20_2036 ();
 sg13g2_fill_1 FILLER_20_2166 ();
 sg13g2_fill_2 FILLER_20_2181 ();
 sg13g2_fill_1 FILLER_20_2183 ();
 sg13g2_fill_1 FILLER_20_2213 ();
 sg13g2_fill_2 FILLER_20_2233 ();
 sg13g2_fill_2 FILLER_20_2277 ();
 sg13g2_fill_1 FILLER_20_2288 ();
 sg13g2_fill_1 FILLER_20_2301 ();
 sg13g2_fill_1 FILLER_20_2362 ();
 sg13g2_fill_2 FILLER_20_2393 ();
 sg13g2_fill_2 FILLER_20_2448 ();
 sg13g2_fill_2 FILLER_20_2471 ();
 sg13g2_fill_1 FILLER_20_2473 ();
 sg13g2_fill_1 FILLER_20_2515 ();
 sg13g2_fill_2 FILLER_20_2568 ();
 sg13g2_decap_8 FILLER_20_2650 ();
 sg13g2_decap_8 FILLER_20_2657 ();
 sg13g2_decap_8 FILLER_20_2664 ();
 sg13g2_fill_2 FILLER_20_2671 ();
 sg13g2_fill_1 FILLER_20_2673 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_53 ();
 sg13g2_fill_1 FILLER_21_55 ();
 sg13g2_fill_2 FILLER_21_82 ();
 sg13g2_fill_1 FILLER_21_101 ();
 sg13g2_fill_2 FILLER_21_121 ();
 sg13g2_fill_1 FILLER_21_128 ();
 sg13g2_fill_2 FILLER_21_156 ();
 sg13g2_fill_1 FILLER_21_158 ();
 sg13g2_fill_2 FILLER_21_164 ();
 sg13g2_fill_1 FILLER_21_252 ();
 sg13g2_fill_1 FILLER_21_266 ();
 sg13g2_fill_2 FILLER_21_272 ();
 sg13g2_fill_1 FILLER_21_312 ();
 sg13g2_fill_2 FILLER_21_318 ();
 sg13g2_fill_2 FILLER_21_346 ();
 sg13g2_fill_2 FILLER_21_386 ();
 sg13g2_fill_1 FILLER_21_388 ();
 sg13g2_fill_2 FILLER_21_415 ();
 sg13g2_fill_2 FILLER_21_457 ();
 sg13g2_fill_1 FILLER_21_459 ();
 sg13g2_fill_2 FILLER_21_478 ();
 sg13g2_fill_1 FILLER_21_480 ();
 sg13g2_fill_1 FILLER_21_503 ();
 sg13g2_fill_2 FILLER_21_546 ();
 sg13g2_fill_2 FILLER_21_562 ();
 sg13g2_fill_2 FILLER_21_570 ();
 sg13g2_fill_1 FILLER_21_572 ();
 sg13g2_fill_2 FILLER_21_608 ();
 sg13g2_fill_2 FILLER_21_619 ();
 sg13g2_fill_1 FILLER_21_634 ();
 sg13g2_fill_1 FILLER_21_664 ();
 sg13g2_fill_1 FILLER_21_742 ();
 sg13g2_fill_2 FILLER_21_801 ();
 sg13g2_fill_2 FILLER_21_938 ();
 sg13g2_fill_2 FILLER_21_953 ();
 sg13g2_fill_2 FILLER_21_1023 ();
 sg13g2_fill_1 FILLER_21_1025 ();
 sg13g2_fill_2 FILLER_21_1031 ();
 sg13g2_fill_1 FILLER_21_1033 ();
 sg13g2_fill_2 FILLER_21_1038 ();
 sg13g2_fill_1 FILLER_21_1040 ();
 sg13g2_fill_2 FILLER_21_1067 ();
 sg13g2_fill_1 FILLER_21_1069 ();
 sg13g2_fill_1 FILLER_21_1128 ();
 sg13g2_fill_1 FILLER_21_1212 ();
 sg13g2_fill_2 FILLER_21_1285 ();
 sg13g2_fill_1 FILLER_21_1316 ();
 sg13g2_fill_2 FILLER_21_1343 ();
 sg13g2_fill_2 FILLER_21_1401 ();
 sg13g2_fill_1 FILLER_21_1403 ();
 sg13g2_fill_2 FILLER_21_1423 ();
 sg13g2_fill_1 FILLER_21_1452 ();
 sg13g2_fill_2 FILLER_21_1478 ();
 sg13g2_fill_1 FILLER_21_1522 ();
 sg13g2_fill_1 FILLER_21_1547 ();
 sg13g2_fill_2 FILLER_21_1556 ();
 sg13g2_fill_1 FILLER_21_1558 ();
 sg13g2_decap_8 FILLER_21_1564 ();
 sg13g2_fill_2 FILLER_21_1571 ();
 sg13g2_fill_1 FILLER_21_1573 ();
 sg13g2_fill_2 FILLER_21_1590 ();
 sg13g2_fill_2 FILLER_21_1598 ();
 sg13g2_fill_1 FILLER_21_1600 ();
 sg13g2_fill_1 FILLER_21_1608 ();
 sg13g2_fill_2 FILLER_21_1648 ();
 sg13g2_fill_1 FILLER_21_1664 ();
 sg13g2_fill_2 FILLER_21_1671 ();
 sg13g2_fill_1 FILLER_21_1673 ();
 sg13g2_fill_2 FILLER_21_1804 ();
 sg13g2_fill_2 FILLER_21_1821 ();
 sg13g2_fill_1 FILLER_21_1823 ();
 sg13g2_fill_1 FILLER_21_1874 ();
 sg13g2_fill_2 FILLER_21_1889 ();
 sg13g2_fill_2 FILLER_21_1909 ();
 sg13g2_fill_1 FILLER_21_1911 ();
 sg13g2_fill_2 FILLER_21_1938 ();
 sg13g2_fill_1 FILLER_21_1940 ();
 sg13g2_fill_2 FILLER_21_1967 ();
 sg13g2_fill_2 FILLER_21_2071 ();
 sg13g2_fill_1 FILLER_21_2117 ();
 sg13g2_fill_1 FILLER_21_2131 ();
 sg13g2_fill_1 FILLER_21_2146 ();
 sg13g2_fill_1 FILLER_21_2217 ();
 sg13g2_fill_1 FILLER_21_2245 ();
 sg13g2_fill_2 FILLER_21_2298 ();
 sg13g2_fill_1 FILLER_21_2300 ();
 sg13g2_fill_1 FILLER_21_2326 ();
 sg13g2_fill_1 FILLER_21_2389 ();
 sg13g2_fill_2 FILLER_21_2400 ();
 sg13g2_fill_1 FILLER_21_2402 ();
 sg13g2_fill_2 FILLER_21_2452 ();
 sg13g2_fill_1 FILLER_21_2454 ();
 sg13g2_fill_2 FILLER_21_2499 ();
 sg13g2_fill_1 FILLER_21_2510 ();
 sg13g2_fill_1 FILLER_21_2551 ();
 sg13g2_fill_2 FILLER_21_2594 ();
 sg13g2_fill_1 FILLER_21_2596 ();
 sg13g2_fill_2 FILLER_21_2612 ();
 sg13g2_decap_8 FILLER_21_2644 ();
 sg13g2_decap_8 FILLER_21_2651 ();
 sg13g2_decap_8 FILLER_21_2658 ();
 sg13g2_decap_8 FILLER_21_2665 ();
 sg13g2_fill_2 FILLER_21_2672 ();
 sg13g2_fill_1 FILLER_22_69 ();
 sg13g2_fill_2 FILLER_22_111 ();
 sg13g2_fill_1 FILLER_22_118 ();
 sg13g2_fill_1 FILLER_22_149 ();
 sg13g2_fill_2 FILLER_22_170 ();
 sg13g2_fill_2 FILLER_22_219 ();
 sg13g2_fill_2 FILLER_22_247 ();
 sg13g2_fill_2 FILLER_22_254 ();
 sg13g2_fill_1 FILLER_22_390 ();
 sg13g2_fill_1 FILLER_22_411 ();
 sg13g2_fill_1 FILLER_22_523 ();
 sg13g2_fill_1 FILLER_22_539 ();
 sg13g2_fill_2 FILLER_22_576 ();
 sg13g2_fill_1 FILLER_22_578 ();
 sg13g2_fill_2 FILLER_22_584 ();
 sg13g2_fill_2 FILLER_22_595 ();
 sg13g2_fill_1 FILLER_22_597 ();
 sg13g2_fill_1 FILLER_22_608 ();
 sg13g2_fill_2 FILLER_22_630 ();
 sg13g2_fill_1 FILLER_22_650 ();
 sg13g2_fill_2 FILLER_22_677 ();
 sg13g2_fill_1 FILLER_22_687 ();
 sg13g2_fill_2 FILLER_22_723 ();
 sg13g2_fill_1 FILLER_22_725 ();
 sg13g2_fill_1 FILLER_22_731 ();
 sg13g2_fill_2 FILLER_22_749 ();
 sg13g2_fill_1 FILLER_22_751 ();
 sg13g2_fill_1 FILLER_22_794 ();
 sg13g2_fill_2 FILLER_22_839 ();
 sg13g2_fill_2 FILLER_22_932 ();
 sg13g2_fill_1 FILLER_22_934 ();
 sg13g2_fill_1 FILLER_22_943 ();
 sg13g2_fill_2 FILLER_22_1032 ();
 sg13g2_fill_1 FILLER_22_1034 ();
 sg13g2_fill_1 FILLER_22_1089 ();
 sg13g2_fill_2 FILLER_22_1099 ();
 sg13g2_fill_1 FILLER_22_1101 ();
 sg13g2_fill_2 FILLER_22_1234 ();
 sg13g2_fill_1 FILLER_22_1293 ();
 sg13g2_decap_4 FILLER_22_1310 ();
 sg13g2_fill_2 FILLER_22_1337 ();
 sg13g2_fill_1 FILLER_22_1339 ();
 sg13g2_fill_1 FILLER_22_1348 ();
 sg13g2_fill_2 FILLER_22_1365 ();
 sg13g2_fill_2 FILLER_22_1379 ();
 sg13g2_fill_2 FILLER_22_1400 ();
 sg13g2_fill_1 FILLER_22_1402 ();
 sg13g2_fill_2 FILLER_22_1416 ();
 sg13g2_fill_1 FILLER_22_1423 ();
 sg13g2_fill_2 FILLER_22_1430 ();
 sg13g2_fill_1 FILLER_22_1432 ();
 sg13g2_decap_4 FILLER_22_1441 ();
 sg13g2_fill_2 FILLER_22_1445 ();
 sg13g2_decap_8 FILLER_22_1453 ();
 sg13g2_fill_2 FILLER_22_1460 ();
 sg13g2_decap_8 FILLER_22_1474 ();
 sg13g2_decap_4 FILLER_22_1481 ();
 sg13g2_fill_1 FILLER_22_1485 ();
 sg13g2_decap_8 FILLER_22_1515 ();
 sg13g2_decap_4 FILLER_22_1522 ();
 sg13g2_fill_2 FILLER_22_1526 ();
 sg13g2_fill_2 FILLER_22_1544 ();
 sg13g2_fill_2 FILLER_22_1559 ();
 sg13g2_fill_2 FILLER_22_1587 ();
 sg13g2_fill_2 FILLER_22_1597 ();
 sg13g2_fill_1 FILLER_22_1599 ();
 sg13g2_fill_2 FILLER_22_1617 ();
 sg13g2_fill_1 FILLER_22_1619 ();
 sg13g2_fill_1 FILLER_22_1624 ();
 sg13g2_fill_1 FILLER_22_1679 ();
 sg13g2_fill_1 FILLER_22_1703 ();
 sg13g2_fill_2 FILLER_22_1731 ();
 sg13g2_fill_1 FILLER_22_1733 ();
 sg13g2_fill_2 FILLER_22_1794 ();
 sg13g2_fill_1 FILLER_22_1796 ();
 sg13g2_decap_8 FILLER_22_1881 ();
 sg13g2_fill_2 FILLER_22_1888 ();
 sg13g2_fill_2 FILLER_22_1925 ();
 sg13g2_fill_1 FILLER_22_1927 ();
 sg13g2_fill_2 FILLER_22_1971 ();
 sg13g2_fill_2 FILLER_22_2023 ();
 sg13g2_fill_2 FILLER_22_2051 ();
 sg13g2_fill_1 FILLER_22_2088 ();
 sg13g2_fill_2 FILLER_22_2195 ();
 sg13g2_fill_1 FILLER_22_2197 ();
 sg13g2_fill_2 FILLER_22_2319 ();
 sg13g2_fill_2 FILLER_22_2372 ();
 sg13g2_fill_2 FILLER_22_2400 ();
 sg13g2_fill_1 FILLER_22_2402 ();
 sg13g2_fill_1 FILLER_22_2474 ();
 sg13g2_fill_1 FILLER_22_2480 ();
 sg13g2_fill_2 FILLER_22_2517 ();
 sg13g2_fill_1 FILLER_22_2540 ();
 sg13g2_fill_2 FILLER_22_2571 ();
 sg13g2_fill_2 FILLER_22_2592 ();
 sg13g2_decap_8 FILLER_22_2641 ();
 sg13g2_decap_8 FILLER_22_2648 ();
 sg13g2_decap_8 FILLER_22_2655 ();
 sg13g2_decap_8 FILLER_22_2662 ();
 sg13g2_decap_4 FILLER_22_2669 ();
 sg13g2_fill_1 FILLER_22_2673 ();
 sg13g2_fill_2 FILLER_23_30 ();
 sg13g2_fill_1 FILLER_23_49 ();
 sg13g2_fill_2 FILLER_23_59 ();
 sg13g2_fill_1 FILLER_23_61 ();
 sg13g2_fill_2 FILLER_23_95 ();
 sg13g2_fill_1 FILLER_23_113 ();
 sg13g2_fill_2 FILLER_23_136 ();
 sg13g2_fill_2 FILLER_23_171 ();
 sg13g2_fill_1 FILLER_23_173 ();
 sg13g2_fill_1 FILLER_23_238 ();
 sg13g2_fill_2 FILLER_23_264 ();
 sg13g2_fill_1 FILLER_23_266 ();
 sg13g2_fill_1 FILLER_23_417 ();
 sg13g2_fill_1 FILLER_23_427 ();
 sg13g2_fill_1 FILLER_23_447 ();
 sg13g2_fill_1 FILLER_23_458 ();
 sg13g2_fill_2 FILLER_23_474 ();
 sg13g2_fill_1 FILLER_23_476 ();
 sg13g2_fill_1 FILLER_23_511 ();
 sg13g2_fill_2 FILLER_23_544 ();
 sg13g2_fill_1 FILLER_23_551 ();
 sg13g2_fill_1 FILLER_23_569 ();
 sg13g2_fill_2 FILLER_23_612 ();
 sg13g2_fill_1 FILLER_23_658 ();
 sg13g2_fill_1 FILLER_23_720 ();
 sg13g2_fill_1 FILLER_23_747 ();
 sg13g2_fill_1 FILLER_23_780 ();
 sg13g2_fill_2 FILLER_23_807 ();
 sg13g2_fill_2 FILLER_23_851 ();
 sg13g2_fill_1 FILLER_23_881 ();
 sg13g2_fill_1 FILLER_23_924 ();
 sg13g2_fill_1 FILLER_23_976 ();
 sg13g2_fill_1 FILLER_23_1003 ();
 sg13g2_fill_2 FILLER_23_1019 ();
 sg13g2_fill_1 FILLER_23_1041 ();
 sg13g2_fill_1 FILLER_23_1116 ();
 sg13g2_fill_2 FILLER_23_1127 ();
 sg13g2_fill_2 FILLER_23_1174 ();
 sg13g2_fill_1 FILLER_23_1176 ();
 sg13g2_fill_1 FILLER_23_1190 ();
 sg13g2_fill_2 FILLER_23_1209 ();
 sg13g2_fill_2 FILLER_23_1227 ();
 sg13g2_fill_1 FILLER_23_1229 ();
 sg13g2_fill_2 FILLER_23_1236 ();
 sg13g2_fill_2 FILLER_23_1279 ();
 sg13g2_fill_1 FILLER_23_1281 ();
 sg13g2_fill_1 FILLER_23_1300 ();
 sg13g2_fill_2 FILLER_23_1324 ();
 sg13g2_decap_4 FILLER_23_1391 ();
 sg13g2_fill_1 FILLER_23_1395 ();
 sg13g2_fill_2 FILLER_23_1420 ();
 sg13g2_fill_2 FILLER_23_1430 ();
 sg13g2_decap_4 FILLER_23_1444 ();
 sg13g2_fill_1 FILLER_23_1448 ();
 sg13g2_fill_2 FILLER_23_1522 ();
 sg13g2_fill_2 FILLER_23_1549 ();
 sg13g2_fill_2 FILLER_23_1556 ();
 sg13g2_fill_1 FILLER_23_1558 ();
 sg13g2_fill_2 FILLER_23_1564 ();
 sg13g2_fill_2 FILLER_23_1640 ();
 sg13g2_fill_2 FILLER_23_1662 ();
 sg13g2_fill_2 FILLER_23_1707 ();
 sg13g2_fill_1 FILLER_23_1766 ();
 sg13g2_fill_1 FILLER_23_1865 ();
 sg13g2_decap_4 FILLER_23_1893 ();
 sg13g2_fill_2 FILLER_23_2028 ();
 sg13g2_fill_2 FILLER_23_2047 ();
 sg13g2_fill_1 FILLER_23_2049 ();
 sg13g2_fill_2 FILLER_23_2069 ();
 sg13g2_fill_1 FILLER_23_2071 ();
 sg13g2_fill_2 FILLER_23_2080 ();
 sg13g2_fill_1 FILLER_23_2082 ();
 sg13g2_fill_1 FILLER_23_2091 ();
 sg13g2_fill_2 FILLER_23_2118 ();
 sg13g2_fill_1 FILLER_23_2138 ();
 sg13g2_fill_2 FILLER_23_2169 ();
 sg13g2_fill_2 FILLER_23_2240 ();
 sg13g2_fill_1 FILLER_23_2242 ();
 sg13g2_fill_2 FILLER_23_2292 ();
 sg13g2_fill_2 FILLER_23_2356 ();
 sg13g2_fill_1 FILLER_23_2358 ();
 sg13g2_fill_1 FILLER_23_2393 ();
 sg13g2_fill_2 FILLER_23_2404 ();
 sg13g2_fill_1 FILLER_23_2406 ();
 sg13g2_fill_1 FILLER_23_2426 ();
 sg13g2_fill_1 FILLER_23_2469 ();
 sg13g2_fill_1 FILLER_23_2530 ();
 sg13g2_decap_8 FILLER_23_2651 ();
 sg13g2_decap_8 FILLER_23_2658 ();
 sg13g2_decap_8 FILLER_23_2665 ();
 sg13g2_fill_2 FILLER_23_2672 ();
 sg13g2_fill_2 FILLER_24_48 ();
 sg13g2_fill_2 FILLER_24_134 ();
 sg13g2_fill_1 FILLER_24_201 ();
 sg13g2_fill_2 FILLER_24_224 ();
 sg13g2_fill_2 FILLER_24_252 ();
 sg13g2_fill_2 FILLER_24_260 ();
 sg13g2_fill_1 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_282 ();
 sg13g2_fill_1 FILLER_24_313 ();
 sg13g2_fill_1 FILLER_24_363 ();
 sg13g2_fill_2 FILLER_24_399 ();
 sg13g2_fill_1 FILLER_24_401 ();
 sg13g2_fill_2 FILLER_24_438 ();
 sg13g2_fill_1 FILLER_24_440 ();
 sg13g2_fill_2 FILLER_24_486 ();
 sg13g2_fill_1 FILLER_24_488 ();
 sg13g2_fill_1 FILLER_24_501 ();
 sg13g2_fill_2 FILLER_24_536 ();
 sg13g2_fill_1 FILLER_24_538 ();
 sg13g2_fill_1 FILLER_24_551 ();
 sg13g2_fill_1 FILLER_24_597 ();
 sg13g2_fill_2 FILLER_24_623 ();
 sg13g2_fill_1 FILLER_24_692 ();
 sg13g2_fill_2 FILLER_24_725 ();
 sg13g2_fill_2 FILLER_24_735 ();
 sg13g2_fill_1 FILLER_24_737 ();
 sg13g2_fill_2 FILLER_24_790 ();
 sg13g2_fill_1 FILLER_24_792 ();
 sg13g2_fill_2 FILLER_24_842 ();
 sg13g2_fill_2 FILLER_24_889 ();
 sg13g2_fill_1 FILLER_24_891 ();
 sg13g2_fill_2 FILLER_24_928 ();
 sg13g2_fill_2 FILLER_24_936 ();
 sg13g2_fill_1 FILLER_24_938 ();
 sg13g2_fill_2 FILLER_24_974 ();
 sg13g2_fill_2 FILLER_24_986 ();
 sg13g2_fill_2 FILLER_24_1016 ();
 sg13g2_fill_1 FILLER_24_1018 ();
 sg13g2_fill_1 FILLER_24_1068 ();
 sg13g2_fill_2 FILLER_24_1082 ();
 sg13g2_fill_2 FILLER_24_1102 ();
 sg13g2_fill_1 FILLER_24_1104 ();
 sg13g2_fill_2 FILLER_24_1110 ();
 sg13g2_fill_2 FILLER_24_1156 ();
 sg13g2_fill_2 FILLER_24_1240 ();
 sg13g2_fill_1 FILLER_24_1242 ();
 sg13g2_decap_8 FILLER_24_1288 ();
 sg13g2_decap_4 FILLER_24_1295 ();
 sg13g2_fill_1 FILLER_24_1299 ();
 sg13g2_decap_4 FILLER_24_1304 ();
 sg13g2_decap_4 FILLER_24_1346 ();
 sg13g2_fill_2 FILLER_24_1350 ();
 sg13g2_fill_2 FILLER_24_1365 ();
 sg13g2_fill_2 FILLER_24_1389 ();
 sg13g2_fill_1 FILLER_24_1391 ();
 sg13g2_fill_1 FILLER_24_1412 ();
 sg13g2_decap_8 FILLER_24_1446 ();
 sg13g2_fill_1 FILLER_24_1453 ();
 sg13g2_decap_8 FILLER_24_1478 ();
 sg13g2_decap_4 FILLER_24_1485 ();
 sg13g2_fill_2 FILLER_24_1503 ();
 sg13g2_fill_2 FILLER_24_1542 ();
 sg13g2_fill_1 FILLER_24_1544 ();
 sg13g2_fill_1 FILLER_24_1559 ();
 sg13g2_fill_2 FILLER_24_1583 ();
 sg13g2_fill_1 FILLER_24_1585 ();
 sg13g2_fill_1 FILLER_24_1592 ();
 sg13g2_fill_1 FILLER_24_1606 ();
 sg13g2_fill_1 FILLER_24_1620 ();
 sg13g2_fill_2 FILLER_24_1647 ();
 sg13g2_fill_1 FILLER_24_1649 ();
 sg13g2_fill_1 FILLER_24_1744 ();
 sg13g2_fill_2 FILLER_24_1812 ();
 sg13g2_fill_2 FILLER_24_1822 ();
 sg13g2_fill_2 FILLER_24_1830 ();
 sg13g2_fill_1 FILLER_24_1840 ();
 sg13g2_decap_4 FILLER_24_1870 ();
 sg13g2_fill_1 FILLER_24_1874 ();
 sg13g2_fill_2 FILLER_24_1890 ();
 sg13g2_fill_1 FILLER_24_1905 ();
 sg13g2_fill_2 FILLER_24_1969 ();
 sg13g2_fill_1 FILLER_24_1971 ();
 sg13g2_fill_1 FILLER_24_2080 ();
 sg13g2_fill_2 FILLER_24_2185 ();
 sg13g2_fill_1 FILLER_24_2313 ();
 sg13g2_fill_1 FILLER_24_2335 ();
 sg13g2_fill_1 FILLER_24_2380 ();
 sg13g2_fill_1 FILLER_24_2439 ();
 sg13g2_fill_1 FILLER_24_2475 ();
 sg13g2_fill_1 FILLER_24_2495 ();
 sg13g2_fill_2 FILLER_24_2548 ();
 sg13g2_fill_1 FILLER_24_2550 ();
 sg13g2_fill_1 FILLER_24_2576 ();
 sg13g2_fill_1 FILLER_24_2582 ();
 sg13g2_fill_1 FILLER_24_2588 ();
 sg13g2_fill_2 FILLER_24_2598 ();
 sg13g2_fill_1 FILLER_24_2600 ();
 sg13g2_fill_1 FILLER_24_2611 ();
 sg13g2_decap_8 FILLER_24_2646 ();
 sg13g2_decap_8 FILLER_24_2653 ();
 sg13g2_decap_8 FILLER_24_2660 ();
 sg13g2_decap_8 FILLER_24_2667 ();
 sg13g2_fill_1 FILLER_25_49 ();
 sg13g2_fill_2 FILLER_25_67 ();
 sg13g2_fill_2 FILLER_25_105 ();
 sg13g2_fill_1 FILLER_25_145 ();
 sg13g2_fill_1 FILLER_25_156 ();
 sg13g2_fill_2 FILLER_25_181 ();
 sg13g2_fill_2 FILLER_25_200 ();
 sg13g2_fill_2 FILLER_25_244 ();
 sg13g2_fill_1 FILLER_25_294 ();
 sg13g2_fill_1 FILLER_25_335 ();
 sg13g2_fill_2 FILLER_25_412 ();
 sg13g2_fill_2 FILLER_25_433 ();
 sg13g2_fill_1 FILLER_25_435 ();
 sg13g2_fill_1 FILLER_25_442 ();
 sg13g2_fill_2 FILLER_25_461 ();
 sg13g2_fill_2 FILLER_25_495 ();
 sg13g2_fill_1 FILLER_25_497 ();
 sg13g2_fill_2 FILLER_25_524 ();
 sg13g2_fill_1 FILLER_25_526 ();
 sg13g2_fill_2 FILLER_25_563 ();
 sg13g2_fill_1 FILLER_25_565 ();
 sg13g2_fill_1 FILLER_25_620 ();
 sg13g2_fill_2 FILLER_25_635 ();
 sg13g2_fill_1 FILLER_25_747 ();
 sg13g2_fill_2 FILLER_25_759 ();
 sg13g2_fill_1 FILLER_25_836 ();
 sg13g2_fill_2 FILLER_25_863 ();
 sg13g2_fill_1 FILLER_25_865 ();
 sg13g2_fill_1 FILLER_25_902 ();
 sg13g2_fill_2 FILLER_25_917 ();
 sg13g2_fill_1 FILLER_25_919 ();
 sg13g2_fill_2 FILLER_25_929 ();
 sg13g2_fill_2 FILLER_25_936 ();
 sg13g2_fill_1 FILLER_25_938 ();
 sg13g2_fill_1 FILLER_25_959 ();
 sg13g2_fill_2 FILLER_25_977 ();
 sg13g2_fill_1 FILLER_25_979 ();
 sg13g2_fill_2 FILLER_25_1052 ();
 sg13g2_fill_1 FILLER_25_1054 ();
 sg13g2_fill_1 FILLER_25_1137 ();
 sg13g2_fill_1 FILLER_25_1178 ();
 sg13g2_fill_2 FILLER_25_1221 ();
 sg13g2_fill_1 FILLER_25_1223 ();
 sg13g2_fill_1 FILLER_25_1238 ();
 sg13g2_fill_2 FILLER_25_1247 ();
 sg13g2_fill_1 FILLER_25_1249 ();
 sg13g2_fill_2 FILLER_25_1267 ();
 sg13g2_fill_1 FILLER_25_1269 ();
 sg13g2_fill_2 FILLER_25_1276 ();
 sg13g2_fill_1 FILLER_25_1278 ();
 sg13g2_fill_1 FILLER_25_1299 ();
 sg13g2_decap_8 FILLER_25_1312 ();
 sg13g2_decap_8 FILLER_25_1319 ();
 sg13g2_fill_1 FILLER_25_1326 ();
 sg13g2_decap_8 FILLER_25_1337 ();
 sg13g2_fill_2 FILLER_25_1344 ();
 sg13g2_fill_2 FILLER_25_1381 ();
 sg13g2_fill_1 FILLER_25_1399 ();
 sg13g2_fill_1 FILLER_25_1426 ();
 sg13g2_decap_4 FILLER_25_1441 ();
 sg13g2_fill_1 FILLER_25_1457 ();
 sg13g2_fill_1 FILLER_25_1461 ();
 sg13g2_fill_1 FILLER_25_1483 ();
 sg13g2_fill_1 FILLER_25_1497 ();
 sg13g2_fill_2 FILLER_25_1502 ();
 sg13g2_fill_1 FILLER_25_1504 ();
 sg13g2_decap_4 FILLER_25_1521 ();
 sg13g2_fill_2 FILLER_25_1545 ();
 sg13g2_fill_1 FILLER_25_1547 ();
 sg13g2_fill_2 FILLER_25_1596 ();
 sg13g2_fill_1 FILLER_25_1598 ();
 sg13g2_fill_2 FILLER_25_1607 ();
 sg13g2_fill_1 FILLER_25_1609 ();
 sg13g2_fill_2 FILLER_25_1618 ();
 sg13g2_fill_1 FILLER_25_1620 ();
 sg13g2_fill_2 FILLER_25_1630 ();
 sg13g2_fill_1 FILLER_25_1632 ();
 sg13g2_fill_1 FILLER_25_1659 ();
 sg13g2_fill_1 FILLER_25_1665 ();
 sg13g2_fill_1 FILLER_25_1729 ();
 sg13g2_fill_1 FILLER_25_1760 ();
 sg13g2_fill_1 FILLER_25_1767 ();
 sg13g2_decap_4 FILLER_25_1827 ();
 sg13g2_fill_1 FILLER_25_1831 ();
 sg13g2_fill_2 FILLER_25_1873 ();
 sg13g2_fill_1 FILLER_25_1891 ();
 sg13g2_fill_2 FILLER_25_1937 ();
 sg13g2_fill_1 FILLER_25_1939 ();
 sg13g2_fill_2 FILLER_25_1970 ();
 sg13g2_fill_1 FILLER_25_1972 ();
 sg13g2_fill_1 FILLER_25_2072 ();
 sg13g2_fill_1 FILLER_25_2160 ();
 sg13g2_fill_1 FILLER_25_2171 ();
 sg13g2_fill_1 FILLER_25_2198 ();
 sg13g2_fill_1 FILLER_25_2204 ();
 sg13g2_fill_2 FILLER_25_2222 ();
 sg13g2_fill_2 FILLER_25_2232 ();
 sg13g2_fill_1 FILLER_25_2254 ();
 sg13g2_fill_2 FILLER_25_2263 ();
 sg13g2_fill_1 FILLER_25_2265 ();
 sg13g2_fill_2 FILLER_25_2281 ();
 sg13g2_fill_1 FILLER_25_2304 ();
 sg13g2_fill_1 FILLER_25_2388 ();
 sg13g2_fill_2 FILLER_25_2399 ();
 sg13g2_fill_1 FILLER_25_2401 ();
 sg13g2_fill_1 FILLER_25_2453 ();
 sg13g2_fill_1 FILLER_25_2514 ();
 sg13g2_fill_2 FILLER_25_2596 ();
 sg13g2_decap_8 FILLER_25_2642 ();
 sg13g2_decap_8 FILLER_25_2649 ();
 sg13g2_decap_8 FILLER_25_2656 ();
 sg13g2_decap_8 FILLER_25_2663 ();
 sg13g2_decap_4 FILLER_25_2670 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_124 ();
 sg13g2_fill_2 FILLER_26_132 ();
 sg13g2_fill_2 FILLER_26_167 ();
 sg13g2_fill_1 FILLER_26_169 ();
 sg13g2_fill_2 FILLER_26_214 ();
 sg13g2_fill_1 FILLER_26_234 ();
 sg13g2_fill_1 FILLER_26_255 ();
 sg13g2_fill_1 FILLER_26_266 ();
 sg13g2_fill_2 FILLER_26_281 ();
 sg13g2_fill_1 FILLER_26_314 ();
 sg13g2_fill_2 FILLER_26_369 ();
 sg13g2_fill_1 FILLER_26_371 ();
 sg13g2_fill_2 FILLER_26_445 ();
 sg13g2_fill_2 FILLER_26_529 ();
 sg13g2_fill_1 FILLER_26_531 ();
 sg13g2_fill_2 FILLER_26_537 ();
 sg13g2_fill_2 FILLER_26_545 ();
 sg13g2_fill_2 FILLER_26_568 ();
 sg13g2_fill_1 FILLER_26_596 ();
 sg13g2_fill_2 FILLER_26_637 ();
 sg13g2_fill_1 FILLER_26_686 ();
 sg13g2_fill_2 FILLER_26_697 ();
 sg13g2_fill_2 FILLER_26_723 ();
 sg13g2_fill_1 FILLER_26_725 ();
 sg13g2_fill_1 FILLER_26_752 ();
 sg13g2_fill_1 FILLER_26_802 ();
 sg13g2_fill_1 FILLER_26_843 ();
 sg13g2_fill_1 FILLER_26_885 ();
 sg13g2_fill_1 FILLER_26_895 ();
 sg13g2_fill_2 FILLER_26_986 ();
 sg13g2_fill_2 FILLER_26_1005 ();
 sg13g2_fill_2 FILLER_26_1062 ();
 sg13g2_fill_1 FILLER_26_1064 ();
 sg13g2_fill_2 FILLER_26_1101 ();
 sg13g2_fill_1 FILLER_26_1116 ();
 sg13g2_fill_2 FILLER_26_1194 ();
 sg13g2_fill_1 FILLER_26_1206 ();
 sg13g2_fill_1 FILLER_26_1238 ();
 sg13g2_fill_1 FILLER_26_1270 ();
 sg13g2_fill_2 FILLER_26_1279 ();
 sg13g2_decap_8 FILLER_26_1301 ();
 sg13g2_decap_4 FILLER_26_1308 ();
 sg13g2_fill_1 FILLER_26_1312 ();
 sg13g2_decap_8 FILLER_26_1317 ();
 sg13g2_decap_4 FILLER_26_1324 ();
 sg13g2_fill_2 FILLER_26_1367 ();
 sg13g2_decap_4 FILLER_26_1377 ();
 sg13g2_fill_2 FILLER_26_1381 ();
 sg13g2_fill_2 FILLER_26_1391 ();
 sg13g2_fill_2 FILLER_26_1414 ();
 sg13g2_fill_1 FILLER_26_1438 ();
 sg13g2_decap_8 FILLER_26_1464 ();
 sg13g2_fill_2 FILLER_26_1471 ();
 sg13g2_fill_1 FILLER_26_1473 ();
 sg13g2_fill_1 FILLER_26_1499 ();
 sg13g2_fill_2 FILLER_26_1514 ();
 sg13g2_fill_1 FILLER_26_1516 ();
 sg13g2_fill_1 FILLER_26_1580 ();
 sg13g2_fill_1 FILLER_26_1589 ();
 sg13g2_fill_2 FILLER_26_1641 ();
 sg13g2_fill_1 FILLER_26_1643 ();
 sg13g2_decap_4 FILLER_26_1656 ();
 sg13g2_fill_1 FILLER_26_1660 ();
 sg13g2_fill_2 FILLER_26_1665 ();
 sg13g2_fill_2 FILLER_26_1722 ();
 sg13g2_fill_1 FILLER_26_1724 ();
 sg13g2_fill_1 FILLER_26_1787 ();
 sg13g2_fill_2 FILLER_26_1807 ();
 sg13g2_fill_1 FILLER_26_1809 ();
 sg13g2_fill_2 FILLER_26_1836 ();
 sg13g2_fill_1 FILLER_26_1838 ();
 sg13g2_decap_4 FILLER_26_1879 ();
 sg13g2_fill_2 FILLER_26_1909 ();
 sg13g2_fill_2 FILLER_26_1930 ();
 sg13g2_fill_2 FILLER_26_1959 ();
 sg13g2_fill_2 FILLER_26_2033 ();
 sg13g2_fill_1 FILLER_26_2035 ();
 sg13g2_fill_2 FILLER_26_2059 ();
 sg13g2_fill_1 FILLER_26_2061 ();
 sg13g2_fill_1 FILLER_26_2122 ();
 sg13g2_fill_1 FILLER_26_2198 ();
 sg13g2_fill_1 FILLER_26_2235 ();
 sg13g2_fill_2 FILLER_26_2245 ();
 sg13g2_fill_1 FILLER_26_2247 ();
 sg13g2_fill_1 FILLER_26_2274 ();
 sg13g2_fill_1 FILLER_26_2311 ();
 sg13g2_fill_1 FILLER_26_2328 ();
 sg13g2_fill_1 FILLER_26_2348 ();
 sg13g2_fill_2 FILLER_26_2359 ();
 sg13g2_fill_1 FILLER_26_2361 ();
 sg13g2_fill_2 FILLER_26_2376 ();
 sg13g2_fill_1 FILLER_26_2434 ();
 sg13g2_fill_2 FILLER_26_2463 ();
 sg13g2_fill_1 FILLER_26_2465 ();
 sg13g2_fill_2 FILLER_26_2484 ();
 sg13g2_fill_1 FILLER_26_2486 ();
 sg13g2_fill_2 FILLER_26_2502 ();
 sg13g2_fill_2 FILLER_26_2525 ();
 sg13g2_fill_1 FILLER_26_2527 ();
 sg13g2_fill_1 FILLER_26_2543 ();
 sg13g2_fill_2 FILLER_26_2574 ();
 sg13g2_fill_1 FILLER_26_2602 ();
 sg13g2_fill_1 FILLER_26_2613 ();
 sg13g2_decap_8 FILLER_26_2648 ();
 sg13g2_decap_8 FILLER_26_2655 ();
 sg13g2_decap_8 FILLER_26_2662 ();
 sg13g2_decap_4 FILLER_26_2669 ();
 sg13g2_fill_1 FILLER_26_2673 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_64 ();
 sg13g2_fill_1 FILLER_27_66 ();
 sg13g2_fill_2 FILLER_27_102 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_fill_1 FILLER_27_186 ();
 sg13g2_fill_2 FILLER_27_192 ();
 sg13g2_fill_1 FILLER_27_208 ();
 sg13g2_fill_2 FILLER_27_244 ();
 sg13g2_fill_1 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_321 ();
 sg13g2_fill_1 FILLER_27_348 ();
 sg13g2_fill_2 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_365 ();
 sg13g2_fill_1 FILLER_27_426 ();
 sg13g2_fill_2 FILLER_27_450 ();
 sg13g2_fill_1 FILLER_27_452 ();
 sg13g2_fill_2 FILLER_27_470 ();
 sg13g2_fill_1 FILLER_27_472 ();
 sg13g2_fill_2 FILLER_27_488 ();
 sg13g2_fill_1 FILLER_27_490 ();
 sg13g2_fill_2 FILLER_27_499 ();
 sg13g2_fill_1 FILLER_27_501 ();
 sg13g2_fill_2 FILLER_27_523 ();
 sg13g2_fill_1 FILLER_27_525 ();
 sg13g2_fill_2 FILLER_27_570 ();
 sg13g2_fill_1 FILLER_27_577 ();
 sg13g2_fill_1 FILLER_27_729 ();
 sg13g2_fill_1 FILLER_27_755 ();
 sg13g2_fill_2 FILLER_27_776 ();
 sg13g2_fill_1 FILLER_27_778 ();
 sg13g2_fill_2 FILLER_27_783 ();
 sg13g2_fill_2 FILLER_27_805 ();
 sg13g2_fill_1 FILLER_27_807 ();
 sg13g2_fill_1 FILLER_27_826 ();
 sg13g2_fill_1 FILLER_27_863 ();
 sg13g2_fill_2 FILLER_27_918 ();
 sg13g2_fill_2 FILLER_27_939 ();
 sg13g2_fill_2 FILLER_27_955 ();
 sg13g2_fill_1 FILLER_27_957 ();
 sg13g2_fill_1 FILLER_27_984 ();
 sg13g2_fill_2 FILLER_27_1030 ();
 sg13g2_fill_1 FILLER_27_1032 ();
 sg13g2_fill_2 FILLER_27_1158 ();
 sg13g2_fill_2 FILLER_27_1173 ();
 sg13g2_fill_1 FILLER_27_1175 ();
 sg13g2_fill_1 FILLER_27_1190 ();
 sg13g2_fill_1 FILLER_27_1209 ();
 sg13g2_fill_1 FILLER_27_1290 ();
 sg13g2_fill_2 FILLER_27_1329 ();
 sg13g2_fill_2 FILLER_27_1340 ();
 sg13g2_fill_1 FILLER_27_1342 ();
 sg13g2_fill_2 FILLER_27_1349 ();
 sg13g2_fill_2 FILLER_27_1357 ();
 sg13g2_fill_1 FILLER_27_1359 ();
 sg13g2_fill_2 FILLER_27_1384 ();
 sg13g2_fill_1 FILLER_27_1386 ();
 sg13g2_fill_1 FILLER_27_1416 ();
 sg13g2_fill_1 FILLER_27_1422 ();
 sg13g2_decap_4 FILLER_27_1428 ();
 sg13g2_fill_1 FILLER_27_1432 ();
 sg13g2_decap_8 FILLER_27_1441 ();
 sg13g2_fill_2 FILLER_27_1448 ();
 sg13g2_fill_2 FILLER_27_1476 ();
 sg13g2_fill_1 FILLER_27_1478 ();
 sg13g2_fill_1 FILLER_27_1502 ();
 sg13g2_decap_4 FILLER_27_1535 ();
 sg13g2_fill_1 FILLER_27_1539 ();
 sg13g2_decap_4 FILLER_27_1564 ();
 sg13g2_fill_1 FILLER_27_1617 ();
 sg13g2_fill_2 FILLER_27_1635 ();
 sg13g2_fill_2 FILLER_27_1645 ();
 sg13g2_fill_1 FILLER_27_1647 ();
 sg13g2_fill_2 FILLER_27_1684 ();
 sg13g2_fill_1 FILLER_27_1765 ();
 sg13g2_fill_1 FILLER_27_1811 ();
 sg13g2_fill_2 FILLER_27_1885 ();
 sg13g2_fill_1 FILLER_27_1887 ();
 sg13g2_decap_4 FILLER_27_1936 ();
 sg13g2_fill_1 FILLER_27_1989 ();
 sg13g2_fill_2 FILLER_27_1999 ();
 sg13g2_fill_1 FILLER_27_2024 ();
 sg13g2_fill_1 FILLER_27_2051 ();
 sg13g2_fill_2 FILLER_27_2083 ();
 sg13g2_fill_1 FILLER_27_2085 ();
 sg13g2_fill_2 FILLER_27_2107 ();
 sg13g2_fill_1 FILLER_27_2109 ();
 sg13g2_fill_2 FILLER_27_2190 ();
 sg13g2_fill_1 FILLER_27_2212 ();
 sg13g2_fill_2 FILLER_27_2388 ();
 sg13g2_fill_1 FILLER_27_2390 ();
 sg13g2_decap_8 FILLER_27_2643 ();
 sg13g2_decap_8 FILLER_27_2650 ();
 sg13g2_decap_8 FILLER_27_2657 ();
 sg13g2_decap_8 FILLER_27_2664 ();
 sg13g2_fill_2 FILLER_27_2671 ();
 sg13g2_fill_1 FILLER_27_2673 ();
 sg13g2_fill_1 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_42 ();
 sg13g2_fill_2 FILLER_28_56 ();
 sg13g2_fill_2 FILLER_28_79 ();
 sg13g2_fill_1 FILLER_28_111 ();
 sg13g2_fill_2 FILLER_28_134 ();
 sg13g2_fill_1 FILLER_28_136 ();
 sg13g2_fill_2 FILLER_28_148 ();
 sg13g2_fill_2 FILLER_28_184 ();
 sg13g2_fill_2 FILLER_28_264 ();
 sg13g2_fill_1 FILLER_28_266 ();
 sg13g2_fill_1 FILLER_28_291 ();
 sg13g2_fill_1 FILLER_28_315 ();
 sg13g2_fill_1 FILLER_28_325 ();
 sg13g2_fill_2 FILLER_28_340 ();
 sg13g2_fill_1 FILLER_28_342 ();
 sg13g2_fill_1 FILLER_28_365 ();
 sg13g2_fill_2 FILLER_28_477 ();
 sg13g2_fill_1 FILLER_28_479 ();
 sg13g2_fill_1 FILLER_28_511 ();
 sg13g2_fill_1 FILLER_28_522 ();
 sg13g2_fill_1 FILLER_28_538 ();
 sg13g2_fill_2 FILLER_28_572 ();
 sg13g2_fill_2 FILLER_28_587 ();
 sg13g2_fill_2 FILLER_28_639 ();
 sg13g2_fill_1 FILLER_28_681 ();
 sg13g2_fill_1 FILLER_28_694 ();
 sg13g2_fill_1 FILLER_28_712 ();
 sg13g2_fill_1 FILLER_28_753 ();
 sg13g2_fill_2 FILLER_28_803 ();
 sg13g2_fill_1 FILLER_28_805 ();
 sg13g2_fill_2 FILLER_28_836 ();
 sg13g2_fill_1 FILLER_28_847 ();
 sg13g2_fill_2 FILLER_28_857 ();
 sg13g2_fill_1 FILLER_28_955 ();
 sg13g2_fill_1 FILLER_28_1037 ();
 sg13g2_fill_2 FILLER_28_1046 ();
 sg13g2_fill_1 FILLER_28_1048 ();
 sg13g2_fill_1 FILLER_28_1122 ();
 sg13g2_fill_2 FILLER_28_1145 ();
 sg13g2_fill_2 FILLER_28_1160 ();
 sg13g2_fill_1 FILLER_28_1214 ();
 sg13g2_decap_4 FILLER_28_1351 ();
 sg13g2_fill_2 FILLER_28_1355 ();
 sg13g2_decap_4 FILLER_28_1402 ();
 sg13g2_fill_2 FILLER_28_1414 ();
 sg13g2_fill_2 FILLER_28_1448 ();
 sg13g2_fill_1 FILLER_28_1450 ();
 sg13g2_fill_2 FILLER_28_1492 ();
 sg13g2_fill_1 FILLER_28_1504 ();
 sg13g2_fill_1 FILLER_28_1517 ();
 sg13g2_decap_4 FILLER_28_1540 ();
 sg13g2_fill_1 FILLER_28_1544 ();
 sg13g2_fill_1 FILLER_28_1576 ();
 sg13g2_fill_2 FILLER_28_1581 ();
 sg13g2_fill_1 FILLER_28_1583 ();
 sg13g2_fill_2 FILLER_28_1589 ();
 sg13g2_fill_1 FILLER_28_1591 ();
 sg13g2_fill_2 FILLER_28_1601 ();
 sg13g2_fill_2 FILLER_28_1661 ();
 sg13g2_fill_1 FILLER_28_1757 ();
 sg13g2_fill_2 FILLER_28_1825 ();
 sg13g2_fill_1 FILLER_28_1848 ();
 sg13g2_fill_2 FILLER_28_1920 ();
 sg13g2_fill_1 FILLER_28_1922 ();
 sg13g2_fill_2 FILLER_28_1928 ();
 sg13g2_fill_1 FILLER_28_1930 ();
 sg13g2_fill_2 FILLER_28_1972 ();
 sg13g2_fill_1 FILLER_28_2014 ();
 sg13g2_fill_1 FILLER_28_2050 ();
 sg13g2_fill_2 FILLER_28_2101 ();
 sg13g2_fill_2 FILLER_28_2181 ();
 sg13g2_fill_1 FILLER_28_2373 ();
 sg13g2_fill_2 FILLER_28_2412 ();
 sg13g2_fill_1 FILLER_28_2414 ();
 sg13g2_fill_2 FILLER_28_2424 ();
 sg13g2_fill_1 FILLER_28_2426 ();
 sg13g2_fill_2 FILLER_28_2447 ();
 sg13g2_fill_1 FILLER_28_2472 ();
 sg13g2_fill_1 FILLER_28_2506 ();
 sg13g2_fill_2 FILLER_28_2517 ();
 sg13g2_fill_1 FILLER_28_2519 ();
 sg13g2_fill_2 FILLER_28_2556 ();
 sg13g2_fill_1 FILLER_28_2558 ();
 sg13g2_fill_2 FILLER_28_2585 ();
 sg13g2_decap_8 FILLER_28_2645 ();
 sg13g2_decap_8 FILLER_28_2652 ();
 sg13g2_decap_8 FILLER_28_2659 ();
 sg13g2_decap_8 FILLER_28_2666 ();
 sg13g2_fill_1 FILLER_28_2673 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_1 FILLER_29_26 ();
 sg13g2_fill_2 FILLER_29_52 ();
 sg13g2_fill_1 FILLER_29_54 ();
 sg13g2_fill_1 FILLER_29_104 ();
 sg13g2_fill_2 FILLER_29_141 ();
 sg13g2_fill_1 FILLER_29_143 ();
 sg13g2_fill_2 FILLER_29_170 ();
 sg13g2_fill_2 FILLER_29_192 ();
 sg13g2_fill_1 FILLER_29_194 ();
 sg13g2_fill_2 FILLER_29_224 ();
 sg13g2_fill_2 FILLER_29_243 ();
 sg13g2_fill_2 FILLER_29_293 ();
 sg13g2_fill_2 FILLER_29_309 ();
 sg13g2_fill_1 FILLER_29_311 ();
 sg13g2_fill_1 FILLER_29_388 ();
 sg13g2_fill_1 FILLER_29_394 ();
 sg13g2_fill_1 FILLER_29_516 ();
 sg13g2_fill_1 FILLER_29_631 ();
 sg13g2_fill_2 FILLER_29_645 ();
 sg13g2_fill_2 FILLER_29_673 ();
 sg13g2_fill_2 FILLER_29_696 ();
 sg13g2_fill_1 FILLER_29_698 ();
 sg13g2_fill_2 FILLER_29_713 ();
 sg13g2_fill_1 FILLER_29_715 ();
 sg13g2_fill_1 FILLER_29_763 ();
 sg13g2_fill_2 FILLER_29_783 ();
 sg13g2_fill_1 FILLER_29_798 ();
 sg13g2_fill_2 FILLER_29_854 ();
 sg13g2_fill_1 FILLER_29_901 ();
 sg13g2_fill_1 FILLER_29_917 ();
 sg13g2_fill_2 FILLER_29_927 ();
 sg13g2_fill_1 FILLER_29_938 ();
 sg13g2_fill_2 FILLER_29_997 ();
 sg13g2_fill_1 FILLER_29_999 ();
 sg13g2_fill_2 FILLER_29_1015 ();
 sg13g2_fill_1 FILLER_29_1017 ();
 sg13g2_fill_1 FILLER_29_1028 ();
 sg13g2_fill_1 FILLER_29_1071 ();
 sg13g2_fill_1 FILLER_29_1082 ();
 sg13g2_fill_2 FILLER_29_1115 ();
 sg13g2_fill_2 FILLER_29_1153 ();
 sg13g2_fill_1 FILLER_29_1183 ();
 sg13g2_fill_1 FILLER_29_1203 ();
 sg13g2_fill_1 FILLER_29_1223 ();
 sg13g2_fill_1 FILLER_29_1248 ();
 sg13g2_fill_1 FILLER_29_1280 ();
 sg13g2_fill_1 FILLER_29_1296 ();
 sg13g2_fill_2 FILLER_29_1382 ();
 sg13g2_fill_1 FILLER_29_1384 ();
 sg13g2_fill_2 FILLER_29_1394 ();
 sg13g2_fill_1 FILLER_29_1396 ();
 sg13g2_fill_2 FILLER_29_1440 ();
 sg13g2_fill_2 FILLER_29_1460 ();
 sg13g2_decap_8 FILLER_29_1466 ();
 sg13g2_fill_1 FILLER_29_1473 ();
 sg13g2_decap_4 FILLER_29_1523 ();
 sg13g2_fill_1 FILLER_29_1527 ();
 sg13g2_decap_8 FILLER_29_1532 ();
 sg13g2_decap_4 FILLER_29_1539 ();
 sg13g2_fill_1 FILLER_29_1543 ();
 sg13g2_fill_2 FILLER_29_1581 ();
 sg13g2_fill_2 FILLER_29_1619 ();
 sg13g2_fill_1 FILLER_29_1663 ();
 sg13g2_fill_2 FILLER_29_1706 ();
 sg13g2_fill_1 FILLER_29_1708 ();
 sg13g2_fill_2 FILLER_29_1749 ();
 sg13g2_fill_1 FILLER_29_1751 ();
 sg13g2_fill_2 FILLER_29_1778 ();
 sg13g2_fill_1 FILLER_29_1810 ();
 sg13g2_fill_2 FILLER_29_1903 ();
 sg13g2_fill_1 FILLER_29_1905 ();
 sg13g2_fill_2 FILLER_29_1932 ();
 sg13g2_fill_1 FILLER_29_1934 ();
 sg13g2_fill_1 FILLER_29_1948 ();
 sg13g2_fill_2 FILLER_29_1967 ();
 sg13g2_fill_2 FILLER_29_1995 ();
 sg13g2_fill_2 FILLER_29_2028 ();
 sg13g2_fill_1 FILLER_29_2030 ();
 sg13g2_fill_2 FILLER_29_2040 ();
 sg13g2_fill_1 FILLER_29_2083 ();
 sg13g2_fill_1 FILLER_29_2110 ();
 sg13g2_fill_2 FILLER_29_2137 ();
 sg13g2_fill_2 FILLER_29_2165 ();
 sg13g2_fill_1 FILLER_29_2167 ();
 sg13g2_fill_1 FILLER_29_2202 ();
 sg13g2_fill_1 FILLER_29_2212 ();
 sg13g2_fill_1 FILLER_29_2273 ();
 sg13g2_fill_1 FILLER_29_2315 ();
 sg13g2_fill_1 FILLER_29_2361 ();
 sg13g2_fill_2 FILLER_29_2476 ();
 sg13g2_fill_2 FILLER_29_2496 ();
 sg13g2_fill_2 FILLER_29_2538 ();
 sg13g2_fill_1 FILLER_29_2540 ();
 sg13g2_fill_2 FILLER_29_2567 ();
 sg13g2_fill_1 FILLER_29_2569 ();
 sg13g2_fill_1 FILLER_29_2619 ();
 sg13g2_decap_8 FILLER_29_2641 ();
 sg13g2_decap_8 FILLER_29_2648 ();
 sg13g2_decap_8 FILLER_29_2655 ();
 sg13g2_decap_8 FILLER_29_2662 ();
 sg13g2_decap_4 FILLER_29_2669 ();
 sg13g2_fill_1 FILLER_29_2673 ();
 sg13g2_fill_1 FILLER_30_46 ();
 sg13g2_fill_1 FILLER_30_60 ();
 sg13g2_fill_2 FILLER_30_65 ();
 sg13g2_fill_1 FILLER_30_93 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_fill_1 FILLER_30_141 ();
 sg13g2_fill_2 FILLER_30_152 ();
 sg13g2_fill_2 FILLER_30_160 ();
 sg13g2_fill_2 FILLER_30_192 ();
 sg13g2_fill_2 FILLER_30_269 ();
 sg13g2_fill_1 FILLER_30_271 ();
 sg13g2_fill_2 FILLER_30_296 ();
 sg13g2_fill_2 FILLER_30_313 ();
 sg13g2_fill_1 FILLER_30_381 ();
 sg13g2_fill_1 FILLER_30_405 ();
 sg13g2_fill_2 FILLER_30_480 ();
 sg13g2_fill_1 FILLER_30_543 ();
 sg13g2_fill_2 FILLER_30_553 ();
 sg13g2_fill_2 FILLER_30_600 ();
 sg13g2_fill_1 FILLER_30_602 ();
 sg13g2_fill_1 FILLER_30_611 ();
 sg13g2_fill_1 FILLER_30_659 ();
 sg13g2_fill_1 FILLER_30_683 ();
 sg13g2_fill_1 FILLER_30_745 ();
 sg13g2_fill_1 FILLER_30_841 ();
 sg13g2_fill_1 FILLER_30_991 ();
 sg13g2_fill_2 FILLER_30_1040 ();
 sg13g2_fill_1 FILLER_30_1048 ();
 sg13g2_fill_2 FILLER_30_1102 ();
 sg13g2_fill_1 FILLER_30_1104 ();
 sg13g2_fill_2 FILLER_30_1146 ();
 sg13g2_fill_2 FILLER_30_1210 ();
 sg13g2_fill_2 FILLER_30_1258 ();
 sg13g2_fill_2 FILLER_30_1293 ();
 sg13g2_fill_1 FILLER_30_1295 ();
 sg13g2_fill_2 FILLER_30_1304 ();
 sg13g2_fill_1 FILLER_30_1340 ();
 sg13g2_fill_1 FILLER_30_1359 ();
 sg13g2_fill_1 FILLER_30_1372 ();
 sg13g2_fill_2 FILLER_30_1401 ();
 sg13g2_decap_8 FILLER_30_1408 ();
 sg13g2_fill_1 FILLER_30_1498 ();
 sg13g2_fill_2 FILLER_30_1515 ();
 sg13g2_fill_1 FILLER_30_1573 ();
 sg13g2_fill_2 FILLER_30_1588 ();
 sg13g2_fill_1 FILLER_30_1599 ();
 sg13g2_fill_1 FILLER_30_1693 ();
 sg13g2_fill_2 FILLER_30_1720 ();
 sg13g2_fill_1 FILLER_30_1722 ();
 sg13g2_fill_2 FILLER_30_1759 ();
 sg13g2_fill_1 FILLER_30_1761 ();
 sg13g2_fill_2 FILLER_30_1803 ();
 sg13g2_fill_1 FILLER_30_1805 ();
 sg13g2_fill_2 FILLER_30_1816 ();
 sg13g2_fill_1 FILLER_30_1827 ();
 sg13g2_fill_2 FILLER_30_1856 ();
 sg13g2_fill_2 FILLER_30_1887 ();
 sg13g2_fill_2 FILLER_30_1946 ();
 sg13g2_fill_1 FILLER_30_1948 ();
 sg13g2_fill_2 FILLER_30_1975 ();
 sg13g2_fill_2 FILLER_30_2055 ();
 sg13g2_fill_1 FILLER_30_2057 ();
 sg13g2_fill_2 FILLER_30_2067 ();
 sg13g2_fill_1 FILLER_30_2069 ();
 sg13g2_fill_2 FILLER_30_2085 ();
 sg13g2_fill_1 FILLER_30_2087 ();
 sg13g2_fill_1 FILLER_30_2101 ();
 sg13g2_fill_2 FILLER_30_2116 ();
 sg13g2_fill_1 FILLER_30_2118 ();
 sg13g2_fill_2 FILLER_30_2145 ();
 sg13g2_fill_1 FILLER_30_2147 ();
 sg13g2_fill_2 FILLER_30_2172 ();
 sg13g2_fill_2 FILLER_30_2225 ();
 sg13g2_fill_1 FILLER_30_2227 ();
 sg13g2_fill_1 FILLER_30_2343 ();
 sg13g2_fill_1 FILLER_30_2392 ();
 sg13g2_fill_1 FILLER_30_2411 ();
 sg13g2_fill_2 FILLER_30_2426 ();
 sg13g2_fill_1 FILLER_30_2428 ();
 sg13g2_fill_1 FILLER_30_2527 ();
 sg13g2_fill_2 FILLER_30_2564 ();
 sg13g2_fill_1 FILLER_30_2566 ();
 sg13g2_fill_2 FILLER_30_2587 ();
 sg13g2_decap_8 FILLER_30_2640 ();
 sg13g2_decap_8 FILLER_30_2647 ();
 sg13g2_decap_8 FILLER_30_2654 ();
 sg13g2_decap_8 FILLER_30_2661 ();
 sg13g2_decap_4 FILLER_30_2668 ();
 sg13g2_fill_2 FILLER_30_2672 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_18 ();
 sg13g2_fill_2 FILLER_31_62 ();
 sg13g2_fill_1 FILLER_31_64 ();
 sg13g2_decap_8 FILLER_31_82 ();
 sg13g2_fill_2 FILLER_31_89 ();
 sg13g2_fill_1 FILLER_31_106 ();
 sg13g2_fill_2 FILLER_31_115 ();
 sg13g2_fill_1 FILLER_31_158 ();
 sg13g2_fill_2 FILLER_31_184 ();
 sg13g2_fill_1 FILLER_31_191 ();
 sg13g2_fill_1 FILLER_31_212 ();
 sg13g2_fill_1 FILLER_31_276 ();
 sg13g2_fill_1 FILLER_31_287 ();
 sg13g2_fill_2 FILLER_31_384 ();
 sg13g2_fill_1 FILLER_31_386 ();
 sg13g2_fill_1 FILLER_31_417 ();
 sg13g2_fill_2 FILLER_31_483 ();
 sg13g2_fill_2 FILLER_31_508 ();
 sg13g2_fill_2 FILLER_31_516 ();
 sg13g2_fill_1 FILLER_31_518 ();
 sg13g2_fill_2 FILLER_31_535 ();
 sg13g2_fill_1 FILLER_31_537 ();
 sg13g2_fill_2 FILLER_31_604 ();
 sg13g2_fill_1 FILLER_31_606 ();
 sg13g2_fill_2 FILLER_31_641 ();
 sg13g2_fill_1 FILLER_31_643 ();
 sg13g2_fill_2 FILLER_31_696 ();
 sg13g2_fill_2 FILLER_31_710 ();
 sg13g2_fill_2 FILLER_31_743 ();
 sg13g2_fill_2 FILLER_31_777 ();
 sg13g2_fill_1 FILLER_31_814 ();
 sg13g2_fill_1 FILLER_31_841 ();
 sg13g2_fill_1 FILLER_31_865 ();
 sg13g2_fill_1 FILLER_31_892 ();
 sg13g2_fill_1 FILLER_31_905 ();
 sg13g2_fill_2 FILLER_31_915 ();
 sg13g2_fill_2 FILLER_31_927 ();
 sg13g2_fill_2 FILLER_31_935 ();
 sg13g2_fill_1 FILLER_31_942 ();
 sg13g2_fill_1 FILLER_31_1059 ();
 sg13g2_fill_2 FILLER_31_1079 ();
 sg13g2_fill_1 FILLER_31_1081 ();
 sg13g2_fill_1 FILLER_31_1091 ();
 sg13g2_fill_1 FILLER_31_1100 ();
 sg13g2_fill_1 FILLER_31_1132 ();
 sg13g2_fill_2 FILLER_31_1166 ();
 sg13g2_fill_1 FILLER_31_1173 ();
 sg13g2_fill_1 FILLER_31_1183 ();
 sg13g2_fill_2 FILLER_31_1194 ();
 sg13g2_fill_1 FILLER_31_1210 ();
 sg13g2_fill_1 FILLER_31_1258 ();
 sg13g2_fill_2 FILLER_31_1265 ();
 sg13g2_fill_1 FILLER_31_1297 ();
 sg13g2_fill_1 FILLER_31_1342 ();
 sg13g2_fill_1 FILLER_31_1348 ();
 sg13g2_fill_1 FILLER_31_1372 ();
 sg13g2_fill_2 FILLER_31_1384 ();
 sg13g2_fill_1 FILLER_31_1436 ();
 sg13g2_fill_1 FILLER_31_1441 ();
 sg13g2_decap_4 FILLER_31_1451 ();
 sg13g2_decap_8 FILLER_31_1468 ();
 sg13g2_fill_1 FILLER_31_1475 ();
 sg13g2_fill_2 FILLER_31_1503 ();
 sg13g2_fill_2 FILLER_31_1526 ();
 sg13g2_fill_1 FILLER_31_1528 ();
 sg13g2_fill_2 FILLER_31_1547 ();
 sg13g2_fill_1 FILLER_31_1549 ();
 sg13g2_fill_1 FILLER_31_1562 ();
 sg13g2_fill_2 FILLER_31_1577 ();
 sg13g2_decap_4 FILLER_31_1596 ();
 sg13g2_decap_4 FILLER_31_1636 ();
 sg13g2_fill_2 FILLER_31_1649 ();
 sg13g2_fill_1 FILLER_31_1651 ();
 sg13g2_fill_2 FILLER_31_1660 ();
 sg13g2_fill_1 FILLER_31_1662 ();
 sg13g2_fill_1 FILLER_31_1682 ();
 sg13g2_fill_2 FILLER_31_1704 ();
 sg13g2_fill_1 FILLER_31_1706 ();
 sg13g2_fill_2 FILLER_31_1717 ();
 sg13g2_fill_1 FILLER_31_1757 ();
 sg13g2_fill_2 FILLER_31_1798 ();
 sg13g2_fill_2 FILLER_31_1873 ();
 sg13g2_fill_2 FILLER_31_1905 ();
 sg13g2_fill_1 FILLER_31_1907 ();
 sg13g2_fill_2 FILLER_31_1943 ();
 sg13g2_fill_1 FILLER_31_1945 ();
 sg13g2_fill_2 FILLER_31_2004 ();
 sg13g2_fill_2 FILLER_31_2042 ();
 sg13g2_fill_1 FILLER_31_2044 ();
 sg13g2_fill_2 FILLER_31_2081 ();
 sg13g2_fill_2 FILLER_31_2218 ();
 sg13g2_fill_2 FILLER_31_2237 ();
 sg13g2_fill_1 FILLER_31_2288 ();
 sg13g2_fill_1 FILLER_31_2329 ();
 sg13g2_fill_1 FILLER_31_2479 ();
 sg13g2_fill_2 FILLER_31_2500 ();
 sg13g2_fill_2 FILLER_31_2599 ();
 sg13g2_fill_2 FILLER_31_2611 ();
 sg13g2_fill_1 FILLER_31_2613 ();
 sg13g2_decap_8 FILLER_31_2644 ();
 sg13g2_decap_8 FILLER_31_2651 ();
 sg13g2_decap_8 FILLER_31_2658 ();
 sg13g2_decap_8 FILLER_31_2665 ();
 sg13g2_fill_2 FILLER_31_2672 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_4 ();
 sg13g2_fill_1 FILLER_32_18 ();
 sg13g2_decap_4 FILLER_32_39 ();
 sg13g2_fill_2 FILLER_32_49 ();
 sg13g2_fill_1 FILLER_32_51 ();
 sg13g2_decap_8 FILLER_32_62 ();
 sg13g2_decap_8 FILLER_32_69 ();
 sg13g2_decap_4 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_120 ();
 sg13g2_fill_2 FILLER_32_132 ();
 sg13g2_fill_2 FILLER_32_197 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_fill_1 FILLER_32_218 ();
 sg13g2_fill_2 FILLER_32_245 ();
 sg13g2_fill_1 FILLER_32_247 ();
 sg13g2_fill_1 FILLER_32_255 ();
 sg13g2_fill_1 FILLER_32_266 ();
 sg13g2_fill_1 FILLER_32_324 ();
 sg13g2_fill_2 FILLER_32_334 ();
 sg13g2_fill_1 FILLER_32_336 ();
 sg13g2_fill_2 FILLER_32_345 ();
 sg13g2_fill_1 FILLER_32_371 ();
 sg13g2_fill_2 FILLER_32_434 ();
 sg13g2_fill_1 FILLER_32_436 ();
 sg13g2_fill_2 FILLER_32_462 ();
 sg13g2_fill_2 FILLER_32_490 ();
 sg13g2_fill_1 FILLER_32_492 ();
 sg13g2_fill_1 FILLER_32_519 ();
 sg13g2_fill_2 FILLER_32_561 ();
 sg13g2_fill_1 FILLER_32_563 ();
 sg13g2_fill_1 FILLER_32_641 ();
 sg13g2_fill_2 FILLER_32_661 ();
 sg13g2_fill_2 FILLER_32_721 ();
 sg13g2_fill_2 FILLER_32_737 ();
 sg13g2_fill_2 FILLER_32_749 ();
 sg13g2_fill_1 FILLER_32_751 ();
 sg13g2_fill_2 FILLER_32_779 ();
 sg13g2_fill_1 FILLER_32_794 ();
 sg13g2_fill_2 FILLER_32_807 ();
 sg13g2_fill_1 FILLER_32_809 ();
 sg13g2_fill_1 FILLER_32_876 ();
 sg13g2_fill_2 FILLER_32_966 ();
 sg13g2_fill_2 FILLER_32_1099 ();
 sg13g2_fill_1 FILLER_32_1111 ();
 sg13g2_fill_1 FILLER_32_1122 ();
 sg13g2_fill_1 FILLER_32_1221 ();
 sg13g2_fill_1 FILLER_32_1236 ();
 sg13g2_fill_1 FILLER_32_1256 ();
 sg13g2_fill_2 FILLER_32_1282 ();
 sg13g2_fill_2 FILLER_32_1293 ();
 sg13g2_fill_1 FILLER_32_1295 ();
 sg13g2_fill_2 FILLER_32_1305 ();
 sg13g2_fill_2 FILLER_32_1316 ();
 sg13g2_fill_1 FILLER_32_1318 ();
 sg13g2_fill_2 FILLER_32_1326 ();
 sg13g2_fill_1 FILLER_32_1333 ();
 sg13g2_fill_2 FILLER_32_1339 ();
 sg13g2_fill_1 FILLER_32_1349 ();
 sg13g2_fill_2 FILLER_32_1400 ();
 sg13g2_fill_1 FILLER_32_1407 ();
 sg13g2_fill_1 FILLER_32_1425 ();
 sg13g2_decap_4 FILLER_32_1452 ();
 sg13g2_decap_4 FILLER_32_1496 ();
 sg13g2_fill_1 FILLER_32_1508 ();
 sg13g2_decap_8 FILLER_32_1529 ();
 sg13g2_decap_8 FILLER_32_1536 ();
 sg13g2_fill_1 FILLER_32_1543 ();
 sg13g2_decap_8 FILLER_32_1581 ();
 sg13g2_fill_1 FILLER_32_1588 ();
 sg13g2_decap_4 FILLER_32_1619 ();
 sg13g2_fill_2 FILLER_32_1720 ();
 sg13g2_fill_1 FILLER_32_1722 ();
 sg13g2_fill_2 FILLER_32_1735 ();
 sg13g2_fill_2 FILLER_32_1750 ();
 sg13g2_fill_1 FILLER_32_1752 ();
 sg13g2_fill_1 FILLER_32_1778 ();
 sg13g2_fill_2 FILLER_32_1789 ();
 sg13g2_fill_1 FILLER_32_1791 ();
 sg13g2_fill_1 FILLER_32_1863 ();
 sg13g2_fill_2 FILLER_32_1902 ();
 sg13g2_fill_1 FILLER_32_1962 ();
 sg13g2_fill_2 FILLER_32_1997 ();
 sg13g2_fill_1 FILLER_32_1999 ();
 sg13g2_fill_2 FILLER_32_2086 ();
 sg13g2_fill_1 FILLER_32_2088 ();
 sg13g2_fill_1 FILLER_32_2135 ();
 sg13g2_fill_1 FILLER_32_2146 ();
 sg13g2_fill_1 FILLER_32_2152 ();
 sg13g2_fill_2 FILLER_32_2181 ();
 sg13g2_fill_2 FILLER_32_2198 ();
 sg13g2_fill_2 FILLER_32_2263 ();
 sg13g2_fill_1 FILLER_32_2265 ();
 sg13g2_fill_2 FILLER_32_2285 ();
 sg13g2_fill_2 FILLER_32_2401 ();
 sg13g2_fill_1 FILLER_32_2403 ();
 sg13g2_fill_1 FILLER_32_2409 ();
 sg13g2_fill_1 FILLER_32_2513 ();
 sg13g2_fill_2 FILLER_32_2577 ();
 sg13g2_decap_8 FILLER_32_2655 ();
 sg13g2_decap_8 FILLER_32_2662 ();
 sg13g2_decap_4 FILLER_32_2669 ();
 sg13g2_fill_1 FILLER_32_2673 ();
 sg13g2_fill_2 FILLER_33_37 ();
 sg13g2_fill_2 FILLER_33_50 ();
 sg13g2_fill_1 FILLER_33_52 ();
 sg13g2_fill_1 FILLER_33_79 ();
 sg13g2_fill_1 FILLER_33_92 ();
 sg13g2_fill_1 FILLER_33_118 ();
 sg13g2_decap_4 FILLER_33_124 ();
 sg13g2_fill_2 FILLER_33_136 ();
 sg13g2_decap_4 FILLER_33_159 ();
 sg13g2_fill_1 FILLER_33_205 ();
 sg13g2_fill_1 FILLER_33_265 ();
 sg13g2_fill_2 FILLER_33_282 ();
 sg13g2_fill_1 FILLER_33_284 ();
 sg13g2_fill_1 FILLER_33_354 ();
 sg13g2_fill_2 FILLER_33_381 ();
 sg13g2_fill_1 FILLER_33_394 ();
 sg13g2_fill_2 FILLER_33_451 ();
 sg13g2_fill_1 FILLER_33_453 ();
 sg13g2_fill_1 FILLER_33_500 ();
 sg13g2_fill_2 FILLER_33_526 ();
 sg13g2_fill_2 FILLER_33_562 ();
 sg13g2_fill_1 FILLER_33_574 ();
 sg13g2_fill_2 FILLER_33_599 ();
 sg13g2_fill_1 FILLER_33_601 ();
 sg13g2_fill_2 FILLER_33_632 ();
 sg13g2_fill_2 FILLER_33_646 ();
 sg13g2_fill_1 FILLER_33_648 ();
 sg13g2_fill_2 FILLER_33_654 ();
 sg13g2_fill_2 FILLER_33_717 ();
 sg13g2_fill_2 FILLER_33_807 ();
 sg13g2_fill_1 FILLER_33_809 ();
 sg13g2_fill_2 FILLER_33_820 ();
 sg13g2_fill_1 FILLER_33_822 ();
 sg13g2_fill_2 FILLER_33_860 ();
 sg13g2_fill_1 FILLER_33_862 ();
 sg13g2_fill_2 FILLER_33_884 ();
 sg13g2_fill_1 FILLER_33_886 ();
 sg13g2_fill_2 FILLER_33_895 ();
 sg13g2_fill_1 FILLER_33_897 ();
 sg13g2_fill_2 FILLER_33_942 ();
 sg13g2_fill_1 FILLER_33_944 ();
 sg13g2_fill_1 FILLER_33_1001 ();
 sg13g2_fill_2 FILLER_33_1017 ();
 sg13g2_fill_2 FILLER_33_1146 ();
 sg13g2_fill_1 FILLER_33_1172 ();
 sg13g2_fill_2 FILLER_33_1288 ();
 sg13g2_fill_2 FILLER_33_1332 ();
 sg13g2_fill_2 FILLER_33_1340 ();
 sg13g2_fill_2 FILLER_33_1353 ();
 sg13g2_fill_1 FILLER_33_1359 ();
 sg13g2_fill_2 FILLER_33_1371 ();
 sg13g2_fill_2 FILLER_33_1378 ();
 sg13g2_decap_4 FILLER_33_1385 ();
 sg13g2_fill_2 FILLER_33_1389 ();
 sg13g2_decap_4 FILLER_33_1419 ();
 sg13g2_decap_8 FILLER_33_1463 ();
 sg13g2_decap_4 FILLER_33_1479 ();
 sg13g2_fill_1 FILLER_33_1514 ();
 sg13g2_fill_2 FILLER_33_1550 ();
 sg13g2_fill_2 FILLER_33_1636 ();
 sg13g2_fill_1 FILLER_33_1638 ();
 sg13g2_fill_1 FILLER_33_1652 ();
 sg13g2_fill_2 FILLER_33_1658 ();
 sg13g2_fill_2 FILLER_33_1739 ();
 sg13g2_fill_1 FILLER_33_1741 ();
 sg13g2_decap_8 FILLER_33_1763 ();
 sg13g2_fill_1 FILLER_33_1786 ();
 sg13g2_fill_2 FILLER_33_1792 ();
 sg13g2_fill_2 FILLER_33_1845 ();
 sg13g2_fill_1 FILLER_33_1847 ();
 sg13g2_fill_1 FILLER_33_1924 ();
 sg13g2_fill_1 FILLER_33_1953 ();
 sg13g2_decap_4 FILLER_33_1990 ();
 sg13g2_fill_2 FILLER_33_2030 ();
 sg13g2_fill_1 FILLER_33_2032 ();
 sg13g2_fill_2 FILLER_33_2065 ();
 sg13g2_fill_1 FILLER_33_2067 ();
 sg13g2_fill_1 FILLER_33_2105 ();
 sg13g2_fill_2 FILLER_33_2111 ();
 sg13g2_fill_2 FILLER_33_2139 ();
 sg13g2_fill_2 FILLER_33_2167 ();
 sg13g2_fill_2 FILLER_33_2174 ();
 sg13g2_fill_1 FILLER_33_2176 ();
 sg13g2_fill_1 FILLER_33_2208 ();
 sg13g2_fill_1 FILLER_33_2292 ();
 sg13g2_fill_2 FILLER_33_2355 ();
 sg13g2_fill_1 FILLER_33_2357 ();
 sg13g2_fill_2 FILLER_33_2373 ();
 sg13g2_fill_1 FILLER_33_2375 ();
 sg13g2_fill_1 FILLER_33_2412 ();
 sg13g2_fill_2 FILLER_33_2421 ();
 sg13g2_fill_2 FILLER_33_2483 ();
 sg13g2_fill_1 FILLER_33_2485 ();
 sg13g2_fill_2 FILLER_33_2565 ();
 sg13g2_fill_1 FILLER_33_2567 ();
 sg13g2_fill_2 FILLER_33_2608 ();
 sg13g2_decap_8 FILLER_33_2645 ();
 sg13g2_decap_8 FILLER_33_2652 ();
 sg13g2_decap_8 FILLER_33_2659 ();
 sg13g2_decap_8 FILLER_33_2666 ();
 sg13g2_fill_1 FILLER_33_2673 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_19 ();
 sg13g2_fill_1 FILLER_34_26 ();
 sg13g2_fill_1 FILLER_34_59 ();
 sg13g2_decap_4 FILLER_34_73 ();
 sg13g2_fill_1 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_108 ();
 sg13g2_fill_2 FILLER_34_147 ();
 sg13g2_fill_2 FILLER_34_165 ();
 sg13g2_fill_1 FILLER_34_167 ();
 sg13g2_fill_2 FILLER_34_193 ();
 sg13g2_fill_2 FILLER_34_209 ();
 sg13g2_fill_1 FILLER_34_258 ();
 sg13g2_fill_2 FILLER_34_270 ();
 sg13g2_fill_1 FILLER_34_284 ();
 sg13g2_fill_2 FILLER_34_296 ();
 sg13g2_fill_1 FILLER_34_298 ();
 sg13g2_fill_1 FILLER_34_309 ();
 sg13g2_fill_2 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_351 ();
 sg13g2_fill_2 FILLER_34_361 ();
 sg13g2_fill_1 FILLER_34_396 ();
 sg13g2_fill_2 FILLER_34_423 ();
 sg13g2_fill_2 FILLER_34_440 ();
 sg13g2_fill_1 FILLER_34_442 ();
 sg13g2_fill_2 FILLER_34_511 ();
 sg13g2_fill_1 FILLER_34_621 ();
 sg13g2_fill_2 FILLER_34_630 ();
 sg13g2_fill_2 FILLER_34_637 ();
 sg13g2_fill_1 FILLER_34_639 ();
 sg13g2_fill_2 FILLER_34_676 ();
 sg13g2_fill_1 FILLER_34_678 ();
 sg13g2_fill_2 FILLER_34_705 ();
 sg13g2_fill_1 FILLER_34_707 ();
 sg13g2_fill_2 FILLER_34_720 ();
 sg13g2_fill_2 FILLER_34_757 ();
 sg13g2_fill_1 FILLER_34_814 ();
 sg13g2_fill_2 FILLER_34_841 ();
 sg13g2_fill_1 FILLER_34_843 ();
 sg13g2_fill_1 FILLER_34_926 ();
 sg13g2_fill_1 FILLER_34_978 ();
 sg13g2_fill_2 FILLER_34_992 ();
 sg13g2_fill_1 FILLER_34_1002 ();
 sg13g2_fill_2 FILLER_34_1089 ();
 sg13g2_fill_1 FILLER_34_1105 ();
 sg13g2_fill_2 FILLER_34_1151 ();
 sg13g2_fill_1 FILLER_34_1153 ();
 sg13g2_fill_1 FILLER_34_1189 ();
 sg13g2_fill_1 FILLER_34_1207 ();
 sg13g2_fill_1 FILLER_34_1223 ();
 sg13g2_fill_1 FILLER_34_1233 ();
 sg13g2_fill_2 FILLER_34_1319 ();
 sg13g2_fill_2 FILLER_34_1329 ();
 sg13g2_fill_1 FILLER_34_1341 ();
 sg13g2_fill_2 FILLER_34_1410 ();
 sg13g2_fill_1 FILLER_34_1495 ();
 sg13g2_decap_8 FILLER_34_1502 ();
 sg13g2_decap_8 FILLER_34_1518 ();
 sg13g2_fill_1 FILLER_34_1525 ();
 sg13g2_decap_4 FILLER_34_1530 ();
 sg13g2_fill_1 FILLER_34_1534 ();
 sg13g2_fill_1 FILLER_34_1565 ();
 sg13g2_fill_1 FILLER_34_1589 ();
 sg13g2_fill_2 FILLER_34_1607 ();
 sg13g2_fill_1 FILLER_34_1640 ();
 sg13g2_fill_1 FILLER_34_1697 ();
 sg13g2_fill_1 FILLER_34_1721 ();
 sg13g2_fill_1 FILLER_34_1789 ();
 sg13g2_fill_2 FILLER_34_1859 ();
 sg13g2_fill_2 FILLER_34_1875 ();
 sg13g2_fill_2 FILLER_34_1898 ();
 sg13g2_fill_2 FILLER_34_1919 ();
 sg13g2_fill_1 FILLER_34_1921 ();
 sg13g2_fill_1 FILLER_34_1962 ();
 sg13g2_fill_2 FILLER_34_1986 ();
 sg13g2_fill_1 FILLER_34_2031 ();
 sg13g2_fill_1 FILLER_34_2058 ();
 sg13g2_fill_2 FILLER_34_2108 ();
 sg13g2_fill_2 FILLER_34_2150 ();
 sg13g2_fill_2 FILLER_34_2160 ();
 sg13g2_fill_2 FILLER_34_2206 ();
 sg13g2_fill_1 FILLER_34_2208 ();
 sg13g2_fill_1 FILLER_34_2227 ();
 sg13g2_fill_2 FILLER_34_2260 ();
 sg13g2_fill_2 FILLER_34_2285 ();
 sg13g2_fill_1 FILLER_34_2297 ();
 sg13g2_fill_2 FILLER_34_2336 ();
 sg13g2_fill_2 FILLER_34_2347 ();
 sg13g2_fill_1 FILLER_34_2372 ();
 sg13g2_fill_2 FILLER_34_2406 ();
 sg13g2_fill_1 FILLER_34_2408 ();
 sg13g2_fill_2 FILLER_34_2503 ();
 sg13g2_fill_2 FILLER_34_2522 ();
 sg13g2_fill_1 FILLER_34_2524 ();
 sg13g2_fill_2 FILLER_34_2555 ();
 sg13g2_fill_1 FILLER_34_2557 ();
 sg13g2_fill_2 FILLER_34_2578 ();
 sg13g2_decap_8 FILLER_34_2636 ();
 sg13g2_decap_8 FILLER_34_2643 ();
 sg13g2_decap_8 FILLER_34_2650 ();
 sg13g2_decap_8 FILLER_34_2657 ();
 sg13g2_decap_8 FILLER_34_2664 ();
 sg13g2_fill_2 FILLER_34_2671 ();
 sg13g2_fill_1 FILLER_34_2673 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_4 ();
 sg13g2_decap_4 FILLER_35_43 ();
 sg13g2_fill_2 FILLER_35_58 ();
 sg13g2_fill_2 FILLER_35_114 ();
 sg13g2_fill_1 FILLER_35_116 ();
 sg13g2_fill_2 FILLER_35_140 ();
 sg13g2_fill_1 FILLER_35_142 ();
 sg13g2_fill_2 FILLER_35_156 ();
 sg13g2_fill_1 FILLER_35_176 ();
 sg13g2_fill_2 FILLER_35_200 ();
 sg13g2_fill_2 FILLER_35_216 ();
 sg13g2_fill_1 FILLER_35_218 ();
 sg13g2_fill_2 FILLER_35_253 ();
 sg13g2_fill_1 FILLER_35_260 ();
 sg13g2_fill_2 FILLER_35_309 ();
 sg13g2_fill_1 FILLER_35_327 ();
 sg13g2_fill_1 FILLER_35_341 ();
 sg13g2_fill_2 FILLER_35_385 ();
 sg13g2_fill_2 FILLER_35_472 ();
 sg13g2_fill_1 FILLER_35_484 ();
 sg13g2_fill_2 FILLER_35_587 ();
 sg13g2_fill_1 FILLER_35_589 ();
 sg13g2_fill_2 FILLER_35_603 ();
 sg13g2_fill_1 FILLER_35_675 ();
 sg13g2_fill_1 FILLER_35_721 ();
 sg13g2_fill_1 FILLER_35_738 ();
 sg13g2_fill_1 FILLER_35_748 ();
 sg13g2_fill_2 FILLER_35_762 ();
 sg13g2_fill_1 FILLER_35_764 ();
 sg13g2_fill_1 FILLER_35_784 ();
 sg13g2_fill_2 FILLER_35_802 ();
 sg13g2_fill_1 FILLER_35_804 ();
 sg13g2_fill_2 FILLER_35_886 ();
 sg13g2_fill_1 FILLER_35_888 ();
 sg13g2_fill_1 FILLER_35_933 ();
 sg13g2_fill_2 FILLER_35_960 ();
 sg13g2_fill_2 FILLER_35_971 ();
 sg13g2_fill_1 FILLER_35_973 ();
 sg13g2_fill_1 FILLER_35_984 ();
 sg13g2_fill_2 FILLER_35_1000 ();
 sg13g2_fill_1 FILLER_35_1018 ();
 sg13g2_fill_2 FILLER_35_1038 ();
 sg13g2_fill_1 FILLER_35_1040 ();
 sg13g2_fill_1 FILLER_35_1065 ();
 sg13g2_fill_2 FILLER_35_1071 ();
 sg13g2_fill_1 FILLER_35_1073 ();
 sg13g2_fill_1 FILLER_35_1095 ();
 sg13g2_fill_2 FILLER_35_1125 ();
 sg13g2_fill_2 FILLER_35_1145 ();
 sg13g2_fill_1 FILLER_35_1147 ();
 sg13g2_decap_4 FILLER_35_1156 ();
 sg13g2_fill_2 FILLER_35_1169 ();
 sg13g2_fill_2 FILLER_35_1178 ();
 sg13g2_fill_2 FILLER_35_1206 ();
 sg13g2_fill_2 FILLER_35_1238 ();
 sg13g2_fill_1 FILLER_35_1240 ();
 sg13g2_fill_1 FILLER_35_1250 ();
 sg13g2_fill_2 FILLER_35_1256 ();
 sg13g2_fill_1 FILLER_35_1258 ();
 sg13g2_fill_2 FILLER_35_1290 ();
 sg13g2_fill_1 FILLER_35_1292 ();
 sg13g2_fill_1 FILLER_35_1326 ();
 sg13g2_fill_1 FILLER_35_1343 ();
 sg13g2_fill_2 FILLER_35_1359 ();
 sg13g2_fill_1 FILLER_35_1365 ();
 sg13g2_fill_2 FILLER_35_1374 ();
 sg13g2_fill_2 FILLER_35_1390 ();
 sg13g2_fill_1 FILLER_35_1392 ();
 sg13g2_fill_2 FILLER_35_1419 ();
 sg13g2_fill_1 FILLER_35_1421 ();
 sg13g2_fill_2 FILLER_35_1435 ();
 sg13g2_decap_8 FILLER_35_1456 ();
 sg13g2_fill_2 FILLER_35_1463 ();
 sg13g2_fill_1 FILLER_35_1465 ();
 sg13g2_decap_8 FILLER_35_1470 ();
 sg13g2_decap_4 FILLER_35_1508 ();
 sg13g2_decap_4 FILLER_35_1516 ();
 sg13g2_fill_1 FILLER_35_1520 ();
 sg13g2_decap_4 FILLER_35_1528 ();
 sg13g2_fill_1 FILLER_35_1532 ();
 sg13g2_decap_4 FILLER_35_1540 ();
 sg13g2_decap_4 FILLER_35_1555 ();
 sg13g2_fill_1 FILLER_35_1563 ();
 sg13g2_fill_2 FILLER_35_1577 ();
 sg13g2_fill_1 FILLER_35_1676 ();
 sg13g2_fill_2 FILLER_35_1702 ();
 sg13g2_fill_2 FILLER_35_1730 ();
 sg13g2_decap_4 FILLER_35_1772 ();
 sg13g2_fill_2 FILLER_35_1776 ();
 sg13g2_decap_8 FILLER_35_1786 ();
 sg13g2_fill_2 FILLER_35_1793 ();
 sg13g2_fill_1 FILLER_35_1868 ();
 sg13g2_fill_1 FILLER_35_1951 ();
 sg13g2_fill_2 FILLER_35_2024 ();
 sg13g2_fill_1 FILLER_35_2026 ();
 sg13g2_fill_2 FILLER_35_2041 ();
 sg13g2_fill_1 FILLER_35_2043 ();
 sg13g2_fill_1 FILLER_35_2069 ();
 sg13g2_fill_1 FILLER_35_2080 ();
 sg13g2_fill_1 FILLER_35_2097 ();
 sg13g2_fill_1 FILLER_35_2112 ();
 sg13g2_fill_1 FILLER_35_2193 ();
 sg13g2_fill_2 FILLER_35_2204 ();
 sg13g2_fill_1 FILLER_35_2206 ();
 sg13g2_fill_2 FILLER_35_2311 ();
 sg13g2_fill_1 FILLER_35_2313 ();
 sg13g2_fill_2 FILLER_35_2453 ();
 sg13g2_fill_2 FILLER_35_2599 ();
 sg13g2_fill_1 FILLER_35_2601 ();
 sg13g2_fill_1 FILLER_35_2620 ();
 sg13g2_decap_8 FILLER_35_2634 ();
 sg13g2_decap_8 FILLER_35_2641 ();
 sg13g2_decap_8 FILLER_35_2648 ();
 sg13g2_decap_8 FILLER_35_2655 ();
 sg13g2_decap_8 FILLER_35_2662 ();
 sg13g2_decap_4 FILLER_35_2669 ();
 sg13g2_fill_1 FILLER_35_2673 ();
 sg13g2_fill_1 FILLER_36_26 ();
 sg13g2_fill_2 FILLER_36_43 ();
 sg13g2_fill_1 FILLER_36_45 ();
 sg13g2_fill_1 FILLER_36_50 ();
 sg13g2_decap_4 FILLER_36_60 ();
 sg13g2_fill_1 FILLER_36_64 ();
 sg13g2_fill_1 FILLER_36_71 ();
 sg13g2_fill_2 FILLER_36_95 ();
 sg13g2_fill_1 FILLER_36_97 ();
 sg13g2_fill_2 FILLER_36_110 ();
 sg13g2_fill_2 FILLER_36_121 ();
 sg13g2_fill_1 FILLER_36_123 ();
 sg13g2_fill_1 FILLER_36_128 ();
 sg13g2_fill_2 FILLER_36_133 ();
 sg13g2_fill_1 FILLER_36_135 ();
 sg13g2_decap_4 FILLER_36_158 ();
 sg13g2_fill_2 FILLER_36_162 ();
 sg13g2_decap_8 FILLER_36_200 ();
 sg13g2_fill_1 FILLER_36_207 ();
 sg13g2_fill_2 FILLER_36_214 ();
 sg13g2_fill_2 FILLER_36_229 ();
 sg13g2_fill_1 FILLER_36_231 ();
 sg13g2_fill_2 FILLER_36_256 ();
 sg13g2_fill_2 FILLER_36_277 ();
 sg13g2_fill_1 FILLER_36_279 ();
 sg13g2_fill_2 FILLER_36_308 ();
 sg13g2_fill_2 FILLER_36_315 ();
 sg13g2_fill_1 FILLER_36_317 ();
 sg13g2_fill_2 FILLER_36_330 ();
 sg13g2_fill_1 FILLER_36_332 ();
 sg13g2_fill_2 FILLER_36_373 ();
 sg13g2_fill_2 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_413 ();
 sg13g2_fill_1 FILLER_36_445 ();
 sg13g2_fill_2 FILLER_36_478 ();
 sg13g2_fill_1 FILLER_36_521 ();
 sg13g2_fill_2 FILLER_36_616 ();
 sg13g2_fill_2 FILLER_36_645 ();
 sg13g2_fill_1 FILLER_36_647 ();
 sg13g2_fill_1 FILLER_36_674 ();
 sg13g2_fill_2 FILLER_36_740 ();
 sg13g2_fill_1 FILLER_36_742 ();
 sg13g2_fill_1 FILLER_36_782 ();
 sg13g2_fill_1 FILLER_36_809 ();
 sg13g2_fill_2 FILLER_36_820 ();
 sg13g2_fill_2 FILLER_36_866 ();
 sg13g2_fill_1 FILLER_36_868 ();
 sg13g2_fill_2 FILLER_36_956 ();
 sg13g2_fill_1 FILLER_36_958 ();
 sg13g2_fill_2 FILLER_36_1052 ();
 sg13g2_fill_1 FILLER_36_1054 ();
 sg13g2_fill_2 FILLER_36_1068 ();
 sg13g2_fill_2 FILLER_36_1078 ();
 sg13g2_fill_1 FILLER_36_1108 ();
 sg13g2_fill_2 FILLER_36_1117 ();
 sg13g2_fill_2 FILLER_36_1158 ();
 sg13g2_fill_1 FILLER_36_1226 ();
 sg13g2_fill_1 FILLER_36_1237 ();
 sg13g2_fill_2 FILLER_36_1264 ();
 sg13g2_fill_1 FILLER_36_1266 ();
 sg13g2_fill_1 FILLER_36_1294 ();
 sg13g2_fill_1 FILLER_36_1305 ();
 sg13g2_fill_1 FILLER_36_1375 ();
 sg13g2_fill_2 FILLER_36_1382 ();
 sg13g2_fill_2 FILLER_36_1394 ();
 sg13g2_fill_1 FILLER_36_1396 ();
 sg13g2_fill_1 FILLER_36_1445 ();
 sg13g2_fill_1 FILLER_36_1454 ();
 sg13g2_decap_4 FILLER_36_1585 ();
 sg13g2_fill_1 FILLER_36_1630 ();
 sg13g2_fill_1 FILLER_36_1650 ();
 sg13g2_fill_1 FILLER_36_1699 ();
 sg13g2_fill_1 FILLER_36_1747 ();
 sg13g2_decap_4 FILLER_36_1778 ();
 sg13g2_fill_2 FILLER_36_1812 ();
 sg13g2_fill_1 FILLER_36_1814 ();
 sg13g2_fill_1 FILLER_36_1847 ();
 sg13g2_fill_2 FILLER_36_1914 ();
 sg13g2_fill_1 FILLER_36_1916 ();
 sg13g2_fill_1 FILLER_36_1998 ();
 sg13g2_fill_2 FILLER_36_2013 ();
 sg13g2_fill_1 FILLER_36_2015 ();
 sg13g2_fill_1 FILLER_36_2051 ();
 sg13g2_fill_2 FILLER_36_2116 ();
 sg13g2_fill_1 FILLER_36_2118 ();
 sg13g2_fill_2 FILLER_36_2123 ();
 sg13g2_fill_2 FILLER_36_2149 ();
 sg13g2_fill_1 FILLER_36_2151 ();
 sg13g2_fill_1 FILLER_36_2175 ();
 sg13g2_fill_2 FILLER_36_2235 ();
 sg13g2_fill_1 FILLER_36_2237 ();
 sg13g2_fill_1 FILLER_36_2252 ();
 sg13g2_fill_2 FILLER_36_2275 ();
 sg13g2_fill_1 FILLER_36_2277 ();
 sg13g2_fill_1 FILLER_36_2411 ();
 sg13g2_fill_1 FILLER_36_2490 ();
 sg13g2_fill_2 FILLER_36_2565 ();
 sg13g2_decap_8 FILLER_36_2636 ();
 sg13g2_decap_8 FILLER_36_2643 ();
 sg13g2_decap_8 FILLER_36_2650 ();
 sg13g2_decap_8 FILLER_36_2657 ();
 sg13g2_decap_8 FILLER_36_2664 ();
 sg13g2_fill_2 FILLER_36_2671 ();
 sg13g2_fill_1 FILLER_36_2673 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_15 ();
 sg13g2_fill_2 FILLER_37_36 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_fill_1 FILLER_37_69 ();
 sg13g2_decap_4 FILLER_37_80 ();
 sg13g2_fill_2 FILLER_37_89 ();
 sg13g2_fill_1 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_97 ();
 sg13g2_fill_1 FILLER_37_107 ();
 sg13g2_fill_1 FILLER_37_113 ();
 sg13g2_fill_2 FILLER_37_133 ();
 sg13g2_fill_1 FILLER_37_135 ();
 sg13g2_fill_2 FILLER_37_155 ();
 sg13g2_fill_1 FILLER_37_157 ();
 sg13g2_fill_2 FILLER_37_170 ();
 sg13g2_fill_1 FILLER_37_172 ();
 sg13g2_fill_2 FILLER_37_203 ();
 sg13g2_fill_2 FILLER_37_250 ();
 sg13g2_fill_2 FILLER_37_270 ();
 sg13g2_fill_1 FILLER_37_272 ();
 sg13g2_fill_2 FILLER_37_281 ();
 sg13g2_fill_1 FILLER_37_283 ();
 sg13g2_fill_2 FILLER_37_294 ();
 sg13g2_fill_2 FILLER_37_303 ();
 sg13g2_fill_1 FILLER_37_314 ();
 sg13g2_fill_1 FILLER_37_328 ();
 sg13g2_fill_1 FILLER_37_391 ();
 sg13g2_fill_2 FILLER_37_452 ();
 sg13g2_fill_2 FILLER_37_463 ();
 sg13g2_fill_1 FILLER_37_570 ();
 sg13g2_fill_2 FILLER_37_706 ();
 sg13g2_fill_1 FILLER_37_708 ();
 sg13g2_fill_2 FILLER_37_760 ();
 sg13g2_fill_1 FILLER_37_762 ();
 sg13g2_fill_2 FILLER_37_785 ();
 sg13g2_fill_2 FILLER_37_806 ();
 sg13g2_fill_1 FILLER_37_808 ();
 sg13g2_fill_1 FILLER_37_892 ();
 sg13g2_fill_2 FILLER_37_908 ();
 sg13g2_fill_1 FILLER_37_910 ();
 sg13g2_fill_1 FILLER_37_927 ();
 sg13g2_fill_2 FILLER_37_931 ();
 sg13g2_fill_1 FILLER_37_942 ();
 sg13g2_fill_1 FILLER_37_974 ();
 sg13g2_fill_1 FILLER_37_989 ();
 sg13g2_fill_1 FILLER_37_1012 ();
 sg13g2_fill_2 FILLER_37_1023 ();
 sg13g2_fill_2 FILLER_37_1038 ();
 sg13g2_fill_1 FILLER_37_1040 ();
 sg13g2_fill_2 FILLER_37_1057 ();
 sg13g2_fill_1 FILLER_37_1059 ();
 sg13g2_fill_2 FILLER_37_1088 ();
 sg13g2_fill_1 FILLER_37_1090 ();
 sg13g2_fill_1 FILLER_37_1134 ();
 sg13g2_fill_1 FILLER_37_1139 ();
 sg13g2_fill_1 FILLER_37_1156 ();
 sg13g2_fill_2 FILLER_37_1188 ();
 sg13g2_fill_1 FILLER_37_1222 ();
 sg13g2_fill_1 FILLER_37_1246 ();
 sg13g2_fill_2 FILLER_37_1251 ();
 sg13g2_fill_1 FILLER_37_1253 ();
 sg13g2_decap_4 FILLER_37_1357 ();
 sg13g2_fill_2 FILLER_37_1408 ();
 sg13g2_fill_2 FILLER_37_1436 ();
 sg13g2_decap_8 FILLER_37_1448 ();
 sg13g2_decap_4 FILLER_37_1455 ();
 sg13g2_fill_2 FILLER_37_1459 ();
 sg13g2_fill_1 FILLER_37_1491 ();
 sg13g2_decap_4 FILLER_37_1505 ();
 sg13g2_decap_8 FILLER_37_1523 ();
 sg13g2_fill_2 FILLER_37_1530 ();
 sg13g2_fill_1 FILLER_37_1532 ();
 sg13g2_decap_4 FILLER_37_1537 ();
 sg13g2_fill_1 FILLER_37_1541 ();
 sg13g2_decap_8 FILLER_37_1590 ();
 sg13g2_fill_2 FILLER_37_1597 ();
 sg13g2_fill_2 FILLER_37_1623 ();
 sg13g2_fill_1 FILLER_37_1625 ();
 sg13g2_fill_2 FILLER_37_1636 ();
 sg13g2_fill_1 FILLER_37_1638 ();
 sg13g2_fill_2 FILLER_37_1816 ();
 sg13g2_fill_1 FILLER_37_1860 ();
 sg13g2_fill_2 FILLER_37_1887 ();
 sg13g2_fill_1 FILLER_37_1889 ();
 sg13g2_fill_2 FILLER_37_1921 ();
 sg13g2_fill_1 FILLER_37_1943 ();
 sg13g2_fill_1 FILLER_37_1958 ();
 sg13g2_fill_2 FILLER_37_2001 ();
 sg13g2_fill_2 FILLER_37_2058 ();
 sg13g2_fill_1 FILLER_37_2134 ();
 sg13g2_fill_2 FILLER_37_2161 ();
 sg13g2_fill_1 FILLER_37_2189 ();
 sg13g2_fill_1 FILLER_37_2205 ();
 sg13g2_fill_1 FILLER_37_2232 ();
 sg13g2_fill_2 FILLER_37_2338 ();
 sg13g2_fill_1 FILLER_37_2340 ();
 sg13g2_decap_8 FILLER_37_2419 ();
 sg13g2_fill_1 FILLER_37_2508 ();
 sg13g2_fill_1 FILLER_37_2525 ();
 sg13g2_fill_1 FILLER_37_2554 ();
 sg13g2_fill_2 FILLER_37_2612 ();
 sg13g2_fill_1 FILLER_37_2614 ();
 sg13g2_decap_8 FILLER_37_2641 ();
 sg13g2_decap_8 FILLER_37_2648 ();
 sg13g2_decap_8 FILLER_37_2655 ();
 sg13g2_decap_8 FILLER_37_2662 ();
 sg13g2_decap_4 FILLER_37_2669 ();
 sg13g2_fill_1 FILLER_37_2673 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_fill_1 FILLER_38_51 ();
 sg13g2_fill_2 FILLER_38_58 ();
 sg13g2_decap_8 FILLER_38_75 ();
 sg13g2_fill_1 FILLER_38_82 ();
 sg13g2_fill_2 FILLER_38_123 ();
 sg13g2_fill_1 FILLER_38_149 ();
 sg13g2_fill_1 FILLER_38_155 ();
 sg13g2_fill_2 FILLER_38_161 ();
 sg13g2_fill_1 FILLER_38_163 ();
 sg13g2_fill_2 FILLER_38_173 ();
 sg13g2_fill_2 FILLER_38_197 ();
 sg13g2_fill_2 FILLER_38_234 ();
 sg13g2_fill_2 FILLER_38_329 ();
 sg13g2_decap_4 FILLER_38_340 ();
 sg13g2_fill_1 FILLER_38_344 ();
 sg13g2_fill_2 FILLER_38_350 ();
 sg13g2_fill_1 FILLER_38_368 ();
 sg13g2_fill_2 FILLER_38_373 ();
 sg13g2_fill_1 FILLER_38_392 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_fill_2 FILLER_38_484 ();
 sg13g2_fill_1 FILLER_38_486 ();
 sg13g2_fill_1 FILLER_38_506 ();
 sg13g2_fill_2 FILLER_38_532 ();
 sg13g2_fill_2 FILLER_38_555 ();
 sg13g2_fill_1 FILLER_38_557 ();
 sg13g2_fill_1 FILLER_38_586 ();
 sg13g2_fill_2 FILLER_38_618 ();
 sg13g2_fill_1 FILLER_38_665 ();
 sg13g2_fill_2 FILLER_38_748 ();
 sg13g2_fill_1 FILLER_38_750 ();
 sg13g2_fill_1 FILLER_38_822 ();
 sg13g2_fill_2 FILLER_38_828 ();
 sg13g2_fill_1 FILLER_38_857 ();
 sg13g2_fill_1 FILLER_38_885 ();
 sg13g2_fill_1 FILLER_38_957 ();
 sg13g2_fill_2 FILLER_38_964 ();
 sg13g2_fill_2 FILLER_38_1068 ();
 sg13g2_fill_1 FILLER_38_1084 ();
 sg13g2_decap_4 FILLER_38_1105 ();
 sg13g2_fill_1 FILLER_38_1195 ();
 sg13g2_fill_1 FILLER_38_1220 ();
 sg13g2_fill_2 FILLER_38_1247 ();
 sg13g2_fill_1 FILLER_38_1288 ();
 sg13g2_fill_2 FILLER_38_1294 ();
 sg13g2_fill_1 FILLER_38_1344 ();
 sg13g2_fill_2 FILLER_38_1360 ();
 sg13g2_fill_1 FILLER_38_1362 ();
 sg13g2_fill_2 FILLER_38_1373 ();
 sg13g2_fill_1 FILLER_38_1375 ();
 sg13g2_fill_2 FILLER_38_1403 ();
 sg13g2_fill_2 FILLER_38_1432 ();
 sg13g2_fill_1 FILLER_38_1480 ();
 sg13g2_fill_2 FILLER_38_1512 ();
 sg13g2_fill_1 FILLER_38_1527 ();
 sg13g2_decap_4 FILLER_38_1545 ();
 sg13g2_fill_2 FILLER_38_1549 ();
 sg13g2_decap_8 FILLER_38_1563 ();
 sg13g2_decap_4 FILLER_38_1570 ();
 sg13g2_fill_1 FILLER_38_1656 ();
 sg13g2_fill_2 FILLER_38_1667 ();
 sg13g2_fill_1 FILLER_38_1669 ();
 sg13g2_fill_1 FILLER_38_1743 ();
 sg13g2_fill_2 FILLER_38_1763 ();
 sg13g2_fill_2 FILLER_38_1793 ();
 sg13g2_fill_1 FILLER_38_1814 ();
 sg13g2_fill_1 FILLER_38_1848 ();
 sg13g2_fill_2 FILLER_38_1960 ();
 sg13g2_fill_1 FILLER_38_1962 ();
 sg13g2_fill_2 FILLER_38_2008 ();
 sg13g2_fill_1 FILLER_38_2038 ();
 sg13g2_fill_2 FILLER_38_2090 ();
 sg13g2_fill_2 FILLER_38_2098 ();
 sg13g2_fill_2 FILLER_38_2132 ();
 sg13g2_fill_1 FILLER_38_2134 ();
 sg13g2_fill_2 FILLER_38_2144 ();
 sg13g2_fill_2 FILLER_38_2183 ();
 sg13g2_fill_1 FILLER_38_2185 ();
 sg13g2_fill_1 FILLER_38_2228 ();
 sg13g2_fill_2 FILLER_38_2261 ();
 sg13g2_fill_1 FILLER_38_2263 ();
 sg13g2_fill_1 FILLER_38_2319 ();
 sg13g2_fill_1 FILLER_38_2346 ();
 sg13g2_fill_2 FILLER_38_2357 ();
 sg13g2_fill_2 FILLER_38_2386 ();
 sg13g2_fill_1 FILLER_38_2448 ();
 sg13g2_fill_2 FILLER_38_2485 ();
 sg13g2_fill_2 FILLER_38_2500 ();
 sg13g2_fill_2 FILLER_38_2506 ();
 sg13g2_fill_1 FILLER_38_2565 ();
 sg13g2_fill_2 FILLER_38_2595 ();
 sg13g2_fill_1 FILLER_38_2597 ();
 sg13g2_fill_1 FILLER_38_2623 ();
 sg13g2_decap_8 FILLER_38_2650 ();
 sg13g2_decap_8 FILLER_38_2657 ();
 sg13g2_decap_8 FILLER_38_2664 ();
 sg13g2_fill_2 FILLER_38_2671 ();
 sg13g2_fill_1 FILLER_38_2673 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_4 ();
 sg13g2_fill_2 FILLER_39_19 ();
 sg13g2_fill_1 FILLER_39_29 ();
 sg13g2_fill_2 FILLER_39_35 ();
 sg13g2_fill_1 FILLER_39_37 ();
 sg13g2_fill_2 FILLER_39_59 ();
 sg13g2_fill_1 FILLER_39_66 ();
 sg13g2_decap_4 FILLER_39_90 ();
 sg13g2_fill_1 FILLER_39_94 ();
 sg13g2_fill_2 FILLER_39_105 ();
 sg13g2_fill_2 FILLER_39_131 ();
 sg13g2_fill_2 FILLER_39_164 ();
 sg13g2_fill_1 FILLER_39_204 ();
 sg13g2_fill_2 FILLER_39_218 ();
 sg13g2_fill_1 FILLER_39_220 ();
 sg13g2_fill_2 FILLER_39_259 ();
 sg13g2_fill_2 FILLER_39_302 ();
 sg13g2_fill_2 FILLER_39_404 ();
 sg13g2_fill_1 FILLER_39_406 ();
 sg13g2_fill_2 FILLER_39_433 ();
 sg13g2_fill_1 FILLER_39_449 ();
 sg13g2_fill_2 FILLER_39_498 ();
 sg13g2_fill_1 FILLER_39_500 ();
 sg13g2_fill_1 FILLER_39_515 ();
 sg13g2_fill_2 FILLER_39_525 ();
 sg13g2_fill_2 FILLER_39_541 ();
 sg13g2_fill_1 FILLER_39_569 ();
 sg13g2_fill_1 FILLER_39_611 ();
 sg13g2_fill_2 FILLER_39_628 ();
 sg13g2_fill_1 FILLER_39_630 ();
 sg13g2_fill_1 FILLER_39_754 ();
 sg13g2_fill_2 FILLER_39_769 ();
 sg13g2_fill_2 FILLER_39_925 ();
 sg13g2_fill_1 FILLER_39_927 ();
 sg13g2_fill_1 FILLER_39_953 ();
 sg13g2_fill_1 FILLER_39_997 ();
 sg13g2_decap_4 FILLER_39_1034 ();
 sg13g2_fill_2 FILLER_39_1046 ();
 sg13g2_fill_1 FILLER_39_1048 ();
 sg13g2_fill_2 FILLER_39_1093 ();
 sg13g2_fill_2 FILLER_39_1103 ();
 sg13g2_fill_1 FILLER_39_1105 ();
 sg13g2_fill_2 FILLER_39_1159 ();
 sg13g2_fill_1 FILLER_39_1161 ();
 sg13g2_fill_1 FILLER_39_1167 ();
 sg13g2_fill_1 FILLER_39_1226 ();
 sg13g2_fill_2 FILLER_39_1240 ();
 sg13g2_fill_2 FILLER_39_1320 ();
 sg13g2_fill_2 FILLER_39_1357 ();
 sg13g2_fill_2 FILLER_39_1368 ();
 sg13g2_fill_1 FILLER_39_1388 ();
 sg13g2_fill_2 FILLER_39_1441 ();
 sg13g2_fill_1 FILLER_39_1443 ();
 sg13g2_fill_2 FILLER_39_1470 ();
 sg13g2_fill_1 FILLER_39_1476 ();
 sg13g2_fill_1 FILLER_39_1531 ();
 sg13g2_fill_1 FILLER_39_1550 ();
 sg13g2_decap_4 FILLER_39_1559 ();
 sg13g2_fill_1 FILLER_39_1563 ();
 sg13g2_fill_2 FILLER_39_1625 ();
 sg13g2_fill_1 FILLER_39_1627 ();
 sg13g2_fill_2 FILLER_39_1658 ();
 sg13g2_fill_1 FILLER_39_1660 ();
 sg13g2_fill_2 FILLER_39_1696 ();
 sg13g2_fill_1 FILLER_39_1698 ();
 sg13g2_fill_2 FILLER_39_1738 ();
 sg13g2_fill_2 FILLER_39_1744 ();
 sg13g2_fill_1 FILLER_39_1746 ();
 sg13g2_fill_2 FILLER_39_1766 ();
 sg13g2_fill_2 FILLER_39_1794 ();
 sg13g2_fill_1 FILLER_39_1800 ();
 sg13g2_fill_1 FILLER_39_1846 ();
 sg13g2_fill_2 FILLER_39_1880 ();
 sg13g2_fill_1 FILLER_39_1882 ();
 sg13g2_fill_2 FILLER_39_1919 ();
 sg13g2_fill_1 FILLER_39_1926 ();
 sg13g2_fill_2 FILLER_39_1942 ();
 sg13g2_fill_2 FILLER_39_1960 ();
 sg13g2_fill_1 FILLER_39_1962 ();
 sg13g2_fill_2 FILLER_39_1987 ();
 sg13g2_fill_1 FILLER_39_1989 ();
 sg13g2_fill_2 FILLER_39_2084 ();
 sg13g2_fill_2 FILLER_39_2122 ();
 sg13g2_fill_1 FILLER_39_2124 ();
 sg13g2_fill_1 FILLER_39_2146 ();
 sg13g2_fill_2 FILLER_39_2182 ();
 sg13g2_fill_1 FILLER_39_2184 ();
 sg13g2_fill_2 FILLER_39_2194 ();
 sg13g2_fill_1 FILLER_39_2196 ();
 sg13g2_fill_2 FILLER_39_2227 ();
 sg13g2_fill_1 FILLER_39_2229 ();
 sg13g2_decap_8 FILLER_39_2238 ();
 sg13g2_fill_1 FILLER_39_2280 ();
 sg13g2_fill_1 FILLER_39_2330 ();
 sg13g2_fill_1 FILLER_39_2376 ();
 sg13g2_fill_2 FILLER_39_2412 ();
 sg13g2_fill_1 FILLER_39_2414 ();
 sg13g2_fill_2 FILLER_39_2424 ();
 sg13g2_fill_2 FILLER_39_2462 ();
 sg13g2_fill_1 FILLER_39_2464 ();
 sg13g2_fill_2 FILLER_39_2551 ();
 sg13g2_fill_2 FILLER_39_2612 ();
 sg13g2_fill_1 FILLER_39_2614 ();
 sg13g2_decap_8 FILLER_39_2641 ();
 sg13g2_decap_8 FILLER_39_2648 ();
 sg13g2_decap_8 FILLER_39_2655 ();
 sg13g2_decap_8 FILLER_39_2662 ();
 sg13g2_decap_4 FILLER_39_2669 ();
 sg13g2_fill_1 FILLER_39_2673 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_7 ();
 sg13g2_decap_4 FILLER_40_54 ();
 sg13g2_fill_1 FILLER_40_58 ();
 sg13g2_fill_2 FILLER_40_68 ();
 sg13g2_fill_1 FILLER_40_90 ();
 sg13g2_decap_8 FILLER_40_111 ();
 sg13g2_fill_2 FILLER_40_118 ();
 sg13g2_fill_1 FILLER_40_120 ();
 sg13g2_fill_2 FILLER_40_154 ();
 sg13g2_fill_1 FILLER_40_156 ();
 sg13g2_fill_2 FILLER_40_205 ();
 sg13g2_fill_2 FILLER_40_242 ();
 sg13g2_fill_1 FILLER_40_244 ();
 sg13g2_fill_1 FILLER_40_267 ();
 sg13g2_fill_1 FILLER_40_324 ();
 sg13g2_fill_1 FILLER_40_391 ();
 sg13g2_fill_1 FILLER_40_423 ();
 sg13g2_fill_1 FILLER_40_448 ();
 sg13g2_fill_1 FILLER_40_484 ();
 sg13g2_fill_2 FILLER_40_537 ();
 sg13g2_fill_1 FILLER_40_539 ();
 sg13g2_fill_1 FILLER_40_555 ();
 sg13g2_fill_1 FILLER_40_570 ();
 sg13g2_fill_2 FILLER_40_585 ();
 sg13g2_fill_1 FILLER_40_587 ();
 sg13g2_fill_1 FILLER_40_601 ();
 sg13g2_decap_4 FILLER_40_618 ();
 sg13g2_fill_2 FILLER_40_638 ();
 sg13g2_fill_1 FILLER_40_640 ();
 sg13g2_fill_2 FILLER_40_682 ();
 sg13g2_fill_1 FILLER_40_684 ();
 sg13g2_fill_1 FILLER_40_693 ();
 sg13g2_fill_1 FILLER_40_698 ();
 sg13g2_fill_2 FILLER_40_707 ();
 sg13g2_fill_2 FILLER_40_732 ();
 sg13g2_fill_1 FILLER_40_734 ();
 sg13g2_fill_2 FILLER_40_784 ();
 sg13g2_fill_1 FILLER_40_786 ();
 sg13g2_decap_4 FILLER_40_795 ();
 sg13g2_fill_2 FILLER_40_833 ();
 sg13g2_fill_2 FILLER_40_839 ();
 sg13g2_decap_8 FILLER_40_854 ();
 sg13g2_fill_2 FILLER_40_861 ();
 sg13g2_decap_4 FILLER_40_867 ();
 sg13g2_fill_2 FILLER_40_891 ();
 sg13g2_fill_1 FILLER_40_893 ();
 sg13g2_fill_2 FILLER_40_939 ();
 sg13g2_fill_1 FILLER_40_941 ();
 sg13g2_fill_1 FILLER_40_947 ();
 sg13g2_fill_1 FILLER_40_961 ();
 sg13g2_fill_1 FILLER_40_981 ();
 sg13g2_decap_4 FILLER_40_991 ();
 sg13g2_fill_1 FILLER_40_995 ();
 sg13g2_fill_2 FILLER_40_1104 ();
 sg13g2_fill_1 FILLER_40_1106 ();
 sg13g2_fill_2 FILLER_40_1117 ();
 sg13g2_fill_1 FILLER_40_1119 ();
 sg13g2_fill_2 FILLER_40_1156 ();
 sg13g2_fill_1 FILLER_40_1158 ();
 sg13g2_fill_2 FILLER_40_1252 ();
 sg13g2_fill_2 FILLER_40_1282 ();
 sg13g2_fill_1 FILLER_40_1289 ();
 sg13g2_fill_2 FILLER_40_1312 ();
 sg13g2_fill_2 FILLER_40_1328 ();
 sg13g2_fill_1 FILLER_40_1359 ();
 sg13g2_fill_2 FILLER_40_1370 ();
 sg13g2_fill_1 FILLER_40_1372 ();
 sg13g2_fill_1 FILLER_40_1397 ();
 sg13g2_fill_2 FILLER_40_1425 ();
 sg13g2_decap_4 FILLER_40_1437 ();
 sg13g2_decap_4 FILLER_40_1449 ();
 sg13g2_fill_2 FILLER_40_1488 ();
 sg13g2_fill_1 FILLER_40_1490 ();
 sg13g2_fill_2 FILLER_40_1510 ();
 sg13g2_fill_1 FILLER_40_1512 ();
 sg13g2_fill_1 FILLER_40_1519 ();
 sg13g2_decap_4 FILLER_40_1525 ();
 sg13g2_fill_2 FILLER_40_1529 ();
 sg13g2_fill_1 FILLER_40_1548 ();
 sg13g2_fill_1 FILLER_40_1554 ();
 sg13g2_decap_8 FILLER_40_1570 ();
 sg13g2_fill_1 FILLER_40_1604 ();
 sg13g2_decap_8 FILLER_40_1631 ();
 sg13g2_fill_1 FILLER_40_1668 ();
 sg13g2_fill_2 FILLER_40_1776 ();
 sg13g2_fill_1 FILLER_40_1778 ();
 sg13g2_fill_1 FILLER_40_1783 ();
 sg13g2_fill_2 FILLER_40_1835 ();
 sg13g2_fill_1 FILLER_40_1951 ();
 sg13g2_fill_2 FILLER_40_1978 ();
 sg13g2_fill_1 FILLER_40_1980 ();
 sg13g2_fill_1 FILLER_40_2033 ();
 sg13g2_decap_8 FILLER_40_2044 ();
 sg13g2_decap_8 FILLER_40_2051 ();
 sg13g2_decap_8 FILLER_40_2066 ();
 sg13g2_fill_2 FILLER_40_2073 ();
 sg13g2_fill_1 FILLER_40_2075 ();
 sg13g2_fill_1 FILLER_40_2093 ();
 sg13g2_fill_1 FILLER_40_2108 ();
 sg13g2_decap_8 FILLER_40_2213 ();
 sg13g2_fill_1 FILLER_40_2220 ();
 sg13g2_fill_2 FILLER_40_2247 ();
 sg13g2_fill_1 FILLER_40_2249 ();
 sg13g2_decap_4 FILLER_40_2255 ();
 sg13g2_fill_2 FILLER_40_2259 ();
 sg13g2_fill_1 FILLER_40_2304 ();
 sg13g2_fill_2 FILLER_40_2360 ();
 sg13g2_fill_2 FILLER_40_2371 ();
 sg13g2_fill_2 FILLER_40_2404 ();
 sg13g2_fill_1 FILLER_40_2406 ();
 sg13g2_fill_1 FILLER_40_2433 ();
 sg13g2_fill_2 FILLER_40_2443 ();
 sg13g2_fill_1 FILLER_40_2445 ();
 sg13g2_decap_4 FILLER_40_2463 ();
 sg13g2_decap_4 FILLER_40_2482 ();
 sg13g2_fill_2 FILLER_40_2490 ();
 sg13g2_fill_2 FILLER_40_2496 ();
 sg13g2_fill_1 FILLER_40_2510 ();
 sg13g2_fill_2 FILLER_40_2585 ();
 sg13g2_fill_1 FILLER_40_2587 ();
 sg13g2_decap_4 FILLER_40_2609 ();
 sg13g2_fill_1 FILLER_40_2613 ();
 sg13g2_decap_8 FILLER_40_2657 ();
 sg13g2_decap_8 FILLER_40_2664 ();
 sg13g2_fill_2 FILLER_40_2671 ();
 sg13g2_fill_1 FILLER_40_2673 ();
 sg13g2_decap_4 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_47 ();
 sg13g2_decap_8 FILLER_41_54 ();
 sg13g2_fill_2 FILLER_41_61 ();
 sg13g2_fill_1 FILLER_41_63 ();
 sg13g2_fill_2 FILLER_41_69 ();
 sg13g2_fill_1 FILLER_41_71 ();
 sg13g2_fill_1 FILLER_41_96 ();
 sg13g2_fill_2 FILLER_41_109 ();
 sg13g2_fill_1 FILLER_41_111 ();
 sg13g2_fill_2 FILLER_41_117 ();
 sg13g2_decap_8 FILLER_41_128 ();
 sg13g2_fill_2 FILLER_41_144 ();
 sg13g2_decap_4 FILLER_41_182 ();
 sg13g2_fill_2 FILLER_41_198 ();
 sg13g2_fill_1 FILLER_41_200 ();
 sg13g2_fill_2 FILLER_41_318 ();
 sg13g2_fill_2 FILLER_41_380 ();
 sg13g2_fill_2 FILLER_41_386 ();
 sg13g2_fill_1 FILLER_41_482 ();
 sg13g2_fill_2 FILLER_41_493 ();
 sg13g2_fill_2 FILLER_41_515 ();
 sg13g2_fill_1 FILLER_41_517 ();
 sg13g2_fill_2 FILLER_41_627 ();
 sg13g2_fill_1 FILLER_41_637 ();
 sg13g2_fill_2 FILLER_41_710 ();
 sg13g2_fill_1 FILLER_41_712 ();
 sg13g2_fill_1 FILLER_41_758 ();
 sg13g2_fill_2 FILLER_41_800 ();
 sg13g2_fill_2 FILLER_41_860 ();
 sg13g2_fill_1 FILLER_41_862 ();
 sg13g2_fill_2 FILLER_41_875 ();
 sg13g2_fill_1 FILLER_41_877 ();
 sg13g2_fill_1 FILLER_41_893 ();
 sg13g2_decap_4 FILLER_41_899 ();
 sg13g2_fill_2 FILLER_41_909 ();
 sg13g2_fill_1 FILLER_41_911 ();
 sg13g2_fill_2 FILLER_41_948 ();
 sg13g2_fill_2 FILLER_41_960 ();
 sg13g2_fill_1 FILLER_41_962 ();
 sg13g2_fill_1 FILLER_41_980 ();
 sg13g2_fill_1 FILLER_41_1015 ();
 sg13g2_fill_1 FILLER_41_1071 ();
 sg13g2_fill_2 FILLER_41_1108 ();
 sg13g2_fill_1 FILLER_41_1110 ();
 sg13g2_fill_1 FILLER_41_1141 ();
 sg13g2_decap_8 FILLER_41_1148 ();
 sg13g2_fill_2 FILLER_41_1155 ();
 sg13g2_fill_1 FILLER_41_1157 ();
 sg13g2_decap_8 FILLER_41_1175 ();
 sg13g2_fill_1 FILLER_41_1237 ();
 sg13g2_fill_2 FILLER_41_1313 ();
 sg13g2_fill_2 FILLER_41_1320 ();
 sg13g2_fill_2 FILLER_41_1336 ();
 sg13g2_fill_1 FILLER_41_1357 ();
 sg13g2_fill_1 FILLER_41_1379 ();
 sg13g2_decap_4 FILLER_41_1388 ();
 sg13g2_fill_2 FILLER_41_1392 ();
 sg13g2_fill_1 FILLER_41_1423 ();
 sg13g2_fill_2 FILLER_41_1447 ();
 sg13g2_fill_1 FILLER_41_1449 ();
 sg13g2_fill_2 FILLER_41_1460 ();
 sg13g2_fill_1 FILLER_41_1462 ();
 sg13g2_fill_1 FILLER_41_1495 ();
 sg13g2_fill_2 FILLER_41_1512 ();
 sg13g2_fill_1 FILLER_41_1524 ();
 sg13g2_decap_4 FILLER_41_1537 ();
 sg13g2_fill_1 FILLER_41_1554 ();
 sg13g2_fill_2 FILLER_41_1563 ();
 sg13g2_fill_1 FILLER_41_1565 ();
 sg13g2_fill_1 FILLER_41_1574 ();
 sg13g2_decap_8 FILLER_41_1592 ();
 sg13g2_decap_4 FILLER_41_1718 ();
 sg13g2_fill_1 FILLER_41_1722 ();
 sg13g2_fill_2 FILLER_41_1759 ();
 sg13g2_fill_1 FILLER_41_1761 ();
 sg13g2_fill_1 FILLER_41_1812 ();
 sg13g2_fill_1 FILLER_41_1840 ();
 sg13g2_fill_2 FILLER_41_1851 ();
 sg13g2_decap_4 FILLER_41_1904 ();
 sg13g2_fill_2 FILLER_41_1912 ();
 sg13g2_decap_4 FILLER_41_1918 ();
 sg13g2_fill_1 FILLER_41_1922 ();
 sg13g2_fill_1 FILLER_41_1934 ();
 sg13g2_fill_2 FILLER_41_1940 ();
 sg13g2_fill_2 FILLER_41_1953 ();
 sg13g2_fill_1 FILLER_41_1979 ();
 sg13g2_fill_2 FILLER_41_2019 ();
 sg13g2_fill_1 FILLER_41_2026 ();
 sg13g2_fill_1 FILLER_41_2067 ();
 sg13g2_fill_2 FILLER_41_2074 ();
 sg13g2_fill_1 FILLER_41_2076 ();
 sg13g2_fill_1 FILLER_41_2083 ();
 sg13g2_fill_1 FILLER_41_2093 ();
 sg13g2_fill_2 FILLER_41_2115 ();
 sg13g2_fill_1 FILLER_41_2117 ();
 sg13g2_fill_2 FILLER_41_2160 ();
 sg13g2_fill_1 FILLER_41_2188 ();
 sg13g2_decap_8 FILLER_41_2216 ();
 sg13g2_fill_1 FILLER_41_2223 ();
 sg13g2_fill_1 FILLER_41_2277 ();
 sg13g2_fill_2 FILLER_41_2290 ();
 sg13g2_fill_1 FILLER_41_2342 ();
 sg13g2_fill_2 FILLER_41_2357 ();
 sg13g2_fill_1 FILLER_41_2379 ();
 sg13g2_fill_2 FILLER_41_2421 ();
 sg13g2_fill_1 FILLER_41_2423 ();
 sg13g2_fill_1 FILLER_41_2450 ();
 sg13g2_decap_4 FILLER_41_2481 ();
 sg13g2_fill_1 FILLER_41_2485 ();
 sg13g2_fill_1 FILLER_41_2512 ();
 sg13g2_fill_2 FILLER_41_2545 ();
 sg13g2_fill_1 FILLER_41_2547 ();
 sg13g2_fill_1 FILLER_41_2558 ();
 sg13g2_fill_2 FILLER_41_2582 ();
 sg13g2_fill_1 FILLER_41_2584 ();
 sg13g2_decap_4 FILLER_41_2612 ();
 sg13g2_decap_8 FILLER_41_2642 ();
 sg13g2_decap_8 FILLER_41_2649 ();
 sg13g2_decap_8 FILLER_41_2656 ();
 sg13g2_decap_8 FILLER_41_2663 ();
 sg13g2_decap_4 FILLER_41_2670 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_16 ();
 sg13g2_fill_2 FILLER_42_27 ();
 sg13g2_fill_1 FILLER_42_29 ();
 sg13g2_decap_8 FILLER_42_62 ();
 sg13g2_fill_1 FILLER_42_69 ();
 sg13g2_fill_2 FILLER_42_80 ();
 sg13g2_fill_1 FILLER_42_93 ();
 sg13g2_decap_8 FILLER_42_108 ();
 sg13g2_fill_1 FILLER_42_115 ();
 sg13g2_decap_4 FILLER_42_130 ();
 sg13g2_fill_2 FILLER_42_162 ();
 sg13g2_fill_1 FILLER_42_164 ();
 sg13g2_decap_4 FILLER_42_193 ();
 sg13g2_fill_2 FILLER_42_257 ();
 sg13g2_fill_2 FILLER_42_298 ();
 sg13g2_fill_2 FILLER_42_385 ();
 sg13g2_fill_2 FILLER_42_391 ();
 sg13g2_fill_1 FILLER_42_393 ();
 sg13g2_fill_1 FILLER_42_419 ();
 sg13g2_fill_2 FILLER_42_450 ();
 sg13g2_fill_2 FILLER_42_519 ();
 sg13g2_fill_1 FILLER_42_521 ();
 sg13g2_fill_2 FILLER_42_527 ();
 sg13g2_fill_1 FILLER_42_538 ();
 sg13g2_fill_1 FILLER_42_550 ();
 sg13g2_fill_2 FILLER_42_556 ();
 sg13g2_fill_1 FILLER_42_558 ();
 sg13g2_fill_2 FILLER_42_580 ();
 sg13g2_decap_8 FILLER_42_598 ();
 sg13g2_fill_2 FILLER_42_605 ();
 sg13g2_decap_4 FILLER_42_617 ();
 sg13g2_fill_2 FILLER_42_621 ();
 sg13g2_fill_2 FILLER_42_641 ();
 sg13g2_fill_1 FILLER_42_643 ();
 sg13g2_fill_2 FILLER_42_679 ();
 sg13g2_fill_1 FILLER_42_681 ();
 sg13g2_fill_1 FILLER_42_729 ();
 sg13g2_fill_2 FILLER_42_750 ();
 sg13g2_fill_1 FILLER_42_752 ();
 sg13g2_fill_2 FILLER_42_758 ();
 sg13g2_decap_8 FILLER_42_790 ();
 sg13g2_fill_1 FILLER_42_815 ();
 sg13g2_fill_2 FILLER_42_843 ();
 sg13g2_fill_1 FILLER_42_845 ();
 sg13g2_fill_2 FILLER_42_860 ();
 sg13g2_decap_8 FILLER_42_888 ();
 sg13g2_fill_1 FILLER_42_908 ();
 sg13g2_fill_1 FILLER_42_949 ();
 sg13g2_fill_1 FILLER_42_1007 ();
 sg13g2_fill_1 FILLER_42_1014 ();
 sg13g2_fill_2 FILLER_42_1029 ();
 sg13g2_fill_1 FILLER_42_1031 ();
 sg13g2_fill_2 FILLER_42_1041 ();
 sg13g2_fill_1 FILLER_42_1043 ();
 sg13g2_fill_1 FILLER_42_1078 ();
 sg13g2_fill_2 FILLER_42_1089 ();
 sg13g2_fill_1 FILLER_42_1091 ();
 sg13g2_fill_1 FILLER_42_1101 ();
 sg13g2_fill_1 FILLER_42_1133 ();
 sg13g2_decap_4 FILLER_42_1178 ();
 sg13g2_fill_2 FILLER_42_1230 ();
 sg13g2_fill_1 FILLER_42_1253 ();
 sg13g2_fill_2 FILLER_42_1259 ();
 sg13g2_fill_2 FILLER_42_1272 ();
 sg13g2_fill_1 FILLER_42_1342 ();
 sg13g2_fill_2 FILLER_42_1352 ();
 sg13g2_fill_1 FILLER_42_1377 ();
 sg13g2_decap_4 FILLER_42_1448 ();
 sg13g2_fill_1 FILLER_42_1478 ();
 sg13g2_fill_1 FILLER_42_1496 ();
 sg13g2_fill_2 FILLER_42_1526 ();
 sg13g2_fill_1 FILLER_42_1528 ();
 sg13g2_fill_2 FILLER_42_1543 ();
 sg13g2_fill_1 FILLER_42_1549 ();
 sg13g2_decap_4 FILLER_42_1570 ();
 sg13g2_decap_4 FILLER_42_1588 ();
 sg13g2_fill_2 FILLER_42_1622 ();
 sg13g2_fill_2 FILLER_42_1664 ();
 sg13g2_fill_1 FILLER_42_1738 ();
 sg13g2_fill_1 FILLER_42_1884 ();
 sg13g2_fill_1 FILLER_42_1895 ();
 sg13g2_fill_1 FILLER_42_1938 ();
 sg13g2_fill_2 FILLER_42_1952 ();
 sg13g2_fill_1 FILLER_42_1954 ();
 sg13g2_fill_2 FILLER_42_1963 ();
 sg13g2_decap_8 FILLER_42_2009 ();
 sg13g2_fill_2 FILLER_42_2016 ();
 sg13g2_fill_1 FILLER_42_2018 ();
 sg13g2_fill_2 FILLER_42_2024 ();
 sg13g2_decap_4 FILLER_42_2043 ();
 sg13g2_fill_2 FILLER_42_2074 ();
 sg13g2_fill_2 FILLER_42_2112 ();
 sg13g2_fill_1 FILLER_42_2114 ();
 sg13g2_fill_2 FILLER_42_2120 ();
 sg13g2_fill_1 FILLER_42_2122 ();
 sg13g2_fill_1 FILLER_42_2143 ();
 sg13g2_fill_2 FILLER_42_2154 ();
 sg13g2_decap_4 FILLER_42_2175 ();
 sg13g2_fill_2 FILLER_42_2179 ();
 sg13g2_fill_2 FILLER_42_2231 ();
 sg13g2_fill_1 FILLER_42_2278 ();
 sg13g2_fill_1 FILLER_42_2287 ();
 sg13g2_fill_1 FILLER_42_2321 ();
 sg13g2_fill_1 FILLER_42_2331 ();
 sg13g2_fill_1 FILLER_42_2387 ();
 sg13g2_fill_1 FILLER_42_2400 ();
 sg13g2_fill_1 FILLER_42_2419 ();
 sg13g2_fill_2 FILLER_42_2436 ();
 sg13g2_decap_4 FILLER_42_2474 ();
 sg13g2_fill_2 FILLER_42_2478 ();
 sg13g2_fill_2 FILLER_42_2484 ();
 sg13g2_fill_2 FILLER_42_2500 ();
 sg13g2_fill_1 FILLER_42_2502 ();
 sg13g2_fill_1 FILLER_42_2602 ();
 sg13g2_fill_1 FILLER_42_2613 ();
 sg13g2_decap_8 FILLER_42_2640 ();
 sg13g2_decap_8 FILLER_42_2647 ();
 sg13g2_decap_8 FILLER_42_2654 ();
 sg13g2_decap_8 FILLER_42_2661 ();
 sg13g2_decap_4 FILLER_42_2668 ();
 sg13g2_fill_2 FILLER_42_2672 ();
 sg13g2_fill_2 FILLER_43_35 ();
 sg13g2_fill_1 FILLER_43_37 ();
 sg13g2_fill_1 FILLER_43_49 ();
 sg13g2_fill_2 FILLER_43_55 ();
 sg13g2_fill_2 FILLER_43_87 ();
 sg13g2_fill_1 FILLER_43_111 ();
 sg13g2_fill_1 FILLER_43_122 ();
 sg13g2_fill_1 FILLER_43_137 ();
 sg13g2_fill_2 FILLER_43_147 ();
 sg13g2_decap_4 FILLER_43_168 ();
 sg13g2_fill_2 FILLER_43_177 ();
 sg13g2_fill_1 FILLER_43_179 ();
 sg13g2_fill_1 FILLER_43_197 ();
 sg13g2_fill_2 FILLER_43_227 ();
 sg13g2_fill_2 FILLER_43_233 ();
 sg13g2_fill_1 FILLER_43_320 ();
 sg13g2_fill_1 FILLER_43_360 ();
 sg13g2_fill_2 FILLER_43_365 ();
 sg13g2_fill_1 FILLER_43_410 ();
 sg13g2_fill_2 FILLER_43_458 ();
 sg13g2_fill_2 FILLER_43_492 ();
 sg13g2_fill_1 FILLER_43_494 ();
 sg13g2_fill_2 FILLER_43_503 ();
 sg13g2_fill_1 FILLER_43_505 ();
 sg13g2_fill_1 FILLER_43_541 ();
 sg13g2_fill_2 FILLER_43_578 ();
 sg13g2_fill_1 FILLER_43_580 ();
 sg13g2_decap_4 FILLER_43_607 ();
 sg13g2_decap_8 FILLER_43_630 ();
 sg13g2_fill_2 FILLER_43_637 ();
 sg13g2_fill_2 FILLER_43_662 ();
 sg13g2_fill_1 FILLER_43_672 ();
 sg13g2_fill_1 FILLER_43_679 ();
 sg13g2_fill_1 FILLER_43_700 ();
 sg13g2_fill_1 FILLER_43_735 ();
 sg13g2_fill_2 FILLER_43_749 ();
 sg13g2_decap_4 FILLER_43_786 ();
 sg13g2_fill_1 FILLER_43_790 ();
 sg13g2_fill_1 FILLER_43_810 ();
 sg13g2_decap_4 FILLER_43_840 ();
 sg13g2_fill_1 FILLER_43_844 ();
 sg13g2_decap_4 FILLER_43_869 ();
 sg13g2_fill_2 FILLER_43_910 ();
 sg13g2_fill_1 FILLER_43_912 ();
 sg13g2_fill_2 FILLER_43_929 ();
 sg13g2_fill_1 FILLER_43_931 ();
 sg13g2_fill_2 FILLER_43_956 ();
 sg13g2_fill_1 FILLER_43_958 ();
 sg13g2_fill_1 FILLER_43_970 ();
 sg13g2_fill_1 FILLER_43_1041 ();
 sg13g2_fill_1 FILLER_43_1202 ();
 sg13g2_fill_2 FILLER_43_1255 ();
 sg13g2_fill_1 FILLER_43_1322 ();
 sg13g2_fill_1 FILLER_43_1331 ();
 sg13g2_fill_2 FILLER_43_1337 ();
 sg13g2_fill_1 FILLER_43_1370 ();
 sg13g2_fill_1 FILLER_43_1391 ();
 sg13g2_decap_8 FILLER_43_1401 ();
 sg13g2_decap_4 FILLER_43_1408 ();
 sg13g2_fill_2 FILLER_43_1412 ();
 sg13g2_fill_1 FILLER_43_1430 ();
 sg13g2_decap_8 FILLER_43_1435 ();
 sg13g2_fill_2 FILLER_43_1442 ();
 sg13g2_fill_1 FILLER_43_1444 ();
 sg13g2_fill_1 FILLER_43_1450 ();
 sg13g2_fill_1 FILLER_43_1477 ();
 sg13g2_decap_4 FILLER_43_1516 ();
 sg13g2_fill_1 FILLER_43_1520 ();
 sg13g2_fill_2 FILLER_43_1526 ();
 sg13g2_fill_2 FILLER_43_1533 ();
 sg13g2_decap_4 FILLER_43_1580 ();
 sg13g2_fill_1 FILLER_43_1592 ();
 sg13g2_fill_2 FILLER_43_1685 ();
 sg13g2_fill_1 FILLER_43_1687 ();
 sg13g2_fill_2 FILLER_43_1779 ();
 sg13g2_fill_2 FILLER_43_1799 ();
 sg13g2_fill_1 FILLER_43_1801 ();
 sg13g2_fill_1 FILLER_43_1859 ();
 sg13g2_fill_2 FILLER_43_1869 ();
 sg13g2_fill_1 FILLER_43_1871 ();
 sg13g2_fill_2 FILLER_43_1929 ();
 sg13g2_fill_1 FILLER_43_1931 ();
 sg13g2_fill_2 FILLER_43_1936 ();
 sg13g2_fill_2 FILLER_43_1985 ();
 sg13g2_decap_4 FILLER_43_2035 ();
 sg13g2_fill_1 FILLER_43_2039 ();
 sg13g2_fill_1 FILLER_43_2110 ();
 sg13g2_fill_1 FILLER_43_2285 ();
 sg13g2_fill_2 FILLER_43_2422 ();
 sg13g2_fill_1 FILLER_43_2424 ();
 sg13g2_fill_1 FILLER_43_2495 ();
 sg13g2_fill_1 FILLER_43_2510 ();
 sg13g2_fill_1 FILLER_43_2551 ();
 sg13g2_fill_2 FILLER_43_2564 ();
 sg13g2_fill_1 FILLER_43_2580 ();
 sg13g2_fill_1 FILLER_43_2585 ();
 sg13g2_fill_1 FILLER_43_2595 ();
 sg13g2_fill_2 FILLER_43_2612 ();
 sg13g2_fill_1 FILLER_43_2614 ();
 sg13g2_decap_8 FILLER_43_2641 ();
 sg13g2_decap_8 FILLER_43_2648 ();
 sg13g2_decap_8 FILLER_43_2655 ();
 sg13g2_decap_8 FILLER_43_2662 ();
 sg13g2_decap_4 FILLER_43_2669 ();
 sg13g2_fill_1 FILLER_43_2673 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_50 ();
 sg13g2_fill_2 FILLER_44_71 ();
 sg13g2_fill_1 FILLER_44_82 ();
 sg13g2_fill_2 FILLER_44_90 ();
 sg13g2_fill_1 FILLER_44_92 ();
 sg13g2_decap_8 FILLER_44_106 ();
 sg13g2_fill_1 FILLER_44_113 ();
 sg13g2_decap_4 FILLER_44_128 ();
 sg13g2_fill_1 FILLER_44_132 ();
 sg13g2_decap_4 FILLER_44_141 ();
 sg13g2_fill_2 FILLER_44_145 ();
 sg13g2_fill_1 FILLER_44_180 ();
 sg13g2_fill_1 FILLER_44_199 ();
 sg13g2_fill_2 FILLER_44_238 ();
 sg13g2_fill_2 FILLER_44_279 ();
 sg13g2_fill_1 FILLER_44_300 ();
 sg13g2_fill_1 FILLER_44_365 ();
 sg13g2_fill_1 FILLER_44_379 ();
 sg13g2_fill_2 FILLER_44_462 ();
 sg13g2_fill_1 FILLER_44_464 ();
 sg13g2_fill_2 FILLER_44_475 ();
 sg13g2_fill_1 FILLER_44_477 ();
 sg13g2_fill_2 FILLER_44_514 ();
 sg13g2_fill_1 FILLER_44_516 ();
 sg13g2_fill_1 FILLER_44_549 ();
 sg13g2_fill_2 FILLER_44_559 ();
 sg13g2_fill_1 FILLER_44_575 ();
 sg13g2_decap_4 FILLER_44_623 ();
 sg13g2_fill_2 FILLER_44_653 ();
 sg13g2_fill_1 FILLER_44_655 ();
 sg13g2_fill_1 FILLER_44_719 ();
 sg13g2_decap_4 FILLER_44_776 ();
 sg13g2_decap_4 FILLER_44_797 ();
 sg13g2_fill_1 FILLER_44_801 ();
 sg13g2_fill_2 FILLER_44_838 ();
 sg13g2_fill_2 FILLER_44_880 ();
 sg13g2_fill_2 FILLER_44_904 ();
 sg13g2_fill_1 FILLER_44_906 ();
 sg13g2_fill_1 FILLER_44_928 ();
 sg13g2_fill_2 FILLER_44_935 ();
 sg13g2_fill_1 FILLER_44_1008 ();
 sg13g2_fill_2 FILLER_44_1015 ();
 sg13g2_fill_1 FILLER_44_1022 ();
 sg13g2_fill_2 FILLER_44_1056 ();
 sg13g2_fill_2 FILLER_44_1072 ();
 sg13g2_fill_2 FILLER_44_1121 ();
 sg13g2_fill_1 FILLER_44_1123 ();
 sg13g2_fill_1 FILLER_44_1201 ();
 sg13g2_fill_1 FILLER_44_1211 ();
 sg13g2_fill_2 FILLER_44_1240 ();
 sg13g2_fill_2 FILLER_44_1255 ();
 sg13g2_fill_1 FILLER_44_1257 ();
 sg13g2_fill_1 FILLER_44_1267 ();
 sg13g2_fill_1 FILLER_44_1276 ();
 sg13g2_fill_2 FILLER_44_1311 ();
 sg13g2_fill_2 FILLER_44_1353 ();
 sg13g2_decap_8 FILLER_44_1359 ();
 sg13g2_fill_2 FILLER_44_1407 ();
 sg13g2_fill_1 FILLER_44_1409 ();
 sg13g2_decap_4 FILLER_44_1446 ();
 sg13g2_decap_8 FILLER_44_1455 ();
 sg13g2_fill_1 FILLER_44_1466 ();
 sg13g2_fill_2 FILLER_44_1471 ();
 sg13g2_fill_2 FILLER_44_1486 ();
 sg13g2_decap_8 FILLER_44_1496 ();
 sg13g2_decap_8 FILLER_44_1503 ();
 sg13g2_fill_2 FILLER_44_1510 ();
 sg13g2_fill_1 FILLER_44_1512 ();
 sg13g2_fill_1 FILLER_44_1529 ();
 sg13g2_fill_2 FILLER_44_1538 ();
 sg13g2_fill_1 FILLER_44_1540 ();
 sg13g2_fill_2 FILLER_44_1549 ();
 sg13g2_fill_1 FILLER_44_1551 ();
 sg13g2_fill_1 FILLER_44_1561 ();
 sg13g2_fill_1 FILLER_44_1598 ();
 sg13g2_fill_2 FILLER_44_1629 ();
 sg13g2_fill_1 FILLER_44_1656 ();
 sg13g2_fill_1 FILLER_44_1683 ();
 sg13g2_fill_2 FILLER_44_1688 ();
 sg13g2_fill_1 FILLER_44_1690 ();
 sg13g2_fill_1 FILLER_44_1736 ();
 sg13g2_fill_2 FILLER_44_1842 ();
 sg13g2_fill_2 FILLER_44_1855 ();
 sg13g2_fill_2 FILLER_44_1869 ();
 sg13g2_fill_2 FILLER_44_1890 ();
 sg13g2_fill_1 FILLER_44_1892 ();
 sg13g2_fill_2 FILLER_44_1919 ();
 sg13g2_fill_2 FILLER_44_1927 ();
 sg13g2_fill_1 FILLER_44_1929 ();
 sg13g2_fill_1 FILLER_44_1946 ();
 sg13g2_fill_2 FILLER_44_1952 ();
 sg13g2_fill_1 FILLER_44_1954 ();
 sg13g2_fill_2 FILLER_44_2054 ();
 sg13g2_fill_1 FILLER_44_2111 ();
 sg13g2_fill_2 FILLER_44_2134 ();
 sg13g2_fill_1 FILLER_44_2193 ();
 sg13g2_fill_2 FILLER_44_2215 ();
 sg13g2_fill_1 FILLER_44_2227 ();
 sg13g2_fill_1 FILLER_44_2258 ();
 sg13g2_fill_2 FILLER_44_2294 ();
 sg13g2_decap_4 FILLER_44_2300 ();
 sg13g2_fill_2 FILLER_44_2304 ();
 sg13g2_fill_2 FILLER_44_2316 ();
 sg13g2_fill_2 FILLER_44_2356 ();
 sg13g2_fill_1 FILLER_44_2358 ();
 sg13g2_fill_2 FILLER_44_2426 ();
 sg13g2_fill_1 FILLER_44_2458 ();
 sg13g2_fill_1 FILLER_44_2482 ();
 sg13g2_fill_2 FILLER_44_2553 ();
 sg13g2_fill_1 FILLER_44_2555 ();
 sg13g2_fill_2 FILLER_44_2571 ();
 sg13g2_fill_1 FILLER_44_2603 ();
 sg13g2_decap_8 FILLER_44_2640 ();
 sg13g2_decap_8 FILLER_44_2647 ();
 sg13g2_decap_8 FILLER_44_2654 ();
 sg13g2_decap_8 FILLER_44_2661 ();
 sg13g2_decap_4 FILLER_44_2668 ();
 sg13g2_fill_2 FILLER_44_2672 ();
 sg13g2_fill_1 FILLER_45_40 ();
 sg13g2_fill_2 FILLER_45_97 ();
 sg13g2_fill_2 FILLER_45_130 ();
 sg13g2_fill_1 FILLER_45_132 ();
 sg13g2_fill_2 FILLER_45_154 ();
 sg13g2_fill_2 FILLER_45_179 ();
 sg13g2_fill_2 FILLER_45_191 ();
 sg13g2_fill_1 FILLER_45_201 ();
 sg13g2_fill_2 FILLER_45_415 ();
 sg13g2_fill_2 FILLER_45_432 ();
 sg13g2_fill_1 FILLER_45_470 ();
 sg13g2_fill_1 FILLER_45_497 ();
 sg13g2_fill_2 FILLER_45_517 ();
 sg13g2_fill_1 FILLER_45_519 ();
 sg13g2_fill_2 FILLER_45_525 ();
 sg13g2_fill_1 FILLER_45_527 ();
 sg13g2_fill_1 FILLER_45_555 ();
 sg13g2_fill_2 FILLER_45_608 ();
 sg13g2_fill_1 FILLER_45_610 ();
 sg13g2_fill_2 FILLER_45_623 ();
 sg13g2_fill_2 FILLER_45_644 ();
 sg13g2_fill_1 FILLER_45_658 ();
 sg13g2_fill_1 FILLER_45_662 ();
 sg13g2_fill_1 FILLER_45_667 ();
 sg13g2_fill_2 FILLER_45_713 ();
 sg13g2_fill_2 FILLER_45_730 ();
 sg13g2_fill_2 FILLER_45_741 ();
 sg13g2_fill_2 FILLER_45_751 ();
 sg13g2_fill_1 FILLER_45_753 ();
 sg13g2_decap_4 FILLER_45_784 ();
 sg13g2_fill_2 FILLER_45_788 ();
 sg13g2_fill_1 FILLER_45_832 ();
 sg13g2_fill_2 FILLER_45_889 ();
 sg13g2_fill_1 FILLER_45_957 ();
 sg13g2_fill_2 FILLER_45_1014 ();
 sg13g2_fill_1 FILLER_45_1016 ();
 sg13g2_fill_2 FILLER_45_1043 ();
 sg13g2_fill_1 FILLER_45_1045 ();
 sg13g2_fill_2 FILLER_45_1076 ();
 sg13g2_fill_1 FILLER_45_1078 ();
 sg13g2_fill_2 FILLER_45_1105 ();
 sg13g2_fill_1 FILLER_45_1179 ();
 sg13g2_fill_2 FILLER_45_1284 ();
 sg13g2_fill_1 FILLER_45_1291 ();
 sg13g2_fill_1 FILLER_45_1302 ();
 sg13g2_fill_2 FILLER_45_1308 ();
 sg13g2_fill_1 FILLER_45_1320 ();
 sg13g2_decap_4 FILLER_45_1325 ();
 sg13g2_fill_2 FILLER_45_1329 ();
 sg13g2_fill_2 FILLER_45_1334 ();
 sg13g2_decap_4 FILLER_45_1340 ();
 sg13g2_fill_2 FILLER_45_1397 ();
 sg13g2_fill_1 FILLER_45_1399 ();
 sg13g2_fill_1 FILLER_45_1455 ();
 sg13g2_fill_2 FILLER_45_1494 ();
 sg13g2_fill_1 FILLER_45_1496 ();
 sg13g2_fill_2 FILLER_45_1521 ();
 sg13g2_decap_4 FILLER_45_1575 ();
 sg13g2_fill_2 FILLER_45_1579 ();
 sg13g2_fill_1 FILLER_45_1589 ();
 sg13g2_decap_4 FILLER_45_1598 ();
 sg13g2_fill_1 FILLER_45_1602 ();
 sg13g2_fill_2 FILLER_45_1757 ();
 sg13g2_fill_1 FILLER_45_1905 ();
 sg13g2_fill_2 FILLER_45_1993 ();
 sg13g2_fill_2 FILLER_45_2020 ();
 sg13g2_fill_2 FILLER_45_2109 ();
 sg13g2_fill_2 FILLER_45_2151 ();
 sg13g2_fill_1 FILLER_45_2153 ();
 sg13g2_fill_2 FILLER_45_2180 ();
 sg13g2_fill_1 FILLER_45_2226 ();
 sg13g2_fill_2 FILLER_45_2261 ();
 sg13g2_fill_2 FILLER_45_2272 ();
 sg13g2_fill_1 FILLER_45_2274 ();
 sg13g2_fill_2 FILLER_45_2311 ();
 sg13g2_fill_2 FILLER_45_2364 ();
 sg13g2_fill_1 FILLER_45_2366 ();
 sg13g2_fill_2 FILLER_45_2377 ();
 sg13g2_fill_1 FILLER_45_2393 ();
 sg13g2_fill_2 FILLER_45_2434 ();
 sg13g2_fill_1 FILLER_45_2436 ();
 sg13g2_fill_1 FILLER_45_2450 ();
 sg13g2_fill_2 FILLER_45_2523 ();
 sg13g2_fill_2 FILLER_45_2561 ();
 sg13g2_fill_2 FILLER_45_2577 ();
 sg13g2_fill_2 FILLER_45_2588 ();
 sg13g2_fill_2 FILLER_45_2621 ();
 sg13g2_fill_1 FILLER_45_2623 ();
 sg13g2_decap_8 FILLER_45_2641 ();
 sg13g2_decap_8 FILLER_45_2648 ();
 sg13g2_decap_8 FILLER_45_2655 ();
 sg13g2_decap_8 FILLER_45_2662 ();
 sg13g2_decap_4 FILLER_45_2669 ();
 sg13g2_fill_1 FILLER_45_2673 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_56 ();
 sg13g2_fill_1 FILLER_46_58 ();
 sg13g2_fill_2 FILLER_46_69 ();
 sg13g2_decap_4 FILLER_46_97 ();
 sg13g2_fill_2 FILLER_46_101 ();
 sg13g2_fill_2 FILLER_46_154 ();
 sg13g2_fill_1 FILLER_46_156 ();
 sg13g2_fill_1 FILLER_46_188 ();
 sg13g2_fill_2 FILLER_46_237 ();
 sg13g2_fill_2 FILLER_46_308 ();
 sg13g2_fill_2 FILLER_46_347 ();
 sg13g2_fill_1 FILLER_46_372 ();
 sg13g2_fill_2 FILLER_46_406 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_fill_2 FILLER_46_451 ();
 sg13g2_fill_1 FILLER_46_453 ();
 sg13g2_fill_2 FILLER_46_469 ();
 sg13g2_fill_2 FILLER_46_500 ();
 sg13g2_fill_1 FILLER_46_502 ();
 sg13g2_fill_2 FILLER_46_529 ();
 sg13g2_fill_1 FILLER_46_531 ();
 sg13g2_fill_2 FILLER_46_563 ();
 sg13g2_fill_2 FILLER_46_615 ();
 sg13g2_fill_1 FILLER_46_655 ();
 sg13g2_fill_1 FILLER_46_669 ();
 sg13g2_fill_1 FILLER_46_679 ();
 sg13g2_fill_1 FILLER_46_706 ();
 sg13g2_fill_2 FILLER_46_743 ();
 sg13g2_fill_1 FILLER_46_745 ();
 sg13g2_decap_4 FILLER_46_836 ();
 sg13g2_fill_2 FILLER_46_853 ();
 sg13g2_fill_2 FILLER_46_900 ();
 sg13g2_fill_1 FILLER_46_902 ();
 sg13g2_decap_4 FILLER_46_907 ();
 sg13g2_fill_1 FILLER_46_911 ();
 sg13g2_fill_1 FILLER_46_920 ();
 sg13g2_fill_1 FILLER_46_969 ();
 sg13g2_fill_2 FILLER_46_1015 ();
 sg13g2_fill_1 FILLER_46_1017 ();
 sg13g2_fill_2 FILLER_46_1048 ();
 sg13g2_fill_1 FILLER_46_1058 ();
 sg13g2_fill_2 FILLER_46_1099 ();
 sg13g2_fill_2 FILLER_46_1137 ();
 sg13g2_fill_1 FILLER_46_1139 ();
 sg13g2_fill_1 FILLER_46_1263 ();
 sg13g2_fill_2 FILLER_46_1277 ();
 sg13g2_fill_2 FILLER_46_1289 ();
 sg13g2_fill_1 FILLER_46_1291 ();
 sg13g2_fill_2 FILLER_46_1345 ();
 sg13g2_fill_1 FILLER_46_1347 ();
 sg13g2_decap_4 FILLER_46_1387 ();
 sg13g2_fill_2 FILLER_46_1398 ();
 sg13g2_fill_1 FILLER_46_1415 ();
 sg13g2_decap_4 FILLER_46_1468 ();
 sg13g2_fill_1 FILLER_46_1477 ();
 sg13g2_fill_1 FILLER_46_1556 ();
 sg13g2_fill_2 FILLER_46_1567 ();
 sg13g2_fill_1 FILLER_46_1574 ();
 sg13g2_fill_2 FILLER_46_1580 ();
 sg13g2_fill_1 FILLER_46_1603 ();
 sg13g2_fill_2 FILLER_46_1690 ();
 sg13g2_fill_1 FILLER_46_1692 ();
 sg13g2_fill_1 FILLER_46_1714 ();
 sg13g2_fill_1 FILLER_46_1750 ();
 sg13g2_fill_2 FILLER_46_1771 ();
 sg13g2_fill_1 FILLER_46_1773 ();
 sg13g2_fill_1 FILLER_46_1788 ();
 sg13g2_fill_2 FILLER_46_1794 ();
 sg13g2_fill_1 FILLER_46_1796 ();
 sg13g2_fill_1 FILLER_46_1842 ();
 sg13g2_fill_2 FILLER_46_1853 ();
 sg13g2_fill_1 FILLER_46_1855 ();
 sg13g2_fill_2 FILLER_46_1891 ();
 sg13g2_fill_1 FILLER_46_1893 ();
 sg13g2_decap_8 FILLER_46_1918 ();
 sg13g2_fill_1 FILLER_46_1930 ();
 sg13g2_fill_1 FILLER_46_1984 ();
 sg13g2_fill_1 FILLER_46_2011 ();
 sg13g2_fill_2 FILLER_46_2054 ();
 sg13g2_fill_2 FILLER_46_2077 ();
 sg13g2_fill_1 FILLER_46_2079 ();
 sg13g2_fill_1 FILLER_46_2094 ();
 sg13g2_fill_2 FILLER_46_2129 ();
 sg13g2_fill_1 FILLER_46_2148 ();
 sg13g2_fill_2 FILLER_46_2170 ();
 sg13g2_fill_1 FILLER_46_2172 ();
 sg13g2_fill_2 FILLER_46_2178 ();
 sg13g2_fill_1 FILLER_46_2180 ();
 sg13g2_fill_1 FILLER_46_2189 ();
 sg13g2_fill_2 FILLER_46_2237 ();
 sg13g2_fill_2 FILLER_46_2248 ();
 sg13g2_decap_4 FILLER_46_2304 ();
 sg13g2_fill_1 FILLER_46_2308 ();
 sg13g2_fill_1 FILLER_46_2319 ();
 sg13g2_fill_1 FILLER_46_2342 ();
 sg13g2_decap_4 FILLER_46_2379 ();
 sg13g2_decap_4 FILLER_46_2409 ();
 sg13g2_fill_1 FILLER_46_2413 ();
 sg13g2_decap_4 FILLER_46_2424 ();
 sg13g2_fill_2 FILLER_46_2454 ();
 sg13g2_fill_1 FILLER_46_2456 ();
 sg13g2_fill_2 FILLER_46_2522 ();
 sg13g2_fill_1 FILLER_46_2524 ();
 sg13g2_fill_2 FILLER_46_2565 ();
 sg13g2_fill_1 FILLER_46_2567 ();
 sg13g2_decap_8 FILLER_46_2648 ();
 sg13g2_decap_8 FILLER_46_2655 ();
 sg13g2_decap_8 FILLER_46_2662 ();
 sg13g2_decap_4 FILLER_46_2669 ();
 sg13g2_fill_1 FILLER_46_2673 ();
 sg13g2_decap_4 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_53 ();
 sg13g2_fill_2 FILLER_47_69 ();
 sg13g2_fill_1 FILLER_47_71 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_fill_1 FILLER_47_112 ();
 sg13g2_fill_1 FILLER_47_130 ();
 sg13g2_fill_2 FILLER_47_143 ();
 sg13g2_fill_1 FILLER_47_155 ();
 sg13g2_fill_2 FILLER_47_161 ();
 sg13g2_fill_2 FILLER_47_230 ();
 sg13g2_fill_2 FILLER_47_371 ();
 sg13g2_fill_1 FILLER_47_382 ();
 sg13g2_fill_1 FILLER_47_418 ();
 sg13g2_fill_1 FILLER_47_438 ();
 sg13g2_fill_2 FILLER_47_481 ();
 sg13g2_fill_2 FILLER_47_509 ();
 sg13g2_fill_2 FILLER_47_530 ();
 sg13g2_fill_1 FILLER_47_532 ();
 sg13g2_fill_2 FILLER_47_542 ();
 sg13g2_fill_1 FILLER_47_597 ();
 sg13g2_fill_2 FILLER_47_623 ();
 sg13g2_fill_2 FILLER_47_680 ();
 sg13g2_fill_1 FILLER_47_682 ();
 sg13g2_fill_1 FILLER_47_693 ();
 sg13g2_decap_8 FILLER_47_780 ();
 sg13g2_fill_2 FILLER_47_797 ();
 sg13g2_fill_1 FILLER_47_799 ();
 sg13g2_fill_1 FILLER_47_871 ();
 sg13g2_fill_1 FILLER_47_914 ();
 sg13g2_fill_2 FILLER_47_920 ();
 sg13g2_fill_1 FILLER_47_922 ();
 sg13g2_fill_2 FILLER_47_942 ();
 sg13g2_fill_1 FILLER_47_944 ();
 sg13g2_fill_2 FILLER_47_1043 ();
 sg13g2_fill_1 FILLER_47_1045 ();
 sg13g2_fill_1 FILLER_47_1072 ();
 sg13g2_fill_2 FILLER_47_1113 ();
 sg13g2_fill_1 FILLER_47_1115 ();
 sg13g2_fill_2 FILLER_47_1152 ();
 sg13g2_fill_1 FILLER_47_1239 ();
 sg13g2_fill_2 FILLER_47_1244 ();
 sg13g2_fill_1 FILLER_47_1268 ();
 sg13g2_decap_4 FILLER_47_1304 ();
 sg13g2_fill_1 FILLER_47_1308 ();
 sg13g2_fill_2 FILLER_47_1318 ();
 sg13g2_fill_1 FILLER_47_1320 ();
 sg13g2_decap_4 FILLER_47_1347 ();
 sg13g2_fill_2 FILLER_47_1397 ();
 sg13g2_fill_2 FILLER_47_1447 ();
 sg13g2_fill_2 FILLER_47_1491 ();
 sg13g2_fill_2 FILLER_47_1525 ();
 sg13g2_fill_1 FILLER_47_1527 ();
 sg13g2_fill_2 FILLER_47_1550 ();
 sg13g2_fill_1 FILLER_47_1552 ();
 sg13g2_fill_2 FILLER_47_1565 ();
 sg13g2_fill_1 FILLER_47_1567 ();
 sg13g2_fill_1 FILLER_47_1573 ();
 sg13g2_fill_1 FILLER_47_1592 ();
 sg13g2_fill_2 FILLER_47_1598 ();
 sg13g2_fill_1 FILLER_47_1654 ();
 sg13g2_fill_2 FILLER_47_1669 ();
 sg13g2_fill_2 FILLER_47_1734 ();
 sg13g2_fill_1 FILLER_47_1736 ();
 sg13g2_fill_2 FILLER_47_1745 ();
 sg13g2_fill_2 FILLER_47_1751 ();
 sg13g2_fill_1 FILLER_47_1753 ();
 sg13g2_fill_2 FILLER_47_1775 ();
 sg13g2_fill_1 FILLER_47_1777 ();
 sg13g2_fill_1 FILLER_47_1789 ();
 sg13g2_decap_8 FILLER_47_1798 ();
 sg13g2_decap_8 FILLER_47_1805 ();
 sg13g2_decap_4 FILLER_47_1812 ();
 sg13g2_fill_2 FILLER_47_1876 ();
 sg13g2_fill_1 FILLER_47_1878 ();
 sg13g2_fill_2 FILLER_47_1958 ();
 sg13g2_fill_2 FILLER_47_2005 ();
 sg13g2_fill_1 FILLER_47_2007 ();
 sg13g2_fill_2 FILLER_47_2064 ();
 sg13g2_fill_1 FILLER_47_2066 ();
 sg13g2_fill_2 FILLER_47_2110 ();
 sg13g2_fill_2 FILLER_47_2148 ();
 sg13g2_fill_2 FILLER_47_2155 ();
 sg13g2_fill_1 FILLER_47_2157 ();
 sg13g2_fill_2 FILLER_47_2176 ();
 sg13g2_fill_1 FILLER_47_2178 ();
 sg13g2_fill_2 FILLER_47_2205 ();
 sg13g2_fill_2 FILLER_47_2256 ();
 sg13g2_fill_1 FILLER_47_2276 ();
 sg13g2_fill_2 FILLER_47_2333 ();
 sg13g2_decap_4 FILLER_47_2363 ();
 sg13g2_fill_1 FILLER_47_2376 ();
 sg13g2_fill_2 FILLER_47_2390 ();
 sg13g2_fill_1 FILLER_47_2463 ();
 sg13g2_fill_1 FILLER_47_2490 ();
 sg13g2_decap_4 FILLER_47_2563 ();
 sg13g2_fill_1 FILLER_47_2601 ();
 sg13g2_fill_1 FILLER_47_2612 ();
 sg13g2_decap_8 FILLER_47_2639 ();
 sg13g2_decap_8 FILLER_47_2646 ();
 sg13g2_decap_8 FILLER_47_2653 ();
 sg13g2_decap_8 FILLER_47_2660 ();
 sg13g2_decap_8 FILLER_47_2667 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_61 ();
 sg13g2_fill_1 FILLER_48_63 ();
 sg13g2_fill_2 FILLER_48_147 ();
 sg13g2_fill_1 FILLER_48_217 ();
 sg13g2_fill_1 FILLER_48_240 ();
 sg13g2_fill_2 FILLER_48_267 ();
 sg13g2_fill_1 FILLER_48_284 ();
 sg13g2_fill_2 FILLER_48_295 ();
 sg13g2_fill_2 FILLER_48_302 ();
 sg13g2_fill_2 FILLER_48_334 ();
 sg13g2_fill_1 FILLER_48_394 ();
 sg13g2_fill_2 FILLER_48_437 ();
 sg13g2_fill_1 FILLER_48_453 ();
 sg13g2_fill_2 FILLER_48_492 ();
 sg13g2_fill_2 FILLER_48_554 ();
 sg13g2_fill_1 FILLER_48_565 ();
 sg13g2_fill_2 FILLER_48_570 ();
 sg13g2_fill_1 FILLER_48_572 ();
 sg13g2_fill_2 FILLER_48_619 ();
 sg13g2_fill_1 FILLER_48_621 ();
 sg13g2_fill_1 FILLER_48_649 ();
 sg13g2_fill_2 FILLER_48_673 ();
 sg13g2_fill_2 FILLER_48_746 ();
 sg13g2_fill_1 FILLER_48_765 ();
 sg13g2_decap_4 FILLER_48_833 ();
 sg13g2_fill_2 FILLER_48_837 ();
 sg13g2_fill_1 FILLER_48_852 ();
 sg13g2_fill_1 FILLER_48_904 ();
 sg13g2_fill_2 FILLER_48_946 ();
 sg13g2_fill_2 FILLER_48_970 ();
 sg13g2_fill_1 FILLER_48_972 ();
 sg13g2_fill_2 FILLER_48_1008 ();
 sg13g2_fill_2 FILLER_48_1061 ();
 sg13g2_fill_1 FILLER_48_1094 ();
 sg13g2_fill_2 FILLER_48_1108 ();
 sg13g2_fill_1 FILLER_48_1110 ();
 sg13g2_fill_1 FILLER_48_1149 ();
 sg13g2_fill_2 FILLER_48_1298 ();
 sg13g2_fill_2 FILLER_48_1335 ();
 sg13g2_fill_1 FILLER_48_1346 ();
 sg13g2_fill_2 FILLER_48_1382 ();
 sg13g2_fill_1 FILLER_48_1384 ();
 sg13g2_fill_1 FILLER_48_1468 ();
 sg13g2_fill_1 FILLER_48_1492 ();
 sg13g2_fill_2 FILLER_48_1512 ();
 sg13g2_fill_1 FILLER_48_1518 ();
 sg13g2_fill_2 FILLER_48_1527 ();
 sg13g2_fill_2 FILLER_48_1533 ();
 sg13g2_fill_1 FILLER_48_1535 ();
 sg13g2_fill_2 FILLER_48_1542 ();
 sg13g2_fill_2 FILLER_48_1550 ();
 sg13g2_fill_1 FILLER_48_1552 ();
 sg13g2_fill_1 FILLER_48_1576 ();
 sg13g2_fill_1 FILLER_48_1590 ();
 sg13g2_fill_2 FILLER_48_1645 ();
 sg13g2_fill_2 FILLER_48_1766 ();
 sg13g2_fill_1 FILLER_48_1768 ();
 sg13g2_fill_1 FILLER_48_1775 ();
 sg13g2_fill_1 FILLER_48_1786 ();
 sg13g2_fill_1 FILLER_48_1836 ();
 sg13g2_fill_2 FILLER_48_1851 ();
 sg13g2_fill_2 FILLER_48_1885 ();
 sg13g2_fill_1 FILLER_48_1933 ();
 sg13g2_fill_2 FILLER_48_1939 ();
 sg13g2_fill_1 FILLER_48_1946 ();
 sg13g2_fill_2 FILLER_48_1974 ();
 sg13g2_fill_1 FILLER_48_1976 ();
 sg13g2_fill_2 FILLER_48_2013 ();
 sg13g2_fill_2 FILLER_48_2030 ();
 sg13g2_fill_1 FILLER_48_2032 ();
 sg13g2_fill_2 FILLER_48_2090 ();
 sg13g2_fill_1 FILLER_48_2114 ();
 sg13g2_fill_2 FILLER_48_2220 ();
 sg13g2_fill_1 FILLER_48_2244 ();
 sg13g2_fill_1 FILLER_48_2322 ();
 sg13g2_fill_2 FILLER_48_2354 ();
 sg13g2_fill_1 FILLER_48_2356 ();
 sg13g2_decap_8 FILLER_48_2393 ();
 sg13g2_fill_1 FILLER_48_2400 ();
 sg13g2_decap_8 FILLER_48_2409 ();
 sg13g2_fill_2 FILLER_48_2430 ();
 sg13g2_fill_1 FILLER_48_2432 ();
 sg13g2_fill_1 FILLER_48_2469 ();
 sg13g2_fill_2 FILLER_48_2531 ();
 sg13g2_fill_1 FILLER_48_2560 ();
 sg13g2_fill_2 FILLER_48_2589 ();
 sg13g2_fill_1 FILLER_48_2621 ();
 sg13g2_decap_8 FILLER_48_2635 ();
 sg13g2_decap_8 FILLER_48_2642 ();
 sg13g2_decap_8 FILLER_48_2649 ();
 sg13g2_decap_8 FILLER_48_2656 ();
 sg13g2_decap_8 FILLER_48_2663 ();
 sg13g2_decap_4 FILLER_48_2670 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_4 FILLER_49_21 ();
 sg13g2_fill_2 FILLER_49_29 ();
 sg13g2_fill_2 FILLER_49_75 ();
 sg13g2_fill_1 FILLER_49_77 ();
 sg13g2_fill_2 FILLER_49_193 ();
 sg13g2_fill_1 FILLER_49_215 ();
 sg13g2_fill_1 FILLER_49_384 ();
 sg13g2_fill_2 FILLER_49_411 ();
 sg13g2_fill_2 FILLER_49_462 ();
 sg13g2_fill_2 FILLER_49_586 ();
 sg13g2_fill_1 FILLER_49_588 ();
 sg13g2_fill_1 FILLER_49_658 ();
 sg13g2_fill_1 FILLER_49_663 ();
 sg13g2_fill_2 FILLER_49_672 ();
 sg13g2_fill_2 FILLER_49_694 ();
 sg13g2_fill_1 FILLER_49_776 ();
 sg13g2_fill_2 FILLER_49_800 ();
 sg13g2_fill_1 FILLER_49_802 ();
 sg13g2_fill_1 FILLER_49_825 ();
 sg13g2_decap_4 FILLER_49_852 ();
 sg13g2_fill_2 FILLER_49_903 ();
 sg13g2_fill_1 FILLER_49_934 ();
 sg13g2_fill_2 FILLER_49_944 ();
 sg13g2_fill_1 FILLER_49_946 ();
 sg13g2_fill_2 FILLER_49_1027 ();
 sg13g2_fill_1 FILLER_49_1029 ();
 sg13g2_fill_1 FILLER_49_1035 ();
 sg13g2_fill_1 FILLER_49_1096 ();
 sg13g2_fill_1 FILLER_49_1143 ();
 sg13g2_fill_1 FILLER_49_1201 ();
 sg13g2_fill_1 FILLER_49_1233 ();
 sg13g2_fill_1 FILLER_49_1243 ();
 sg13g2_fill_1 FILLER_49_1290 ();
 sg13g2_fill_1 FILLER_49_1518 ();
 sg13g2_fill_1 FILLER_49_1534 ();
 sg13g2_fill_1 FILLER_49_1540 ();
 sg13g2_fill_2 FILLER_49_1555 ();
 sg13g2_fill_1 FILLER_49_1557 ();
 sg13g2_fill_2 FILLER_49_1564 ();
 sg13g2_fill_2 FILLER_49_1584 ();
 sg13g2_fill_2 FILLER_49_1624 ();
 sg13g2_fill_1 FILLER_49_1626 ();
 sg13g2_fill_2 FILLER_49_1656 ();
 sg13g2_fill_1 FILLER_49_1658 ();
 sg13g2_fill_2 FILLER_49_1669 ();
 sg13g2_fill_1 FILLER_49_1671 ();
 sg13g2_fill_1 FILLER_49_1681 ();
 sg13g2_fill_1 FILLER_49_1738 ();
 sg13g2_fill_1 FILLER_49_1753 ();
 sg13g2_fill_1 FILLER_49_1809 ();
 sg13g2_fill_2 FILLER_49_1824 ();
 sg13g2_fill_1 FILLER_49_1826 ();
 sg13g2_fill_2 FILLER_49_1908 ();
 sg13g2_fill_1 FILLER_49_1924 ();
 sg13g2_fill_1 FILLER_49_1950 ();
 sg13g2_fill_2 FILLER_49_2053 ();
 sg13g2_fill_2 FILLER_49_2098 ();
 sg13g2_fill_1 FILLER_49_2112 ();
 sg13g2_fill_2 FILLER_49_2139 ();
 sg13g2_fill_2 FILLER_49_2169 ();
 sg13g2_fill_1 FILLER_49_2171 ();
 sg13g2_fill_1 FILLER_49_2200 ();
 sg13g2_fill_2 FILLER_49_2228 ();
 sg13g2_fill_2 FILLER_49_2251 ();
 sg13g2_fill_2 FILLER_49_2306 ();
 sg13g2_fill_1 FILLER_49_2308 ();
 sg13g2_fill_2 FILLER_49_2330 ();
 sg13g2_fill_1 FILLER_49_2380 ();
 sg13g2_fill_2 FILLER_49_2472 ();
 sg13g2_fill_1 FILLER_49_2474 ();
 sg13g2_fill_1 FILLER_49_2508 ();
 sg13g2_fill_2 FILLER_49_2519 ();
 sg13g2_fill_1 FILLER_49_2521 ();
 sg13g2_decap_8 FILLER_49_2640 ();
 sg13g2_decap_8 FILLER_49_2647 ();
 sg13g2_decap_8 FILLER_49_2654 ();
 sg13g2_decap_8 FILLER_49_2661 ();
 sg13g2_decap_4 FILLER_49_2668 ();
 sg13g2_fill_2 FILLER_49_2672 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_fill_2 FILLER_50_42 ();
 sg13g2_fill_1 FILLER_50_44 ();
 sg13g2_fill_2 FILLER_50_156 ();
 sg13g2_fill_2 FILLER_50_178 ();
 sg13g2_fill_2 FILLER_50_206 ();
 sg13g2_fill_1 FILLER_50_328 ();
 sg13g2_fill_2 FILLER_50_338 ();
 sg13g2_fill_2 FILLER_50_373 ();
 sg13g2_fill_1 FILLER_50_379 ();
 sg13g2_fill_2 FILLER_50_406 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_fill_2 FILLER_50_505 ();
 sg13g2_fill_1 FILLER_50_507 ();
 sg13g2_fill_2 FILLER_50_548 ();
 sg13g2_fill_1 FILLER_50_550 ();
 sg13g2_fill_1 FILLER_50_578 ();
 sg13g2_fill_2 FILLER_50_600 ();
 sg13g2_fill_1 FILLER_50_602 ();
 sg13g2_fill_2 FILLER_50_651 ();
 sg13g2_fill_1 FILLER_50_653 ();
 sg13g2_fill_2 FILLER_50_722 ();
 sg13g2_fill_1 FILLER_50_724 ();
 sg13g2_fill_2 FILLER_50_756 ();
 sg13g2_fill_1 FILLER_50_758 ();
 sg13g2_fill_2 FILLER_50_915 ();
 sg13g2_fill_1 FILLER_50_960 ();
 sg13g2_fill_2 FILLER_50_967 ();
 sg13g2_fill_2 FILLER_50_993 ();
 sg13g2_fill_1 FILLER_50_995 ();
 sg13g2_fill_2 FILLER_50_1005 ();
 sg13g2_fill_1 FILLER_50_1007 ();
 sg13g2_fill_1 FILLER_50_1122 ();
 sg13g2_fill_2 FILLER_50_1161 ();
 sg13g2_fill_1 FILLER_50_1163 ();
 sg13g2_fill_1 FILLER_50_1208 ();
 sg13g2_fill_1 FILLER_50_1219 ();
 sg13g2_fill_2 FILLER_50_1225 ();
 sg13g2_fill_1 FILLER_50_1271 ();
 sg13g2_fill_2 FILLER_50_1322 ();
 sg13g2_fill_1 FILLER_50_1324 ();
 sg13g2_fill_2 FILLER_50_1348 ();
 sg13g2_fill_2 FILLER_50_1390 ();
 sg13g2_fill_2 FILLER_50_1405 ();
 sg13g2_fill_1 FILLER_50_1527 ();
 sg13g2_fill_1 FILLER_50_1536 ();
 sg13g2_fill_1 FILLER_50_1548 ();
 sg13g2_fill_1 FILLER_50_1559 ();
 sg13g2_decap_4 FILLER_50_1589 ();
 sg13g2_fill_2 FILLER_50_1603 ();
 sg13g2_fill_1 FILLER_50_1605 ();
 sg13g2_fill_2 FILLER_50_1702 ();
 sg13g2_fill_1 FILLER_50_1704 ();
 sg13g2_fill_2 FILLER_50_1726 ();
 sg13g2_fill_1 FILLER_50_1728 ();
 sg13g2_decap_4 FILLER_50_1733 ();
 sg13g2_fill_1 FILLER_50_1737 ();
 sg13g2_fill_2 FILLER_50_1773 ();
 sg13g2_fill_2 FILLER_50_1779 ();
 sg13g2_fill_1 FILLER_50_1781 ();
 sg13g2_fill_2 FILLER_50_1820 ();
 sg13g2_fill_1 FILLER_50_1822 ();
 sg13g2_decap_4 FILLER_50_1831 ();
 sg13g2_fill_2 FILLER_50_1840 ();
 sg13g2_fill_2 FILLER_50_1881 ();
 sg13g2_fill_1 FILLER_50_1893 ();
 sg13g2_fill_2 FILLER_50_1937 ();
 sg13g2_decap_4 FILLER_50_1961 ();
 sg13g2_fill_2 FILLER_50_1975 ();
 sg13g2_fill_2 FILLER_50_1991 ();
 sg13g2_fill_2 FILLER_50_2042 ();
 sg13g2_fill_2 FILLER_50_2081 ();
 sg13g2_fill_1 FILLER_50_2083 ();
 sg13g2_fill_1 FILLER_50_2094 ();
 sg13g2_fill_1 FILLER_50_2128 ();
 sg13g2_fill_1 FILLER_50_2162 ();
 sg13g2_fill_1 FILLER_50_2272 ();
 sg13g2_fill_2 FILLER_50_2286 ();
 sg13g2_fill_2 FILLER_50_2314 ();
 sg13g2_fill_2 FILLER_50_2342 ();
 sg13g2_fill_1 FILLER_50_2344 ();
 sg13g2_fill_1 FILLER_50_2410 ();
 sg13g2_fill_2 FILLER_50_2431 ();
 sg13g2_fill_1 FILLER_50_2433 ();
 sg13g2_fill_1 FILLER_50_2481 ();
 sg13g2_fill_2 FILLER_50_2512 ();
 sg13g2_fill_2 FILLER_50_2616 ();
 sg13g2_fill_1 FILLER_50_2618 ();
 sg13g2_decap_8 FILLER_50_2632 ();
 sg13g2_decap_8 FILLER_50_2639 ();
 sg13g2_decap_8 FILLER_50_2646 ();
 sg13g2_decap_8 FILLER_50_2653 ();
 sg13g2_decap_8 FILLER_50_2660 ();
 sg13g2_decap_8 FILLER_50_2667 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_4 FILLER_51_63 ();
 sg13g2_fill_2 FILLER_51_118 ();
 sg13g2_fill_2 FILLER_51_139 ();
 sg13g2_fill_2 FILLER_51_187 ();
 sg13g2_fill_1 FILLER_51_223 ();
 sg13g2_fill_1 FILLER_51_287 ();
 sg13g2_fill_1 FILLER_51_383 ();
 sg13g2_fill_2 FILLER_51_433 ();
 sg13g2_fill_1 FILLER_51_463 ();
 sg13g2_fill_2 FILLER_51_519 ();
 sg13g2_fill_1 FILLER_51_521 ();
 sg13g2_fill_1 FILLER_51_552 ();
 sg13g2_fill_1 FILLER_51_591 ();
 sg13g2_fill_1 FILLER_51_601 ();
 sg13g2_fill_1 FILLER_51_636 ();
 sg13g2_fill_2 FILLER_51_643 ();
 sg13g2_fill_1 FILLER_51_651 ();
 sg13g2_fill_2 FILLER_51_729 ();
 sg13g2_fill_1 FILLER_51_740 ();
 sg13g2_fill_1 FILLER_51_779 ();
 sg13g2_fill_1 FILLER_51_822 ();
 sg13g2_fill_1 FILLER_51_921 ();
 sg13g2_fill_2 FILLER_51_931 ();
 sg13g2_fill_1 FILLER_51_933 ();
 sg13g2_fill_1 FILLER_51_948 ();
 sg13g2_fill_1 FILLER_51_974 ();
 sg13g2_decap_4 FILLER_51_1022 ();
 sg13g2_fill_2 FILLER_51_1055 ();
 sg13g2_fill_2 FILLER_51_1071 ();
 sg13g2_fill_2 FILLER_51_1089 ();
 sg13g2_fill_1 FILLER_51_1091 ();
 sg13g2_fill_1 FILLER_51_1178 ();
 sg13g2_fill_2 FILLER_51_1193 ();
 sg13g2_fill_1 FILLER_51_1218 ();
 sg13g2_fill_1 FILLER_51_1264 ();
 sg13g2_decap_8 FILLER_51_1276 ();
 sg13g2_fill_1 FILLER_51_1287 ();
 sg13g2_fill_1 FILLER_51_1293 ();
 sg13g2_decap_8 FILLER_51_1303 ();
 sg13g2_fill_1 FILLER_51_1310 ();
 sg13g2_fill_2 FILLER_51_1337 ();
 sg13g2_fill_1 FILLER_51_1339 ();
 sg13g2_fill_1 FILLER_51_1435 ();
 sg13g2_fill_1 FILLER_51_1451 ();
 sg13g2_fill_1 FILLER_51_1456 ();
 sg13g2_fill_2 FILLER_51_1506 ();
 sg13g2_fill_1 FILLER_51_1508 ();
 sg13g2_decap_4 FILLER_51_1523 ();
 sg13g2_fill_2 FILLER_51_1553 ();
 sg13g2_fill_1 FILLER_51_1565 ();
 sg13g2_fill_1 FILLER_51_1585 ();
 sg13g2_decap_8 FILLER_51_1594 ();
 sg13g2_decap_4 FILLER_51_1601 ();
 sg13g2_decap_4 FILLER_51_1608 ();
 sg13g2_fill_1 FILLER_51_1612 ();
 sg13g2_fill_1 FILLER_51_1621 ();
 sg13g2_fill_1 FILLER_51_1650 ();
 sg13g2_fill_2 FILLER_51_1670 ();
 sg13g2_fill_1 FILLER_51_1672 ();
 sg13g2_decap_4 FILLER_51_1713 ();
 sg13g2_fill_1 FILLER_51_1717 ();
 sg13g2_fill_2 FILLER_51_1754 ();
 sg13g2_fill_1 FILLER_51_1756 ();
 sg13g2_fill_2 FILLER_51_1835 ();
 sg13g2_fill_1 FILLER_51_1837 ();
 sg13g2_fill_1 FILLER_51_1869 ();
 sg13g2_decap_8 FILLER_51_1914 ();
 sg13g2_fill_1 FILLER_51_1921 ();
 sg13g2_fill_2 FILLER_51_1948 ();
 sg13g2_fill_1 FILLER_51_1950 ();
 sg13g2_fill_2 FILLER_51_1981 ();
 sg13g2_fill_1 FILLER_51_1983 ();
 sg13g2_fill_2 FILLER_51_2014 ();
 sg13g2_fill_2 FILLER_51_2047 ();
 sg13g2_fill_1 FILLER_51_2049 ();
 sg13g2_fill_2 FILLER_51_2142 ();
 sg13g2_fill_1 FILLER_51_2144 ();
 sg13g2_fill_2 FILLER_51_2171 ();
 sg13g2_fill_2 FILLER_51_2196 ();
 sg13g2_fill_2 FILLER_51_2234 ();
 sg13g2_fill_1 FILLER_51_2302 ();
 sg13g2_fill_2 FILLER_51_2312 ();
 sg13g2_fill_1 FILLER_51_2314 ();
 sg13g2_fill_2 FILLER_51_2334 ();
 sg13g2_fill_2 FILLER_51_2447 ();
 sg13g2_fill_1 FILLER_51_2468 ();
 sg13g2_fill_2 FILLER_51_2573 ();
 sg13g2_decap_8 FILLER_51_2627 ();
 sg13g2_decap_8 FILLER_51_2634 ();
 sg13g2_decap_8 FILLER_51_2641 ();
 sg13g2_decap_8 FILLER_51_2648 ();
 sg13g2_decap_8 FILLER_51_2655 ();
 sg13g2_decap_8 FILLER_51_2662 ();
 sg13g2_decap_4 FILLER_51_2669 ();
 sg13g2_fill_1 FILLER_51_2673 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_4 FILLER_52_56 ();
 sg13g2_fill_2 FILLER_52_64 ();
 sg13g2_fill_1 FILLER_52_66 ();
 sg13g2_fill_1 FILLER_52_127 ();
 sg13g2_fill_1 FILLER_52_147 ();
 sg13g2_fill_1 FILLER_52_169 ();
 sg13g2_fill_2 FILLER_52_183 ();
 sg13g2_fill_1 FILLER_52_193 ();
 sg13g2_fill_1 FILLER_52_252 ();
 sg13g2_fill_1 FILLER_52_346 ();
 sg13g2_fill_2 FILLER_52_383 ();
 sg13g2_fill_2 FILLER_52_412 ();
 sg13g2_fill_1 FILLER_52_424 ();
 sg13g2_fill_2 FILLER_52_547 ();
 sg13g2_fill_1 FILLER_52_549 ();
 sg13g2_fill_1 FILLER_52_556 ();
 sg13g2_fill_2 FILLER_52_566 ();
 sg13g2_fill_2 FILLER_52_594 ();
 sg13g2_fill_2 FILLER_52_631 ();
 sg13g2_fill_1 FILLER_52_633 ();
 sg13g2_fill_2 FILLER_52_662 ();
 sg13g2_fill_2 FILLER_52_709 ();
 sg13g2_fill_2 FILLER_52_746 ();
 sg13g2_fill_2 FILLER_52_788 ();
 sg13g2_fill_1 FILLER_52_790 ();
 sg13g2_fill_2 FILLER_52_829 ();
 sg13g2_fill_1 FILLER_52_831 ();
 sg13g2_fill_2 FILLER_52_845 ();
 sg13g2_fill_2 FILLER_52_853 ();
 sg13g2_fill_1 FILLER_52_855 ();
 sg13g2_fill_2 FILLER_52_894 ();
 sg13g2_fill_1 FILLER_52_896 ();
 sg13g2_fill_1 FILLER_52_927 ();
 sg13g2_fill_2 FILLER_52_936 ();
 sg13g2_fill_1 FILLER_52_947 ();
 sg13g2_fill_1 FILLER_52_952 ();
 sg13g2_fill_1 FILLER_52_970 ();
 sg13g2_fill_2 FILLER_52_981 ();
 sg13g2_fill_2 FILLER_52_1060 ();
 sg13g2_fill_2 FILLER_52_1105 ();
 sg13g2_fill_1 FILLER_52_1107 ();
 sg13g2_fill_2 FILLER_52_1144 ();
 sg13g2_fill_2 FILLER_52_1172 ();
 sg13g2_fill_2 FILLER_52_1205 ();
 sg13g2_fill_2 FILLER_52_1219 ();
 sg13g2_fill_1 FILLER_52_1253 ();
 sg13g2_fill_2 FILLER_52_1305 ();
 sg13g2_fill_1 FILLER_52_1376 ();
 sg13g2_fill_1 FILLER_52_1402 ();
 sg13g2_fill_2 FILLER_52_1449 ();
 sg13g2_fill_2 FILLER_52_1459 ();
 sg13g2_fill_1 FILLER_52_1461 ();
 sg13g2_decap_4 FILLER_52_1528 ();
 sg13g2_fill_2 FILLER_52_1532 ();
 sg13g2_fill_2 FILLER_52_1546 ();
 sg13g2_fill_2 FILLER_52_1565 ();
 sg13g2_fill_1 FILLER_52_1580 ();
 sg13g2_fill_1 FILLER_52_1593 ();
 sg13g2_decap_8 FILLER_52_1606 ();
 sg13g2_fill_1 FILLER_52_1613 ();
 sg13g2_fill_2 FILLER_52_1641 ();
 sg13g2_fill_1 FILLER_52_1643 ();
 sg13g2_fill_2 FILLER_52_1679 ();
 sg13g2_fill_1 FILLER_52_1681 ();
 sg13g2_decap_4 FILLER_52_1713 ();
 sg13g2_fill_1 FILLER_52_1808 ();
 sg13g2_fill_2 FILLER_52_1843 ();
 sg13g2_fill_1 FILLER_52_1850 ();
 sg13g2_fill_2 FILLER_52_1883 ();
 sg13g2_fill_2 FILLER_52_1953 ();
 sg13g2_fill_2 FILLER_52_2013 ();
 sg13g2_fill_1 FILLER_52_2015 ();
 sg13g2_fill_2 FILLER_52_2041 ();
 sg13g2_fill_2 FILLER_52_2056 ();
 sg13g2_fill_2 FILLER_52_2068 ();
 sg13g2_fill_1 FILLER_52_2070 ();
 sg13g2_fill_1 FILLER_52_2107 ();
 sg13g2_fill_1 FILLER_52_2138 ();
 sg13g2_fill_1 FILLER_52_2173 ();
 sg13g2_fill_1 FILLER_52_2198 ();
 sg13g2_fill_1 FILLER_52_2240 ();
 sg13g2_fill_2 FILLER_52_2321 ();
 sg13g2_fill_2 FILLER_52_2358 ();
 sg13g2_fill_1 FILLER_52_2360 ();
 sg13g2_fill_2 FILLER_52_2376 ();
 sg13g2_fill_1 FILLER_52_2378 ();
 sg13g2_fill_2 FILLER_52_2419 ();
 sg13g2_fill_1 FILLER_52_2421 ();
 sg13g2_fill_1 FILLER_52_2483 ();
 sg13g2_fill_1 FILLER_52_2527 ();
 sg13g2_fill_2 FILLER_52_2568 ();
 sg13g2_fill_1 FILLER_52_2570 ();
 sg13g2_fill_1 FILLER_52_2611 ();
 sg13g2_decap_8 FILLER_52_2625 ();
 sg13g2_decap_8 FILLER_52_2632 ();
 sg13g2_decap_8 FILLER_52_2639 ();
 sg13g2_decap_8 FILLER_52_2646 ();
 sg13g2_decap_8 FILLER_52_2653 ();
 sg13g2_decap_8 FILLER_52_2660 ();
 sg13g2_decap_8 FILLER_52_2667 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_fill_1 FILLER_53_49 ();
 sg13g2_fill_2 FILLER_53_85 ();
 sg13g2_fill_1 FILLER_53_111 ();
 sg13g2_fill_1 FILLER_53_282 ();
 sg13g2_fill_1 FILLER_53_300 ();
 sg13g2_fill_2 FILLER_53_444 ();
 sg13g2_fill_2 FILLER_53_452 ();
 sg13g2_fill_1 FILLER_53_505 ();
 sg13g2_fill_1 FILLER_53_518 ();
 sg13g2_fill_1 FILLER_53_664 ();
 sg13g2_fill_2 FILLER_53_757 ();
 sg13g2_fill_2 FILLER_53_858 ();
 sg13g2_fill_1 FILLER_53_892 ();
 sg13g2_fill_1 FILLER_53_919 ();
 sg13g2_fill_2 FILLER_53_1023 ();
 sg13g2_fill_1 FILLER_53_1025 ();
 sg13g2_fill_1 FILLER_53_1059 ();
 sg13g2_fill_2 FILLER_53_1090 ();
 sg13g2_fill_1 FILLER_53_1092 ();
 sg13g2_fill_2 FILLER_53_1137 ();
 sg13g2_fill_1 FILLER_53_1139 ();
 sg13g2_fill_2 FILLER_53_1146 ();
 sg13g2_fill_1 FILLER_53_1169 ();
 sg13g2_fill_1 FILLER_53_1192 ();
 sg13g2_fill_2 FILLER_53_1218 ();
 sg13g2_fill_1 FILLER_53_1249 ();
 sg13g2_fill_1 FILLER_53_1258 ();
 sg13g2_fill_1 FILLER_53_1276 ();
 sg13g2_fill_2 FILLER_53_1281 ();
 sg13g2_fill_1 FILLER_53_1283 ();
 sg13g2_fill_2 FILLER_53_1293 ();
 sg13g2_fill_1 FILLER_53_1352 ();
 sg13g2_fill_2 FILLER_53_1374 ();
 sg13g2_fill_2 FILLER_53_1382 ();
 sg13g2_fill_1 FILLER_53_1384 ();
 sg13g2_fill_2 FILLER_53_1478 ();
 sg13g2_fill_1 FILLER_53_1510 ();
 sg13g2_fill_2 FILLER_53_1518 ();
 sg13g2_decap_8 FILLER_53_1532 ();
 sg13g2_fill_2 FILLER_53_1551 ();
 sg13g2_decap_8 FILLER_53_1561 ();
 sg13g2_fill_2 FILLER_53_1568 ();
 sg13g2_decap_4 FILLER_53_1583 ();
 sg13g2_fill_1 FILLER_53_1630 ();
 sg13g2_fill_2 FILLER_53_1657 ();
 sg13g2_fill_1 FILLER_53_1659 ();
 sg13g2_fill_1 FILLER_53_1686 ();
 sg13g2_fill_2 FILLER_53_1717 ();
 sg13g2_fill_1 FILLER_53_1719 ();
 sg13g2_fill_1 FILLER_53_1772 ();
 sg13g2_fill_2 FILLER_53_1777 ();
 sg13g2_fill_2 FILLER_53_1847 ();
 sg13g2_fill_1 FILLER_53_1849 ();
 sg13g2_fill_2 FILLER_53_1912 ();
 sg13g2_fill_1 FILLER_53_1914 ();
 sg13g2_fill_2 FILLER_53_1929 ();
 sg13g2_fill_1 FILLER_53_1931 ();
 sg13g2_fill_2 FILLER_53_1966 ();
 sg13g2_fill_1 FILLER_53_1968 ();
 sg13g2_fill_1 FILLER_53_2045 ();
 sg13g2_fill_1 FILLER_53_2081 ();
 sg13g2_fill_1 FILLER_53_2133 ();
 sg13g2_fill_2 FILLER_53_2143 ();
 sg13g2_fill_1 FILLER_53_2257 ();
 sg13g2_fill_2 FILLER_53_2385 ();
 sg13g2_fill_1 FILLER_53_2427 ();
 sg13g2_fill_1 FILLER_53_2454 ();
 sg13g2_decap_8 FILLER_53_2636 ();
 sg13g2_decap_8 FILLER_53_2643 ();
 sg13g2_decap_8 FILLER_53_2650 ();
 sg13g2_decap_8 FILLER_53_2657 ();
 sg13g2_decap_8 FILLER_53_2664 ();
 sg13g2_fill_2 FILLER_53_2671 ();
 sg13g2_fill_1 FILLER_53_2673 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_fill_2 FILLER_54_42 ();
 sg13g2_fill_1 FILLER_54_44 ();
 sg13g2_fill_1 FILLER_54_145 ();
 sg13g2_fill_1 FILLER_54_183 ();
 sg13g2_fill_2 FILLER_54_197 ();
 sg13g2_fill_1 FILLER_54_204 ();
 sg13g2_fill_1 FILLER_54_215 ();
 sg13g2_fill_2 FILLER_54_247 ();
 sg13g2_fill_2 FILLER_54_428 ();
 sg13g2_fill_2 FILLER_54_445 ();
 sg13g2_fill_1 FILLER_54_447 ();
 sg13g2_fill_2 FILLER_54_458 ();
 sg13g2_fill_1 FILLER_54_460 ();
 sg13g2_fill_2 FILLER_54_480 ();
 sg13g2_fill_1 FILLER_54_694 ();
 sg13g2_fill_1 FILLER_54_710 ();
 sg13g2_fill_1 FILLER_54_730 ();
 sg13g2_fill_1 FILLER_54_793 ();
 sg13g2_fill_1 FILLER_54_803 ();
 sg13g2_fill_2 FILLER_54_863 ();
 sg13g2_fill_1 FILLER_54_865 ();
 sg13g2_fill_1 FILLER_54_891 ();
 sg13g2_fill_1 FILLER_54_972 ();
 sg13g2_fill_2 FILLER_54_978 ();
 sg13g2_fill_2 FILLER_54_1045 ();
 sg13g2_fill_2 FILLER_54_1094 ();
 sg13g2_fill_1 FILLER_54_1096 ();
 sg13g2_fill_2 FILLER_54_1254 ();
 sg13g2_fill_1 FILLER_54_1256 ();
 sg13g2_fill_1 FILLER_54_1270 ();
 sg13g2_fill_1 FILLER_54_1284 ();
 sg13g2_fill_1 FILLER_54_1330 ();
 sg13g2_fill_1 FILLER_54_1429 ();
 sg13g2_fill_1 FILLER_54_1439 ();
 sg13g2_fill_2 FILLER_54_1449 ();
 sg13g2_fill_1 FILLER_54_1451 ();
 sg13g2_fill_1 FILLER_54_1493 ();
 sg13g2_fill_1 FILLER_54_1516 ();
 sg13g2_decap_4 FILLER_54_1541 ();
 sg13g2_fill_2 FILLER_54_1554 ();
 sg13g2_decap_4 FILLER_54_1581 ();
 sg13g2_fill_1 FILLER_54_1585 ();
 sg13g2_fill_1 FILLER_54_1615 ();
 sg13g2_fill_1 FILLER_54_1624 ();
 sg13g2_fill_2 FILLER_54_1644 ();
 sg13g2_fill_1 FILLER_54_1734 ();
 sg13g2_fill_1 FILLER_54_1763 ();
 sg13g2_fill_2 FILLER_54_1874 ();
 sg13g2_fill_2 FILLER_54_1931 ();
 sg13g2_fill_1 FILLER_54_1933 ();
 sg13g2_fill_2 FILLER_54_1942 ();
 sg13g2_fill_1 FILLER_54_1944 ();
 sg13g2_fill_1 FILLER_54_1989 ();
 sg13g2_fill_1 FILLER_54_2052 ();
 sg13g2_fill_2 FILLER_54_2093 ();
 sg13g2_fill_1 FILLER_54_2184 ();
 sg13g2_fill_2 FILLER_54_2194 ();
 sg13g2_fill_2 FILLER_54_2202 ();
 sg13g2_fill_1 FILLER_54_2242 ();
 sg13g2_fill_1 FILLER_54_2276 ();
 sg13g2_fill_1 FILLER_54_2287 ();
 sg13g2_fill_1 FILLER_54_2298 ();
 sg13g2_fill_1 FILLER_54_2313 ();
 sg13g2_fill_2 FILLER_54_2364 ();
 sg13g2_fill_2 FILLER_54_2445 ();
 sg13g2_fill_2 FILLER_54_2491 ();
 sg13g2_fill_1 FILLER_54_2575 ();
 sg13g2_fill_2 FILLER_54_2594 ();
 sg13g2_fill_1 FILLER_54_2596 ();
 sg13g2_decap_8 FILLER_54_2635 ();
 sg13g2_decap_8 FILLER_54_2642 ();
 sg13g2_decap_8 FILLER_54_2649 ();
 sg13g2_decap_8 FILLER_54_2656 ();
 sg13g2_decap_8 FILLER_54_2663 ();
 sg13g2_decap_4 FILLER_54_2670 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_4 FILLER_55_28 ();
 sg13g2_fill_2 FILLER_55_32 ();
 sg13g2_fill_1 FILLER_55_86 ();
 sg13g2_fill_1 FILLER_55_112 ();
 sg13g2_fill_2 FILLER_55_122 ();
 sg13g2_fill_2 FILLER_55_129 ();
 sg13g2_fill_1 FILLER_55_139 ();
 sg13g2_fill_2 FILLER_55_292 ();
 sg13g2_fill_2 FILLER_55_308 ();
 sg13g2_fill_1 FILLER_55_324 ();
 sg13g2_fill_1 FILLER_55_346 ();
 sg13g2_fill_2 FILLER_55_445 ();
 sg13g2_fill_1 FILLER_55_447 ();
 sg13g2_fill_2 FILLER_55_483 ();
 sg13g2_fill_2 FILLER_55_514 ();
 sg13g2_fill_1 FILLER_55_516 ();
 sg13g2_fill_2 FILLER_55_522 ();
 sg13g2_fill_2 FILLER_55_529 ();
 sg13g2_fill_2 FILLER_55_555 ();
 sg13g2_fill_2 FILLER_55_566 ();
 sg13g2_fill_1 FILLER_55_624 ();
 sg13g2_fill_1 FILLER_55_640 ();
 sg13g2_fill_2 FILLER_55_677 ();
 sg13g2_fill_2 FILLER_55_742 ();
 sg13g2_fill_1 FILLER_55_744 ();
 sg13g2_fill_2 FILLER_55_750 ();
 sg13g2_fill_1 FILLER_55_760 ();
 sg13g2_fill_2 FILLER_55_782 ();
 sg13g2_fill_2 FILLER_55_829 ();
 sg13g2_fill_1 FILLER_55_831 ();
 sg13g2_fill_1 FILLER_55_882 ();
 sg13g2_fill_2 FILLER_55_909 ();
 sg13g2_fill_1 FILLER_55_911 ();
 sg13g2_fill_2 FILLER_55_921 ();
 sg13g2_fill_2 FILLER_55_955 ();
 sg13g2_fill_1 FILLER_55_957 ();
 sg13g2_fill_2 FILLER_55_1059 ();
 sg13g2_fill_1 FILLER_55_1061 ();
 sg13g2_fill_2 FILLER_55_1144 ();
 sg13g2_fill_2 FILLER_55_1158 ();
 sg13g2_fill_1 FILLER_55_1250 ();
 sg13g2_decap_4 FILLER_55_1293 ();
 sg13g2_fill_1 FILLER_55_1300 ();
 sg13g2_fill_1 FILLER_55_1378 ();
 sg13g2_fill_2 FILLER_55_1393 ();
 sg13g2_fill_2 FILLER_55_1459 ();
 sg13g2_fill_1 FILLER_55_1474 ();
 sg13g2_fill_2 FILLER_55_1503 ();
 sg13g2_fill_2 FILLER_55_1518 ();
 sg13g2_fill_1 FILLER_55_1520 ();
 sg13g2_fill_2 FILLER_55_1556 ();
 sg13g2_decap_4 FILLER_55_1566 ();
 sg13g2_fill_2 FILLER_55_1586 ();
 sg13g2_decap_4 FILLER_55_1593 ();
 sg13g2_fill_2 FILLER_55_1662 ();
 sg13g2_fill_2 FILLER_55_1777 ();
 sg13g2_fill_1 FILLER_55_1779 ();
 sg13g2_fill_1 FILLER_55_1811 ();
 sg13g2_fill_2 FILLER_55_1860 ();
 sg13g2_decap_4 FILLER_55_1926 ();
 sg13g2_fill_1 FILLER_55_1930 ();
 sg13g2_fill_1 FILLER_55_1939 ();
 sg13g2_fill_1 FILLER_55_1971 ();
 sg13g2_fill_1 FILLER_55_2024 ();
 sg13g2_fill_2 FILLER_55_2145 ();
 sg13g2_fill_2 FILLER_55_2162 ();
 sg13g2_fill_1 FILLER_55_2164 ();
 sg13g2_fill_1 FILLER_55_2195 ();
 sg13g2_fill_2 FILLER_55_2229 ();
 sg13g2_fill_1 FILLER_55_2231 ();
 sg13g2_fill_2 FILLER_55_2280 ();
 sg13g2_fill_1 FILLER_55_2282 ();
 sg13g2_fill_1 FILLER_55_2364 ();
 sg13g2_fill_2 FILLER_55_2379 ();
 sg13g2_fill_2 FILLER_55_2406 ();
 sg13g2_fill_1 FILLER_55_2421 ();
 sg13g2_fill_2 FILLER_55_2566 ();
 sg13g2_fill_1 FILLER_55_2568 ();
 sg13g2_fill_2 FILLER_55_2595 ();
 sg13g2_decap_8 FILLER_55_2633 ();
 sg13g2_decap_8 FILLER_55_2640 ();
 sg13g2_decap_8 FILLER_55_2647 ();
 sg13g2_decap_8 FILLER_55_2654 ();
 sg13g2_decap_8 FILLER_55_2661 ();
 sg13g2_decap_4 FILLER_55_2668 ();
 sg13g2_fill_2 FILLER_55_2672 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_4 FILLER_56_35 ();
 sg13g2_fill_1 FILLER_56_65 ();
 sg13g2_fill_2 FILLER_56_170 ();
 sg13g2_fill_2 FILLER_56_272 ();
 sg13g2_fill_1 FILLER_56_310 ();
 sg13g2_fill_2 FILLER_56_350 ();
 sg13g2_fill_1 FILLER_56_383 ();
 sg13g2_fill_1 FILLER_56_435 ();
 sg13g2_fill_2 FILLER_56_441 ();
 sg13g2_fill_1 FILLER_56_443 ();
 sg13g2_fill_2 FILLER_56_453 ();
 sg13g2_fill_1 FILLER_56_455 ();
 sg13g2_fill_2 FILLER_56_519 ();
 sg13g2_fill_1 FILLER_56_521 ();
 sg13g2_fill_1 FILLER_56_575 ();
 sg13g2_fill_1 FILLER_56_650 ();
 sg13g2_fill_1 FILLER_56_676 ();
 sg13g2_fill_1 FILLER_56_694 ();
 sg13g2_fill_1 FILLER_56_701 ();
 sg13g2_fill_2 FILLER_56_757 ();
 sg13g2_fill_2 FILLER_56_785 ();
 sg13g2_fill_1 FILLER_56_787 ();
 sg13g2_fill_2 FILLER_56_877 ();
 sg13g2_fill_1 FILLER_56_879 ();
 sg13g2_fill_2 FILLER_56_890 ();
 sg13g2_fill_1 FILLER_56_1017 ();
 sg13g2_fill_1 FILLER_56_1027 ();
 sg13g2_fill_1 FILLER_56_1072 ();
 sg13g2_fill_1 FILLER_56_1126 ();
 sg13g2_fill_2 FILLER_56_1198 ();
 sg13g2_fill_1 FILLER_56_1261 ();
 sg13g2_fill_1 FILLER_56_1289 ();
 sg13g2_fill_2 FILLER_56_1376 ();
 sg13g2_fill_1 FILLER_56_1385 ();
 sg13g2_fill_2 FILLER_56_1405 ();
 sg13g2_fill_1 FILLER_56_1416 ();
 sg13g2_fill_2 FILLER_56_1502 ();
 sg13g2_fill_1 FILLER_56_1504 ();
 sg13g2_fill_2 FILLER_56_1521 ();
 sg13g2_fill_2 FILLER_56_1541 ();
 sg13g2_fill_1 FILLER_56_1543 ();
 sg13g2_fill_2 FILLER_56_1558 ();
 sg13g2_fill_1 FILLER_56_1560 ();
 sg13g2_decap_8 FILLER_56_1566 ();
 sg13g2_decap_8 FILLER_56_1573 ();
 sg13g2_fill_2 FILLER_56_1580 ();
 sg13g2_fill_1 FILLER_56_1582 ();
 sg13g2_decap_4 FILLER_56_1606 ();
 sg13g2_fill_1 FILLER_56_1622 ();
 sg13g2_fill_1 FILLER_56_1692 ();
 sg13g2_fill_1 FILLER_56_1734 ();
 sg13g2_fill_1 FILLER_56_1748 ();
 sg13g2_fill_1 FILLER_56_1785 ();
 sg13g2_fill_2 FILLER_56_1857 ();
 sg13g2_fill_1 FILLER_56_1859 ();
 sg13g2_decap_4 FILLER_56_1883 ();
 sg13g2_fill_1 FILLER_56_1887 ();
 sg13g2_fill_1 FILLER_56_1908 ();
 sg13g2_decap_4 FILLER_56_1931 ();
 sg13g2_fill_2 FILLER_56_1935 ();
 sg13g2_fill_1 FILLER_56_2030 ();
 sg13g2_fill_1 FILLER_56_2075 ();
 sg13g2_fill_1 FILLER_56_2097 ();
 sg13g2_fill_2 FILLER_56_2163 ();
 sg13g2_fill_1 FILLER_56_2258 ();
 sg13g2_fill_2 FILLER_56_2289 ();
 sg13g2_fill_2 FILLER_56_2343 ();
 sg13g2_fill_2 FILLER_56_2392 ();
 sg13g2_fill_1 FILLER_56_2436 ();
 sg13g2_fill_1 FILLER_56_2457 ();
 sg13g2_fill_1 FILLER_56_2537 ();
 sg13g2_fill_2 FILLER_56_2552 ();
 sg13g2_fill_1 FILLER_56_2564 ();
 sg13g2_fill_2 FILLER_56_2596 ();
 sg13g2_decap_8 FILLER_56_2637 ();
 sg13g2_decap_8 FILLER_56_2644 ();
 sg13g2_decap_8 FILLER_56_2651 ();
 sg13g2_decap_8 FILLER_56_2658 ();
 sg13g2_decap_8 FILLER_56_2665 ();
 sg13g2_fill_2 FILLER_56_2672 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_fill_1 FILLER_57_42 ();
 sg13g2_fill_2 FILLER_57_108 ();
 sg13g2_fill_2 FILLER_57_119 ();
 sg13g2_fill_1 FILLER_57_148 ();
 sg13g2_fill_2 FILLER_57_175 ();
 sg13g2_fill_1 FILLER_57_187 ();
 sg13g2_fill_2 FILLER_57_219 ();
 sg13g2_fill_2 FILLER_57_334 ();
 sg13g2_fill_2 FILLER_57_396 ();
 sg13g2_fill_1 FILLER_57_463 ();
 sg13g2_fill_1 FILLER_57_505 ();
 sg13g2_fill_1 FILLER_57_538 ();
 sg13g2_fill_2 FILLER_57_627 ();
 sg13g2_fill_2 FILLER_57_641 ();
 sg13g2_fill_1 FILLER_57_643 ();
 sg13g2_fill_2 FILLER_57_649 ();
 sg13g2_fill_1 FILLER_57_660 ();
 sg13g2_fill_2 FILLER_57_667 ();
 sg13g2_fill_1 FILLER_57_669 ();
 sg13g2_fill_2 FILLER_57_688 ();
 sg13g2_fill_1 FILLER_57_690 ();
 sg13g2_fill_2 FILLER_57_743 ();
 sg13g2_fill_2 FILLER_57_796 ();
 sg13g2_fill_1 FILLER_57_813 ();
 sg13g2_fill_1 FILLER_57_829 ();
 sg13g2_fill_2 FILLER_57_866 ();
 sg13g2_fill_1 FILLER_57_868 ();
 sg13g2_fill_1 FILLER_57_895 ();
 sg13g2_fill_1 FILLER_57_930 ();
 sg13g2_fill_2 FILLER_57_983 ();
 sg13g2_fill_1 FILLER_57_985 ();
 sg13g2_fill_1 FILLER_57_1003 ();
 sg13g2_fill_1 FILLER_57_1031 ();
 sg13g2_fill_2 FILLER_57_1056 ();
 sg13g2_fill_1 FILLER_57_1103 ();
 sg13g2_fill_1 FILLER_57_1121 ();
 sg13g2_fill_1 FILLER_57_1132 ();
 sg13g2_fill_1 FILLER_57_1190 ();
 sg13g2_fill_2 FILLER_57_1232 ();
 sg13g2_decap_4 FILLER_57_1563 ();
 sg13g2_fill_2 FILLER_57_1605 ();
 sg13g2_fill_1 FILLER_57_1633 ();
 sg13g2_fill_1 FILLER_57_1664 ();
 sg13g2_fill_2 FILLER_57_1704 ();
 sg13g2_fill_1 FILLER_57_1706 ();
 sg13g2_fill_2 FILLER_57_1745 ();
 sg13g2_fill_1 FILLER_57_1768 ();
 sg13g2_fill_2 FILLER_57_1827 ();
 sg13g2_decap_4 FILLER_57_1871 ();
 sg13g2_fill_2 FILLER_57_1894 ();
 sg13g2_fill_1 FILLER_57_1896 ();
 sg13g2_decap_4 FILLER_57_1907 ();
 sg13g2_fill_1 FILLER_57_1911 ();
 sg13g2_decap_4 FILLER_57_1923 ();
 sg13g2_fill_1 FILLER_57_1927 ();
 sg13g2_decap_8 FILLER_57_1934 ();
 sg13g2_decap_4 FILLER_57_1941 ();
 sg13g2_fill_1 FILLER_57_1945 ();
 sg13g2_fill_2 FILLER_57_2039 ();
 sg13g2_fill_1 FILLER_57_2041 ();
 sg13g2_fill_2 FILLER_57_2139 ();
 sg13g2_fill_1 FILLER_57_2141 ();
 sg13g2_fill_2 FILLER_57_2190 ();
 sg13g2_fill_2 FILLER_57_2279 ();
 sg13g2_fill_1 FILLER_57_2360 ();
 sg13g2_fill_1 FILLER_57_2397 ();
 sg13g2_fill_1 FILLER_57_2443 ();
 sg13g2_fill_2 FILLER_57_2526 ();
 sg13g2_fill_1 FILLER_57_2554 ();
 sg13g2_fill_1 FILLER_57_2565 ();
 sg13g2_fill_2 FILLER_57_2606 ();
 sg13g2_fill_1 FILLER_57_2608 ();
 sg13g2_decap_8 FILLER_57_2639 ();
 sg13g2_decap_8 FILLER_57_2646 ();
 sg13g2_decap_8 FILLER_57_2653 ();
 sg13g2_decap_8 FILLER_57_2660 ();
 sg13g2_decap_8 FILLER_57_2667 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_4 FILLER_58_35 ();
 sg13g2_fill_2 FILLER_58_39 ();
 sg13g2_fill_1 FILLER_58_96 ();
 sg13g2_fill_1 FILLER_58_170 ();
 sg13g2_fill_1 FILLER_58_176 ();
 sg13g2_fill_2 FILLER_58_259 ();
 sg13g2_fill_1 FILLER_58_287 ();
 sg13g2_fill_2 FILLER_58_342 ();
 sg13g2_fill_1 FILLER_58_380 ();
 sg13g2_fill_1 FILLER_58_390 ();
 sg13g2_fill_2 FILLER_58_401 ();
 sg13g2_fill_1 FILLER_58_403 ();
 sg13g2_fill_2 FILLER_58_436 ();
 sg13g2_fill_1 FILLER_58_438 ();
 sg13g2_fill_1 FILLER_58_634 ();
 sg13g2_fill_2 FILLER_58_665 ();
 sg13g2_fill_2 FILLER_58_750 ();
 sg13g2_fill_2 FILLER_58_788 ();
 sg13g2_fill_2 FILLER_58_809 ();
 sg13g2_fill_1 FILLER_58_811 ();
 sg13g2_fill_2 FILLER_58_935 ();
 sg13g2_fill_2 FILLER_58_967 ();
 sg13g2_fill_1 FILLER_58_1009 ();
 sg13g2_fill_2 FILLER_58_1061 ();
 sg13g2_fill_1 FILLER_58_1063 ();
 sg13g2_fill_2 FILLER_58_1119 ();
 sg13g2_fill_1 FILLER_58_1121 ();
 sg13g2_fill_1 FILLER_58_1165 ();
 sg13g2_fill_2 FILLER_58_1188 ();
 sg13g2_fill_1 FILLER_58_1283 ();
 sg13g2_fill_1 FILLER_58_1357 ();
 sg13g2_fill_1 FILLER_58_1459 ();
 sg13g2_fill_2 FILLER_58_1476 ();
 sg13g2_fill_1 FILLER_58_1478 ();
 sg13g2_fill_2 FILLER_58_1506 ();
 sg13g2_fill_1 FILLER_58_1524 ();
 sg13g2_fill_2 FILLER_58_1557 ();
 sg13g2_fill_2 FILLER_58_1577 ();
 sg13g2_fill_1 FILLER_58_1579 ();
 sg13g2_fill_2 FILLER_58_1587 ();
 sg13g2_fill_1 FILLER_58_1589 ();
 sg13g2_fill_2 FILLER_58_1620 ();
 sg13g2_fill_2 FILLER_58_1667 ();
 sg13g2_fill_1 FILLER_58_1702 ();
 sg13g2_fill_2 FILLER_58_1755 ();
 sg13g2_fill_2 FILLER_58_1793 ();
 sg13g2_fill_1 FILLER_58_1799 ();
 sg13g2_fill_2 FILLER_58_1838 ();
 sg13g2_fill_2 FILLER_58_1852 ();
 sg13g2_fill_1 FILLER_58_1854 ();
 sg13g2_fill_2 FILLER_58_1861 ();
 sg13g2_fill_1 FILLER_58_1872 ();
 sg13g2_fill_2 FILLER_58_1892 ();
 sg13g2_fill_2 FILLER_58_1899 ();
 sg13g2_fill_1 FILLER_58_1901 ();
 sg13g2_decap_4 FILLER_58_1915 ();
 sg13g2_decap_4 FILLER_58_1924 ();
 sg13g2_fill_2 FILLER_58_1928 ();
 sg13g2_fill_2 FILLER_58_1994 ();
 sg13g2_fill_1 FILLER_58_1996 ();
 sg13g2_fill_2 FILLER_58_2006 ();
 sg13g2_fill_1 FILLER_58_2008 ();
 sg13g2_fill_1 FILLER_58_2013 ();
 sg13g2_fill_2 FILLER_58_2024 ();
 sg13g2_fill_1 FILLER_58_2026 ();
 sg13g2_fill_2 FILLER_58_2068 ();
 sg13g2_fill_1 FILLER_58_2070 ();
 sg13g2_fill_1 FILLER_58_2106 ();
 sg13g2_fill_2 FILLER_58_2131 ();
 sg13g2_fill_2 FILLER_58_2159 ();
 sg13g2_fill_1 FILLER_58_2167 ();
 sg13g2_fill_2 FILLER_58_2194 ();
 sg13g2_fill_1 FILLER_58_2196 ();
 sg13g2_fill_2 FILLER_58_2207 ();
 sg13g2_fill_1 FILLER_58_2209 ();
 sg13g2_fill_1 FILLER_58_2219 ();
 sg13g2_fill_1 FILLER_58_2264 ();
 sg13g2_fill_2 FILLER_58_2288 ();
 sg13g2_fill_1 FILLER_58_2290 ();
 sg13g2_fill_2 FILLER_58_2352 ();
 sg13g2_fill_2 FILLER_58_2390 ();
 sg13g2_fill_2 FILLER_58_2431 ();
 sg13g2_fill_2 FILLER_58_2546 ();
 sg13g2_fill_1 FILLER_58_2587 ();
 sg13g2_decap_8 FILLER_58_2641 ();
 sg13g2_decap_8 FILLER_58_2648 ();
 sg13g2_decap_8 FILLER_58_2655 ();
 sg13g2_decap_8 FILLER_58_2662 ();
 sg13g2_decap_4 FILLER_58_2669 ();
 sg13g2_fill_1 FILLER_58_2673 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_fill_2 FILLER_59_35 ();
 sg13g2_fill_1 FILLER_59_37 ();
 sg13g2_fill_1 FILLER_59_151 ();
 sg13g2_fill_1 FILLER_59_157 ();
 sg13g2_fill_2 FILLER_59_178 ();
 sg13g2_fill_2 FILLER_59_227 ();
 sg13g2_fill_1 FILLER_59_314 ();
 sg13g2_fill_1 FILLER_59_376 ();
 sg13g2_fill_2 FILLER_59_435 ();
 sg13g2_fill_1 FILLER_59_473 ();
 sg13g2_fill_2 FILLER_59_509 ();
 sg13g2_fill_1 FILLER_59_511 ();
 sg13g2_fill_1 FILLER_59_538 ();
 sg13g2_fill_2 FILLER_59_621 ();
 sg13g2_fill_2 FILLER_59_640 ();
 sg13g2_fill_1 FILLER_59_642 ();
 sg13g2_fill_1 FILLER_59_679 ();
 sg13g2_fill_2 FILLER_59_692 ();
 sg13g2_fill_2 FILLER_59_819 ();
 sg13g2_fill_1 FILLER_59_821 ();
 sg13g2_fill_2 FILLER_59_848 ();
 sg13g2_fill_1 FILLER_59_881 ();
 sg13g2_fill_2 FILLER_59_914 ();
 sg13g2_fill_2 FILLER_59_929 ();
 sg13g2_fill_1 FILLER_59_931 ();
 sg13g2_fill_1 FILLER_59_972 ();
 sg13g2_fill_2 FILLER_59_983 ();
 sg13g2_fill_2 FILLER_59_1073 ();
 sg13g2_fill_1 FILLER_59_1085 ();
 sg13g2_fill_1 FILLER_59_1095 ();
 sg13g2_fill_2 FILLER_59_1101 ();
 sg13g2_fill_1 FILLER_59_1103 ();
 sg13g2_fill_1 FILLER_59_1137 ();
 sg13g2_fill_2 FILLER_59_1148 ();
 sg13g2_fill_1 FILLER_59_1150 ();
 sg13g2_fill_1 FILLER_59_1213 ();
 sg13g2_fill_1 FILLER_59_1297 ();
 sg13g2_fill_1 FILLER_59_1411 ();
 sg13g2_fill_2 FILLER_59_1537 ();
 sg13g2_fill_1 FILLER_59_1559 ();
 sg13g2_fill_2 FILLER_59_1576 ();
 sg13g2_fill_1 FILLER_59_1638 ();
 sg13g2_fill_2 FILLER_59_1649 ();
 sg13g2_fill_1 FILLER_59_1660 ();
 sg13g2_fill_2 FILLER_59_1726 ();
 sg13g2_fill_1 FILLER_59_1728 ();
 sg13g2_fill_2 FILLER_59_1753 ();
 sg13g2_fill_1 FILLER_59_1755 ();
 sg13g2_decap_4 FILLER_59_1868 ();
 sg13g2_fill_1 FILLER_59_1884 ();
 sg13g2_fill_1 FILLER_59_1890 ();
 sg13g2_fill_2 FILLER_59_1897 ();
 sg13g2_fill_1 FILLER_59_1933 ();
 sg13g2_decap_4 FILLER_59_1955 ();
 sg13g2_fill_1 FILLER_59_1959 ();
 sg13g2_decap_4 FILLER_59_1964 ();
 sg13g2_fill_1 FILLER_59_1968 ();
 sg13g2_fill_1 FILLER_59_2014 ();
 sg13g2_fill_2 FILLER_59_2033 ();
 sg13g2_fill_1 FILLER_59_2104 ();
 sg13g2_fill_1 FILLER_59_2145 ();
 sg13g2_fill_2 FILLER_59_2159 ();
 sg13g2_fill_1 FILLER_59_2191 ();
 sg13g2_fill_2 FILLER_59_2228 ();
 sg13g2_fill_2 FILLER_59_2246 ();
 sg13g2_fill_1 FILLER_59_2248 ();
 sg13g2_fill_1 FILLER_59_2343 ();
 sg13g2_fill_2 FILLER_59_2390 ();
 sg13g2_fill_1 FILLER_59_2425 ();
 sg13g2_fill_1 FILLER_59_2473 ();
 sg13g2_fill_2 FILLER_59_2601 ();
 sg13g2_fill_1 FILLER_59_2603 ();
 sg13g2_decap_8 FILLER_59_2630 ();
 sg13g2_decap_8 FILLER_59_2637 ();
 sg13g2_decap_8 FILLER_59_2644 ();
 sg13g2_decap_8 FILLER_59_2651 ();
 sg13g2_decap_8 FILLER_59_2658 ();
 sg13g2_decap_8 FILLER_59_2665 ();
 sg13g2_fill_2 FILLER_59_2672 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_fill_2 FILLER_60_28 ();
 sg13g2_fill_2 FILLER_60_79 ();
 sg13g2_fill_2 FILLER_60_89 ();
 sg13g2_fill_2 FILLER_60_160 ();
 sg13g2_fill_1 FILLER_60_192 ();
 sg13g2_fill_2 FILLER_60_219 ();
 sg13g2_fill_1 FILLER_60_347 ();
 sg13g2_fill_1 FILLER_60_358 ();
 sg13g2_fill_2 FILLER_60_388 ();
 sg13g2_fill_2 FILLER_60_398 ();
 sg13g2_fill_2 FILLER_60_422 ();
 sg13g2_fill_2 FILLER_60_449 ();
 sg13g2_fill_1 FILLER_60_451 ();
 sg13g2_fill_2 FILLER_60_466 ();
 sg13g2_fill_1 FILLER_60_468 ();
 sg13g2_fill_2 FILLER_60_475 ();
 sg13g2_fill_1 FILLER_60_500 ();
 sg13g2_fill_2 FILLER_60_510 ();
 sg13g2_fill_2 FILLER_60_521 ();
 sg13g2_fill_1 FILLER_60_523 ();
 sg13g2_fill_2 FILLER_60_581 ();
 sg13g2_fill_1 FILLER_60_583 ();
 sg13g2_fill_1 FILLER_60_649 ();
 sg13g2_fill_1 FILLER_60_672 ();
 sg13g2_fill_2 FILLER_60_711 ();
 sg13g2_fill_1 FILLER_60_765 ();
 sg13g2_fill_2 FILLER_60_797 ();
 sg13g2_fill_2 FILLER_60_837 ();
 sg13g2_fill_2 FILLER_60_896 ();
 sg13g2_fill_2 FILLER_60_932 ();
 sg13g2_fill_2 FILLER_60_938 ();
 sg13g2_fill_1 FILLER_60_940 ();
 sg13g2_fill_1 FILLER_60_979 ();
 sg13g2_fill_2 FILLER_60_991 ();
 sg13g2_fill_2 FILLER_60_1015 ();
 sg13g2_fill_1 FILLER_60_1178 ();
 sg13g2_fill_1 FILLER_60_1197 ();
 sg13g2_fill_2 FILLER_60_1238 ();
 sg13g2_fill_1 FILLER_60_1240 ();
 sg13g2_fill_1 FILLER_60_1249 ();
 sg13g2_fill_1 FILLER_60_1263 ();
 sg13g2_fill_2 FILLER_60_1349 ();
 sg13g2_fill_1 FILLER_60_1360 ();
 sg13g2_fill_1 FILLER_60_1411 ();
 sg13g2_fill_1 FILLER_60_1429 ();
 sg13g2_fill_1 FILLER_60_1444 ();
 sg13g2_fill_2 FILLER_60_1476 ();
 sg13g2_fill_2 FILLER_60_1517 ();
 sg13g2_fill_1 FILLER_60_1519 ();
 sg13g2_fill_2 FILLER_60_1560 ();
 sg13g2_decap_4 FILLER_60_1583 ();
 sg13g2_decap_4 FILLER_60_1591 ();
 sg13g2_fill_2 FILLER_60_1595 ();
 sg13g2_fill_1 FILLER_60_1680 ();
 sg13g2_fill_2 FILLER_60_1710 ();
 sg13g2_fill_1 FILLER_60_1712 ();
 sg13g2_fill_1 FILLER_60_1722 ();
 sg13g2_fill_2 FILLER_60_1811 ();
 sg13g2_fill_1 FILLER_60_1855 ();
 sg13g2_fill_1 FILLER_60_1877 ();
 sg13g2_fill_1 FILLER_60_1888 ();
 sg13g2_fill_2 FILLER_60_1899 ();
 sg13g2_fill_1 FILLER_60_1901 ();
 sg13g2_fill_2 FILLER_60_1914 ();
 sg13g2_fill_1 FILLER_60_1916 ();
 sg13g2_decap_4 FILLER_60_1931 ();
 sg13g2_fill_1 FILLER_60_1935 ();
 sg13g2_fill_2 FILLER_60_1941 ();
 sg13g2_fill_1 FILLER_60_1959 ();
 sg13g2_fill_1 FILLER_60_1965 ();
 sg13g2_decap_4 FILLER_60_1975 ();
 sg13g2_fill_1 FILLER_60_2014 ();
 sg13g2_fill_2 FILLER_60_2118 ();
 sg13g2_fill_1 FILLER_60_2187 ();
 sg13g2_fill_2 FILLER_60_2194 ();
 sg13g2_fill_1 FILLER_60_2237 ();
 sg13g2_fill_2 FILLER_60_2276 ();
 sg13g2_fill_2 FILLER_60_2354 ();
 sg13g2_fill_1 FILLER_60_2356 ();
 sg13g2_fill_1 FILLER_60_2398 ();
 sg13g2_fill_2 FILLER_60_2435 ();
 sg13g2_fill_2 FILLER_60_2443 ();
 sg13g2_fill_1 FILLER_60_2454 ();
 sg13g2_fill_2 FILLER_60_2465 ();
 sg13g2_fill_1 FILLER_60_2475 ();
 sg13g2_fill_1 FILLER_60_2538 ();
 sg13g2_fill_1 FILLER_60_2567 ();
 sg13g2_fill_2 FILLER_60_2582 ();
 sg13g2_fill_1 FILLER_60_2584 ();
 sg13g2_decap_8 FILLER_60_2635 ();
 sg13g2_decap_8 FILLER_60_2642 ();
 sg13g2_decap_8 FILLER_60_2649 ();
 sg13g2_decap_8 FILLER_60_2656 ();
 sg13g2_decap_8 FILLER_60_2663 ();
 sg13g2_decap_4 FILLER_60_2670 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_4 FILLER_61_35 ();
 sg13g2_fill_1 FILLER_61_39 ();
 sg13g2_fill_1 FILLER_61_60 ();
 sg13g2_fill_1 FILLER_61_87 ();
 sg13g2_fill_1 FILLER_61_157 ();
 sg13g2_fill_1 FILLER_61_163 ();
 sg13g2_fill_1 FILLER_61_182 ();
 sg13g2_fill_2 FILLER_61_188 ();
 sg13g2_fill_1 FILLER_61_249 ();
 sg13g2_fill_2 FILLER_61_276 ();
 sg13g2_fill_2 FILLER_61_326 ();
 sg13g2_fill_1 FILLER_61_328 ();
 sg13g2_fill_2 FILLER_61_333 ();
 sg13g2_fill_1 FILLER_61_335 ();
 sg13g2_fill_2 FILLER_61_367 ();
 sg13g2_fill_2 FILLER_61_388 ();
 sg13g2_fill_1 FILLER_61_425 ();
 sg13g2_fill_2 FILLER_61_452 ();
 sg13g2_fill_2 FILLER_61_480 ();
 sg13g2_fill_2 FILLER_61_516 ();
 sg13g2_fill_1 FILLER_61_518 ();
 sg13g2_fill_1 FILLER_61_529 ();
 sg13g2_fill_1 FILLER_61_559 ();
 sg13g2_fill_1 FILLER_61_579 ();
 sg13g2_fill_2 FILLER_61_590 ();
 sg13g2_fill_1 FILLER_61_592 ();
 sg13g2_fill_1 FILLER_61_615 ();
 sg13g2_fill_2 FILLER_61_636 ();
 sg13g2_fill_1 FILLER_61_638 ();
 sg13g2_fill_1 FILLER_61_683 ();
 sg13g2_fill_1 FILLER_61_690 ();
 sg13g2_fill_2 FILLER_61_717 ();
 sg13g2_fill_1 FILLER_61_729 ();
 sg13g2_fill_2 FILLER_61_748 ();
 sg13g2_fill_1 FILLER_61_750 ();
 sg13g2_fill_1 FILLER_61_795 ();
 sg13g2_fill_2 FILLER_61_822 ();
 sg13g2_fill_2 FILLER_61_873 ();
 sg13g2_fill_1 FILLER_61_875 ();
 sg13g2_fill_2 FILLER_61_922 ();
 sg13g2_fill_2 FILLER_61_983 ();
 sg13g2_fill_1 FILLER_61_985 ();
 sg13g2_fill_2 FILLER_61_1039 ();
 sg13g2_fill_1 FILLER_61_1041 ();
 sg13g2_fill_2 FILLER_61_1072 ();
 sg13g2_fill_1 FILLER_61_1103 ();
 sg13g2_fill_1 FILLER_61_1121 ();
 sg13g2_fill_1 FILLER_61_1191 ();
 sg13g2_fill_2 FILLER_61_1245 ();
 sg13g2_fill_2 FILLER_61_1270 ();
 sg13g2_fill_1 FILLER_61_1286 ();
 sg13g2_fill_2 FILLER_61_1330 ();
 sg13g2_decap_4 FILLER_61_1342 ();
 sg13g2_fill_1 FILLER_61_1346 ();
 sg13g2_fill_1 FILLER_61_1372 ();
 sg13g2_fill_2 FILLER_61_1412 ();
 sg13g2_fill_2 FILLER_61_1423 ();
 sg13g2_fill_2 FILLER_61_1434 ();
 sg13g2_fill_2 FILLER_61_1461 ();
 sg13g2_fill_2 FILLER_61_1526 ();
 sg13g2_fill_1 FILLER_61_1575 ();
 sg13g2_fill_2 FILLER_61_1729 ();
 sg13g2_fill_1 FILLER_61_1840 ();
 sg13g2_fill_1 FILLER_61_1852 ();
 sg13g2_fill_1 FILLER_61_1876 ();
 sg13g2_fill_1 FILLER_61_1882 ();
 sg13g2_decap_4 FILLER_61_1935 ();
 sg13g2_fill_1 FILLER_61_1962 ();
 sg13g2_decap_4 FILLER_61_1980 ();
 sg13g2_fill_1 FILLER_61_1988 ();
 sg13g2_fill_2 FILLER_61_2015 ();
 sg13g2_fill_1 FILLER_61_2017 ();
 sg13g2_fill_1 FILLER_61_2072 ();
 sg13g2_fill_2 FILLER_61_2086 ();
 sg13g2_fill_1 FILLER_61_2088 ();
 sg13g2_fill_2 FILLER_61_2130 ();
 sg13g2_fill_2 FILLER_61_2161 ();
 sg13g2_fill_1 FILLER_61_2163 ();
 sg13g2_fill_1 FILLER_61_2173 ();
 sg13g2_fill_2 FILLER_61_2187 ();
 sg13g2_fill_1 FILLER_61_2189 ();
 sg13g2_fill_1 FILLER_61_2207 ();
 sg13g2_fill_1 FILLER_61_2246 ();
 sg13g2_fill_1 FILLER_61_2273 ();
 sg13g2_fill_2 FILLER_61_2278 ();
 sg13g2_fill_1 FILLER_61_2288 ();
 sg13g2_fill_2 FILLER_61_2314 ();
 sg13g2_fill_1 FILLER_61_2326 ();
 sg13g2_fill_2 FILLER_61_2385 ();
 sg13g2_fill_1 FILLER_61_2435 ();
 sg13g2_fill_1 FILLER_61_2472 ();
 sg13g2_fill_2 FILLER_61_2539 ();
 sg13g2_fill_1 FILLER_61_2541 ();
 sg13g2_fill_2 FILLER_61_2572 ();
 sg13g2_fill_1 FILLER_61_2574 ();
 sg13g2_fill_2 FILLER_61_2596 ();
 sg13g2_fill_1 FILLER_61_2598 ();
 sg13g2_decap_8 FILLER_61_2625 ();
 sg13g2_decap_8 FILLER_61_2632 ();
 sg13g2_decap_8 FILLER_61_2639 ();
 sg13g2_decap_8 FILLER_61_2646 ();
 sg13g2_decap_8 FILLER_61_2653 ();
 sg13g2_decap_8 FILLER_61_2660 ();
 sg13g2_decap_8 FILLER_61_2667 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_4 FILLER_62_21 ();
 sg13g2_fill_1 FILLER_62_25 ();
 sg13g2_fill_1 FILLER_62_66 ();
 sg13g2_fill_1 FILLER_62_90 ();
 sg13g2_fill_1 FILLER_62_101 ();
 sg13g2_fill_1 FILLER_62_173 ();
 sg13g2_fill_1 FILLER_62_204 ();
 sg13g2_fill_2 FILLER_62_218 ();
 sg13g2_fill_2 FILLER_62_230 ();
 sg13g2_fill_1 FILLER_62_246 ();
 sg13g2_fill_2 FILLER_62_275 ();
 sg13g2_fill_1 FILLER_62_296 ();
 sg13g2_fill_1 FILLER_62_316 ();
 sg13g2_fill_2 FILLER_62_396 ();
 sg13g2_fill_1 FILLER_62_398 ();
 sg13g2_fill_1 FILLER_62_417 ();
 sg13g2_fill_2 FILLER_62_443 ();
 sg13g2_fill_1 FILLER_62_454 ();
 sg13g2_fill_2 FILLER_62_517 ();
 sg13g2_fill_2 FILLER_62_580 ();
 sg13g2_fill_1 FILLER_62_612 ();
 sg13g2_fill_2 FILLER_62_631 ();
 sg13g2_fill_1 FILLER_62_633 ();
 sg13g2_fill_2 FILLER_62_673 ();
 sg13g2_fill_1 FILLER_62_675 ();
 sg13g2_fill_2 FILLER_62_705 ();
 sg13g2_fill_1 FILLER_62_707 ();
 sg13g2_fill_1 FILLER_62_719 ();
 sg13g2_fill_1 FILLER_62_827 ();
 sg13g2_fill_1 FILLER_62_837 ();
 sg13g2_fill_2 FILLER_62_847 ();
 sg13g2_fill_1 FILLER_62_891 ();
 sg13g2_fill_2 FILLER_62_909 ();
 sg13g2_fill_1 FILLER_62_958 ();
 sg13g2_fill_2 FILLER_62_980 ();
 sg13g2_fill_2 FILLER_62_1022 ();
 sg13g2_fill_1 FILLER_62_1059 ();
 sg13g2_fill_2 FILLER_62_1138 ();
 sg13g2_fill_1 FILLER_62_1140 ();
 sg13g2_fill_1 FILLER_62_1180 ();
 sg13g2_decap_4 FILLER_62_1225 ();
 sg13g2_fill_2 FILLER_62_1308 ();
 sg13g2_fill_1 FILLER_62_1325 ();
 sg13g2_fill_2 FILLER_62_1338 ();
 sg13g2_fill_1 FILLER_62_1406 ();
 sg13g2_fill_2 FILLER_62_1456 ();
 sg13g2_fill_2 FILLER_62_1468 ();
 sg13g2_fill_2 FILLER_62_1481 ();
 sg13g2_fill_2 FILLER_62_1534 ();
 sg13g2_fill_2 FILLER_62_1554 ();
 sg13g2_fill_2 FILLER_62_1669 ();
 sg13g2_fill_1 FILLER_62_1671 ();
 sg13g2_fill_2 FILLER_62_1702 ();
 sg13g2_fill_1 FILLER_62_1704 ();
 sg13g2_fill_2 FILLER_62_1754 ();
 sg13g2_fill_1 FILLER_62_1756 ();
 sg13g2_fill_2 FILLER_62_1772 ();
 sg13g2_fill_1 FILLER_62_1774 ();
 sg13g2_fill_2 FILLER_62_1823 ();
 sg13g2_fill_2 FILLER_62_1835 ();
 sg13g2_fill_1 FILLER_62_1837 ();
 sg13g2_decap_4 FILLER_62_1887 ();
 sg13g2_fill_1 FILLER_62_1899 ();
 sg13g2_fill_1 FILLER_62_1920 ();
 sg13g2_fill_2 FILLER_62_1950 ();
 sg13g2_fill_1 FILLER_62_1952 ();
 sg13g2_decap_4 FILLER_62_1958 ();
 sg13g2_decap_4 FILLER_62_1978 ();
 sg13g2_fill_2 FILLER_62_2008 ();
 sg13g2_fill_1 FILLER_62_2020 ();
 sg13g2_fill_1 FILLER_62_2118 ();
 sg13g2_fill_2 FILLER_62_2170 ();
 sg13g2_fill_1 FILLER_62_2277 ();
 sg13g2_fill_1 FILLER_62_2334 ();
 sg13g2_fill_2 FILLER_62_2368 ();
 sg13g2_fill_1 FILLER_62_2370 ();
 sg13g2_fill_1 FILLER_62_2380 ();
 sg13g2_fill_1 FILLER_62_2399 ();
 sg13g2_fill_1 FILLER_62_2410 ();
 sg13g2_fill_2 FILLER_62_2434 ();
 sg13g2_fill_2 FILLER_62_2484 ();
 sg13g2_fill_1 FILLER_62_2491 ();
 sg13g2_fill_2 FILLER_62_2501 ();
 sg13g2_fill_1 FILLER_62_2503 ();
 sg13g2_fill_2 FILLER_62_2527 ();
 sg13g2_fill_1 FILLER_62_2529 ();
 sg13g2_fill_2 FILLER_62_2581 ();
 sg13g2_decap_8 FILLER_62_2622 ();
 sg13g2_decap_8 FILLER_62_2629 ();
 sg13g2_decap_8 FILLER_62_2636 ();
 sg13g2_decap_8 FILLER_62_2643 ();
 sg13g2_decap_8 FILLER_62_2650 ();
 sg13g2_decap_8 FILLER_62_2657 ();
 sg13g2_decap_8 FILLER_62_2664 ();
 sg13g2_fill_2 FILLER_62_2671 ();
 sg13g2_fill_1 FILLER_62_2673 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_fill_1 FILLER_63_35 ();
 sg13g2_fill_1 FILLER_63_94 ();
 sg13g2_fill_1 FILLER_63_179 ();
 sg13g2_fill_2 FILLER_63_238 ();
 sg13g2_fill_1 FILLER_63_266 ();
 sg13g2_fill_1 FILLER_63_298 ();
 sg13g2_fill_2 FILLER_63_339 ();
 sg13g2_fill_1 FILLER_63_421 ();
 sg13g2_fill_1 FILLER_63_441 ();
 sg13g2_fill_2 FILLER_63_472 ();
 sg13g2_fill_1 FILLER_63_474 ();
 sg13g2_fill_1 FILLER_63_485 ();
 sg13g2_fill_2 FILLER_63_520 ();
 sg13g2_fill_2 FILLER_63_532 ();
 sg13g2_fill_1 FILLER_63_534 ();
 sg13g2_fill_1 FILLER_63_587 ();
 sg13g2_fill_2 FILLER_63_598 ();
 sg13g2_fill_1 FILLER_63_600 ();
 sg13g2_fill_2 FILLER_63_624 ();
 sg13g2_fill_1 FILLER_63_626 ();
 sg13g2_fill_1 FILLER_63_650 ();
 sg13g2_fill_1 FILLER_63_900 ();
 sg13g2_fill_1 FILLER_63_962 ();
 sg13g2_fill_2 FILLER_63_968 ();
 sg13g2_fill_1 FILLER_63_970 ();
 sg13g2_fill_2 FILLER_63_976 ();
 sg13g2_fill_1 FILLER_63_978 ();
 sg13g2_fill_1 FILLER_63_1046 ();
 sg13g2_fill_2 FILLER_63_1052 ();
 sg13g2_fill_1 FILLER_63_1068 ();
 sg13g2_fill_1 FILLER_63_1090 ();
 sg13g2_fill_2 FILLER_63_1096 ();
 sg13g2_fill_1 FILLER_63_1115 ();
 sg13g2_fill_1 FILLER_63_1121 ();
 sg13g2_fill_2 FILLER_63_1145 ();
 sg13g2_fill_1 FILLER_63_1147 ();
 sg13g2_fill_2 FILLER_63_1154 ();
 sg13g2_fill_2 FILLER_63_1175 ();
 sg13g2_fill_2 FILLER_63_1191 ();
 sg13g2_fill_1 FILLER_63_1193 ();
 sg13g2_fill_2 FILLER_63_1235 ();
 sg13g2_fill_1 FILLER_63_1237 ();
 sg13g2_fill_2 FILLER_63_1248 ();
 sg13g2_fill_2 FILLER_63_1275 ();
 sg13g2_fill_1 FILLER_63_1317 ();
 sg13g2_fill_1 FILLER_63_1329 ();
 sg13g2_fill_1 FILLER_63_1348 ();
 sg13g2_fill_2 FILLER_63_1367 ();
 sg13g2_decap_8 FILLER_63_1385 ();
 sg13g2_fill_1 FILLER_63_1392 ();
 sg13g2_fill_2 FILLER_63_1396 ();
 sg13g2_fill_1 FILLER_63_1398 ();
 sg13g2_fill_2 FILLER_63_1403 ();
 sg13g2_fill_1 FILLER_63_1415 ();
 sg13g2_fill_1 FILLER_63_1437 ();
 sg13g2_fill_1 FILLER_63_1486 ();
 sg13g2_fill_1 FILLER_63_1584 ();
 sg13g2_fill_2 FILLER_63_1590 ();
 sg13g2_fill_1 FILLER_63_1623 ();
 sg13g2_fill_2 FILLER_63_1637 ();
 sg13g2_fill_1 FILLER_63_1639 ();
 sg13g2_fill_2 FILLER_63_1722 ();
 sg13g2_fill_1 FILLER_63_1798 ();
 sg13g2_fill_2 FILLER_63_1817 ();
 sg13g2_fill_2 FILLER_63_1833 ();
 sg13g2_fill_1 FILLER_63_1835 ();
 sg13g2_fill_2 FILLER_63_1840 ();
 sg13g2_fill_2 FILLER_63_1847 ();
 sg13g2_fill_1 FILLER_63_1849 ();
 sg13g2_fill_2 FILLER_63_1861 ();
 sg13g2_fill_1 FILLER_63_1863 ();
 sg13g2_decap_8 FILLER_63_1869 ();
 sg13g2_fill_2 FILLER_63_1876 ();
 sg13g2_fill_2 FILLER_63_1901 ();
 sg13g2_fill_2 FILLER_63_1949 ();
 sg13g2_fill_2 FILLER_63_1979 ();
 sg13g2_fill_1 FILLER_63_1981 ();
 sg13g2_fill_2 FILLER_63_2008 ();
 sg13g2_decap_4 FILLER_63_2020 ();
 sg13g2_fill_1 FILLER_63_2024 ();
 sg13g2_fill_1 FILLER_63_2049 ();
 sg13g2_fill_2 FILLER_63_2110 ();
 sg13g2_fill_2 FILLER_63_2139 ();
 sg13g2_fill_1 FILLER_63_2177 ();
 sg13g2_fill_1 FILLER_63_2210 ();
 sg13g2_fill_2 FILLER_63_2238 ();
 sg13g2_fill_1 FILLER_63_2250 ();
 sg13g2_fill_2 FILLER_63_2291 ();
 sg13g2_fill_1 FILLER_63_2333 ();
 sg13g2_fill_1 FILLER_63_2419 ();
 sg13g2_fill_2 FILLER_63_2471 ();
 sg13g2_fill_1 FILLER_63_2499 ();
 sg13g2_fill_2 FILLER_63_2540 ();
 sg13g2_fill_1 FILLER_63_2560 ();
 sg13g2_fill_1 FILLER_63_2575 ();
 sg13g2_fill_1 FILLER_63_2603 ();
 sg13g2_decap_8 FILLER_63_2625 ();
 sg13g2_decap_8 FILLER_63_2632 ();
 sg13g2_decap_8 FILLER_63_2639 ();
 sg13g2_decap_8 FILLER_63_2646 ();
 sg13g2_decap_8 FILLER_63_2653 ();
 sg13g2_decap_8 FILLER_63_2660 ();
 sg13g2_decap_8 FILLER_63_2667 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_fill_1 FILLER_64_107 ();
 sg13g2_fill_1 FILLER_64_174 ();
 sg13g2_fill_2 FILLER_64_194 ();
 sg13g2_fill_1 FILLER_64_210 ();
 sg13g2_fill_1 FILLER_64_278 ();
 sg13g2_fill_2 FILLER_64_296 ();
 sg13g2_fill_1 FILLER_64_298 ();
 sg13g2_fill_2 FILLER_64_309 ();
 sg13g2_fill_1 FILLER_64_311 ();
 sg13g2_fill_1 FILLER_64_320 ();
 sg13g2_fill_2 FILLER_64_339 ();
 sg13g2_fill_1 FILLER_64_341 ();
 sg13g2_fill_1 FILLER_64_419 ();
 sg13g2_fill_2 FILLER_64_455 ();
 sg13g2_fill_1 FILLER_64_457 ();
 sg13g2_fill_2 FILLER_64_467 ();
 sg13g2_fill_1 FILLER_64_593 ();
 sg13g2_fill_2 FILLER_64_655 ();
 sg13g2_fill_2 FILLER_64_676 ();
 sg13g2_fill_2 FILLER_64_766 ();
 sg13g2_fill_2 FILLER_64_789 ();
 sg13g2_fill_1 FILLER_64_806 ();
 sg13g2_fill_2 FILLER_64_826 ();
 sg13g2_fill_2 FILLER_64_854 ();
 sg13g2_fill_1 FILLER_64_865 ();
 sg13g2_fill_1 FILLER_64_881 ();
 sg13g2_fill_2 FILLER_64_898 ();
 sg13g2_fill_2 FILLER_64_915 ();
 sg13g2_fill_2 FILLER_64_1004 ();
 sg13g2_fill_1 FILLER_64_1006 ();
 sg13g2_fill_2 FILLER_64_1064 ();
 sg13g2_fill_2 FILLER_64_1071 ();
 sg13g2_fill_1 FILLER_64_1084 ();
 sg13g2_fill_2 FILLER_64_1095 ();
 sg13g2_fill_1 FILLER_64_1097 ();
 sg13g2_fill_2 FILLER_64_1113 ();
 sg13g2_fill_2 FILLER_64_1167 ();
 sg13g2_fill_1 FILLER_64_1175 ();
 sg13g2_fill_1 FILLER_64_1206 ();
 sg13g2_decap_4 FILLER_64_1233 ();
 sg13g2_fill_1 FILLER_64_1237 ();
 sg13g2_fill_1 FILLER_64_1249 ();
 sg13g2_decap_4 FILLER_64_1259 ();
 sg13g2_fill_1 FILLER_64_1263 ();
 sg13g2_fill_1 FILLER_64_1272 ();
 sg13g2_fill_1 FILLER_64_1287 ();
 sg13g2_fill_2 FILLER_64_1319 ();
 sg13g2_fill_2 FILLER_64_1329 ();
 sg13g2_fill_2 FILLER_64_1346 ();
 sg13g2_decap_8 FILLER_64_1362 ();
 sg13g2_fill_2 FILLER_64_1374 ();
 sg13g2_fill_1 FILLER_64_1376 ();
 sg13g2_fill_1 FILLER_64_1423 ();
 sg13g2_fill_1 FILLER_64_1429 ();
 sg13g2_fill_1 FILLER_64_1446 ();
 sg13g2_fill_1 FILLER_64_1486 ();
 sg13g2_fill_1 FILLER_64_1517 ();
 sg13g2_fill_1 FILLER_64_1524 ();
 sg13g2_fill_1 FILLER_64_1547 ();
 sg13g2_fill_1 FILLER_64_1575 ();
 sg13g2_fill_1 FILLER_64_1581 ();
 sg13g2_fill_2 FILLER_64_1608 ();
 sg13g2_fill_2 FILLER_64_1636 ();
 sg13g2_fill_1 FILLER_64_1638 ();
 sg13g2_fill_2 FILLER_64_1718 ();
 sg13g2_decap_4 FILLER_64_1787 ();
 sg13g2_fill_2 FILLER_64_1811 ();
 sg13g2_fill_2 FILLER_64_1867 ();
 sg13g2_fill_1 FILLER_64_1869 ();
 sg13g2_decap_4 FILLER_64_1880 ();
 sg13g2_fill_1 FILLER_64_1913 ();
 sg13g2_fill_1 FILLER_64_1928 ();
 sg13g2_fill_2 FILLER_64_1939 ();
 sg13g2_fill_2 FILLER_64_1963 ();
 sg13g2_fill_2 FILLER_64_1984 ();
 sg13g2_fill_2 FILLER_64_2179 ();
 sg13g2_fill_2 FILLER_64_2205 ();
 sg13g2_fill_1 FILLER_64_2299 ();
 sg13g2_fill_1 FILLER_64_2330 ();
 sg13g2_fill_2 FILLER_64_2466 ();
 sg13g2_fill_1 FILLER_64_2482 ();
 sg13g2_fill_2 FILLER_64_2539 ();
 sg13g2_fill_1 FILLER_64_2541 ();
 sg13g2_fill_2 FILLER_64_2546 ();
 sg13g2_decap_8 FILLER_64_2620 ();
 sg13g2_decap_8 FILLER_64_2627 ();
 sg13g2_decap_8 FILLER_64_2634 ();
 sg13g2_decap_8 FILLER_64_2641 ();
 sg13g2_decap_8 FILLER_64_2648 ();
 sg13g2_decap_8 FILLER_64_2655 ();
 sg13g2_decap_8 FILLER_64_2662 ();
 sg13g2_decap_4 FILLER_64_2669 ();
 sg13g2_fill_1 FILLER_64_2673 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_fill_1 FILLER_65_59 ();
 sg13g2_fill_2 FILLER_65_95 ();
 sg13g2_fill_2 FILLER_65_177 ();
 sg13g2_fill_1 FILLER_65_238 ();
 sg13g2_fill_1 FILLER_65_262 ();
 sg13g2_fill_2 FILLER_65_351 ();
 sg13g2_fill_1 FILLER_65_353 ();
 sg13g2_fill_1 FILLER_65_363 ();
 sg13g2_fill_2 FILLER_65_425 ();
 sg13g2_fill_1 FILLER_65_427 ();
 sg13g2_fill_2 FILLER_65_445 ();
 sg13g2_fill_1 FILLER_65_463 ();
 sg13g2_fill_2 FILLER_65_470 ();
 sg13g2_fill_1 FILLER_65_477 ();
 sg13g2_fill_2 FILLER_65_492 ();
 sg13g2_fill_1 FILLER_65_494 ();
 sg13g2_fill_1 FILLER_65_521 ();
 sg13g2_fill_1 FILLER_65_543 ();
 sg13g2_fill_2 FILLER_65_562 ();
 sg13g2_fill_2 FILLER_65_620 ();
 sg13g2_fill_2 FILLER_65_653 ();
 sg13g2_fill_2 FILLER_65_695 ();
 sg13g2_fill_1 FILLER_65_697 ();
 sg13g2_fill_2 FILLER_65_720 ();
 sg13g2_fill_2 FILLER_65_752 ();
 sg13g2_fill_1 FILLER_65_754 ();
 sg13g2_fill_1 FILLER_65_781 ();
 sg13g2_fill_2 FILLER_65_887 ();
 sg13g2_fill_1 FILLER_65_898 ();
 sg13g2_fill_2 FILLER_65_916 ();
 sg13g2_fill_2 FILLER_65_944 ();
 sg13g2_fill_1 FILLER_65_946 ();
 sg13g2_fill_1 FILLER_65_952 ();
 sg13g2_fill_2 FILLER_65_966 ();
 sg13g2_fill_2 FILLER_65_974 ();
 sg13g2_fill_1 FILLER_65_1012 ();
 sg13g2_fill_2 FILLER_65_1022 ();
 sg13g2_fill_1 FILLER_65_1024 ();
 sg13g2_fill_1 FILLER_65_1031 ();
 sg13g2_fill_2 FILLER_65_1074 ();
 sg13g2_fill_1 FILLER_65_1076 ();
 sg13g2_fill_2 FILLER_65_1083 ();
 sg13g2_fill_1 FILLER_65_1085 ();
 sg13g2_fill_1 FILLER_65_1121 ();
 sg13g2_fill_1 FILLER_65_1150 ();
 sg13g2_fill_2 FILLER_65_1172 ();
 sg13g2_fill_1 FILLER_65_1174 ();
 sg13g2_fill_2 FILLER_65_1180 ();
 sg13g2_fill_1 FILLER_65_1269 ();
 sg13g2_decap_4 FILLER_65_1275 ();
 sg13g2_fill_1 FILLER_65_1283 ();
 sg13g2_decap_4 FILLER_65_1303 ();
 sg13g2_fill_1 FILLER_65_1307 ();
 sg13g2_decap_4 FILLER_65_1353 ();
 sg13g2_fill_2 FILLER_65_1357 ();
 sg13g2_decap_8 FILLER_65_1386 ();
 sg13g2_fill_2 FILLER_65_1393 ();
 sg13g2_fill_1 FILLER_65_1395 ();
 sg13g2_fill_2 FILLER_65_1404 ();
 sg13g2_fill_1 FILLER_65_1406 ();
 sg13g2_fill_2 FILLER_65_1418 ();
 sg13g2_fill_2 FILLER_65_1492 ();
 sg13g2_fill_2 FILLER_65_1499 ();
 sg13g2_fill_1 FILLER_65_1518 ();
 sg13g2_fill_1 FILLER_65_1541 ();
 sg13g2_fill_1 FILLER_65_1564 ();
 sg13g2_fill_2 FILLER_65_1591 ();
 sg13g2_fill_1 FILLER_65_1593 ();
 sg13g2_fill_2 FILLER_65_1599 ();
 sg13g2_fill_1 FILLER_65_1601 ();
 sg13g2_decap_8 FILLER_65_1646 ();
 sg13g2_fill_2 FILLER_65_1653 ();
 sg13g2_fill_2 FILLER_65_1673 ();
 sg13g2_fill_2 FILLER_65_1688 ();
 sg13g2_fill_2 FILLER_65_1725 ();
 sg13g2_fill_1 FILLER_65_1727 ();
 sg13g2_fill_2 FILLER_65_1767 ();
 sg13g2_decap_8 FILLER_65_1782 ();
 sg13g2_fill_2 FILLER_65_1789 ();
 sg13g2_fill_1 FILLER_65_1838 ();
 sg13g2_fill_2 FILLER_65_1872 ();
 sg13g2_fill_1 FILLER_65_1874 ();
 sg13g2_fill_2 FILLER_65_1880 ();
 sg13g2_fill_1 FILLER_65_1886 ();
 sg13g2_fill_1 FILLER_65_1917 ();
 sg13g2_decap_4 FILLER_65_1923 ();
 sg13g2_fill_2 FILLER_65_1932 ();
 sg13g2_fill_2 FILLER_65_1939 ();
 sg13g2_fill_1 FILLER_65_1961 ();
 sg13g2_fill_1 FILLER_65_1967 ();
 sg13g2_decap_8 FILLER_65_1986 ();
 sg13g2_fill_1 FILLER_65_1993 ();
 sg13g2_decap_4 FILLER_65_2017 ();
 sg13g2_fill_2 FILLER_65_2021 ();
 sg13g2_decap_8 FILLER_65_2027 ();
 sg13g2_fill_1 FILLER_65_2053 ();
 sg13g2_fill_1 FILLER_65_2135 ();
 sg13g2_fill_2 FILLER_65_2146 ();
 sg13g2_fill_1 FILLER_65_2148 ();
 sg13g2_fill_2 FILLER_65_2191 ();
 sg13g2_fill_2 FILLER_65_2224 ();
 sg13g2_fill_1 FILLER_65_2226 ();
 sg13g2_fill_2 FILLER_65_2236 ();
 sg13g2_fill_1 FILLER_65_2257 ();
 sg13g2_fill_2 FILLER_65_2292 ();
 sg13g2_fill_1 FILLER_65_2294 ();
 sg13g2_fill_1 FILLER_65_2309 ();
 sg13g2_fill_2 FILLER_65_2350 ();
 sg13g2_fill_1 FILLER_65_2352 ();
 sg13g2_fill_1 FILLER_65_2431 ();
 sg13g2_fill_1 FILLER_65_2442 ();
 sg13g2_fill_2 FILLER_65_2527 ();
 sg13g2_fill_1 FILLER_65_2529 ();
 sg13g2_fill_1 FILLER_65_2574 ();
 sg13g2_decap_8 FILLER_65_2601 ();
 sg13g2_decap_8 FILLER_65_2608 ();
 sg13g2_decap_8 FILLER_65_2615 ();
 sg13g2_decap_8 FILLER_65_2622 ();
 sg13g2_decap_8 FILLER_65_2629 ();
 sg13g2_decap_8 FILLER_65_2636 ();
 sg13g2_decap_8 FILLER_65_2643 ();
 sg13g2_decap_8 FILLER_65_2650 ();
 sg13g2_decap_8 FILLER_65_2657 ();
 sg13g2_decap_8 FILLER_65_2664 ();
 sg13g2_fill_2 FILLER_65_2671 ();
 sg13g2_fill_1 FILLER_65_2673 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_fill_1 FILLER_66_42 ();
 sg13g2_fill_1 FILLER_66_120 ();
 sg13g2_fill_2 FILLER_66_206 ();
 sg13g2_fill_2 FILLER_66_285 ();
 sg13g2_fill_1 FILLER_66_314 ();
 sg13g2_fill_1 FILLER_66_320 ();
 sg13g2_fill_2 FILLER_66_375 ();
 sg13g2_fill_1 FILLER_66_377 ();
 sg13g2_fill_2 FILLER_66_398 ();
 sg13g2_fill_2 FILLER_66_426 ();
 sg13g2_fill_1 FILLER_66_428 ();
 sg13g2_fill_2 FILLER_66_507 ();
 sg13g2_fill_1 FILLER_66_509 ();
 sg13g2_fill_2 FILLER_66_546 ();
 sg13g2_fill_2 FILLER_66_584 ();
 sg13g2_fill_1 FILLER_66_596 ();
 sg13g2_fill_2 FILLER_66_614 ();
 sg13g2_fill_2 FILLER_66_657 ();
 sg13g2_fill_1 FILLER_66_727 ();
 sg13g2_fill_1 FILLER_66_737 ();
 sg13g2_fill_1 FILLER_66_748 ();
 sg13g2_fill_2 FILLER_66_795 ();
 sg13g2_fill_1 FILLER_66_797 ();
 sg13g2_fill_1 FILLER_66_812 ();
 sg13g2_fill_2 FILLER_66_839 ();
 sg13g2_fill_2 FILLER_66_873 ();
 sg13g2_fill_1 FILLER_66_875 ();
 sg13g2_fill_2 FILLER_66_937 ();
 sg13g2_fill_1 FILLER_66_1001 ();
 sg13g2_fill_2 FILLER_66_1088 ();
 sg13g2_fill_1 FILLER_66_1090 ();
 sg13g2_fill_2 FILLER_66_1096 ();
 sg13g2_fill_1 FILLER_66_1098 ();
 sg13g2_fill_2 FILLER_66_1176 ();
 sg13g2_fill_1 FILLER_66_1192 ();
 sg13g2_decap_4 FILLER_66_1213 ();
 sg13g2_fill_1 FILLER_66_1217 ();
 sg13g2_fill_1 FILLER_66_1222 ();
 sg13g2_fill_2 FILLER_66_1239 ();
 sg13g2_fill_1 FILLER_66_1241 ();
 sg13g2_fill_1 FILLER_66_1251 ();
 sg13g2_fill_2 FILLER_66_1272 ();
 sg13g2_fill_1 FILLER_66_1301 ();
 sg13g2_fill_2 FILLER_66_1319 ();
 sg13g2_fill_1 FILLER_66_1334 ();
 sg13g2_fill_1 FILLER_66_1345 ();
 sg13g2_fill_2 FILLER_66_1355 ();
 sg13g2_fill_1 FILLER_66_1370 ();
 sg13g2_decap_4 FILLER_66_1381 ();
 sg13g2_fill_2 FILLER_66_1391 ();
 sg13g2_fill_2 FILLER_66_1427 ();
 sg13g2_fill_1 FILLER_66_1433 ();
 sg13g2_fill_2 FILLER_66_1500 ();
 sg13g2_fill_1 FILLER_66_1502 ();
 sg13g2_fill_2 FILLER_66_1546 ();
 sg13g2_fill_2 FILLER_66_1609 ();
 sg13g2_fill_1 FILLER_66_1628 ();
 sg13g2_fill_1 FILLER_66_1754 ();
 sg13g2_fill_1 FILLER_66_1794 ();
 sg13g2_fill_1 FILLER_66_1839 ();
 sg13g2_fill_2 FILLER_66_1851 ();
 sg13g2_fill_2 FILLER_66_1868 ();
 sg13g2_fill_2 FILLER_66_1875 ();
 sg13g2_fill_1 FILLER_66_1877 ();
 sg13g2_decap_4 FILLER_66_1893 ();
 sg13g2_fill_2 FILLER_66_1913 ();
 sg13g2_fill_1 FILLER_66_1915 ();
 sg13g2_fill_2 FILLER_66_1921 ();
 sg13g2_fill_1 FILLER_66_1923 ();
 sg13g2_decap_4 FILLER_66_1944 ();
 sg13g2_fill_2 FILLER_66_1956 ();
 sg13g2_fill_2 FILLER_66_1963 ();
 sg13g2_fill_1 FILLER_66_1965 ();
 sg13g2_fill_2 FILLER_66_1971 ();
 sg13g2_fill_1 FILLER_66_1986 ();
 sg13g2_fill_2 FILLER_66_2065 ();
 sg13g2_fill_2 FILLER_66_2101 ();
 sg13g2_fill_2 FILLER_66_2113 ();
 sg13g2_fill_2 FILLER_66_2147 ();
 sg13g2_fill_2 FILLER_66_2190 ();
 sg13g2_fill_2 FILLER_66_2271 ();
 sg13g2_fill_2 FILLER_66_2327 ();
 sg13g2_fill_2 FILLER_66_2379 ();
 sg13g2_fill_1 FILLER_66_2381 ();
 sg13g2_fill_2 FILLER_66_2418 ();
 sg13g2_fill_1 FILLER_66_2420 ();
 sg13g2_fill_2 FILLER_66_2568 ();
 sg13g2_decap_8 FILLER_66_2578 ();
 sg13g2_decap_8 FILLER_66_2598 ();
 sg13g2_decap_8 FILLER_66_2605 ();
 sg13g2_decap_8 FILLER_66_2612 ();
 sg13g2_decap_8 FILLER_66_2619 ();
 sg13g2_decap_8 FILLER_66_2626 ();
 sg13g2_decap_8 FILLER_66_2633 ();
 sg13g2_decap_8 FILLER_66_2640 ();
 sg13g2_decap_8 FILLER_66_2647 ();
 sg13g2_decap_8 FILLER_66_2654 ();
 sg13g2_decap_8 FILLER_66_2661 ();
 sg13g2_decap_4 FILLER_66_2668 ();
 sg13g2_fill_2 FILLER_66_2672 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_4 FILLER_67_42 ();
 sg13g2_fill_1 FILLER_67_98 ();
 sg13g2_fill_2 FILLER_67_141 ();
 sg13g2_fill_2 FILLER_67_157 ();
 sg13g2_fill_2 FILLER_67_190 ();
 sg13g2_fill_1 FILLER_67_219 ();
 sg13g2_fill_2 FILLER_67_290 ();
 sg13g2_fill_2 FILLER_67_375 ();
 sg13g2_fill_1 FILLER_67_377 ();
 sg13g2_fill_1 FILLER_67_411 ();
 sg13g2_fill_1 FILLER_67_438 ();
 sg13g2_fill_2 FILLER_67_457 ();
 sg13g2_fill_1 FILLER_67_459 ();
 sg13g2_fill_1 FILLER_67_470 ();
 sg13g2_fill_1 FILLER_67_476 ();
 sg13g2_fill_2 FILLER_67_483 ();
 sg13g2_fill_1 FILLER_67_485 ();
 sg13g2_fill_1 FILLER_67_521 ();
 sg13g2_fill_2 FILLER_67_527 ();
 sg13g2_fill_1 FILLER_67_529 ();
 sg13g2_fill_1 FILLER_67_539 ();
 sg13g2_fill_2 FILLER_67_608 ();
 sg13g2_fill_1 FILLER_67_610 ();
 sg13g2_fill_2 FILLER_67_639 ();
 sg13g2_fill_2 FILLER_67_646 ();
 sg13g2_fill_1 FILLER_67_648 ();
 sg13g2_fill_2 FILLER_67_675 ();
 sg13g2_fill_2 FILLER_67_691 ();
 sg13g2_fill_2 FILLER_67_714 ();
 sg13g2_fill_1 FILLER_67_716 ();
 sg13g2_fill_2 FILLER_67_767 ();
 sg13g2_fill_1 FILLER_67_814 ();
 sg13g2_fill_2 FILLER_67_820 ();
 sg13g2_fill_1 FILLER_67_822 ();
 sg13g2_fill_1 FILLER_67_856 ();
 sg13g2_fill_1 FILLER_67_866 ();
 sg13g2_fill_1 FILLER_67_888 ();
 sg13g2_fill_1 FILLER_67_893 ();
 sg13g2_fill_2 FILLER_67_939 ();
 sg13g2_fill_1 FILLER_67_941 ();
 sg13g2_fill_2 FILLER_67_977 ();
 sg13g2_fill_1 FILLER_67_979 ();
 sg13g2_fill_2 FILLER_67_1002 ();
 sg13g2_fill_1 FILLER_67_1012 ();
 sg13g2_fill_1 FILLER_67_1022 ();
 sg13g2_fill_2 FILLER_67_1042 ();
 sg13g2_fill_1 FILLER_67_1044 ();
 sg13g2_fill_2 FILLER_67_1049 ();
 sg13g2_fill_1 FILLER_67_1051 ();
 sg13g2_fill_2 FILLER_67_1083 ();
 sg13g2_fill_1 FILLER_67_1085 ();
 sg13g2_fill_1 FILLER_67_1145 ();
 sg13g2_fill_2 FILLER_67_1166 ();
 sg13g2_decap_8 FILLER_67_1209 ();
 sg13g2_fill_2 FILLER_67_1220 ();
 sg13g2_fill_1 FILLER_67_1222 ();
 sg13g2_fill_2 FILLER_67_1262 ();
 sg13g2_fill_1 FILLER_67_1264 ();
 sg13g2_decap_8 FILLER_67_1275 ();
 sg13g2_fill_1 FILLER_67_1282 ();
 sg13g2_fill_2 FILLER_67_1296 ();
 sg13g2_decap_4 FILLER_67_1302 ();
 sg13g2_fill_1 FILLER_67_1306 ();
 sg13g2_decap_4 FILLER_67_1316 ();
 sg13g2_decap_4 FILLER_67_1334 ();
 sg13g2_fill_2 FILLER_67_1338 ();
 sg13g2_decap_8 FILLER_67_1360 ();
 sg13g2_fill_2 FILLER_67_1367 ();
 sg13g2_fill_1 FILLER_67_1369 ();
 sg13g2_decap_4 FILLER_67_1379 ();
 sg13g2_fill_2 FILLER_67_1383 ();
 sg13g2_fill_2 FILLER_67_1407 ();
 sg13g2_fill_2 FILLER_67_1418 ();
 sg13g2_fill_1 FILLER_67_1420 ();
 sg13g2_fill_1 FILLER_67_1441 ();
 sg13g2_fill_1 FILLER_67_1450 ();
 sg13g2_fill_2 FILLER_67_1497 ();
 sg13g2_fill_2 FILLER_67_1519 ();
 sg13g2_fill_2 FILLER_67_1536 ();
 sg13g2_fill_1 FILLER_67_1579 ();
 sg13g2_fill_2 FILLER_67_1631 ();
 sg13g2_fill_1 FILLER_67_1641 ();
 sg13g2_fill_2 FILLER_67_1657 ();
 sg13g2_fill_1 FILLER_67_1659 ();
 sg13g2_fill_1 FILLER_67_1674 ();
 sg13g2_fill_2 FILLER_67_1685 ();
 sg13g2_fill_2 FILLER_67_1769 ();
 sg13g2_fill_2 FILLER_67_1792 ();
 sg13g2_fill_1 FILLER_67_1794 ();
 sg13g2_decap_4 FILLER_67_1831 ();
 sg13g2_fill_1 FILLER_67_1835 ();
 sg13g2_fill_1 FILLER_67_1861 ();
 sg13g2_fill_2 FILLER_67_1884 ();
 sg13g2_fill_2 FILLER_67_1896 ();
 sg13g2_fill_2 FILLER_67_1906 ();
 sg13g2_fill_1 FILLER_67_1908 ();
 sg13g2_fill_2 FILLER_67_1983 ();
 sg13g2_fill_1 FILLER_67_1985 ();
 sg13g2_fill_1 FILLER_67_2026 ();
 sg13g2_fill_2 FILLER_67_2079 ();
 sg13g2_fill_1 FILLER_67_2081 ();
 sg13g2_fill_2 FILLER_67_2118 ();
 sg13g2_fill_1 FILLER_67_2120 ();
 sg13g2_fill_2 FILLER_67_2152 ();
 sg13g2_fill_2 FILLER_67_2229 ();
 sg13g2_fill_1 FILLER_67_2267 ();
 sg13g2_fill_2 FILLER_67_2299 ();
 sg13g2_fill_2 FILLER_67_2337 ();
 sg13g2_fill_1 FILLER_67_2348 ();
 sg13g2_fill_2 FILLER_67_2367 ();
 sg13g2_fill_2 FILLER_67_2418 ();
 sg13g2_fill_1 FILLER_67_2465 ();
 sg13g2_decap_4 FILLER_67_2559 ();
 sg13g2_fill_1 FILLER_67_2563 ();
 sg13g2_decap_8 FILLER_67_2568 ();
 sg13g2_decap_8 FILLER_67_2575 ();
 sg13g2_decap_8 FILLER_67_2582 ();
 sg13g2_decap_8 FILLER_67_2589 ();
 sg13g2_decap_8 FILLER_67_2596 ();
 sg13g2_decap_8 FILLER_67_2603 ();
 sg13g2_decap_8 FILLER_67_2610 ();
 sg13g2_decap_8 FILLER_67_2617 ();
 sg13g2_decap_8 FILLER_67_2624 ();
 sg13g2_decap_8 FILLER_67_2631 ();
 sg13g2_decap_8 FILLER_67_2638 ();
 sg13g2_decap_8 FILLER_67_2645 ();
 sg13g2_decap_8 FILLER_67_2652 ();
 sg13g2_decap_8 FILLER_67_2659 ();
 sg13g2_decap_8 FILLER_67_2666 ();
 sg13g2_fill_1 FILLER_67_2673 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_fill_1 FILLER_68_49 ();
 sg13g2_fill_1 FILLER_68_128 ();
 sg13g2_fill_2 FILLER_68_207 ();
 sg13g2_fill_1 FILLER_68_233 ();
 sg13g2_fill_1 FILLER_68_243 ();
 sg13g2_fill_1 FILLER_68_275 ();
 sg13g2_fill_2 FILLER_68_302 ();
 sg13g2_fill_2 FILLER_68_314 ();
 sg13g2_fill_2 FILLER_68_342 ();
 sg13g2_fill_1 FILLER_68_344 ();
 sg13g2_fill_2 FILLER_68_379 ();
 sg13g2_fill_1 FILLER_68_420 ();
 sg13g2_fill_2 FILLER_68_434 ();
 sg13g2_fill_2 FILLER_68_441 ();
 sg13g2_fill_1 FILLER_68_443 ();
 sg13g2_fill_2 FILLER_68_449 ();
 sg13g2_fill_1 FILLER_68_477 ();
 sg13g2_fill_1 FILLER_68_513 ();
 sg13g2_fill_2 FILLER_68_580 ();
 sg13g2_fill_1 FILLER_68_639 ();
 sg13g2_fill_1 FILLER_68_699 ();
 sg13g2_fill_1 FILLER_68_798 ();
 sg13g2_fill_1 FILLER_68_862 ();
 sg13g2_fill_1 FILLER_68_893 ();
 sg13g2_fill_2 FILLER_68_945 ();
 sg13g2_fill_1 FILLER_68_1020 ();
 sg13g2_fill_1 FILLER_68_1037 ();
 sg13g2_fill_1 FILLER_68_1047 ();
 sg13g2_fill_1 FILLER_68_1074 ();
 sg13g2_fill_2 FILLER_68_1099 ();
 sg13g2_fill_1 FILLER_68_1101 ();
 sg13g2_fill_1 FILLER_68_1173 ();
 sg13g2_fill_1 FILLER_68_1231 ();
 sg13g2_decap_4 FILLER_68_1273 ();
 sg13g2_fill_2 FILLER_68_1277 ();
 sg13g2_decap_8 FILLER_68_1309 ();
 sg13g2_fill_2 FILLER_68_1316 ();
 sg13g2_fill_2 FILLER_68_1336 ();
 sg13g2_fill_2 FILLER_68_1358 ();
 sg13g2_fill_2 FILLER_68_1368 ();
 sg13g2_fill_1 FILLER_68_1390 ();
 sg13g2_fill_2 FILLER_68_1407 ();
 sg13g2_fill_2 FILLER_68_1419 ();
 sg13g2_fill_1 FILLER_68_1440 ();
 sg13g2_fill_2 FILLER_68_1453 ();
 sg13g2_fill_1 FILLER_68_1455 ();
 sg13g2_fill_2 FILLER_68_1486 ();
 sg13g2_fill_2 FILLER_68_1507 ();
 sg13g2_fill_2 FILLER_68_1525 ();
 sg13g2_fill_1 FILLER_68_1554 ();
 sg13g2_fill_2 FILLER_68_1564 ();
 sg13g2_fill_1 FILLER_68_1566 ();
 sg13g2_fill_1 FILLER_68_1613 ();
 sg13g2_fill_1 FILLER_68_1658 ();
 sg13g2_fill_2 FILLER_68_1682 ();
 sg13g2_fill_1 FILLER_68_1684 ();
 sg13g2_fill_2 FILLER_68_1691 ();
 sg13g2_fill_1 FILLER_68_1693 ();
 sg13g2_fill_2 FILLER_68_1703 ();
 sg13g2_fill_2 FILLER_68_1749 ();
 sg13g2_fill_1 FILLER_68_1751 ();
 sg13g2_fill_1 FILLER_68_1834 ();
 sg13g2_fill_1 FILLER_68_1839 ();
 sg13g2_fill_2 FILLER_68_1853 ();
 sg13g2_decap_4 FILLER_68_1859 ();
 sg13g2_fill_1 FILLER_68_1867 ();
 sg13g2_fill_1 FILLER_68_1884 ();
 sg13g2_fill_1 FILLER_68_1898 ();
 sg13g2_decap_4 FILLER_68_1916 ();
 sg13g2_fill_2 FILLER_68_1920 ();
 sg13g2_fill_2 FILLER_68_1959 ();
 sg13g2_fill_1 FILLER_68_1961 ();
 sg13g2_fill_2 FILLER_68_1986 ();
 sg13g2_fill_1 FILLER_68_2044 ();
 sg13g2_fill_1 FILLER_68_2089 ();
 sg13g2_fill_2 FILLER_68_2099 ();
 sg13g2_fill_1 FILLER_68_2101 ();
 sg13g2_fill_2 FILLER_68_2107 ();
 sg13g2_fill_2 FILLER_68_2144 ();
 sg13g2_fill_2 FILLER_68_2208 ();
 sg13g2_fill_1 FILLER_68_2210 ();
 sg13g2_fill_2 FILLER_68_2232 ();
 sg13g2_fill_1 FILLER_68_2234 ();
 sg13g2_fill_1 FILLER_68_2245 ();
 sg13g2_fill_1 FILLER_68_2268 ();
 sg13g2_fill_2 FILLER_68_2292 ();
 sg13g2_fill_2 FILLER_68_2324 ();
 sg13g2_fill_2 FILLER_68_2335 ();
 sg13g2_fill_2 FILLER_68_2434 ();
 sg13g2_fill_2 FILLER_68_2544 ();
 sg13g2_decap_8 FILLER_68_2558 ();
 sg13g2_decap_8 FILLER_68_2565 ();
 sg13g2_decap_8 FILLER_68_2572 ();
 sg13g2_decap_8 FILLER_68_2579 ();
 sg13g2_decap_8 FILLER_68_2586 ();
 sg13g2_decap_8 FILLER_68_2593 ();
 sg13g2_decap_8 FILLER_68_2600 ();
 sg13g2_decap_8 FILLER_68_2607 ();
 sg13g2_decap_8 FILLER_68_2614 ();
 sg13g2_decap_8 FILLER_68_2621 ();
 sg13g2_decap_8 FILLER_68_2628 ();
 sg13g2_decap_8 FILLER_68_2635 ();
 sg13g2_decap_8 FILLER_68_2642 ();
 sg13g2_decap_8 FILLER_68_2649 ();
 sg13g2_decap_8 FILLER_68_2656 ();
 sg13g2_decap_8 FILLER_68_2663 ();
 sg13g2_decap_4 FILLER_68_2670 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_4 FILLER_69_49 ();
 sg13g2_fill_2 FILLER_69_53 ();
 sg13g2_fill_1 FILLER_69_118 ();
 sg13g2_fill_1 FILLER_69_148 ();
 sg13g2_fill_1 FILLER_69_206 ();
 sg13g2_fill_2 FILLER_69_237 ();
 sg13g2_fill_1 FILLER_69_249 ();
 sg13g2_fill_2 FILLER_69_309 ();
 sg13g2_fill_2 FILLER_69_321 ();
 sg13g2_fill_1 FILLER_69_436 ();
 sg13g2_fill_2 FILLER_69_451 ();
 sg13g2_fill_1 FILLER_69_468 ();
 sg13g2_fill_2 FILLER_69_503 ();
 sg13g2_fill_1 FILLER_69_505 ();
 sg13g2_fill_2 FILLER_69_515 ();
 sg13g2_fill_2 FILLER_69_590 ();
 sg13g2_fill_2 FILLER_69_615 ();
 sg13g2_fill_1 FILLER_69_617 ();
 sg13g2_fill_2 FILLER_69_634 ();
 sg13g2_fill_1 FILLER_69_716 ();
 sg13g2_fill_1 FILLER_69_777 ();
 sg13g2_fill_2 FILLER_69_786 ();
 sg13g2_fill_1 FILLER_69_871 ();
 sg13g2_fill_1 FILLER_69_944 ();
 sg13g2_fill_2 FILLER_69_968 ();
 sg13g2_fill_2 FILLER_69_1048 ();
 sg13g2_fill_2 FILLER_69_1121 ();
 sg13g2_fill_1 FILLER_69_1215 ();
 sg13g2_decap_8 FILLER_69_1270 ();
 sg13g2_fill_1 FILLER_69_1277 ();
 sg13g2_fill_2 FILLER_69_1320 ();
 sg13g2_decap_4 FILLER_69_1341 ();
 sg13g2_fill_1 FILLER_69_1345 ();
 sg13g2_fill_2 FILLER_69_1350 ();
 sg13g2_fill_1 FILLER_69_1352 ();
 sg13g2_decap_4 FILLER_69_1362 ();
 sg13g2_fill_2 FILLER_69_1366 ();
 sg13g2_decap_4 FILLER_69_1372 ();
 sg13g2_decap_4 FILLER_69_1394 ();
 sg13g2_fill_2 FILLER_69_1398 ();
 sg13g2_fill_2 FILLER_69_1413 ();
 sg13g2_fill_2 FILLER_69_1442 ();
 sg13g2_fill_1 FILLER_69_1482 ();
 sg13g2_fill_2 FILLER_69_1518 ();
 sg13g2_fill_1 FILLER_69_1525 ();
 sg13g2_fill_2 FILLER_69_1539 ();
 sg13g2_fill_2 FILLER_69_1546 ();
 sg13g2_fill_1 FILLER_69_1581 ();
 sg13g2_fill_1 FILLER_69_1609 ();
 sg13g2_fill_1 FILLER_69_1702 ();
 sg13g2_decap_4 FILLER_69_1790 ();
 sg13g2_decap_4 FILLER_69_1810 ();
 sg13g2_decap_4 FILLER_69_1824 ();
 sg13g2_fill_2 FILLER_69_1840 ();
 sg13g2_fill_1 FILLER_69_1877 ();
 sg13g2_fill_2 FILLER_69_1907 ();
 sg13g2_fill_1 FILLER_69_1909 ();
 sg13g2_fill_1 FILLER_69_1919 ();
 sg13g2_decap_4 FILLER_69_1934 ();
 sg13g2_fill_2 FILLER_69_2171 ();
 sg13g2_fill_1 FILLER_69_2173 ();
 sg13g2_fill_2 FILLER_69_2212 ();
 sg13g2_fill_2 FILLER_69_2284 ();
 sg13g2_fill_1 FILLER_69_2400 ();
 sg13g2_fill_2 FILLER_69_2429 ();
 sg13g2_fill_2 FILLER_69_2463 ();
 sg13g2_fill_1 FILLER_69_2475 ();
 sg13g2_fill_1 FILLER_69_2495 ();
 sg13g2_fill_1 FILLER_69_2506 ();
 sg13g2_decap_8 FILLER_69_2542 ();
 sg13g2_decap_8 FILLER_69_2549 ();
 sg13g2_decap_8 FILLER_69_2556 ();
 sg13g2_decap_8 FILLER_69_2563 ();
 sg13g2_decap_8 FILLER_69_2570 ();
 sg13g2_decap_8 FILLER_69_2577 ();
 sg13g2_decap_8 FILLER_69_2584 ();
 sg13g2_decap_8 FILLER_69_2591 ();
 sg13g2_decap_8 FILLER_69_2598 ();
 sg13g2_decap_8 FILLER_69_2605 ();
 sg13g2_decap_8 FILLER_69_2612 ();
 sg13g2_decap_8 FILLER_69_2619 ();
 sg13g2_decap_8 FILLER_69_2626 ();
 sg13g2_decap_8 FILLER_69_2633 ();
 sg13g2_decap_8 FILLER_69_2640 ();
 sg13g2_decap_8 FILLER_69_2647 ();
 sg13g2_decap_8 FILLER_69_2654 ();
 sg13g2_decap_8 FILLER_69_2661 ();
 sg13g2_decap_4 FILLER_69_2668 ();
 sg13g2_fill_2 FILLER_69_2672 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_4 FILLER_70_49 ();
 sg13g2_fill_2 FILLER_70_53 ();
 sg13g2_fill_1 FILLER_70_100 ();
 sg13g2_fill_2 FILLER_70_177 ();
 sg13g2_fill_1 FILLER_70_217 ();
 sg13g2_fill_1 FILLER_70_323 ();
 sg13g2_fill_1 FILLER_70_352 ();
 sg13g2_fill_1 FILLER_70_420 ();
 sg13g2_fill_1 FILLER_70_443 ();
 sg13g2_fill_2 FILLER_70_488 ();
 sg13g2_fill_1 FILLER_70_520 ();
 sg13g2_fill_2 FILLER_70_547 ();
 sg13g2_fill_1 FILLER_70_549 ();
 sg13g2_fill_2 FILLER_70_555 ();
 sg13g2_fill_2 FILLER_70_566 ();
 sg13g2_fill_1 FILLER_70_568 ();
 sg13g2_fill_2 FILLER_70_579 ();
 sg13g2_fill_1 FILLER_70_581 ();
 sg13g2_fill_1 FILLER_70_643 ();
 sg13g2_fill_2 FILLER_70_649 ();
 sg13g2_fill_1 FILLER_70_651 ();
 sg13g2_fill_2 FILLER_70_661 ();
 sg13g2_fill_2 FILLER_70_703 ();
 sg13g2_fill_1 FILLER_70_705 ();
 sg13g2_fill_2 FILLER_70_737 ();
 sg13g2_fill_2 FILLER_70_814 ();
 sg13g2_fill_2 FILLER_70_830 ();
 sg13g2_fill_2 FILLER_70_868 ();
 sg13g2_fill_1 FILLER_70_870 ();
 sg13g2_fill_2 FILLER_70_910 ();
 sg13g2_fill_2 FILLER_70_921 ();
 sg13g2_fill_1 FILLER_70_923 ();
 sg13g2_fill_2 FILLER_70_959 ();
 sg13g2_fill_2 FILLER_70_987 ();
 sg13g2_fill_1 FILLER_70_989 ();
 sg13g2_fill_2 FILLER_70_1002 ();
 sg13g2_fill_1 FILLER_70_1046 ();
 sg13g2_fill_1 FILLER_70_1056 ();
 sg13g2_fill_2 FILLER_70_1074 ();
 sg13g2_fill_1 FILLER_70_1076 ();
 sg13g2_fill_2 FILLER_70_1109 ();
 sg13g2_fill_1 FILLER_70_1111 ();
 sg13g2_fill_1 FILLER_70_1144 ();
 sg13g2_fill_2 FILLER_70_1204 ();
 sg13g2_fill_2 FILLER_70_1237 ();
 sg13g2_fill_1 FILLER_70_1294 ();
 sg13g2_decap_4 FILLER_70_1307 ();
 sg13g2_fill_1 FILLER_70_1311 ();
 sg13g2_fill_1 FILLER_70_1337 ();
 sg13g2_fill_2 FILLER_70_1368 ();
 sg13g2_fill_1 FILLER_70_1370 ();
 sg13g2_fill_2 FILLER_70_1392 ();
 sg13g2_decap_4 FILLER_70_1399 ();
 sg13g2_decap_4 FILLER_70_1422 ();
 sg13g2_fill_1 FILLER_70_1426 ();
 sg13g2_decap_4 FILLER_70_1436 ();
 sg13g2_fill_1 FILLER_70_1440 ();
 sg13g2_fill_2 FILLER_70_1445 ();
 sg13g2_fill_2 FILLER_70_1496 ();
 sg13g2_fill_1 FILLER_70_1511 ();
 sg13g2_fill_2 FILLER_70_1521 ();
 sg13g2_fill_1 FILLER_70_1523 ();
 sg13g2_fill_1 FILLER_70_1619 ();
 sg13g2_fill_1 FILLER_70_1638 ();
 sg13g2_fill_1 FILLER_70_1655 ();
 sg13g2_fill_1 FILLER_70_1680 ();
 sg13g2_fill_1 FILLER_70_1700 ();
 sg13g2_fill_2 FILLER_70_1710 ();
 sg13g2_fill_1 FILLER_70_1733 ();
 sg13g2_fill_1 FILLER_70_1750 ();
 sg13g2_fill_2 FILLER_70_1760 ();
 sg13g2_fill_2 FILLER_70_1783 ();
 sg13g2_decap_4 FILLER_70_1796 ();
 sg13g2_decap_8 FILLER_70_1805 ();
 sg13g2_fill_1 FILLER_70_1812 ();
 sg13g2_decap_4 FILLER_70_1831 ();
 sg13g2_fill_1 FILLER_70_1835 ();
 sg13g2_fill_2 FILLER_70_1845 ();
 sg13g2_fill_1 FILLER_70_1874 ();
 sg13g2_fill_2 FILLER_70_1911 ();
 sg13g2_fill_1 FILLER_70_1913 ();
 sg13g2_fill_1 FILLER_70_1920 ();
 sg13g2_fill_1 FILLER_70_1972 ();
 sg13g2_decap_8 FILLER_70_1977 ();
 sg13g2_fill_1 FILLER_70_1984 ();
 sg13g2_fill_2 FILLER_70_2052 ();
 sg13g2_fill_2 FILLER_70_2125 ();
 sg13g2_fill_2 FILLER_70_2156 ();
 sg13g2_fill_1 FILLER_70_2198 ();
 sg13g2_fill_1 FILLER_70_2256 ();
 sg13g2_fill_2 FILLER_70_2280 ();
 sg13g2_fill_1 FILLER_70_2298 ();
 sg13g2_fill_2 FILLER_70_2321 ();
 sg13g2_fill_2 FILLER_70_2364 ();
 sg13g2_fill_2 FILLER_70_2386 ();
 sg13g2_fill_1 FILLER_70_2445 ();
 sg13g2_fill_1 FILLER_70_2497 ();
 sg13g2_decap_8 FILLER_70_2543 ();
 sg13g2_decap_8 FILLER_70_2550 ();
 sg13g2_decap_8 FILLER_70_2557 ();
 sg13g2_decap_8 FILLER_70_2564 ();
 sg13g2_decap_8 FILLER_70_2571 ();
 sg13g2_decap_8 FILLER_70_2578 ();
 sg13g2_decap_8 FILLER_70_2585 ();
 sg13g2_decap_8 FILLER_70_2592 ();
 sg13g2_decap_8 FILLER_70_2599 ();
 sg13g2_decap_8 FILLER_70_2606 ();
 sg13g2_decap_8 FILLER_70_2613 ();
 sg13g2_decap_8 FILLER_70_2620 ();
 sg13g2_decap_8 FILLER_70_2627 ();
 sg13g2_decap_8 FILLER_70_2634 ();
 sg13g2_decap_8 FILLER_70_2641 ();
 sg13g2_decap_8 FILLER_70_2648 ();
 sg13g2_decap_8 FILLER_70_2655 ();
 sg13g2_decap_8 FILLER_70_2662 ();
 sg13g2_decap_4 FILLER_70_2669 ();
 sg13g2_fill_1 FILLER_70_2673 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_4 FILLER_71_56 ();
 sg13g2_fill_2 FILLER_71_60 ();
 sg13g2_fill_1 FILLER_71_132 ();
 sg13g2_fill_2 FILLER_71_188 ();
 sg13g2_fill_1 FILLER_71_190 ();
 sg13g2_fill_2 FILLER_71_196 ();
 sg13g2_fill_1 FILLER_71_198 ();
 sg13g2_fill_1 FILLER_71_252 ();
 sg13g2_fill_1 FILLER_71_279 ();
 sg13g2_fill_2 FILLER_71_312 ();
 sg13g2_fill_1 FILLER_71_314 ();
 sg13g2_fill_1 FILLER_71_320 ();
 sg13g2_fill_1 FILLER_71_367 ();
 sg13g2_fill_2 FILLER_71_427 ();
 sg13g2_fill_1 FILLER_71_442 ();
 sg13g2_fill_2 FILLER_71_473 ();
 sg13g2_fill_1 FILLER_71_489 ();
 sg13g2_fill_1 FILLER_71_508 ();
 sg13g2_fill_1 FILLER_71_532 ();
 sg13g2_fill_2 FILLER_71_548 ();
 sg13g2_fill_2 FILLER_71_618 ();
 sg13g2_fill_1 FILLER_71_620 ();
 sg13g2_fill_1 FILLER_71_627 ();
 sg13g2_fill_2 FILLER_71_648 ();
 sg13g2_fill_2 FILLER_71_753 ();
 sg13g2_fill_1 FILLER_71_764 ();
 sg13g2_fill_2 FILLER_71_790 ();
 sg13g2_fill_1 FILLER_71_792 ();
 sg13g2_fill_2 FILLER_71_806 ();
 sg13g2_fill_1 FILLER_71_808 ();
 sg13g2_fill_1 FILLER_71_858 ();
 sg13g2_fill_1 FILLER_71_867 ();
 sg13g2_fill_2 FILLER_71_928 ();
 sg13g2_fill_1 FILLER_71_930 ();
 sg13g2_fill_1 FILLER_71_939 ();
 sg13g2_fill_2 FILLER_71_975 ();
 sg13g2_fill_1 FILLER_71_994 ();
 sg13g2_fill_2 FILLER_71_1059 ();
 sg13g2_fill_2 FILLER_71_1071 ();
 sg13g2_fill_1 FILLER_71_1073 ();
 sg13g2_fill_1 FILLER_71_1099 ();
 sg13g2_fill_2 FILLER_71_1108 ();
 sg13g2_fill_2 FILLER_71_1158 ();
 sg13g2_fill_2 FILLER_71_1175 ();
 sg13g2_fill_1 FILLER_71_1177 ();
 sg13g2_fill_2 FILLER_71_1204 ();
 sg13g2_fill_1 FILLER_71_1232 ();
 sg13g2_decap_4 FILLER_71_1276 ();
 sg13g2_fill_2 FILLER_71_1280 ();
 sg13g2_decap_4 FILLER_71_1308 ();
 sg13g2_fill_2 FILLER_71_1312 ();
 sg13g2_decap_8 FILLER_71_1342 ();
 sg13g2_fill_1 FILLER_71_1355 ();
 sg13g2_fill_1 FILLER_71_1386 ();
 sg13g2_fill_2 FILLER_71_1395 ();
 sg13g2_fill_1 FILLER_71_1397 ();
 sg13g2_fill_1 FILLER_71_1429 ();
 sg13g2_fill_1 FILLER_71_1490 ();
 sg13g2_fill_2 FILLER_71_1563 ();
 sg13g2_fill_2 FILLER_71_1591 ();
 sg13g2_fill_1 FILLER_71_1612 ();
 sg13g2_fill_2 FILLER_71_1656 ();
 sg13g2_fill_2 FILLER_71_1675 ();
 sg13g2_fill_2 FILLER_71_1690 ();
 sg13g2_fill_1 FILLER_71_1692 ();
 sg13g2_fill_2 FILLER_71_1735 ();
 sg13g2_decap_4 FILLER_71_1766 ();
 sg13g2_fill_2 FILLER_71_1770 ();
 sg13g2_fill_2 FILLER_71_1784 ();
 sg13g2_fill_1 FILLER_71_1786 ();
 sg13g2_fill_2 FILLER_71_1795 ();
 sg13g2_fill_1 FILLER_71_1797 ();
 sg13g2_fill_2 FILLER_71_1804 ();
 sg13g2_fill_1 FILLER_71_1806 ();
 sg13g2_fill_1 FILLER_71_1834 ();
 sg13g2_fill_2 FILLER_71_1857 ();
 sg13g2_fill_2 FILLER_71_1875 ();
 sg13g2_fill_2 FILLER_71_1882 ();
 sg13g2_fill_2 FILLER_71_1892 ();
 sg13g2_fill_2 FILLER_71_1914 ();
 sg13g2_decap_8 FILLER_71_1943 ();
 sg13g2_decap_8 FILLER_71_1950 ();
 sg13g2_fill_1 FILLER_71_1962 ();
 sg13g2_fill_1 FILLER_71_1993 ();
 sg13g2_fill_2 FILLER_71_2023 ();
 sg13g2_fill_1 FILLER_71_2025 ();
 sg13g2_fill_2 FILLER_71_2061 ();
 sg13g2_fill_1 FILLER_71_2063 ();
 sg13g2_fill_2 FILLER_71_2107 ();
 sg13g2_fill_1 FILLER_71_2109 ();
 sg13g2_fill_2 FILLER_71_2136 ();
 sg13g2_fill_1 FILLER_71_2138 ();
 sg13g2_fill_2 FILLER_71_2165 ();
 sg13g2_fill_1 FILLER_71_2177 ();
 sg13g2_fill_1 FILLER_71_2191 ();
 sg13g2_fill_1 FILLER_71_2237 ();
 sg13g2_fill_1 FILLER_71_2248 ();
 sg13g2_fill_2 FILLER_71_2303 ();
 sg13g2_fill_1 FILLER_71_2331 ();
 sg13g2_fill_1 FILLER_71_2342 ();
 sg13g2_fill_2 FILLER_71_2392 ();
 sg13g2_fill_1 FILLER_71_2394 ();
 sg13g2_fill_2 FILLER_71_2431 ();
 sg13g2_fill_2 FILLER_71_2463 ();
 sg13g2_fill_2 FILLER_71_2479 ();
 sg13g2_fill_1 FILLER_71_2481 ();
 sg13g2_decap_8 FILLER_71_2534 ();
 sg13g2_decap_8 FILLER_71_2541 ();
 sg13g2_decap_8 FILLER_71_2548 ();
 sg13g2_decap_8 FILLER_71_2555 ();
 sg13g2_decap_8 FILLER_71_2562 ();
 sg13g2_decap_8 FILLER_71_2569 ();
 sg13g2_decap_8 FILLER_71_2576 ();
 sg13g2_decap_8 FILLER_71_2583 ();
 sg13g2_decap_8 FILLER_71_2590 ();
 sg13g2_decap_8 FILLER_71_2597 ();
 sg13g2_decap_8 FILLER_71_2604 ();
 sg13g2_decap_8 FILLER_71_2611 ();
 sg13g2_decap_8 FILLER_71_2618 ();
 sg13g2_decap_8 FILLER_71_2625 ();
 sg13g2_decap_8 FILLER_71_2632 ();
 sg13g2_decap_8 FILLER_71_2639 ();
 sg13g2_decap_8 FILLER_71_2646 ();
 sg13g2_decap_8 FILLER_71_2653 ();
 sg13g2_decap_8 FILLER_71_2660 ();
 sg13g2_decap_8 FILLER_71_2667 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_fill_2 FILLER_72_56 ();
 sg13g2_fill_1 FILLER_72_58 ();
 sg13g2_fill_1 FILLER_72_237 ();
 sg13g2_fill_1 FILLER_72_247 ();
 sg13g2_fill_2 FILLER_72_282 ();
 sg13g2_fill_1 FILLER_72_352 ();
 sg13g2_fill_1 FILLER_72_369 ();
 sg13g2_fill_2 FILLER_72_418 ();
 sg13g2_fill_1 FILLER_72_501 ();
 sg13g2_fill_2 FILLER_72_555 ();
 sg13g2_fill_1 FILLER_72_557 ();
 sg13g2_fill_1 FILLER_72_622 ();
 sg13g2_fill_2 FILLER_72_659 ();
 sg13g2_fill_1 FILLER_72_661 ();
 sg13g2_fill_2 FILLER_72_727 ();
 sg13g2_fill_2 FILLER_72_769 ();
 sg13g2_fill_2 FILLER_72_797 ();
 sg13g2_fill_1 FILLER_72_799 ();
 sg13g2_fill_2 FILLER_72_805 ();
 sg13g2_fill_1 FILLER_72_807 ();
 sg13g2_fill_2 FILLER_72_920 ();
 sg13g2_fill_2 FILLER_72_957 ();
 sg13g2_fill_2 FILLER_72_996 ();
 sg13g2_fill_2 FILLER_72_1025 ();
 sg13g2_fill_1 FILLER_72_1081 ();
 sg13g2_fill_2 FILLER_72_1153 ();
 sg13g2_fill_2 FILLER_72_1227 ();
 sg13g2_fill_1 FILLER_72_1229 ();
 sg13g2_fill_1 FILLER_72_1287 ();
 sg13g2_fill_2 FILLER_72_1296 ();
 sg13g2_decap_4 FILLER_72_1302 ();
 sg13g2_fill_2 FILLER_72_1325 ();
 sg13g2_fill_1 FILLER_72_1327 ();
 sg13g2_fill_2 FILLER_72_1333 ();
 sg13g2_fill_1 FILLER_72_1344 ();
 sg13g2_fill_2 FILLER_72_1349 ();
 sg13g2_fill_1 FILLER_72_1351 ();
 sg13g2_decap_4 FILLER_72_1375 ();
 sg13g2_fill_1 FILLER_72_1379 ();
 sg13g2_fill_2 FILLER_72_1385 ();
 sg13g2_fill_1 FILLER_72_1395 ();
 sg13g2_fill_1 FILLER_72_1414 ();
 sg13g2_decap_4 FILLER_72_1420 ();
 sg13g2_fill_1 FILLER_72_1424 ();
 sg13g2_decap_4 FILLER_72_1429 ();
 sg13g2_decap_4 FILLER_72_1438 ();
 sg13g2_fill_1 FILLER_72_1442 ();
 sg13g2_fill_2 FILLER_72_1450 ();
 sg13g2_fill_1 FILLER_72_1582 ();
 sg13g2_fill_1 FILLER_72_1593 ();
 sg13g2_fill_2 FILLER_72_1653 ();
 sg13g2_fill_1 FILLER_72_1712 ();
 sg13g2_fill_2 FILLER_72_1726 ();
 sg13g2_fill_1 FILLER_72_1728 ();
 sg13g2_decap_4 FILLER_72_1760 ();
 sg13g2_fill_1 FILLER_72_1764 ();
 sg13g2_fill_1 FILLER_72_1791 ();
 sg13g2_fill_2 FILLER_72_1804 ();
 sg13g2_fill_1 FILLER_72_1806 ();
 sg13g2_fill_2 FILLER_72_1812 ();
 sg13g2_fill_1 FILLER_72_1814 ();
 sg13g2_fill_2 FILLER_72_1839 ();
 sg13g2_fill_1 FILLER_72_1841 ();
 sg13g2_decap_4 FILLER_72_1851 ();
 sg13g2_fill_1 FILLER_72_1860 ();
 sg13g2_fill_1 FILLER_72_1873 ();
 sg13g2_fill_2 FILLER_72_1881 ();
 sg13g2_decap_8 FILLER_72_1896 ();
 sg13g2_fill_2 FILLER_72_1921 ();
 sg13g2_decap_4 FILLER_72_1927 ();
 sg13g2_fill_1 FILLER_72_1931 ();
 sg13g2_fill_2 FILLER_72_1969 ();
 sg13g2_fill_1 FILLER_72_2040 ();
 sg13g2_fill_1 FILLER_72_2141 ();
 sg13g2_fill_2 FILLER_72_2170 ();
 sg13g2_fill_2 FILLER_72_2198 ();
 sg13g2_fill_2 FILLER_72_2236 ();
 sg13g2_fill_2 FILLER_72_2297 ();
 sg13g2_fill_1 FILLER_72_2366 ();
 sg13g2_fill_1 FILLER_72_2407 ();
 sg13g2_fill_2 FILLER_72_2450 ();
 sg13g2_decap_8 FILLER_72_2537 ();
 sg13g2_decap_8 FILLER_72_2544 ();
 sg13g2_decap_8 FILLER_72_2551 ();
 sg13g2_decap_8 FILLER_72_2558 ();
 sg13g2_decap_8 FILLER_72_2565 ();
 sg13g2_decap_8 FILLER_72_2572 ();
 sg13g2_decap_8 FILLER_72_2579 ();
 sg13g2_decap_8 FILLER_72_2586 ();
 sg13g2_decap_8 FILLER_72_2593 ();
 sg13g2_decap_8 FILLER_72_2600 ();
 sg13g2_decap_8 FILLER_72_2607 ();
 sg13g2_decap_8 FILLER_72_2614 ();
 sg13g2_decap_8 FILLER_72_2621 ();
 sg13g2_decap_8 FILLER_72_2628 ();
 sg13g2_decap_8 FILLER_72_2635 ();
 sg13g2_decap_8 FILLER_72_2642 ();
 sg13g2_decap_8 FILLER_72_2649 ();
 sg13g2_decap_8 FILLER_72_2656 ();
 sg13g2_decap_8 FILLER_72_2663 ();
 sg13g2_decap_4 FILLER_72_2670 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_4 FILLER_73_70 ();
 sg13g2_fill_1 FILLER_73_132 ();
 sg13g2_fill_1 FILLER_73_142 ();
 sg13g2_fill_2 FILLER_73_183 ();
 sg13g2_fill_1 FILLER_73_185 ();
 sg13g2_fill_1 FILLER_73_196 ();
 sg13g2_fill_2 FILLER_73_206 ();
 sg13g2_fill_1 FILLER_73_215 ();
 sg13g2_fill_1 FILLER_73_229 ();
 sg13g2_fill_1 FILLER_73_296 ();
 sg13g2_fill_2 FILLER_73_421 ();
 sg13g2_fill_2 FILLER_73_569 ();
 sg13g2_fill_1 FILLER_73_580 ();
 sg13g2_fill_2 FILLER_73_590 ();
 sg13g2_fill_2 FILLER_73_711 ();
 sg13g2_fill_1 FILLER_73_713 ();
 sg13g2_fill_1 FILLER_73_771 ();
 sg13g2_fill_1 FILLER_73_778 ();
 sg13g2_fill_1 FILLER_73_797 ();
 sg13g2_fill_1 FILLER_73_833 ();
 sg13g2_fill_1 FILLER_73_848 ();
 sg13g2_fill_2 FILLER_73_858 ();
 sg13g2_fill_1 FILLER_73_860 ();
 sg13g2_fill_1 FILLER_73_885 ();
 sg13g2_fill_2 FILLER_73_914 ();
 sg13g2_fill_1 FILLER_73_916 ();
 sg13g2_fill_2 FILLER_73_934 ();
 sg13g2_fill_1 FILLER_73_940 ();
 sg13g2_fill_1 FILLER_73_976 ();
 sg13g2_fill_2 FILLER_73_1016 ();
 sg13g2_fill_2 FILLER_73_1058 ();
 sg13g2_fill_1 FILLER_73_1060 ();
 sg13g2_fill_1 FILLER_73_1086 ();
 sg13g2_fill_2 FILLER_73_1174 ();
 sg13g2_fill_1 FILLER_73_1176 ();
 sg13g2_fill_2 FILLER_73_1191 ();
 sg13g2_fill_2 FILLER_73_1307 ();
 sg13g2_decap_4 FILLER_73_1313 ();
 sg13g2_fill_2 FILLER_73_1338 ();
 sg13g2_fill_1 FILLER_73_1340 ();
 sg13g2_fill_2 FILLER_73_1361 ();
 sg13g2_fill_2 FILLER_73_1390 ();
 sg13g2_fill_1 FILLER_73_1392 ();
 sg13g2_fill_1 FILLER_73_1407 ();
 sg13g2_fill_1 FILLER_73_1433 ();
 sg13g2_fill_1 FILLER_73_1521 ();
 sg13g2_fill_1 FILLER_73_1561 ();
 sg13g2_fill_1 FILLER_73_1598 ();
 sg13g2_fill_2 FILLER_73_1639 ();
 sg13g2_fill_2 FILLER_73_1660 ();
 sg13g2_fill_1 FILLER_73_1687 ();
 sg13g2_fill_2 FILLER_73_1734 ();
 sg13g2_decap_4 FILLER_73_1753 ();
 sg13g2_decap_8 FILLER_73_1774 ();
 sg13g2_fill_1 FILLER_73_1781 ();
 sg13g2_fill_2 FILLER_73_1800 ();
 sg13g2_fill_1 FILLER_73_1836 ();
 sg13g2_decap_8 FILLER_73_1849 ();
 sg13g2_decap_8 FILLER_73_1856 ();
 sg13g2_fill_2 FILLER_73_1863 ();
 sg13g2_decap_4 FILLER_73_1882 ();
 sg13g2_fill_1 FILLER_73_1886 ();
 sg13g2_decap_8 FILLER_73_1891 ();
 sg13g2_fill_1 FILLER_73_1898 ();
 sg13g2_decap_8 FILLER_73_1903 ();
 sg13g2_fill_2 FILLER_73_1910 ();
 sg13g2_fill_1 FILLER_73_1912 ();
 sg13g2_fill_1 FILLER_73_1917 ();
 sg13g2_decap_8 FILLER_73_1938 ();
 sg13g2_decap_4 FILLER_73_1945 ();
 sg13g2_fill_2 FILLER_73_1958 ();
 sg13g2_fill_1 FILLER_73_1960 ();
 sg13g2_fill_1 FILLER_73_1975 ();
 sg13g2_fill_2 FILLER_73_1989 ();
 sg13g2_fill_1 FILLER_73_1991 ();
 sg13g2_fill_1 FILLER_73_2017 ();
 sg13g2_fill_2 FILLER_73_2036 ();
 sg13g2_fill_2 FILLER_73_2043 ();
 sg13g2_fill_1 FILLER_73_2045 ();
 sg13g2_fill_2 FILLER_73_2209 ();
 sg13g2_fill_1 FILLER_73_2211 ();
 sg13g2_fill_1 FILLER_73_2363 ();
 sg13g2_fill_2 FILLER_73_2409 ();
 sg13g2_fill_1 FILLER_73_2420 ();
 sg13g2_fill_2 FILLER_73_2434 ();
 sg13g2_fill_1 FILLER_73_2436 ();
 sg13g2_fill_2 FILLER_73_2454 ();
 sg13g2_decap_8 FILLER_73_2536 ();
 sg13g2_decap_8 FILLER_73_2543 ();
 sg13g2_decap_8 FILLER_73_2550 ();
 sg13g2_decap_8 FILLER_73_2557 ();
 sg13g2_decap_8 FILLER_73_2564 ();
 sg13g2_decap_8 FILLER_73_2571 ();
 sg13g2_decap_8 FILLER_73_2578 ();
 sg13g2_decap_8 FILLER_73_2585 ();
 sg13g2_decap_8 FILLER_73_2592 ();
 sg13g2_decap_8 FILLER_73_2599 ();
 sg13g2_decap_8 FILLER_73_2606 ();
 sg13g2_decap_8 FILLER_73_2613 ();
 sg13g2_decap_8 FILLER_73_2620 ();
 sg13g2_decap_8 FILLER_73_2627 ();
 sg13g2_decap_8 FILLER_73_2634 ();
 sg13g2_decap_8 FILLER_73_2641 ();
 sg13g2_decap_8 FILLER_73_2648 ();
 sg13g2_decap_8 FILLER_73_2655 ();
 sg13g2_decap_8 FILLER_73_2662 ();
 sg13g2_decap_4 FILLER_73_2669 ();
 sg13g2_fill_1 FILLER_73_2673 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_fill_2 FILLER_74_77 ();
 sg13g2_fill_1 FILLER_74_79 ();
 sg13g2_fill_1 FILLER_74_171 ();
 sg13g2_fill_2 FILLER_74_212 ();
 sg13g2_fill_1 FILLER_74_229 ();
 sg13g2_fill_2 FILLER_74_235 ();
 sg13g2_fill_2 FILLER_74_242 ();
 sg13g2_fill_2 FILLER_74_311 ();
 sg13g2_fill_1 FILLER_74_319 ();
 sg13g2_fill_1 FILLER_74_329 ();
 sg13g2_fill_1 FILLER_74_446 ();
 sg13g2_fill_2 FILLER_74_506 ();
 sg13g2_fill_2 FILLER_74_541 ();
 sg13g2_fill_2 FILLER_74_566 ();
 sg13g2_fill_2 FILLER_74_602 ();
 sg13g2_fill_1 FILLER_74_604 ();
 sg13g2_fill_2 FILLER_74_647 ();
 sg13g2_fill_1 FILLER_74_649 ();
 sg13g2_fill_1 FILLER_74_676 ();
 sg13g2_fill_2 FILLER_74_897 ();
 sg13g2_fill_2 FILLER_74_909 ();
 sg13g2_fill_1 FILLER_74_911 ();
 sg13g2_fill_1 FILLER_74_942 ();
 sg13g2_fill_1 FILLER_74_952 ();
 sg13g2_fill_2 FILLER_74_1029 ();
 sg13g2_fill_2 FILLER_74_1040 ();
 sg13g2_fill_1 FILLER_74_1042 ();
 sg13g2_fill_2 FILLER_74_1074 ();
 sg13g2_fill_1 FILLER_74_1076 ();
 sg13g2_fill_1 FILLER_74_1094 ();
 sg13g2_fill_1 FILLER_74_1115 ();
 sg13g2_fill_2 FILLER_74_1126 ();
 sg13g2_fill_1 FILLER_74_1128 ();
 sg13g2_fill_2 FILLER_74_1142 ();
 sg13g2_fill_2 FILLER_74_1154 ();
 sg13g2_fill_1 FILLER_74_1156 ();
 sg13g2_fill_1 FILLER_74_1214 ();
 sg13g2_fill_2 FILLER_74_1247 ();
 sg13g2_fill_2 FILLER_74_1254 ();
 sg13g2_fill_1 FILLER_74_1282 ();
 sg13g2_fill_1 FILLER_74_1292 ();
 sg13g2_fill_1 FILLER_74_1322 ();
 sg13g2_decap_4 FILLER_74_1340 ();
 sg13g2_fill_1 FILLER_74_1344 ();
 sg13g2_decap_4 FILLER_74_1354 ();
 sg13g2_fill_2 FILLER_74_1358 ();
 sg13g2_fill_2 FILLER_74_1377 ();
 sg13g2_fill_1 FILLER_74_1379 ();
 sg13g2_fill_1 FILLER_74_1394 ();
 sg13g2_fill_2 FILLER_74_1415 ();
 sg13g2_decap_8 FILLER_74_1431 ();
 sg13g2_fill_2 FILLER_74_1438 ();
 sg13g2_decap_4 FILLER_74_1448 ();
 sg13g2_fill_2 FILLER_74_1452 ();
 sg13g2_fill_1 FILLER_74_1468 ();
 sg13g2_fill_2 FILLER_74_1491 ();
 sg13g2_fill_2 FILLER_74_1506 ();
 sg13g2_fill_2 FILLER_74_1573 ();
 sg13g2_fill_2 FILLER_74_1584 ();
 sg13g2_fill_1 FILLER_74_1594 ();
 sg13g2_fill_2 FILLER_74_1631 ();
 sg13g2_fill_2 FILLER_74_1716 ();
 sg13g2_fill_2 FILLER_74_1741 ();
 sg13g2_fill_2 FILLER_74_1783 ();
 sg13g2_decap_4 FILLER_74_1809 ();
 sg13g2_decap_4 FILLER_74_1817 ();
 sg13g2_fill_2 FILLER_74_1821 ();
 sg13g2_fill_1 FILLER_74_1841 ();
 sg13g2_fill_2 FILLER_74_1868 ();
 sg13g2_fill_1 FILLER_74_1870 ();
 sg13g2_fill_1 FILLER_74_1887 ();
 sg13g2_fill_2 FILLER_74_1914 ();
 sg13g2_fill_1 FILLER_74_1916 ();
 sg13g2_fill_2 FILLER_74_1922 ();
 sg13g2_fill_1 FILLER_74_1924 ();
 sg13g2_fill_2 FILLER_74_1942 ();
 sg13g2_fill_2 FILLER_74_1957 ();
 sg13g2_fill_1 FILLER_74_1959 ();
 sg13g2_fill_2 FILLER_74_1968 ();
 sg13g2_fill_1 FILLER_74_1970 ();
 sg13g2_fill_1 FILLER_74_1981 ();
 sg13g2_fill_2 FILLER_74_2123 ();
 sg13g2_fill_1 FILLER_74_2125 ();
 sg13g2_fill_2 FILLER_74_2174 ();
 sg13g2_fill_1 FILLER_74_2186 ();
 sg13g2_fill_2 FILLER_74_2220 ();
 sg13g2_fill_1 FILLER_74_2222 ();
 sg13g2_fill_2 FILLER_74_2253 ();
 sg13g2_fill_1 FILLER_74_2255 ();
 sg13g2_fill_1 FILLER_74_2290 ();
 sg13g2_fill_1 FILLER_74_2374 ();
 sg13g2_fill_2 FILLER_74_2388 ();
 sg13g2_fill_1 FILLER_74_2390 ();
 sg13g2_fill_2 FILLER_74_2427 ();
 sg13g2_fill_2 FILLER_74_2465 ();
 sg13g2_fill_2 FILLER_74_2503 ();
 sg13g2_fill_1 FILLER_74_2505 ();
 sg13g2_decap_8 FILLER_74_2541 ();
 sg13g2_decap_8 FILLER_74_2548 ();
 sg13g2_decap_8 FILLER_74_2555 ();
 sg13g2_decap_8 FILLER_74_2562 ();
 sg13g2_decap_8 FILLER_74_2569 ();
 sg13g2_decap_8 FILLER_74_2576 ();
 sg13g2_decap_8 FILLER_74_2583 ();
 sg13g2_decap_8 FILLER_74_2590 ();
 sg13g2_decap_8 FILLER_74_2597 ();
 sg13g2_decap_8 FILLER_74_2604 ();
 sg13g2_decap_8 FILLER_74_2611 ();
 sg13g2_decap_8 FILLER_74_2618 ();
 sg13g2_decap_8 FILLER_74_2625 ();
 sg13g2_decap_8 FILLER_74_2632 ();
 sg13g2_decap_8 FILLER_74_2639 ();
 sg13g2_decap_8 FILLER_74_2646 ();
 sg13g2_decap_8 FILLER_74_2653 ();
 sg13g2_decap_8 FILLER_74_2660 ();
 sg13g2_decap_8 FILLER_74_2667 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_4 FILLER_75_84 ();
 sg13g2_fill_1 FILLER_75_147 ();
 sg13g2_fill_2 FILLER_75_153 ();
 sg13g2_fill_2 FILLER_75_177 ();
 sg13g2_fill_1 FILLER_75_179 ();
 sg13g2_fill_1 FILLER_75_243 ();
 sg13g2_fill_2 FILLER_75_279 ();
 sg13g2_fill_2 FILLER_75_346 ();
 sg13g2_fill_2 FILLER_75_383 ();
 sg13g2_fill_1 FILLER_75_407 ();
 sg13g2_fill_1 FILLER_75_474 ();
 sg13g2_fill_2 FILLER_75_501 ();
 sg13g2_fill_1 FILLER_75_570 ();
 sg13g2_fill_1 FILLER_75_623 ();
 sg13g2_fill_2 FILLER_75_654 ();
 sg13g2_fill_1 FILLER_75_656 ();
 sg13g2_fill_2 FILLER_75_773 ();
 sg13g2_fill_1 FILLER_75_849 ();
 sg13g2_fill_1 FILLER_75_911 ();
 sg13g2_fill_2 FILLER_75_1022 ();
 sg13g2_fill_1 FILLER_75_1032 ();
 sg13g2_fill_2 FILLER_75_1039 ();
 sg13g2_fill_1 FILLER_75_1041 ();
 sg13g2_fill_1 FILLER_75_1055 ();
 sg13g2_fill_1 FILLER_75_1101 ();
 sg13g2_fill_2 FILLER_75_1116 ();
 sg13g2_fill_2 FILLER_75_1187 ();
 sg13g2_fill_1 FILLER_75_1254 ();
 sg13g2_fill_1 FILLER_75_1316 ();
 sg13g2_fill_2 FILLER_75_1325 ();
 sg13g2_fill_2 FILLER_75_1339 ();
 sg13g2_fill_1 FILLER_75_1341 ();
 sg13g2_decap_4 FILLER_75_1358 ();
 sg13g2_fill_1 FILLER_75_1362 ();
 sg13g2_decap_4 FILLER_75_1376 ();
 sg13g2_fill_1 FILLER_75_1401 ();
 sg13g2_fill_2 FILLER_75_1418 ();
 sg13g2_fill_2 FILLER_75_1428 ();
 sg13g2_fill_2 FILLER_75_1443 ();
 sg13g2_decap_4 FILLER_75_1449 ();
 sg13g2_fill_1 FILLER_75_1498 ();
 sg13g2_fill_2 FILLER_75_1533 ();
 sg13g2_fill_2 FILLER_75_1542 ();
 sg13g2_fill_2 FILLER_75_1628 ();
 sg13g2_decap_4 FILLER_75_1660 ();
 sg13g2_fill_2 FILLER_75_1664 ();
 sg13g2_decap_8 FILLER_75_1670 ();
 sg13g2_fill_2 FILLER_75_1677 ();
 sg13g2_fill_1 FILLER_75_1679 ();
 sg13g2_decap_8 FILLER_75_1717 ();
 sg13g2_fill_1 FILLER_75_1724 ();
 sg13g2_decap_4 FILLER_75_1757 ();
 sg13g2_fill_1 FILLER_75_1761 ();
 sg13g2_fill_2 FILLER_75_1776 ();
 sg13g2_fill_2 FILLER_75_1783 ();
 sg13g2_decap_4 FILLER_75_1812 ();
 sg13g2_fill_1 FILLER_75_1816 ();
 sg13g2_decap_4 FILLER_75_1821 ();
 sg13g2_fill_2 FILLER_75_1825 ();
 sg13g2_fill_2 FILLER_75_1831 ();
 sg13g2_fill_2 FILLER_75_1863 ();
 sg13g2_fill_2 FILLER_75_1873 ();
 sg13g2_decap_4 FILLER_75_1883 ();
 sg13g2_fill_1 FILLER_75_1887 ();
 sg13g2_fill_1 FILLER_75_1905 ();
 sg13g2_decap_4 FILLER_75_1918 ();
 sg13g2_fill_1 FILLER_75_1922 ();
 sg13g2_fill_2 FILLER_75_1939 ();
 sg13g2_fill_1 FILLER_75_1941 ();
 sg13g2_fill_2 FILLER_75_1955 ();
 sg13g2_fill_2 FILLER_75_1965 ();
 sg13g2_fill_2 FILLER_75_1971 ();
 sg13g2_decap_8 FILLER_75_1982 ();
 sg13g2_fill_2 FILLER_75_1989 ();
 sg13g2_fill_1 FILLER_75_2008 ();
 sg13g2_fill_2 FILLER_75_2014 ();
 sg13g2_fill_2 FILLER_75_2042 ();
 sg13g2_fill_1 FILLER_75_2044 ();
 sg13g2_fill_2 FILLER_75_2055 ();
 sg13g2_fill_1 FILLER_75_2057 ();
 sg13g2_fill_1 FILLER_75_2062 ();
 sg13g2_fill_1 FILLER_75_2085 ();
 sg13g2_fill_2 FILLER_75_2095 ();
 sg13g2_fill_2 FILLER_75_2138 ();
 sg13g2_fill_1 FILLER_75_2140 ();
 sg13g2_fill_2 FILLER_75_2167 ();
 sg13g2_fill_1 FILLER_75_2208 ();
 sg13g2_fill_1 FILLER_75_2278 ();
 sg13g2_fill_1 FILLER_75_2314 ();
 sg13g2_fill_2 FILLER_75_2341 ();
 sg13g2_fill_2 FILLER_75_2384 ();
 sg13g2_fill_2 FILLER_75_2407 ();
 sg13g2_fill_2 FILLER_75_2469 ();
 sg13g2_decap_8 FILLER_75_2502 ();
 sg13g2_decap_8 FILLER_75_2509 ();
 sg13g2_fill_1 FILLER_75_2516 ();
 sg13g2_decap_8 FILLER_75_2521 ();
 sg13g2_decap_8 FILLER_75_2528 ();
 sg13g2_decap_8 FILLER_75_2535 ();
 sg13g2_decap_8 FILLER_75_2542 ();
 sg13g2_decap_8 FILLER_75_2549 ();
 sg13g2_decap_8 FILLER_75_2556 ();
 sg13g2_decap_8 FILLER_75_2563 ();
 sg13g2_decap_8 FILLER_75_2570 ();
 sg13g2_decap_8 FILLER_75_2577 ();
 sg13g2_decap_8 FILLER_75_2584 ();
 sg13g2_decap_8 FILLER_75_2591 ();
 sg13g2_decap_8 FILLER_75_2598 ();
 sg13g2_decap_8 FILLER_75_2605 ();
 sg13g2_decap_8 FILLER_75_2612 ();
 sg13g2_decap_8 FILLER_75_2619 ();
 sg13g2_decap_8 FILLER_75_2626 ();
 sg13g2_decap_8 FILLER_75_2633 ();
 sg13g2_decap_8 FILLER_75_2640 ();
 sg13g2_decap_8 FILLER_75_2647 ();
 sg13g2_decap_8 FILLER_75_2654 ();
 sg13g2_decap_8 FILLER_75_2661 ();
 sg13g2_decap_4 FILLER_75_2668 ();
 sg13g2_fill_2 FILLER_75_2672 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_fill_1 FILLER_76_91 ();
 sg13g2_fill_2 FILLER_76_129 ();
 sg13g2_fill_2 FILLER_76_236 ();
 sg13g2_fill_1 FILLER_76_238 ();
 sg13g2_fill_1 FILLER_76_312 ();
 sg13g2_fill_1 FILLER_76_364 ();
 sg13g2_fill_2 FILLER_76_406 ();
 sg13g2_fill_1 FILLER_76_439 ();
 sg13g2_fill_2 FILLER_76_576 ();
 sg13g2_fill_2 FILLER_76_614 ();
 sg13g2_fill_1 FILLER_76_616 ();
 sg13g2_fill_1 FILLER_76_638 ();
 sg13g2_fill_2 FILLER_76_649 ();
 sg13g2_fill_2 FILLER_76_693 ();
 sg13g2_fill_2 FILLER_76_714 ();
 sg13g2_fill_1 FILLER_76_716 ();
 sg13g2_fill_1 FILLER_76_752 ();
 sg13g2_fill_2 FILLER_76_762 ();
 sg13g2_fill_2 FILLER_76_773 ();
 sg13g2_fill_1 FILLER_76_775 ();
 sg13g2_fill_2 FILLER_76_782 ();
 sg13g2_fill_1 FILLER_76_784 ();
 sg13g2_fill_1 FILLER_76_830 ();
 sg13g2_fill_1 FILLER_76_850 ();
 sg13g2_fill_1 FILLER_76_905 ();
 sg13g2_fill_1 FILLER_76_932 ();
 sg13g2_fill_2 FILLER_76_1047 ();
 sg13g2_fill_1 FILLER_76_1049 ();
 sg13g2_fill_2 FILLER_76_1076 ();
 sg13g2_fill_1 FILLER_76_1078 ();
 sg13g2_fill_2 FILLER_76_1088 ();
 sg13g2_fill_2 FILLER_76_1095 ();
 sg13g2_fill_1 FILLER_76_1097 ();
 sg13g2_fill_2 FILLER_76_1108 ();
 sg13g2_fill_1 FILLER_76_1110 ();
 sg13g2_fill_1 FILLER_76_1138 ();
 sg13g2_fill_2 FILLER_76_1154 ();
 sg13g2_fill_1 FILLER_76_1156 ();
 sg13g2_fill_2 FILLER_76_1183 ();
 sg13g2_fill_1 FILLER_76_1185 ();
 sg13g2_fill_1 FILLER_76_1190 ();
 sg13g2_fill_2 FILLER_76_1226 ();
 sg13g2_fill_1 FILLER_76_1228 ();
 sg13g2_fill_2 FILLER_76_1318 ();
 sg13g2_decap_4 FILLER_76_1340 ();
 sg13g2_fill_2 FILLER_76_1344 ();
 sg13g2_fill_2 FILLER_76_1405 ();
 sg13g2_fill_1 FILLER_76_1407 ();
 sg13g2_fill_1 FILLER_76_1418 ();
 sg13g2_fill_1 FILLER_76_1424 ();
 sg13g2_fill_2 FILLER_76_1502 ();
 sg13g2_fill_1 FILLER_76_1538 ();
 sg13g2_decap_4 FILLER_76_1654 ();
 sg13g2_fill_1 FILLER_76_1658 ();
 sg13g2_fill_1 FILLER_76_1685 ();
 sg13g2_fill_1 FILLER_76_1695 ();
 sg13g2_fill_1 FILLER_76_1742 ();
 sg13g2_fill_2 FILLER_76_1765 ();
 sg13g2_fill_1 FILLER_76_1767 ();
 sg13g2_fill_2 FILLER_76_1776 ();
 sg13g2_fill_2 FILLER_76_1793 ();
 sg13g2_fill_1 FILLER_76_1795 ();
 sg13g2_fill_2 FILLER_76_1804 ();
 sg13g2_fill_1 FILLER_76_1832 ();
 sg13g2_decap_4 FILLER_76_1841 ();
 sg13g2_fill_2 FILLER_76_1875 ();
 sg13g2_fill_2 FILLER_76_1889 ();
 sg13g2_fill_2 FILLER_76_1899 ();
 sg13g2_fill_1 FILLER_76_1901 ();
 sg13g2_decap_8 FILLER_76_1928 ();
 sg13g2_fill_2 FILLER_76_1935 ();
 sg13g2_fill_2 FILLER_76_1947 ();
 sg13g2_fill_2 FILLER_76_1957 ();
 sg13g2_fill_1 FILLER_76_1959 ();
 sg13g2_fill_2 FILLER_76_1965 ();
 sg13g2_fill_1 FILLER_76_2028 ();
 sg13g2_fill_2 FILLER_76_2071 ();
 sg13g2_fill_1 FILLER_76_2078 ();
 sg13g2_fill_1 FILLER_76_2089 ();
 sg13g2_fill_2 FILLER_76_2120 ();
 sg13g2_fill_1 FILLER_76_2122 ();
 sg13g2_fill_2 FILLER_76_2217 ();
 sg13g2_fill_1 FILLER_76_2219 ();
 sg13g2_fill_2 FILLER_76_2289 ();
 sg13g2_fill_1 FILLER_76_2291 ();
 sg13g2_fill_2 FILLER_76_2351 ();
 sg13g2_fill_1 FILLER_76_2353 ();
 sg13g2_fill_2 FILLER_76_2403 ();
 sg13g2_fill_1 FILLER_76_2405 ();
 sg13g2_decap_8 FILLER_76_2493 ();
 sg13g2_decap_8 FILLER_76_2500 ();
 sg13g2_decap_8 FILLER_76_2507 ();
 sg13g2_decap_8 FILLER_76_2514 ();
 sg13g2_decap_8 FILLER_76_2521 ();
 sg13g2_decap_8 FILLER_76_2528 ();
 sg13g2_decap_8 FILLER_76_2535 ();
 sg13g2_decap_8 FILLER_76_2542 ();
 sg13g2_decap_8 FILLER_76_2549 ();
 sg13g2_decap_8 FILLER_76_2556 ();
 sg13g2_decap_8 FILLER_76_2563 ();
 sg13g2_decap_8 FILLER_76_2570 ();
 sg13g2_decap_8 FILLER_76_2577 ();
 sg13g2_decap_8 FILLER_76_2584 ();
 sg13g2_decap_8 FILLER_76_2591 ();
 sg13g2_decap_8 FILLER_76_2598 ();
 sg13g2_decap_8 FILLER_76_2605 ();
 sg13g2_decap_8 FILLER_76_2612 ();
 sg13g2_decap_8 FILLER_76_2619 ();
 sg13g2_decap_8 FILLER_76_2626 ();
 sg13g2_decap_8 FILLER_76_2633 ();
 sg13g2_decap_8 FILLER_76_2640 ();
 sg13g2_decap_8 FILLER_76_2647 ();
 sg13g2_decap_8 FILLER_76_2654 ();
 sg13g2_decap_8 FILLER_76_2661 ();
 sg13g2_decap_4 FILLER_76_2668 ();
 sg13g2_fill_2 FILLER_76_2672 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_4 FILLER_77_91 ();
 sg13g2_fill_2 FILLER_77_95 ();
 sg13g2_fill_1 FILLER_77_204 ();
 sg13g2_fill_2 FILLER_77_427 ();
 sg13g2_fill_1 FILLER_77_444 ();
 sg13g2_fill_1 FILLER_77_454 ();
 sg13g2_fill_1 FILLER_77_482 ();
 sg13g2_fill_2 FILLER_77_600 ();
 sg13g2_fill_1 FILLER_77_602 ();
 sg13g2_fill_2 FILLER_77_711 ();
 sg13g2_fill_1 FILLER_77_713 ();
 sg13g2_fill_2 FILLER_77_750 ();
 sg13g2_fill_1 FILLER_77_752 ();
 sg13g2_fill_1 FILLER_77_762 ();
 sg13g2_fill_2 FILLER_77_822 ();
 sg13g2_fill_1 FILLER_77_824 ();
 sg13g2_fill_2 FILLER_77_859 ();
 sg13g2_fill_1 FILLER_77_887 ();
 sg13g2_fill_2 FILLER_77_897 ();
 sg13g2_fill_1 FILLER_77_924 ();
 sg13g2_fill_2 FILLER_77_969 ();
 sg13g2_fill_1 FILLER_77_971 ();
 sg13g2_fill_2 FILLER_77_983 ();
 sg13g2_fill_1 FILLER_77_985 ();
 sg13g2_fill_1 FILLER_77_1010 ();
 sg13g2_fill_1 FILLER_77_1030 ();
 sg13g2_fill_1 FILLER_77_1074 ();
 sg13g2_fill_1 FILLER_77_1080 ();
 sg13g2_fill_2 FILLER_77_1113 ();
 sg13g2_fill_1 FILLER_77_1115 ();
 sg13g2_fill_2 FILLER_77_1125 ();
 sg13g2_fill_2 FILLER_77_1158 ();
 sg13g2_fill_1 FILLER_77_1160 ();
 sg13g2_fill_2 FILLER_77_1167 ();
 sg13g2_fill_1 FILLER_77_1169 ();
 sg13g2_fill_1 FILLER_77_1201 ();
 sg13g2_fill_1 FILLER_77_1233 ();
 sg13g2_fill_2 FILLER_77_1239 ();
 sg13g2_fill_1 FILLER_77_1241 ();
 sg13g2_decap_4 FILLER_77_1293 ();
 sg13g2_fill_2 FILLER_77_1297 ();
 sg13g2_decap_8 FILLER_77_1315 ();
 sg13g2_decap_4 FILLER_77_1322 ();
 sg13g2_fill_2 FILLER_77_1326 ();
 sg13g2_decap_8 FILLER_77_1341 ();
 sg13g2_fill_1 FILLER_77_1353 ();
 sg13g2_decap_4 FILLER_77_1365 ();
 sg13g2_fill_2 FILLER_77_1369 ();
 sg13g2_fill_2 FILLER_77_1393 ();
 sg13g2_fill_2 FILLER_77_1400 ();
 sg13g2_decap_4 FILLER_77_1406 ();
 sg13g2_fill_1 FILLER_77_1410 ();
 sg13g2_fill_2 FILLER_77_1418 ();
 sg13g2_decap_8 FILLER_77_1428 ();
 sg13g2_fill_1 FILLER_77_1446 ();
 sg13g2_fill_1 FILLER_77_1474 ();
 sg13g2_fill_2 FILLER_77_1508 ();
 sg13g2_fill_1 FILLER_77_1559 ();
 sg13g2_fill_2 FILLER_77_1578 ();
 sg13g2_fill_1 FILLER_77_1599 ();
 sg13g2_fill_1 FILLER_77_1614 ();
 sg13g2_decap_8 FILLER_77_1656 ();
 sg13g2_decap_8 FILLER_77_1663 ();
 sg13g2_decap_4 FILLER_77_1674 ();
 sg13g2_fill_1 FILLER_77_1678 ();
 sg13g2_fill_2 FILLER_77_1700 ();
 sg13g2_fill_2 FILLER_77_1715 ();
 sg13g2_decap_8 FILLER_77_1722 ();
 sg13g2_fill_1 FILLER_77_1729 ();
 sg13g2_fill_2 FILLER_77_1735 ();
 sg13g2_decap_4 FILLER_77_1742 ();
 sg13g2_fill_1 FILLER_77_1776 ();
 sg13g2_decap_4 FILLER_77_1788 ();
 sg13g2_fill_1 FILLER_77_1792 ();
 sg13g2_fill_1 FILLER_77_1812 ();
 sg13g2_fill_1 FILLER_77_1829 ();
 sg13g2_fill_2 FILLER_77_1834 ();
 sg13g2_fill_2 FILLER_77_1852 ();
 sg13g2_fill_1 FILLER_77_1854 ();
 sg13g2_decap_4 FILLER_77_1881 ();
 sg13g2_fill_1 FILLER_77_1885 ();
 sg13g2_decap_8 FILLER_77_1890 ();
 sg13g2_decap_4 FILLER_77_1902 ();
 sg13g2_fill_1 FILLER_77_1906 ();
 sg13g2_fill_2 FILLER_77_1942 ();
 sg13g2_fill_2 FILLER_77_1948 ();
 sg13g2_decap_4 FILLER_77_1983 ();
 sg13g2_fill_2 FILLER_77_1987 ();
 sg13g2_decap_4 FILLER_77_1993 ();
 sg13g2_fill_2 FILLER_77_1997 ();
 sg13g2_fill_1 FILLER_77_2013 ();
 sg13g2_decap_4 FILLER_77_2017 ();
 sg13g2_fill_2 FILLER_77_2026 ();
 sg13g2_fill_1 FILLER_77_2038 ();
 sg13g2_fill_1 FILLER_77_2144 ();
 sg13g2_fill_2 FILLER_77_2164 ();
 sg13g2_fill_1 FILLER_77_2166 ();
 sg13g2_fill_2 FILLER_77_2238 ();
 sg13g2_fill_1 FILLER_77_2240 ();
 sg13g2_fill_2 FILLER_77_2322 ();
 sg13g2_fill_2 FILLER_77_2342 ();
 sg13g2_fill_1 FILLER_77_2344 ();
 sg13g2_fill_2 FILLER_77_2355 ();
 sg13g2_fill_1 FILLER_77_2357 ();
 sg13g2_fill_2 FILLER_77_2377 ();
 sg13g2_fill_1 FILLER_77_2379 ();
 sg13g2_fill_2 FILLER_77_2399 ();
 sg13g2_fill_1 FILLER_77_2401 ();
 sg13g2_fill_1 FILLER_77_2425 ();
 sg13g2_decap_8 FILLER_77_2478 ();
 sg13g2_decap_8 FILLER_77_2485 ();
 sg13g2_decap_8 FILLER_77_2492 ();
 sg13g2_decap_8 FILLER_77_2499 ();
 sg13g2_decap_8 FILLER_77_2506 ();
 sg13g2_decap_8 FILLER_77_2513 ();
 sg13g2_decap_8 FILLER_77_2520 ();
 sg13g2_decap_8 FILLER_77_2527 ();
 sg13g2_decap_8 FILLER_77_2534 ();
 sg13g2_decap_8 FILLER_77_2541 ();
 sg13g2_decap_8 FILLER_77_2548 ();
 sg13g2_decap_8 FILLER_77_2555 ();
 sg13g2_decap_8 FILLER_77_2562 ();
 sg13g2_decap_8 FILLER_77_2569 ();
 sg13g2_decap_8 FILLER_77_2576 ();
 sg13g2_decap_8 FILLER_77_2583 ();
 sg13g2_decap_8 FILLER_77_2590 ();
 sg13g2_decap_8 FILLER_77_2597 ();
 sg13g2_decap_8 FILLER_77_2604 ();
 sg13g2_decap_8 FILLER_77_2611 ();
 sg13g2_decap_8 FILLER_77_2618 ();
 sg13g2_decap_8 FILLER_77_2625 ();
 sg13g2_decap_8 FILLER_77_2632 ();
 sg13g2_decap_8 FILLER_77_2639 ();
 sg13g2_decap_8 FILLER_77_2646 ();
 sg13g2_decap_8 FILLER_77_2653 ();
 sg13g2_decap_8 FILLER_77_2660 ();
 sg13g2_decap_8 FILLER_77_2667 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_fill_1 FILLER_78_98 ();
 sg13g2_fill_2 FILLER_78_103 ();
 sg13g2_fill_1 FILLER_78_196 ();
 sg13g2_fill_2 FILLER_78_246 ();
 sg13g2_fill_2 FILLER_78_274 ();
 sg13g2_fill_1 FILLER_78_294 ();
 sg13g2_fill_1 FILLER_78_334 ();
 sg13g2_fill_2 FILLER_78_349 ();
 sg13g2_fill_2 FILLER_78_406 ();
 sg13g2_fill_1 FILLER_78_422 ();
 sg13g2_fill_1 FILLER_78_431 ();
 sg13g2_fill_2 FILLER_78_441 ();
 sg13g2_fill_1 FILLER_78_452 ();
 sg13g2_fill_1 FILLER_78_613 ();
 sg13g2_fill_2 FILLER_78_623 ();
 sg13g2_fill_2 FILLER_78_631 ();
 sg13g2_fill_1 FILLER_78_649 ();
 sg13g2_fill_2 FILLER_78_744 ();
 sg13g2_fill_2 FILLER_78_777 ();
 sg13g2_fill_1 FILLER_78_831 ();
 sg13g2_fill_2 FILLER_78_856 ();
 sg13g2_fill_2 FILLER_78_884 ();
 sg13g2_fill_1 FILLER_78_886 ();
 sg13g2_fill_1 FILLER_78_911 ();
 sg13g2_fill_1 FILLER_78_928 ();
 sg13g2_fill_1 FILLER_78_937 ();
 sg13g2_fill_2 FILLER_78_964 ();
 sg13g2_fill_1 FILLER_78_966 ();
 sg13g2_fill_1 FILLER_78_1002 ();
 sg13g2_fill_1 FILLER_78_1100 ();
 sg13g2_fill_1 FILLER_78_1110 ();
 sg13g2_fill_2 FILLER_78_1137 ();
 sg13g2_fill_2 FILLER_78_1152 ();
 sg13g2_fill_1 FILLER_78_1154 ();
 sg13g2_fill_2 FILLER_78_1166 ();
 sg13g2_fill_1 FILLER_78_1168 ();
 sg13g2_fill_2 FILLER_78_1174 ();
 sg13g2_fill_2 FILLER_78_1328 ();
 sg13g2_decap_4 FILLER_78_1343 ();
 sg13g2_fill_1 FILLER_78_1365 ();
 sg13g2_fill_2 FILLER_78_1372 ();
 sg13g2_fill_1 FILLER_78_1374 ();
 sg13g2_fill_1 FILLER_78_1384 ();
 sg13g2_fill_2 FILLER_78_1393 ();
 sg13g2_fill_1 FILLER_78_1395 ();
 sg13g2_fill_2 FILLER_78_1411 ();
 sg13g2_decap_4 FILLER_78_1430 ();
 sg13g2_decap_8 FILLER_78_1442 ();
 sg13g2_fill_1 FILLER_78_1511 ();
 sg13g2_decap_8 FILLER_78_1650 ();
 sg13g2_decap_8 FILLER_78_1657 ();
 sg13g2_decap_8 FILLER_78_1664 ();
 sg13g2_decap_8 FILLER_78_1671 ();
 sg13g2_decap_4 FILLER_78_1678 ();
 sg13g2_fill_1 FILLER_78_1682 ();
 sg13g2_fill_2 FILLER_78_1693 ();
 sg13g2_fill_2 FILLER_78_1729 ();
 sg13g2_fill_2 FILLER_78_1747 ();
 sg13g2_fill_1 FILLER_78_1749 ();
 sg13g2_fill_2 FILLER_78_1767 ();
 sg13g2_fill_1 FILLER_78_1769 ();
 sg13g2_decap_4 FILLER_78_1782 ();
 sg13g2_fill_2 FILLER_78_1811 ();
 sg13g2_fill_1 FILLER_78_1813 ();
 sg13g2_fill_1 FILLER_78_1819 ();
 sg13g2_fill_2 FILLER_78_1828 ();
 sg13g2_fill_2 FILLER_78_1851 ();
 sg13g2_decap_8 FILLER_78_1858 ();
 sg13g2_fill_1 FILLER_78_1865 ();
 sg13g2_fill_1 FILLER_78_1870 ();
 sg13g2_fill_1 FILLER_78_1907 ();
 sg13g2_fill_2 FILLER_78_1925 ();
 sg13g2_fill_2 FILLER_78_1959 ();
 sg13g2_fill_1 FILLER_78_1981 ();
 sg13g2_decap_8 FILLER_78_1990 ();
 sg13g2_fill_2 FILLER_78_1997 ();
 sg13g2_fill_1 FILLER_78_1999 ();
 sg13g2_fill_2 FILLER_78_2025 ();
 sg13g2_fill_1 FILLER_78_2050 ();
 sg13g2_fill_2 FILLER_78_2070 ();
 sg13g2_fill_1 FILLER_78_2072 ();
 sg13g2_fill_2 FILLER_78_2091 ();
 sg13g2_fill_1 FILLER_78_2093 ();
 sg13g2_fill_1 FILLER_78_2103 ();
 sg13g2_fill_2 FILLER_78_2187 ();
 sg13g2_fill_2 FILLER_78_2213 ();
 sg13g2_fill_1 FILLER_78_2215 ();
 sg13g2_fill_2 FILLER_78_2314 ();
 sg13g2_fill_1 FILLER_78_2316 ();
 sg13g2_fill_1 FILLER_78_2343 ();
 sg13g2_fill_2 FILLER_78_2370 ();
 sg13g2_decap_8 FILLER_78_2474 ();
 sg13g2_decap_8 FILLER_78_2481 ();
 sg13g2_decap_8 FILLER_78_2488 ();
 sg13g2_decap_8 FILLER_78_2495 ();
 sg13g2_decap_8 FILLER_78_2502 ();
 sg13g2_decap_8 FILLER_78_2509 ();
 sg13g2_decap_8 FILLER_78_2516 ();
 sg13g2_decap_8 FILLER_78_2523 ();
 sg13g2_decap_8 FILLER_78_2530 ();
 sg13g2_decap_8 FILLER_78_2537 ();
 sg13g2_decap_8 FILLER_78_2544 ();
 sg13g2_decap_8 FILLER_78_2551 ();
 sg13g2_decap_8 FILLER_78_2558 ();
 sg13g2_decap_8 FILLER_78_2565 ();
 sg13g2_decap_8 FILLER_78_2572 ();
 sg13g2_decap_8 FILLER_78_2579 ();
 sg13g2_decap_8 FILLER_78_2586 ();
 sg13g2_decap_8 FILLER_78_2593 ();
 sg13g2_decap_8 FILLER_78_2600 ();
 sg13g2_decap_8 FILLER_78_2607 ();
 sg13g2_decap_8 FILLER_78_2614 ();
 sg13g2_decap_8 FILLER_78_2621 ();
 sg13g2_decap_8 FILLER_78_2628 ();
 sg13g2_decap_8 FILLER_78_2635 ();
 sg13g2_decap_8 FILLER_78_2642 ();
 sg13g2_decap_8 FILLER_78_2649 ();
 sg13g2_decap_8 FILLER_78_2656 ();
 sg13g2_decap_8 FILLER_78_2663 ();
 sg13g2_decap_4 FILLER_78_2670 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_4 FILLER_79_91 ();
 sg13g2_fill_2 FILLER_79_226 ();
 sg13g2_fill_2 FILLER_79_263 ();
 sg13g2_fill_1 FILLER_79_508 ();
 sg13g2_fill_2 FILLER_79_554 ();
 sg13g2_fill_1 FILLER_79_556 ();
 sg13g2_fill_2 FILLER_79_627 ();
 sg13g2_fill_1 FILLER_79_669 ();
 sg13g2_fill_2 FILLER_79_679 ();
 sg13g2_fill_1 FILLER_79_681 ();
 sg13g2_fill_2 FILLER_79_688 ();
 sg13g2_fill_2 FILLER_79_703 ();
 sg13g2_fill_1 FILLER_79_705 ();
 sg13g2_fill_2 FILLER_79_757 ();
 sg13g2_fill_1 FILLER_79_759 ();
 sg13g2_fill_2 FILLER_79_804 ();
 sg13g2_fill_2 FILLER_79_858 ();
 sg13g2_fill_1 FILLER_79_860 ();
 sg13g2_fill_2 FILLER_79_904 ();
 sg13g2_fill_2 FILLER_79_974 ();
 sg13g2_fill_1 FILLER_79_976 ();
 sg13g2_fill_1 FILLER_79_986 ();
 sg13g2_fill_2 FILLER_79_1022 ();
 sg13g2_fill_2 FILLER_79_1052 ();
 sg13g2_fill_1 FILLER_79_1054 ();
 sg13g2_fill_1 FILLER_79_1081 ();
 sg13g2_fill_1 FILLER_79_1209 ();
 sg13g2_fill_1 FILLER_79_1280 ();
 sg13g2_fill_2 FILLER_79_1289 ();
 sg13g2_fill_1 FILLER_79_1295 ();
 sg13g2_fill_1 FILLER_79_1304 ();
 sg13g2_fill_2 FILLER_79_1316 ();
 sg13g2_fill_2 FILLER_79_1352 ();
 sg13g2_fill_1 FILLER_79_1354 ();
 sg13g2_fill_1 FILLER_79_1388 ();
 sg13g2_decap_8 FILLER_79_1400 ();
 sg13g2_fill_2 FILLER_79_1407 ();
 sg13g2_fill_1 FILLER_79_1409 ();
 sg13g2_fill_1 FILLER_79_1471 ();
 sg13g2_fill_1 FILLER_79_1491 ();
 sg13g2_fill_2 FILLER_79_1509 ();
 sg13g2_fill_2 FILLER_79_1541 ();
 sg13g2_fill_2 FILLER_79_1595 ();
 sg13g2_fill_2 FILLER_79_1616 ();
 sg13g2_decap_8 FILLER_79_1644 ();
 sg13g2_decap_8 FILLER_79_1651 ();
 sg13g2_decap_8 FILLER_79_1658 ();
 sg13g2_decap_8 FILLER_79_1665 ();
 sg13g2_decap_8 FILLER_79_1672 ();
 sg13g2_fill_2 FILLER_79_1679 ();
 sg13g2_fill_1 FILLER_79_1681 ();
 sg13g2_decap_8 FILLER_79_1722 ();
 sg13g2_decap_4 FILLER_79_1729 ();
 sg13g2_fill_2 FILLER_79_1733 ();
 sg13g2_fill_2 FILLER_79_1739 ();
 sg13g2_fill_1 FILLER_79_1791 ();
 sg13g2_fill_2 FILLER_79_1811 ();
 sg13g2_decap_8 FILLER_79_1817 ();
 sg13g2_decap_4 FILLER_79_1824 ();
 sg13g2_fill_2 FILLER_79_1832 ();
 sg13g2_fill_1 FILLER_79_1851 ();
 sg13g2_fill_2 FILLER_79_1878 ();
 sg13g2_fill_1 FILLER_79_1880 ();
 sg13g2_fill_2 FILLER_79_1908 ();
 sg13g2_fill_1 FILLER_79_1910 ();
 sg13g2_fill_1 FILLER_79_1923 ();
 sg13g2_fill_1 FILLER_79_1932 ();
 sg13g2_decap_4 FILLER_79_1958 ();
 sg13g2_fill_2 FILLER_79_1962 ();
 sg13g2_decap_4 FILLER_79_1968 ();
 sg13g2_fill_1 FILLER_79_1972 ();
 sg13g2_fill_1 FILLER_79_1977 ();
 sg13g2_fill_2 FILLER_79_2002 ();
 sg13g2_fill_2 FILLER_79_2013 ();
 sg13g2_fill_2 FILLER_79_2089 ();
 sg13g2_fill_1 FILLER_79_2091 ();
 sg13g2_fill_1 FILLER_79_2131 ();
 sg13g2_fill_1 FILLER_79_2158 ();
 sg13g2_fill_2 FILLER_79_2199 ();
 sg13g2_fill_1 FILLER_79_2227 ();
 sg13g2_fill_2 FILLER_79_2277 ();
 sg13g2_fill_1 FILLER_79_2279 ();
 sg13g2_fill_2 FILLER_79_2294 ();
 sg13g2_fill_1 FILLER_79_2339 ();
 sg13g2_fill_1 FILLER_79_2349 ();
 sg13g2_fill_2 FILLER_79_2355 ();
 sg13g2_fill_1 FILLER_79_2357 ();
 sg13g2_fill_2 FILLER_79_2382 ();
 sg13g2_fill_2 FILLER_79_2397 ();
 sg13g2_fill_1 FILLER_79_2399 ();
 sg13g2_decap_8 FILLER_79_2466 ();
 sg13g2_decap_8 FILLER_79_2473 ();
 sg13g2_decap_8 FILLER_79_2480 ();
 sg13g2_decap_8 FILLER_79_2487 ();
 sg13g2_decap_8 FILLER_79_2494 ();
 sg13g2_decap_8 FILLER_79_2501 ();
 sg13g2_decap_8 FILLER_79_2508 ();
 sg13g2_decap_8 FILLER_79_2515 ();
 sg13g2_decap_8 FILLER_79_2522 ();
 sg13g2_decap_8 FILLER_79_2529 ();
 sg13g2_decap_8 FILLER_79_2536 ();
 sg13g2_decap_8 FILLER_79_2543 ();
 sg13g2_decap_8 FILLER_79_2550 ();
 sg13g2_decap_8 FILLER_79_2557 ();
 sg13g2_decap_8 FILLER_79_2564 ();
 sg13g2_decap_8 FILLER_79_2571 ();
 sg13g2_decap_8 FILLER_79_2578 ();
 sg13g2_decap_8 FILLER_79_2585 ();
 sg13g2_decap_8 FILLER_79_2592 ();
 sg13g2_decap_8 FILLER_79_2599 ();
 sg13g2_decap_8 FILLER_79_2606 ();
 sg13g2_decap_8 FILLER_79_2613 ();
 sg13g2_decap_8 FILLER_79_2620 ();
 sg13g2_decap_8 FILLER_79_2627 ();
 sg13g2_decap_8 FILLER_79_2634 ();
 sg13g2_decap_8 FILLER_79_2641 ();
 sg13g2_decap_8 FILLER_79_2648 ();
 sg13g2_decap_8 FILLER_79_2655 ();
 sg13g2_decap_8 FILLER_79_2662 ();
 sg13g2_decap_4 FILLER_79_2669 ();
 sg13g2_fill_1 FILLER_79_2673 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_8 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_75 ();
 sg13g2_fill_1 FILLER_80_79 ();
 sg13g2_fill_2 FILLER_80_333 ();
 sg13g2_fill_1 FILLER_80_428 ();
 sg13g2_fill_1 FILLER_80_455 ();
 sg13g2_fill_1 FILLER_80_465 ();
 sg13g2_fill_2 FILLER_80_536 ();
 sg13g2_fill_2 FILLER_80_567 ();
 sg13g2_fill_1 FILLER_80_569 ();
 sg13g2_fill_2 FILLER_80_589 ();
 sg13g2_fill_1 FILLER_80_591 ();
 sg13g2_fill_1 FILLER_80_601 ();
 sg13g2_fill_2 FILLER_80_650 ();
 sg13g2_fill_1 FILLER_80_652 ();
 sg13g2_fill_2 FILLER_80_662 ();
 sg13g2_fill_2 FILLER_80_793 ();
 sg13g2_fill_1 FILLER_80_795 ();
 sg13g2_fill_1 FILLER_80_861 ();
 sg13g2_fill_2 FILLER_80_966 ();
 sg13g2_fill_2 FILLER_80_1020 ();
 sg13g2_fill_1 FILLER_80_1060 ();
 sg13g2_fill_2 FILLER_80_1087 ();
 sg13g2_fill_2 FILLER_80_1185 ();
 sg13g2_fill_1 FILLER_80_1187 ();
 sg13g2_fill_1 FILLER_80_1238 ();
 sg13g2_fill_1 FILLER_80_1278 ();
 sg13g2_decap_8 FILLER_80_1334 ();
 sg13g2_decap_8 FILLER_80_1341 ();
 sg13g2_fill_1 FILLER_80_1348 ();
 sg13g2_decap_8 FILLER_80_1369 ();
 sg13g2_fill_2 FILLER_80_1376 ();
 sg13g2_fill_2 FILLER_80_1383 ();
 sg13g2_decap_8 FILLER_80_1395 ();
 sg13g2_decap_8 FILLER_80_1402 ();
 sg13g2_decap_8 FILLER_80_1409 ();
 sg13g2_decap_8 FILLER_80_1416 ();
 sg13g2_decap_8 FILLER_80_1423 ();
 sg13g2_decap_4 FILLER_80_1430 ();
 sg13g2_fill_1 FILLER_80_1434 ();
 sg13g2_fill_1 FILLER_80_1447 ();
 sg13g2_fill_2 FILLER_80_1475 ();
 sg13g2_fill_1 FILLER_80_1512 ();
 sg13g2_decap_8 FILLER_80_1549 ();
 sg13g2_fill_1 FILLER_80_1556 ();
 sg13g2_fill_1 FILLER_80_1586 ();
 sg13g2_fill_2 FILLER_80_1596 ();
 sg13g2_decap_8 FILLER_80_1633 ();
 sg13g2_decap_8 FILLER_80_1640 ();
 sg13g2_decap_8 FILLER_80_1647 ();
 sg13g2_decap_8 FILLER_80_1654 ();
 sg13g2_decap_8 FILLER_80_1661 ();
 sg13g2_decap_8 FILLER_80_1668 ();
 sg13g2_decap_8 FILLER_80_1675 ();
 sg13g2_decap_8 FILLER_80_1682 ();
 sg13g2_decap_8 FILLER_80_1689 ();
 sg13g2_fill_1 FILLER_80_1696 ();
 sg13g2_fill_2 FILLER_80_1714 ();
 sg13g2_fill_1 FILLER_80_1716 ();
 sg13g2_decap_8 FILLER_80_1726 ();
 sg13g2_decap_8 FILLER_80_1733 ();
 sg13g2_decap_8 FILLER_80_1740 ();
 sg13g2_fill_2 FILLER_80_1747 ();
 sg13g2_fill_1 FILLER_80_1749 ();
 sg13g2_decap_8 FILLER_80_1765 ();
 sg13g2_decap_4 FILLER_80_1772 ();
 sg13g2_decap_8 FILLER_80_1780 ();
 sg13g2_decap_8 FILLER_80_1787 ();
 sg13g2_decap_4 FILLER_80_1798 ();
 sg13g2_fill_1 FILLER_80_1802 ();
 sg13g2_decap_8 FILLER_80_1829 ();
 sg13g2_fill_1 FILLER_80_1836 ();
 sg13g2_fill_2 FILLER_80_1850 ();
 sg13g2_fill_2 FILLER_80_1861 ();
 sg13g2_fill_1 FILLER_80_1867 ();
 sg13g2_decap_4 FILLER_80_1876 ();
 sg13g2_fill_2 FILLER_80_1880 ();
 sg13g2_fill_1 FILLER_80_1887 ();
 sg13g2_fill_1 FILLER_80_1919 ();
 sg13g2_decap_4 FILLER_80_1932 ();
 sg13g2_fill_2 FILLER_80_1945 ();
 sg13g2_fill_1 FILLER_80_1947 ();
 sg13g2_decap_4 FILLER_80_1979 ();
 sg13g2_fill_1 FILLER_80_1983 ();
 sg13g2_fill_1 FILLER_80_2104 ();
 sg13g2_fill_2 FILLER_80_2208 ();
 sg13g2_fill_1 FILLER_80_2210 ();
 sg13g2_fill_2 FILLER_80_2287 ();
 sg13g2_fill_1 FILLER_80_2289 ();
 sg13g2_fill_2 FILLER_80_2343 ();
 sg13g2_fill_1 FILLER_80_2354 ();
 sg13g2_fill_2 FILLER_80_2360 ();
 sg13g2_fill_1 FILLER_80_2362 ();
 sg13g2_fill_2 FILLER_80_2402 ();
 sg13g2_decap_8 FILLER_80_2464 ();
 sg13g2_decap_8 FILLER_80_2471 ();
 sg13g2_decap_8 FILLER_80_2478 ();
 sg13g2_decap_8 FILLER_80_2485 ();
 sg13g2_decap_8 FILLER_80_2492 ();
 sg13g2_decap_8 FILLER_80_2499 ();
 sg13g2_decap_8 FILLER_80_2506 ();
 sg13g2_decap_8 FILLER_80_2513 ();
 sg13g2_decap_8 FILLER_80_2520 ();
 sg13g2_decap_8 FILLER_80_2527 ();
 sg13g2_decap_8 FILLER_80_2534 ();
 sg13g2_decap_8 FILLER_80_2541 ();
 sg13g2_decap_8 FILLER_80_2548 ();
 sg13g2_decap_8 FILLER_80_2555 ();
 sg13g2_decap_8 FILLER_80_2562 ();
 sg13g2_decap_8 FILLER_80_2569 ();
 sg13g2_decap_8 FILLER_80_2576 ();
 sg13g2_decap_8 FILLER_80_2583 ();
 sg13g2_decap_8 FILLER_80_2590 ();
 sg13g2_decap_8 FILLER_80_2597 ();
 sg13g2_decap_8 FILLER_80_2604 ();
 sg13g2_decap_8 FILLER_80_2611 ();
 sg13g2_decap_8 FILLER_80_2618 ();
 sg13g2_decap_8 FILLER_80_2625 ();
 sg13g2_decap_8 FILLER_80_2632 ();
 sg13g2_decap_8 FILLER_80_2639 ();
 sg13g2_decap_8 FILLER_80_2646 ();
 sg13g2_decap_8 FILLER_80_2653 ();
 sg13g2_decap_8 FILLER_80_2660 ();
 sg13g2_decap_8 FILLER_80_2667 ();
 assign uio_oe[0] = net2886;
 assign uio_oe[3] = net2887;
 assign uio_oe[6] = net2888;
 assign uio_oe[7] = net2889;
 assign uio_out[6] = net2890;
endmodule

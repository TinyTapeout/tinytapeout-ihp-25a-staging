module tt_um_tinysynth (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \ChiselTop.tinySynth.io_pwmOut ;
 wire \ChiselTop.tinySynth.midi._GEN_0[0] ;
 wire \ChiselTop.tinySynth.midi._GEN_0[1] ;
 wire \ChiselTop.tinySynth.midi._GEN_0[2] ;
 wire \ChiselTop.tinySynth.midi._GEN_0[4] ;
 wire \ChiselTop.tinySynth.midi._GEN_0[5] ;
 wire \ChiselTop.tinySynth.midi._GEN_0[6] ;
 wire \ChiselTop.tinySynth.midi.hdr_channel[3] ;
 wire \ChiselTop.tinySynth.midi.hdr_msgType[3] ;
 wire \ChiselTop.tinySynth.midi.io_midiOut_bits_hdr_channel[0] ;
 wire \ChiselTop.tinySynth.midi.io_midiOut_bits_hdr_channel[1] ;
 wire \ChiselTop.tinySynth.midi.io_midiOut_bits_hdr_channel[2] ;
 wire \ChiselTop.tinySynth.midi.io_midiOut_bits_hdr_channel[3] ;
 wire \ChiselTop.tinySynth.midi.io_midiOut_bits_note[0] ;
 wire \ChiselTop.tinySynth.midi.io_midiOut_bits_note[1] ;
 wire \ChiselTop.tinySynth.midi.io_midiOut_bits_note[2] ;
 wire \ChiselTop.tinySynth.midi.io_midiOut_bits_note[3] ;
 wire \ChiselTop.tinySynth.midi.io_midiOut_bits_note[4] ;
 wire \ChiselTop.tinySynth.midi.io_midiOut_bits_note[5] ;
 wire \ChiselTop.tinySynth.midi.io_midiOut_bits_note[6] ;
 wire \ChiselTop.tinySynth.midi.io_uartIn_valid ;
 wire \ChiselTop.tinySynth.midi.regState[0] ;
 wire \ChiselTop.tinySynth.midi.regState[1] ;
 wire \ChiselTop.tinySynth.midi.regState[2] ;
 wire \ChiselTop.tinySynth.midi.regState[3] ;
 wire \ChiselTop.tinySynth.osc.square._cnt_T_1[0] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[0] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[10] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[11] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[12] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[13] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[14] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[15] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[16] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[17] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[18] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[19] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[1] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[20] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[21] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[22] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[23] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[24] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[25] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[26] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[27] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[28] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[29] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[2] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[30] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[31] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[3] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[4] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[5] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[6] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[7] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[8] ;
 wire \ChiselTop.tinySynth.osc.square.cnt[9] ;
 wire \ChiselTop.tinySynth.pwm._counter_T_1[0] ;
 wire \ChiselTop.tinySynth.pwm.counter[0] ;
 wire \ChiselTop.tinySynth.pwm.counter[1] ;
 wire \ChiselTop.tinySynth.pwm.counter[2] ;
 wire \ChiselTop.tinySynth.pwm.counter[3] ;
 wire \ChiselTop.tinySynth.pwm.counter[4] ;
 wire \ChiselTop.tinySynth.pwm.counter[5] ;
 wire \ChiselTop.tinySynth.pwm.counter[6] ;
 wire \ChiselTop.tinySynth.pwm.counter[7] ;
 wire \ChiselTop.tinySynth.uart.rx.bitsReg[0] ;
 wire \ChiselTop.tinySynth.uart.rx.bitsReg[1] ;
 wire \ChiselTop.tinySynth.uart.rx.bitsReg[2] ;
 wire \ChiselTop.tinySynth.uart.rx.bitsReg[3] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[0] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[10] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[11] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[12] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[13] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[14] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[15] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[16] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[17] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[18] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[19] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[1] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[2] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[3] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[4] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[5] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[6] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[7] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[8] ;
 wire \ChiselTop.tinySynth.uart.rx.cntReg[9] ;
 wire \ChiselTop.tinySynth.uart.rx.falling_REG ;
 wire \ChiselTop.tinySynth.uart.rx.rxReg ;
 wire \ChiselTop.tinySynth.uart.rx.rxReg_REG ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire clknet_0_clk;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net1;
 wire net2;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;

 sg13g2_inv_1 _0713_ (.Y(_0111_),
    .A(net170));
 sg13g2_inv_1 _0714_ (.Y(_0112_),
    .A(net175));
 sg13g2_inv_1 _0715_ (.Y(_0113_),
    .A(net184));
 sg13g2_inv_1 _0716_ (.Y(_0114_),
    .A(net168));
 sg13g2_inv_2 _0717_ (.Y(_0115_),
    .A(net129));
 sg13g2_inv_1 _0718_ (.Y(_0116_),
    .A(net296));
 sg13g2_inv_1 _0719_ (.Y(_0117_),
    .A(net210));
 sg13g2_inv_1 _0720_ (.Y(_0118_),
    .A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[3] ));
 sg13g2_inv_1 _0721_ (.Y(_0119_),
    .A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[2] ));
 sg13g2_inv_1 _0722_ (.Y(_0120_),
    .A(net260));
 sg13g2_inv_1 _0723_ (.Y(_0121_),
    .A(net290));
 sg13g2_inv_1 _0724_ (.Y(_0122_),
    .A(net230));
 sg13g2_inv_1 _0725_ (.Y(_0123_),
    .A(net232));
 sg13g2_inv_1 _0726_ (.Y(_0124_),
    .A(net245));
 sg13g2_inv_1 _0727_ (.Y(_0125_),
    .A(net270));
 sg13g2_inv_1 _0728_ (.Y(_0126_),
    .A(net213));
 sg13g2_inv_1 _0729_ (.Y(_0127_),
    .A(net152));
 sg13g2_inv_1 _0730_ (.Y(_0128_),
    .A(net202));
 sg13g2_inv_1 _0731_ (.Y(_0129_),
    .A(_0012_));
 sg13g2_inv_1 _0732_ (.Y(_0130_),
    .A(_0011_));
 sg13g2_inv_1 _0733_ (.Y(_0131_),
    .A(_0010_));
 sg13g2_inv_1 _0734_ (.Y(_0132_),
    .A(_0009_));
 sg13g2_inv_1 _0735_ (.Y(_0133_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[19] ));
 sg13g2_inv_1 _0736_ (.Y(_0134_),
    .A(net305));
 sg13g2_inv_1 _0737_ (.Y(_0135_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[21] ));
 sg13g2_inv_1 _0738_ (.Y(_0136_),
    .A(net309));
 sg13g2_inv_1 _0739_ (.Y(_0137_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[31] ));
 sg13g2_inv_1 _0740_ (.Y(_0138_),
    .A(net134));
 sg13g2_inv_1 _0741_ (.Y(_0139_),
    .A(net132));
 sg13g2_inv_1 _0742_ (.Y(_0140_),
    .A(\ChiselTop.tinySynth.uart.rx.falling_REG ));
 sg13g2_inv_1 _0743_ (.Y(_0141_),
    .A(net162));
 sg13g2_inv_1 _0744_ (.Y(_0142_),
    .A(net157));
 sg13g2_inv_1 _0745_ (.Y(_0143_),
    .A(net179));
 sg13g2_inv_1 _0746_ (.Y(_0144_),
    .A(net302));
 sg13g2_inv_1 _0747_ (.Y(_0145_),
    .A(net310));
 sg13g2_inv_1 _0748_ (.Y(_0146_),
    .A(net153));
 sg13g2_nor2_1 _0749_ (.A(\ChiselTop.tinySynth.midi.regState[1] ),
    .B(\ChiselTop.tinySynth.midi.regState[2] ),
    .Y(_0147_));
 sg13g2_nand2_1 _0750_ (.Y(_0148_),
    .A(_0024_),
    .B(_0147_));
 sg13g2_nand2_1 _0751_ (.Y(_0149_),
    .A(net245),
    .B(_0148_));
 sg13g2_nand2_1 _0752_ (.Y(_0150_),
    .A(net137),
    .B(_0149_));
 sg13g2_nand3_1 _0753_ (.B(net286),
    .C(_0149_),
    .A(net136),
    .Y(_0151_));
 sg13g2_nor2_1 _0754_ (.A(net260),
    .B(net230),
    .Y(_0152_));
 sg13g2_nand2_1 _0755_ (.Y(_0153_),
    .A(\ChiselTop.tinySynth.midi.hdr_msgType[3] ),
    .B(_0152_));
 sg13g2_nand3_1 _0756_ (.B(\ChiselTop.tinySynth.midi.regState[0] ),
    .C(_0153_),
    .A(net202),
    .Y(_0154_));
 sg13g2_nand4_1 _0757_ (.B(_0139_),
    .C(_0151_),
    .A(net139),
    .Y(_0001_),
    .D(_0154_));
 sg13g2_nand3_1 _0758_ (.B(net136),
    .C(net234),
    .A(_0124_),
    .Y(_0155_));
 sg13g2_nand3_1 _0759_ (.B(net136),
    .C(_0148_),
    .A(net245),
    .Y(_0156_));
 sg13g2_nand3_1 _0760_ (.B(net286),
    .C(_0152_),
    .A(net202),
    .Y(_0157_));
 sg13g2_o21ai_1 _0761_ (.B1(_0155_),
    .Y(_0003_),
    .A1(_0156_),
    .A2(_0157_));
 sg13g2_nand3_1 _0762_ (.B(net136),
    .C(net208),
    .A(_0124_),
    .Y(_0158_));
 sg13g2_a21oi_1 _0763_ (.A1(_0128_),
    .A2(\ChiselTop.tinySynth.midi.regState[0] ),
    .Y(_0159_),
    .B1(net234));
 sg13g2_o21ai_1 _0764_ (.B1(_0158_),
    .Y(_0002_),
    .A1(_0156_),
    .A2(net235));
 sg13g2_nor2_1 _0765_ (.A(\ChiselTop.tinySynth.osc.square.cnt[22] ),
    .B(\ChiselTop.tinySynth.osc.square.cnt[23] ),
    .Y(_0160_));
 sg13g2_nor3_2 _0766_ (.A(\ChiselTop.tinySynth.midi.io_midiOut_bits_hdr_channel[1] ),
    .B(\ChiselTop.tinySynth.midi.io_midiOut_bits_hdr_channel[0] ),
    .C(\ChiselTop.tinySynth.midi.regState[0] ),
    .Y(_0161_));
 sg13g2_nor4_2 _0767_ (.A(\ChiselTop.tinySynth.midi.io_midiOut_bits_hdr_channel[3] ),
    .B(\ChiselTop.tinySynth.midi.io_midiOut_bits_hdr_channel[2] ),
    .C(\ChiselTop.tinySynth.midi.regState[1] ),
    .Y(_0162_),
    .D(\ChiselTop.tinySynth.midi.regState[2] ));
 sg13g2_and3_1 _0768_ (.X(_0163_),
    .A(net131),
    .B(net128),
    .C(_0162_));
 sg13g2_nand3_1 _0769_ (.B(net128),
    .C(_0162_),
    .A(net131),
    .Y(_0164_));
 sg13g2_nand4_1 _0770_ (.B(net131),
    .C(_0161_),
    .A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[4] ),
    .Y(_0165_),
    .D(net127));
 sg13g2_nor3_2 _0771_ (.A(_0115_),
    .B(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[5] ),
    .C(_0165_),
    .Y(_0166_));
 sg13g2_nor3_1 _0772_ (.A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[2] ),
    .B(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[1] ),
    .C(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[0] ),
    .Y(_0167_));
 sg13g2_or4_1 _0773_ (.A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[3] ),
    .B(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[2] ),
    .C(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[1] ),
    .D(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[0] ),
    .X(_0168_));
 sg13g2_and4_1 _0774_ (.A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[3] ),
    .B(net131),
    .C(net128),
    .D(net127),
    .X(_0169_));
 sg13g2_nand4_1 _0775_ (.B(net132),
    .C(net128),
    .A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[3] ),
    .Y(_0170_),
    .D(net127));
 sg13g2_nand4_1 _0776_ (.B(net128),
    .C(net127),
    .A(net131),
    .Y(_0171_),
    .D(_0168_));
 sg13g2_nand4_1 _0777_ (.B(net131),
    .C(_0161_),
    .A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[5] ),
    .Y(_0172_),
    .D(net127));
 sg13g2_and2_1 _0778_ (.A(_0165_),
    .B(_0172_),
    .X(_0173_));
 sg13g2_nand4_1 _0779_ (.B(net131),
    .C(net128),
    .A(net129),
    .Y(_0174_),
    .D(net127));
 sg13g2_nor4_1 _0780_ (.A(_0115_),
    .B(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[5] ),
    .C(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[4] ),
    .D(net123),
    .Y(_0175_));
 sg13g2_nor2_1 _0781_ (.A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[2] ),
    .B(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[1] ),
    .Y(_0176_));
 sg13g2_nor2_1 _0782_ (.A(_0170_),
    .B(_0176_),
    .Y(_0177_));
 sg13g2_nand2b_1 _0783_ (.Y(_0178_),
    .B(_0169_),
    .A_N(_0176_));
 sg13g2_nor2_1 _0784_ (.A(_0117_),
    .B(_0172_),
    .Y(_0179_));
 sg13g2_nor3_1 _0785_ (.A(net129),
    .B(_0116_),
    .C(_0165_),
    .Y(_0180_));
 sg13g2_a221oi_1 _0786_ (.B2(_0180_),
    .C1(_0175_),
    .B1(_0177_),
    .A1(_0166_),
    .Y(_0181_),
    .A2(_0171_));
 sg13g2_nor3_2 _0787_ (.A(net129),
    .B(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[4] ),
    .C(_0172_),
    .Y(_0182_));
 sg13g2_nor3_1 _0788_ (.A(_0119_),
    .B(_0121_),
    .C(_0170_),
    .Y(_0183_));
 sg13g2_a22oi_1 _0789_ (.Y(_0184_),
    .B1(_0182_),
    .B2(_0183_),
    .A2(_0180_),
    .A1(_0178_));
 sg13g2_nand2_1 _0790_ (.Y(_0185_),
    .A(net121),
    .B(_0184_));
 sg13g2_a21o_1 _0791_ (.A2(_0176_),
    .A1(_0118_),
    .B1(net123),
    .X(_0186_));
 sg13g2_nand3_1 _0792_ (.B(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[2] ),
    .C(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[1] ),
    .A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[3] ),
    .Y(_0187_));
 sg13g2_nand3b_1 _0793_ (.B(_0187_),
    .C(_0182_),
    .Y(_0188_),
    .A_N(_0186_));
 sg13g2_inv_1 _0794_ (.Y(_0189_),
    .A(_0188_));
 sg13g2_nor3_1 _0795_ (.A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[6] ),
    .B(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[5] ),
    .C(_0165_),
    .Y(_0190_));
 sg13g2_a21o_1 _0796_ (.A2(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[1] ),
    .A1(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[2] ),
    .B1(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[3] ),
    .X(_0191_));
 sg13g2_and4_1 _0797_ (.A(net131),
    .B(net128),
    .C(net127),
    .D(_0191_),
    .X(_0192_));
 sg13g2_nand4_1 _0798_ (.B(net128),
    .C(net127),
    .A(net132),
    .Y(_0193_),
    .D(_0191_));
 sg13g2_nor4_2 _0799_ (.A(net129),
    .B(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[5] ),
    .C(_0165_),
    .Y(_0194_),
    .D(_0193_));
 sg13g2_a21oi_1 _0800_ (.A1(_0182_),
    .A2(_0186_),
    .Y(_0195_),
    .B1(_0194_));
 sg13g2_nor4_2 _0801_ (.A(net129),
    .B(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[5] ),
    .C(_0165_),
    .Y(_0196_),
    .D(_0192_));
 sg13g2_nor3_1 _0802_ (.A(net129),
    .B(_0170_),
    .C(_0176_),
    .Y(_0197_));
 sg13g2_a21oi_1 _0803_ (.A1(_0173_),
    .A2(_0197_),
    .Y(_0198_),
    .B1(_0196_));
 sg13g2_a221oi_1 _0804_ (.B2(_0173_),
    .C1(_0190_),
    .B1(_0197_),
    .A1(_0182_),
    .Y(_0199_),
    .A2(_0186_));
 sg13g2_and4_1 _0805_ (.A(net120),
    .B(_0184_),
    .C(net119),
    .D(_0199_),
    .X(_0200_));
 sg13g2_nand4_1 _0806_ (.B(_0184_),
    .C(net119),
    .A(net120),
    .Y(_0201_),
    .D(_0199_));
 sg13g2_nor3_2 _0807_ (.A(_0115_),
    .B(_0116_),
    .C(_0165_),
    .Y(_0202_));
 sg13g2_nor3_2 _0808_ (.A(_0115_),
    .B(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[4] ),
    .C(_0172_),
    .Y(_0203_));
 sg13g2_nor2_2 _0809_ (.A(_0167_),
    .B(_0170_),
    .Y(_0204_));
 sg13g2_nand2b_1 _0810_ (.Y(_0205_),
    .B(_0169_),
    .A_N(_0167_));
 sg13g2_a21oi_2 _0811_ (.B1(_0202_),
    .Y(_0206_),
    .A2(_0204_),
    .A1(_0203_));
 sg13g2_a21oi_1 _0812_ (.A1(_0121_),
    .A2(_0123_),
    .Y(_0207_),
    .B1(_0119_));
 sg13g2_o21ai_1 _0813_ (.B1(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[2] ),
    .Y(_0208_),
    .A1(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[1] ),
    .A2(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[0] ));
 sg13g2_nor2_2 _0814_ (.A(_0170_),
    .B(_0208_),
    .Y(_0209_));
 sg13g2_a22oi_1 _0815_ (.Y(_0210_),
    .B1(_0209_),
    .B2(_0166_),
    .A2(_0205_),
    .A1(_0203_));
 sg13g2_a221oi_1 _0816_ (.B2(_0166_),
    .C1(_0203_),
    .B1(_0209_),
    .A1(net129),
    .Y(_0211_),
    .A2(_0179_));
 sg13g2_a21oi_2 _0817_ (.B1(_0171_),
    .Y(_0212_),
    .A2(_0207_),
    .A1(_0169_));
 sg13g2_nand2_2 _0818_ (.Y(_0213_),
    .A(_0166_),
    .B(_0212_));
 sg13g2_a221oi_1 _0819_ (.B2(_0166_),
    .C1(_0194_),
    .B1(_0212_),
    .A1(_0182_),
    .Y(_0214_),
    .A2(_0186_));
 sg13g2_and3_1 _0820_ (.X(_0215_),
    .A(net120),
    .B(_0211_),
    .C(_0214_));
 sg13g2_and4_1 _0821_ (.A(net125),
    .B(net120),
    .C(_0211_),
    .D(_0214_),
    .X(_0216_));
 sg13g2_nand4_1 _0822_ (.B(net120),
    .C(_0211_),
    .A(net126),
    .Y(_0217_),
    .D(_0214_));
 sg13g2_a221oi_1 _0823_ (.B2(_0166_),
    .C1(_0202_),
    .B1(_0212_),
    .A1(_0203_),
    .Y(_0218_),
    .A2(_0204_));
 sg13g2_and2_1 _0824_ (.A(net119),
    .B(_0210_),
    .X(_0219_));
 sg13g2_nand4_1 _0825_ (.B(net119),
    .C(_0210_),
    .A(net126),
    .Y(_0220_),
    .D(_0218_));
 sg13g2_a21oi_2 _0826_ (.B1(_0201_),
    .Y(_0221_),
    .A2(_0220_),
    .A1(_0217_));
 sg13g2_nand3_1 _0827_ (.B(_0210_),
    .C(_0218_),
    .A(net119),
    .Y(_0222_));
 sg13g2_and3_1 _0828_ (.X(_0223_),
    .A(_0165_),
    .B(_0172_),
    .C(_0174_));
 sg13g2_a21oi_2 _0829_ (.B1(_0196_),
    .Y(_0224_),
    .A2(_0223_),
    .A1(_0177_));
 sg13g2_nand2_1 _0830_ (.Y(_0225_),
    .A(_0195_),
    .B(_0224_));
 sg13g2_xnor2_1 _0831_ (.Y(_0226_),
    .A(_0134_),
    .B(_0221_));
 sg13g2_nor4_2 _0832_ (.A(\ChiselTop.tinySynth.osc.square.cnt[21] ),
    .B(\ChiselTop.tinySynth.osc.square.cnt[22] ),
    .C(\ChiselTop.tinySynth.osc.square.cnt[23] ),
    .Y(_0227_),
    .D(_0226_));
 sg13g2_nand2_1 _0833_ (.Y(_0228_),
    .A(_0118_),
    .B(_0208_));
 sg13g2_nand2_1 _0834_ (.Y(_0229_),
    .A(net126),
    .B(_0228_));
 sg13g2_nand3_1 _0835_ (.B(_0202_),
    .C(_0228_),
    .A(net126),
    .Y(_0230_));
 sg13g2_a21oi_2 _0836_ (.B1(net123),
    .Y(_0231_),
    .A2(_0228_),
    .A1(_0202_));
 sg13g2_a22oi_1 _0837_ (.Y(_0232_),
    .B1(_0229_),
    .B2(_0202_),
    .A2(_0204_),
    .A1(_0203_));
 sg13g2_a221oi_1 _0838_ (.B2(_0202_),
    .C1(_0203_),
    .B1(_0229_),
    .A1(_0166_),
    .Y(_0233_),
    .A2(_0209_));
 sg13g2_nand2_1 _0839_ (.Y(_0234_),
    .A(_0210_),
    .B(_0232_));
 sg13g2_nand2_1 _0840_ (.Y(_0235_),
    .A(_0231_),
    .B(_0233_));
 sg13g2_nand4_1 _0841_ (.B(_0184_),
    .C(_0195_),
    .A(net121),
    .Y(_0236_),
    .D(_0213_));
 sg13g2_nor3_2 _0842_ (.A(_0189_),
    .B(_0235_),
    .C(_0236_),
    .Y(_0237_));
 sg13g2_nand2b_1 _0843_ (.Y(_0238_),
    .B(\ChiselTop.tinySynth.osc.square.cnt[19] ),
    .A_N(_0237_));
 sg13g2_and4_1 _0844_ (.A(net121),
    .B(_0184_),
    .C(_0198_),
    .D(_0213_),
    .X(_0239_));
 sg13g2_nand4_1 _0845_ (.B(_0184_),
    .C(_0198_),
    .A(net121),
    .Y(_0240_),
    .D(_0213_));
 sg13g2_nor2_1 _0846_ (.A(_0235_),
    .B(_0240_),
    .Y(_0241_));
 sg13g2_nand2b_1 _0847_ (.Y(_0242_),
    .B(_0239_),
    .A_N(_0235_));
 sg13g2_nor2_1 _0848_ (.A(_0234_),
    .B(_0240_),
    .Y(_0243_));
 sg13g2_nand2_1 _0849_ (.Y(_0244_),
    .A(net125),
    .B(_0243_));
 sg13g2_xnor2_1 _0850_ (.Y(_0245_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[18] ),
    .B(_0199_));
 sg13g2_and2_1 _0851_ (.A(_0133_),
    .B(_0237_),
    .X(_0246_));
 sg13g2_a221oi_1 _0852_ (.B2(_0132_),
    .C1(_0245_),
    .B1(_0242_),
    .A1(_0133_),
    .Y(_0247_),
    .A2(_0237_));
 sg13g2_a22oi_1 _0853_ (.Y(_0248_),
    .B1(_0220_),
    .B2(_0130_),
    .A2(_0217_),
    .A1(_0131_));
 sg13g2_nand3_1 _0854_ (.B(_0247_),
    .C(_0248_),
    .A(_0238_),
    .Y(_0249_));
 sg13g2_nand3_1 _0855_ (.B(_0206_),
    .C(_0224_),
    .A(net121),
    .Y(_0250_));
 sg13g2_or2_1 _0856_ (.X(_0251_),
    .B(_0250_),
    .A(net124));
 sg13g2_and4_2 _0857_ (.A(net120),
    .B(net119),
    .C(_0199_),
    .D(_0213_),
    .X(_0252_));
 sg13g2_nand4_1 _0858_ (.B(net119),
    .C(_0199_),
    .A(net120),
    .Y(_0253_),
    .D(_0213_));
 sg13g2_xnor2_1 _0859_ (.Y(_0254_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[14] ),
    .B(_0252_));
 sg13g2_a21oi_1 _0860_ (.A1(\ChiselTop.tinySynth.osc.square.cnt[13] ),
    .A2(_0251_),
    .Y(_0255_),
    .B1(_0254_));
 sg13g2_nand2_1 _0861_ (.Y(_0256_),
    .A(_0214_),
    .B(_0231_));
 sg13g2_or2_1 _0862_ (.X(_0257_),
    .B(_0256_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[12] ));
 sg13g2_o21ai_1 _0863_ (.B1(_0257_),
    .Y(_0258_),
    .A1(\ChiselTop.tinySynth.osc.square.cnt[13] ),
    .A2(_0251_));
 sg13g2_nand2_1 _0864_ (.Y(_0259_),
    .A(_0184_),
    .B(_0232_));
 sg13g2_nor2_1 _0865_ (.A(net124),
    .B(_0259_),
    .Y(_0260_));
 sg13g2_xor2_1 _0866_ (.B(_0260_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[10] ),
    .X(_0261_));
 sg13g2_and2_1 _0867_ (.A(net120),
    .B(_0231_),
    .X(_0262_));
 sg13g2_a21oi_1 _0868_ (.A1(_0200_),
    .A2(_0211_),
    .Y(_0263_),
    .B1(\ChiselTop.tinySynth.osc.square.cnt[8] ));
 sg13g2_xnor2_1 _0869_ (.Y(_0264_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[9] ),
    .B(_0262_));
 sg13g2_a22oi_1 _0870_ (.Y(_0265_),
    .B1(_0263_),
    .B2(_0264_),
    .A2(_0262_),
    .A1(_0016_));
 sg13g2_and3_1 _0871_ (.X(_0266_),
    .A(_0014_),
    .B(net125),
    .C(_0219_));
 sg13g2_a21oi_1 _0872_ (.A1(_0015_),
    .A2(_0260_),
    .Y(_0267_),
    .B1(_0266_));
 sg13g2_o21ai_1 _0873_ (.B1(_0267_),
    .Y(_0268_),
    .A1(_0261_),
    .A2(_0265_));
 sg13g2_a21oi_1 _0874_ (.A1(net125),
    .A2(_0219_),
    .Y(_0269_),
    .B1(_0014_));
 sg13g2_a21oi_1 _0875_ (.A1(\ChiselTop.tinySynth.osc.square.cnt[12] ),
    .A2(_0256_),
    .Y(_0270_),
    .B1(_0269_));
 sg13g2_a21o_1 _0876_ (.A2(_0270_),
    .A1(_0268_),
    .B1(_0258_),
    .X(_0271_));
 sg13g2_nor3_1 _0877_ (.A(_0130_),
    .B(net124),
    .C(_0222_),
    .Y(_0272_));
 sg13g2_a221oi_1 _0878_ (.B2(_0271_),
    .C1(_0272_),
    .B1(_0255_),
    .A1(_0012_),
    .Y(_0273_),
    .A2(_0253_));
 sg13g2_nor2_1 _0879_ (.A(_0249_),
    .B(_0273_),
    .Y(_0274_));
 sg13g2_and3_1 _0880_ (.X(_0275_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[8] ),
    .B(_0200_),
    .C(_0211_));
 sg13g2_or4_1 _0881_ (.A(_0258_),
    .B(_0261_),
    .C(_0263_),
    .D(_0275_),
    .X(_0276_));
 sg13g2_nor2_1 _0882_ (.A(_0266_),
    .B(_0272_),
    .Y(_0277_));
 sg13g2_nand4_1 _0883_ (.B(_0264_),
    .C(_0270_),
    .A(_0255_),
    .Y(_0278_),
    .D(_0277_));
 sg13g2_nand2_1 _0884_ (.Y(_0279_),
    .A(_0010_),
    .B(_0216_));
 sg13g2_o21ai_1 _0885_ (.B1(_0279_),
    .Y(_0280_),
    .A1(_0132_),
    .A2(_0242_));
 sg13g2_nor4_1 _0886_ (.A(_0249_),
    .B(_0276_),
    .C(_0278_),
    .D(_0280_),
    .Y(_0281_));
 sg13g2_nand3b_1 _0887_ (.B(_0188_),
    .C(_0206_),
    .Y(_0282_),
    .A_N(_0236_));
 sg13g2_and2_1 _0888_ (.A(_0018_),
    .B(_0282_),
    .X(_0283_));
 sg13g2_nor2_1 _0889_ (.A(_0164_),
    .B(_0225_),
    .Y(_0284_));
 sg13g2_nand2_2 _0890_ (.Y(_0285_),
    .A(net125),
    .B(_0206_));
 sg13g2_o21ai_1 _0891_ (.B1(_0230_),
    .Y(_0286_),
    .A1(_0225_),
    .A2(_0285_));
 sg13g2_xor2_1 _0892_ (.B(_0286_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[6] ),
    .X(_0287_));
 sg13g2_nor2_1 _0893_ (.A(_0018_),
    .B(_0282_),
    .Y(_0288_));
 sg13g2_or3_1 _0894_ (.A(_0283_),
    .B(_0287_),
    .C(_0288_),
    .X(_0289_));
 sg13g2_nand3_1 _0895_ (.B(net119),
    .C(_0224_),
    .A(net126),
    .Y(_0290_));
 sg13g2_nor3_2 _0896_ (.A(_0185_),
    .B(_0234_),
    .C(_0290_),
    .Y(_0291_));
 sg13g2_nand2_1 _0897_ (.Y(_0292_),
    .A(_0023_),
    .B(_0250_));
 sg13g2_nand3b_1 _0898_ (.B(_0292_),
    .C(\ChiselTop.tinySynth.osc.square.cnt[0] ),
    .Y(_0293_),
    .A_N(_0291_));
 sg13g2_nor2_1 _0899_ (.A(\ChiselTop.tinySynth.osc.square.cnt[4] ),
    .B(_0215_),
    .Y(_0294_));
 sg13g2_a21oi_1 _0900_ (.A1(_0233_),
    .A2(_0239_),
    .Y(_0295_),
    .B1(net130));
 sg13g2_or2_1 _0901_ (.X(_0296_),
    .B(_0295_),
    .A(_0294_));
 sg13g2_and3_1 _0902_ (.X(_0297_),
    .A(net130),
    .B(_0233_),
    .C(_0239_));
 sg13g2_nand2_1 _0903_ (.Y(_0298_),
    .A(net130),
    .B(_0243_));
 sg13g2_and2_1 _0904_ (.A(\ChiselTop.tinySynth.osc.square.cnt[4] ),
    .B(_0215_),
    .X(_0299_));
 sg13g2_nor4_2 _0905_ (.A(_0294_),
    .B(_0295_),
    .C(_0297_),
    .Y(_0300_),
    .D(_0299_));
 sg13g2_nand2_1 _0906_ (.Y(_0301_),
    .A(net125),
    .B(_0252_));
 sg13g2_nor3_1 _0907_ (.A(\ChiselTop.tinySynth.osc.square.cnt[2] ),
    .B(net124),
    .C(_0253_),
    .Y(_0302_));
 sg13g2_a21oi_1 _0908_ (.A1(net125),
    .A2(_0252_),
    .Y(_0303_),
    .B1(_0145_));
 sg13g2_nor2_1 _0909_ (.A(_0023_),
    .B(_0250_),
    .Y(_0304_));
 sg13g2_nand2_1 _0910_ (.Y(_0305_),
    .A(_0021_),
    .B(_0222_));
 sg13g2_xnor2_1 _0911_ (.Y(_0306_),
    .A(_0021_),
    .B(_0222_));
 sg13g2_nor4_1 _0912_ (.A(_0302_),
    .B(_0303_),
    .C(_0304_),
    .D(_0306_),
    .Y(_0307_));
 sg13g2_nand2_1 _0913_ (.Y(_0308_),
    .A(_0300_),
    .B(_0307_));
 sg13g2_nand3_1 _0914_ (.B(_0300_),
    .C(_0307_),
    .A(_0293_),
    .Y(_0309_));
 sg13g2_o21ai_1 _0915_ (.B1(_0022_),
    .Y(_0310_),
    .A1(_0021_),
    .A2(_0222_));
 sg13g2_o21ai_1 _0916_ (.B1(_0305_),
    .Y(_0311_),
    .A1(_0301_),
    .A2(_0310_));
 sg13g2_a22oi_1 _0917_ (.Y(_0312_),
    .B1(_0300_),
    .B2(_0311_),
    .A2(_0298_),
    .A1(_0296_));
 sg13g2_a21oi_1 _0918_ (.A1(_0309_),
    .A2(_0312_),
    .Y(_0313_),
    .B1(_0289_));
 sg13g2_a22oi_1 _0919_ (.Y(_0314_),
    .B1(_0286_),
    .B2(_0019_),
    .A2(_0282_),
    .A1(_0018_));
 sg13g2_nor2_1 _0920_ (.A(_0288_),
    .B(_0314_),
    .Y(_0315_));
 sg13g2_o21ai_1 _0921_ (.B1(_0281_),
    .Y(_0316_),
    .A1(_0313_),
    .A2(_0315_));
 sg13g2_nand3_1 _0922_ (.B(_0247_),
    .C(_0280_),
    .A(_0238_),
    .Y(_0317_));
 sg13g2_nor2b_1 _0923_ (.A(_0199_),
    .B_N(_0008_),
    .Y(_0318_));
 sg13g2_o21ai_1 _0924_ (.B1(_0238_),
    .Y(_0319_),
    .A1(_0246_),
    .A2(_0318_));
 sg13g2_nand3_1 _0925_ (.B(_0317_),
    .C(_0319_),
    .A(_0316_),
    .Y(_0320_));
 sg13g2_o21ai_1 _0926_ (.B1(_0227_),
    .Y(_0321_),
    .A1(_0274_),
    .A2(_0320_));
 sg13g2_nand4_1 _0927_ (.B(_0135_),
    .C(_0160_),
    .A(_0007_),
    .Y(_0322_),
    .D(_0221_));
 sg13g2_nor4_1 _0928_ (.A(\ChiselTop.tinySynth.osc.square.cnt[28] ),
    .B(\ChiselTop.tinySynth.osc.square.cnt[29] ),
    .C(\ChiselTop.tinySynth.osc.square.cnt[30] ),
    .D(\ChiselTop.tinySynth.osc.square.cnt[31] ),
    .Y(_0323_));
 sg13g2_nor4_1 _0929_ (.A(\ChiselTop.tinySynth.osc.square.cnt[24] ),
    .B(\ChiselTop.tinySynth.osc.square.cnt[25] ),
    .C(\ChiselTop.tinySynth.osc.square.cnt[26] ),
    .D(\ChiselTop.tinySynth.osc.square.cnt[27] ),
    .Y(_0324_));
 sg13g2_and2_1 _0930_ (.A(_0323_),
    .B(_0324_),
    .X(_0325_));
 sg13g2_nor4_1 _0931_ (.A(\ChiselTop.tinySynth.pwm.counter[5] ),
    .B(\ChiselTop.tinySynth.pwm.counter[4] ),
    .C(\ChiselTop.tinySynth.pwm.counter[3] ),
    .D(\ChiselTop.tinySynth.pwm.counter[2] ),
    .Y(_0326_));
 sg13g2_nor4_1 _0932_ (.A(\ChiselTop.tinySynth.pwm.counter[0] ),
    .B(\ChiselTop.tinySynth.pwm.counter[6] ),
    .C(\ChiselTop.tinySynth.pwm.counter[7] ),
    .D(\ChiselTop.tinySynth.pwm.counter[1] ),
    .Y(_0327_));
 sg13g2_nand3_1 _0933_ (.B(_0326_),
    .C(_0327_),
    .A(_0325_),
    .Y(_0328_));
 sg13g2_xnor2_1 _0934_ (.Y(_0329_),
    .A(_0146_),
    .B(_0291_));
 sg13g2_nand3_1 _0935_ (.B(_0292_),
    .C(_0329_),
    .A(_0227_),
    .Y(_0330_));
 sg13g2_nor3_1 _0936_ (.A(_0289_),
    .B(_0308_),
    .C(_0330_),
    .Y(_0331_));
 sg13g2_a221oi_1 _0937_ (.B2(_0281_),
    .C1(_0328_),
    .B1(_0331_),
    .A1(_0321_),
    .Y(\ChiselTop.tinySynth.io_pwmOut ),
    .A2(_0322_));
 sg13g2_and3_1 _0938_ (.X(_0000_),
    .A(\ChiselTop.tinySynth.midi.io_uartIn_valid ),
    .B(net136),
    .C(net208));
 sg13g2_and2_1 _0939_ (.A(net140),
    .B(net154),
    .X(_0025_));
 sg13g2_nor2_1 _0940_ (.A(_0236_),
    .B(_0285_),
    .Y(_0332_));
 sg13g2_nand2_1 _0941_ (.Y(_0333_),
    .A(_0188_),
    .B(_0332_));
 sg13g2_xor2_1 _0942_ (.B(_0333_),
    .A(_0017_),
    .X(_0334_));
 sg13g2_xor2_1 _0943_ (.B(_0244_),
    .A(_0019_),
    .X(_0335_));
 sg13g2_o21ai_1 _0944_ (.B1(_0008_),
    .Y(_0336_),
    .A1(_0164_),
    .A2(_0241_));
 sg13g2_and3_1 _0945_ (.X(_0337_),
    .A(net126),
    .B(_0200_),
    .C(_0211_));
 sg13g2_xnor2_1 _0946_ (.Y(_0338_),
    .A(_0016_),
    .B(_0337_));
 sg13g2_nand4_1 _0947_ (.B(_0335_),
    .C(_0336_),
    .A(_0334_),
    .Y(_0339_),
    .D(_0338_));
 sg13g2_or3_1 _0948_ (.A(_0250_),
    .B(_0291_),
    .C(_0332_),
    .X(_0340_));
 sg13g2_o21ai_1 _0949_ (.B1(_0250_),
    .Y(_0341_),
    .A1(_0291_),
    .A2(_0332_));
 sg13g2_and2_1 _0950_ (.A(_0340_),
    .B(_0341_),
    .X(_0342_));
 sg13g2_xor2_1 _0951_ (.B(_0342_),
    .A(_0022_),
    .X(_0343_));
 sg13g2_a21oi_1 _0952_ (.A1(_0252_),
    .A2(_0340_),
    .Y(_0344_),
    .B1(_0164_));
 sg13g2_xnor2_1 _0953_ (.Y(_0345_),
    .A(_0021_),
    .B(_0344_));
 sg13g2_o21ai_1 _0954_ (.B1(_0007_),
    .Y(_0346_),
    .A1(net123),
    .A2(_0237_));
 sg13g2_xor2_1 _0955_ (.B(_0291_),
    .A(_0023_),
    .X(_0347_));
 sg13g2_o21ai_1 _0956_ (.B1(\ChiselTop.tinySynth.osc.square.cnt[0] ),
    .Y(_0348_),
    .A1(_0236_),
    .A2(_0285_));
 sg13g2_nand2b_1 _0957_ (.Y(_0349_),
    .B(_0332_),
    .A_N(\ChiselTop.tinySynth.osc.square.cnt[0] ));
 sg13g2_mux2_1 _0958_ (.A0(_0348_),
    .A1(_0349_),
    .S(_0347_),
    .X(_0350_));
 sg13g2_nor3_1 _0959_ (.A(_0007_),
    .B(net123),
    .C(_0237_),
    .Y(_0351_));
 sg13g2_nor2_1 _0960_ (.A(_0350_),
    .B(_0351_),
    .Y(_0352_));
 sg13g2_nor2_1 _0961_ (.A(net124),
    .B(_0221_),
    .Y(_0353_));
 sg13g2_xnor2_1 _0962_ (.Y(_0354_),
    .A(_0135_),
    .B(_0353_));
 sg13g2_a21oi_1 _0963_ (.A1(_0214_),
    .A2(_0231_),
    .Y(_0355_),
    .B1(net123));
 sg13g2_xor2_1 _0964_ (.B(_0355_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[13] ),
    .X(_0356_));
 sg13g2_xnor2_1 _0965_ (.Y(_0357_),
    .A(_0130_),
    .B(net125));
 sg13g2_a22oi_1 _0966_ (.Y(_0358_),
    .B1(_0252_),
    .B2(_0357_),
    .A2(_0220_),
    .A1(_0020_));
 sg13g2_nand2_1 _0967_ (.Y(_0359_),
    .A(_0356_),
    .B(_0358_));
 sg13g2_xor2_1 _0968_ (.B(_0259_),
    .A(_0014_),
    .X(_0360_));
 sg13g2_xnor2_1 _0969_ (.Y(_0361_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[19] ),
    .B(_0284_));
 sg13g2_nor2_1 _0970_ (.A(_0252_),
    .B(_0357_),
    .Y(_0362_));
 sg13g2_or2_1 _0971_ (.X(_0363_),
    .B(_0219_),
    .A(_0013_));
 sg13g2_a21oi_1 _0972_ (.A1(_0160_),
    .A2(_0325_),
    .Y(_0364_),
    .B1(net124));
 sg13g2_nand4_1 _0973_ (.B(net199),
    .C(net237),
    .A(\ChiselTop.tinySynth.osc.square.cnt[24] ),
    .Y(_0365_),
    .D(net225));
 sg13g2_nand2_1 _0974_ (.Y(_0366_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[22] ),
    .B(net282));
 sg13g2_nor3_1 _0975_ (.A(_0137_),
    .B(_0365_),
    .C(_0366_),
    .Y(_0367_));
 sg13g2_nand4_1 _0976_ (.B(\ChiselTop.tinySynth.osc.square.cnt[29] ),
    .C(\ChiselTop.tinySynth.osc.square.cnt[30] ),
    .A(\ChiselTop.tinySynth.osc.square.cnt[28] ),
    .Y(_0368_),
    .D(_0367_));
 sg13g2_a221oi_1 _0977_ (.B2(net124),
    .C1(_0364_),
    .B1(_0368_),
    .A1(_0013_),
    .Y(_0369_),
    .A2(_0219_));
 sg13g2_nand3b_1 _0978_ (.B(_0363_),
    .C(_0369_),
    .Y(_0370_),
    .A_N(_0362_));
 sg13g2_nor4_1 _0979_ (.A(_0359_),
    .B(_0360_),
    .C(_0361_),
    .D(_0370_),
    .Y(_0371_));
 sg13g2_o21ai_1 _0980_ (.B1(_0231_),
    .Y(_0372_),
    .A1(_0225_),
    .A2(_0285_));
 sg13g2_xnor2_1 _0981_ (.Y(_0373_),
    .A(_0018_),
    .B(_0372_));
 sg13g2_nor2_1 _0982_ (.A(_0009_),
    .B(_0215_),
    .Y(_0374_));
 sg13g2_nand2_1 _0983_ (.Y(_0375_),
    .A(_0009_),
    .B(_0215_));
 sg13g2_o21ai_1 _0984_ (.B1(_0375_),
    .Y(_0376_),
    .A1(_0020_),
    .A2(_0220_));
 sg13g2_nor3_1 _0985_ (.A(_0373_),
    .B(_0374_),
    .C(_0376_),
    .Y(_0377_));
 sg13g2_nor3_1 _0986_ (.A(_0008_),
    .B(net123),
    .C(_0241_),
    .Y(_0378_));
 sg13g2_nand2_1 _0987_ (.Y(_0379_),
    .A(net130),
    .B(_0216_));
 sg13g2_or2_1 _0988_ (.X(_0380_),
    .B(_0222_),
    .A(_0131_));
 sg13g2_or2_1 _0989_ (.X(_0381_),
    .B(_0250_),
    .A(_0129_));
 sg13g2_a22oi_1 _0990_ (.Y(_0382_),
    .B1(_0250_),
    .B2(_0129_),
    .A2(_0222_),
    .A1(_0131_));
 sg13g2_nand4_1 _0991_ (.B(_0380_),
    .C(_0381_),
    .A(_0379_),
    .Y(_0383_),
    .D(_0382_));
 sg13g2_nor2_1 _0992_ (.A(net130),
    .B(_0216_),
    .Y(_0384_));
 sg13g2_nor2_1 _0993_ (.A(net123),
    .B(_0262_),
    .Y(_0385_));
 sg13g2_xor2_1 _0994_ (.B(_0385_),
    .A(_0015_),
    .X(_0386_));
 sg13g2_nor4_1 _0995_ (.A(_0378_),
    .B(_0383_),
    .C(_0384_),
    .D(_0386_),
    .Y(_0387_));
 sg13g2_and4_1 _0996_ (.A(_0354_),
    .B(_0371_),
    .C(_0377_),
    .D(_0387_),
    .X(_0388_));
 sg13g2_nand4_1 _0997_ (.B(_0346_),
    .C(_0352_),
    .A(_0345_),
    .Y(_0389_),
    .D(_0388_));
 sg13g2_nor3_1 _0998_ (.A(_0339_),
    .B(_0343_),
    .C(_0389_),
    .Y(_0390_));
 sg13g2_nand2b_1 _0999_ (.Y(_0391_),
    .B(net140),
    .A_N(_0390_));
 sg13g2_nor2_1 _1000_ (.A(_0146_),
    .B(net109),
    .Y(_0026_));
 sg13g2_nand2_1 _1001_ (.Y(_0392_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[0] ),
    .B(net217));
 sg13g2_xnor2_1 _1002_ (.Y(_0393_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[0] ),
    .B(net217));
 sg13g2_nor2_1 _1003_ (.A(net110),
    .B(net218),
    .Y(_0027_));
 sg13g2_xnor2_1 _1004_ (.Y(_0394_),
    .A(_0145_),
    .B(_0392_));
 sg13g2_nor2_1 _1005_ (.A(net110),
    .B(net311),
    .Y(_0028_));
 sg13g2_nor2_1 _1006_ (.A(_0022_),
    .B(_0392_),
    .Y(_0395_));
 sg13g2_xnor2_1 _1007_ (.Y(_0396_),
    .A(net211),
    .B(_0395_));
 sg13g2_nor2_1 _1008_ (.A(net110),
    .B(net212),
    .Y(_0029_));
 sg13g2_and4_2 _1009_ (.A(\ChiselTop.tinySynth.osc.square.cnt[2] ),
    .B(\ChiselTop.tinySynth.osc.square.cnt[0] ),
    .C(net217),
    .D(net211),
    .X(_0397_));
 sg13g2_and2_1 _1010_ (.A(net280),
    .B(_0397_),
    .X(_0398_));
 sg13g2_nor2_1 _1011_ (.A(net280),
    .B(_0397_),
    .Y(_0399_));
 sg13g2_nor3_1 _1012_ (.A(net110),
    .B(_0398_),
    .C(net281),
    .Y(_0030_));
 sg13g2_nor2b_1 _1013_ (.A(_0020_),
    .B_N(_0397_),
    .Y(_0400_));
 sg13g2_xnor2_1 _1014_ (.Y(_0401_),
    .A(net203),
    .B(_0400_));
 sg13g2_nor2_1 _1015_ (.A(net110),
    .B(net204),
    .Y(_0031_));
 sg13g2_and4_1 _1016_ (.A(net189),
    .B(net130),
    .C(\ChiselTop.tinySynth.osc.square.cnt[4] ),
    .D(_0397_),
    .X(_0402_));
 sg13g2_a21oi_1 _1017_ (.A1(net130),
    .A2(_0398_),
    .Y(_0403_),
    .B1(net189));
 sg13g2_nor3_1 _1018_ (.A(net110),
    .B(_0402_),
    .C(net190),
    .Y(_0032_));
 sg13g2_nand3b_1 _1019_ (.B(net130),
    .C(_0398_),
    .Y(_0404_),
    .A_N(_0019_));
 sg13g2_xor2_1 _1020_ (.B(_0404_),
    .A(net257),
    .X(_0405_));
 sg13g2_nor2_1 _1021_ (.A(net110),
    .B(net258),
    .Y(_0033_));
 sg13g2_and2_1 _1022_ (.A(net257),
    .B(_0402_),
    .X(_0406_));
 sg13g2_xnor2_1 _1023_ (.Y(_0407_),
    .A(net297),
    .B(_0406_));
 sg13g2_nor2_1 _1024_ (.A(_0391_),
    .B(_0407_),
    .Y(_0034_));
 sg13g2_nor2b_1 _1025_ (.A(net255),
    .B_N(_0406_),
    .Y(_0408_));
 sg13g2_xnor2_1 _1026_ (.Y(_0409_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[9] ),
    .B(_0408_));
 sg13g2_nor2_1 _1027_ (.A(net110),
    .B(net256),
    .Y(_0035_));
 sg13g2_and4_2 _1028_ (.A(\ChiselTop.tinySynth.osc.square.cnt[9] ),
    .B(\ChiselTop.tinySynth.osc.square.cnt[8] ),
    .C(net257),
    .D(_0402_),
    .X(_0410_));
 sg13g2_and2_1 _1029_ (.A(net265),
    .B(_0410_),
    .X(_0411_));
 sg13g2_nor2_1 _1030_ (.A(net265),
    .B(_0410_),
    .Y(_0412_));
 sg13g2_nor3_1 _1031_ (.A(net108),
    .B(_0411_),
    .C(net266),
    .Y(_0036_));
 sg13g2_nand2b_1 _1032_ (.Y(_0413_),
    .B(_0410_),
    .A_N(_0015_));
 sg13g2_xor2_1 _1033_ (.B(_0413_),
    .A(net288),
    .X(_0414_));
 sg13g2_nor2_1 _1034_ (.A(net108),
    .B(net289),
    .Y(_0037_));
 sg13g2_nand2_1 _1035_ (.Y(_0415_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[11] ),
    .B(_0411_));
 sg13g2_and4_1 _1036_ (.A(net181),
    .B(\ChiselTop.tinySynth.osc.square.cnt[10] ),
    .C(\ChiselTop.tinySynth.osc.square.cnt[11] ),
    .D(_0410_),
    .X(_0416_));
 sg13g2_a21oi_1 _1037_ (.A1(\ChiselTop.tinySynth.osc.square.cnt[11] ),
    .A2(_0411_),
    .Y(_0417_),
    .B1(net181));
 sg13g2_nor3_1 _1038_ (.A(net108),
    .B(_0416_),
    .C(net182),
    .Y(_0038_));
 sg13g2_nor2_1 _1039_ (.A(net219),
    .B(_0415_),
    .Y(_0418_));
 sg13g2_xnor2_1 _1040_ (.Y(_0419_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[13] ),
    .B(net220));
 sg13g2_nor2_1 _1041_ (.A(net108),
    .B(net221),
    .Y(_0039_));
 sg13g2_and2_1 _1042_ (.A(\ChiselTop.tinySynth.osc.square.cnt[13] ),
    .B(_0416_),
    .X(_0420_));
 sg13g2_xnor2_1 _1043_ (.Y(_0421_),
    .A(net294),
    .B(_0420_));
 sg13g2_nor2_1 _1044_ (.A(net108),
    .B(_0421_),
    .Y(_0040_));
 sg13g2_nand2_1 _1045_ (.Y(_0422_),
    .A(_0129_),
    .B(_0420_));
 sg13g2_xor2_1 _1046_ (.B(_0422_),
    .A(net261),
    .X(_0423_));
 sg13g2_nor2_1 _1047_ (.A(net108),
    .B(net262),
    .Y(_0041_));
 sg13g2_and4_1 _1048_ (.A(\ChiselTop.tinySynth.osc.square.cnt[14] ),
    .B(\ChiselTop.tinySynth.osc.square.cnt[15] ),
    .C(net205),
    .D(_0420_),
    .X(_0424_));
 sg13g2_and3_1 _1049_ (.X(_0425_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[14] ),
    .B(\ChiselTop.tinySynth.osc.square.cnt[15] ),
    .C(_0420_));
 sg13g2_nor2_1 _1050_ (.A(net205),
    .B(_0425_),
    .Y(_0426_));
 sg13g2_nor3_1 _1051_ (.A(net108),
    .B(_0424_),
    .C(net206),
    .Y(_0042_));
 sg13g2_and2_1 _1052_ (.A(_0131_),
    .B(_0425_),
    .X(_0427_));
 sg13g2_xnor2_1 _1053_ (.Y(_0428_),
    .A(net253),
    .B(_0427_));
 sg13g2_nor2_1 _1054_ (.A(net109),
    .B(net254),
    .Y(_0043_));
 sg13g2_nand3_1 _1055_ (.B(net253),
    .C(_0425_),
    .A(net205),
    .Y(_0429_));
 sg13g2_xnor2_1 _1056_ (.Y(_0430_),
    .A(net308),
    .B(_0429_));
 sg13g2_nor2b_1 _1057_ (.A(net109),
    .B_N(_0430_),
    .Y(_0044_));
 sg13g2_nor2_1 _1058_ (.A(net300),
    .B(_0429_),
    .Y(_0431_));
 sg13g2_xnor2_1 _1059_ (.Y(_0432_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[19] ),
    .B(_0431_));
 sg13g2_nor2_1 _1060_ (.A(net108),
    .B(net301),
    .Y(_0045_));
 sg13g2_nand4_1 _1061_ (.B(\ChiselTop.tinySynth.osc.square.cnt[18] ),
    .C(\ChiselTop.tinySynth.osc.square.cnt[19] ),
    .A(net253),
    .Y(_0433_),
    .D(_0424_));
 sg13g2_xnor2_1 _1062_ (.Y(_0434_),
    .A(_0134_),
    .B(_0433_));
 sg13g2_nor2_1 _1063_ (.A(net106),
    .B(net306),
    .Y(_0046_));
 sg13g2_nor2_1 _1064_ (.A(_0007_),
    .B(_0433_),
    .Y(_0435_));
 sg13g2_xnor2_1 _1065_ (.Y(_0436_),
    .A(net276),
    .B(_0435_));
 sg13g2_nor2_1 _1066_ (.A(net107),
    .B(net277),
    .Y(_0047_));
 sg13g2_or3_2 _1067_ (.A(_0134_),
    .B(_0135_),
    .C(_0433_),
    .X(_0437_));
 sg13g2_nor2_1 _1068_ (.A(_0136_),
    .B(_0437_),
    .Y(_0438_));
 sg13g2_and2_1 _1069_ (.A(_0136_),
    .B(_0437_),
    .X(_0439_));
 sg13g2_nor3_1 _1070_ (.A(net107),
    .B(_0438_),
    .C(_0439_),
    .Y(_0048_));
 sg13g2_nor2_1 _1071_ (.A(net282),
    .B(_0438_),
    .Y(_0440_));
 sg13g2_nor2_2 _1072_ (.A(_0366_),
    .B(_0437_),
    .Y(_0441_));
 sg13g2_nor3_1 _1073_ (.A(net107),
    .B(net283),
    .C(_0441_),
    .Y(_0049_));
 sg13g2_xnor2_1 _1074_ (.Y(_0442_),
    .A(net291),
    .B(_0441_));
 sg13g2_nor2_1 _1075_ (.A(net107),
    .B(net292),
    .Y(_0050_));
 sg13g2_a21oi_1 _1076_ (.A1(\ChiselTop.tinySynth.osc.square.cnt[24] ),
    .A2(_0441_),
    .Y(_0443_),
    .B1(net199));
 sg13g2_and3_1 _1077_ (.X(_0444_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[24] ),
    .B(net199),
    .C(_0441_));
 sg13g2_nor3_1 _1078_ (.A(net106),
    .B(net200),
    .C(_0444_),
    .Y(_0051_));
 sg13g2_nor2_1 _1079_ (.A(net237),
    .B(_0444_),
    .Y(_0445_));
 sg13g2_and2_1 _1080_ (.A(net237),
    .B(_0444_),
    .X(_0446_));
 sg13g2_nor3_1 _1081_ (.A(net106),
    .B(net238),
    .C(_0446_),
    .Y(_0052_));
 sg13g2_nor2_1 _1082_ (.A(net225),
    .B(_0446_),
    .Y(_0447_));
 sg13g2_nor3_1 _1083_ (.A(_0365_),
    .B(_0366_),
    .C(_0437_),
    .Y(_0448_));
 sg13g2_nor3_1 _1084_ (.A(net106),
    .B(net226),
    .C(_0448_),
    .Y(_0053_));
 sg13g2_nor2_1 _1085_ (.A(net263),
    .B(_0448_),
    .Y(_0449_));
 sg13g2_and2_1 _1086_ (.A(net263),
    .B(_0448_),
    .X(_0450_));
 sg13g2_nor3_1 _1087_ (.A(net106),
    .B(net264),
    .C(_0450_),
    .Y(_0054_));
 sg13g2_nor2_1 _1088_ (.A(net269),
    .B(_0450_),
    .Y(_0451_));
 sg13g2_and2_1 _1089_ (.A(net269),
    .B(_0450_),
    .X(_0452_));
 sg13g2_nor3_1 _1090_ (.A(net106),
    .B(_0451_),
    .C(_0452_),
    .Y(_0055_));
 sg13g2_nor2_1 _1091_ (.A(net248),
    .B(_0452_),
    .Y(_0453_));
 sg13g2_and3_1 _1092_ (.X(_0454_),
    .A(\ChiselTop.tinySynth.osc.square.cnt[29] ),
    .B(net248),
    .C(_0450_));
 sg13g2_nor3_1 _1093_ (.A(net106),
    .B(net249),
    .C(_0454_),
    .Y(_0056_));
 sg13g2_nor2_1 _1094_ (.A(net214),
    .B(_0454_),
    .Y(_0455_));
 sg13g2_nor2_1 _1095_ (.A(_0368_),
    .B(_0437_),
    .Y(_0456_));
 sg13g2_nor3_1 _1096_ (.A(net106),
    .B(net215),
    .C(_0456_),
    .Y(_0057_));
 sg13g2_and2_1 _1097_ (.A(net135),
    .B(net151),
    .X(_0058_));
 sg13g2_o21ai_1 _1098_ (.B1(net135),
    .Y(_0457_),
    .A1(net166),
    .A2(\ChiselTop.tinySynth.pwm.counter[1] ));
 sg13g2_a21oi_1 _1099_ (.A1(net166),
    .A2(\ChiselTop.tinySynth.pwm.counter[1] ),
    .Y(_0059_),
    .B1(_0457_));
 sg13g2_a21oi_1 _1100_ (.A1(\ChiselTop.tinySynth.pwm.counter[0] ),
    .A2(\ChiselTop.tinySynth.pwm.counter[1] ),
    .Y(_0458_),
    .B1(net159));
 sg13g2_nand3_1 _1101_ (.B(net159),
    .C(\ChiselTop.tinySynth.pwm.counter[1] ),
    .A(net166),
    .Y(_0459_));
 sg13g2_nand2_1 _1102_ (.Y(_0460_),
    .A(net135),
    .B(_0459_));
 sg13g2_nor2_1 _1103_ (.A(net160),
    .B(_0460_),
    .Y(_0060_));
 sg13g2_and2_1 _1104_ (.A(_0144_),
    .B(_0459_),
    .X(_0461_));
 sg13g2_nor2_1 _1105_ (.A(_0144_),
    .B(_0459_),
    .Y(_0462_));
 sg13g2_nor3_1 _1106_ (.A(net133),
    .B(net303),
    .C(_0462_),
    .Y(_0061_));
 sg13g2_and2_1 _1107_ (.A(net274),
    .B(_0462_),
    .X(_0463_));
 sg13g2_o21ai_1 _1108_ (.B1(net135),
    .Y(_0464_),
    .A1(net274),
    .A2(_0462_));
 sg13g2_nor2_1 _1109_ (.A(_0463_),
    .B(net275),
    .Y(_0062_));
 sg13g2_xnor2_1 _1110_ (.Y(_0465_),
    .A(net272),
    .B(_0463_));
 sg13g2_nor2_1 _1111_ (.A(net133),
    .B(net273),
    .Y(_0063_));
 sg13g2_a21oi_1 _1112_ (.A1(\ChiselTop.tinySynth.pwm.counter[5] ),
    .A2(_0463_),
    .Y(_0466_),
    .B1(net172));
 sg13g2_nand3_1 _1113_ (.B(\ChiselTop.tinySynth.pwm.counter[5] ),
    .C(_0463_),
    .A(net172),
    .Y(_0467_));
 sg13g2_nand2_1 _1114_ (.Y(_0468_),
    .A(net134),
    .B(_0467_));
 sg13g2_nor2_1 _1115_ (.A(net173),
    .B(_0468_),
    .Y(_0064_));
 sg13g2_o21ai_1 _1116_ (.B1(net134),
    .Y(_0469_),
    .A1(_0143_),
    .A2(_0467_));
 sg13g2_a21oi_1 _1117_ (.A1(_0143_),
    .A2(_0467_),
    .Y(_0065_),
    .B1(_0469_));
 sg13g2_and2_1 _1118_ (.A(net140),
    .B(net1),
    .X(_0066_));
 sg13g2_nor3_1 _1119_ (.A(net304),
    .B(net293),
    .C(net241),
    .Y(_0470_));
 sg13g2_or4_2 _1120_ (.A(net176),
    .B(\ChiselTop.tinySynth.uart.rx.cntReg[2] ),
    .C(\ChiselTop.tinySynth.uart.rx.cntReg[1] ),
    .D(\ChiselTop.tinySynth.uart.rx.cntReg[0] ),
    .X(_0471_));
 sg13g2_nor3_1 _1121_ (.A(net312),
    .B(net307),
    .C(_0471_),
    .Y(_0472_));
 sg13g2_nor4_2 _1122_ (.A(\ChiselTop.tinySynth.uart.rx.cntReg[6] ),
    .B(\ChiselTop.tinySynth.uart.rx.cntReg[5] ),
    .C(\ChiselTop.tinySynth.uart.rx.cntReg[4] ),
    .Y(_0473_),
    .D(_0471_));
 sg13g2_nand2b_1 _1123_ (.Y(_0474_),
    .B(_0473_),
    .A_N(\ChiselTop.tinySynth.uart.rx.cntReg[7] ));
 sg13g2_or3_2 _1124_ (.A(net193),
    .B(\ChiselTop.tinySynth.uart.rx.cntReg[8] ),
    .C(_0474_),
    .X(_0475_));
 sg13g2_nor3_1 _1125_ (.A(\ChiselTop.tinySynth.uart.rx.cntReg[11] ),
    .B(\ChiselTop.tinySynth.uart.rx.cntReg[10] ),
    .C(_0475_),
    .Y(_0476_));
 sg13g2_nor4_2 _1126_ (.A(net228),
    .B(\ChiselTop.tinySynth.uart.rx.cntReg[11] ),
    .C(\ChiselTop.tinySynth.uart.rx.cntReg[10] ),
    .Y(_0477_),
    .D(_0475_));
 sg13g2_nand2b_2 _1127_ (.Y(_0478_),
    .B(_0477_),
    .A_N(net186));
 sg13g2_nor3_1 _1128_ (.A(\ChiselTop.tinySynth.uart.rx.cntReg[15] ),
    .B(\ChiselTop.tinySynth.uart.rx.cntReg[14] ),
    .C(_0478_),
    .Y(_0479_));
 sg13g2_nor4_2 _1129_ (.A(\ChiselTop.tinySynth.uart.rx.cntReg[16] ),
    .B(\ChiselTop.tinySynth.uart.rx.cntReg[15] ),
    .C(\ChiselTop.tinySynth.uart.rx.cntReg[14] ),
    .Y(_0480_),
    .D(_0478_));
 sg13g2_nand2b_1 _1130_ (.Y(_0481_),
    .B(_0480_),
    .A_N(net196));
 sg13g2_nor3_1 _1131_ (.A(\ChiselTop.tinySynth.uart.rx.cntReg[19] ),
    .B(\ChiselTop.tinySynth.uart.rx.cntReg[18] ),
    .C(_0481_),
    .Y(_0482_));
 sg13g2_nor2_1 _1132_ (.A(\ChiselTop.tinySynth.uart.rx.bitsReg[1] ),
    .B(net222),
    .Y(_0483_));
 sg13g2_nor4_2 _1133_ (.A(net191),
    .B(\ChiselTop.tinySynth.uart.rx.bitsReg[2] ),
    .C(\ChiselTop.tinySynth.uart.rx.bitsReg[1] ),
    .Y(_0484_),
    .D(\ChiselTop.tinySynth.uart.rx.bitsReg[0] ));
 sg13g2_nor2b_1 _1134_ (.A(_0484_),
    .B_N(net116),
    .Y(_0485_));
 sg13g2_o21ai_1 _1135_ (.B1(net134),
    .Y(_0486_),
    .A1(\ChiselTop.tinySynth.midi._GEN_0[0] ),
    .A2(net113));
 sg13g2_a21oi_1 _1136_ (.A1(_0122_),
    .A2(net113),
    .Y(_0067_),
    .B1(_0486_));
 sg13g2_o21ai_1 _1137_ (.B1(net134),
    .Y(_0487_),
    .A1(net230),
    .A2(net113));
 sg13g2_a21oi_1 _1138_ (.A1(_0120_),
    .A2(net113),
    .Y(_0068_),
    .B1(_0487_));
 sg13g2_o21ai_1 _1139_ (.B1(net137),
    .Y(_0488_),
    .A1(net260),
    .A2(net115));
 sg13g2_a21oi_1 _1140_ (.A1(_0128_),
    .A2(net115),
    .Y(_0069_),
    .B1(_0488_));
 sg13g2_o21ai_1 _1141_ (.B1(net137),
    .Y(_0489_),
    .A1(net202),
    .A2(net113));
 sg13g2_a21oi_1 _1142_ (.A1(_0114_),
    .A2(net113),
    .Y(_0070_),
    .B1(_0489_));
 sg13g2_o21ai_1 _1143_ (.B1(net134),
    .Y(_0490_),
    .A1(net168),
    .A2(net113));
 sg13g2_a21oi_1 _1144_ (.A1(_0113_),
    .A2(net113),
    .Y(_0071_),
    .B1(_0490_));
 sg13g2_o21ai_1 _1145_ (.B1(net138),
    .Y(_0491_),
    .A1(net184),
    .A2(net114));
 sg13g2_a21oi_1 _1146_ (.A1(_0112_),
    .A2(net114),
    .Y(_0072_),
    .B1(_0491_));
 sg13g2_o21ai_1 _1147_ (.B1(net137),
    .Y(_0492_),
    .A1(net175),
    .A2(net114));
 sg13g2_a21oi_1 _1148_ (.A1(_0111_),
    .A2(net115),
    .Y(_0073_),
    .B1(_0492_));
 sg13g2_o21ai_1 _1149_ (.B1(net137),
    .Y(_0493_),
    .A1(net170),
    .A2(net115));
 sg13g2_a21oi_1 _1150_ (.A1(_0127_),
    .A2(net115),
    .Y(_0074_),
    .B1(_0493_));
 sg13g2_o21ai_1 _1151_ (.B1(_0484_),
    .Y(_0494_),
    .A1(\ChiselTop.tinySynth.uart.rx.rxReg ),
    .A2(_0140_));
 sg13g2_inv_1 _1152_ (.Y(_0495_),
    .A(_0494_));
 sg13g2_nand2_1 _1153_ (.Y(_0496_),
    .A(_0482_),
    .B(_0495_));
 sg13g2_inv_1 _1154_ (.Y(_0497_),
    .A(_0496_));
 sg13g2_o21ai_1 _1155_ (.B1(net134),
    .Y(_0075_),
    .A1(net241),
    .A2(_0497_));
 sg13g2_nand2b_1 _1156_ (.Y(_0498_),
    .B(net134),
    .A_N(net116));
 sg13g2_xor2_1 _1157_ (.B(net241),
    .A(net293),
    .X(_0499_));
 sg13g2_nor2_1 _1158_ (.A(net112),
    .B(_0499_),
    .Y(_0076_));
 sg13g2_o21ai_1 _1159_ (.B1(net304),
    .Y(_0500_),
    .A1(net293),
    .A2(net241));
 sg13g2_nor2b_1 _1160_ (.A(_0470_),
    .B_N(_0500_),
    .Y(_0501_));
 sg13g2_nor2_1 _1161_ (.A(net112),
    .B(_0501_),
    .Y(_0077_));
 sg13g2_nor2_2 _1162_ (.A(net133),
    .B(net114),
    .Y(_0502_));
 sg13g2_nand2_1 _1163_ (.Y(_0503_),
    .A(_0496_),
    .B(_0502_));
 sg13g2_nand2b_1 _1164_ (.Y(_0504_),
    .B(net176),
    .A_N(_0470_));
 sg13g2_a21oi_1 _1165_ (.A1(_0471_),
    .A2(net177),
    .Y(_0078_),
    .B1(_0503_));
 sg13g2_xor2_1 _1166_ (.B(_0471_),
    .A(net307),
    .X(_0505_));
 sg13g2_o21ai_1 _1167_ (.B1(_0502_),
    .Y(_0079_),
    .A1(net116),
    .A2(_0505_));
 sg13g2_o21ai_1 _1168_ (.B1(net312),
    .Y(_0506_),
    .A1(\ChiselTop.tinySynth.uart.rx.cntReg[4] ),
    .A2(_0471_));
 sg13g2_nor2b_1 _1169_ (.A(_0472_),
    .B_N(net313),
    .Y(_0507_));
 sg13g2_o21ai_1 _1170_ (.B1(_0502_),
    .Y(_0080_),
    .A1(net116),
    .A2(_0507_));
 sg13g2_xnor2_1 _1171_ (.Y(_0508_),
    .A(net223),
    .B(_0472_));
 sg13g2_nor2_1 _1172_ (.A(net112),
    .B(net224),
    .Y(_0081_));
 sg13g2_nand2_1 _1173_ (.Y(_0509_),
    .A(_0473_),
    .B(_0496_));
 sg13g2_a21oi_1 _1174_ (.A1(net155),
    .A2(_0509_),
    .Y(_0510_),
    .B1(net133));
 sg13g2_o21ai_1 _1175_ (.B1(_0510_),
    .Y(_0082_),
    .A1(net155),
    .A2(_0509_));
 sg13g2_xor2_1 _1176_ (.B(_0474_),
    .A(net298),
    .X(_0511_));
 sg13g2_o21ai_1 _1177_ (.B1(_0502_),
    .Y(_0083_),
    .A1(net116),
    .A2(net299));
 sg13g2_o21ai_1 _1178_ (.B1(net193),
    .Y(_0512_),
    .A1(\ChiselTop.tinySynth.uart.rx.cntReg[8] ),
    .A2(_0474_));
 sg13g2_a21oi_1 _1179_ (.A1(_0475_),
    .A2(net194),
    .Y(_0084_),
    .B1(_0503_));
 sg13g2_nor2_1 _1180_ (.A(_0141_),
    .B(_0475_),
    .Y(_0513_));
 sg13g2_xnor2_1 _1181_ (.Y(_0514_),
    .A(net162),
    .B(_0475_));
 sg13g2_nor2_1 _1182_ (.A(net111),
    .B(net163),
    .Y(_0085_));
 sg13g2_xnor2_1 _1183_ (.Y(_0515_),
    .A(net259),
    .B(_0513_));
 sg13g2_nor2_1 _1184_ (.A(net112),
    .B(_0515_),
    .Y(_0086_));
 sg13g2_xnor2_1 _1185_ (.Y(_0516_),
    .A(net228),
    .B(_0476_));
 sg13g2_nor2_1 _1186_ (.A(net111),
    .B(net229),
    .Y(_0087_));
 sg13g2_nand2b_1 _1187_ (.Y(_0517_),
    .B(net186),
    .A_N(_0477_));
 sg13g2_a21oi_1 _1188_ (.A1(_0478_),
    .A2(net187),
    .Y(_0088_),
    .B1(net111));
 sg13g2_nor2_1 _1189_ (.A(_0142_),
    .B(_0478_),
    .Y(_0518_));
 sg13g2_xnor2_1 _1190_ (.Y(_0519_),
    .A(net157),
    .B(_0478_));
 sg13g2_nor2_1 _1191_ (.A(net111),
    .B(net158),
    .Y(_0089_));
 sg13g2_xnor2_1 _1192_ (.Y(_0520_),
    .A(net267),
    .B(_0518_));
 sg13g2_nor2_1 _1193_ (.A(net111),
    .B(net268),
    .Y(_0090_));
 sg13g2_xnor2_1 _1194_ (.Y(_0521_),
    .A(net243),
    .B(_0479_));
 sg13g2_nor2_1 _1195_ (.A(net111),
    .B(net244),
    .Y(_0091_));
 sg13g2_nand2b_1 _1196_ (.Y(_0522_),
    .B(net196),
    .A_N(_0480_));
 sg13g2_a21oi_1 _1197_ (.A1(_0481_),
    .A2(net197),
    .Y(_0092_),
    .B1(net111));
 sg13g2_nand3b_1 _1198_ (.B(net164),
    .C(_0480_),
    .Y(_0523_),
    .A_N(net196));
 sg13g2_xnor2_1 _1199_ (.Y(_0524_),
    .A(net164),
    .B(_0481_));
 sg13g2_nor2_1 _1200_ (.A(net111),
    .B(net165),
    .Y(_0093_));
 sg13g2_xor2_1 _1201_ (.B(_0523_),
    .A(net239),
    .X(_0525_));
 sg13g2_nor2_1 _1202_ (.A(net112),
    .B(net240),
    .Y(_0094_));
 sg13g2_nand2_1 _1203_ (.Y(_0526_),
    .A(_0126_),
    .B(net115));
 sg13g2_nand2_1 _1204_ (.Y(_0527_),
    .A(net116),
    .B(_0494_));
 sg13g2_inv_1 _1205_ (.Y(_0528_),
    .A(_0527_));
 sg13g2_nand2_1 _1206_ (.Y(_0529_),
    .A(net213),
    .B(_0527_));
 sg13g2_a21oi_1 _1207_ (.A1(_0526_),
    .A2(_0529_),
    .Y(_0095_),
    .B1(_0138_));
 sg13g2_o21ai_1 _1208_ (.B1(net136),
    .Y(_0530_),
    .A1(_0125_),
    .A2(_0526_));
 sg13g2_a21oi_1 _1209_ (.A1(_0125_),
    .A2(_0526_),
    .Y(_0096_),
    .B1(_0530_));
 sg13g2_xor2_1 _1210_ (.B(_0483_),
    .A(net295),
    .X(_0531_));
 sg13g2_a22oi_1 _1211_ (.Y(_0532_),
    .B1(_0531_),
    .B2(net115),
    .A2(_0527_),
    .A1(net295));
 sg13g2_nor2_1 _1212_ (.A(net133),
    .B(_0532_),
    .Y(_0097_));
 sg13g2_nand3b_1 _1213_ (.B(net116),
    .C(_0483_),
    .Y(_0533_),
    .A_N(\ChiselTop.tinySynth.uart.rx.bitsReg[2] ));
 sg13g2_a22oi_1 _1214_ (.Y(_0534_),
    .B1(_0533_),
    .B2(net191),
    .A2(_0528_),
    .A1(_0484_));
 sg13g2_nor2_1 _1215_ (.A(net133),
    .B(net192),
    .Y(_0098_));
 sg13g2_nor4_1 _1216_ (.A(net191),
    .B(\ChiselTop.tinySynth.uart.rx.bitsReg[2] ),
    .C(\ChiselTop.tinySynth.uart.rx.bitsReg[1] ),
    .D(_0126_),
    .Y(_0535_));
 sg13g2_a21oi_1 _1217_ (.A1(net116),
    .A2(_0535_),
    .Y(_0536_),
    .B1(net245));
 sg13g2_nor2_1 _1218_ (.A(_0150_),
    .B(net246),
    .Y(_0099_));
 sg13g2_nor3_1 _1219_ (.A(_0124_),
    .B(_0024_),
    .C(_0153_),
    .Y(_0537_));
 sg13g2_o21ai_1 _1220_ (.B1(net245),
    .Y(_0538_),
    .A1(\ChiselTop.tinySynth.midi.regState[0] ),
    .A2(\ChiselTop.tinySynth.midi.regState[2] ));
 sg13g2_nor2_1 _1221_ (.A(_0537_),
    .B(_0538_),
    .Y(_0539_));
 sg13g2_nand2_1 _1222_ (.Y(_0540_),
    .A(_0154_),
    .B(_0539_));
 sg13g2_o21ai_1 _1223_ (.B1(net138),
    .Y(_0541_),
    .A1(\ChiselTop.tinySynth.midi._GEN_0[0] ),
    .A2(net117));
 sg13g2_a21oi_1 _1224_ (.A1(_0123_),
    .A2(net117),
    .Y(_0100_),
    .B1(_0541_));
 sg13g2_o21ai_1 _1225_ (.B1(net138),
    .Y(_0542_),
    .A1(net230),
    .A2(net118));
 sg13g2_a21oi_1 _1226_ (.A1(_0121_),
    .A2(net118),
    .Y(_0101_),
    .B1(_0542_));
 sg13g2_nor2_1 _1227_ (.A(net260),
    .B(net118),
    .Y(_0543_));
 sg13g2_a21oi_1 _1228_ (.A1(_0154_),
    .A2(_0539_),
    .Y(_0544_),
    .B1(net285));
 sg13g2_nor3_1 _1229_ (.A(net133),
    .B(_0543_),
    .C(_0544_),
    .Y(_0102_));
 sg13g2_nor3_1 _1230_ (.A(\ChiselTop.tinySynth.midi.regState[0] ),
    .B(_0537_),
    .C(_0538_),
    .Y(_0545_));
 sg13g2_a22oi_1 _1231_ (.Y(_0546_),
    .B1(_0545_),
    .B2(net202),
    .A2(net118),
    .A1(net278));
 sg13g2_nor2_1 _1232_ (.A(net133),
    .B(net279),
    .Y(_0103_));
 sg13g2_o21ai_1 _1233_ (.B1(net138),
    .Y(_0547_),
    .A1(net168),
    .A2(net117));
 sg13g2_a21oi_1 _1234_ (.A1(_0117_),
    .A2(net117),
    .Y(_0104_),
    .B1(_0547_));
 sg13g2_o21ai_1 _1235_ (.B1(net138),
    .Y(_0548_),
    .A1(net184),
    .A2(net117));
 sg13g2_a21oi_1 _1236_ (.A1(_0116_),
    .A2(net117),
    .Y(_0105_),
    .B1(_0548_));
 sg13g2_o21ai_1 _1237_ (.B1(net138),
    .Y(_0549_),
    .A1(net175),
    .A2(net117));
 sg13g2_a21oi_1 _1238_ (.A1(_0115_),
    .A2(net117),
    .Y(_0106_),
    .B1(_0549_));
 sg13g2_o21ai_1 _1239_ (.B1(net138),
    .Y(_0550_),
    .A1(\ChiselTop.tinySynth.midi.io_midiOut_bits_hdr_channel[0] ),
    .A2(net122));
 sg13g2_a21oi_1 _1240_ (.A1(_0114_),
    .A2(net122),
    .Y(_0107_),
    .B1(_0550_));
 sg13g2_o21ai_1 _1241_ (.B1(net138),
    .Y(_0551_),
    .A1(\ChiselTop.tinySynth.midi.io_midiOut_bits_hdr_channel[1] ),
    .A2(net122));
 sg13g2_a21oi_1 _1242_ (.A1(_0113_),
    .A2(net122),
    .Y(_0108_),
    .B1(_0551_));
 sg13g2_o21ai_1 _1243_ (.B1(net136),
    .Y(_0552_),
    .A1(net251),
    .A2(net122));
 sg13g2_a21oi_1 _1244_ (.A1(_0112_),
    .A2(net122),
    .Y(_0109_),
    .B1(_0552_));
 sg13g2_o21ai_1 _1245_ (.B1(net136),
    .Y(_0553_),
    .A1(\ChiselTop.tinySynth.midi.io_midiOut_bits_hdr_channel[3] ),
    .A2(net122));
 sg13g2_a21oi_1 _1246_ (.A1(_0111_),
    .A2(net122),
    .Y(_0110_),
    .B1(_0553_));
 sg13g2_dfrbp_1 _1247_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net27),
    .D(net315),
    .Q_N(_0024_),
    .Q(\ChiselTop.tinySynth.midi.regState[0] ));
 sg13g2_dfrbp_1 _1248_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net28),
    .D(net236),
    .Q_N(_0619_),
    .Q(\ChiselTop.tinySynth.midi.regState[1] ));
 sg13g2_dfrbp_1 _1249_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net71),
    .D(net287),
    .Q_N(_0620_),
    .Q(\ChiselTop.tinySynth.midi.regState[2] ));
 sg13g2_dfrbp_1 _1250_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net26),
    .D(net209),
    .Q_N(_0618_),
    .Q(\ChiselTop.tinySynth.midi.regState[3] ));
 sg13g2_dfrbp_1 _1251_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net39),
    .D(_0025_),
    .Q_N(_0617_),
    .Q(\ChiselTop.tinySynth.uart.rx.rxReg ));
 sg13g2_dfrbp_1 _1252_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net38),
    .D(_0026_),
    .Q_N(\ChiselTop.tinySynth.osc.square._cnt_T_1[0] ),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[0] ));
 sg13g2_dfrbp_1 _1253_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net37),
    .D(_0027_),
    .Q_N(_0023_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[1] ));
 sg13g2_dfrbp_1 _1254_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net36),
    .D(_0028_),
    .Q_N(_0022_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[2] ));
 sg13g2_dfrbp_1 _1255_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net35),
    .D(_0029_),
    .Q_N(_0021_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[3] ));
 sg13g2_dfrbp_1 _1256_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net34),
    .D(_0030_),
    .Q_N(_0020_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[4] ));
 sg13g2_dfrbp_1 _1257_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net33),
    .D(_0031_),
    .Q_N(_0616_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[5] ));
 sg13g2_dfrbp_1 _1258_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net32),
    .D(_0032_),
    .Q_N(_0019_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[6] ));
 sg13g2_dfrbp_1 _1259_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net31),
    .D(_0033_),
    .Q_N(_0018_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[7] ));
 sg13g2_dfrbp_1 _1260_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net30),
    .D(_0034_),
    .Q_N(_0017_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[8] ));
 sg13g2_dfrbp_1 _1261_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net29),
    .D(_0035_),
    .Q_N(_0016_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[9] ));
 sg13g2_dfrbp_1 _1262_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net25),
    .D(_0036_),
    .Q_N(_0015_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[10] ));
 sg13g2_dfrbp_1 _1263_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net150),
    .D(_0037_),
    .Q_N(_0014_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[11] ));
 sg13g2_dfrbp_1 _1264_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net149),
    .D(net183),
    .Q_N(_0013_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[12] ));
 sg13g2_dfrbp_1 _1265_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net148),
    .D(_0039_),
    .Q_N(_0615_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[13] ));
 sg13g2_dfrbp_1 _1266_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net147),
    .D(_0040_),
    .Q_N(_0012_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[14] ));
 sg13g2_dfrbp_1 _1267_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net146),
    .D(_0041_),
    .Q_N(_0011_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[15] ));
 sg13g2_dfrbp_1 _1268_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net145),
    .D(net207),
    .Q_N(_0010_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[16] ));
 sg13g2_dfrbp_1 _1269_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net144),
    .D(_0043_),
    .Q_N(_0009_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[17] ));
 sg13g2_dfrbp_1 _1270_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net143),
    .D(_0044_),
    .Q_N(_0008_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[18] ));
 sg13g2_dfrbp_1 _1271_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net142),
    .D(_0045_),
    .Q_N(_0614_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[19] ));
 sg13g2_dfrbp_1 _1272_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net141),
    .D(_0046_),
    .Q_N(_0007_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[20] ));
 sg13g2_dfrbp_1 _1273_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net105),
    .D(_0047_),
    .Q_N(_0613_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[21] ));
 sg13g2_dfrbp_1 _1274_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net104),
    .D(_0048_),
    .Q_N(_0612_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[22] ));
 sg13g2_dfrbp_1 _1275_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net103),
    .D(net284),
    .Q_N(_0611_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[23] ));
 sg13g2_dfrbp_1 _1276_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net102),
    .D(_0050_),
    .Q_N(_0610_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[24] ));
 sg13g2_dfrbp_1 _1277_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net101),
    .D(net201),
    .Q_N(_0609_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[25] ));
 sg13g2_dfrbp_1 _1278_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net100),
    .D(_0052_),
    .Q_N(_0608_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[26] ));
 sg13g2_dfrbp_1 _1279_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net99),
    .D(net227),
    .Q_N(_0607_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[27] ));
 sg13g2_dfrbp_1 _1280_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net98),
    .D(_0054_),
    .Q_N(_0606_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[28] ));
 sg13g2_dfrbp_1 _1281_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net97),
    .D(_0055_),
    .Q_N(_0605_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[29] ));
 sg13g2_dfrbp_1 _1282_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net96),
    .D(net250),
    .Q_N(_0604_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[30] ));
 sg13g2_dfrbp_1 _1283_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net95),
    .D(net216),
    .Q_N(_0603_),
    .Q(\ChiselTop.tinySynth.osc.square.cnt[31] ));
 sg13g2_dfrbp_1 _1284_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net94),
    .D(_0058_),
    .Q_N(\ChiselTop.tinySynth.pwm._counter_T_1[0] ),
    .Q(\ChiselTop.tinySynth.pwm.counter[0] ));
 sg13g2_dfrbp_1 _1285_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net93),
    .D(net167),
    .Q_N(_0602_),
    .Q(\ChiselTop.tinySynth.pwm.counter[1] ));
 sg13g2_dfrbp_1 _1286_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net92),
    .D(net161),
    .Q_N(_0601_),
    .Q(\ChiselTop.tinySynth.pwm.counter[2] ));
 sg13g2_dfrbp_1 _1287_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net91),
    .D(_0061_),
    .Q_N(_0600_),
    .Q(\ChiselTop.tinySynth.pwm.counter[3] ));
 sg13g2_dfrbp_1 _1288_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net90),
    .D(_0062_),
    .Q_N(_0599_),
    .Q(\ChiselTop.tinySynth.pwm.counter[4] ));
 sg13g2_dfrbp_1 _1289_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net89),
    .D(_0063_),
    .Q_N(_0598_),
    .Q(\ChiselTop.tinySynth.pwm.counter[5] ));
 sg13g2_dfrbp_1 _1290_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net88),
    .D(net174),
    .Q_N(_0597_),
    .Q(\ChiselTop.tinySynth.pwm.counter[6] ));
 sg13g2_dfrbp_1 _1291_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net87),
    .D(net180),
    .Q_N(_0596_),
    .Q(\ChiselTop.tinySynth.pwm.counter[7] ));
 sg13g2_dfrbp_1 _1292_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net59),
    .D(_0066_),
    .Q_N(_0621_),
    .Q(\ChiselTop.tinySynth.uart.rx.rxReg_REG ));
 sg13g2_dfrbp_1 _1293_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net86),
    .D(net152),
    .Q_N(_0595_),
    .Q(\ChiselTop.tinySynth.uart.rx.falling_REG ));
 sg13g2_dfrbp_1 _1294_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net85),
    .D(net231),
    .Q_N(_0594_),
    .Q(\ChiselTop.tinySynth.midi._GEN_0[0] ));
 sg13g2_dfrbp_1 _1295_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net83),
    .D(_0068_),
    .Q_N(_0593_),
    .Q(\ChiselTop.tinySynth.midi._GEN_0[1] ));
 sg13g2_dfrbp_1 _1296_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net81),
    .D(_0069_),
    .Q_N(_0592_),
    .Q(\ChiselTop.tinySynth.midi._GEN_0[2] ));
 sg13g2_dfrbp_1 _1297_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net79),
    .D(_0070_),
    .Q_N(_0591_),
    .Q(\ChiselTop.tinySynth.midi.hdr_msgType[3] ));
 sg13g2_dfrbp_1 _1298_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net77),
    .D(_0071_),
    .Q_N(_0590_),
    .Q(\ChiselTop.tinySynth.midi._GEN_0[4] ));
 sg13g2_dfrbp_1 _1299_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net75),
    .D(_0072_),
    .Q_N(_0589_),
    .Q(\ChiselTop.tinySynth.midi._GEN_0[5] ));
 sg13g2_dfrbp_1 _1300_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net73),
    .D(_0073_),
    .Q_N(_0588_),
    .Q(\ChiselTop.tinySynth.midi._GEN_0[6] ));
 sg13g2_dfrbp_1 _1301_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net70),
    .D(_0074_),
    .Q_N(_0587_),
    .Q(\ChiselTop.tinySynth.midi.hdr_channel[3] ));
 sg13g2_dfrbp_1 _1302_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net68),
    .D(net242),
    .Q_N(_0586_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[0] ));
 sg13g2_dfrbp_1 _1303_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net66),
    .D(_0076_),
    .Q_N(_0585_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[1] ));
 sg13g2_dfrbp_1 _1304_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net64),
    .D(_0077_),
    .Q_N(_0584_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[2] ));
 sg13g2_dfrbp_1 _1305_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net62),
    .D(net178),
    .Q_N(_0583_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[3] ));
 sg13g2_dfrbp_1 _1306_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net60),
    .D(_0079_),
    .Q_N(_0582_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[4] ));
 sg13g2_dfrbp_1 _1307_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net58),
    .D(_0080_),
    .Q_N(_0581_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[5] ));
 sg13g2_dfrbp_1 _1308_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net56),
    .D(_0081_),
    .Q_N(_0580_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[6] ));
 sg13g2_dfrbp_1 _1309_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net54),
    .D(net156),
    .Q_N(_0579_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[7] ));
 sg13g2_dfrbp_1 _1310_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net52),
    .D(_0083_),
    .Q_N(_0578_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[8] ));
 sg13g2_dfrbp_1 _1311_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net50),
    .D(net195),
    .Q_N(_0577_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[9] ));
 sg13g2_dfrbp_1 _1312_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net48),
    .D(_0085_),
    .Q_N(_0006_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[10] ));
 sg13g2_dfrbp_1 _1313_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net46),
    .D(_0086_),
    .Q_N(_0576_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[11] ));
 sg13g2_dfrbp_1 _1314_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net44),
    .D(_0087_),
    .Q_N(_0575_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[12] ));
 sg13g2_dfrbp_1 _1315_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net42),
    .D(net188),
    .Q_N(_0574_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[13] ));
 sg13g2_dfrbp_1 _1316_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net40),
    .D(_0089_),
    .Q_N(_0005_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[14] ));
 sg13g2_dfrbp_1 _1317_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net82),
    .D(_0090_),
    .Q_N(_0573_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[15] ));
 sg13g2_dfrbp_1 _1318_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net78),
    .D(_0091_),
    .Q_N(_0572_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[16] ));
 sg13g2_dfrbp_1 _1319_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net74),
    .D(net198),
    .Q_N(_0571_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[17] ));
 sg13g2_dfrbp_1 _1320_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net69),
    .D(_0093_),
    .Q_N(_0004_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[18] ));
 sg13g2_dfrbp_1 _1321_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net65),
    .D(_0094_),
    .Q_N(_0570_),
    .Q(\ChiselTop.tinySynth.uart.rx.cntReg[19] ));
 sg13g2_dfrbp_1 _1322_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net61),
    .D(_0095_),
    .Q_N(_0569_),
    .Q(\ChiselTop.tinySynth.uart.rx.bitsReg[0] ));
 sg13g2_dfrbp_1 _1323_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net57),
    .D(_0096_),
    .Q_N(_0568_),
    .Q(\ChiselTop.tinySynth.uart.rx.bitsReg[1] ));
 sg13g2_dfrbp_1 _1324_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net53),
    .D(_0097_),
    .Q_N(_0567_),
    .Q(\ChiselTop.tinySynth.uart.rx.bitsReg[2] ));
 sg13g2_dfrbp_1 _1325_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net49),
    .D(_0098_),
    .Q_N(_0566_),
    .Q(\ChiselTop.tinySynth.uart.rx.bitsReg[3] ));
 sg13g2_dfrbp_1 _1326_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net45),
    .D(net247),
    .Q_N(_0565_),
    .Q(\ChiselTop.tinySynth.midi.io_uartIn_valid ));
 sg13g2_dfrbp_1 _1327_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net41),
    .D(net233),
    .Q_N(_0564_),
    .Q(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[0] ));
 sg13g2_dfrbp_1 _1328_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net80),
    .D(_0101_),
    .Q_N(_0563_),
    .Q(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[1] ));
 sg13g2_dfrbp_1 _1329_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net72),
    .D(_0102_),
    .Q_N(_0562_),
    .Q(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[2] ));
 sg13g2_dfrbp_1 _1330_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net63),
    .D(_0103_),
    .Q_N(_0561_),
    .Q(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[3] ));
 sg13g2_dfrbp_1 _1331_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net55),
    .D(_0104_),
    .Q_N(_0560_),
    .Q(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[4] ));
 sg13g2_dfrbp_1 _1332_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net47),
    .D(_0105_),
    .Q_N(_0559_),
    .Q(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[5] ));
 sg13g2_dfrbp_1 _1333_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net84),
    .D(_0106_),
    .Q_N(_0558_),
    .Q(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[6] ));
 sg13g2_dfrbp_1 _1334_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net67),
    .D(net169),
    .Q_N(_0557_),
    .Q(\ChiselTop.tinySynth.midi.io_midiOut_bits_hdr_channel[0] ));
 sg13g2_dfrbp_1 _1335_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net51),
    .D(net185),
    .Q_N(_0556_),
    .Q(\ChiselTop.tinySynth.midi.io_midiOut_bits_hdr_channel[1] ));
 sg13g2_dfrbp_1 _1336_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net76),
    .D(net252),
    .Q_N(_0555_),
    .Q(\ChiselTop.tinySynth.midi.io_midiOut_bits_hdr_channel[2] ));
 sg13g2_dfrbp_1 _1337_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net43),
    .D(net171),
    .Q_N(_0554_),
    .Q(\ChiselTop.tinySynth.midi.io_midiOut_bits_hdr_channel[3] ));
 sg13g2_tiehi _1250__26 (.L_HI(net26));
 sg13g2_tiehi _1247__27 (.L_HI(net27));
 sg13g2_tiehi _1248__28 (.L_HI(net28));
 sg13g2_tiehi _1261__29 (.L_HI(net29));
 sg13g2_tiehi _1260__30 (.L_HI(net30));
 sg13g2_tiehi _1259__31 (.L_HI(net31));
 sg13g2_tiehi _1258__32 (.L_HI(net32));
 sg13g2_tiehi _1257__33 (.L_HI(net33));
 sg13g2_tiehi _1256__34 (.L_HI(net34));
 sg13g2_tiehi _1255__35 (.L_HI(net35));
 sg13g2_tiehi _1254__36 (.L_HI(net36));
 sg13g2_tiehi _1253__37 (.L_HI(net37));
 sg13g2_tiehi _1252__38 (.L_HI(net38));
 sg13g2_tiehi _1251__39 (.L_HI(net39));
 sg13g2_tiehi _1316__40 (.L_HI(net40));
 sg13g2_tiehi _1327__41 (.L_HI(net41));
 sg13g2_tiehi _1315__42 (.L_HI(net42));
 sg13g2_tiehi _1337__43 (.L_HI(net43));
 sg13g2_tiehi _1314__44 (.L_HI(net44));
 sg13g2_tiehi _1326__45 (.L_HI(net45));
 sg13g2_tiehi _1313__46 (.L_HI(net46));
 sg13g2_tiehi _1332__47 (.L_HI(net47));
 sg13g2_tiehi _1312__48 (.L_HI(net48));
 sg13g2_tiehi _1325__49 (.L_HI(net49));
 sg13g2_tiehi _1311__50 (.L_HI(net50));
 sg13g2_tiehi _1335__51 (.L_HI(net51));
 sg13g2_tiehi _1310__52 (.L_HI(net52));
 sg13g2_tiehi _1324__53 (.L_HI(net53));
 sg13g2_tiehi _1309__54 (.L_HI(net54));
 sg13g2_tiehi _1331__55 (.L_HI(net55));
 sg13g2_tiehi _1308__56 (.L_HI(net56));
 sg13g2_tiehi _1323__57 (.L_HI(net57));
 sg13g2_tiehi _1307__58 (.L_HI(net58));
 sg13g2_tiehi _1292__59 (.L_HI(net59));
 sg13g2_tiehi _1306__60 (.L_HI(net60));
 sg13g2_tiehi _1322__61 (.L_HI(net61));
 sg13g2_tiehi _1305__62 (.L_HI(net62));
 sg13g2_tiehi _1330__63 (.L_HI(net63));
 sg13g2_tiehi _1304__64 (.L_HI(net64));
 sg13g2_tiehi _1321__65 (.L_HI(net65));
 sg13g2_tiehi _1303__66 (.L_HI(net66));
 sg13g2_tiehi _1334__67 (.L_HI(net67));
 sg13g2_tiehi _1302__68 (.L_HI(net68));
 sg13g2_tiehi _1320__69 (.L_HI(net69));
 sg13g2_tiehi _1301__70 (.L_HI(net70));
 sg13g2_tiehi _1249__71 (.L_HI(net71));
 sg13g2_tiehi _1329__72 (.L_HI(net72));
 sg13g2_tiehi _1300__73 (.L_HI(net73));
 sg13g2_tiehi _1319__74 (.L_HI(net74));
 sg13g2_tiehi _1299__75 (.L_HI(net75));
 sg13g2_tiehi _1336__76 (.L_HI(net76));
 sg13g2_tiehi _1298__77 (.L_HI(net77));
 sg13g2_tiehi _1318__78 (.L_HI(net78));
 sg13g2_tiehi _1297__79 (.L_HI(net79));
 sg13g2_tiehi _1328__80 (.L_HI(net80));
 sg13g2_tiehi _1296__81 (.L_HI(net81));
 sg13g2_tiehi _1317__82 (.L_HI(net82));
 sg13g2_tiehi _1295__83 (.L_HI(net83));
 sg13g2_tiehi _1333__84 (.L_HI(net84));
 sg13g2_tiehi _1294__85 (.L_HI(net85));
 sg13g2_tiehi _1293__86 (.L_HI(net86));
 sg13g2_tiehi _1291__87 (.L_HI(net87));
 sg13g2_tiehi _1290__88 (.L_HI(net88));
 sg13g2_tiehi _1289__89 (.L_HI(net89));
 sg13g2_tiehi _1288__90 (.L_HI(net90));
 sg13g2_tiehi _1287__91 (.L_HI(net91));
 sg13g2_tiehi _1286__92 (.L_HI(net92));
 sg13g2_tiehi _1285__93 (.L_HI(net93));
 sg13g2_tiehi _1284__94 (.L_HI(net94));
 sg13g2_tiehi _1283__95 (.L_HI(net95));
 sg13g2_tiehi _1282__96 (.L_HI(net96));
 sg13g2_tiehi _1281__97 (.L_HI(net97));
 sg13g2_tiehi _1280__98 (.L_HI(net98));
 sg13g2_tiehi _1279__99 (.L_HI(net99));
 sg13g2_tiehi _1278__100 (.L_HI(net100));
 sg13g2_tiehi _1277__101 (.L_HI(net101));
 sg13g2_tiehi _1276__102 (.L_HI(net102));
 sg13g2_tiehi _1275__103 (.L_HI(net103));
 sg13g2_tiehi _1274__104 (.L_HI(net104));
 sg13g2_tiehi _1273__105 (.L_HI(net105));
 sg13g2_tiehi _1272__106 (.L_HI(net141));
 sg13g2_tiehi _1271__107 (.L_HI(net142));
 sg13g2_tiehi _1270__108 (.L_HI(net143));
 sg13g2_tiehi _1269__109 (.L_HI(net144));
 sg13g2_tiehi _1268__110 (.L_HI(net145));
 sg13g2_tiehi _1267__111 (.L_HI(net146));
 sg13g2_tiehi _1266__112 (.L_HI(net147));
 sg13g2_tiehi _1265__113 (.L_HI(net148));
 sg13g2_tiehi _1264__114 (.L_HI(net149));
 sg13g2_tiehi _1263__115 (.L_HI(net150));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_tinysynth_3 (.L_LO(net3));
 sg13g2_tielo tt_um_tinysynth_4 (.L_LO(net4));
 sg13g2_tielo tt_um_tinysynth_5 (.L_LO(net5));
 sg13g2_tielo tt_um_tinysynth_6 (.L_LO(net6));
 sg13g2_tielo tt_um_tinysynth_7 (.L_LO(net7));
 sg13g2_tielo tt_um_tinysynth_8 (.L_LO(net8));
 sg13g2_tielo tt_um_tinysynth_9 (.L_LO(net9));
 sg13g2_tielo tt_um_tinysynth_10 (.L_LO(net10));
 sg13g2_tielo tt_um_tinysynth_11 (.L_LO(net11));
 sg13g2_tielo tt_um_tinysynth_12 (.L_LO(net12));
 sg13g2_tielo tt_um_tinysynth_13 (.L_LO(net13));
 sg13g2_tielo tt_um_tinysynth_14 (.L_LO(net14));
 sg13g2_tielo tt_um_tinysynth_15 (.L_LO(net15));
 sg13g2_tielo tt_um_tinysynth_16 (.L_LO(net16));
 sg13g2_tielo tt_um_tinysynth_17 (.L_LO(net17));
 sg13g2_tielo tt_um_tinysynth_18 (.L_LO(net18));
 sg13g2_tielo tt_um_tinysynth_19 (.L_LO(net19));
 sg13g2_tielo tt_um_tinysynth_20 (.L_LO(net20));
 sg13g2_tielo tt_um_tinysynth_21 (.L_LO(net21));
 sg13g2_tielo tt_um_tinysynth_22 (.L_LO(net22));
 sg13g2_tielo tt_um_tinysynth_23 (.L_LO(net23));
 sg13g2_tielo tt_um_tinysynth_24 (.L_LO(net24));
 sg13g2_tiehi _1262__25 (.L_HI(net25));
 sg13g2_buf_1 _1452_ (.A(\ChiselTop.tinySynth.io_pwmOut ),
    .X(uo_out[0]));
 sg13g2_buf_2 fanout106 (.A(net109),
    .X(net106));
 sg13g2_buf_1 fanout107 (.A(net109),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(net109),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_0391_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_0391_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(net112),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_0498_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(net114),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(net115),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_0485_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_0482_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_0540_),
    .X(net117));
 sg13g2_buf_1 fanout118 (.A(_0540_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_0188_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_0181_),
    .X(net120));
 sg13g2_buf_1 fanout121 (.A(_0181_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_0537_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(net124),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_0164_),
    .X(net124));
 sg13g2_buf_4 fanout125 (.X(net125),
    .A(_0163_));
 sg13g2_buf_2 fanout126 (.A(_0163_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_0162_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_0161_),
    .X(net128));
 sg13g2_buf_4 fanout129 (.X(net129),
    .A(net271));
 sg13g2_buf_2 fanout130 (.A(\ChiselTop.tinySynth.osc.square.cnt[5] ),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_1 fanout132 (.A(net314),
    .X(net132));
 sg13g2_buf_4 fanout133 (.X(net133),
    .A(_0138_));
 sg13g2_buf_2 fanout134 (.A(net139),
    .X(net134));
 sg13g2_buf_1 fanout135 (.A(net139),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(net137),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(net139),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(net139),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(rst_n),
    .X(net140));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_tielo tt_um_tinysynth_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\ChiselTop.tinySynth.pwm._counter_T_1[0] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold2 (.A(\ChiselTop.tinySynth.uart.rx.rxReg ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold3 (.A(\ChiselTop.tinySynth.osc.square._cnt_T_1[0] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold4 (.A(\ChiselTop.tinySynth.uart.rx.rxReg_REG ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold5 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[7] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0082_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0005_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0519_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold9 (.A(\ChiselTop.tinySynth.pwm.counter[2] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0458_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0060_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0006_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0514_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0004_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0524_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold16 (.A(\ChiselTop.tinySynth.pwm.counter[0] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0059_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold18 (.A(\ChiselTop.tinySynth.midi._GEN_0[4] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0107_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold20 (.A(\ChiselTop.tinySynth.midi.hdr_channel[3] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0110_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold22 (.A(\ChiselTop.tinySynth.pwm.counter[6] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0466_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0064_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold25 (.A(\ChiselTop.tinySynth.midi._GEN_0[6] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold26 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[3] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0504_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0078_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold29 (.A(\ChiselTop.tinySynth.pwm.counter[7] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0065_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold31 (.A(\ChiselTop.tinySynth.osc.square.cnt[12] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0417_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0038_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold34 (.A(\ChiselTop.tinySynth.midi._GEN_0[5] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0108_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold36 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[13] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0517_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0088_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold39 (.A(\ChiselTop.tinySynth.osc.square.cnt[6] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0403_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold41 (.A(\ChiselTop.tinySynth.uart.rx.bitsReg[3] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0534_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold43 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[9] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0512_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0084_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold46 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[17] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0522_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0092_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold49 (.A(\ChiselTop.tinySynth.osc.square.cnt[25] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0443_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0051_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold52 (.A(\ChiselTop.tinySynth.midi.hdr_msgType[3] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold53 (.A(\ChiselTop.tinySynth.osc.square.cnt[5] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0401_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold55 (.A(\ChiselTop.tinySynth.osc.square.cnt[16] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0426_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0042_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold58 (.A(\ChiselTop.tinySynth.midi.regState[1] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0000_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold60 (.A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[4] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold61 (.A(\ChiselTop.tinySynth.osc.square.cnt[3] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0396_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold63 (.A(\ChiselTop.tinySynth.uart.rx.bitsReg[0] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold64 (.A(\ChiselTop.tinySynth.osc.square.cnt[31] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0455_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0057_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold67 (.A(\ChiselTop.tinySynth.osc.square.cnt[1] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0393_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0013_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0418_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0419_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold72 (.A(\ChiselTop.tinySynth.uart.rx.bitsReg[0] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold73 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[6] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0508_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold75 (.A(\ChiselTop.tinySynth.osc.square.cnt[27] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0447_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0053_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold78 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[12] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0516_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold80 (.A(\ChiselTop.tinySynth.midi._GEN_0[1] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0067_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold82 (.A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[0] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0100_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold84 (.A(\ChiselTop.tinySynth.midi.regState[2] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0159_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0002_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold87 (.A(\ChiselTop.tinySynth.osc.square.cnt[26] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0445_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold89 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[19] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0525_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold91 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[0] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0075_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold93 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[16] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0521_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold95 (.A(\ChiselTop.tinySynth.midi.io_uartIn_valid ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0536_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0099_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold98 (.A(\ChiselTop.tinySynth.osc.square.cnt[30] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0453_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0056_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold101 (.A(\ChiselTop.tinySynth.midi.io_midiOut_bits_hdr_channel[2] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0109_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold103 (.A(\ChiselTop.tinySynth.osc.square.cnt[17] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0428_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0017_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0409_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold107 (.A(\ChiselTop.tinySynth.osc.square.cnt[7] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0405_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold109 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[11] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold110 (.A(\ChiselTop.tinySynth.midi._GEN_0[2] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold111 (.A(\ChiselTop.tinySynth.osc.square.cnt[15] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0423_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold113 (.A(\ChiselTop.tinySynth.osc.square.cnt[28] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0449_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold115 (.A(\ChiselTop.tinySynth.osc.square.cnt[10] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0412_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold117 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[15] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0520_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold119 (.A(\ChiselTop.tinySynth.osc.square.cnt[29] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold120 (.A(\ChiselTop.tinySynth.uart.rx.bitsReg[1] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold121 (.A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[6] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold122 (.A(\ChiselTop.tinySynth.pwm.counter[5] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0465_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold124 (.A(\ChiselTop.tinySynth.pwm.counter[4] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0464_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold126 (.A(\ChiselTop.tinySynth.osc.square.cnt[21] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0436_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold128 (.A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[3] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0546_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold130 (.A(\ChiselTop.tinySynth.osc.square.cnt[4] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0399_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold132 (.A(\ChiselTop.tinySynth.osc.square.cnt[23] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0440_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0049_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold135 (.A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[2] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold136 (.A(\ChiselTop.tinySynth.midi.regState[0] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0003_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold138 (.A(\ChiselTop.tinySynth.osc.square.cnt[11] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0414_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold140 (.A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[1] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold141 (.A(\ChiselTop.tinySynth.osc.square.cnt[24] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0442_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold143 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[1] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold144 (.A(\ChiselTop.tinySynth.osc.square.cnt[14] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold145 (.A(\ChiselTop.tinySynth.uart.rx.bitsReg[2] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold146 (.A(\ChiselTop.tinySynth.midi.io_midiOut_bits_note[5] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold147 (.A(\ChiselTop.tinySynth.osc.square.cnt[8] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold148 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[8] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0511_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0008_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0432_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold152 (.A(\ChiselTop.tinySynth.pwm.counter[3] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0461_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold154 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[2] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold155 (.A(\ChiselTop.tinySynth.osc.square.cnt[20] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0434_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold157 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[4] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold158 (.A(\ChiselTop.tinySynth.osc.square.cnt[18] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold159 (.A(\ChiselTop.tinySynth.osc.square.cnt[22] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold160 (.A(\ChiselTop.tinySynth.osc.square.cnt[2] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0394_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold162 (.A(\ChiselTop.tinySynth.uart.rx.cntReg[5] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0506_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold164 (.A(\ChiselTop.tinySynth.midi.regState[3] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0001_),
    .X(net315));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_fill_2 FILLER_4_231 ();
 sg13g2_fill_2 FILLER_4_237 ();
 sg13g2_decap_8 FILLER_4_247 ();
 sg13g2_decap_4 FILLER_4_254 ();
 sg13g2_fill_2 FILLER_4_258 ();
 sg13g2_decap_8 FILLER_4_265 ();
 sg13g2_decap_8 FILLER_4_272 ();
 sg13g2_decap_8 FILLER_4_279 ();
 sg13g2_decap_8 FILLER_4_286 ();
 sg13g2_decap_8 FILLER_4_293 ();
 sg13g2_decap_8 FILLER_4_300 ();
 sg13g2_decap_8 FILLER_4_307 ();
 sg13g2_decap_8 FILLER_4_314 ();
 sg13g2_decap_8 FILLER_4_321 ();
 sg13g2_decap_8 FILLER_4_328 ();
 sg13g2_decap_8 FILLER_4_335 ();
 sg13g2_decap_8 FILLER_4_342 ();
 sg13g2_decap_8 FILLER_4_349 ();
 sg13g2_decap_8 FILLER_4_356 ();
 sg13g2_decap_8 FILLER_4_363 ();
 sg13g2_decap_8 FILLER_4_370 ();
 sg13g2_decap_8 FILLER_4_377 ();
 sg13g2_decap_8 FILLER_4_384 ();
 sg13g2_decap_8 FILLER_4_391 ();
 sg13g2_decap_8 FILLER_4_398 ();
 sg13g2_decap_4 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_4 FILLER_5_133 ();
 sg13g2_fill_2 FILLER_5_137 ();
 sg13g2_fill_1 FILLER_5_157 ();
 sg13g2_decap_4 FILLER_5_173 ();
 sg13g2_fill_1 FILLER_5_177 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_4 FILLER_5_203 ();
 sg13g2_fill_1 FILLER_5_207 ();
 sg13g2_fill_2 FILLER_5_260 ();
 sg13g2_decap_8 FILLER_5_276 ();
 sg13g2_decap_8 FILLER_5_283 ();
 sg13g2_decap_8 FILLER_5_290 ();
 sg13g2_decap_8 FILLER_5_297 ();
 sg13g2_decap_8 FILLER_5_304 ();
 sg13g2_decap_8 FILLER_5_311 ();
 sg13g2_decap_8 FILLER_5_318 ();
 sg13g2_decap_8 FILLER_5_325 ();
 sg13g2_decap_8 FILLER_5_332 ();
 sg13g2_decap_8 FILLER_5_339 ();
 sg13g2_decap_8 FILLER_5_346 ();
 sg13g2_decap_8 FILLER_5_353 ();
 sg13g2_decap_8 FILLER_5_360 ();
 sg13g2_decap_8 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_374 ();
 sg13g2_decap_8 FILLER_5_381 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_4 FILLER_6_126 ();
 sg13g2_fill_1 FILLER_6_130 ();
 sg13g2_decap_8 FILLER_6_191 ();
 sg13g2_fill_2 FILLER_6_198 ();
 sg13g2_fill_1 FILLER_6_242 ();
 sg13g2_fill_2 FILLER_6_262 ();
 sg13g2_decap_8 FILLER_6_290 ();
 sg13g2_decap_8 FILLER_6_297 ();
 sg13g2_decap_4 FILLER_6_304 ();
 sg13g2_fill_1 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_313 ();
 sg13g2_decap_4 FILLER_6_320 ();
 sg13g2_fill_2 FILLER_6_329 ();
 sg13g2_fill_2 FILLER_6_335 ();
 sg13g2_decap_8 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_356 ();
 sg13g2_decap_8 FILLER_6_363 ();
 sg13g2_decap_8 FILLER_6_370 ();
 sg13g2_decap_8 FILLER_6_377 ();
 sg13g2_decap_8 FILLER_6_384 ();
 sg13g2_decap_8 FILLER_6_391 ();
 sg13g2_decap_8 FILLER_6_398 ();
 sg13g2_decap_4 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_fill_2 FILLER_7_119 ();
 sg13g2_fill_1 FILLER_7_152 ();
 sg13g2_fill_2 FILLER_7_255 ();
 sg13g2_fill_1 FILLER_7_262 ();
 sg13g2_fill_1 FILLER_7_297 ();
 sg13g2_decap_8 FILLER_7_358 ();
 sg13g2_decap_8 FILLER_7_365 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_4 FILLER_8_119 ();
 sg13g2_fill_1 FILLER_8_123 ();
 sg13g2_fill_2 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_186 ();
 sg13g2_decap_4 FILLER_8_193 ();
 sg13g2_fill_1 FILLER_8_197 ();
 sg13g2_fill_1 FILLER_8_257 ();
 sg13g2_fill_2 FILLER_8_284 ();
 sg13g2_decap_4 FILLER_8_294 ();
 sg13g2_fill_1 FILLER_8_305 ();
 sg13g2_fill_2 FILLER_8_327 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_fill_2 FILLER_9_160 ();
 sg13g2_fill_1 FILLER_9_241 ();
 sg13g2_fill_2 FILLER_9_251 ();
 sg13g2_fill_2 FILLER_9_309 ();
 sg13g2_fill_1 FILLER_9_320 ();
 sg13g2_fill_1 FILLER_9_341 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_fill_2 FILLER_10_119 ();
 sg13g2_fill_1 FILLER_10_121 ();
 sg13g2_fill_1 FILLER_10_171 ();
 sg13g2_fill_2 FILLER_10_211 ();
 sg13g2_fill_1 FILLER_10_253 ();
 sg13g2_fill_1 FILLER_10_290 ();
 sg13g2_fill_1 FILLER_10_308 ();
 sg13g2_fill_2 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_390 ();
 sg13g2_decap_8 FILLER_10_397 ();
 sg13g2_decap_4 FILLER_10_404 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_4 FILLER_11_119 ();
 sg13g2_fill_2 FILLER_11_123 ();
 sg13g2_fill_2 FILLER_11_207 ();
 sg13g2_fill_1 FILLER_11_209 ();
 sg13g2_fill_2 FILLER_11_215 ();
 sg13g2_fill_1 FILLER_11_226 ();
 sg13g2_fill_2 FILLER_11_331 ();
 sg13g2_fill_2 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_384 ();
 sg13g2_decap_8 FILLER_11_391 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_4 FILLER_12_119 ();
 sg13g2_decap_4 FILLER_12_198 ();
 sg13g2_fill_1 FILLER_12_258 ();
 sg13g2_fill_2 FILLER_12_327 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_4 FILLER_13_112 ();
 sg13g2_fill_2 FILLER_13_116 ();
 sg13g2_fill_1 FILLER_13_153 ();
 sg13g2_fill_2 FILLER_13_180 ();
 sg13g2_fill_2 FILLER_13_217 ();
 sg13g2_fill_2 FILLER_13_229 ();
 sg13g2_fill_2 FILLER_13_236 ();
 sg13g2_decap_4 FILLER_13_245 ();
 sg13g2_fill_1 FILLER_13_249 ();
 sg13g2_fill_1 FILLER_13_276 ();
 sg13g2_fill_1 FILLER_13_335 ();
 sg13g2_fill_2 FILLER_13_365 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_fill_2 FILLER_14_126 ();
 sg13g2_fill_1 FILLER_14_128 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_4 FILLER_14_140 ();
 sg13g2_fill_1 FILLER_14_144 ();
 sg13g2_fill_2 FILLER_14_171 ();
 sg13g2_fill_1 FILLER_14_173 ();
 sg13g2_fill_1 FILLER_14_197 ();
 sg13g2_decap_4 FILLER_14_215 ();
 sg13g2_fill_2 FILLER_14_219 ();
 sg13g2_decap_4 FILLER_14_250 ();
 sg13g2_fill_1 FILLER_14_254 ();
 sg13g2_fill_1 FILLER_14_282 ();
 sg13g2_fill_1 FILLER_14_293 ();
 sg13g2_fill_1 FILLER_14_320 ();
 sg13g2_fill_1 FILLER_14_330 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_4 FILLER_15_147 ();
 sg13g2_fill_1 FILLER_15_151 ();
 sg13g2_decap_4 FILLER_15_156 ();
 sg13g2_decap_4 FILLER_15_168 ();
 sg13g2_fill_1 FILLER_15_172 ();
 sg13g2_fill_2 FILLER_15_213 ();
 sg13g2_fill_1 FILLER_15_215 ();
 sg13g2_fill_2 FILLER_15_242 ();
 sg13g2_fill_2 FILLER_15_283 ();
 sg13g2_decap_4 FILLER_15_300 ();
 sg13g2_fill_1 FILLER_15_304 ();
 sg13g2_fill_1 FILLER_15_309 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_4 FILLER_16_161 ();
 sg13g2_fill_1 FILLER_16_165 ();
 sg13g2_decap_8 FILLER_16_268 ();
 sg13g2_decap_4 FILLER_16_314 ();
 sg13g2_fill_2 FILLER_16_318 ();
 sg13g2_fill_1 FILLER_16_329 ();
 sg13g2_fill_2 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_fill_2 FILLER_17_154 ();
 sg13g2_fill_1 FILLER_17_156 ();
 sg13g2_fill_1 FILLER_17_187 ();
 sg13g2_fill_2 FILLER_17_199 ();
 sg13g2_fill_2 FILLER_17_229 ();
 sg13g2_fill_1 FILLER_17_240 ();
 sg13g2_decap_4 FILLER_17_327 ();
 sg13g2_fill_2 FILLER_17_331 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_fill_2 FILLER_18_147 ();
 sg13g2_fill_1 FILLER_18_203 ();
 sg13g2_fill_1 FILLER_18_223 ();
 sg13g2_fill_2 FILLER_18_233 ();
 sg13g2_fill_1 FILLER_18_287 ();
 sg13g2_fill_2 FILLER_18_317 ();
 sg13g2_fill_1 FILLER_18_319 ();
 sg13g2_decap_4 FILLER_18_339 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_fill_2 FILLER_19_154 ();
 sg13g2_fill_1 FILLER_19_156 ();
 sg13g2_fill_1 FILLER_19_187 ();
 sg13g2_decap_8 FILLER_19_261 ();
 sg13g2_decap_8 FILLER_19_268 ();
 sg13g2_fill_2 FILLER_19_290 ();
 sg13g2_fill_1 FILLER_19_292 ();
 sg13g2_fill_2 FILLER_19_315 ();
 sg13g2_fill_1 FILLER_19_332 ();
 sg13g2_decap_4 FILLER_19_338 ();
 sg13g2_fill_1 FILLER_19_348 ();
 sg13g2_fill_1 FILLER_19_354 ();
 sg13g2_fill_2 FILLER_19_381 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_fill_1 FILLER_20_161 ();
 sg13g2_fill_1 FILLER_20_201 ();
 sg13g2_fill_2 FILLER_20_223 ();
 sg13g2_fill_1 FILLER_20_225 ();
 sg13g2_fill_1 FILLER_20_243 ();
 sg13g2_fill_2 FILLER_20_291 ();
 sg13g2_decap_4 FILLER_20_301 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_decap_4 FILLER_20_322 ();
 sg13g2_decap_4 FILLER_20_333 ();
 sg13g2_fill_2 FILLER_20_366 ();
 sg13g2_fill_2 FILLER_20_377 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_4 FILLER_21_168 ();
 sg13g2_fill_1 FILLER_21_172 ();
 sg13g2_fill_2 FILLER_21_199 ();
 sg13g2_fill_1 FILLER_21_201 ();
 sg13g2_decap_8 FILLER_21_241 ();
 sg13g2_decap_8 FILLER_21_248 ();
 sg13g2_fill_2 FILLER_21_269 ();
 sg13g2_fill_1 FILLER_21_271 ();
 sg13g2_fill_1 FILLER_21_293 ();
 sg13g2_fill_2 FILLER_21_308 ();
 sg13g2_decap_4 FILLER_21_334 ();
 sg13g2_fill_2 FILLER_21_366 ();
 sg13g2_fill_2 FILLER_21_376 ();
 sg13g2_fill_1 FILLER_21_378 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_4 FILLER_22_175 ();
 sg13g2_fill_1 FILLER_22_179 ();
 sg13g2_fill_2 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_208 ();
 sg13g2_fill_2 FILLER_22_244 ();
 sg13g2_fill_1 FILLER_22_276 ();
 sg13g2_fill_2 FILLER_22_314 ();
 sg13g2_fill_1 FILLER_22_316 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_fill_2 FILLER_22_343 ();
 sg13g2_decap_4 FILLER_22_366 ();
 sg13g2_fill_2 FILLER_22_370 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_fill_1 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_141 ();
 sg13g2_fill_1 FILLER_23_148 ();
 sg13g2_decap_8 FILLER_23_158 ();
 sg13g2_decap_4 FILLER_23_165 ();
 sg13g2_fill_1 FILLER_23_169 ();
 sg13g2_fill_2 FILLER_23_196 ();
 sg13g2_fill_1 FILLER_23_224 ();
 sg13g2_fill_1 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_261 ();
 sg13g2_decap_8 FILLER_23_268 ();
 sg13g2_decap_8 FILLER_23_275 ();
 sg13g2_fill_1 FILLER_23_282 ();
 sg13g2_fill_2 FILLER_23_291 ();
 sg13g2_fill_1 FILLER_23_293 ();
 sg13g2_fill_2 FILLER_23_300 ();
 sg13g2_fill_1 FILLER_23_302 ();
 sg13g2_fill_1 FILLER_23_351 ();
 sg13g2_fill_1 FILLER_23_356 ();
 sg13g2_fill_1 FILLER_23_362 ();
 sg13g2_decap_4 FILLER_23_373 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_4 FILLER_24_119 ();
 sg13g2_fill_2 FILLER_24_123 ();
 sg13g2_fill_2 FILLER_24_151 ();
 sg13g2_fill_1 FILLER_24_153 ();
 sg13g2_decap_8 FILLER_24_163 ();
 sg13g2_fill_1 FILLER_24_170 ();
 sg13g2_fill_2 FILLER_24_223 ();
 sg13g2_fill_1 FILLER_24_225 ();
 sg13g2_fill_2 FILLER_24_264 ();
 sg13g2_fill_2 FILLER_24_275 ();
 sg13g2_fill_1 FILLER_24_277 ();
 sg13g2_decap_4 FILLER_24_282 ();
 sg13g2_fill_1 FILLER_24_286 ();
 sg13g2_decap_8 FILLER_24_293 ();
 sg13g2_decap_4 FILLER_24_300 ();
 sg13g2_fill_2 FILLER_24_304 ();
 sg13g2_decap_4 FILLER_24_324 ();
 sg13g2_fill_2 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_362 ();
 sg13g2_decap_4 FILLER_24_369 ();
 sg13g2_fill_2 FILLER_24_373 ();
 sg13g2_fill_1 FILLER_24_383 ();
 sg13g2_decap_4 FILLER_24_389 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_4 FILLER_25_105 ();
 sg13g2_fill_2 FILLER_25_109 ();
 sg13g2_fill_2 FILLER_25_129 ();
 sg13g2_fill_1 FILLER_25_206 ();
 sg13g2_fill_2 FILLER_25_264 ();
 sg13g2_fill_2 FILLER_25_271 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_fill_1 FILLER_25_332 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_4 FILLER_26_98 ();
 sg13g2_fill_2 FILLER_26_102 ();
 sg13g2_fill_1 FILLER_26_130 ();
 sg13g2_fill_1 FILLER_26_159 ();
 sg13g2_fill_1 FILLER_26_164 ();
 sg13g2_decap_4 FILLER_26_178 ();
 sg13g2_fill_2 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_207 ();
 sg13g2_fill_2 FILLER_26_217 ();
 sg13g2_fill_1 FILLER_26_236 ();
 sg13g2_fill_1 FILLER_26_251 ();
 sg13g2_fill_2 FILLER_26_265 ();
 sg13g2_decap_8 FILLER_26_272 ();
 sg13g2_decap_4 FILLER_26_291 ();
 sg13g2_fill_2 FILLER_26_295 ();
 sg13g2_fill_2 FILLER_26_312 ();
 sg13g2_fill_2 FILLER_26_320 ();
 sg13g2_decap_4 FILLER_26_327 ();
 sg13g2_fill_2 FILLER_26_331 ();
 sg13g2_decap_4 FILLER_26_343 ();
 sg13g2_fill_2 FILLER_26_347 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_4 FILLER_27_91 ();
 sg13g2_fill_1 FILLER_27_144 ();
 sg13g2_decap_4 FILLER_27_187 ();
 sg13g2_fill_2 FILLER_27_191 ();
 sg13g2_fill_1 FILLER_27_246 ();
 sg13g2_decap_4 FILLER_27_268 ();
 sg13g2_decap_4 FILLER_27_339 ();
 sg13g2_fill_1 FILLER_27_343 ();
 sg13g2_fill_1 FILLER_27_356 ();
 sg13g2_fill_2 FILLER_27_367 ();
 sg13g2_decap_4 FILLER_27_378 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_fill_2 FILLER_28_170 ();
 sg13g2_fill_2 FILLER_28_185 ();
 sg13g2_fill_1 FILLER_28_213 ();
 sg13g2_fill_1 FILLER_28_223 ();
 sg13g2_fill_2 FILLER_28_245 ();
 sg13g2_fill_1 FILLER_28_261 ();
 sg13g2_fill_1 FILLER_28_284 ();
 sg13g2_decap_8 FILLER_28_292 ();
 sg13g2_decap_8 FILLER_28_299 ();
 sg13g2_decap_8 FILLER_28_306 ();
 sg13g2_fill_2 FILLER_28_313 ();
 sg13g2_fill_2 FILLER_28_351 ();
 sg13g2_fill_1 FILLER_28_353 ();
 sg13g2_fill_2 FILLER_28_371 ();
 sg13g2_fill_1 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_fill_1 FILLER_29_180 ();
 sg13g2_decap_4 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_197 ();
 sg13g2_decap_4 FILLER_29_202 ();
 sg13g2_fill_2 FILLER_29_206 ();
 sg13g2_decap_4 FILLER_29_220 ();
 sg13g2_decap_8 FILLER_29_227 ();
 sg13g2_decap_8 FILLER_29_234 ();
 sg13g2_fill_1 FILLER_29_241 ();
 sg13g2_fill_2 FILLER_29_251 ();
 sg13g2_fill_1 FILLER_29_253 ();
 sg13g2_decap_4 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_272 ();
 sg13g2_decap_4 FILLER_29_291 ();
 sg13g2_decap_8 FILLER_29_328 ();
 sg13g2_fill_2 FILLER_29_362 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_91 ();
 sg13g2_fill_1 FILLER_30_150 ();
 sg13g2_fill_1 FILLER_30_161 ();
 sg13g2_fill_1 FILLER_30_191 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_4 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_228 ();
 sg13g2_fill_2 FILLER_30_235 ();
 sg13g2_fill_1 FILLER_30_237 ();
 sg13g2_fill_1 FILLER_30_246 ();
 sg13g2_fill_2 FILLER_30_259 ();
 sg13g2_fill_1 FILLER_30_261 ();
 sg13g2_fill_2 FILLER_30_271 ();
 sg13g2_fill_1 FILLER_30_278 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_fill_2 FILLER_30_294 ();
 sg13g2_fill_1 FILLER_30_313 ();
 sg13g2_decap_4 FILLER_30_327 ();
 sg13g2_decap_4 FILLER_30_335 ();
 sg13g2_fill_2 FILLER_30_339 ();
 sg13g2_fill_2 FILLER_30_360 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_fill_1 FILLER_31_98 ();
 sg13g2_fill_2 FILLER_31_166 ();
 sg13g2_fill_2 FILLER_31_177 ();
 sg13g2_fill_1 FILLER_31_179 ();
 sg13g2_fill_2 FILLER_31_192 ();
 sg13g2_decap_4 FILLER_31_232 ();
 sg13g2_fill_2 FILLER_31_267 ();
 sg13g2_decap_8 FILLER_31_277 ();
 sg13g2_fill_2 FILLER_31_284 ();
 sg13g2_fill_1 FILLER_31_286 ();
 sg13g2_decap_4 FILLER_31_297 ();
 sg13g2_fill_1 FILLER_31_307 ();
 sg13g2_decap_8 FILLER_31_313 ();
 sg13g2_fill_2 FILLER_31_337 ();
 sg13g2_fill_1 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_348 ();
 sg13g2_fill_2 FILLER_31_369 ();
 sg13g2_fill_1 FILLER_31_371 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_4 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_128 ();
 sg13g2_fill_1 FILLER_32_181 ();
 sg13g2_decap_8 FILLER_32_198 ();
 sg13g2_fill_2 FILLER_32_205 ();
 sg13g2_fill_1 FILLER_32_236 ();
 sg13g2_fill_1 FILLER_32_242 ();
 sg13g2_fill_1 FILLER_32_246 ();
 sg13g2_fill_1 FILLER_32_251 ();
 sg13g2_fill_1 FILLER_32_285 ();
 sg13g2_fill_2 FILLER_32_312 ();
 sg13g2_fill_2 FILLER_32_356 ();
 sg13g2_fill_1 FILLER_32_358 ();
 sg13g2_fill_2 FILLER_32_364 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_fill_2 FILLER_33_116 ();
 sg13g2_fill_1 FILLER_33_127 ();
 sg13g2_fill_2 FILLER_33_141 ();
 sg13g2_fill_2 FILLER_33_147 ();
 sg13g2_fill_2 FILLER_33_158 ();
 sg13g2_fill_2 FILLER_33_193 ();
 sg13g2_fill_2 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_263 ();
 sg13g2_decap_8 FILLER_33_277 ();
 sg13g2_decap_8 FILLER_33_284 ();
 sg13g2_fill_2 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_308 ();
 sg13g2_fill_1 FILLER_33_318 ();
 sg13g2_fill_1 FILLER_33_332 ();
 sg13g2_fill_2 FILLER_33_351 ();
 sg13g2_fill_1 FILLER_33_353 ();
 sg13g2_fill_2 FILLER_33_378 ();
 sg13g2_fill_1 FILLER_33_380 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_fill_2 FILLER_34_133 ();
 sg13g2_fill_1 FILLER_34_135 ();
 sg13g2_fill_2 FILLER_34_140 ();
 sg13g2_fill_2 FILLER_34_146 ();
 sg13g2_fill_1 FILLER_34_148 ();
 sg13g2_decap_8 FILLER_34_153 ();
 sg13g2_fill_2 FILLER_34_160 ();
 sg13g2_decap_4 FILLER_34_197 ();
 sg13g2_fill_1 FILLER_34_201 ();
 sg13g2_decap_8 FILLER_34_270 ();
 sg13g2_decap_8 FILLER_34_290 ();
 sg13g2_fill_2 FILLER_34_318 ();
 sg13g2_fill_1 FILLER_34_320 ();
 sg13g2_decap_8 FILLER_34_325 ();
 sg13g2_fill_2 FILLER_34_355 ();
 sg13g2_fill_2 FILLER_34_366 ();
 sg13g2_fill_1 FILLER_34_368 ();
 sg13g2_fill_2 FILLER_34_378 ();
 sg13g2_fill_1 FILLER_34_380 ();
 sg13g2_decap_4 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_4 FILLER_35_182 ();
 sg13g2_fill_1 FILLER_35_186 ();
 sg13g2_decap_4 FILLER_35_190 ();
 sg13g2_fill_2 FILLER_35_246 ();
 sg13g2_fill_2 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_302 ();
 sg13g2_fill_1 FILLER_35_306 ();
 sg13g2_fill_2 FILLER_35_328 ();
 sg13g2_decap_8 FILLER_35_395 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_fill_2 FILLER_36_210 ();
 sg13g2_fill_1 FILLER_36_212 ();
 sg13g2_decap_4 FILLER_36_222 ();
 sg13g2_fill_2 FILLER_36_226 ();
 sg13g2_decap_4 FILLER_36_272 ();
 sg13g2_fill_2 FILLER_36_280 ();
 sg13g2_fill_1 FILLER_36_282 ();
 sg13g2_fill_2 FILLER_36_290 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_fill_2 FILLER_36_308 ();
 sg13g2_fill_1 FILLER_36_310 ();
 sg13g2_decap_4 FILLER_36_337 ();
 sg13g2_decap_8 FILLER_36_345 ();
 sg13g2_fill_2 FILLER_36_352 ();
 sg13g2_fill_1 FILLER_36_354 ();
 sg13g2_fill_2 FILLER_36_363 ();
 sg13g2_fill_2 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_384 ();
 sg13g2_decap_8 FILLER_36_391 ();
 sg13g2_decap_8 FILLER_36_398 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_fill_1 FILLER_37_231 ();
 sg13g2_fill_2 FILLER_37_236 ();
 sg13g2_fill_1 FILLER_37_238 ();
 sg13g2_decap_4 FILLER_37_243 ();
 sg13g2_fill_1 FILLER_37_247 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_4 FILLER_37_315 ();
 sg13g2_fill_1 FILLER_37_319 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_decap_4 FILLER_38_220 ();
 sg13g2_decap_4 FILLER_38_228 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_decap_8 FILLER_38_257 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_decap_8 FILLER_38_278 ();
 sg13g2_decap_8 FILLER_38_285 ();
 sg13g2_decap_8 FILLER_38_292 ();
 sg13g2_decap_8 FILLER_38_299 ();
 sg13g2_decap_8 FILLER_38_306 ();
 sg13g2_decap_8 FILLER_38_313 ();
 sg13g2_decap_8 FILLER_38_320 ();
 sg13g2_decap_8 FILLER_38_327 ();
 sg13g2_decap_8 FILLER_38_334 ();
 sg13g2_decap_8 FILLER_38_341 ();
 sg13g2_decap_8 FILLER_38_348 ();
 sg13g2_decap_8 FILLER_38_355 ();
 sg13g2_decap_4 FILLER_38_362 ();
 sg13g2_fill_2 FILLER_38_366 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
 assign uo_out[1] = net18;
 assign uo_out[2] = net19;
 assign uo_out[3] = net20;
 assign uo_out[4] = net21;
 assign uo_out[5] = net22;
 assign uo_out[6] = net23;
 assign uo_out[7] = net24;
endmodule

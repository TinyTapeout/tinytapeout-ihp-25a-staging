module tt_um_tt08_wirecube (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire clk_regs;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire hsync;
 wire rst_n_sync;
 wire net11;
 wire net12;
 wire net73;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire vsync;
 wire \wirecube_top_inst.any_line_set ;
 wire \wirecube_top_inst.any_line_set2 ;
 wire \wirecube_top_inst.counter_h[0] ;
 wire \wirecube_top_inst.counter_h[10] ;
 wire \wirecube_top_inst.counter_h[1] ;
 wire \wirecube_top_inst.counter_h[2] ;
 wire \wirecube_top_inst.counter_h[3] ;
 wire \wirecube_top_inst.counter_h[4] ;
 wire \wirecube_top_inst.counter_h[5] ;
 wire \wirecube_top_inst.counter_h[6] ;
 wire \wirecube_top_inst.counter_h[7] ;
 wire \wirecube_top_inst.counter_h[8] ;
 wire \wirecube_top_inst.counter_h[9] ;
 wire \wirecube_top_inst.counter_v[0] ;
 wire \wirecube_top_inst.counter_v[10] ;
 wire \wirecube_top_inst.counter_v[1] ;
 wire \wirecube_top_inst.counter_v[2] ;
 wire \wirecube_top_inst.counter_v[3] ;
 wire \wirecube_top_inst.counter_v[4] ;
 wire \wirecube_top_inst.counter_v[5] ;
 wire \wirecube_top_inst.counter_v[6] ;
 wire \wirecube_top_inst.counter_v[7] ;
 wire \wirecube_top_inst.counter_v[8] ;
 wire \wirecube_top_inst.counter_v[9] ;
 wire \wirecube_top_inst.cur_state_background[0] ;
 wire \wirecube_top_inst.cur_state_background[1] ;
 wire \wirecube_top_inst.cur_state_background[2] ;
 wire \wirecube_top_inst.cur_state_background[3] ;
 wire \wirecube_top_inst.delay_inst_hsync.in_i ;
 wire \wirecube_top_inst.delay_inst_hsync.pipe[0] ;
 wire \wirecube_top_inst.delay_inst_vsync.in_i ;
 wire \wirecube_top_inst.delay_inst_vsync.pipe[0] ;
 wire \wirecube_top_inst.edge_function_inst.absolute[0] ;
 wire \wirecube_top_inst.edge_function_inst.absolute[10] ;
 wire \wirecube_top_inst.edge_function_inst.absolute[11] ;
 wire \wirecube_top_inst.edge_function_inst.absolute[12] ;
 wire \wirecube_top_inst.edge_function_inst.absolute[13] ;
 wire \wirecube_top_inst.edge_function_inst.absolute[1] ;
 wire \wirecube_top_inst.edge_function_inst.absolute[2] ;
 wire \wirecube_top_inst.edge_function_inst.absolute[3] ;
 wire \wirecube_top_inst.edge_function_inst.absolute[4] ;
 wire \wirecube_top_inst.edge_function_inst.absolute[5] ;
 wire \wirecube_top_inst.edge_function_inst.absolute[6] ;
 wire \wirecube_top_inst.edge_function_inst.absolute[7] ;
 wire \wirecube_top_inst.edge_function_inst.absolute[8] ;
 wire \wirecube_top_inst.edge_function_inst.absolute[9] ;
 wire \wirecube_top_inst.edge_function_inst.pixel_x_i[0] ;
 wire \wirecube_top_inst.edge_function_inst.pixel_x_i[1] ;
 wire \wirecube_top_inst.edge_function_inst.pixel_x_i[2] ;
 wire \wirecube_top_inst.edge_function_inst.pixel_x_i[3] ;
 wire \wirecube_top_inst.edge_function_inst.pixel_x_i[4] ;
 wire \wirecube_top_inst.edge_function_inst.pixel_x_i[5] ;
 wire \wirecube_top_inst.edge_function_inst.pixel_x_i[6] ;
 wire \wirecube_top_inst.edge_function_inst.pixel_y_i[0] ;
 wire \wirecube_top_inst.edge_function_inst.pixel_y_i[1] ;
 wire \wirecube_top_inst.edge_function_inst.pixel_y_i[2] ;
 wire \wirecube_top_inst.edge_function_inst.pixel_y_i[3] ;
 wire \wirecube_top_inst.edge_function_inst.pixel_y_i[4] ;
 wire \wirecube_top_inst.edge_function_inst.pixel_y_i[5] ;
 wire \wirecube_top_inst.edge_function_inst.pixel_y_i[6] ;
 wire \wirecube_top_inst.edge_function_inst.term0[0] ;
 wire \wirecube_top_inst.edge_function_inst.term0[1] ;
 wire \wirecube_top_inst.edge_function_inst.term0[2] ;
 wire \wirecube_top_inst.edge_function_inst.term0[3] ;
 wire \wirecube_top_inst.edge_function_inst.term0[4] ;
 wire \wirecube_top_inst.edge_function_inst.term0[5] ;
 wire \wirecube_top_inst.edge_function_inst.term0[6] ;
 wire \wirecube_top_inst.edge_function_inst.term1[0] ;
 wire \wirecube_top_inst.edge_function_inst.term1[1] ;
 wire \wirecube_top_inst.edge_function_inst.term1[2] ;
 wire \wirecube_top_inst.edge_function_inst.term1[3] ;
 wire \wirecube_top_inst.edge_function_inst.term1[4] ;
 wire \wirecube_top_inst.edge_function_inst.term1[5] ;
 wire \wirecube_top_inst.edge_function_inst.term1[6] ;
 wire \wirecube_top_inst.edge_function_inst.term2[0] ;
 wire \wirecube_top_inst.edge_function_inst.term2[1] ;
 wire \wirecube_top_inst.edge_function_inst.term2[2] ;
 wire \wirecube_top_inst.edge_function_inst.term2[3] ;
 wire \wirecube_top_inst.edge_function_inst.term2[4] ;
 wire \wirecube_top_inst.edge_function_inst.term2[5] ;
 wire \wirecube_top_inst.edge_function_inst.term2[6] ;
 wire \wirecube_top_inst.edge_function_inst.term3[0] ;
 wire \wirecube_top_inst.edge_function_inst.term3[1] ;
 wire \wirecube_top_inst.edge_function_inst.term3[2] ;
 wire \wirecube_top_inst.edge_function_inst.term3[3] ;
 wire \wirecube_top_inst.edge_function_inst.term3[4] ;
 wire \wirecube_top_inst.edge_function_inst.term3[5] ;
 wire \wirecube_top_inst.edge_function_inst.term3[6] ;
 wire \wirecube_top_inst.edge_function_inst.visible ;
 wire \wirecube_top_inst.edge_function_inst.visible_2 ;
 wire \wirecube_top_inst.final_pixel ;
 wire \wirecube_top_inst.final_pixel2 ;
 wire \wirecube_top_inst.frame_cnt[0] ;
 wire \wirecube_top_inst.frame_cnt[12] ;
 wire \wirecube_top_inst.frame_cnt[1] ;
 wire \wirecube_top_inst.frame_cnt[2] ;
 wire \wirecube_top_inst.frame_cnt[3] ;
 wire \wirecube_top_inst.frame_cnt[4] ;
 wire \wirecube_top_inst.frame_cnt[5] ;
 wire \wirecube_top_inst.frame_cnt[6] ;
 wire \wirecube_top_inst.frame_cnt[7] ;
 wire \wirecube_top_inst.line_rom_inst.line_i[0] ;
 wire \wirecube_top_inst.line_rom_inst.line_i[1] ;
 wire \wirecube_top_inst.line_rom_inst.line_i[2] ;
 wire \wirecube_top_inst.line_rom_inst.line_i[3] ;
 wire \wirecube_top_inst.linecounter_h[0] ;
 wire \wirecube_top_inst.linecounter_h[1] ;
 wire \wirecube_top_inst.linecounter_h[2] ;
 wire \wirecube_top_inst.linecounter_h[3] ;
 wire \wirecube_top_inst.subcounter_v[0] ;
 wire \wirecube_top_inst.subcounter_v[1] ;
 wire \wirecube_top_inst.subcounter_v[2] ;
 wire \wirecube_top_inst.timing_hor.counter[11] ;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire delaynet_0_clk;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;

 sg13g2_inv_2 _2677_ (.Y(_1793_),
    .A(net691));
 sg13g2_inv_2 _2678_ (.Y(_1804_),
    .A(net692));
 sg13g2_inv_2 _2679_ (.Y(_1813_),
    .A(net685));
 sg13g2_inv_1 _2680_ (.Y(_1821_),
    .A(net684));
 sg13g2_inv_1 _2681_ (.Y(_1829_),
    .A(net9));
 sg13g2_inv_1 _2682_ (.Y(_1834_),
    .A(_0069_));
 sg13g2_inv_1 _2683_ (.Y(_1835_),
    .A(_0070_));
 sg13g2_inv_1 _2684_ (.Y(_1836_),
    .A(_0072_));
 sg13g2_inv_1 _2685_ (.Y(_1837_),
    .A(net160));
 sg13g2_inv_1 _2686_ (.Y(_1838_),
    .A(net700));
 sg13g2_inv_1 _2687_ (.Y(_1839_),
    .A(net175));
 sg13g2_inv_1 _2688_ (.Y(_1840_),
    .A(\wirecube_top_inst.counter_v[8] ));
 sg13g2_inv_1 _2689_ (.Y(_1841_),
    .A(\wirecube_top_inst.subcounter_v[0] ));
 sg13g2_inv_1 _2690_ (.Y(_1842_),
    .A(\wirecube_top_inst.edge_function_inst.pixel_y_i[5] ));
 sg13g2_inv_1 _2691_ (.Y(_1843_),
    .A(\wirecube_top_inst.edge_function_inst.pixel_y_i[3] ));
 sg13g2_inv_1 _2692_ (.Y(_1844_),
    .A(\wirecube_top_inst.edge_function_inst.pixel_y_i[2] ));
 sg13g2_inv_2 _2693_ (.Y(_1845_),
    .A(\wirecube_top_inst.edge_function_inst.pixel_y_i[1] ));
 sg13g2_inv_1 _2694_ (.Y(_1846_),
    .A(\wirecube_top_inst.edge_function_inst.pixel_x_i[6] ));
 sg13g2_inv_1 _2695_ (.Y(_1847_),
    .A(\wirecube_top_inst.edge_function_inst.pixel_x_i[4] ));
 sg13g2_inv_2 _2696_ (.Y(_1848_),
    .A(\wirecube_top_inst.edge_function_inst.pixel_x_i[3] ));
 sg13g2_inv_1 _2697_ (.Y(_1849_),
    .A(net681));
 sg13g2_inv_2 _2698_ (.Y(_1850_),
    .A(net168));
 sg13g2_inv_1 _2699_ (.Y(_1851_),
    .A(_0064_));
 sg13g2_inv_1 _2700_ (.Y(_1852_),
    .A(net105));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_nor2b_1 _2702_ (.A(\wirecube_top_inst.timing_hor.counter[11] ),
    .B_N(\wirecube_top_inst.counter_h[10] ),
    .Y(_1853_));
 sg13g2_and2_1 _2703_ (.A(net159),
    .B(net113),
    .X(_1854_));
 sg13g2_nand2_1 _2704_ (.Y(_1855_),
    .A(net202),
    .B(net113));
 sg13g2_and3_1 _2705_ (.X(_1856_),
    .A(\wirecube_top_inst.counter_h[3] ),
    .B(\wirecube_top_inst.counter_h[2] ),
    .C(_1854_));
 sg13g2_and2_1 _2706_ (.A(net143),
    .B(_1856_),
    .X(_1857_));
 sg13g2_and3_2 _2707_ (.X(_1858_),
    .A(\wirecube_top_inst.counter_h[6] ),
    .B(\wirecube_top_inst.counter_h[5] ),
    .C(_1857_));
 sg13g2_a21oi_1 _2708_ (.A1(\wirecube_top_inst.counter_h[7] ),
    .A2(_1858_),
    .Y(_1859_),
    .B1(net119));
 sg13g2_nand2b_1 _2709_ (.Y(_1860_),
    .B(_1859_),
    .A_N(\wirecube_top_inst.counter_h[9] ));
 sg13g2_and2_1 _2710_ (.A(_1853_),
    .B(_1860_),
    .X(_1861_));
 sg13g2_nand2_1 _2711_ (.Y(_1862_),
    .A(_1853_),
    .B(_1860_));
 sg13g2_and4_1 _2712_ (.A(net119),
    .B(net141),
    .C(net128),
    .D(\wirecube_top_inst.counter_h[7] ),
    .X(_1863_));
 sg13g2_nand2_1 _2713_ (.Y(_1864_),
    .A(_1858_),
    .B(_1863_));
 sg13g2_xnor2_1 _2714_ (.Y(_1865_),
    .A(net125),
    .B(_1864_));
 sg13g2_nor2_1 _2715_ (.A(net627),
    .B(_1865_),
    .Y(_0107_));
 sg13g2_and3_1 _2716_ (.X(_1866_),
    .A(net119),
    .B(net172),
    .C(_1858_));
 sg13g2_a21o_1 _2717_ (.A2(_1866_),
    .A1(\wirecube_top_inst.counter_h[9] ),
    .B1(net128),
    .X(_1867_));
 sg13g2_a21oi_1 _2718_ (.A1(_1864_),
    .A2(net129),
    .Y(_0106_),
    .B1(net627));
 sg13g2_xor2_1 _2719_ (.B(_1866_),
    .A(net135),
    .X(_1868_));
 sg13g2_nor2_1 _2720_ (.A(net627),
    .B(_1868_),
    .Y(_0105_));
 sg13g2_xor2_1 _2721_ (.B(_1858_),
    .A(net163),
    .X(_1869_));
 sg13g2_nor2_1 _2722_ (.A(net627),
    .B(_1869_),
    .Y(_0104_));
 sg13g2_a21oi_1 _2723_ (.A1(\wirecube_top_inst.counter_h[5] ),
    .A2(_1857_),
    .Y(_1870_),
    .B1(net173));
 sg13g2_o21ai_1 _2724_ (.B1(net626),
    .Y(_1871_),
    .A1(_1858_),
    .A2(net174));
 sg13g2_inv_1 _2725_ (.Y(_0103_),
    .A(_1871_));
 sg13g2_nand2_2 _2726_ (.Y(_1872_),
    .A(\wirecube_top_inst.frame_cnt[0] ),
    .B(\wirecube_top_inst.counter_v[0] ));
 sg13g2_or2_1 _2727_ (.X(_1873_),
    .B(\wirecube_top_inst.counter_v[0] ),
    .A(\wirecube_top_inst.frame_cnt[0] ));
 sg13g2_xor2_1 _2728_ (.B(\wirecube_top_inst.counter_v[0] ),
    .A(\wirecube_top_inst.frame_cnt[0] ),
    .X(_1874_));
 sg13g2_nand2_2 _2729_ (.Y(_1875_),
    .A(_1872_),
    .B(_1873_));
 sg13g2_nor3_2 _2730_ (.A(net684),
    .B(\wirecube_top_inst.cur_state_background[3] ),
    .C(_0062_),
    .Y(_1876_));
 sg13g2_or3_2 _2731_ (.A(\wirecube_top_inst.cur_state_background[2] ),
    .B(\wirecube_top_inst.cur_state_background[3] ),
    .C(_0062_),
    .X(_1877_));
 sg13g2_and2_2 _2732_ (.A(net688),
    .B(net686),
    .X(_1878_));
 sg13g2_nand2_2 _2733_ (.Y(_1879_),
    .A(net688),
    .B(net686));
 sg13g2_nor2_2 _2734_ (.A(net687),
    .B(net685),
    .Y(_1880_));
 sg13g2_or2_2 _2735_ (.X(_1881_),
    .B(net685),
    .A(net687));
 sg13g2_nor2_2 _2736_ (.A(net687),
    .B(_1813_),
    .Y(_1882_));
 sg13g2_nand2b_1 _2737_ (.Y(_1883_),
    .B(net685),
    .A_N(net688));
 sg13g2_nor2b_1 _2738_ (.A(net685),
    .B_N(net687),
    .Y(_1884_));
 sg13g2_nand2b_2 _2739_ (.Y(_1885_),
    .B(net687),
    .A_N(net685));
 sg13g2_nor3_1 _2740_ (.A(_1877_),
    .B(_1878_),
    .C(_1880_),
    .Y(_1886_));
 sg13g2_nand2b_1 _2741_ (.Y(_1887_),
    .B(net683),
    .A_N(net684));
 sg13g2_nand3b_1 _2742_ (.B(net683),
    .C(net682),
    .Y(_1888_),
    .A_N(\wirecube_top_inst.cur_state_background[2] ));
 sg13g2_nor2_1 _2743_ (.A(_1879_),
    .B(_1888_),
    .Y(_1889_));
 sg13g2_nand2_2 _2744_ (.Y(_1890_),
    .A(net684),
    .B(net683));
 sg13g2_nor2_2 _2745_ (.A(_0062_),
    .B(_1890_),
    .Y(_1891_));
 sg13g2_nand3b_1 _2746_ (.B(\wirecube_top_inst.cur_state_background[3] ),
    .C(net684),
    .Y(_1892_),
    .A_N(_0062_));
 sg13g2_nor3_1 _2747_ (.A(_1886_),
    .B(_1889_),
    .C(_1891_),
    .Y(_1893_));
 sg13g2_nor2_1 _2748_ (.A(_1883_),
    .B(_1888_),
    .Y(_1894_));
 sg13g2_nand2b_1 _2749_ (.Y(_1895_),
    .B(_1893_),
    .A_N(_1894_));
 sg13g2_nand2b_2 _2750_ (.Y(_1896_),
    .B(net684),
    .A_N(net683));
 sg13g2_nor2_2 _2751_ (.A(_0062_),
    .B(_1896_),
    .Y(_1897_));
 sg13g2_or2_2 _2752_ (.X(_1898_),
    .B(_1896_),
    .A(_0062_));
 sg13g2_nand2_1 _2753_ (.Y(_1899_),
    .A(\wirecube_top_inst.cur_state_background[1] ),
    .B(_1897_));
 sg13g2_nand2b_1 _2754_ (.Y(_1900_),
    .B(_1883_),
    .A_N(_1888_));
 sg13g2_o21ai_1 _2755_ (.B1(_1900_),
    .Y(_1901_),
    .A1(_1879_),
    .A2(_1898_));
 sg13g2_nand2_1 _2756_ (.Y(_1902_),
    .A(_1893_),
    .B(_1901_));
 sg13g2_nor2_1 _2757_ (.A(_1878_),
    .B(_1898_),
    .Y(_1903_));
 sg13g2_nor2_2 _2758_ (.A(net682),
    .B(_1890_),
    .Y(_1904_));
 sg13g2_nand3b_1 _2759_ (.B(net683),
    .C(net684),
    .Y(_1905_),
    .A_N(net682));
 sg13g2_nor2_1 _2760_ (.A(net689),
    .B(net692),
    .Y(_1906_));
 sg13g2_or2_1 _2761_ (.X(_1907_),
    .B(net692),
    .A(net689));
 sg13g2_nor3_2 _2762_ (.A(_1881_),
    .B(_1905_),
    .C(_1907_),
    .Y(_1908_));
 sg13g2_nor2_2 _2763_ (.A(net682),
    .B(_1887_),
    .Y(_1909_));
 sg13g2_nor3_1 _2764_ (.A(_1903_),
    .B(_1908_),
    .C(_1909_),
    .Y(_1910_));
 sg13g2_nor2_1 _2765_ (.A(net683),
    .B(net682),
    .Y(_1911_));
 sg13g2_nor2_1 _2766_ (.A(_1881_),
    .B(_1906_),
    .Y(_1912_));
 sg13g2_a21oi_2 _2767_ (.B1(_1911_),
    .Y(_1913_),
    .A2(_1912_),
    .A1(_1904_));
 sg13g2_nor2_1 _2768_ (.A(_1877_),
    .B(_1879_),
    .Y(_1914_));
 sg13g2_nor3_1 _2769_ (.A(_1874_),
    .B(_1877_),
    .C(_1879_),
    .Y(_1915_));
 sg13g2_o21ai_1 _2770_ (.B1(_1875_),
    .Y(_1916_),
    .A1(_1895_),
    .A2(_1914_));
 sg13g2_and4_1 _2771_ (.A(_1902_),
    .B(_1910_),
    .C(_1913_),
    .D(_1916_),
    .X(_1917_));
 sg13g2_nand4_1 _2772_ (.B(_1910_),
    .C(_1913_),
    .A(_1902_),
    .Y(_1918_),
    .D(_1916_));
 sg13g2_nor3_2 _2773_ (.A(net682),
    .B(_1881_),
    .C(_1887_),
    .Y(_1919_));
 sg13g2_nor2_2 _2774_ (.A(_1885_),
    .B(_1905_),
    .Y(_1920_));
 sg13g2_o21ai_1 _2775_ (.B1(_1906_),
    .Y(_1921_),
    .A1(_1919_),
    .A2(_1920_));
 sg13g2_nor2_1 _2776_ (.A(_1793_),
    .B(_1804_),
    .Y(_1922_));
 sg13g2_nand2_1 _2777_ (.Y(_1923_),
    .A(net689),
    .B(net692));
 sg13g2_a21oi_2 _2778_ (.B1(_1908_),
    .Y(_1924_),
    .A2(_1922_),
    .A1(_1919_));
 sg13g2_nor3_2 _2779_ (.A(net684),
    .B(net683),
    .C(net682),
    .Y(_1925_));
 sg13g2_a22oi_1 _2780_ (.Y(_1926_),
    .B1(_1925_),
    .B2(_1813_),
    .A2(_1920_),
    .A1(_1907_));
 sg13g2_and3_1 _2781_ (.X(_1927_),
    .A(_1921_),
    .B(_1924_),
    .C(_1926_));
 sg13g2_nand3_1 _2782_ (.B(_1924_),
    .C(_1926_),
    .A(_1921_),
    .Y(_1928_));
 sg13g2_nor2_1 _2783_ (.A(_1881_),
    .B(_1892_),
    .Y(_1929_));
 sg13g2_nor2_1 _2784_ (.A(_1877_),
    .B(_1885_),
    .Y(_1930_));
 sg13g2_o21ai_1 _2785_ (.B1(_1874_),
    .Y(_1931_),
    .A1(_1929_),
    .A2(_1930_));
 sg13g2_nor2_2 _2786_ (.A(net682),
    .B(_1896_),
    .Y(_1932_));
 sg13g2_a221oi_1 _2787_ (.B2(_1884_),
    .C1(_1915_),
    .B1(_1932_),
    .A1(_1878_),
    .Y(_1933_),
    .A2(_1909_));
 sg13g2_o21ai_1 _2788_ (.B1(_1880_),
    .Y(_1934_),
    .A1(_1876_),
    .A2(_1932_));
 sg13g2_and3_1 _2789_ (.X(_1935_),
    .A(_1931_),
    .B(_1933_),
    .C(_1934_));
 sg13g2_nand3_1 _2790_ (.B(_1933_),
    .C(_1934_),
    .A(_1931_),
    .Y(_1936_));
 sg13g2_nor3_1 _2791_ (.A(net9),
    .B(_1928_),
    .C(_1936_),
    .Y(_1937_));
 sg13g2_a21oi_2 _2792_ (.B1(_1829_),
    .Y(_1938_),
    .A2(_1935_),
    .A1(_1927_));
 sg13g2_o21ai_1 _2793_ (.B1(net9),
    .Y(_1939_),
    .A1(_1928_),
    .A2(_1936_));
 sg13g2_nand2b_1 _2794_ (.Y(_1940_),
    .B(_1939_),
    .A_N(net644));
 sg13g2_nor2_2 _2795_ (.A(_1793_),
    .B(_1879_),
    .Y(_1941_));
 sg13g2_nand2_1 _2796_ (.Y(_1942_),
    .A(_1904_),
    .B(_1941_));
 sg13g2_nand2_1 _2797_ (.Y(_1943_),
    .A(net690),
    .B(_1882_));
 sg13g2_nand3_1 _2798_ (.B(_1882_),
    .C(_1909_),
    .A(net689),
    .Y(_1944_));
 sg13g2_o21ai_1 _2799_ (.B1(_1882_),
    .Y(_1945_),
    .A1(_1876_),
    .A2(_1932_));
 sg13g2_a21oi_1 _2800_ (.A1(_1885_),
    .A2(_1891_),
    .Y(_1946_),
    .B1(_1894_));
 sg13g2_nor2_1 _2801_ (.A(_1874_),
    .B(_1946_),
    .Y(_1947_));
 sg13g2_nand2_1 _2802_ (.Y(_1948_),
    .A(_1884_),
    .B(_1891_));
 sg13g2_nor2_2 _2803_ (.A(net689),
    .B(_1883_),
    .Y(_1949_));
 sg13g2_nand2_1 _2804_ (.Y(_1950_),
    .A(_1909_),
    .B(_1949_));
 sg13g2_nor2_1 _2805_ (.A(net689),
    .B(_1905_),
    .Y(_1951_));
 sg13g2_o21ai_1 _2806_ (.B1(_1878_),
    .Y(_1952_),
    .A1(_1925_),
    .A2(_1951_));
 sg13g2_nand4_1 _2807_ (.B(_1944_),
    .C(_1945_),
    .A(_1942_),
    .Y(_1953_),
    .D(_1952_));
 sg13g2_nand4_1 _2808_ (.B(_1900_),
    .C(_1948_),
    .A(_1898_),
    .Y(_1954_),
    .D(_1950_));
 sg13g2_nor4_2 _2809_ (.A(_1928_),
    .B(_1947_),
    .C(_1953_),
    .Y(_1955_),
    .D(_1954_));
 sg13g2_xor2_1 _2810_ (.B(_1955_),
    .A(net8),
    .X(_1956_));
 sg13g2_xnor2_1 _2811_ (.Y(_1957_),
    .A(net8),
    .B(_1955_));
 sg13g2_and2_1 _2812_ (.A(net630),
    .B(net629),
    .X(_1958_));
 sg13g2_and3_1 _2813_ (.X(_1959_),
    .A(_0060_),
    .B(net630),
    .C(net629));
 sg13g2_nand2_1 _2814_ (.Y(_1960_),
    .A(net693),
    .B(net630));
 sg13g2_o21ai_1 _2815_ (.B1(_1956_),
    .Y(_1961_),
    .A1(_1834_),
    .A2(net630));
 sg13g2_a21oi_1 _2816_ (.A1(_1960_),
    .A2(_1961_),
    .Y(_1962_),
    .B1(_1959_));
 sg13g2_a21o_1 _2817_ (.A2(_1961_),
    .A1(_1960_),
    .B1(_1959_),
    .X(_1963_));
 sg13g2_nand3_1 _2818_ (.B(net630),
    .C(net629),
    .A(_0069_),
    .Y(_1964_));
 sg13g2_o21ai_1 _2819_ (.B1(net695),
    .Y(_1965_),
    .A1(net644),
    .A2(net643));
 sg13g2_nor3_1 _2820_ (.A(_1835_),
    .B(net644),
    .C(net643),
    .Y(_1966_));
 sg13g2_nand3b_1 _2821_ (.B(_1939_),
    .C(_0070_),
    .Y(_1967_),
    .A_N(net644));
 sg13g2_a22oi_1 _2822_ (.Y(_1968_),
    .B1(_1956_),
    .B2(_1967_),
    .A2(net631),
    .A1(net695));
 sg13g2_o21ai_1 _2823_ (.B1(_1965_),
    .Y(_1969_),
    .A1(_1957_),
    .A2(_1966_));
 sg13g2_nand2_1 _2824_ (.Y(_1970_),
    .A(_1964_),
    .B(_1969_));
 sg13g2_nand3_1 _2825_ (.B(net630),
    .C(net629),
    .A(_0071_),
    .Y(_1971_));
 sg13g2_o21ai_1 _2826_ (.B1(net694),
    .Y(_1972_),
    .A1(net644),
    .A2(_1938_));
 sg13g2_nor3_1 _2827_ (.A(_1836_),
    .B(net645),
    .C(net643),
    .Y(_1973_));
 sg13g2_nand3b_1 _2828_ (.B(_1939_),
    .C(_0072_),
    .Y(_1974_),
    .A_N(net644));
 sg13g2_a22oi_1 _2829_ (.Y(_1975_),
    .B1(net629),
    .B2(_1974_),
    .A2(net631),
    .A1(net694));
 sg13g2_o21ai_1 _2830_ (.B1(_1972_),
    .Y(_1976_),
    .A1(_1957_),
    .A2(_1973_));
 sg13g2_a221oi_1 _2831_ (.B2(_1976_),
    .C1(_1968_),
    .B1(_1971_),
    .A1(_0069_),
    .Y(_1977_),
    .A2(_1958_));
 sg13g2_nand3_1 _2832_ (.B(net630),
    .C(net629),
    .A(_0072_),
    .Y(_1978_));
 sg13g2_o21ai_1 _2833_ (.B1(net696),
    .Y(_1979_),
    .A1(net644),
    .A2(net643));
 sg13g2_nor3_1 _2834_ (.A(_1837_),
    .B(net645),
    .C(net643),
    .Y(_1980_));
 sg13g2_nand3b_1 _2835_ (.B(_1939_),
    .C(_0073_),
    .Y(_1981_),
    .A_N(net645));
 sg13g2_a22oi_1 _2836_ (.Y(_1982_),
    .B1(_1956_),
    .B2(_1981_),
    .A2(net631),
    .A1(net696));
 sg13g2_o21ai_1 _2837_ (.B1(_1979_),
    .Y(_1983_),
    .A1(_1957_),
    .A2(_1980_));
 sg13g2_and2_1 _2838_ (.A(_1978_),
    .B(_1983_),
    .X(_1984_));
 sg13g2_nand2_1 _2839_ (.Y(_1985_),
    .A(_1978_),
    .B(_1983_));
 sg13g2_nand3_1 _2840_ (.B(net630),
    .C(net629),
    .A(_0070_),
    .Y(_1986_));
 sg13g2_o21ai_1 _2841_ (.B1(net697),
    .Y(_1987_),
    .A1(net645),
    .A2(net643));
 sg13g2_nor3_1 _2842_ (.A(net698),
    .B(net644),
    .C(net643),
    .Y(_1988_));
 sg13g2_or3_1 _2843_ (.A(net698),
    .B(net645),
    .C(net643),
    .X(_1989_));
 sg13g2_a22oi_1 _2844_ (.Y(_1990_),
    .B1(net629),
    .B2(_1989_),
    .A2(net631),
    .A1(net697));
 sg13g2_o21ai_1 _2845_ (.B1(_1987_),
    .Y(_1991_),
    .A1(_1957_),
    .A2(_1988_));
 sg13g2_and2_2 _2846_ (.A(_1986_),
    .B(_1991_),
    .X(_1992_));
 sg13g2_nand2_2 _2847_ (.Y(_1993_),
    .A(_1986_),
    .B(_1991_));
 sg13g2_a221oi_1 _2848_ (.B2(_1983_),
    .C1(_1990_),
    .B1(_1978_),
    .A1(_0070_),
    .Y(_1994_),
    .A2(_1958_));
 sg13g2_and3_2 _2849_ (.X(_1995_),
    .A(net622),
    .B(net609),
    .C(net601));
 sg13g2_nand3_1 _2850_ (.B(net609),
    .C(net601),
    .A(net623),
    .Y(_1996_));
 sg13g2_a221oi_1 _2851_ (.B2(_1991_),
    .C1(_1982_),
    .B1(_1986_),
    .A1(_0072_),
    .Y(_1997_),
    .A2(_1958_));
 sg13g2_a22oi_1 _2852_ (.Y(_1998_),
    .B1(_1971_),
    .B2(_1976_),
    .A2(_1969_),
    .A1(_1964_));
 sg13g2_and2_2 _2853_ (.A(net624),
    .B(net596),
    .X(_1999_));
 sg13g2_nand2_2 _2854_ (.Y(_2000_),
    .A(net622),
    .B(net594));
 sg13g2_nand2_2 _2855_ (.Y(_2001_),
    .A(net599),
    .B(net595));
 sg13g2_and3_1 _2856_ (.X(_2002_),
    .A(net621),
    .B(net597),
    .C(net593));
 sg13g2_nand3_1 _2857_ (.B(net597),
    .C(net594),
    .A(net621),
    .Y(_2003_));
 sg13g2_and4_1 _2858_ (.A(_1964_),
    .B(_1969_),
    .C(_1971_),
    .D(_1976_),
    .X(_2004_));
 sg13g2_nand4_1 _2859_ (.B(_1969_),
    .C(_1971_),
    .A(_1964_),
    .Y(_2005_),
    .D(_1976_));
 sg13g2_nor2_2 _2860_ (.A(net614),
    .B(net590),
    .Y(_2006_));
 sg13g2_nand2_2 _2861_ (.Y(_2007_),
    .A(net624),
    .B(net592));
 sg13g2_nor3_2 _2862_ (.A(net614),
    .B(_1993_),
    .C(net590),
    .Y(_2008_));
 sg13g2_nand2_2 _2863_ (.Y(_2009_),
    .A(_1992_),
    .B(_2006_));
 sg13g2_and2_2 _2864_ (.A(net601),
    .B(_2006_),
    .X(_2010_));
 sg13g2_nand3_1 _2865_ (.B(net600),
    .C(net592),
    .A(net618),
    .Y(_2011_));
 sg13g2_nand3_1 _2866_ (.B(net574),
    .C(_2011_),
    .A(_1996_),
    .Y(_2012_));
 sg13g2_and4_1 _2867_ (.A(_1978_),
    .B(_1983_),
    .C(_1986_),
    .D(_1991_),
    .X(_2013_));
 sg13g2_a22oi_1 _2868_ (.Y(_2014_),
    .B1(_1986_),
    .B2(_1991_),
    .A2(_1983_),
    .A1(_1978_));
 sg13g2_nor2_2 _2869_ (.A(net624),
    .B(net589),
    .Y(_2015_));
 sg13g2_nand2_2 _2870_ (.Y(_2016_),
    .A(net612),
    .B(net592));
 sg13g2_nor3_2 _2871_ (.A(net619),
    .B(net589),
    .C(net583),
    .Y(_2017_));
 sg13g2_nor2b_2 _2872_ (.A(net586),
    .B_N(_2017_),
    .Y(_2018_));
 sg13g2_or4_2 _2873_ (.A(net619),
    .B(net589),
    .C(net586),
    .D(net581),
    .X(_2019_));
 sg13g2_a221oi_1 _2874_ (.B2(_1969_),
    .C1(_1975_),
    .B1(_1964_),
    .A1(_0071_),
    .Y(_2020_),
    .A2(_1958_));
 sg13g2_nand2_2 _2875_ (.Y(_2021_),
    .A(net602),
    .B(net579));
 sg13g2_nand2_2 _2876_ (.Y(_2022_),
    .A(net598),
    .B(net578));
 sg13g2_and3_2 _2877_ (.X(_2023_),
    .A(net611),
    .B(net600),
    .C(net577));
 sg13g2_nand3_1 _2878_ (.B(net600),
    .C(net576),
    .A(net612),
    .Y(_2024_));
 sg13g2_and3_1 _2879_ (.X(_2025_),
    .A(net612),
    .B(net599),
    .C(net576));
 sg13g2_nand3_1 _2880_ (.B(net597),
    .C(net578),
    .A(net614),
    .Y(_2026_));
 sg13g2_nor2_2 _2881_ (.A(_2023_),
    .B(net570),
    .Y(_2027_));
 sg13g2_nand3_1 _2882_ (.B(_2024_),
    .C(_2026_),
    .A(_2019_),
    .Y(_2028_));
 sg13g2_nor3_2 _2883_ (.A(net614),
    .B(net603),
    .C(net590),
    .Y(_2029_));
 sg13g2_nand3_1 _2884_ (.B(net605),
    .C(net591),
    .A(net621),
    .Y(_2030_));
 sg13g2_nor4_2 _2885_ (.A(net616),
    .B(net603),
    .C(_1993_),
    .Y(_2031_),
    .D(net589));
 sg13g2_nand2_2 _2886_ (.Y(_2032_),
    .A(net573),
    .B(net585));
 sg13g2_and3_2 _2887_ (.X(_2033_),
    .A(net612),
    .B(net608),
    .C(net600));
 sg13g2_nand3_1 _2888_ (.B(net607),
    .C(net600),
    .A(net612),
    .Y(_2034_));
 sg13g2_nand2b_1 _2889_ (.Y(_2035_),
    .B(net568),
    .A_N(_2031_));
 sg13g2_and3_1 _2890_ (.X(_2036_),
    .A(net615),
    .B(net609),
    .C(net583));
 sg13g2_nand3_1 _2891_ (.B(net607),
    .C(net581),
    .A(net611),
    .Y(_2037_));
 sg13g2_and3_2 _2892_ (.X(_2038_),
    .A(net611),
    .B(net607),
    .C(net585));
 sg13g2_nand3_1 _2893_ (.B(net607),
    .C(net585),
    .A(net611),
    .Y(_2039_));
 sg13g2_nor2_1 _2894_ (.A(net566),
    .B(_2038_),
    .Y(_2040_));
 sg13g2_nand2_1 _2895_ (.Y(_2041_),
    .A(net565),
    .B(net564));
 sg13g2_and3_2 _2896_ (.X(_2042_),
    .A(net615),
    .B(net598),
    .C(net595));
 sg13g2_nand3_1 _2897_ (.B(net597),
    .C(net593),
    .A(net613),
    .Y(_2043_));
 sg13g2_and3_2 _2898_ (.X(_2044_),
    .A(net613),
    .B(net593),
    .C(net587));
 sg13g2_nand3_1 _2899_ (.B(net596),
    .C(net586),
    .A(net617),
    .Y(_2045_));
 sg13g2_and3_2 _2900_ (.X(_2046_),
    .A(net614),
    .B(net605),
    .C(net594));
 sg13g2_nand3_1 _2901_ (.B(net606),
    .C(net596),
    .A(net612),
    .Y(_2047_));
 sg13g2_nor2_2 _2902_ (.A(_1993_),
    .B(_2000_),
    .Y(_2048_));
 sg13g2_and3_1 _2903_ (.X(_2049_),
    .A(net623),
    .B(net601),
    .C(net593));
 sg13g2_nand3_1 _2904_ (.B(net601),
    .C(net593),
    .A(net621),
    .Y(_2050_));
 sg13g2_nor2_2 _2905_ (.A(_2046_),
    .B(net562),
    .Y(_2051_));
 sg13g2_and3_1 _2906_ (.X(_2052_),
    .A(net618),
    .B(net599),
    .C(net576));
 sg13g2_and3_2 _2907_ (.X(_2053_),
    .A(net618),
    .B(net600),
    .C(net577));
 sg13g2_nand3_1 _2908_ (.B(net601),
    .C(net578),
    .A(net622),
    .Y(_2054_));
 sg13g2_nor2_2 _2909_ (.A(_2052_),
    .B(_2053_),
    .Y(_2055_));
 sg13g2_nor3_1 _2910_ (.A(_2012_),
    .B(_2028_),
    .C(_2035_),
    .Y(_2056_));
 sg13g2_nand4_1 _2911_ (.B(_2051_),
    .C(_2055_),
    .A(_2040_),
    .Y(_2057_),
    .D(_2056_));
 sg13g2_nor2b_2 _2912_ (.A(\wirecube_top_inst.line_rom_inst.line_i[0] ),
    .B_N(\wirecube_top_inst.line_rom_inst.line_i[1] ),
    .Y(_2058_));
 sg13g2_nor2b_2 _2913_ (.A(net679),
    .B_N(net678),
    .Y(_2059_));
 sg13g2_nand2b_2 _2914_ (.Y(_2060_),
    .B(net678),
    .A_N(net679));
 sg13g2_and2_2 _2915_ (.A(_2058_),
    .B(_2059_),
    .X(_2061_));
 sg13g2_nand2_2 _2916_ (.Y(_2062_),
    .A(_2058_),
    .B(_2059_));
 sg13g2_nor2b_2 _2917_ (.A(net678),
    .B_N(net680),
    .Y(_2063_));
 sg13g2_and2_1 _2918_ (.A(_2058_),
    .B(_2063_),
    .X(_2064_));
 sg13g2_nand2_1 _2919_ (.Y(_2065_),
    .A(_2058_),
    .B(_2063_));
 sg13g2_nand2_1 _2920_ (.Y(_2066_),
    .A(_2062_),
    .B(_2065_));
 sg13g2_nand2_1 _2921_ (.Y(_2067_),
    .A(\wirecube_top_inst.line_rom_inst.line_i[3] ),
    .B(net679));
 sg13g2_nor2_2 _2922_ (.A(net201),
    .B(\wirecube_top_inst.line_rom_inst.line_i[0] ),
    .Y(_2068_));
 sg13g2_inv_1 _2923_ (.Y(_2069_),
    .A(_2068_));
 sg13g2_o21ai_1 _2924_ (.B1(_2060_),
    .Y(_2070_),
    .A1(net678),
    .A2(_2068_));
 sg13g2_o21ai_1 _2925_ (.B1(_2067_),
    .Y(_2071_),
    .A1(net678),
    .A2(_2069_));
 sg13g2_nor2_1 _2926_ (.A(_2063_),
    .B(_2070_),
    .Y(_2072_));
 sg13g2_or2_1 _2927_ (.X(_2073_),
    .B(_2070_),
    .A(_2063_));
 sg13g2_nand2b_1 _2928_ (.Y(_2074_),
    .B(net649),
    .A_N(net654));
 sg13g2_nor2_2 _2929_ (.A(net603),
    .B(_2000_),
    .Y(_2075_));
 sg13g2_nor2_1 _2930_ (.A(_2048_),
    .B(_2075_),
    .Y(_2076_));
 sg13g2_nand2_2 _2931_ (.Y(_2077_),
    .A(net574),
    .B(net561));
 sg13g2_a221oi_1 _2932_ (.B2(net604),
    .C1(net562),
    .B1(_2015_),
    .A1(net599),
    .Y(_2078_),
    .A2(_1999_));
 sg13g2_nand2_2 _2933_ (.Y(_2079_),
    .A(net591),
    .B(net583));
 sg13g2_nor4_2 _2934_ (.A(net622),
    .B(net605),
    .C(_1992_),
    .Y(_2080_),
    .D(net590));
 sg13g2_nand3_1 _2935_ (.B(net591),
    .C(net583),
    .A(net613),
    .Y(_2081_));
 sg13g2_and3_1 _2936_ (.X(_2082_),
    .A(net615),
    .B(net601),
    .C(net595));
 sg13g2_nand3_1 _2937_ (.B(net601),
    .C(net593),
    .A(net613),
    .Y(_2083_));
 sg13g2_nor2_2 _2938_ (.A(_2038_),
    .B(net558),
    .Y(_2084_));
 sg13g2_nor3_1 _2939_ (.A(_2038_),
    .B(_2080_),
    .C(net558),
    .Y(_2085_));
 sg13g2_nor2_2 _2940_ (.A(net566),
    .B(_2044_),
    .Y(_2086_));
 sg13g2_nand2_2 _2941_ (.Y(_2087_),
    .A(net565),
    .B(_2045_));
 sg13g2_nor2_2 _2942_ (.A(net567),
    .B(_2046_),
    .Y(_2088_));
 sg13g2_and2_1 _2943_ (.A(net588),
    .B(net579),
    .X(_2089_));
 sg13g2_nand3_1 _2944_ (.B(net587),
    .C(net578),
    .A(net621),
    .Y(_2090_));
 sg13g2_nand3_1 _2945_ (.B(net606),
    .C(net576),
    .A(net618),
    .Y(_2091_));
 sg13g2_and3_1 _2946_ (.X(_2092_),
    .A(net623),
    .B(net604),
    .C(net578));
 sg13g2_nor2_1 _2947_ (.A(_2023_),
    .B(net555),
    .Y(_2093_));
 sg13g2_nand4_1 _2948_ (.B(_2085_),
    .C(_2088_),
    .A(_2078_),
    .Y(_2094_),
    .D(_2093_));
 sg13g2_nor2_1 _2949_ (.A(\wirecube_top_inst.line_rom_inst.line_i[3] ),
    .B(net679),
    .Y(_2095_));
 sg13g2_nor3_1 _2950_ (.A(\wirecube_top_inst.line_rom_inst.line_i[0] ),
    .B(net678),
    .C(net679),
    .Y(_2096_));
 sg13g2_and2_1 _2951_ (.A(\wirecube_top_inst.line_rom_inst.line_i[1] ),
    .B(_2096_),
    .X(_2097_));
 sg13g2_nand2_2 _2952_ (.Y(_2098_),
    .A(\wirecube_top_inst.line_rom_inst.line_i[1] ),
    .B(net677));
 sg13g2_nor2_2 _2953_ (.A(_2060_),
    .B(_2069_),
    .Y(_2099_));
 sg13g2_nand2_1 _2954_ (.Y(_2100_),
    .A(_2059_),
    .B(_2068_));
 sg13g2_nand2b_2 _2955_ (.Y(_2101_),
    .B(\wirecube_top_inst.line_rom_inst.line_i[0] ),
    .A_N(\wirecube_top_inst.line_rom_inst.line_i[1] ));
 sg13g2_nor2_2 _2956_ (.A(net678),
    .B(_2101_),
    .Y(_2102_));
 sg13g2_or2_2 _2957_ (.X(_2103_),
    .B(_2101_),
    .A(net678));
 sg13g2_nand2_2 _2958_ (.Y(_2104_),
    .A(net680),
    .B(_2102_));
 sg13g2_and2_2 _2959_ (.A(net661),
    .B(_2104_),
    .X(_2105_));
 sg13g2_nand2_2 _2960_ (.Y(_2106_),
    .A(net661),
    .B(_2104_));
 sg13g2_o21ai_1 _2961_ (.B1(_2094_),
    .Y(_2107_),
    .A1(net663),
    .A2(_2106_));
 sg13g2_a22oi_1 _2962_ (.Y(_2108_),
    .B1(net585),
    .B2(net576),
    .A2(net592),
    .A1(net611));
 sg13g2_and3_1 _2963_ (.X(_2109_),
    .A(net623),
    .B(net595),
    .C(net587));
 sg13g2_nand3_1 _2964_ (.B(net596),
    .C(net585),
    .A(net618),
    .Y(_2110_));
 sg13g2_and2_1 _2965_ (.A(net608),
    .B(net599),
    .X(_2111_));
 sg13g2_and3_2 _2966_ (.X(_2112_),
    .A(net622),
    .B(net610),
    .C(net597));
 sg13g2_nand3_1 _2967_ (.B(net610),
    .C(net598),
    .A(net621),
    .Y(_2113_));
 sg13g2_and3_2 _2968_ (.X(_2114_),
    .A(net619),
    .B(net608),
    .C(net582));
 sg13g2_nand3_1 _2969_ (.B(net607),
    .C(net582),
    .A(net619),
    .Y(_2115_));
 sg13g2_nand3_1 _2970_ (.B(net609),
    .C(_1993_),
    .A(net623),
    .Y(_2116_));
 sg13g2_nand3_1 _2971_ (.B(_1970_),
    .C(net602),
    .A(net616),
    .Y(_2117_));
 sg13g2_and2_1 _2972_ (.A(_2047_),
    .B(_2117_),
    .X(_2118_));
 sg13g2_and4_1 _2973_ (.A(_2079_),
    .B(_2108_),
    .C(_2110_),
    .D(_2116_),
    .X(_2119_));
 sg13g2_and3_1 _2974_ (.X(_2120_),
    .A(net615),
    .B(net587),
    .C(net578));
 sg13g2_nand3_1 _2975_ (.B(net587),
    .C(net578),
    .A(net615),
    .Y(_2121_));
 sg13g2_nand2_1 _2976_ (.Y(_2122_),
    .A(_2118_),
    .B(_2119_));
 sg13g2_and2_2 _2977_ (.A(\wirecube_top_inst.line_rom_inst.line_i[1] ),
    .B(\wirecube_top_inst.line_rom_inst.line_i[0] ),
    .X(_2123_));
 sg13g2_nand2_2 _2978_ (.Y(_2124_),
    .A(\wirecube_top_inst.line_rom_inst.line_i[1] ),
    .B(\wirecube_top_inst.line_rom_inst.line_i[0] ));
 sg13g2_and2_2 _2979_ (.A(_2095_),
    .B(_2123_),
    .X(_2125_));
 sg13g2_nand2_2 _2980_ (.Y(_2126_),
    .A(_2095_),
    .B(_2123_));
 sg13g2_nand2_1 _2981_ (.Y(_2127_),
    .A(_2063_),
    .B(_2123_));
 sg13g2_nor2_2 _2982_ (.A(_2060_),
    .B(_2101_),
    .Y(_2128_));
 sg13g2_or2_2 _2983_ (.X(_2129_),
    .B(_2101_),
    .A(_2060_));
 sg13g2_and2_2 _2984_ (.A(net658),
    .B(_2129_),
    .X(_2130_));
 sg13g2_nand2_1 _2985_ (.Y(_2131_),
    .A(net658),
    .B(_2129_));
 sg13g2_o21ai_1 _2986_ (.B1(_2122_),
    .Y(_2132_),
    .A1(net659),
    .A2(net648));
 sg13g2_nor2_2 _2987_ (.A(_2053_),
    .B(net555),
    .Y(_2133_));
 sg13g2_nand2_1 _2988_ (.Y(_2134_),
    .A(net560),
    .B(_2091_));
 sg13g2_and3_2 _2989_ (.X(_2135_),
    .A(net623),
    .B(net609),
    .C(net587));
 sg13g2_nand3_1 _2990_ (.B(net610),
    .C(net587),
    .A(net621),
    .Y(_2136_));
 sg13g2_nand3_1 _2991_ (.B(net607),
    .C(net606),
    .A(net618),
    .Y(_2137_));
 sg13g2_and3_2 _2992_ (.X(_2138_),
    .A(net619),
    .B(net608),
    .C(net606));
 sg13g2_nand2_1 _2993_ (.Y(_2139_),
    .A(net560),
    .B(_2136_));
 sg13g2_nor3_2 _2994_ (.A(_2053_),
    .B(net555),
    .C(_2138_),
    .Y(_2140_));
 sg13g2_nor3_2 _2995_ (.A(net615),
    .B(net604),
    .C(net589),
    .Y(_2141_));
 sg13g2_nand2_1 _2996_ (.Y(_2142_),
    .A(net603),
    .B(net573));
 sg13g2_nor2_2 _2997_ (.A(net598),
    .B(_2007_),
    .Y(_2143_));
 sg13g2_nor4_1 _2998_ (.A(_2008_),
    .B(_2017_),
    .C(net571),
    .D(_2141_),
    .Y(_2144_));
 sg13g2_nor2_2 _2999_ (.A(_1995_),
    .B(_2114_),
    .Y(_2145_));
 sg13g2_and3_2 _3000_ (.X(_2146_),
    .A(net622),
    .B(net609),
    .C(_1985_));
 sg13g2_nand4_1 _3001_ (.B(_2140_),
    .C(_2144_),
    .A(_2051_),
    .Y(_2147_),
    .D(_2145_));
 sg13g2_nor2_2 _3002_ (.A(net680),
    .B(_2103_),
    .Y(_2148_));
 sg13g2_nand2b_2 _3003_ (.Y(_2149_),
    .B(_2102_),
    .A_N(net679));
 sg13g2_nor2_2 _3004_ (.A(_2060_),
    .B(_2124_),
    .Y(_2150_));
 sg13g2_nand2_2 _3005_ (.Y(_2151_),
    .A(_2059_),
    .B(_2123_));
 sg13g2_nand2_2 _3006_ (.Y(_2152_),
    .A(_2063_),
    .B(_2068_));
 sg13g2_and2_2 _3007_ (.A(_2151_),
    .B(_2152_),
    .X(_2153_));
 sg13g2_nand2_2 _3008_ (.Y(_2154_),
    .A(_2151_),
    .B(_2152_));
 sg13g2_o21ai_1 _3009_ (.B1(_2147_),
    .Y(_2155_),
    .A1(_2148_),
    .A2(_2154_));
 sg13g2_nand3_1 _3010_ (.B(_2132_),
    .C(_2155_),
    .A(_2107_),
    .Y(_2156_));
 sg13g2_a21oi_2 _3011_ (.B1(_2156_),
    .Y(_2157_),
    .A2(_2074_),
    .A1(_2057_));
 sg13g2_a21o_1 _3012_ (.A2(_2074_),
    .A1(_2057_),
    .B1(_2156_),
    .X(_2158_));
 sg13g2_nor2_1 _3013_ (.A(net634),
    .B(_2157_),
    .Y(_2159_));
 sg13g2_and2_2 _3014_ (.A(net596),
    .B(net581),
    .X(_2160_));
 sg13g2_nand2_1 _3015_ (.Y(_2161_),
    .A(net596),
    .B(net581));
 sg13g2_nand2_2 _3016_ (.Y(_2162_),
    .A(_2043_),
    .B(_2083_));
 sg13g2_nor2_2 _3017_ (.A(net604),
    .B(_2000_),
    .Y(_2163_));
 sg13g2_or2_2 _3018_ (.X(_2164_),
    .B(_2141_),
    .A(net575));
 sg13g2_nor3_1 _3019_ (.A(net575),
    .B(net573),
    .C(_2163_),
    .Y(_2165_));
 sg13g2_nand2_2 _3020_ (.Y(_2166_),
    .A(net584),
    .B(net579));
 sg13g2_and3_2 _3021_ (.X(_2167_),
    .A(net618),
    .B(net581),
    .C(net576));
 sg13g2_nand3_1 _3022_ (.B(net581),
    .C(net576),
    .A(net618),
    .Y(_2168_));
 sg13g2_and3_2 _3023_ (.X(_2169_),
    .A(net619),
    .B(net603),
    .C(net577));
 sg13g2_and3_2 _3024_ (.X(_2170_),
    .A(net611),
    .B(net582),
    .C(net577));
 sg13g2_nand3_1 _3025_ (.B(net581),
    .C(net576),
    .A(net611),
    .Y(_2171_));
 sg13g2_nor2_1 _3026_ (.A(_2023_),
    .B(_2170_),
    .Y(_2172_));
 sg13g2_and3_2 _3027_ (.X(_2173_),
    .A(net614),
    .B(net603),
    .C(net578));
 sg13g2_nand3_1 _3028_ (.B(_2145_),
    .C(_2166_),
    .A(_2021_),
    .Y(_2174_));
 sg13g2_and3_1 _3029_ (.X(_2175_),
    .A(net613),
    .B(net609),
    .C(net597));
 sg13g2_nand3_1 _3030_ (.B(net609),
    .C(net597),
    .A(net613),
    .Y(_2176_));
 sg13g2_nand3_1 _3031_ (.B(_2090_),
    .C(_2176_),
    .A(_2022_),
    .Y(_2177_));
 sg13g2_nand2_2 _3032_ (.Y(_2178_),
    .A(net568),
    .B(net551));
 sg13g2_nor2_2 _3033_ (.A(net553),
    .B(_2138_),
    .Y(_2179_));
 sg13g2_nand4_1 _3034_ (.B(net564),
    .C(net550),
    .A(_2034_),
    .Y(_2180_),
    .D(_2179_));
 sg13g2_nor3_2 _3035_ (.A(_2174_),
    .B(_2177_),
    .C(_2180_),
    .Y(_2181_));
 sg13g2_nand4_1 _3036_ (.B(_2086_),
    .C(_2165_),
    .A(_2016_),
    .Y(_2182_),
    .D(_2181_));
 sg13g2_and3_1 _3037_ (.X(_2183_),
    .A(net613),
    .B(net593),
    .C(net583));
 sg13g2_nand3_1 _3038_ (.B(net593),
    .C(net583),
    .A(net613),
    .Y(_2184_));
 sg13g2_nor3_2 _3039_ (.A(net623),
    .B(net604),
    .C(net589),
    .Y(_2185_));
 sg13g2_nand3_1 _3040_ (.B(net603),
    .C(net591),
    .A(net616),
    .Y(_2186_));
 sg13g2_nor2_2 _3041_ (.A(_1993_),
    .B(_2186_),
    .Y(_2187_));
 sg13g2_nand3_1 _3042_ (.B(net602),
    .C(net591),
    .A(net616),
    .Y(_2188_));
 sg13g2_nor2_1 _3043_ (.A(_2044_),
    .B(_2170_),
    .Y(_2189_));
 sg13g2_nand2_2 _3044_ (.Y(_2190_),
    .A(_2045_),
    .B(_2171_));
 sg13g2_nand4_1 _3045_ (.B(net564),
    .C(net556),
    .A(_2022_),
    .Y(_2191_),
    .D(_2113_));
 sg13g2_or4_2 _3046_ (.A(_2035_),
    .B(_2187_),
    .C(_2190_),
    .D(_2191_),
    .X(_2192_));
 sg13g2_o21ai_1 _3047_ (.B1(net653),
    .Y(_2193_),
    .A1(net545),
    .A2(_2192_));
 sg13g2_nor2_2 _3048_ (.A(_2031_),
    .B(_2146_),
    .Y(_2194_));
 sg13g2_nor3_2 _3049_ (.A(net600),
    .B(net599),
    .C(_2016_),
    .Y(_2195_));
 sg13g2_a21oi_1 _3050_ (.A1(net587),
    .A2(_2015_),
    .Y(_2196_),
    .B1(_2080_));
 sg13g2_nor2_1 _3051_ (.A(net570),
    .B(_2195_),
    .Y(_2197_));
 sg13g2_nand2_2 _3052_ (.Y(_2198_),
    .A(_2026_),
    .B(_2196_));
 sg13g2_and3_2 _3053_ (.X(_2199_),
    .A(net611),
    .B(net607),
    .C(net606));
 sg13g2_nor2_1 _3054_ (.A(net566),
    .B(_2170_),
    .Y(_2200_));
 sg13g2_nand2_1 _3055_ (.Y(_2201_),
    .A(net565),
    .B(_2171_));
 sg13g2_nor4_2 _3056_ (.A(_2139_),
    .B(net544),
    .C(_2199_),
    .Y(_2202_),
    .D(_2201_));
 sg13g2_nand4_1 _3057_ (.B(_2194_),
    .C(_2197_),
    .A(_2051_),
    .Y(_2203_),
    .D(_2202_));
 sg13g2_nand2_1 _3058_ (.Y(_2204_),
    .A(net648),
    .B(_2203_));
 sg13g2_nand2_1 _3059_ (.Y(_2205_),
    .A(_1996_),
    .B(_2027_));
 sg13g2_nor4_2 _3060_ (.A(net622),
    .B(net603),
    .C(_1993_),
    .Y(_2206_),
    .D(net589));
 sg13g2_nand4_1 _3061_ (.B(net605),
    .C(_1992_),
    .A(net614),
    .Y(_2207_),
    .D(net591));
 sg13g2_nand3_1 _3062_ (.B(_2001_),
    .C(_2207_),
    .A(_2000_),
    .Y(_2208_));
 sg13g2_nand2_2 _3063_ (.Y(_2209_),
    .A(_2113_),
    .B(_2168_));
 sg13g2_nor4_2 _3064_ (.A(net615),
    .B(net604),
    .C(_1992_),
    .Y(_2210_),
    .D(net589));
 sg13g2_nor4_1 _3065_ (.A(net566),
    .B(_2208_),
    .C(_2209_),
    .D(_2210_),
    .Y(_2211_));
 sg13g2_nor2b_1 _3066_ (.A(_2205_),
    .B_N(_2211_),
    .Y(_2212_));
 sg13g2_and2_1 _3067_ (.A(net542),
    .B(_2212_),
    .X(_2213_));
 sg13g2_nand2_2 _3068_ (.Y(_2214_),
    .A(net551),
    .B(_2188_));
 sg13g2_nand2_2 _3069_ (.Y(_2215_),
    .A(net574),
    .B(net568));
 sg13g2_nor4_1 _3070_ (.A(_2169_),
    .B(_2199_),
    .C(_2214_),
    .D(_2215_),
    .Y(_2216_));
 sg13g2_nor2_2 _3071_ (.A(_1992_),
    .B(net569),
    .Y(_2217_));
 sg13g2_nand3_1 _3072_ (.B(net597),
    .C(net591),
    .A(net621),
    .Y(_2218_));
 sg13g2_nor3_1 _3073_ (.A(_2087_),
    .B(_2160_),
    .C(_2217_),
    .Y(_2219_));
 sg13g2_nand4_1 _3074_ (.B(_2116_),
    .C(_2216_),
    .A(_2091_),
    .Y(_2220_),
    .D(_2219_));
 sg13g2_nor2_1 _3075_ (.A(net554),
    .B(net546),
    .Y(_2221_));
 sg13g2_nand2_1 _3076_ (.Y(_2222_),
    .A(_2110_),
    .B(net541));
 sg13g2_nor2_1 _3077_ (.A(_1995_),
    .B(_2143_),
    .Y(_2223_));
 sg13g2_o21ai_1 _3078_ (.B1(_2223_),
    .Y(_2224_),
    .A1(net600),
    .A2(_2016_));
 sg13g2_nand4_1 _3079_ (.B(_2026_),
    .C(_2043_),
    .A(_2024_),
    .Y(_2225_),
    .D(net561));
 sg13g2_nand3_1 _3080_ (.B(_2136_),
    .C(_2171_),
    .A(net557),
    .Y(_2226_));
 sg13g2_nor4_2 _3081_ (.A(_2222_),
    .B(_2224_),
    .C(_2225_),
    .Y(_2227_),
    .D(_2226_));
 sg13g2_nor2_1 _3082_ (.A(_2153_),
    .B(_2227_),
    .Y(_2228_));
 sg13g2_nor2_1 _3083_ (.A(_2160_),
    .B(_2178_),
    .Y(_2229_));
 sg13g2_nor3_2 _3084_ (.A(net553),
    .B(_2112_),
    .C(_2217_),
    .Y(_2230_));
 sg13g2_nand2_1 _3085_ (.Y(_2231_),
    .A(net556),
    .B(_2168_));
 sg13g2_nand2_2 _3086_ (.Y(_2232_),
    .A(_2091_),
    .B(_2168_));
 sg13g2_nand2_1 _3087_ (.Y(_2233_),
    .A(_2019_),
    .B(_2024_));
 sg13g2_nor4_2 _3088_ (.A(net558),
    .B(_2164_),
    .C(_2232_),
    .Y(_2234_),
    .D(_2233_));
 sg13g2_nand3_1 _3089_ (.B(_2230_),
    .C(_2234_),
    .A(_2229_),
    .Y(_2235_));
 sg13g2_nand2_1 _3090_ (.Y(_2236_),
    .A(_2106_),
    .B(_2212_));
 sg13g2_a22oi_1 _3091_ (.Y(_2237_),
    .B1(_2235_),
    .B2(net659),
    .A2(_2220_),
    .A1(net647));
 sg13g2_nand2_1 _3092_ (.Y(_2238_),
    .A(_2236_),
    .B(_2237_));
 sg13g2_o21ai_1 _3093_ (.B1(_2193_),
    .Y(_2239_),
    .A1(_2098_),
    .A2(_2213_));
 sg13g2_o21ai_1 _3094_ (.B1(_2204_),
    .Y(_2240_),
    .A1(net649),
    .A2(_2192_));
 sg13g2_nor4_2 _3095_ (.A(_2228_),
    .B(_2238_),
    .C(_2239_),
    .Y(_2241_),
    .D(_2240_));
 sg13g2_a21oi_2 _3096_ (.B1(_2159_),
    .Y(_2242_),
    .A2(_2241_),
    .A1(net634));
 sg13g2_nor2_2 _3097_ (.A(_2064_),
    .B(_2125_),
    .Y(_2243_));
 sg13g2_nand2_2 _3098_ (.Y(_2244_),
    .A(_2065_),
    .B(_2126_));
 sg13g2_or4_2 _3099_ (.A(net553),
    .B(_2138_),
    .C(_2146_),
    .D(_2169_),
    .X(_2245_));
 sg13g2_inv_1 _3100_ (.Y(_2246_),
    .A(_2245_));
 sg13g2_nor2_2 _3101_ (.A(_2033_),
    .B(net567),
    .Y(_2247_));
 sg13g2_nand2_1 _3102_ (.Y(_2248_),
    .A(net568),
    .B(net565));
 sg13g2_nand2b_1 _3103_ (.Y(_2249_),
    .B(_2171_),
    .A_N(_2199_));
 sg13g2_a21oi_1 _3104_ (.A1(net617),
    .A2(net608),
    .Y(_2250_),
    .B1(_2170_));
 sg13g2_nor2_1 _3105_ (.A(_2062_),
    .B(_2250_),
    .Y(_2251_));
 sg13g2_nand2_2 _3106_ (.Y(_2252_),
    .A(_2076_),
    .B(_2145_));
 sg13g2_a21oi_1 _3107_ (.A1(net652),
    .A2(_2252_),
    .Y(_2253_),
    .B1(_2251_));
 sg13g2_and2_2 _3108_ (.A(_2098_),
    .B(net658),
    .X(_2254_));
 sg13g2_nand2_2 _3109_ (.Y(_2255_),
    .A(_2098_),
    .B(net658));
 sg13g2_and3_2 _3110_ (.X(_2256_),
    .A(net624),
    .B(_1993_),
    .C(net579));
 sg13g2_nand2_2 _3111_ (.Y(_2257_),
    .A(_2055_),
    .B(_2168_));
 sg13g2_nand2_2 _3112_ (.Y(_2258_),
    .A(net620),
    .B(net580));
 sg13g2_nor2_2 _3113_ (.A(net572),
    .B(net588),
    .Y(_2259_));
 sg13g2_o21ai_1 _3114_ (.B1(_2258_),
    .Y(_2260_),
    .A1(net572),
    .A2(net586));
 sg13g2_nand2_1 _3115_ (.Y(_2261_),
    .A(_2255_),
    .B(_2260_));
 sg13g2_nor2_1 _3116_ (.A(net571),
    .B(net552),
    .Y(_2262_));
 sg13g2_nand2_2 _3117_ (.Y(_2263_),
    .A(_2026_),
    .B(net550));
 sg13g2_nand2_2 _3118_ (.Y(_2264_),
    .A(_2024_),
    .B(_2262_));
 sg13g2_nor2_2 _3119_ (.A(_2080_),
    .B(net552),
    .Y(_2265_));
 sg13g2_nand2_1 _3120_ (.Y(_2266_),
    .A(_2081_),
    .B(net550));
 sg13g2_nor3_2 _3121_ (.A(_2080_),
    .B(net552),
    .C(_2170_),
    .Y(_2267_));
 sg13g2_nand4_1 _3122_ (.B(_2027_),
    .C(net551),
    .A(_2016_),
    .Y(_2268_),
    .D(_2171_));
 sg13g2_a22oi_1 _3123_ (.Y(_2269_),
    .B1(_2268_),
    .B2(net656),
    .A2(_2245_),
    .A1(_2244_));
 sg13g2_nand3_1 _3124_ (.B(_2261_),
    .C(_2269_),
    .A(_2253_),
    .Y(_2270_));
 sg13g2_nand2_1 _3125_ (.Y(_2271_),
    .A(net635),
    .B(_2270_));
 sg13g2_or2_1 _3126_ (.X(_2272_),
    .B(_2250_),
    .A(_2130_));
 sg13g2_a22oi_1 _3127_ (.Y(_2273_),
    .B1(_2268_),
    .B2(net654),
    .A2(_2245_),
    .A1(net663));
 sg13g2_a22oi_1 _3128_ (.Y(_2274_),
    .B1(_2260_),
    .B2(_2148_),
    .A2(_2252_),
    .A1(net659));
 sg13g2_nand3_1 _3129_ (.B(_2273_),
    .C(_2274_),
    .A(_2272_),
    .Y(_2275_));
 sg13g2_nor2_1 _3130_ (.A(_2271_),
    .B(_2275_),
    .Y(_2276_));
 sg13g2_nand3_1 _3131_ (.B(_2270_),
    .C(_2275_),
    .A(net635),
    .Y(_2277_));
 sg13g2_o21ai_1 _3132_ (.B1(net635),
    .Y(_2278_),
    .A1(_2270_),
    .A2(_2275_));
 sg13g2_nand2b_2 _3133_ (.Y(_2279_),
    .B(_2277_),
    .A_N(_2278_));
 sg13g2_nor2_2 _3134_ (.A(_1995_),
    .B(_2112_),
    .Y(_2280_));
 sg13g2_nor2_2 _3135_ (.A(net554),
    .B(_2210_),
    .Y(_2281_));
 sg13g2_and2_1 _3136_ (.A(_2090_),
    .B(_2136_),
    .X(_2282_));
 sg13g2_nand2_1 _3137_ (.Y(_2283_),
    .A(net556),
    .B(_2136_));
 sg13g2_nand4_1 _3138_ (.B(_2280_),
    .C(_2281_),
    .A(_2115_),
    .Y(_2284_),
    .D(_2282_));
 sg13g2_nor2_2 _3139_ (.A(net553),
    .B(_2114_),
    .Y(_2285_));
 sg13g2_nor2_1 _3140_ (.A(_2257_),
    .B(_2284_),
    .Y(_2286_));
 sg13g2_nand2_1 _3141_ (.Y(_2287_),
    .A(net574),
    .B(_2037_));
 sg13g2_nor3_1 _3142_ (.A(_1995_),
    .B(_2002_),
    .C(net567),
    .Y(_2288_));
 sg13g2_nand3_1 _3143_ (.B(net574),
    .C(net565),
    .A(_1996_),
    .Y(_2289_));
 sg13g2_nor4_2 _3144_ (.A(net573),
    .B(net554),
    .C(_2114_),
    .Y(_2290_),
    .D(_2167_));
 sg13g2_nand3_1 _3145_ (.B(_2288_),
    .C(_2290_),
    .A(_2140_),
    .Y(_2291_));
 sg13g2_nor2b_1 _3146_ (.A(_2287_),
    .B_N(_2291_),
    .Y(_2292_));
 sg13g2_a21oi_1 _3147_ (.A1(_2285_),
    .A2(_2292_),
    .Y(_2293_),
    .B1(_2153_));
 sg13g2_nand2_1 _3148_ (.Y(_2294_),
    .A(net572),
    .B(net556));
 sg13g2_and3_1 _3149_ (.X(_2295_),
    .A(net619),
    .B(net595),
    .C(net583));
 sg13g2_nand2_2 _3150_ (.Y(_2296_),
    .A(_1999_),
    .B(net584));
 sg13g2_nor3_2 _3151_ (.A(net573),
    .B(_2092_),
    .C(_2295_),
    .Y(_2297_));
 sg13g2_and4_1 _3152_ (.A(_2078_),
    .B(_2186_),
    .C(_2262_),
    .D(_2297_),
    .X(_2298_));
 sg13g2_nor2_1 _3153_ (.A(_2033_),
    .B(_2087_),
    .Y(_2299_));
 sg13g2_nor2_2 _3154_ (.A(_2042_),
    .B(net546),
    .Y(_2300_));
 sg13g2_nand2_2 _3155_ (.Y(_2301_),
    .A(net568),
    .B(net541));
 sg13g2_nand4_1 _3156_ (.B(net565),
    .C(_2047_),
    .A(net568),
    .Y(_2302_),
    .D(net541));
 sg13g2_or4_1 _3157_ (.A(_2173_),
    .B(_2199_),
    .C(_2263_),
    .D(_2302_),
    .X(_2303_));
 sg13g2_a21oi_1 _3158_ (.A1(_2246_),
    .A2(_2298_),
    .Y(_2304_),
    .B1(_2303_));
 sg13g2_nor2_1 _3159_ (.A(_2105_),
    .B(_2304_),
    .Y(_2305_));
 sg13g2_nand3_1 _3160_ (.B(_2084_),
    .C(_2088_),
    .A(net561),
    .Y(_2306_));
 sg13g2_nand2_1 _3161_ (.Y(_2307_),
    .A(net569),
    .B(net568));
 sg13g2_nor3_1 _3162_ (.A(_2029_),
    .B(_2033_),
    .C(_2160_),
    .Y(_2308_));
 sg13g2_nor2_2 _3163_ (.A(_2114_),
    .B(net548),
    .Y(_2309_));
 sg13g2_nand2_2 _3164_ (.Y(_2310_),
    .A(_2115_),
    .B(_2176_));
 sg13g2_a21oi_1 _3165_ (.A1(net606),
    .A2(_1999_),
    .Y(_2311_),
    .B1(_2141_));
 sg13g2_nand4_1 _3166_ (.B(_2308_),
    .C(_2309_),
    .A(net556),
    .Y(_2312_),
    .D(_2311_));
 sg13g2_nor2_2 _3167_ (.A(_2033_),
    .B(_2114_),
    .Y(_2313_));
 sg13g2_nand2_1 _3168_ (.Y(_2314_),
    .A(net568),
    .B(_2115_));
 sg13g2_o21ai_1 _3169_ (.B1(net654),
    .Y(_2315_),
    .A1(_2306_),
    .A2(_2312_));
 sg13g2_nand2_1 _3170_ (.Y(_2316_),
    .A(_2179_),
    .B(_2194_));
 sg13g2_nor2_1 _3171_ (.A(_2138_),
    .B(net540),
    .Y(_2317_));
 sg13g2_nor3_1 _3172_ (.A(_2017_),
    .B(_2053_),
    .C(_2256_),
    .Y(_2318_));
 sg13g2_nand2_1 _3173_ (.Y(_2319_),
    .A(_2317_),
    .B(_2318_));
 sg13g2_nor2_1 _3174_ (.A(net573),
    .B(net547),
    .Y(_2320_));
 sg13g2_nor3_1 _3175_ (.A(net573),
    .B(net552),
    .C(net546),
    .Y(_2321_));
 sg13g2_nor3_1 _3176_ (.A(_2023_),
    .B(net571),
    .C(_2046_),
    .Y(_2322_));
 sg13g2_nor4_1 _3177_ (.A(_2053_),
    .B(net559),
    .C(net555),
    .D(_2185_),
    .Y(_2323_));
 sg13g2_nand3_1 _3178_ (.B(_2322_),
    .C(_2323_),
    .A(_2321_),
    .Y(_2324_));
 sg13g2_nand2_1 _3179_ (.Y(_2325_),
    .A(net648),
    .B(_2324_));
 sg13g2_o21ai_1 _3180_ (.B1(net649),
    .Y(_2326_),
    .A1(_2098_),
    .A2(_2298_));
 sg13g2_a22oi_1 _3181_ (.Y(_2327_),
    .B1(_2319_),
    .B2(_2125_),
    .A2(_2316_),
    .A1(net647));
 sg13g2_nand3_1 _3182_ (.B(_2325_),
    .C(_2327_),
    .A(_2315_),
    .Y(_2328_));
 sg13g2_nor4_1 _3183_ (.A(_2293_),
    .B(_2305_),
    .C(_2326_),
    .D(_2328_),
    .Y(_2329_));
 sg13g2_a21oi_2 _3184_ (.B1(_2329_),
    .Y(_2330_),
    .A2(_2286_),
    .A1(net651));
 sg13g2_nor2_1 _3185_ (.A(net562),
    .B(_2135_),
    .Y(_2331_));
 sg13g2_nand2_2 _3186_ (.Y(_2332_),
    .A(_2050_),
    .B(_2136_));
 sg13g2_nor4_2 _3187_ (.A(_2160_),
    .B(net548),
    .C(_2209_),
    .Y(_2333_),
    .D(_2332_));
 sg13g2_nor3_1 _3188_ (.A(net575),
    .B(_2010_),
    .C(_2307_),
    .Y(_2334_));
 sg13g2_nand4_1 _3189_ (.B(_2088_),
    .C(_2333_),
    .A(net557),
    .Y(_2335_),
    .D(_2334_));
 sg13g2_nor2_1 _3190_ (.A(net649),
    .B(_2335_),
    .Y(_2336_));
 sg13g2_a221oi_1 _3191_ (.B2(_2290_),
    .C1(_2289_),
    .B1(_2140_),
    .A1(net620),
    .Y(_2337_),
    .A2(_2111_));
 sg13g2_nor2_1 _3192_ (.A(_2153_),
    .B(_2337_),
    .Y(_2338_));
 sg13g2_nand4_1 _3193_ (.B(net550),
    .C(_2137_),
    .A(net572),
    .Y(_2339_),
    .D(_2161_));
 sg13g2_nor4_2 _3194_ (.A(net570),
    .B(_2195_),
    .C(_2231_),
    .Y(_2340_),
    .D(_2339_));
 sg13g2_o21ai_1 _3195_ (.B1(net649),
    .Y(_2341_),
    .A1(_2126_),
    .A2(_2340_));
 sg13g2_nor3_1 _3196_ (.A(_2135_),
    .B(_2167_),
    .C(_2295_),
    .Y(_2342_));
 sg13g2_a21oi_1 _3197_ (.A1(net604),
    .A2(_2015_),
    .Y(_2343_),
    .B1(net559));
 sg13g2_nand4_1 _3198_ (.B(_2322_),
    .C(_2342_),
    .A(_2321_),
    .Y(_2344_),
    .D(_2343_));
 sg13g2_and2_1 _3199_ (.A(net648),
    .B(_2344_),
    .X(_2345_));
 sg13g2_nor3_1 _3200_ (.A(_2033_),
    .B(_2173_),
    .C(_2199_),
    .Y(_2346_));
 sg13g2_and2_1 _3201_ (.A(net543),
    .B(_2188_),
    .X(_2347_));
 sg13g2_and4_1 _3202_ (.A(_2078_),
    .B(_2297_),
    .C(_2346_),
    .D(_2347_),
    .X(_2348_));
 sg13g2_inv_1 _3203_ (.Y(_2349_),
    .A(_2348_));
 sg13g2_nor3_2 _3204_ (.A(_2033_),
    .B(_2190_),
    .C(_2199_),
    .Y(_2350_));
 sg13g2_nand3b_1 _3205_ (.B(net557),
    .C(_2161_),
    .Y(_2351_),
    .A_N(_2031_));
 sg13g2_nand3_1 _3206_ (.B(net565),
    .C(_2137_),
    .A(net574),
    .Y(_2352_));
 sg13g2_nor4_2 _3207_ (.A(_2225_),
    .B(_2266_),
    .C(_2351_),
    .Y(_2353_),
    .D(_2352_));
 sg13g2_nand2_1 _3208_ (.Y(_2354_),
    .A(_2032_),
    .B(net550));
 sg13g2_a21oi_1 _3209_ (.A1(_2350_),
    .A2(_2353_),
    .Y(_2355_),
    .B1(_2149_));
 sg13g2_nor4_1 _3210_ (.A(_2135_),
    .B(_2167_),
    .C(net548),
    .D(net540),
    .Y(_2356_));
 sg13g2_nand3_1 _3211_ (.B(_2280_),
    .C(_2356_),
    .A(_2055_),
    .Y(_2357_));
 sg13g2_or4_1 _3212_ (.A(net545),
    .B(_2306_),
    .C(_2307_),
    .D(_2357_),
    .X(_2358_));
 sg13g2_nor2_2 _3213_ (.A(net558),
    .B(_2302_),
    .Y(_2359_));
 sg13g2_nor3_1 _3214_ (.A(net592),
    .B(_2249_),
    .C(net540),
    .Y(_2360_));
 sg13g2_a21oi_1 _3215_ (.A1(_2359_),
    .A2(_2360_),
    .Y(_2361_),
    .B1(_2105_));
 sg13g2_a221oi_1 _3216_ (.B2(net654),
    .C1(_2341_),
    .B1(_2358_),
    .A1(_2097_),
    .Y(_2362_),
    .A2(_2349_));
 sg13g2_nor4_2 _3217_ (.A(_2338_),
    .B(_2345_),
    .C(_2355_),
    .Y(_2363_),
    .D(_2361_));
 sg13g2_a21oi_1 _3218_ (.A1(_2362_),
    .A2(_2363_),
    .Y(_2364_),
    .B1(_2336_));
 sg13g2_nand2_2 _3219_ (.Y(_2365_),
    .A(_2115_),
    .B(_2207_));
 sg13g2_nand3_1 _3220_ (.B(_2171_),
    .C(_2218_),
    .A(net564),
    .Y(_2366_));
 sg13g2_nor4_2 _3221_ (.A(_2012_),
    .B(_2134_),
    .C(_2365_),
    .Y(_2367_),
    .D(_2366_));
 sg13g2_and2_1 _3222_ (.A(net651),
    .B(_2367_),
    .X(_2368_));
 sg13g2_nand4_1 _3223_ (.B(net561),
    .C(_2117_),
    .A(net574),
    .Y(_2369_),
    .D(_2186_));
 sg13g2_nor4_2 _3224_ (.A(_2177_),
    .B(_2245_),
    .C(_2302_),
    .Y(_2370_),
    .D(_2369_));
 sg13g2_or2_1 _3225_ (.X(_2371_),
    .B(_2370_),
    .A(_2105_));
 sg13g2_nor2_2 _3226_ (.A(_2029_),
    .B(net558),
    .Y(_2372_));
 sg13g2_o21ai_1 _3227_ (.B1(_2047_),
    .Y(_2373_),
    .A1(_1992_),
    .A2(_2016_));
 sg13g2_nand3_1 _3228_ (.B(_2011_),
    .C(_2113_),
    .A(_1996_),
    .Y(_2374_));
 sg13g2_nor3_2 _3229_ (.A(_2023_),
    .B(net570),
    .C(net544),
    .Y(_2375_));
 sg13g2_nor3_2 _3230_ (.A(_2077_),
    .B(_2232_),
    .C(_2373_),
    .Y(_2376_));
 sg13g2_and4_1 _3231_ (.A(_2011_),
    .B(_2280_),
    .C(_2372_),
    .D(_2375_),
    .X(_2377_));
 sg13g2_a21o_1 _3232_ (.A2(_2377_),
    .A1(_2376_),
    .B1(_2130_),
    .X(_2378_));
 sg13g2_nor4_1 _3233_ (.A(_1995_),
    .B(_2017_),
    .C(_2029_),
    .D(net559),
    .Y(_2379_));
 sg13g2_nand4_1 _3234_ (.B(_2265_),
    .C(_2342_),
    .A(_2221_),
    .Y(_2380_),
    .D(_2379_));
 sg13g2_nand2_1 _3235_ (.Y(_2381_),
    .A(_2154_),
    .B(_2380_));
 sg13g2_and2_1 _3236_ (.A(net620),
    .B(net608),
    .X(_2382_));
 sg13g2_nor2_1 _3237_ (.A(_1999_),
    .B(_2015_),
    .Y(_2383_));
 sg13g2_nor4_1 _3238_ (.A(net573),
    .B(net552),
    .C(net546),
    .D(_2382_),
    .Y(_2384_));
 sg13g2_and4_1 _3239_ (.A(_2027_),
    .B(_2258_),
    .C(_2383_),
    .D(_2384_),
    .X(_2385_));
 sg13g2_a221oi_1 _3240_ (.B2(net624),
    .C1(_2046_),
    .B1(_2089_),
    .A1(_1993_),
    .Y(_2386_),
    .A2(_2015_));
 sg13g2_nand4_1 _3241_ (.B(_2250_),
    .C(_2317_),
    .A(_2021_),
    .Y(_2387_),
    .D(_2386_));
 sg13g2_o21ai_1 _3242_ (.B1(net659),
    .Y(_2388_),
    .A1(_2385_),
    .A2(_2387_));
 sg13g2_nor3_1 _3243_ (.A(_2017_),
    .B(_2031_),
    .C(_2135_),
    .Y(_2389_));
 sg13g2_nand3_1 _3244_ (.B(_2346_),
    .C(_2389_),
    .A(_2288_),
    .Y(_2390_));
 sg13g2_nor2_1 _3245_ (.A(_2077_),
    .B(_2173_),
    .Y(_2391_));
 sg13g2_nor4_1 _3246_ (.A(net567),
    .B(_2042_),
    .C(_2044_),
    .D(net559),
    .Y(_2392_));
 sg13g2_nor3_1 _3247_ (.A(_2002_),
    .B(net563),
    .C(_2170_),
    .Y(_2393_));
 sg13g2_nor3_2 _3248_ (.A(_2023_),
    .B(_2080_),
    .C(net552),
    .Y(_2394_));
 sg13g2_nand4_1 _3249_ (.B(_2392_),
    .C(_2393_),
    .A(_2297_),
    .Y(_2395_),
    .D(_2394_));
 sg13g2_a22oi_1 _3250_ (.Y(_2396_),
    .B1(_2395_),
    .B2(net663),
    .A2(_2390_),
    .A1(net647));
 sg13g2_nand4_1 _3251_ (.B(net550),
    .C(net543),
    .A(_2085_),
    .Y(_2397_),
    .D(_2311_));
 sg13g2_o21ai_1 _3252_ (.B1(net654),
    .Y(_2398_),
    .A1(_2357_),
    .A2(_2397_));
 sg13g2_and3_1 _3253_ (.X(_2399_),
    .A(_2381_),
    .B(_2396_),
    .C(_2398_));
 sg13g2_and4_1 _3254_ (.A(_2073_),
    .B(_2371_),
    .C(_2378_),
    .D(_2388_),
    .X(_2400_));
 sg13g2_a22oi_1 _3255_ (.Y(_2401_),
    .B1(_2399_),
    .B2(_2400_),
    .A2(_2367_),
    .A1(net651));
 sg13g2_a21o_1 _3256_ (.A2(_2400_),
    .A1(_2399_),
    .B1(_2368_),
    .X(_2402_));
 sg13g2_a221oi_1 _3257_ (.B2(_2157_),
    .C1(_2336_),
    .B1(_2402_),
    .A1(_2362_),
    .Y(_2403_),
    .A2(_2363_));
 sg13g2_nor3_1 _3258_ (.A(_2275_),
    .B(_2330_),
    .C(_2403_),
    .Y(_2404_));
 sg13g2_mux2_2 _3259_ (.A0(_2364_),
    .A1(_2404_),
    .S(net639),
    .X(_2405_));
 sg13g2_a21oi_1 _3260_ (.A1(_2285_),
    .A2(_2292_),
    .Y(_2406_),
    .B1(net661));
 sg13g2_nor2_1 _3261_ (.A(_2129_),
    .B(_2304_),
    .Y(_2407_));
 sg13g2_a22oi_1 _3262_ (.Y(_2408_),
    .B1(_2324_),
    .B2(_2061_),
    .A2(_2319_),
    .A1(_2071_));
 sg13g2_o21ai_1 _3263_ (.B1(_2408_),
    .Y(_2409_),
    .A1(_2243_),
    .A2(_2298_));
 sg13g2_o21ai_1 _3264_ (.B1(net656),
    .Y(_2410_),
    .A1(_2306_),
    .A2(_2312_));
 sg13g2_nand2_1 _3265_ (.Y(_2411_),
    .A(_2255_),
    .B(_2316_));
 sg13g2_o21ai_1 _3266_ (.B1(_2102_),
    .Y(_2412_),
    .A1(_2257_),
    .A2(_2284_));
 sg13g2_nand3_1 _3267_ (.B(_2411_),
    .C(_2412_),
    .A(_2410_),
    .Y(_2413_));
 sg13g2_nor4_2 _3268_ (.A(_2406_),
    .B(_2407_),
    .C(_2409_),
    .Y(_2414_),
    .D(_2413_));
 sg13g2_nor2_1 _3269_ (.A(net661),
    .B(_2337_),
    .Y(_2415_));
 sg13g2_a21o_1 _3270_ (.A2(_2360_),
    .A1(_2359_),
    .B1(_2129_),
    .X(_2416_));
 sg13g2_nor2_1 _3271_ (.A(_2070_),
    .B(_2340_),
    .Y(_2417_));
 sg13g2_and2_1 _3272_ (.A(_2061_),
    .B(_2344_),
    .X(_2418_));
 sg13g2_a22oi_1 _3273_ (.Y(_2419_),
    .B1(_2358_),
    .B2(net656),
    .A2(_2335_),
    .A1(_2102_));
 sg13g2_a21oi_1 _3274_ (.A1(_2350_),
    .A2(_2353_),
    .Y(_2420_),
    .B1(_2254_));
 sg13g2_nand2_1 _3275_ (.Y(_2421_),
    .A(_2244_),
    .B(_2349_));
 sg13g2_nor4_1 _3276_ (.A(_2415_),
    .B(_2417_),
    .C(_2418_),
    .D(_2420_),
    .Y(_2422_));
 sg13g2_and4_2 _3277_ (.A(_2416_),
    .B(_2419_),
    .C(_2421_),
    .D(_2422_),
    .X(_2423_));
 sg13g2_nand2_1 _3278_ (.Y(_2424_),
    .A(_2103_),
    .B(_2151_));
 sg13g2_nand2_1 _3279_ (.Y(_2425_),
    .A(net662),
    .B(_2254_));
 sg13g2_a22oi_1 _3280_ (.Y(_2426_),
    .B1(_2118_),
    .B2(_2119_),
    .A2(_2070_),
    .A1(_2062_));
 sg13g2_nand2_1 _3281_ (.Y(_2427_),
    .A(_2129_),
    .B(_2243_));
 sg13g2_a21o_1 _3282_ (.A2(_2427_),
    .A1(_2094_),
    .B1(_2426_),
    .X(_2428_));
 sg13g2_a221oi_1 _3283_ (.B2(_2147_),
    .C1(_2428_),
    .B1(_2425_),
    .A1(_2057_),
    .Y(_2429_),
    .A2(_2424_));
 sg13g2_a21oi_1 _3284_ (.A1(_2376_),
    .A2(_2377_),
    .Y(_2430_),
    .B1(_2062_));
 sg13g2_nor2_1 _3285_ (.A(net660),
    .B(_2367_),
    .Y(_2431_));
 sg13g2_nor2_1 _3286_ (.A(_2129_),
    .B(_2370_),
    .Y(_2432_));
 sg13g2_nor3_1 _3287_ (.A(_2430_),
    .B(_2431_),
    .C(_2432_),
    .Y(_2433_));
 sg13g2_o21ai_1 _3288_ (.B1(_2071_),
    .Y(_2434_),
    .A1(_2385_),
    .A2(_2387_));
 sg13g2_a22oi_1 _3289_ (.Y(_2435_),
    .B1(_2390_),
    .B2(_2255_),
    .A2(_2380_),
    .A1(_2099_));
 sg13g2_o21ai_1 _3290_ (.B1(net656),
    .Y(_2436_),
    .A1(_2357_),
    .A2(_2397_));
 sg13g2_nand2_1 _3291_ (.Y(_2437_),
    .A(_2244_),
    .B(_2395_));
 sg13g2_and4_1 _3292_ (.A(_2434_),
    .B(_2435_),
    .C(_2436_),
    .D(_2437_),
    .X(_2438_));
 sg13g2_and2_1 _3293_ (.A(_2433_),
    .B(_2438_),
    .X(_2439_));
 sg13g2_and3_1 _3294_ (.X(_2440_),
    .A(_2429_),
    .B(_2433_),
    .C(_2438_));
 sg13g2_o21ai_1 _3295_ (.B1(_2414_),
    .Y(_2441_),
    .A1(_2423_),
    .A2(_2440_));
 sg13g2_o21ai_1 _3296_ (.B1(net640),
    .Y(_2442_),
    .A1(_2270_),
    .A2(_2441_));
 sg13g2_nand2_1 _3297_ (.Y(_2443_),
    .A(net635),
    .B(_2423_));
 sg13g2_nand2_2 _3298_ (.Y(_2444_),
    .A(_2442_),
    .B(_2443_));
 sg13g2_nor2_1 _3299_ (.A(_2405_),
    .B(_2444_),
    .Y(_2445_));
 sg13g2_nand2_1 _3300_ (.Y(_2446_),
    .A(_2414_),
    .B(_2442_));
 sg13g2_nor2_1 _3301_ (.A(net640),
    .B(_2330_),
    .Y(_2447_));
 sg13g2_nor2_1 _3302_ (.A(_2404_),
    .B(_2447_),
    .Y(_2448_));
 sg13g2_nor2b_1 _3303_ (.A(_2448_),
    .B_N(_2446_),
    .Y(_2449_));
 sg13g2_nand2b_1 _3304_ (.Y(_2450_),
    .B(_2448_),
    .A_N(_2446_));
 sg13g2_xor2_1 _3305_ (.B(_2444_),
    .A(_2405_),
    .X(_2451_));
 sg13g2_nand3b_1 _3306_ (.B(_2450_),
    .C(_2451_),
    .Y(_2452_),
    .A_N(_2449_));
 sg13g2_nor2_1 _3307_ (.A(net641),
    .B(_2402_),
    .Y(_2453_));
 sg13g2_xor2_1 _3308_ (.B(_2403_),
    .A(_2330_),
    .X(_2454_));
 sg13g2_xnor2_1 _3309_ (.Y(_2455_),
    .A(_2330_),
    .B(_2403_));
 sg13g2_nor2_1 _3310_ (.A(net639),
    .B(_2401_),
    .Y(_2456_));
 sg13g2_a21oi_2 _3311_ (.B1(_2453_),
    .Y(_2457_),
    .A2(_2455_),
    .A1(net639));
 sg13g2_or2_1 _3312_ (.X(_2458_),
    .B(_2439_),
    .A(net639));
 sg13g2_or3_1 _3313_ (.A(_2414_),
    .B(_2423_),
    .C(_2440_),
    .X(_2459_));
 sg13g2_a21o_1 _3314_ (.A2(_2459_),
    .A1(_2441_),
    .B1(net635),
    .X(_2460_));
 sg13g2_nand2_1 _3315_ (.Y(_2461_),
    .A(net636),
    .B(_2439_));
 sg13g2_nand3_1 _3316_ (.B(_2441_),
    .C(_2459_),
    .A(net640),
    .Y(_2462_));
 sg13g2_nand2_1 _3317_ (.Y(_2463_),
    .A(_2461_),
    .B(_2462_));
 sg13g2_a221oi_1 _3318_ (.B2(_2462_),
    .C1(_2456_),
    .B1(_2461_),
    .A1(net639),
    .Y(_2464_),
    .A2(_2454_));
 sg13g2_nand2b_1 _3319_ (.Y(_2465_),
    .B(_2463_),
    .A_N(_2457_));
 sg13g2_a221oi_1 _3320_ (.B2(_2460_),
    .C1(_2453_),
    .B1(_2458_),
    .A1(net640),
    .Y(_2466_),
    .A2(_2455_));
 sg13g2_nor3_1 _3321_ (.A(net635),
    .B(_2423_),
    .C(_2440_),
    .Y(_2467_));
 sg13g2_a21o_1 _3322_ (.A2(_2439_),
    .A1(_2423_),
    .B1(net635),
    .X(_2468_));
 sg13g2_a21o_2 _3323_ (.A2(_2468_),
    .A1(_2429_),
    .B1(_2467_),
    .X(_2469_));
 sg13g2_and2_1 _3324_ (.A(net639),
    .B(_2403_),
    .X(_2470_));
 sg13g2_o21ai_1 _3325_ (.B1(net639),
    .Y(_2471_),
    .A1(_2364_),
    .A2(_2401_));
 sg13g2_a22oi_1 _3326_ (.Y(_2472_),
    .B1(_2471_),
    .B2(_2157_),
    .A2(_2403_),
    .A1(net639));
 sg13g2_a21o_1 _3327_ (.A2(_2471_),
    .A1(_2157_),
    .B1(_2470_),
    .X(_2473_));
 sg13g2_nor2_1 _3328_ (.A(_2469_),
    .B(_2472_),
    .Y(_2474_));
 sg13g2_xnor2_1 _3329_ (.Y(_2475_),
    .A(_2469_),
    .B(_2472_));
 sg13g2_nor3_1 _3330_ (.A(_2464_),
    .B(_2466_),
    .C(_2475_),
    .Y(_2476_));
 sg13g2_or3_1 _3331_ (.A(_2464_),
    .B(_2466_),
    .C(_2475_),
    .X(_2477_));
 sg13g2_a21oi_1 _3332_ (.A1(_2433_),
    .A2(_2438_),
    .Y(_2478_),
    .B1(_2429_));
 sg13g2_nor3_1 _3333_ (.A(net635),
    .B(_2440_),
    .C(_2478_),
    .Y(_2479_));
 sg13g2_nor2_2 _3334_ (.A(net555),
    .B(_2210_),
    .Y(_2480_));
 sg13g2_nor3_1 _3335_ (.A(_2017_),
    .B(net558),
    .C(_2263_),
    .Y(_2481_));
 sg13g2_nand4_1 _3336_ (.B(_2350_),
    .C(_2480_),
    .A(_2194_),
    .Y(_2482_),
    .D(_2481_));
 sg13g2_nand2_1 _3337_ (.Y(_2483_),
    .A(_2255_),
    .B(_2482_));
 sg13g2_o21ai_1 _3338_ (.B1(_2483_),
    .Y(_2484_),
    .A1(net661),
    .A2(_2482_));
 sg13g2_nand2_2 _3339_ (.Y(_2485_),
    .A(_2207_),
    .B(_2296_));
 sg13g2_nand4_1 _3340_ (.B(net557),
    .C(_2207_),
    .A(net574),
    .Y(_2486_),
    .D(_2296_));
 sg13g2_nand3_1 _3341_ (.B(_2022_),
    .C(_2172_),
    .A(net572),
    .Y(_2487_));
 sg13g2_or4_2 _3342_ (.A(_2199_),
    .B(_2382_),
    .C(_2486_),
    .D(_2487_),
    .X(_2488_));
 sg13g2_nand2_1 _3343_ (.Y(_2489_),
    .A(_2244_),
    .B(_2488_));
 sg13g2_o21ai_1 _3344_ (.B1(_2489_),
    .Y(_2490_),
    .A1(_2129_),
    .A2(_2488_));
 sg13g2_nor2_1 _3345_ (.A(_2044_),
    .B(_2206_),
    .Y(_2491_));
 sg13g2_nand2_2 _3346_ (.Y(_2492_),
    .A(net564),
    .B(_2491_));
 sg13g2_and2_2 _3347_ (.A(net599),
    .B(_2015_),
    .X(_2493_));
 sg13g2_nand4_1 _3348_ (.B(_2083_),
    .C(_2267_),
    .A(_2021_),
    .Y(_2494_),
    .D(_2281_));
 sg13g2_nor4_2 _3349_ (.A(net562),
    .B(_2492_),
    .C(_2493_),
    .Y(_2495_),
    .D(_2494_));
 sg13g2_nand2_1 _3350_ (.Y(_2496_),
    .A(_2055_),
    .B(_2142_));
 sg13g2_nor2_1 _3351_ (.A(net571),
    .B(net540),
    .Y(_2497_));
 sg13g2_nand2_2 _3352_ (.Y(_2498_),
    .A(_1996_),
    .B(net557));
 sg13g2_nand4_1 _3353_ (.B(net565),
    .C(_2267_),
    .A(_2001_),
    .Y(_2499_),
    .D(_2497_));
 sg13g2_nor3_2 _3354_ (.A(_2496_),
    .B(_2498_),
    .C(_2499_),
    .Y(_2500_));
 sg13g2_mux2_1 _3355_ (.A0(net652),
    .A1(_2061_),
    .S(_2500_),
    .X(_2501_));
 sg13g2_a21o_1 _3356_ (.A2(_2495_),
    .A1(_2150_),
    .B1(_2501_),
    .X(_2502_));
 sg13g2_o21ai_1 _3357_ (.B1(net634),
    .Y(_2503_),
    .A1(net660),
    .A2(_2495_));
 sg13g2_nor4_1 _3358_ (.A(_2484_),
    .B(_2490_),
    .C(_2502_),
    .D(_2503_),
    .Y(_2504_));
 sg13g2_nor2_1 _3359_ (.A(_2479_),
    .B(_2504_),
    .Y(_2505_));
 sg13g2_inv_1 _3360_ (.Y(_2506_),
    .A(_2505_));
 sg13g2_xnor2_1 _3361_ (.Y(_2507_),
    .A(_2158_),
    .B(_2401_));
 sg13g2_nand2_1 _3362_ (.Y(_2508_),
    .A(net663),
    .B(_2488_));
 sg13g2_nand2_1 _3363_ (.Y(_2509_),
    .A(net647),
    .B(_2482_));
 sg13g2_o21ai_1 _3364_ (.B1(_2509_),
    .Y(_2510_),
    .A1(_2153_),
    .A2(_2482_));
 sg13g2_nor2_1 _3365_ (.A(_2126_),
    .B(_2500_),
    .Y(_2511_));
 sg13g2_a22oi_1 _3366_ (.Y(_2512_),
    .B1(_2500_),
    .B2(_2131_),
    .A2(_2495_),
    .A1(net654));
 sg13g2_nand2_1 _3367_ (.Y(_2513_),
    .A(_2508_),
    .B(_2512_));
 sg13g2_o21ai_1 _3368_ (.B1(net649),
    .Y(_2514_),
    .A1(_2105_),
    .A2(_2488_));
 sg13g2_or4_1 _3369_ (.A(_2510_),
    .B(_2511_),
    .C(_2513_),
    .D(_2514_),
    .X(_2515_));
 sg13g2_a21oi_1 _3370_ (.A1(net651),
    .A2(_2495_),
    .Y(_2516_),
    .B1(net638));
 sg13g2_a22oi_1 _3371_ (.Y(_2517_),
    .B1(_2515_),
    .B2(_2516_),
    .A2(_2507_),
    .A1(net638));
 sg13g2_nand2_1 _3372_ (.Y(_2518_),
    .A(_2505_),
    .B(_2517_));
 sg13g2_nor2_1 _3373_ (.A(net634),
    .B(_2429_),
    .Y(_2519_));
 sg13g2_nor2_1 _3374_ (.A(_2213_),
    .B(_2243_),
    .Y(_2520_));
 sg13g2_o21ai_1 _3375_ (.B1(net655),
    .Y(_2521_),
    .A1(net544),
    .A2(_2192_));
 sg13g2_nand2_1 _3376_ (.Y(_2522_),
    .A(_2061_),
    .B(_2203_));
 sg13g2_nor2_1 _3377_ (.A(net660),
    .B(_2192_),
    .Y(_2523_));
 sg13g2_a21oi_1 _3378_ (.A1(net657),
    .A2(_2212_),
    .Y(_2524_),
    .B1(_2523_));
 sg13g2_o21ai_1 _3379_ (.B1(_2524_),
    .Y(_2525_),
    .A1(net661),
    .A2(_2227_));
 sg13g2_a22oi_1 _3380_ (.Y(_2526_),
    .B1(_2255_),
    .B2(_2220_),
    .A2(_2235_),
    .A1(net652));
 sg13g2_nand3_1 _3381_ (.B(_2522_),
    .C(_2526_),
    .A(_2521_),
    .Y(_2527_));
 sg13g2_nor4_2 _3382_ (.A(net637),
    .B(_2520_),
    .C(_2525_),
    .Y(_2528_),
    .D(_2527_));
 sg13g2_nor2_2 _3383_ (.A(_2519_),
    .B(_2528_),
    .Y(_2529_));
 sg13g2_nor2b_1 _3384_ (.A(_2529_),
    .B_N(_2242_),
    .Y(_2530_));
 sg13g2_xnor2_1 _3385_ (.Y(_2531_),
    .A(_2505_),
    .B(_2517_));
 sg13g2_nor2_1 _3386_ (.A(_2530_),
    .B(_2531_),
    .Y(_2532_));
 sg13g2_o21ai_1 _3387_ (.B1(_2518_),
    .Y(_2533_),
    .A1(_2530_),
    .A2(_2531_));
 sg13g2_a221oi_1 _3388_ (.B2(_2533_),
    .C1(_2466_),
    .B1(_2476_),
    .A1(_2465_),
    .Y(_2534_),
    .A2(_2474_));
 sg13g2_a21oi_1 _3389_ (.A1(_2445_),
    .A2(_2450_),
    .Y(_2535_),
    .B1(_2449_));
 sg13g2_o21ai_1 _3390_ (.B1(_2535_),
    .Y(_2536_),
    .A1(_2452_),
    .A2(_2534_));
 sg13g2_a21oi_2 _3391_ (.B1(_2276_),
    .Y(_2537_),
    .A2(_2536_),
    .A1(_2279_));
 sg13g2_a21o_1 _3392_ (.A2(_2536_),
    .A1(_2279_),
    .B1(_2276_),
    .X(_2538_));
 sg13g2_nand2b_1 _3393_ (.Y(_2539_),
    .B(_2529_),
    .A_N(_2242_));
 sg13g2_nand3_1 _3394_ (.B(_2532_),
    .C(_2539_),
    .A(_2279_),
    .Y(_2540_));
 sg13g2_nor3_2 _3395_ (.A(_2452_),
    .B(_2477_),
    .C(_2540_),
    .Y(_2541_));
 sg13g2_or3_1 _3396_ (.A(_2452_),
    .B(_2477_),
    .C(_2540_),
    .X(_2542_));
 sg13g2_nand2_1 _3397_ (.Y(_2543_),
    .A(_2538_),
    .B(_2542_));
 sg13g2_mux2_1 _3398_ (.A0(_2529_),
    .A1(_2242_),
    .S(net537),
    .X(_2544_));
 sg13g2_nand2_1 _3399_ (.Y(_2545_),
    .A(_0059_),
    .B(_2544_));
 sg13g2_nor2_1 _3400_ (.A(net144),
    .B(_2544_),
    .Y(_2546_));
 sg13g2_xnor2_1 _3401_ (.Y(_0074_),
    .A(net144),
    .B(_2544_));
 sg13g2_nor3_1 _3402_ (.A(_2242_),
    .B(_2537_),
    .C(_2541_),
    .Y(_2547_));
 sg13g2_a21o_1 _3403_ (.A2(net539),
    .A1(net538),
    .B1(_2529_),
    .X(_0153_));
 sg13g2_nor2b_1 _3404_ (.A(_2547_),
    .B_N(_0153_),
    .Y(_0154_));
 sg13g2_nand3b_1 _3405_ (.B(_0153_),
    .C(net165),
    .Y(_0155_),
    .A_N(_2547_));
 sg13g2_xnor2_1 _3406_ (.Y(_0081_),
    .A(net144),
    .B(_0154_));
 sg13g2_nor3_2 _3407_ (.A(_2033_),
    .B(_2135_),
    .C(_2210_),
    .Y(_0156_));
 sg13g2_nand3_1 _3408_ (.B(_2176_),
    .C(_0156_),
    .A(_2009_),
    .Y(_0157_));
 sg13g2_nand2_1 _3409_ (.Y(_0158_),
    .A(_2116_),
    .B(_2375_));
 sg13g2_or3_1 _3410_ (.A(_2486_),
    .B(_0157_),
    .C(_0158_),
    .X(_0159_));
 sg13g2_nor2_2 _3411_ (.A(_2018_),
    .B(_2120_),
    .Y(_0160_));
 sg13g2_nor2_2 _3412_ (.A(_2007_),
    .B(net583),
    .Y(_0161_));
 sg13g2_nor3_1 _3413_ (.A(net572),
    .B(net585),
    .C(net581),
    .Y(_0162_));
 sg13g2_nor3_2 _3414_ (.A(_2018_),
    .B(net552),
    .C(_0162_),
    .Y(_0163_));
 sg13g2_nor2_2 _3415_ (.A(net554),
    .B(_2162_),
    .Y(_0164_));
 sg13g2_and3_1 _3416_ (.X(_0165_),
    .A(_2022_),
    .B(_2171_),
    .C(_2207_));
 sg13g2_nor4_1 _3417_ (.A(net562),
    .B(_2053_),
    .C(_2112_),
    .D(_2114_),
    .Y(_0166_));
 sg13g2_nand4_1 _3418_ (.B(_0164_),
    .C(_0165_),
    .A(_0163_),
    .Y(_0167_),
    .D(_0166_));
 sg13g2_and2_1 _3419_ (.A(_2106_),
    .B(_0167_),
    .X(_0168_));
 sg13g2_nor4_2 _3420_ (.A(net562),
    .B(_2075_),
    .C(net548),
    .Y(_0169_),
    .D(_2493_));
 sg13g2_nand2_2 _3421_ (.Y(_0170_),
    .A(net557),
    .B(net542));
 sg13g2_a21oi_1 _3422_ (.A1(net608),
    .A2(net602),
    .Y(_0171_),
    .B1(_0170_));
 sg13g2_and3_1 _3423_ (.X(_0172_),
    .A(_2055_),
    .B(_2142_),
    .C(_2491_));
 sg13g2_nand4_1 _3424_ (.B(_0169_),
    .C(_0171_),
    .A(_2200_),
    .Y(_0173_),
    .D(_0172_));
 sg13g2_a221oi_1 _3425_ (.B2(_2154_),
    .C1(_0168_),
    .B1(_0173_),
    .A1(net663),
    .Y(_0174_),
    .A2(_0159_));
 sg13g2_nor2_2 _3426_ (.A(_2038_),
    .B(net540),
    .Y(_0175_));
 sg13g2_nand2_1 _3427_ (.Y(_0176_),
    .A(_2039_),
    .B(_2296_));
 sg13g2_and4_1 _3428_ (.A(_2043_),
    .B(_2115_),
    .C(_2117_),
    .D(_2480_),
    .X(_0177_));
 sg13g2_nand4_1 _3429_ (.B(_0169_),
    .C(_0175_),
    .A(net569),
    .Y(_0178_),
    .D(_0177_));
 sg13g2_nor2_1 _3430_ (.A(_2215_),
    .B(_2365_),
    .Y(_0179_));
 sg13g2_nand2_2 _3431_ (.Y(_0180_),
    .A(net569),
    .B(net560));
 sg13g2_nor3_1 _3432_ (.A(_2041_),
    .B(_2210_),
    .C(_0180_),
    .Y(_0181_));
 sg13g2_nand4_1 _3433_ (.B(_2386_),
    .C(_0179_),
    .A(net541),
    .Y(_0182_),
    .D(_0181_));
 sg13g2_nor4_2 _3434_ (.A(_2038_),
    .B(_2048_),
    .C(_2195_),
    .Y(_0183_),
    .D(_2232_));
 sg13g2_nor2_2 _3435_ (.A(net575),
    .B(_2210_),
    .Y(_0184_));
 sg13g2_nor3_1 _3436_ (.A(net570),
    .B(_2138_),
    .C(_2301_),
    .Y(_0185_));
 sg13g2_nand4_1 _3437_ (.B(_0183_),
    .C(_0184_),
    .A(net569),
    .Y(_0186_),
    .D(_0185_));
 sg13g2_nand2_1 _3438_ (.Y(_0187_),
    .A(net659),
    .B(_0186_));
 sg13g2_nor2_1 _3439_ (.A(_2195_),
    .B(_2310_),
    .Y(_0188_));
 sg13g2_nand2_1 _3440_ (.Y(_0189_),
    .A(_2047_),
    .B(net560));
 sg13g2_nor4_1 _3441_ (.A(_2008_),
    .B(net553),
    .C(_2112_),
    .D(_2164_),
    .Y(_0190_));
 sg13g2_nand4_1 _3442_ (.B(_2027_),
    .C(_2309_),
    .A(_2016_),
    .Y(_0191_),
    .D(_0190_));
 sg13g2_nor2_1 _3443_ (.A(_0189_),
    .B(_0191_),
    .Y(_0192_));
 sg13g2_o21ai_1 _3444_ (.B1(net648),
    .Y(_0193_),
    .A1(_0189_),
    .A2(_0191_));
 sg13g2_nand3_1 _3445_ (.B(_0187_),
    .C(_0193_),
    .A(net649),
    .Y(_0194_));
 sg13g2_a221oi_1 _3446_ (.B2(net653),
    .C1(_0194_),
    .B1(_0182_),
    .A1(net647),
    .Y(_0195_),
    .A2(_0178_));
 sg13g2_nor4_1 _3447_ (.A(_2038_),
    .B(_2167_),
    .C(_2493_),
    .D(_0180_),
    .Y(_0196_));
 sg13g2_and4_2 _3448_ (.A(_2045_),
    .B(_2265_),
    .C(_0164_),
    .D(_0196_),
    .X(_0197_));
 sg13g2_a22oi_1 _3449_ (.Y(_0198_),
    .B1(_0197_),
    .B2(net650),
    .A2(_0195_),
    .A1(_0174_));
 sg13g2_nor2_1 _3450_ (.A(_2010_),
    .B(_2044_),
    .Y(_0199_));
 sg13g2_nand3_1 _3451_ (.B(_0183_),
    .C(_0199_),
    .A(_0160_),
    .Y(_0200_));
 sg13g2_nor4_1 _3452_ (.A(_2042_),
    .B(_2173_),
    .C(_2498_),
    .D(_0200_),
    .Y(_0201_));
 sg13g2_nor2_1 _3453_ (.A(_2126_),
    .B(_0201_),
    .Y(_0202_));
 sg13g2_nor3_1 _3454_ (.A(_2042_),
    .B(_2146_),
    .C(_2206_),
    .Y(_0203_));
 sg13g2_nand3_1 _3455_ (.B(_2145_),
    .C(_2207_),
    .A(_2043_),
    .Y(_0204_));
 sg13g2_nor3_2 _3456_ (.A(net570),
    .B(_2138_),
    .C(_2187_),
    .Y(_0205_));
 sg13g2_nor4_1 _3457_ (.A(_2023_),
    .B(_2075_),
    .C(net558),
    .D(net548),
    .Y(_0206_));
 sg13g2_nand4_1 _3458_ (.B(_2247_),
    .C(_0205_),
    .A(_2218_),
    .Y(_0207_),
    .D(_0206_));
 sg13g2_nor3_1 _3459_ (.A(net555),
    .B(_0204_),
    .C(_0207_),
    .Y(_0208_));
 sg13g2_inv_1 _3460_ (.Y(_0209_),
    .A(_0208_));
 sg13g2_nand2_2 _3461_ (.Y(_0210_),
    .A(_1996_),
    .B(_2166_));
 sg13g2_nor3_1 _3462_ (.A(net563),
    .B(_2146_),
    .C(_2485_),
    .Y(_0211_));
 sg13g2_nand3_1 _3463_ (.B(_2386_),
    .C(_0211_),
    .A(_2166_),
    .Y(_0212_));
 sg13g2_or2_1 _3464_ (.X(_0213_),
    .B(_0212_),
    .A(_0157_));
 sg13g2_a221oi_1 _3465_ (.B2(_2106_),
    .C1(_0202_),
    .B1(_0213_),
    .A1(net647),
    .Y(_0214_),
    .A2(_0209_));
 sg13g2_nand3_1 _3466_ (.B(_2022_),
    .C(_2084_),
    .A(_2021_),
    .Y(_0215_));
 sg13g2_nor3_2 _3467_ (.A(_2214_),
    .B(_2287_),
    .C(_0215_),
    .Y(_0216_));
 sg13g2_and2_1 _3468_ (.A(_2230_),
    .B(_0216_),
    .X(_0217_));
 sg13g2_nor4_1 _3469_ (.A(_2143_),
    .B(_2169_),
    .C(_2493_),
    .D(_0176_),
    .Y(_0218_));
 sg13g2_nand4_1 _3470_ (.B(net561),
    .C(_2267_),
    .A(_2045_),
    .Y(_0219_),
    .D(_0218_));
 sg13g2_nand3_1 _3471_ (.B(_2027_),
    .C(_2040_),
    .A(_1996_),
    .Y(_0220_));
 sg13g2_nand4_1 _3472_ (.B(_2115_),
    .C(net550),
    .A(_2032_),
    .Y(_0221_),
    .D(_2296_));
 sg13g2_or4_1 _3473_ (.A(_2162_),
    .B(_2493_),
    .C(_0220_),
    .D(_0221_),
    .X(_0222_));
 sg13g2_a22oi_1 _3474_ (.Y(_0223_),
    .B1(_0222_),
    .B2(net653),
    .A2(_0219_),
    .A1(_2154_));
 sg13g2_o21ai_1 _3475_ (.B1(_0223_),
    .Y(_0224_),
    .A1(_2098_),
    .A2(_0217_));
 sg13g2_o21ai_1 _3476_ (.B1(_2207_),
    .Y(_0225_),
    .A1(net604),
    .A2(_2000_));
 sg13g2_or2_2 _3477_ (.X(_0226_),
    .B(_0225_),
    .A(_2215_));
 sg13g2_nor4_2 _3478_ (.A(_2053_),
    .B(net548),
    .C(_2185_),
    .Y(_0227_),
    .D(_2217_));
 sg13g2_nor2_1 _3479_ (.A(net555),
    .B(_2141_),
    .Y(_0228_));
 sg13g2_and4_1 _3480_ (.A(_2168_),
    .B(_2179_),
    .C(_2189_),
    .D(_0228_),
    .X(_0229_));
 sg13g2_nand3b_1 _3481_ (.B(_0227_),
    .C(_0229_),
    .Y(_0230_),
    .A_N(_0226_));
 sg13g2_nor4_1 _3482_ (.A(net570),
    .B(_2248_),
    .C(net540),
    .D(_0180_),
    .Y(_0231_));
 sg13g2_nand4_1 _3483_ (.B(_2309_),
    .C(_0184_),
    .A(_2137_),
    .Y(_0232_),
    .D(_0231_));
 sg13g2_a221oi_1 _3484_ (.B2(net648),
    .C1(net637),
    .B1(_0232_),
    .A1(net650),
    .Y(_0233_),
    .A2(_0230_));
 sg13g2_nor2b_1 _3485_ (.A(_0224_),
    .B_N(_0233_),
    .Y(_0234_));
 sg13g2_a22oi_1 _3486_ (.Y(_0235_),
    .B1(_0214_),
    .B2(_0234_),
    .A2(_0198_),
    .A1(net637));
 sg13g2_nand2_1 _3487_ (.Y(_0236_),
    .A(net656),
    .B(_0182_));
 sg13g2_nand2_1 _3488_ (.Y(_0237_),
    .A(net652),
    .B(_0186_));
 sg13g2_o21ai_1 _3489_ (.B1(_0237_),
    .Y(_0238_),
    .A1(net660),
    .A2(_0197_));
 sg13g2_a22oi_1 _3490_ (.Y(_0239_),
    .B1(_0178_),
    .B2(_2255_),
    .A2(_0159_),
    .A1(_2244_));
 sg13g2_nand2_1 _3491_ (.Y(_0240_),
    .A(_0236_),
    .B(_0239_));
 sg13g2_a22oi_1 _3492_ (.Y(_0241_),
    .B1(_0173_),
    .B2(_2099_),
    .A2(_0167_),
    .A1(net657));
 sg13g2_o21ai_1 _3493_ (.B1(_0241_),
    .Y(_0242_),
    .A1(_2062_),
    .A2(_0192_));
 sg13g2_nor3_2 _3494_ (.A(_0238_),
    .B(_0240_),
    .C(_0242_),
    .Y(_0243_));
 sg13g2_or2_1 _3495_ (.X(_0244_),
    .B(_0201_),
    .A(_2070_));
 sg13g2_a22oi_1 _3496_ (.Y(_0245_),
    .B1(_0222_),
    .B2(net655),
    .A2(_0213_),
    .A1(net657));
 sg13g2_a22oi_1 _3497_ (.Y(_0246_),
    .B1(_0232_),
    .B2(_2061_),
    .A2(_0230_),
    .A1(_2102_));
 sg13g2_o21ai_1 _3498_ (.B1(_0246_),
    .Y(_0247_),
    .A1(_2243_),
    .A2(_0217_));
 sg13g2_a221oi_1 _3499_ (.B2(_2099_),
    .C1(_0247_),
    .B1(_0219_),
    .A1(_2255_),
    .Y(_0248_),
    .A2(_0209_));
 sg13g2_nand3_1 _3500_ (.B(_0245_),
    .C(_0248_),
    .A(_0244_),
    .Y(_0249_));
 sg13g2_mux2_1 _3501_ (.A0(_0243_),
    .A1(_0249_),
    .S(net632),
    .X(_0250_));
 sg13g2_mux2_1 _3502_ (.A0(_0235_),
    .A1(_0250_),
    .S(net534),
    .X(_0251_));
 sg13g2_nand2_1 _3503_ (.Y(_0252_),
    .A(net182),
    .B(_0251_));
 sg13g2_or2_1 _3504_ (.X(_0253_),
    .B(_0251_),
    .A(net182));
 sg13g2_nand2_1 _3505_ (.Y(_0028_),
    .A(_0252_),
    .B(_0253_));
 sg13g2_mux2_2 _3506_ (.A0(_0250_),
    .A1(_0235_),
    .S(net537),
    .X(_0254_));
 sg13g2_nand2_1 _3507_ (.Y(_0255_),
    .A(net182),
    .B(_0254_));
 sg13g2_nor2_1 _3508_ (.A(_0058_),
    .B(_0254_),
    .Y(_0256_));
 sg13g2_or2_1 _3509_ (.X(_0257_),
    .B(_0254_),
    .A(net185));
 sg13g2_nand2_1 _3510_ (.Y(_0035_),
    .A(_0255_),
    .B(_0257_));
 sg13g2_nor2_2 _3511_ (.A(_2042_),
    .B(net549),
    .Y(_0258_));
 sg13g2_nand2_2 _3512_ (.Y(_0259_),
    .A(_2372_),
    .B(_0258_));
 sg13g2_nand3_1 _3513_ (.B(_2115_),
    .C(_2200_),
    .A(net561),
    .Y(_0260_));
 sg13g2_or4_1 _3514_ (.A(_2205_),
    .B(_2485_),
    .C(_0259_),
    .D(_0260_),
    .X(_0261_));
 sg13g2_nor4_2 _3515_ (.A(_1999_),
    .B(_2135_),
    .C(_2249_),
    .Y(_0262_),
    .D(_2496_));
 sg13g2_a21oi_1 _3516_ (.A1(_0203_),
    .A2(_0262_),
    .Y(_0263_),
    .B1(_2149_));
 sg13g2_nor2_2 _3517_ (.A(_2041_),
    .B(_2112_),
    .Y(_0264_));
 sg13g2_nor2b_1 _3518_ (.A(_2162_),
    .B_N(_2285_),
    .Y(_0265_));
 sg13g2_nand4_1 _3519_ (.B(_0227_),
    .C(_0264_),
    .A(_2168_),
    .Y(_0266_),
    .D(_0265_));
 sg13g2_nor3_2 _3520_ (.A(_2029_),
    .B(net548),
    .C(_2374_),
    .Y(_0267_));
 sg13g2_nor4_2 _3521_ (.A(net566),
    .B(_2042_),
    .C(_2163_),
    .Y(_0268_),
    .D(_2173_));
 sg13g2_and2_1 _3522_ (.A(_0267_),
    .B(_0268_),
    .X(_0269_));
 sg13g2_nor2_1 _3523_ (.A(_2105_),
    .B(_0269_),
    .Y(_0270_));
 sg13g2_nor2_2 _3524_ (.A(_2053_),
    .B(_0176_),
    .Y(_0271_));
 sg13g2_nor4_2 _3525_ (.A(_2010_),
    .B(_2226_),
    .C(_2493_),
    .Y(_0272_),
    .D(_0204_));
 sg13g2_a21oi_1 _3526_ (.A1(_0271_),
    .A2(_0272_),
    .Y(_0273_),
    .B1(_2153_));
 sg13g2_nand3_1 _3527_ (.B(net556),
    .C(_2168_),
    .A(net564),
    .Y(_0274_));
 sg13g2_nor3_1 _3528_ (.A(_2233_),
    .B(_2332_),
    .C(_0274_),
    .Y(_0275_));
 sg13g2_and4_1 _3529_ (.A(net569),
    .B(_0184_),
    .C(_0188_),
    .D(_0275_),
    .X(_0276_));
 sg13g2_nor2_1 _3530_ (.A(_2130_),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_nand3_1 _3531_ (.B(_2218_),
    .C(_2309_),
    .A(_2137_),
    .Y(_0278_));
 sg13g2_nor4_2 _3532_ (.A(_2028_),
    .B(_2048_),
    .C(_0274_),
    .Y(_0279_),
    .D(_0278_));
 sg13g2_o21ai_1 _3533_ (.B1(net649),
    .Y(_0280_),
    .A1(_2126_),
    .A2(_0279_));
 sg13g2_a221oi_1 _3534_ (.B2(net653),
    .C1(_0273_),
    .B1(_0266_),
    .A1(net663),
    .Y(_0281_),
    .A2(_0261_));
 sg13g2_nor4_1 _3535_ (.A(_0263_),
    .B(_0270_),
    .C(_0277_),
    .D(_0280_),
    .Y(_0282_));
 sg13g2_a21oi_1 _3536_ (.A1(net596),
    .A2(net585),
    .Y(_0283_),
    .B1(net566));
 sg13g2_nand4_1 _3537_ (.B(_2032_),
    .C(net557),
    .A(_2019_),
    .Y(_0284_),
    .D(_0283_));
 sg13g2_nor3_2 _3538_ (.A(_2209_),
    .B(_2310_),
    .C(_0284_),
    .Y(_0285_));
 sg13g2_a22oi_1 _3539_ (.Y(_0286_),
    .B1(_0285_),
    .B2(net650),
    .A2(_0282_),
    .A1(_0281_));
 sg13g2_or2_1 _3540_ (.X(_0287_),
    .B(_0286_),
    .A(_0198_));
 sg13g2_nor4_2 _3541_ (.A(_2087_),
    .B(_2138_),
    .C(net544),
    .Y(_0288_),
    .D(_0226_));
 sg13g2_nand4_1 _3542_ (.B(_2081_),
    .C(_2176_),
    .A(_2019_),
    .Y(_0289_),
    .D(_2296_));
 sg13g2_nor4_2 _3543_ (.A(_2048_),
    .B(_2215_),
    .C(_2365_),
    .Y(_0290_),
    .D(_0289_));
 sg13g2_nor3_2 _3544_ (.A(_2135_),
    .B(_2167_),
    .C(_0180_),
    .Y(_0291_));
 sg13g2_nand4_1 _3545_ (.B(_2300_),
    .C(_0290_),
    .A(_2084_),
    .Y(_0292_),
    .D(_0291_));
 sg13g2_nor4_1 _3546_ (.A(net575),
    .B(_2135_),
    .C(_2257_),
    .D(net540),
    .Y(_0293_));
 sg13g2_nor4_2 _3547_ (.A(net563),
    .B(_2112_),
    .C(_2143_),
    .Y(_0294_),
    .D(_2264_));
 sg13g2_nand4_1 _3548_ (.B(_0171_),
    .C(_0293_),
    .A(_2088_),
    .Y(_0295_),
    .D(_0294_));
 sg13g2_nand3_1 _3549_ (.B(net560),
    .C(_2091_),
    .A(net564),
    .Y(_0296_));
 sg13g2_nor3_1 _3550_ (.A(_2080_),
    .B(net553),
    .C(_2485_),
    .Y(_0297_));
 sg13g2_nor4_1 _3551_ (.A(_2302_),
    .B(_2310_),
    .C(_2498_),
    .D(_0296_),
    .Y(_0298_));
 sg13g2_nand3_1 _3552_ (.B(_0297_),
    .C(_0298_),
    .A(_0163_),
    .Y(_0299_));
 sg13g2_and4_1 _3553_ (.A(_2054_),
    .B(_2113_),
    .C(_2117_),
    .D(_2320_),
    .X(_0300_));
 sg13g2_nand4_1 _3554_ (.B(_0169_),
    .C(_0175_),
    .A(_2267_),
    .Y(_0301_),
    .D(_0300_));
 sg13g2_nor4_2 _3555_ (.A(net570),
    .B(_2187_),
    .C(_0204_),
    .Y(_0302_),
    .D(_0301_));
 sg13g2_nor3_1 _3556_ (.A(_2029_),
    .B(_2052_),
    .C(net545),
    .Y(_0303_));
 sg13g2_nand3_1 _3557_ (.B(_0205_),
    .C(_0303_),
    .A(_2394_),
    .Y(_0304_));
 sg13g2_a21oi_1 _3558_ (.A1(net606),
    .A2(net596),
    .Y(_0305_),
    .B1(_2114_));
 sg13g2_nand4_1 _3559_ (.B(net541),
    .C(_0267_),
    .A(net564),
    .Y(_0306_),
    .D(_0305_));
 sg13g2_nand2_1 _3560_ (.Y(_0307_),
    .A(_2106_),
    .B(_0306_));
 sg13g2_nor4_1 _3561_ (.A(_2077_),
    .B(net553),
    .C(_2170_),
    .D(_2485_),
    .Y(_0308_));
 sg13g2_nand4_1 _3562_ (.B(_2086_),
    .C(_2375_),
    .A(_2084_),
    .Y(_0309_),
    .D(_0308_));
 sg13g2_o21ai_1 _3563_ (.B1(_0307_),
    .Y(_0310_),
    .A1(_2149_),
    .A2(_0302_));
 sg13g2_a221oi_1 _3564_ (.B2(_2154_),
    .C1(_0310_),
    .B1(_0304_),
    .A1(net653),
    .Y(_0311_),
    .A2(_0292_));
 sg13g2_a21o_1 _3565_ (.A2(_0299_),
    .A1(net659),
    .B1(net650),
    .X(_0312_));
 sg13g2_a221oi_1 _3566_ (.B2(net663),
    .C1(_0312_),
    .B1(_0309_),
    .A1(net648),
    .Y(_0313_),
    .A2(_0295_));
 sg13g2_a22oi_1 _3567_ (.Y(_0314_),
    .B1(_0311_),
    .B2(_0313_),
    .A2(_0288_),
    .A1(net650));
 sg13g2_or2_1 _3568_ (.X(_0315_),
    .B(_0314_),
    .A(_0287_));
 sg13g2_nor2_2 _3569_ (.A(_2018_),
    .B(_2266_),
    .Y(_0316_));
 sg13g2_a21oi_1 _3570_ (.A1(_2088_),
    .A2(_0316_),
    .Y(_0317_),
    .B1(_2098_));
 sg13g2_nand2_1 _3571_ (.Y(_0318_),
    .A(_2133_),
    .B(_2299_));
 sg13g2_nor2_1 _3572_ (.A(_2000_),
    .B(net588),
    .Y(_0319_));
 sg13g2_nor4_2 _3573_ (.A(_2015_),
    .B(_2259_),
    .C(_2264_),
    .Y(_0320_),
    .D(_0319_));
 sg13g2_and3_1 _3574_ (.X(_0321_),
    .A(_2088_),
    .B(_2258_),
    .C(_0156_));
 sg13g2_nor2_1 _3575_ (.A(_2105_),
    .B(_0321_),
    .Y(_0322_));
 sg13g2_a22oi_1 _3576_ (.Y(_0323_),
    .B1(_0318_),
    .B2(net647),
    .A2(_2257_),
    .A1(_2154_));
 sg13g2_o21ai_1 _3577_ (.B1(_0323_),
    .Y(_0324_),
    .A1(_2130_),
    .A2(_0320_));
 sg13g2_nor4_1 _3578_ (.A(net650),
    .B(_0317_),
    .C(_0322_),
    .D(_0324_),
    .Y(_0325_));
 sg13g2_nand2_1 _3579_ (.Y(_0326_),
    .A(_2171_),
    .B(_0320_));
 sg13g2_and4_1 _3580_ (.A(_2040_),
    .B(_2480_),
    .C(_0199_),
    .D(_0290_),
    .X(_0327_));
 sg13g2_inv_1 _3581_ (.Y(_0328_),
    .A(_0327_));
 sg13g2_a22oi_1 _3582_ (.Y(_0329_),
    .B1(_0328_),
    .B2(net653),
    .A2(_0326_),
    .A1(net659));
 sg13g2_nand4_1 _3583_ (.B(_2189_),
    .C(_2309_),
    .A(_2110_),
    .Y(_0330_),
    .D(_0316_));
 sg13g2_nor3_2 _3584_ (.A(_0220_),
    .B(_0226_),
    .C(_0330_),
    .Y(_0331_));
 sg13g2_a22oi_1 _3585_ (.Y(_0332_),
    .B1(_0331_),
    .B2(net650),
    .A2(_0329_),
    .A1(_0325_));
 sg13g2_nand2_1 _3586_ (.Y(_0333_),
    .A(_0315_),
    .B(_0332_));
 sg13g2_a21oi_1 _3587_ (.A1(_0315_),
    .A2(_0332_),
    .Y(_0334_),
    .B1(net632));
 sg13g2_or3_2 _3588_ (.A(net591),
    .B(_2264_),
    .C(_0319_),
    .X(_0335_));
 sg13g2_nand2b_1 _3589_ (.Y(_0336_),
    .B(_2131_),
    .A_N(_0335_));
 sg13g2_nand4_1 _3590_ (.B(_0156_),
    .C(_0160_),
    .A(_2391_),
    .Y(_0337_),
    .D(_0267_));
 sg13g2_nand4_1 _3591_ (.B(_2258_),
    .C(_2285_),
    .A(_2197_),
    .Y(_0338_),
    .D(_0175_));
 sg13g2_nor2_1 _3592_ (.A(_0337_),
    .B(_0338_),
    .Y(_0339_));
 sg13g2_nor2_1 _3593_ (.A(_2098_),
    .B(_0339_),
    .Y(_0340_));
 sg13g2_and2_2 _3594_ (.A(_2262_),
    .B(_2280_),
    .X(_0341_));
 sg13g2_nand4_1 _3595_ (.B(_0228_),
    .C(_0291_),
    .A(_2172_),
    .Y(_0342_),
    .D(_0341_));
 sg13g2_nand3_1 _3596_ (.B(_2133_),
    .C(net647),
    .A(net572),
    .Y(_0343_));
 sg13g2_a22oi_1 _3597_ (.Y(_0344_),
    .B1(_0170_),
    .B2(_2106_),
    .A2(_2294_),
    .A1(_2154_));
 sg13g2_a221oi_1 _3598_ (.B2(net653),
    .C1(net651),
    .B1(_0342_),
    .A1(_2031_),
    .Y(_0345_),
    .A2(net659));
 sg13g2_nand4_1 _3599_ (.B(_0343_),
    .C(_0344_),
    .A(_0336_),
    .Y(_0346_),
    .D(_0345_));
 sg13g2_nand2_1 _3600_ (.Y(_0347_),
    .A(net651),
    .B(_2182_));
 sg13g2_o21ai_1 _3601_ (.B1(_0347_),
    .Y(_0348_),
    .A1(_0340_),
    .A2(_0346_));
 sg13g2_or2_1 _3602_ (.X(_0349_),
    .B(_0348_),
    .A(_0334_));
 sg13g2_or2_1 _3603_ (.X(_0350_),
    .B(_2182_),
    .A(net660));
 sg13g2_nor2_1 _3604_ (.A(_2062_),
    .B(_0335_),
    .Y(_0351_));
 sg13g2_nor2_1 _3605_ (.A(_2243_),
    .B(_0339_),
    .Y(_0352_));
 sg13g2_nand3_1 _3606_ (.B(_2133_),
    .C(_2255_),
    .A(net572),
    .Y(_0353_));
 sg13g2_a22oi_1 _3607_ (.Y(_0354_),
    .B1(_0342_),
    .B2(_2150_),
    .A2(_2294_),
    .A1(_2099_));
 sg13g2_nor2_1 _3608_ (.A(_0351_),
    .B(_0352_),
    .Y(_0355_));
 sg13g2_nand4_1 _3609_ (.B(_0353_),
    .C(_0354_),
    .A(_0350_),
    .Y(_0356_),
    .D(_0355_));
 sg13g2_a221oi_1 _3610_ (.B2(_0170_),
    .C1(_0356_),
    .B1(net657),
    .A1(_2031_),
    .Y(_0357_),
    .A2(net652));
 sg13g2_inv_1 _3611_ (.Y(_0358_),
    .A(_0357_));
 sg13g2_nor2_1 _3612_ (.A(net660),
    .B(_0285_),
    .Y(_0359_));
 sg13g2_nand2b_1 _3613_ (.Y(_0360_),
    .B(net657),
    .A_N(_0269_));
 sg13g2_a21o_1 _3614_ (.A2(_0262_),
    .A1(_0203_),
    .B1(_2254_),
    .X(_0361_));
 sg13g2_a21oi_1 _3615_ (.A1(_0271_),
    .A2(_0272_),
    .Y(_0362_),
    .B1(net661));
 sg13g2_nand2b_1 _3616_ (.Y(_0363_),
    .B(_2061_),
    .A_N(_0276_));
 sg13g2_nor2_1 _3617_ (.A(_2070_),
    .B(_0279_),
    .Y(_0364_));
 sg13g2_a22oi_1 _3618_ (.Y(_0365_),
    .B1(_0266_),
    .B2(net655),
    .A2(_0261_),
    .A1(_2244_));
 sg13g2_nand4_1 _3619_ (.B(_0361_),
    .C(_0363_),
    .A(_0360_),
    .Y(_0366_),
    .D(_0365_));
 sg13g2_nor4_2 _3620_ (.A(_0359_),
    .B(_0362_),
    .C(_0364_),
    .Y(_0367_),
    .D(_0366_));
 sg13g2_nand2_1 _3621_ (.Y(_0368_),
    .A(_0243_),
    .B(_0367_));
 sg13g2_nand2_1 _3622_ (.Y(_0369_),
    .A(_2061_),
    .B(_0295_));
 sg13g2_and2_1 _3623_ (.A(net652),
    .B(_0299_),
    .X(_0370_));
 sg13g2_nor2_1 _3624_ (.A(_2254_),
    .B(_0302_),
    .Y(_0371_));
 sg13g2_a22oi_1 _3625_ (.Y(_0372_),
    .B1(_0309_),
    .B2(_2244_),
    .A2(_0306_),
    .A1(net657));
 sg13g2_nor2_1 _3626_ (.A(net660),
    .B(_0288_),
    .Y(_0373_));
 sg13g2_a22oi_1 _3627_ (.Y(_0374_),
    .B1(_0304_),
    .B2(_2099_),
    .A2(_0292_),
    .A1(net655));
 sg13g2_nand3_1 _3628_ (.B(_0372_),
    .C(_0374_),
    .A(_0369_),
    .Y(_0375_));
 sg13g2_nor4_2 _3629_ (.A(_0370_),
    .B(_0371_),
    .C(_0373_),
    .Y(_0376_),
    .D(_0375_));
 sg13g2_nor2b_1 _3630_ (.A(_0368_),
    .B_N(_0376_),
    .Y(_0377_));
 sg13g2_nand2b_1 _3631_ (.Y(_0378_),
    .B(net657),
    .A_N(_0321_));
 sg13g2_o21ai_1 _3632_ (.B1(_0378_),
    .Y(_0379_),
    .A1(_2062_),
    .A2(_0320_));
 sg13g2_a21oi_1 _3633_ (.A1(_2133_),
    .A2(_2299_),
    .Y(_0380_),
    .B1(_2254_));
 sg13g2_a21oi_1 _3634_ (.A1(_2088_),
    .A2(_0316_),
    .Y(_0381_),
    .B1(_2243_));
 sg13g2_a21o_1 _3635_ (.A2(_2257_),
    .A1(_2099_),
    .B1(_0380_),
    .X(_0382_));
 sg13g2_a22oi_1 _3636_ (.Y(_0383_),
    .B1(_0328_),
    .B2(net656),
    .A2(_0326_),
    .A1(net652));
 sg13g2_o21ai_1 _3637_ (.B1(_0383_),
    .Y(_0384_),
    .A1(net660),
    .A2(_0331_));
 sg13g2_nor4_2 _3638_ (.A(_0379_),
    .B(_0381_),
    .C(_0382_),
    .Y(_0385_),
    .D(_0384_));
 sg13g2_nor2_1 _3639_ (.A(_0377_),
    .B(_0385_),
    .Y(_0386_));
 sg13g2_nor2_1 _3640_ (.A(net632),
    .B(_0386_),
    .Y(_0387_));
 sg13g2_nor2_1 _3641_ (.A(_0357_),
    .B(_0387_),
    .Y(_0388_));
 sg13g2_nand2_1 _3642_ (.Y(_0389_),
    .A(net533),
    .B(_0388_));
 sg13g2_o21ai_1 _3643_ (.B1(_0389_),
    .Y(_0390_),
    .A1(net533),
    .A2(_0349_));
 sg13g2_or2_1 _3644_ (.X(_0391_),
    .B(_0390_),
    .A(_0061_));
 sg13g2_and2_1 _3645_ (.A(_0061_),
    .B(_0390_),
    .X(_0392_));
 sg13g2_a21o_1 _3646_ (.A2(_0348_),
    .A1(net638),
    .B1(_0334_),
    .X(_0393_));
 sg13g2_a21oi_1 _3647_ (.A1(net633),
    .A2(_0332_),
    .Y(_0394_),
    .B1(_0393_));
 sg13g2_nor2_1 _3648_ (.A(net637),
    .B(_0385_),
    .Y(_0395_));
 sg13g2_a21oi_1 _3649_ (.A1(_0358_),
    .A2(_0386_),
    .Y(_0396_),
    .B1(net632));
 sg13g2_nor2_1 _3650_ (.A(_0395_),
    .B(_0396_),
    .Y(_0397_));
 sg13g2_mux2_2 _3651_ (.A0(_0394_),
    .A1(_0397_),
    .S(net533),
    .X(_0398_));
 sg13g2_or2_1 _3652_ (.X(_0399_),
    .B(_0398_),
    .A(\wirecube_top_inst.edge_function_inst.pixel_x_i[5] ));
 sg13g2_o21ai_1 _3653_ (.B1(_0334_),
    .Y(_0400_),
    .A1(_0315_),
    .A2(_0332_));
 sg13g2_nand2_1 _3654_ (.Y(_0401_),
    .A(net632),
    .B(_0286_));
 sg13g2_nand2_1 _3655_ (.Y(_0402_),
    .A(_0400_),
    .B(_0401_));
 sg13g2_nand2_1 _3656_ (.Y(_0403_),
    .A(_0377_),
    .B(_0385_));
 sg13g2_nand2_1 _3657_ (.Y(_0404_),
    .A(_0387_),
    .B(_0403_));
 sg13g2_o21ai_1 _3658_ (.B1(_0404_),
    .Y(_0405_),
    .A1(net638),
    .A2(_0367_));
 sg13g2_mux2_2 _3659_ (.A0(_0402_),
    .A1(_0405_),
    .S(net534),
    .X(_0406_));
 sg13g2_nand2b_1 _3660_ (.Y(_0407_),
    .B(\wirecube_top_inst.edge_function_inst.pixel_x_i[3] ),
    .A_N(_0406_));
 sg13g2_inv_1 _3661_ (.Y(_0408_),
    .A(_0407_));
 sg13g2_nand2_1 _3662_ (.Y(_0409_),
    .A(_1848_),
    .B(_0406_));
 sg13g2_inv_1 _3663_ (.Y(_0410_),
    .A(_0409_));
 sg13g2_nand2_1 _3664_ (.Y(_0411_),
    .A(_0287_),
    .B(_0314_));
 sg13g2_a21oi_1 _3665_ (.A1(_0315_),
    .A2(_0411_),
    .Y(_0412_),
    .B1(net632));
 sg13g2_a21oi_1 _3666_ (.A1(net633),
    .A2(_0198_),
    .Y(_0413_),
    .B1(_0412_));
 sg13g2_and3_1 _3667_ (.X(_0414_),
    .A(net538),
    .B(net539),
    .C(_0413_));
 sg13g2_nor2_1 _3668_ (.A(net637),
    .B(_0243_),
    .Y(_0415_));
 sg13g2_xor2_1 _3669_ (.B(_0376_),
    .A(_0368_),
    .X(_0416_));
 sg13g2_a21oi_2 _3670_ (.B1(_0415_),
    .Y(_0417_),
    .A2(_0416_),
    .A1(net638));
 sg13g2_a21oi_2 _3671_ (.B1(_0414_),
    .Y(_0418_),
    .A2(_0417_),
    .A1(net534));
 sg13g2_a21o_1 _3672_ (.A2(_0417_),
    .A1(net533),
    .B1(_0414_),
    .X(_0419_));
 sg13g2_nand4_1 _3673_ (.B(_2086_),
    .C(_2115_),
    .A(_2084_),
    .Y(_0420_),
    .D(net541));
 sg13g2_nor4_2 _3674_ (.A(_2198_),
    .B(_2231_),
    .C(_2374_),
    .Y(_0421_),
    .D(_0420_));
 sg13g2_a21oi_1 _3675_ (.A1(_2106_),
    .A2(net542),
    .Y(_0422_),
    .B1(net663));
 sg13g2_a21oi_1 _3676_ (.A1(net607),
    .A2(net585),
    .Y(_0423_),
    .B1(_2052_));
 sg13g2_nand4_1 _3677_ (.B(net560),
    .C(_2189_),
    .A(net569),
    .Y(_0424_),
    .D(_0423_));
 sg13g2_nor4_2 _3678_ (.A(_2225_),
    .B(_2374_),
    .C(_0289_),
    .Y(_0425_),
    .D(_0424_));
 sg13g2_inv_1 _3679_ (.Y(_0426_),
    .A(_0425_));
 sg13g2_nor3_2 _3680_ (.A(net575),
    .B(_2031_),
    .C(_2210_),
    .Y(_0427_));
 sg13g2_nor4_1 _3681_ (.A(_2112_),
    .B(_2201_),
    .C(_2263_),
    .D(_2498_),
    .Y(_0428_));
 sg13g2_nand3_1 _3682_ (.B(_0427_),
    .C(_0428_),
    .A(_0297_),
    .Y(_0429_));
 sg13g2_a22oi_1 _3683_ (.Y(_0430_),
    .B1(_0429_),
    .B2(net648),
    .A2(_0426_),
    .A1(net650));
 sg13g2_o21ai_1 _3684_ (.B1(_0430_),
    .Y(_0431_),
    .A1(_0421_),
    .A2(_0422_));
 sg13g2_nor2_1 _3685_ (.A(net544),
    .B(_0429_),
    .Y(_0432_));
 sg13g2_nand2_1 _3686_ (.Y(_0433_),
    .A(net541),
    .B(_0425_));
 sg13g2_nand2_1 _3687_ (.Y(_0434_),
    .A(_2079_),
    .B(net550));
 sg13g2_nor3_1 _3688_ (.A(_2256_),
    .B(_0170_),
    .C(_0434_),
    .Y(_0435_));
 sg13g2_nand3_1 _3689_ (.B(_0205_),
    .C(_0435_),
    .A(_0169_),
    .Y(_0436_));
 sg13g2_o21ai_1 _3690_ (.B1(_2153_),
    .Y(_0437_),
    .A1(_2149_),
    .A2(net544));
 sg13g2_a221oi_1 _3691_ (.B2(_0437_),
    .C1(net637),
    .B1(_0436_),
    .A1(net653),
    .Y(_0438_),
    .A2(_0433_));
 sg13g2_o21ai_1 _3692_ (.B1(_0438_),
    .Y(_0439_),
    .A1(_2126_),
    .A2(_0432_));
 sg13g2_nand2_1 _3693_ (.Y(_0440_),
    .A(_0198_),
    .B(_0286_));
 sg13g2_nand3_1 _3694_ (.B(_0287_),
    .C(_0440_),
    .A(net637),
    .Y(_0441_));
 sg13g2_o21ai_1 _3695_ (.B1(_0441_),
    .Y(_0442_),
    .A1(_0431_),
    .A2(_0439_));
 sg13g2_inv_1 _3696_ (.Y(_0443_),
    .A(_0442_));
 sg13g2_a21oi_1 _3697_ (.A1(net657),
    .A2(net541),
    .Y(_0444_),
    .B1(_2244_));
 sg13g2_nor2_1 _3698_ (.A(_0421_),
    .B(_0444_),
    .Y(_0445_));
 sg13g2_o21ai_1 _3699_ (.B1(net661),
    .Y(_0446_),
    .A1(net544),
    .A2(_2254_));
 sg13g2_o21ai_1 _3700_ (.B1(net652),
    .Y(_0447_),
    .A1(net544),
    .A2(_0429_));
 sg13g2_a221oi_1 _3701_ (.B2(_2061_),
    .C1(_0445_),
    .B1(_0429_),
    .A1(_2102_),
    .Y(_0448_),
    .A2(_0426_));
 sg13g2_a22oi_1 _3702_ (.Y(_0449_),
    .B1(_0436_),
    .B2(_0446_),
    .A2(_0433_),
    .A1(net656));
 sg13g2_nand4_1 _3703_ (.B(_0447_),
    .C(_0448_),
    .A(net633),
    .Y(_0450_),
    .D(_0449_));
 sg13g2_xnor2_1 _3704_ (.Y(_0451_),
    .A(_0243_),
    .B(_0367_));
 sg13g2_o21ai_1 _3705_ (.B1(_0450_),
    .Y(_0452_),
    .A1(net632),
    .A2(_0451_));
 sg13g2_inv_1 _3706_ (.Y(_0453_),
    .A(_0452_));
 sg13g2_o21ai_1 _3707_ (.B1(_0453_),
    .Y(_0454_),
    .A1(_2537_),
    .A2(_2541_));
 sg13g2_nand3_1 _3708_ (.B(net539),
    .C(_0443_),
    .A(net538),
    .Y(_0455_));
 sg13g2_nand2_2 _3709_ (.Y(_0456_),
    .A(_0454_),
    .B(_0455_));
 sg13g2_and2_1 _3710_ (.A(_0454_),
    .B(_0455_),
    .X(_0457_));
 sg13g2_nor2_1 _3711_ (.A(_1850_),
    .B(_0456_),
    .Y(_0458_));
 sg13g2_xnor2_1 _3712_ (.Y(_0459_),
    .A(_0057_),
    .B(_0457_));
 sg13g2_xnor2_1 _3713_ (.Y(_0460_),
    .A(net196),
    .B(_0456_));
 sg13g2_a21o_1 _3714_ (.A2(_0459_),
    .A1(_0252_),
    .B1(_0458_),
    .X(_0461_));
 sg13g2_xnor2_1 _3715_ (.Y(_0462_),
    .A(_0056_),
    .B(_0419_));
 sg13g2_a22oi_1 _3716_ (.Y(_0463_),
    .B1(_0461_),
    .B2(_0462_),
    .A2(_0419_),
    .A1(net681));
 sg13g2_a221oi_1 _3717_ (.B2(_0462_),
    .C1(_0408_),
    .B1(_0461_),
    .A1(net681),
    .Y(_0464_),
    .A2(_0419_));
 sg13g2_nor2_1 _3718_ (.A(_0410_),
    .B(_0464_),
    .Y(_0465_));
 sg13g2_nand2_1 _3719_ (.Y(_0466_),
    .A(_0333_),
    .B(_0348_));
 sg13g2_and2_1 _3720_ (.A(net632),
    .B(_0314_),
    .X(_0467_));
 sg13g2_a21o_1 _3721_ (.A2(_0466_),
    .A1(_0393_),
    .B1(_0467_),
    .X(_0468_));
 sg13g2_o21ai_1 _3722_ (.B1(_0396_),
    .Y(_0469_),
    .A1(_0358_),
    .A2(_0386_));
 sg13g2_o21ai_1 _3723_ (.B1(_0469_),
    .Y(_0470_),
    .A1(net637),
    .A2(_0376_));
 sg13g2_mux2_2 _3724_ (.A0(_0468_),
    .A1(_0470_),
    .S(net533),
    .X(_0471_));
 sg13g2_xnor2_1 _3725_ (.Y(_0472_),
    .A(net203),
    .B(_0471_));
 sg13g2_xor2_1 _3726_ (.B(_0471_),
    .A(_0055_),
    .X(_0473_));
 sg13g2_nor2_1 _3727_ (.A(_1847_),
    .B(_0471_),
    .Y(_0474_));
 sg13g2_and2_1 _3728_ (.A(\wirecube_top_inst.edge_function_inst.pixel_x_i[5] ),
    .B(_0398_),
    .X(_0475_));
 sg13g2_inv_1 _3729_ (.Y(_0476_),
    .A(_0475_));
 sg13g2_nand2_1 _3730_ (.Y(_0477_),
    .A(_0399_),
    .B(_0474_));
 sg13g2_nand2_1 _3731_ (.Y(_0478_),
    .A(_0399_),
    .B(_0476_));
 sg13g2_nor2_1 _3732_ (.A(_0472_),
    .B(_0478_),
    .Y(_0479_));
 sg13g2_or4_1 _3733_ (.A(_0410_),
    .B(_0464_),
    .C(_0472_),
    .D(_0478_),
    .X(_0480_));
 sg13g2_nand3_1 _3734_ (.B(_0477_),
    .C(_0480_),
    .A(_0476_),
    .Y(_0481_));
 sg13g2_nand4_1 _3735_ (.B(_0476_),
    .C(_0477_),
    .A(_0391_),
    .Y(_0482_),
    .D(_0480_));
 sg13g2_nor2b_1 _3736_ (.A(_0392_),
    .B_N(_0482_),
    .Y(_0483_));
 sg13g2_nand2_1 _3737_ (.Y(_0484_),
    .A(_0407_),
    .B(_0409_));
 sg13g2_xnor2_1 _3738_ (.Y(_0485_),
    .A(net189),
    .B(_0390_));
 sg13g2_nor2_1 _3739_ (.A(_0484_),
    .B(_0485_),
    .Y(_0486_));
 sg13g2_nor2_1 _3740_ (.A(_0028_),
    .B(_0460_),
    .Y(_0487_));
 sg13g2_nand4_1 _3741_ (.B(_0479_),
    .C(_0486_),
    .A(_0462_),
    .Y(_0488_),
    .D(_0487_));
 sg13g2_nand3b_1 _3742_ (.B(_0482_),
    .C(_0488_),
    .Y(_0489_),
    .A_N(_0392_));
 sg13g2_nor2_1 _3743_ (.A(net533),
    .B(_0388_),
    .Y(_0490_));
 sg13g2_a21oi_1 _3744_ (.A1(net534),
    .A2(_0349_),
    .Y(_0491_),
    .B1(_0490_));
 sg13g2_a21o_2 _3745_ (.A2(_0349_),
    .A1(net534),
    .B1(_0490_),
    .X(_0492_));
 sg13g2_mux2_1 _3746_ (.A0(_0397_),
    .A1(_0394_),
    .S(net533),
    .X(_0493_));
 sg13g2_and2_1 _3747_ (.A(\wirecube_top_inst.edge_function_inst.pixel_x_i[5] ),
    .B(_0493_),
    .X(_0494_));
 sg13g2_inv_1 _3748_ (.Y(_0495_),
    .A(_0494_));
 sg13g2_nor2_1 _3749_ (.A(\wirecube_top_inst.edge_function_inst.pixel_x_i[5] ),
    .B(_0493_),
    .Y(_0496_));
 sg13g2_or2_1 _3750_ (.X(_0497_),
    .B(_0496_),
    .A(_0494_));
 sg13g2_mux2_1 _3751_ (.A0(_0470_),
    .A1(_0468_),
    .S(net533),
    .X(_0498_));
 sg13g2_inv_1 _3752_ (.Y(_0499_),
    .A(_0498_));
 sg13g2_xnor2_1 _3753_ (.Y(_0500_),
    .A(_0055_),
    .B(_0498_));
 sg13g2_inv_1 _3754_ (.Y(_0501_),
    .A(_0500_));
 sg13g2_nor2_1 _3755_ (.A(_0497_),
    .B(_0500_),
    .Y(_0502_));
 sg13g2_a22oi_1 _3756_ (.Y(_0503_),
    .B1(_0400_),
    .B2(_0401_),
    .A2(net539),
    .A1(net538));
 sg13g2_o21ai_1 _3757_ (.B1(_0402_),
    .Y(_0504_),
    .A1(_2537_),
    .A2(_2541_));
 sg13g2_and3_1 _3758_ (.X(_0505_),
    .A(net538),
    .B(net539),
    .C(_0405_));
 sg13g2_nand3_1 _3759_ (.B(net539),
    .C(_0405_),
    .A(net538),
    .Y(_0506_));
 sg13g2_nor2_1 _3760_ (.A(_0503_),
    .B(_0505_),
    .Y(_0507_));
 sg13g2_nor3_2 _3761_ (.A(_1848_),
    .B(_0503_),
    .C(_0505_),
    .Y(_0508_));
 sg13g2_a21oi_1 _3762_ (.A1(_0504_),
    .A2(_0506_),
    .Y(_0509_),
    .B1(\wirecube_top_inst.edge_function_inst.pixel_x_i[3] ));
 sg13g2_o21ai_1 _3763_ (.B1(_1848_),
    .Y(_0510_),
    .A1(_0503_),
    .A2(_0505_));
 sg13g2_nand3_1 _3764_ (.B(net539),
    .C(_0417_),
    .A(net538),
    .Y(_0511_));
 sg13g2_o21ai_1 _3765_ (.B1(_0413_),
    .Y(_0512_),
    .A1(_2537_),
    .A2(_2541_));
 sg13g2_nand2_2 _3766_ (.Y(_0513_),
    .A(_0511_),
    .B(_0512_));
 sg13g2_o21ai_1 _3767_ (.B1(_0443_),
    .Y(_0514_),
    .A1(_2537_),
    .A2(_2541_));
 sg13g2_nand3_1 _3768_ (.B(net539),
    .C(_0453_),
    .A(net538),
    .Y(_0515_));
 sg13g2_nand2_1 _3769_ (.Y(_0516_),
    .A(_0514_),
    .B(_0515_));
 sg13g2_and2_1 _3770_ (.A(_0514_),
    .B(_0515_),
    .X(_0517_));
 sg13g2_nand3_1 _3771_ (.B(_0514_),
    .C(_0515_),
    .A(_0057_),
    .Y(_0518_));
 sg13g2_a21o_1 _3772_ (.A2(_0515_),
    .A1(_0514_),
    .B1(_0057_),
    .X(_0519_));
 sg13g2_and2_1 _3773_ (.A(_0518_),
    .B(_0519_),
    .X(_0520_));
 sg13g2_a22oi_1 _3774_ (.Y(_0521_),
    .B1(_0518_),
    .B2(_0519_),
    .A2(_0254_),
    .A1(_0058_));
 sg13g2_nand2b_1 _3775_ (.Y(_0522_),
    .B(_0255_),
    .A_N(_0520_));
 sg13g2_nor2_1 _3776_ (.A(_1850_),
    .B(_0516_),
    .Y(_0523_));
 sg13g2_or2_1 _3777_ (.X(_0524_),
    .B(_0523_),
    .A(_0521_));
 sg13g2_a21oi_2 _3778_ (.B1(_0056_),
    .Y(_0525_),
    .A2(_0512_),
    .A1(_0511_));
 sg13g2_and3_1 _3779_ (.X(_0526_),
    .A(_0056_),
    .B(_0511_),
    .C(_0512_));
 sg13g2_nor2_2 _3780_ (.A(_0525_),
    .B(_0526_),
    .Y(_0527_));
 sg13g2_a22oi_1 _3781_ (.Y(_0528_),
    .B1(_0524_),
    .B2(_0527_),
    .A2(_0513_),
    .A1(net681));
 sg13g2_nand3_1 _3782_ (.B(_0510_),
    .C(_0513_),
    .A(net681),
    .Y(_0529_));
 sg13g2_nor2_1 _3783_ (.A(_0508_),
    .B(_0509_),
    .Y(_0530_));
 sg13g2_nor4_2 _3784_ (.A(_0508_),
    .B(_0509_),
    .C(_0525_),
    .Y(_0531_),
    .D(_0526_));
 sg13g2_o21ai_1 _3785_ (.B1(_0531_),
    .Y(_0532_),
    .A1(_0521_),
    .A2(_0523_));
 sg13g2_nand3b_1 _3786_ (.B(_0529_),
    .C(_0532_),
    .Y(_0533_),
    .A_N(_0508_));
 sg13g2_nor2_1 _3787_ (.A(_1847_),
    .B(_0498_),
    .Y(_0534_));
 sg13g2_nor2b_1 _3788_ (.A(_0496_),
    .B_N(_0534_),
    .Y(_0535_));
 sg13g2_or2_1 _3789_ (.X(_0536_),
    .B(_0535_),
    .A(_0494_));
 sg13g2_a21oi_1 _3790_ (.A1(_0502_),
    .A2(_0533_),
    .Y(_0537_),
    .B1(_0536_));
 sg13g2_a221oi_1 _3791_ (.B2(_0533_),
    .C1(_0536_),
    .B1(_0502_),
    .A1(\wirecube_top_inst.edge_function_inst.pixel_x_i[6] ),
    .Y(_0538_),
    .A2(_0492_));
 sg13g2_a21oi_1 _3792_ (.A1(_1846_),
    .A2(_0491_),
    .Y(_0539_),
    .B1(_0538_));
 sg13g2_nor2_1 _3793_ (.A(_0456_),
    .B(_0517_),
    .Y(_0540_));
 sg13g2_nand2b_1 _3794_ (.Y(_0541_),
    .B(_0251_),
    .A_N(_0254_));
 sg13g2_a22oi_1 _3795_ (.Y(_0542_),
    .B1(_0517_),
    .B2(_0456_),
    .A2(_0513_),
    .A1(_0418_));
 sg13g2_o21ai_1 _3796_ (.B1(_0542_),
    .Y(_0543_),
    .A1(_0540_),
    .A2(_0541_));
 sg13g2_nor2_1 _3797_ (.A(_0418_),
    .B(_0513_),
    .Y(_0544_));
 sg13g2_nor2_1 _3798_ (.A(_0471_),
    .B(_0499_),
    .Y(_0545_));
 sg13g2_nor2_1 _3799_ (.A(_0406_),
    .B(_0507_),
    .Y(_0546_));
 sg13g2_nor2_1 _3800_ (.A(_0544_),
    .B(_0546_),
    .Y(_0547_));
 sg13g2_a22oi_1 _3801_ (.Y(_0548_),
    .B1(_0543_),
    .B2(_0547_),
    .A2(_0507_),
    .A1(_0406_));
 sg13g2_or2_1 _3802_ (.X(_0549_),
    .B(_0548_),
    .A(_0545_));
 sg13g2_nor2b_1 _3803_ (.A(_0398_),
    .B_N(_0493_),
    .Y(_0550_));
 sg13g2_a21oi_1 _3804_ (.A1(_0471_),
    .A2(_0499_),
    .Y(_0551_),
    .B1(_0550_));
 sg13g2_nand2b_1 _3805_ (.Y(_0552_),
    .B(_0398_),
    .A_N(_0493_));
 sg13g2_o21ai_1 _3806_ (.B1(_0552_),
    .Y(_0553_),
    .A1(_0390_),
    .A2(_0492_));
 sg13g2_a21oi_1 _3807_ (.A1(_0549_),
    .A2(_0551_),
    .Y(_0554_),
    .B1(_0553_));
 sg13g2_a21o_2 _3808_ (.A2(_0492_),
    .A1(_0390_),
    .B1(_0554_),
    .X(_0555_));
 sg13g2_a21oi_2 _3809_ (.B1(_0554_),
    .Y(_0556_),
    .A2(_0492_),
    .A1(_0390_));
 sg13g2_a21oi_2 _3810_ (.B1(_0556_),
    .Y(_0557_),
    .A2(_0539_),
    .A1(_0489_));
 sg13g2_xnor2_1 _3811_ (.Y(_0558_),
    .A(net133),
    .B(_0491_));
 sg13g2_nand4_1 _3812_ (.B(_0502_),
    .C(_0531_),
    .A(_0257_),
    .Y(_0559_),
    .D(_0558_));
 sg13g2_o21ai_1 _3813_ (.B1(_0539_),
    .Y(_0560_),
    .A1(_0522_),
    .A2(_0559_));
 sg13g2_a21oi_2 _3814_ (.B1(_0555_),
    .Y(_0561_),
    .A2(_0560_),
    .A1(_0483_));
 sg13g2_mux2_1 _3815_ (.A0(_2448_),
    .A1(_2446_),
    .S(net535),
    .X(_0562_));
 sg13g2_nor2_1 _3816_ (.A(_1842_),
    .B(_0562_),
    .Y(_0563_));
 sg13g2_nand2_1 _3817_ (.Y(_0564_),
    .A(_2444_),
    .B(net535));
 sg13g2_o21ai_1 _3818_ (.B1(_0564_),
    .Y(_0565_),
    .A1(_2405_),
    .A2(net535));
 sg13g2_nand2_1 _3819_ (.Y(_0566_),
    .A(net153),
    .B(_0565_));
 sg13g2_mux2_1 _3820_ (.A0(_2457_),
    .A1(_2463_),
    .S(net535),
    .X(_0567_));
 sg13g2_and2_1 _3821_ (.A(\wirecube_top_inst.edge_function_inst.pixel_y_i[3] ),
    .B(_0567_),
    .X(_0568_));
 sg13g2_mux2_1 _3822_ (.A0(_2473_),
    .A1(_2469_),
    .S(net536),
    .X(_0569_));
 sg13g2_nand2_1 _3823_ (.Y(_0570_),
    .A(net204),
    .B(_0569_));
 sg13g2_nand3_1 _3824_ (.B(_2538_),
    .C(_2542_),
    .A(_2517_),
    .Y(_0571_));
 sg13g2_o21ai_1 _3825_ (.B1(_2506_),
    .Y(_0572_),
    .A1(_2537_),
    .A2(_2541_));
 sg13g2_a21oi_1 _3826_ (.A1(_0571_),
    .A2(_0572_),
    .Y(_0573_),
    .B1(_1845_));
 sg13g2_nand3_1 _3827_ (.B(_0571_),
    .C(_0572_),
    .A(_1845_),
    .Y(_0574_));
 sg13g2_nand2b_1 _3828_ (.Y(_0575_),
    .B(_0574_),
    .A_N(_0573_));
 sg13g2_a21oi_2 _3829_ (.B1(_0573_),
    .Y(_0576_),
    .A2(_0574_),
    .A1(_0155_));
 sg13g2_xor2_1 _3830_ (.B(_0569_),
    .A(net193),
    .X(_0577_));
 sg13g2_o21ai_1 _3831_ (.B1(_0570_),
    .Y(_0578_),
    .A1(_0576_),
    .A2(_0577_));
 sg13g2_xnor2_1 _3832_ (.Y(_0579_),
    .A(_1843_),
    .B(_0567_));
 sg13g2_a21oi_1 _3833_ (.A1(_0578_),
    .A2(_0579_),
    .Y(_0580_),
    .B1(_0568_));
 sg13g2_xor2_1 _3834_ (.B(_0565_),
    .A(net195),
    .X(_0581_));
 sg13g2_o21ai_1 _3835_ (.B1(_0566_),
    .Y(_0582_),
    .A1(_0580_),
    .A2(_0581_));
 sg13g2_xor2_1 _3836_ (.B(_0562_),
    .A(net166),
    .X(_0583_));
 sg13g2_a21oi_1 _3837_ (.A1(_0582_),
    .A2(_0583_),
    .Y(_0584_),
    .B1(_0563_));
 sg13g2_xor2_1 _3838_ (.B(_2277_),
    .A(net191),
    .X(_0585_));
 sg13g2_nor2_1 _3839_ (.A(_0584_),
    .B(_0585_),
    .Y(_0586_));
 sg13g2_a21oi_1 _3840_ (.A1(net107),
    .A2(_2277_),
    .Y(_0587_),
    .B1(_0586_));
 sg13g2_xor2_1 _3841_ (.B(_2278_),
    .A(_0051_),
    .X(_0588_));
 sg13g2_inv_1 _3842_ (.Y(_0589_),
    .A(_0588_));
 sg13g2_mux2_1 _3843_ (.A0(_2463_),
    .A1(_2457_),
    .S(net535),
    .X(_0590_));
 sg13g2_nand2_1 _3844_ (.Y(_0591_),
    .A(\wirecube_top_inst.edge_function_inst.pixel_y_i[3] ),
    .B(_0590_));
 sg13g2_nor2_1 _3845_ (.A(_2469_),
    .B(net535),
    .Y(_0592_));
 sg13g2_a21oi_2 _3846_ (.B1(_0592_),
    .Y(_0593_),
    .A2(net535),
    .A1(_2472_));
 sg13g2_xnor2_1 _3847_ (.Y(_0594_),
    .A(_0053_),
    .B(_0593_));
 sg13g2_mux2_1 _3848_ (.A0(_2446_),
    .A1(_2448_),
    .S(net535),
    .X(_0595_));
 sg13g2_nor2_1 _3849_ (.A(_1842_),
    .B(_0595_),
    .Y(_0596_));
 sg13g2_inv_1 _3850_ (.Y(_0597_),
    .A(_0596_));
 sg13g2_and2_1 _3851_ (.A(_1842_),
    .B(_0595_),
    .X(_0598_));
 sg13g2_nor2_1 _3852_ (.A(_0596_),
    .B(_0598_),
    .Y(_0599_));
 sg13g2_and3_1 _3853_ (.X(_0600_),
    .A(_2545_),
    .B(_0589_),
    .C(_0594_));
 sg13g2_mux2_2 _3854_ (.A0(_2506_),
    .A1(_2517_),
    .S(net537),
    .X(_0601_));
 sg13g2_nor2_1 _3855_ (.A(\wirecube_top_inst.edge_function_inst.pixel_y_i[1] ),
    .B(_0601_),
    .Y(_0602_));
 sg13g2_xnor2_1 _3856_ (.Y(_0603_),
    .A(\wirecube_top_inst.edge_function_inst.pixel_y_i[1] ),
    .B(_0601_));
 sg13g2_nor2_1 _3857_ (.A(_2546_),
    .B(_0603_),
    .Y(_0604_));
 sg13g2_nor2_1 _3858_ (.A(\wirecube_top_inst.edge_function_inst.pixel_y_i[3] ),
    .B(_0590_),
    .Y(_0605_));
 sg13g2_inv_1 _3859_ (.Y(_0606_),
    .A(_0605_));
 sg13g2_nor2_1 _3860_ (.A(_2444_),
    .B(net536),
    .Y(_0607_));
 sg13g2_a21oi_2 _3861_ (.B1(_0607_),
    .Y(_0608_),
    .A2(net536),
    .A1(_2405_));
 sg13g2_xor2_1 _3862_ (.B(_0608_),
    .A(_0052_),
    .X(_0609_));
 sg13g2_nor2_1 _3863_ (.A(_0605_),
    .B(_0609_),
    .Y(_0610_));
 sg13g2_and4_1 _3864_ (.A(_0591_),
    .B(_0599_),
    .C(_0600_),
    .D(_0610_),
    .X(_0611_));
 sg13g2_nand2_1 _3865_ (.Y(_0612_),
    .A(_0591_),
    .B(_0606_));
 sg13g2_nand2_1 _3866_ (.Y(_0613_),
    .A(net107),
    .B(_2278_));
 sg13g2_a21oi_1 _3867_ (.A1(\wirecube_top_inst.edge_function_inst.pixel_y_i[1] ),
    .A2(_0601_),
    .Y(_0614_),
    .B1(_2545_));
 sg13g2_o21ai_1 _3868_ (.B1(_0594_),
    .Y(_0615_),
    .A1(\wirecube_top_inst.edge_function_inst.pixel_y_i[1] ),
    .A2(_0601_));
 sg13g2_a22oi_1 _3869_ (.Y(_0616_),
    .B1(_0593_),
    .B2(\wirecube_top_inst.edge_function_inst.pixel_y_i[2] ),
    .A2(_0590_),
    .A1(\wirecube_top_inst.edge_function_inst.pixel_y_i[3] ));
 sg13g2_o21ai_1 _3870_ (.B1(_0616_),
    .Y(_0617_),
    .A1(_0614_),
    .A2(_0615_));
 sg13g2_a221oi_1 _3871_ (.B2(_0617_),
    .C1(_0596_),
    .B1(_0610_),
    .A1(\wirecube_top_inst.edge_function_inst.pixel_y_i[4] ),
    .Y(_0618_),
    .A2(_0608_));
 sg13g2_or3_1 _3872_ (.A(_0588_),
    .B(_0598_),
    .C(_0618_),
    .X(_0619_));
 sg13g2_a22oi_1 _3873_ (.Y(_0620_),
    .B1(_0613_),
    .B2(_0619_),
    .A2(_0611_),
    .A1(_0604_));
 sg13g2_nor4_2 _3874_ (.A(_0557_),
    .B(_0561_),
    .C(_0587_),
    .Y(_0042_),
    .D(_0620_));
 sg13g2_a21oi_1 _3875_ (.A1(\wirecube_top_inst.counter_h[7] ),
    .A2(\wirecube_top_inst.counter_h[6] ),
    .Y(_0621_),
    .B1(net119));
 sg13g2_nand3_1 _3876_ (.B(net128),
    .C(net125),
    .A(net135),
    .Y(_0622_));
 sg13g2_nor2_1 _3877_ (.A(_0621_),
    .B(_0622_),
    .Y(_0623_));
 sg13g2_nand2_1 _3878_ (.Y(_0624_),
    .A(_1838_),
    .B(net701));
 sg13g2_nor2_1 _3879_ (.A(\wirecube_top_inst.counter_v[3] ),
    .B(\wirecube_top_inst.counter_v[2] ),
    .Y(_0625_));
 sg13g2_and2_1 _3880_ (.A(\wirecube_top_inst.counter_v[0] ),
    .B(net116),
    .X(_0626_));
 sg13g2_nor4_1 _3881_ (.A(net702),
    .B(\wirecube_top_inst.counter_v[2] ),
    .C(_0624_),
    .D(_0626_),
    .Y(_0627_));
 sg13g2_nand3_1 _3882_ (.B(net699),
    .C(\wirecube_top_inst.counter_v[8] ),
    .A(\wirecube_top_inst.counter_v[7] ),
    .Y(_0628_));
 sg13g2_inv_1 _3883_ (.Y(_0629_),
    .A(_0628_));
 sg13g2_nor2_1 _3884_ (.A(net700),
    .B(net701),
    .Y(_0630_));
 sg13g2_nand2_1 _3885_ (.Y(_0631_),
    .A(\wirecube_top_inst.counter_v[10] ),
    .B(\wirecube_top_inst.counter_v[9] ));
 sg13g2_nor4_1 _3886_ (.A(_0627_),
    .B(_0628_),
    .C(_0630_),
    .D(_0631_),
    .Y(_0632_));
 sg13g2_or2_2 _3887_ (.X(_0633_),
    .B(_0632_),
    .A(_0623_));
 sg13g2_o21ai_1 _3888_ (.B1(_1891_),
    .Y(_0634_),
    .A1(_1804_),
    .A2(_1875_));
 sg13g2_a21oi_1 _3889_ (.A1(_1804_),
    .A2(_1875_),
    .Y(_0635_),
    .B1(_0634_));
 sg13g2_nor3_2 _3890_ (.A(net686),
    .B(_1875_),
    .C(_1892_),
    .Y(_0636_));
 sg13g2_nor2_1 _3891_ (.A(net690),
    .B(_1899_),
    .Y(_0637_));
 sg13g2_nor3_1 _3892_ (.A(net690),
    .B(net685),
    .C(_1888_),
    .Y(_0638_));
 sg13g2_nor2_1 _3893_ (.A(_0637_),
    .B(_0638_),
    .Y(_0639_));
 sg13g2_nand2b_1 _3894_ (.Y(_0640_),
    .B(_0639_),
    .A_N(_0636_));
 sg13g2_a21oi_1 _3895_ (.A1(_1882_),
    .A2(_0635_),
    .Y(_0641_),
    .B1(_0640_));
 sg13g2_xnor2_1 _3896_ (.Y(_0642_),
    .A(net4),
    .B(_0641_));
 sg13g2_nand2_1 _3897_ (.Y(_0643_),
    .A(_1878_),
    .B(_0635_));
 sg13g2_nor2_1 _3898_ (.A(_1885_),
    .B(_1898_),
    .Y(_0644_));
 sg13g2_a21o_1 _3899_ (.A2(_0644_),
    .A1(_1793_),
    .B1(_0638_),
    .X(_0645_));
 sg13g2_a21oi_1 _3900_ (.A1(net688),
    .A2(_0636_),
    .Y(_0646_),
    .B1(_0645_));
 sg13g2_nand2_1 _3901_ (.Y(_0647_),
    .A(_0643_),
    .B(_0646_));
 sg13g2_xor2_1 _3902_ (.B(_0647_),
    .A(net3),
    .X(_0648_));
 sg13g2_inv_1 _3903_ (.Y(_0649_),
    .A(_0648_));
 sg13g2_nor2_1 _3904_ (.A(_0642_),
    .B(_0648_),
    .Y(_0650_));
 sg13g2_o21ai_1 _3905_ (.B1(_1943_),
    .Y(_0651_),
    .A1(net690),
    .A2(_1879_));
 sg13g2_o21ai_1 _3906_ (.B1(_0651_),
    .Y(_0652_),
    .A1(_1876_),
    .A2(_1904_));
 sg13g2_a22oi_1 _3907_ (.Y(_0653_),
    .B1(_1949_),
    .B2(_1904_),
    .A2(_1920_),
    .A1(_1907_));
 sg13g2_nor2_1 _3908_ (.A(_1793_),
    .B(_1899_),
    .Y(_0654_));
 sg13g2_nand2_1 _3909_ (.Y(_0655_),
    .A(_1897_),
    .B(_1941_));
 sg13g2_nand4_1 _3910_ (.B(_0652_),
    .C(_0653_),
    .A(_0639_),
    .Y(_0656_),
    .D(_0655_));
 sg13g2_nand2b_1 _3911_ (.Y(_0657_),
    .B(_0654_),
    .A_N(net688));
 sg13g2_nor3_2 _3912_ (.A(_1793_),
    .B(net686),
    .C(_1888_),
    .Y(_0658_));
 sg13g2_a21oi_1 _3913_ (.A1(net690),
    .A2(_0644_),
    .Y(_0659_),
    .B1(_0658_));
 sg13g2_a22oi_1 _3914_ (.Y(_0660_),
    .B1(_1904_),
    .B2(_1941_),
    .A2(_1897_),
    .A1(_1880_));
 sg13g2_a21oi_1 _3915_ (.A1(net690),
    .A2(net687),
    .Y(_0661_),
    .B1(net685));
 sg13g2_o21ai_1 _3916_ (.B1(_1876_),
    .Y(_0662_),
    .A1(_1941_),
    .A2(_0661_));
 sg13g2_nand3_1 _3917_ (.B(_1912_),
    .C(_1923_),
    .A(_1909_),
    .Y(_0663_));
 sg13g2_nand3_1 _3918_ (.B(net692),
    .C(_1920_),
    .A(_1793_),
    .Y(_0664_));
 sg13g2_nand4_1 _3919_ (.B(_0657_),
    .C(_0659_),
    .A(_1921_),
    .Y(_0665_),
    .D(_0660_));
 sg13g2_nand4_1 _3920_ (.B(_0662_),
    .C(_0663_),
    .A(_1913_),
    .Y(_0666_),
    .D(_0664_));
 sg13g2_nor4_2 _3921_ (.A(_1895_),
    .B(_0656_),
    .C(_0665_),
    .Y(_0667_),
    .D(_0666_));
 sg13g2_nor3_1 _3922_ (.A(net690),
    .B(_1879_),
    .C(_1898_),
    .Y(_0668_));
 sg13g2_a22oi_1 _3923_ (.Y(_0669_),
    .B1(_0645_),
    .B2(net688),
    .A2(_1889_),
    .A1(_1875_));
 sg13g2_nand2_1 _3924_ (.Y(_0670_),
    .A(_0643_),
    .B(_0669_));
 sg13g2_nor4_2 _3925_ (.A(_0636_),
    .B(_0667_),
    .C(_0668_),
    .Y(_0671_),
    .D(_0670_));
 sg13g2_xnor2_1 _3926_ (.Y(_0672_),
    .A(net2),
    .B(_0671_));
 sg13g2_inv_2 _3927_ (.Y(_0673_),
    .A(_0672_));
 sg13g2_a21oi_1 _3928_ (.A1(_0650_),
    .A2(_0673_),
    .Y(_0674_),
    .B1(net105));
 sg13g2_nor2b_2 _3929_ (.A(net138),
    .B_N(_0674_),
    .Y(_0675_));
 sg13g2_nor3_2 _3930_ (.A(_0642_),
    .B(_0649_),
    .C(_0673_),
    .Y(_0676_));
 sg13g2_and2_1 _3931_ (.A(\wirecube_top_inst.counter_h[5] ),
    .B(net700),
    .X(_0677_));
 sg13g2_xor2_1 _3932_ (.B(net700),
    .A(\wirecube_top_inst.counter_h[5] ),
    .X(_0678_));
 sg13g2_a21oi_1 _3933_ (.A1(\wirecube_top_inst.frame_cnt[5] ),
    .A2(_0678_),
    .Y(_0679_),
    .B1(_0677_));
 sg13g2_and2_1 _3934_ (.A(\wirecube_top_inst.counter_h[6] ),
    .B(net699),
    .X(_0680_));
 sg13g2_xor2_1 _3935_ (.B(net699),
    .A(\wirecube_top_inst.counter_h[6] ),
    .X(_0681_));
 sg13g2_xnor2_1 _3936_ (.Y(_0682_),
    .A(net693),
    .B(_0681_));
 sg13g2_nor2_1 _3937_ (.A(_0679_),
    .B(_0682_),
    .Y(_0683_));
 sg13g2_xor2_1 _3938_ (.B(_0682_),
    .A(_0679_),
    .X(_0684_));
 sg13g2_and2_1 _3939_ (.A(\wirecube_top_inst.counter_h[4] ),
    .B(net701),
    .X(_0685_));
 sg13g2_xor2_1 _3940_ (.B(net701),
    .A(\wirecube_top_inst.counter_h[4] ),
    .X(_0686_));
 sg13g2_a21oi_1 _3941_ (.A1(\wirecube_top_inst.frame_cnt[4] ),
    .A2(_0686_),
    .Y(_0687_),
    .B1(_0685_));
 sg13g2_xnor2_1 _3942_ (.Y(_0688_),
    .A(\wirecube_top_inst.frame_cnt[5] ),
    .B(_0678_));
 sg13g2_and2_1 _3943_ (.A(\wirecube_top_inst.counter_h[3] ),
    .B(net702),
    .X(_0689_));
 sg13g2_xor2_1 _3944_ (.B(net702),
    .A(\wirecube_top_inst.counter_h[3] ),
    .X(_0690_));
 sg13g2_xnor2_1 _3945_ (.Y(_0691_),
    .A(\wirecube_top_inst.frame_cnt[3] ),
    .B(_0690_));
 sg13g2_and2_1 _3946_ (.A(\wirecube_top_inst.counter_h[2] ),
    .B(net703),
    .X(_0692_));
 sg13g2_xor2_1 _3947_ (.B(net703),
    .A(\wirecube_top_inst.counter_h[2] ),
    .X(_0693_));
 sg13g2_a21oi_1 _3948_ (.A1(\wirecube_top_inst.frame_cnt[2] ),
    .A2(_0693_),
    .Y(_0694_),
    .B1(_0692_));
 sg13g2_xnor2_1 _3949_ (.Y(_0695_),
    .A(\wirecube_top_inst.frame_cnt[2] ),
    .B(_0693_));
 sg13g2_nand2b_1 _3950_ (.Y(_0696_),
    .B(_1872_),
    .A_N(\wirecube_top_inst.counter_h[0] ));
 sg13g2_nand2_1 _3951_ (.Y(_0697_),
    .A(_1873_),
    .B(_0696_));
 sg13g2_nand2_1 _3952_ (.Y(_0698_),
    .A(\wirecube_top_inst.frame_cnt[1] ),
    .B(net704));
 sg13g2_nand3_1 _3953_ (.B(\wirecube_top_inst.counter_h[1] ),
    .C(net704),
    .A(net698),
    .Y(_0699_));
 sg13g2_o21ai_1 _3954_ (.B1(_0695_),
    .Y(_0700_),
    .A1(_0697_),
    .A2(_0699_));
 sg13g2_nor2_1 _3955_ (.A(net698),
    .B(net704),
    .Y(_0701_));
 sg13g2_nand2_1 _3956_ (.Y(_0702_),
    .A(_0697_),
    .B(_0701_));
 sg13g2_a21oi_1 _3957_ (.A1(net698),
    .A2(net704),
    .Y(_0703_),
    .B1(\wirecube_top_inst.counter_h[1] ));
 sg13g2_o21ai_1 _3958_ (.B1(_0703_),
    .Y(_0704_),
    .A1(_0697_),
    .A2(_0701_));
 sg13g2_nand3_1 _3959_ (.B(_0702_),
    .C(_0704_),
    .A(_0700_),
    .Y(_0705_));
 sg13g2_o21ai_1 _3960_ (.B1(_0705_),
    .Y(_0706_),
    .A1(_0691_),
    .A2(_0694_));
 sg13g2_xnor2_1 _3961_ (.Y(_0707_),
    .A(\wirecube_top_inst.frame_cnt[4] ),
    .B(_0686_));
 sg13g2_a21oi_1 _3962_ (.A1(\wirecube_top_inst.frame_cnt[3] ),
    .A2(_0690_),
    .Y(_0708_),
    .B1(_0689_));
 sg13g2_a22oi_1 _3963_ (.Y(_0709_),
    .B1(_0707_),
    .B2(_0708_),
    .A2(_0694_),
    .A1(_0691_));
 sg13g2_nand2_1 _3964_ (.Y(_0710_),
    .A(_0706_),
    .B(_0709_));
 sg13g2_nor2_1 _3965_ (.A(_0687_),
    .B(_0688_),
    .Y(_0711_));
 sg13g2_nor2_1 _3966_ (.A(_0707_),
    .B(_0708_),
    .Y(_0712_));
 sg13g2_nor2_1 _3967_ (.A(_0711_),
    .B(_0712_),
    .Y(_0713_));
 sg13g2_a22oi_1 _3968_ (.Y(_0714_),
    .B1(_0710_),
    .B2(_0713_),
    .A2(_0688_),
    .A1(_0687_));
 sg13g2_a21oi_1 _3969_ (.A1(_0684_),
    .A2(_0714_),
    .Y(_0715_),
    .B1(_0683_));
 sg13g2_a21oi_1 _3970_ (.A1(net693),
    .A2(_0681_),
    .Y(_0716_),
    .B1(_0680_));
 sg13g2_xnor2_1 _3971_ (.Y(_0717_),
    .A(_0060_),
    .B(\wirecube_top_inst.counter_h[7] ));
 sg13g2_xnor2_1 _3972_ (.Y(_0718_),
    .A(\wirecube_top_inst.counter_v[7] ),
    .B(_0717_));
 sg13g2_xnor2_1 _3973_ (.Y(_0719_),
    .A(_0716_),
    .B(_0718_));
 sg13g2_xnor2_1 _3974_ (.Y(_0720_),
    .A(_0715_),
    .B(_0719_));
 sg13g2_and2_1 _3975_ (.A(_0650_),
    .B(_0672_),
    .X(_0721_));
 sg13g2_inv_1 _3976_ (.Y(_0722_),
    .A(_0721_));
 sg13g2_nand2_1 _3977_ (.Y(_0723_),
    .A(_0642_),
    .B(_0649_));
 sg13g2_nor2_2 _3978_ (.A(_0672_),
    .B(_0723_),
    .Y(_0724_));
 sg13g2_and2_1 _3979_ (.A(net694),
    .B(\wirecube_top_inst.counter_v[5] ),
    .X(_0725_));
 sg13g2_xor2_1 _3980_ (.B(\wirecube_top_inst.counter_v[5] ),
    .A(net694),
    .X(_0726_));
 sg13g2_and2_1 _3981_ (.A(net695),
    .B(net701),
    .X(_0727_));
 sg13g2_and2_1 _3982_ (.A(\wirecube_top_inst.frame_cnt[3] ),
    .B(net702),
    .X(_0728_));
 sg13g2_and2_1 _3983_ (.A(net697),
    .B(net703),
    .X(_0729_));
 sg13g2_xor2_1 _3984_ (.B(net703),
    .A(net697),
    .X(_0730_));
 sg13g2_xnor2_1 _3985_ (.Y(_0731_),
    .A(net698),
    .B(net704));
 sg13g2_o21ai_1 _3986_ (.B1(_0698_),
    .Y(_0732_),
    .A1(_1872_),
    .A2(_0701_));
 sg13g2_a21o_1 _3987_ (.A2(_0732_),
    .A1(_0730_),
    .B1(_0729_),
    .X(_0733_));
 sg13g2_xor2_1 _3988_ (.B(net702),
    .A(net696),
    .X(_0734_));
 sg13g2_a21o_1 _3989_ (.A2(_0734_),
    .A1(_0733_),
    .B1(_0728_),
    .X(_0735_));
 sg13g2_xor2_1 _3990_ (.B(net701),
    .A(net695),
    .X(_0736_));
 sg13g2_a21o_1 _3991_ (.A2(_0736_),
    .A1(_0735_),
    .B1(_0727_),
    .X(_0737_));
 sg13g2_a21oi_1 _3992_ (.A1(_0726_),
    .A2(_0737_),
    .Y(_0738_),
    .B1(_0725_));
 sg13g2_xnor2_1 _3993_ (.Y(_0739_),
    .A(net693),
    .B(net699));
 sg13g2_xnor2_1 _3994_ (.Y(_0740_),
    .A(_0738_),
    .B(_0739_));
 sg13g2_inv_1 _3995_ (.Y(_0741_),
    .A(_0740_));
 sg13g2_a221oi_1 _3996_ (.B2(_0740_),
    .C1(_0721_),
    .B1(_0724_),
    .A1(_0676_),
    .Y(_0742_),
    .A2(_0720_));
 sg13g2_inv_1 _3997_ (.Y(_0743_),
    .A(_0742_));
 sg13g2_nand2_1 _3998_ (.Y(_0744_),
    .A(_0648_),
    .B(_0673_));
 sg13g2_nand3_1 _3999_ (.B(_0648_),
    .C(_0673_),
    .A(_0642_),
    .Y(_0745_));
 sg13g2_nand3_1 _4000_ (.B(_0648_),
    .C(_0672_),
    .A(_0642_),
    .Y(_0746_));
 sg13g2_inv_1 _4001_ (.Y(_0747_),
    .A(_0746_));
 sg13g2_nor2_2 _4002_ (.A(_0673_),
    .B(_0723_),
    .Y(_0748_));
 sg13g2_xor2_1 _4003_ (.B(\wirecube_top_inst.edge_function_inst.pixel_x_i[0] ),
    .A(\wirecube_top_inst.edge_function_inst.pixel_y_i[0] ),
    .X(_0749_));
 sg13g2_xnor2_1 _4004_ (.Y(_0750_),
    .A(_0073_),
    .B(_0749_));
 sg13g2_a22oi_1 _4005_ (.Y(_0751_),
    .B1(_0748_),
    .B2(_0750_),
    .A2(_0747_),
    .A1(_1874_));
 sg13g2_o21ai_1 _4006_ (.B1(_0751_),
    .Y(_0752_),
    .A1(_0073_),
    .A2(_0745_));
 sg13g2_o21ai_1 _4007_ (.B1(_0675_),
    .Y(_0753_),
    .A1(_0743_),
    .A2(_0752_));
 sg13g2_a21oi_1 _4008_ (.A1(net686),
    .A2(_1923_),
    .Y(_0754_),
    .B1(_1892_));
 sg13g2_nand2_1 _4009_ (.Y(_0755_),
    .A(_1881_),
    .B(_0754_));
 sg13g2_or2_1 _4010_ (.X(_0756_),
    .B(_1929_),
    .A(_1889_));
 sg13g2_nor3_1 _4011_ (.A(net691),
    .B(_1804_),
    .C(_1892_),
    .Y(_0757_));
 sg13g2_a22oi_1 _4012_ (.Y(_0758_),
    .B1(_0757_),
    .B2(net686),
    .A2(_0756_),
    .A1(_1804_));
 sg13g2_nand2_1 _4013_ (.Y(_0759_),
    .A(net692),
    .B(_0756_));
 sg13g2_nor2_1 _4014_ (.A(_1793_),
    .B(net692),
    .Y(_0760_));
 sg13g2_nand3_1 _4015_ (.B(_1891_),
    .C(_0760_),
    .A(net686),
    .Y(_0761_));
 sg13g2_nand2_1 _4016_ (.Y(_0762_),
    .A(_0759_),
    .B(_0761_));
 sg13g2_nor3_1 _4017_ (.A(_1813_),
    .B(_1892_),
    .C(_1907_),
    .Y(_0763_));
 sg13g2_nor2_1 _4018_ (.A(_1894_),
    .B(_0763_),
    .Y(_0764_));
 sg13g2_nor2_1 _4019_ (.A(_1874_),
    .B(_0764_),
    .Y(_0765_));
 sg13g2_nor4_1 _4020_ (.A(_0654_),
    .B(_0658_),
    .C(_0762_),
    .D(_0765_),
    .Y(_0766_));
 sg13g2_and3_1 _4021_ (.X(_0767_),
    .A(_0755_),
    .B(_0758_),
    .C(_0766_));
 sg13g2_xor2_1 _4022_ (.B(_0767_),
    .A(net7),
    .X(_0768_));
 sg13g2_nor2b_1 _4023_ (.A(_0762_),
    .B_N(_0764_),
    .Y(_0769_));
 sg13g2_nor2_1 _4024_ (.A(_1874_),
    .B(_0758_),
    .Y(_0770_));
 sg13g2_a221oi_1 _4025_ (.B2(_1904_),
    .C1(_1932_),
    .B1(_1941_),
    .A1(_1882_),
    .Y(_0771_),
    .A2(_1909_));
 sg13g2_o21ai_1 _4026_ (.B1(net688),
    .Y(_0772_),
    .A1(_1909_),
    .A2(_0658_));
 sg13g2_nor3_1 _4027_ (.A(_1881_),
    .B(_1898_),
    .C(_0760_),
    .Y(_0773_));
 sg13g2_a21oi_1 _4028_ (.A1(net689),
    .A2(_1914_),
    .Y(_0774_),
    .B1(_0773_));
 sg13g2_nand4_1 _4029_ (.B(_1924_),
    .C(_0755_),
    .A(_1921_),
    .Y(_0775_),
    .D(_0774_));
 sg13g2_a221oi_1 _4030_ (.B2(_1925_),
    .C1(_0644_),
    .B1(_1881_),
    .A1(_1813_),
    .Y(_0776_),
    .A2(_1876_));
 sg13g2_a21oi_1 _4031_ (.A1(_1876_),
    .A2(_1949_),
    .Y(_0777_),
    .B1(_1897_));
 sg13g2_a221oi_1 _4032_ (.B2(_1923_),
    .C1(_1949_),
    .B1(_1912_),
    .A1(_1878_),
    .Y(_0778_),
    .A2(_1906_));
 sg13g2_or2_1 _4033_ (.X(_0779_),
    .B(_0778_),
    .A(_0777_));
 sg13g2_nand4_1 _4034_ (.B(_0772_),
    .C(_0776_),
    .A(_0771_),
    .Y(_0780_),
    .D(_0779_));
 sg13g2_nor4_1 _4035_ (.A(_0656_),
    .B(_0770_),
    .C(_0775_),
    .D(_0780_),
    .Y(_0781_));
 sg13g2_o21ai_1 _4036_ (.B1(_0781_),
    .Y(_0782_),
    .A1(_1875_),
    .A2(_0769_));
 sg13g2_xor2_1 _4037_ (.B(_0782_),
    .A(net5),
    .X(_0783_));
 sg13g2_nand3_1 _4038_ (.B(_0758_),
    .C(_0764_),
    .A(_0755_),
    .Y(_0784_));
 sg13g2_and2_1 _4039_ (.A(_1874_),
    .B(_0784_),
    .X(_0785_));
 sg13g2_a21oi_1 _4040_ (.A1(_1875_),
    .A2(_0762_),
    .Y(_0786_),
    .B1(_0785_));
 sg13g2_and2_1 _4041_ (.A(_0659_),
    .B(_0786_),
    .X(_0787_));
 sg13g2_xnor2_1 _4042_ (.Y(_0788_),
    .A(net6),
    .B(_0787_));
 sg13g2_inv_1 _4043_ (.Y(_0789_),
    .A(_0788_));
 sg13g2_or2_1 _4044_ (.X(_0790_),
    .B(_0788_),
    .A(_0783_));
 sg13g2_nand2b_1 _4045_ (.Y(_0791_),
    .B(_0768_),
    .A_N(_0790_));
 sg13g2_and2_1 _4046_ (.A(net171),
    .B(_0791_),
    .X(_0792_));
 sg13g2_nor2_2 _4047_ (.A(_0768_),
    .B(_0790_),
    .Y(_0793_));
 sg13g2_nand2_1 _4048_ (.Y(_0794_),
    .A(_0740_),
    .B(_0793_));
 sg13g2_nand2_1 _4049_ (.Y(_0795_),
    .A(_0768_),
    .B(_0783_));
 sg13g2_nor2_1 _4050_ (.A(_0720_),
    .B(_0789_),
    .Y(_0796_));
 sg13g2_or2_1 _4051_ (.X(_0797_),
    .B(_0795_),
    .A(_0788_));
 sg13g2_o21ai_1 _4052_ (.B1(_0794_),
    .Y(_0798_),
    .A1(_0795_),
    .A2(_0796_));
 sg13g2_nand3b_1 _4053_ (.B(_0783_),
    .C(_0789_),
    .Y(_0799_),
    .A_N(_0768_));
 sg13g2_nand2b_1 _4054_ (.Y(_0800_),
    .B(_0750_),
    .A_N(_0799_));
 sg13g2_nand2_1 _4055_ (.Y(_0801_),
    .A(_0783_),
    .B(_0788_));
 sg13g2_or2_2 _4056_ (.X(_0802_),
    .B(_0801_),
    .A(_0768_));
 sg13g2_inv_1 _4057_ (.Y(_0803_),
    .A(_0802_));
 sg13g2_nor3_2 _4058_ (.A(_0768_),
    .B(_0783_),
    .C(_0789_),
    .Y(_0804_));
 sg13g2_a22oi_1 _4059_ (.Y(_0805_),
    .B1(_0804_),
    .B2(net697),
    .A2(_0803_),
    .A1(_1874_));
 sg13g2_nand2_1 _4060_ (.Y(_0806_),
    .A(_0800_),
    .B(_0805_));
 sg13g2_o21ai_1 _4061_ (.B1(_0792_),
    .Y(_0807_),
    .A1(_0798_),
    .A2(_0806_));
 sg13g2_a21oi_1 _4062_ (.A1(_0753_),
    .A2(_0807_),
    .Y(_0004_),
    .B1(_0633_));
 sg13g2_xnor2_1 _4063_ (.Y(_0808_),
    .A(_1872_),
    .B(_0731_));
 sg13g2_xor2_1 _4064_ (.B(\wirecube_top_inst.edge_function_inst.pixel_x_i[1] ),
    .A(\wirecube_top_inst.edge_function_inst.pixel_y_i[1] ),
    .X(_0809_));
 sg13g2_nand2_1 _4065_ (.Y(_0810_),
    .A(net696),
    .B(_0809_));
 sg13g2_xnor2_1 _4066_ (.Y(_0811_),
    .A(net696),
    .B(_0809_));
 sg13g2_nand2_1 _4067_ (.Y(_0812_),
    .A(net697),
    .B(_0749_));
 sg13g2_xor2_1 _4068_ (.B(_0812_),
    .A(_0811_),
    .X(_0813_));
 sg13g2_inv_1 _4069_ (.Y(_0814_),
    .A(_0813_));
 sg13g2_o21ai_1 _4070_ (.B1(_0797_),
    .Y(_0815_),
    .A1(_0799_),
    .A2(_0814_));
 sg13g2_a21oi_1 _4071_ (.A1(net696),
    .A2(_0804_),
    .Y(_0816_),
    .B1(_0815_));
 sg13g2_o21ai_1 _4072_ (.B1(_0816_),
    .Y(_0817_),
    .A1(_0802_),
    .A2(_0808_));
 sg13g2_nor2_1 _4073_ (.A(_0070_),
    .B(_0745_),
    .Y(_0818_));
 sg13g2_a221oi_1 _4074_ (.B2(_0813_),
    .C1(_0818_),
    .B1(_0748_),
    .A1(_0650_),
    .Y(_0819_),
    .A2(_0672_));
 sg13g2_o21ai_1 _4075_ (.B1(_0819_),
    .Y(_0820_),
    .A1(_0746_),
    .A2(_0808_));
 sg13g2_a22oi_1 _4076_ (.Y(_0821_),
    .B1(_0820_),
    .B2(_0675_),
    .A2(_0817_),
    .A1(_0792_));
 sg13g2_nor2_1 _4077_ (.A(_0633_),
    .B(_0821_),
    .Y(_0005_));
 sg13g2_xnor2_1 _4078_ (.Y(_0822_),
    .A(_0684_),
    .B(_0714_));
 sg13g2_nand2_1 _4079_ (.Y(_0823_),
    .A(_0720_),
    .B(_0822_));
 sg13g2_o21ai_1 _4080_ (.B1(_0810_),
    .Y(_0824_),
    .A1(_0811_),
    .A2(_0812_));
 sg13g2_xor2_1 _4081_ (.B(\wirecube_top_inst.edge_function_inst.pixel_x_i[2] ),
    .A(\wirecube_top_inst.edge_function_inst.pixel_y_i[2] ),
    .X(_0825_));
 sg13g2_xor2_1 _4082_ (.B(_0825_),
    .A(net695),
    .X(_0826_));
 sg13g2_xor2_1 _4083_ (.B(_0826_),
    .A(_0824_),
    .X(_0827_));
 sg13g2_nand2b_1 _4084_ (.Y(_0828_),
    .B(_1836_),
    .A_N(_0745_));
 sg13g2_o21ai_1 _4085_ (.B1(_0722_),
    .Y(_0829_),
    .A1(_0642_),
    .A2(_0744_));
 sg13g2_xnor2_1 _4086_ (.Y(_0830_),
    .A(_0730_),
    .B(_0732_));
 sg13g2_or2_1 _4087_ (.X(_0831_),
    .B(_0830_),
    .A(_0746_));
 sg13g2_a21oi_1 _4088_ (.A1(_0748_),
    .A2(_0827_),
    .Y(_0832_),
    .B1(_0829_));
 sg13g2_xnor2_1 _4089_ (.Y(_0833_),
    .A(_0726_),
    .B(_0737_));
 sg13g2_nand2_1 _4090_ (.Y(_0834_),
    .A(_0740_),
    .B(_0833_));
 sg13g2_a22oi_1 _4091_ (.Y(_0835_),
    .B1(_0834_),
    .B2(_0724_),
    .A2(_0823_),
    .A1(_0676_));
 sg13g2_nand4_1 _4092_ (.B(_0831_),
    .C(_0832_),
    .A(_0828_),
    .Y(_0836_),
    .D(_0835_));
 sg13g2_a21oi_1 _4093_ (.A1(_0674_),
    .A2(_0836_),
    .Y(_0837_),
    .B1(net138));
 sg13g2_nand3_1 _4094_ (.B(_0783_),
    .C(_0788_),
    .A(_0768_),
    .Y(_0838_));
 sg13g2_a21oi_1 _4095_ (.A1(_0720_),
    .A2(_0822_),
    .Y(_0839_),
    .B1(_0838_));
 sg13g2_nand2b_1 _4096_ (.Y(_0840_),
    .B(_0827_),
    .A_N(_0799_));
 sg13g2_nand3_1 _4097_ (.B(_0790_),
    .C(_0801_),
    .A(_0768_),
    .Y(_0841_));
 sg13g2_nand2_1 _4098_ (.Y(_0842_),
    .A(net171),
    .B(_0841_));
 sg13g2_o21ai_1 _4099_ (.B1(_0840_),
    .Y(_0843_),
    .A1(_0802_),
    .A2(_0830_));
 sg13g2_a22oi_1 _4100_ (.Y(_0844_),
    .B1(_0834_),
    .B2(_0793_),
    .A2(_0804_),
    .A1(net695));
 sg13g2_inv_1 _4101_ (.Y(_0845_),
    .A(_0844_));
 sg13g2_nor4_1 _4102_ (.A(_0839_),
    .B(_0842_),
    .C(_0843_),
    .D(_0845_),
    .Y(_0846_));
 sg13g2_nor3_1 _4103_ (.A(_0633_),
    .B(_0837_),
    .C(_0846_),
    .Y(_0006_));
 sg13g2_xnor2_1 _4104_ (.Y(_0847_),
    .A(_0733_),
    .B(_0734_));
 sg13g2_nor2_1 _4105_ (.A(_0746_),
    .B(_0847_),
    .Y(_0848_));
 sg13g2_nand2b_1 _4106_ (.Y(_0849_),
    .B(_1834_),
    .A_N(_0745_));
 sg13g2_a22oi_1 _4107_ (.Y(_0850_),
    .B1(_0826_),
    .B2(_0824_),
    .A2(_0825_),
    .A1(_1836_));
 sg13g2_xor2_1 _4108_ (.B(\wirecube_top_inst.edge_function_inst.pixel_x_i[3] ),
    .A(\wirecube_top_inst.edge_function_inst.pixel_y_i[3] ),
    .X(_0851_));
 sg13g2_xnor2_1 _4109_ (.Y(_0852_),
    .A(net694),
    .B(_0851_));
 sg13g2_xor2_1 _4110_ (.B(_0852_),
    .A(_0850_),
    .X(_0853_));
 sg13g2_a21oi_1 _4111_ (.A1(_0748_),
    .A2(_0853_),
    .Y(_0854_),
    .B1(_0829_));
 sg13g2_nand2b_1 _4112_ (.Y(_0855_),
    .B(_0676_),
    .A_N(_0720_));
 sg13g2_a21oi_1 _4113_ (.A1(_0724_),
    .A2(_0741_),
    .Y(_0856_),
    .B1(_0848_));
 sg13g2_nand4_1 _4114_ (.B(_0854_),
    .C(_0855_),
    .A(_0849_),
    .Y(_0857_),
    .D(_0856_));
 sg13g2_a21oi_1 _4115_ (.A1(_0674_),
    .A2(_0857_),
    .Y(_0858_),
    .B1(net138));
 sg13g2_nor2_1 _4116_ (.A(_0720_),
    .B(_0838_),
    .Y(_0859_));
 sg13g2_a22oi_1 _4117_ (.Y(_0860_),
    .B1(_0804_),
    .B2(net694),
    .A2(_0793_),
    .A1(_0741_));
 sg13g2_nand2b_1 _4118_ (.Y(_0861_),
    .B(_0853_),
    .A_N(_0799_));
 sg13g2_or2_1 _4119_ (.X(_0862_),
    .B(_0847_),
    .A(_0802_));
 sg13g2_nand3_1 _4120_ (.B(_0861_),
    .C(_0862_),
    .A(_0860_),
    .Y(_0863_));
 sg13g2_nor3_1 _4121_ (.A(_0842_),
    .B(_0859_),
    .C(_0863_),
    .Y(_0864_));
 sg13g2_nor3_1 _4122_ (.A(_0633_),
    .B(_0858_),
    .C(_0864_),
    .Y(_0007_));
 sg13g2_xnor2_1 _4123_ (.Y(_0865_),
    .A(_0735_),
    .B(_0736_));
 sg13g2_nor2_1 _4124_ (.A(_0746_),
    .B(_0865_),
    .Y(_0866_));
 sg13g2_nand2_1 _4125_ (.Y(_0867_),
    .A(_1834_),
    .B(_0851_));
 sg13g2_o21ai_1 _4126_ (.B1(_0867_),
    .Y(_0868_),
    .A1(_0850_),
    .A2(_0852_));
 sg13g2_xnor2_1 _4127_ (.Y(_0869_),
    .A(\wirecube_top_inst.edge_function_inst.pixel_y_i[4] ),
    .B(\wirecube_top_inst.edge_function_inst.pixel_x_i[4] ));
 sg13g2_nor2_1 _4128_ (.A(_0071_),
    .B(_0869_),
    .Y(_0870_));
 sg13g2_xor2_1 _4129_ (.B(_0869_),
    .A(_0071_),
    .X(_0871_));
 sg13g2_xor2_1 _4130_ (.B(_0871_),
    .A(_0868_),
    .X(_0872_));
 sg13g2_a21oi_1 _4131_ (.A1(_0748_),
    .A2(_0872_),
    .Y(_0873_),
    .B1(_0866_));
 sg13g2_o21ai_1 _4132_ (.B1(_0873_),
    .Y(_0874_),
    .A1(_0071_),
    .A2(_0745_));
 sg13g2_o21ai_1 _4133_ (.B1(_0675_),
    .Y(_0875_),
    .A1(_0743_),
    .A2(_0874_));
 sg13g2_nor2b_1 _4134_ (.A(_0799_),
    .B_N(_0872_),
    .Y(_0876_));
 sg13g2_a21oi_1 _4135_ (.A1(net693),
    .A2(_0804_),
    .Y(_0877_),
    .B1(_0876_));
 sg13g2_o21ai_1 _4136_ (.B1(_0877_),
    .Y(_0878_),
    .A1(_0802_),
    .A2(_0865_));
 sg13g2_o21ai_1 _4137_ (.B1(_0792_),
    .Y(_0879_),
    .A1(_0798_),
    .A2(_0878_));
 sg13g2_a21oi_1 _4138_ (.A1(_0875_),
    .A2(_0879_),
    .Y(_0008_),
    .B1(_0633_));
 sg13g2_xnor2_1 _4139_ (.Y(_0880_),
    .A(_0720_),
    .B(_0822_));
 sg13g2_o21ai_1 _4140_ (.B1(_0722_),
    .Y(_0881_),
    .A1(_0060_),
    .A2(_0745_));
 sg13g2_a21oi_1 _4141_ (.A1(_0868_),
    .A2(_0871_),
    .Y(_0882_),
    .B1(_0870_));
 sg13g2_xnor2_1 _4142_ (.Y(_0883_),
    .A(\wirecube_top_inst.edge_function_inst.pixel_y_i[5] ),
    .B(\wirecube_top_inst.edge_function_inst.pixel_x_i[5] ));
 sg13g2_xnor2_1 _4143_ (.Y(_0884_),
    .A(_0060_),
    .B(_0883_));
 sg13g2_xnor2_1 _4144_ (.Y(_0885_),
    .A(_0882_),
    .B(_0884_));
 sg13g2_nand2b_1 _4145_ (.Y(_0886_),
    .B(_0748_),
    .A_N(_0885_));
 sg13g2_o21ai_1 _4146_ (.B1(_0886_),
    .Y(_0887_),
    .A1(_0746_),
    .A2(_0833_));
 sg13g2_nor2_1 _4147_ (.A(_0881_),
    .B(_0887_),
    .Y(_0888_));
 sg13g2_xnor2_1 _4148_ (.Y(_0889_),
    .A(_0740_),
    .B(_0833_));
 sg13g2_a22oi_1 _4149_ (.Y(_0890_),
    .B1(_0889_),
    .B2(_0724_),
    .A2(_0880_),
    .A1(_0676_));
 sg13g2_nand2_1 _4150_ (.Y(_0891_),
    .A(_0888_),
    .B(_0890_));
 sg13g2_nor2b_1 _4151_ (.A(_0838_),
    .B_N(_0880_),
    .Y(_0892_));
 sg13g2_o21ai_1 _4152_ (.B1(_0797_),
    .Y(_0893_),
    .A1(_0799_),
    .A2(_0885_));
 sg13g2_nor2_1 _4153_ (.A(_0802_),
    .B(_0833_),
    .Y(_0894_));
 sg13g2_a21oi_1 _4154_ (.A1(net691),
    .A2(_0804_),
    .Y(_0895_),
    .B1(_0894_));
 sg13g2_a21oi_1 _4155_ (.A1(_0793_),
    .A2(_0889_),
    .Y(_0896_),
    .B1(_0892_));
 sg13g2_nand3b_1 _4156_ (.B(_0895_),
    .C(_0896_),
    .Y(_0897_),
    .A_N(_0893_));
 sg13g2_a22oi_1 _4157_ (.Y(_0898_),
    .B1(_0897_),
    .B2(net138),
    .A2(_0891_),
    .A1(_0675_));
 sg13g2_nor2_1 _4158_ (.A(_0633_),
    .B(_0898_),
    .Y(_0009_));
 sg13g2_nand2_1 _4159_ (.Y(_0899_),
    .A(\wirecube_top_inst.edge_function_inst.term3[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term2[0] ));
 sg13g2_nand2_2 _4160_ (.Y(_0900_),
    .A(\wirecube_top_inst.edge_function_inst.term1[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[0] ));
 sg13g2_nand2b_1 _4161_ (.Y(_0901_),
    .B(_0900_),
    .A_N(_0899_));
 sg13g2_nand2b_1 _4162_ (.Y(_0902_),
    .B(_0899_),
    .A_N(_0900_));
 sg13g2_nand2_1 _4163_ (.Y(_0014_),
    .A(_0901_),
    .B(_0902_));
 sg13g2_nand2_2 _4164_ (.Y(_0903_),
    .A(\wirecube_top_inst.edge_function_inst.term2[1] ),
    .B(net705));
 sg13g2_nor2_2 _4165_ (.A(_0899_),
    .B(_0903_),
    .Y(_0904_));
 sg13g2_a22oi_1 _4166_ (.Y(_0905_),
    .B1(net705),
    .B2(\wirecube_top_inst.edge_function_inst.term2[0] ),
    .A2(\wirecube_top_inst.edge_function_inst.term2[1] ),
    .A1(\wirecube_top_inst.edge_function_inst.term3[0] ));
 sg13g2_nor2_1 _4167_ (.A(_0904_),
    .B(_0905_),
    .Y(_0906_));
 sg13g2_nand2_1 _4168_ (.Y(_0907_),
    .A(\wirecube_top_inst.edge_function_inst.term0[1] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[1] ));
 sg13g2_nor2_2 _4169_ (.A(_0900_),
    .B(_0907_),
    .Y(_0908_));
 sg13g2_a22oi_1 _4170_ (.Y(_0909_),
    .B1(\wirecube_top_inst.edge_function_inst.term1[1] ),
    .B2(\wirecube_top_inst.edge_function_inst.term0[0] ),
    .A2(\wirecube_top_inst.edge_function_inst.term0[1] ),
    .A1(\wirecube_top_inst.edge_function_inst.term1[0] ));
 sg13g2_nor2_2 _4171_ (.A(_0908_),
    .B(_0909_),
    .Y(_0910_));
 sg13g2_nor2b_1 _4172_ (.A(_0906_),
    .B_N(_0910_),
    .Y(_0911_));
 sg13g2_inv_1 _4173_ (.Y(_0912_),
    .A(_0911_));
 sg13g2_nor2b_1 _4174_ (.A(_0910_),
    .B_N(_0906_),
    .Y(_0913_));
 sg13g2_inv_1 _4175_ (.Y(_0914_),
    .A(_0913_));
 sg13g2_nor2_1 _4176_ (.A(_0911_),
    .B(_0913_),
    .Y(_0915_));
 sg13g2_nand2_1 _4177_ (.Y(_0916_),
    .A(\wirecube_top_inst.edge_function_inst.term0[6] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[4] ));
 sg13g2_nand2_1 _4178_ (.Y(_0917_),
    .A(\wirecube_top_inst.edge_function_inst.term1[5] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[4] ));
 sg13g2_nand2_2 _4179_ (.Y(_0918_),
    .A(\wirecube_top_inst.edge_function_inst.term0[5] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[5] ));
 sg13g2_nand2_1 _4180_ (.Y(_0919_),
    .A(\wirecube_top_inst.edge_function_inst.term1[6] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[4] ));
 sg13g2_or2_1 _4181_ (.X(_0920_),
    .B(_0919_),
    .A(_0918_));
 sg13g2_xor2_1 _4182_ (.B(_0919_),
    .A(_0918_),
    .X(_0921_));
 sg13g2_nand2b_1 _4183_ (.Y(_0922_),
    .B(_0921_),
    .A_N(_0916_));
 sg13g2_xor2_1 _4184_ (.B(_0921_),
    .A(_0916_),
    .X(_0923_));
 sg13g2_nand2_1 _4185_ (.Y(_0924_),
    .A(\wirecube_top_inst.edge_function_inst.term1[5] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[3] ));
 sg13g2_nand2_1 _4186_ (.Y(_0925_),
    .A(\wirecube_top_inst.edge_function_inst.term1[6] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[3] ));
 sg13g2_or2_1 _4187_ (.X(_0926_),
    .B(_0924_),
    .A(_0919_));
 sg13g2_nand2_1 _4188_ (.Y(_0927_),
    .A(\wirecube_top_inst.edge_function_inst.term0[5] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[4] ));
 sg13g2_xor2_1 _4189_ (.B(_0925_),
    .A(_0917_),
    .X(_0928_));
 sg13g2_nand2b_1 _4190_ (.Y(_0929_),
    .B(_0928_),
    .A_N(_0927_));
 sg13g2_a21oi_1 _4191_ (.A1(_0926_),
    .A2(_0929_),
    .Y(_0930_),
    .B1(_0923_));
 sg13g2_inv_1 _4192_ (.Y(_0931_),
    .A(_0930_));
 sg13g2_nand3_1 _4193_ (.B(_0926_),
    .C(_0929_),
    .A(_0923_),
    .Y(_0932_));
 sg13g2_nor2b_1 _4194_ (.A(_0930_),
    .B_N(_0932_),
    .Y(_0933_));
 sg13g2_nand2_1 _4195_ (.Y(_0934_),
    .A(\wirecube_top_inst.edge_function_inst.term1[5] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[2] ));
 sg13g2_nand2_1 _4196_ (.Y(_0935_),
    .A(\wirecube_top_inst.edge_function_inst.term1[6] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[2] ));
 sg13g2_or2_1 _4197_ (.X(_0936_),
    .B(_0934_),
    .A(_0925_));
 sg13g2_nand2_1 _4198_ (.Y(_0937_),
    .A(\wirecube_top_inst.edge_function_inst.term0[4] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[4] ));
 sg13g2_xnor2_1 _4199_ (.Y(_0938_),
    .A(_0924_),
    .B(_0935_));
 sg13g2_o21ai_1 _4200_ (.B1(_0936_),
    .Y(_0939_),
    .A1(_0937_),
    .A2(_0938_));
 sg13g2_xnor2_1 _4201_ (.Y(_0940_),
    .A(_0927_),
    .B(_0928_));
 sg13g2_and2_1 _4202_ (.A(_0939_),
    .B(_0940_),
    .X(_0941_));
 sg13g2_nand2_1 _4203_ (.Y(_0942_),
    .A(\wirecube_top_inst.edge_function_inst.term0[6] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[3] ));
 sg13g2_xnor2_1 _4204_ (.Y(_0943_),
    .A(_0939_),
    .B(_0940_));
 sg13g2_nor2_1 _4205_ (.A(_0942_),
    .B(_0943_),
    .Y(_0944_));
 sg13g2_o21ai_1 _4206_ (.B1(_0933_),
    .Y(_0945_),
    .A1(_0941_),
    .A2(_0944_));
 sg13g2_or3_1 _4207_ (.A(_0933_),
    .B(_0941_),
    .C(_0944_),
    .X(_0946_));
 sg13g2_and2_1 _4208_ (.A(_0945_),
    .B(_0946_),
    .X(_0947_));
 sg13g2_nand2_2 _4209_ (.Y(_0948_),
    .A(\wirecube_top_inst.edge_function_inst.term1[5] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[1] ));
 sg13g2_nand2_1 _4210_ (.Y(_0949_),
    .A(\wirecube_top_inst.edge_function_inst.term1[6] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[1] ));
 sg13g2_nand2_1 _4211_ (.Y(_0950_),
    .A(\wirecube_top_inst.edge_function_inst.term1[4] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[3] ));
 sg13g2_xor2_1 _4212_ (.B(_0949_),
    .A(_0934_),
    .X(_0951_));
 sg13g2_nand2b_1 _4213_ (.Y(_0952_),
    .B(_0951_),
    .A_N(_0950_));
 sg13g2_o21ai_1 _4214_ (.B1(_0952_),
    .Y(_0953_),
    .A1(_0935_),
    .A2(_0948_));
 sg13g2_xor2_1 _4215_ (.B(_0938_),
    .A(_0937_),
    .X(_0954_));
 sg13g2_nand2_1 _4216_ (.Y(_0955_),
    .A(_0953_),
    .B(_0954_));
 sg13g2_a22oi_1 _4217_ (.Y(_0956_),
    .B1(\wirecube_top_inst.edge_function_inst.term1[2] ),
    .B2(\wirecube_top_inst.edge_function_inst.term0[6] ),
    .A2(\wirecube_top_inst.edge_function_inst.term1[3] ),
    .A1(\wirecube_top_inst.edge_function_inst.term0[5] ));
 sg13g2_nand2_1 _4218_ (.Y(_0957_),
    .A(\wirecube_top_inst.edge_function_inst.term0[5] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[2] ));
 sg13g2_or2_1 _4219_ (.X(_0958_),
    .B(_0957_),
    .A(_0942_));
 sg13g2_nand2b_1 _4220_ (.Y(_0959_),
    .B(_0958_),
    .A_N(_0956_));
 sg13g2_xnor2_1 _4221_ (.Y(_0960_),
    .A(_0953_),
    .B(_0954_));
 sg13g2_o21ai_1 _4222_ (.B1(_0955_),
    .Y(_0961_),
    .A1(_0959_),
    .A2(_0960_));
 sg13g2_xor2_1 _4223_ (.B(_0943_),
    .A(_0942_),
    .X(_0962_));
 sg13g2_nand2_1 _4224_ (.Y(_0963_),
    .A(_0961_),
    .B(_0962_));
 sg13g2_xnor2_1 _4225_ (.Y(_0964_),
    .A(_0961_),
    .B(_0962_));
 sg13g2_o21ai_1 _4226_ (.B1(_0963_),
    .Y(_0965_),
    .A1(_0958_),
    .A2(_0964_));
 sg13g2_nand2_1 _4227_ (.Y(_0966_),
    .A(_0947_),
    .B(_0965_));
 sg13g2_nand2_1 _4228_ (.Y(_0967_),
    .A(\wirecube_top_inst.edge_function_inst.term1[6] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[6] ));
 sg13g2_nor2_1 _4229_ (.A(_0918_),
    .B(_0967_),
    .Y(_0968_));
 sg13g2_a22oi_1 _4230_ (.Y(_0969_),
    .B1(\wirecube_top_inst.edge_function_inst.term1[5] ),
    .B2(\wirecube_top_inst.edge_function_inst.term0[6] ),
    .A2(\wirecube_top_inst.edge_function_inst.term0[5] ),
    .A1(\wirecube_top_inst.edge_function_inst.term1[6] ));
 sg13g2_nor2_1 _4231_ (.A(_0968_),
    .B(_0969_),
    .Y(_0970_));
 sg13g2_and2_1 _4232_ (.A(_0920_),
    .B(_0922_),
    .X(_0971_));
 sg13g2_nand2b_1 _4233_ (.Y(_0972_),
    .B(_0970_),
    .A_N(_0971_));
 sg13g2_xor2_1 _4234_ (.B(_0971_),
    .A(_0970_),
    .X(_0973_));
 sg13g2_nand2_1 _4235_ (.Y(_0974_),
    .A(_0931_),
    .B(_0945_));
 sg13g2_or2_1 _4236_ (.X(_0975_),
    .B(_0973_),
    .A(_0945_));
 sg13g2_xor2_1 _4237_ (.B(_0974_),
    .A(_0973_),
    .X(_0976_));
 sg13g2_or2_1 _4238_ (.X(_0977_),
    .B(_0976_),
    .A(_0966_));
 sg13g2_xnor2_1 _4239_ (.Y(_0978_),
    .A(_0947_),
    .B(_0965_));
 sg13g2_xor2_1 _4240_ (.B(_0964_),
    .A(_0958_),
    .X(_0979_));
 sg13g2_nand2_1 _4241_ (.Y(_0980_),
    .A(\wirecube_top_inst.edge_function_inst.term0[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[6] ));
 sg13g2_nand2_1 _4242_ (.Y(_0981_),
    .A(\wirecube_top_inst.edge_function_inst.term1[4] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[2] ));
 sg13g2_xor2_1 _4243_ (.B(_0980_),
    .A(_0948_),
    .X(_0982_));
 sg13g2_nand2b_1 _4244_ (.Y(_0983_),
    .B(_0982_),
    .A_N(_0981_));
 sg13g2_o21ai_1 _4245_ (.B1(_0983_),
    .Y(_0984_),
    .A1(_0948_),
    .A2(_0980_));
 sg13g2_xnor2_1 _4246_ (.Y(_0985_),
    .A(_0950_),
    .B(_0951_));
 sg13g2_nand2_1 _4247_ (.Y(_0986_),
    .A(_0984_),
    .B(_0985_));
 sg13g2_nand2_1 _4248_ (.Y(_0987_),
    .A(\wirecube_top_inst.edge_function_inst.term0[6] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[1] ));
 sg13g2_nand2_1 _4249_ (.Y(_0988_),
    .A(\wirecube_top_inst.edge_function_inst.term0[4] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[2] ));
 sg13g2_nand2_1 _4250_ (.Y(_0989_),
    .A(\wirecube_top_inst.edge_function_inst.term0[4] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[3] ));
 sg13g2_xor2_1 _4251_ (.B(_0989_),
    .A(_0957_),
    .X(_0990_));
 sg13g2_nand2b_1 _4252_ (.Y(_0991_),
    .B(_0990_),
    .A_N(_0987_));
 sg13g2_xnor2_1 _4253_ (.Y(_0992_),
    .A(_0987_),
    .B(_0990_));
 sg13g2_inv_1 _4254_ (.Y(_0993_),
    .A(_0992_));
 sg13g2_xnor2_1 _4255_ (.Y(_0994_),
    .A(_0984_),
    .B(_0985_));
 sg13g2_o21ai_1 _4256_ (.B1(_0986_),
    .Y(_0995_),
    .A1(_0993_),
    .A2(_0994_));
 sg13g2_xor2_1 _4257_ (.B(_0960_),
    .A(_0959_),
    .X(_0996_));
 sg13g2_nand2_1 _4258_ (.Y(_0997_),
    .A(_0995_),
    .B(_0996_));
 sg13g2_o21ai_1 _4259_ (.B1(_0991_),
    .Y(_0998_),
    .A1(_0957_),
    .A2(_0989_));
 sg13g2_inv_1 _4260_ (.Y(_0999_),
    .A(_0998_));
 sg13g2_xnor2_1 _4261_ (.Y(_1000_),
    .A(_0995_),
    .B(_0996_));
 sg13g2_o21ai_1 _4262_ (.B1(_0997_),
    .Y(_1001_),
    .A1(_0999_),
    .A2(_1000_));
 sg13g2_nand2_1 _4263_ (.Y(_1002_),
    .A(_0979_),
    .B(_1001_));
 sg13g2_nor2_1 _4264_ (.A(_0978_),
    .B(_1002_),
    .Y(_1003_));
 sg13g2_xor2_1 _4265_ (.B(_1001_),
    .A(_0979_),
    .X(_1004_));
 sg13g2_xnor2_1 _4266_ (.Y(_1005_),
    .A(_0999_),
    .B(_1000_));
 sg13g2_nand2_2 _4267_ (.Y(_1006_),
    .A(\wirecube_top_inst.edge_function_inst.term0[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[4] ));
 sg13g2_nor2_1 _4268_ (.A(_0948_),
    .B(_1006_),
    .Y(_1007_));
 sg13g2_xnor2_1 _4269_ (.Y(_1008_),
    .A(_0981_),
    .B(_0982_));
 sg13g2_and2_1 _4270_ (.A(_1007_),
    .B(_1008_),
    .X(_1009_));
 sg13g2_xor2_1 _4271_ (.B(_1008_),
    .A(_1007_),
    .X(_1010_));
 sg13g2_nand2_1 _4272_ (.Y(_1011_),
    .A(\wirecube_top_inst.edge_function_inst.term0[5] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[1] ));
 sg13g2_nand2_1 _4273_ (.Y(_1012_),
    .A(\wirecube_top_inst.edge_function_inst.term0[3] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[2] ));
 sg13g2_nand2_1 _4274_ (.Y(_1013_),
    .A(\wirecube_top_inst.edge_function_inst.term0[3] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[3] ));
 sg13g2_xor2_1 _4275_ (.B(_1013_),
    .A(_0988_),
    .X(_1014_));
 sg13g2_nand2b_1 _4276_ (.Y(_1015_),
    .B(_1014_),
    .A_N(_1011_));
 sg13g2_xnor2_1 _4277_ (.Y(_1016_),
    .A(_1011_),
    .B(_1014_));
 sg13g2_a21o_1 _4278_ (.A2(_1016_),
    .A1(_1010_),
    .B1(_1009_),
    .X(_1017_));
 sg13g2_xnor2_1 _4279_ (.Y(_1018_),
    .A(_0993_),
    .B(_0994_));
 sg13g2_nand2b_1 _4280_ (.Y(_1019_),
    .B(_1017_),
    .A_N(_1018_));
 sg13g2_o21ai_1 _4281_ (.B1(_1015_),
    .Y(_1020_),
    .A1(_0988_),
    .A2(_1013_));
 sg13g2_inv_1 _4282_ (.Y(_1021_),
    .A(_1020_));
 sg13g2_xor2_1 _4283_ (.B(_1018_),
    .A(_1017_),
    .X(_1022_));
 sg13g2_o21ai_1 _4284_ (.B1(_1019_),
    .Y(_1023_),
    .A1(_1021_),
    .A2(_1022_));
 sg13g2_nand2b_1 _4285_ (.Y(_1024_),
    .B(_1023_),
    .A_N(_1005_));
 sg13g2_inv_1 _4286_ (.Y(_1025_),
    .A(_1024_));
 sg13g2_nand2_1 _4287_ (.Y(_1026_),
    .A(_1004_),
    .B(_1025_));
 sg13g2_xor2_1 _4288_ (.B(_1023_),
    .A(_1005_),
    .X(_1027_));
 sg13g2_xnor2_1 _4289_ (.Y(_1028_),
    .A(_1021_),
    .B(_1022_));
 sg13g2_nand2_1 _4290_ (.Y(_1029_),
    .A(\wirecube_top_inst.edge_function_inst.term0[4] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[1] ));
 sg13g2_nand2_2 _4291_ (.Y(_1030_),
    .A(\wirecube_top_inst.edge_function_inst.term0[2] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[2] ));
 sg13g2_nand2_1 _4292_ (.Y(_1031_),
    .A(\wirecube_top_inst.edge_function_inst.term0[2] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[3] ));
 sg13g2_or2_1 _4293_ (.X(_1032_),
    .B(_1030_),
    .A(_1013_));
 sg13g2_xor2_1 _4294_ (.B(_1031_),
    .A(_1012_),
    .X(_1033_));
 sg13g2_nand2b_1 _4295_ (.Y(_1034_),
    .B(_1033_),
    .A_N(_1029_));
 sg13g2_xnor2_1 _4296_ (.Y(_1035_),
    .A(_1029_),
    .B(_1033_));
 sg13g2_a22oi_1 _4297_ (.Y(_1036_),
    .B1(\wirecube_top_inst.edge_function_inst.term1[4] ),
    .B2(\wirecube_top_inst.edge_function_inst.term0[1] ),
    .A2(\wirecube_top_inst.edge_function_inst.term1[5] ),
    .A1(\wirecube_top_inst.edge_function_inst.term0[0] ));
 sg13g2_nor2_1 _4298_ (.A(_1007_),
    .B(_1036_),
    .Y(_1037_));
 sg13g2_nand2_1 _4299_ (.Y(_1038_),
    .A(_1035_),
    .B(_1037_));
 sg13g2_xnor2_1 _4300_ (.Y(_1039_),
    .A(_1010_),
    .B(_1016_));
 sg13g2_nor2_1 _4301_ (.A(_1038_),
    .B(_1039_),
    .Y(_1040_));
 sg13g2_and2_1 _4302_ (.A(_1032_),
    .B(_1034_),
    .X(_1041_));
 sg13g2_inv_1 _4303_ (.Y(_1042_),
    .A(_1041_));
 sg13g2_xor2_1 _4304_ (.B(_1039_),
    .A(_1038_),
    .X(_1043_));
 sg13g2_a21oi_1 _4305_ (.A1(_1042_),
    .A2(_1043_),
    .Y(_1044_),
    .B1(_1040_));
 sg13g2_nor2_1 _4306_ (.A(_1028_),
    .B(_1044_),
    .Y(_1045_));
 sg13g2_nor2b_1 _4307_ (.A(_1027_),
    .B_N(_1045_),
    .Y(_1046_));
 sg13g2_xnor2_1 _4308_ (.Y(_1047_),
    .A(_1028_),
    .B(_1044_));
 sg13g2_xor2_1 _4309_ (.B(_1037_),
    .A(_1035_),
    .X(_1048_));
 sg13g2_nand2_1 _4310_ (.Y(_1049_),
    .A(\wirecube_top_inst.edge_function_inst.term0[3] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[1] ));
 sg13g2_nand2_1 _4311_ (.Y(_1050_),
    .A(\wirecube_top_inst.edge_function_inst.term1[3] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[1] ));
 sg13g2_or2_1 _4312_ (.X(_1051_),
    .B(_1050_),
    .A(_1030_));
 sg13g2_and2_1 _4313_ (.A(_1030_),
    .B(_1050_),
    .X(_1052_));
 sg13g2_xor2_1 _4314_ (.B(_1050_),
    .A(_1030_),
    .X(_1053_));
 sg13g2_xnor2_1 _4315_ (.Y(_1054_),
    .A(_1049_),
    .B(_1053_));
 sg13g2_nand2b_1 _4316_ (.Y(_1055_),
    .B(_1054_),
    .A_N(_1006_));
 sg13g2_inv_1 _4317_ (.Y(_1056_),
    .A(_1055_));
 sg13g2_o21ai_1 _4318_ (.B1(_1051_),
    .Y(_1057_),
    .A1(_1049_),
    .A2(_1052_));
 sg13g2_xor2_1 _4319_ (.B(_1055_),
    .A(_1048_),
    .X(_1058_));
 sg13g2_nor2b_1 _4320_ (.A(_1058_),
    .B_N(_1057_),
    .Y(_1059_));
 sg13g2_a21oi_1 _4321_ (.A1(_1048_),
    .A2(_1056_),
    .Y(_1060_),
    .B1(_1059_));
 sg13g2_xnor2_1 _4322_ (.Y(_1061_),
    .A(_1041_),
    .B(_1043_));
 sg13g2_nor2b_1 _4323_ (.A(_1060_),
    .B_N(_1061_),
    .Y(_1062_));
 sg13g2_and2_1 _4324_ (.A(\wirecube_top_inst.edge_function_inst.term1[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[6] ),
    .X(_1063_));
 sg13g2_xnor2_1 _4325_ (.Y(_1064_),
    .A(_1060_),
    .B(_1061_));
 sg13g2_a21oi_1 _4326_ (.A1(_1063_),
    .A2(_1064_),
    .Y(_1065_),
    .B1(_1062_));
 sg13g2_or2_1 _4327_ (.X(_1066_),
    .B(_1065_),
    .A(_1047_));
 sg13g2_nand2_1 _4328_ (.Y(_1067_),
    .A(\wirecube_top_inst.edge_function_inst.term0[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[2] ));
 sg13g2_or2_1 _4329_ (.X(_1068_),
    .B(_1067_),
    .A(_1050_));
 sg13g2_nand2_1 _4330_ (.Y(_1069_),
    .A(\wirecube_top_inst.edge_function_inst.term0[2] ),
    .B(\wirecube_top_inst.edge_function_inst.term1[1] ));
 sg13g2_a22oi_1 _4331_ (.Y(_1070_),
    .B1(\wirecube_top_inst.edge_function_inst.term0[1] ),
    .B2(\wirecube_top_inst.edge_function_inst.term1[2] ),
    .A2(\wirecube_top_inst.edge_function_inst.term1[3] ),
    .A1(\wirecube_top_inst.edge_function_inst.term0[0] ));
 sg13g2_inv_1 _4332_ (.Y(_1071_),
    .A(_1070_));
 sg13g2_and2_1 _4333_ (.A(_1068_),
    .B(_1071_),
    .X(_1072_));
 sg13g2_o21ai_1 _4334_ (.B1(_1068_),
    .Y(_1073_),
    .A1(_1069_),
    .A2(_1070_));
 sg13g2_xor2_1 _4335_ (.B(_1054_),
    .A(_1006_),
    .X(_1074_));
 sg13g2_nor2b_1 _4336_ (.A(_1074_),
    .B_N(_1073_),
    .Y(_1075_));
 sg13g2_xnor2_1 _4337_ (.Y(_1076_),
    .A(_1057_),
    .B(_1058_));
 sg13g2_nand2_1 _4338_ (.Y(_1077_),
    .A(_1075_),
    .B(_1076_));
 sg13g2_nand2_1 _4339_ (.Y(_1078_),
    .A(\wirecube_top_inst.edge_function_inst.term1[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[5] ));
 sg13g2_xnor2_1 _4340_ (.Y(_1079_),
    .A(_1075_),
    .B(_1076_));
 sg13g2_o21ai_1 _4341_ (.B1(_1077_),
    .Y(_1080_),
    .A1(_1078_),
    .A2(_1079_));
 sg13g2_xor2_1 _4342_ (.B(_1064_),
    .A(_1063_),
    .X(_1081_));
 sg13g2_nand2_1 _4343_ (.Y(_1082_),
    .A(_1080_),
    .B(_1081_));
 sg13g2_xor2_1 _4344_ (.B(_1074_),
    .A(_1073_),
    .X(_1083_));
 sg13g2_nand4_1 _4345_ (.B(\wirecube_top_inst.edge_function_inst.term0[1] ),
    .C(\wirecube_top_inst.edge_function_inst.term1[2] ),
    .A(\wirecube_top_inst.edge_function_inst.term0[0] ),
    .Y(_1084_),
    .D(\wirecube_top_inst.edge_function_inst.term1[1] ));
 sg13g2_xnor2_1 _4346_ (.Y(_1085_),
    .A(_1069_),
    .B(_1072_));
 sg13g2_nand2b_1 _4347_ (.Y(_1086_),
    .B(_1085_),
    .A_N(_1084_));
 sg13g2_nand2_1 _4348_ (.Y(_1087_),
    .A(\wirecube_top_inst.edge_function_inst.term1[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[4] ));
 sg13g2_xor2_1 _4349_ (.B(_1086_),
    .A(_1083_),
    .X(_1088_));
 sg13g2_nand2b_1 _4350_ (.Y(_1089_),
    .B(_1088_),
    .A_N(_1087_));
 sg13g2_o21ai_1 _4351_ (.B1(_1089_),
    .Y(_1090_),
    .A1(_1083_),
    .A2(_1086_));
 sg13g2_xor2_1 _4352_ (.B(_1079_),
    .A(_1078_),
    .X(_1091_));
 sg13g2_and2_1 _4353_ (.A(_1090_),
    .B(_1091_),
    .X(_1092_));
 sg13g2_nand2_1 _4354_ (.Y(_1093_),
    .A(\wirecube_top_inst.edge_function_inst.term1[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[3] ));
 sg13g2_xnor2_1 _4355_ (.Y(_1094_),
    .A(_1084_),
    .B(_1085_));
 sg13g2_nor2b_1 _4356_ (.A(_1093_),
    .B_N(_1094_),
    .Y(_1095_));
 sg13g2_xnor2_1 _4357_ (.Y(_1096_),
    .A(_1087_),
    .B(_1088_));
 sg13g2_xnor2_1 _4358_ (.Y(_1097_),
    .A(_1093_),
    .B(_1094_));
 sg13g2_nand2_1 _4359_ (.Y(_1098_),
    .A(_0907_),
    .B(_1067_));
 sg13g2_and4_1 _4360_ (.A(\wirecube_top_inst.edge_function_inst.term1[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term0[2] ),
    .C(_1084_),
    .D(_1098_),
    .X(_1099_));
 sg13g2_nand2_1 _4361_ (.Y(_1100_),
    .A(_1097_),
    .B(_1099_));
 sg13g2_a22oi_1 _4362_ (.Y(_1101_),
    .B1(_1084_),
    .B2(_1098_),
    .A2(\wirecube_top_inst.edge_function_inst.term0[2] ),
    .A1(\wirecube_top_inst.edge_function_inst.term1[0] ));
 sg13g2_nor2_1 _4363_ (.A(_1099_),
    .B(_1101_),
    .Y(_1102_));
 sg13g2_nand2_1 _4364_ (.Y(_1103_),
    .A(_0908_),
    .B(_1102_));
 sg13g2_xnor2_1 _4365_ (.Y(_1104_),
    .A(_1097_),
    .B(_1099_));
 sg13g2_o21ai_1 _4366_ (.B1(_1100_),
    .Y(_1105_),
    .A1(_1103_),
    .A2(_1104_));
 sg13g2_xnor2_1 _4367_ (.Y(_1106_),
    .A(_1095_),
    .B(_1096_));
 sg13g2_nor2b_1 _4368_ (.A(_1106_),
    .B_N(_1105_),
    .Y(_1107_));
 sg13g2_a21oi_1 _4369_ (.A1(_1095_),
    .A2(_1096_),
    .Y(_1108_),
    .B1(_1107_));
 sg13g2_xnor2_1 _4370_ (.Y(_1109_),
    .A(_1090_),
    .B(_1091_));
 sg13g2_nor2_1 _4371_ (.A(_1108_),
    .B(_1109_),
    .Y(_1110_));
 sg13g2_xnor2_1 _4372_ (.Y(_1111_),
    .A(_1080_),
    .B(_1081_));
 sg13g2_inv_1 _4373_ (.Y(_1112_),
    .A(_1111_));
 sg13g2_o21ai_1 _4374_ (.B1(_1112_),
    .Y(_1113_),
    .A1(_1092_),
    .A2(_1110_));
 sg13g2_xnor2_1 _4375_ (.Y(_1114_),
    .A(_1047_),
    .B(_1065_));
 sg13g2_a21o_1 _4376_ (.A2(_1113_),
    .A1(_1082_),
    .B1(_1114_),
    .X(_1115_));
 sg13g2_xor2_1 _4377_ (.B(_1045_),
    .A(_1027_),
    .X(_1116_));
 sg13g2_a21oi_1 _4378_ (.A1(_1066_),
    .A2(_1115_),
    .Y(_1117_),
    .B1(_1116_));
 sg13g2_xnor2_1 _4379_ (.Y(_1118_),
    .A(_1004_),
    .B(_1024_));
 sg13g2_o21ai_1 _4380_ (.B1(_1118_),
    .Y(_1119_),
    .A1(_1046_),
    .A2(_1117_));
 sg13g2_xnor2_1 _4381_ (.Y(_1120_),
    .A(_0978_),
    .B(_1002_));
 sg13g2_a21oi_1 _4382_ (.A1(_1026_),
    .A2(_1119_),
    .Y(_1121_),
    .B1(_1120_));
 sg13g2_xor2_1 _4383_ (.B(_0976_),
    .A(_0966_),
    .X(_1122_));
 sg13g2_o21ai_1 _4384_ (.B1(_1122_),
    .Y(_1123_),
    .A1(_1003_),
    .A2(_1121_));
 sg13g2_nand2b_1 _4385_ (.Y(_1124_),
    .B(_0918_),
    .A_N(_0967_));
 sg13g2_o21ai_1 _4386_ (.B1(_0972_),
    .Y(_1125_),
    .A1(_0931_),
    .A2(_0973_));
 sg13g2_inv_1 _4387_ (.Y(_1126_),
    .A(_1125_));
 sg13g2_xnor2_1 _4388_ (.Y(_1127_),
    .A(_1124_),
    .B(_1125_));
 sg13g2_nor2b_1 _4389_ (.A(_0975_),
    .B_N(_1127_),
    .Y(_1128_));
 sg13g2_xor2_1 _4390_ (.B(_1127_),
    .A(_0975_),
    .X(_1129_));
 sg13g2_a21oi_1 _4391_ (.A1(_0977_),
    .A2(_1123_),
    .Y(_1130_),
    .B1(_1129_));
 sg13g2_a21oi_1 _4392_ (.A1(_0918_),
    .A2(_1126_),
    .Y(_1131_),
    .B1(_0967_));
 sg13g2_nor3_2 _4393_ (.A(_1128_),
    .B(_1130_),
    .C(_1131_),
    .Y(_1132_));
 sg13g2_nand2_1 _4394_ (.Y(_1133_),
    .A(\wirecube_top_inst.edge_function_inst.term2[5] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[4] ));
 sg13g2_nand2_1 _4395_ (.Y(_1134_),
    .A(\wirecube_top_inst.edge_function_inst.term3[6] ),
    .B(\wirecube_top_inst.edge_function_inst.term2[4] ));
 sg13g2_nand2_1 _4396_ (.Y(_1135_),
    .A(\wirecube_top_inst.edge_function_inst.term3[5] ),
    .B(net706));
 sg13g2_nand2_1 _4397_ (.Y(_1136_),
    .A(\wirecube_top_inst.edge_function_inst.term3[5] ),
    .B(\wirecube_top_inst.edge_function_inst.term2[4] ));
 sg13g2_nand2_1 _4398_ (.Y(_1137_),
    .A(\wirecube_top_inst.edge_function_inst.term3[6] ),
    .B(net706));
 sg13g2_or2_1 _4399_ (.X(_1138_),
    .B(_1135_),
    .A(_1134_));
 sg13g2_xor2_1 _4400_ (.B(_1137_),
    .A(_1136_),
    .X(_1139_));
 sg13g2_nand2b_1 _4401_ (.Y(_1140_),
    .B(_1139_),
    .A_N(_1133_));
 sg13g2_xnor2_1 _4402_ (.Y(_1141_),
    .A(_1133_),
    .B(_1139_));
 sg13g2_nand2_2 _4403_ (.Y(_1142_),
    .A(\wirecube_top_inst.edge_function_inst.term3[6] ),
    .B(\wirecube_top_inst.edge_function_inst.term2[2] ));
 sg13g2_nand2_1 _4404_ (.Y(_1143_),
    .A(\wirecube_top_inst.edge_function_inst.term2[4] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[4] ));
 sg13g2_xor2_1 _4405_ (.B(_1142_),
    .A(_1135_),
    .X(_1144_));
 sg13g2_nand2b_1 _4406_ (.Y(_1145_),
    .B(_1144_),
    .A_N(_1143_));
 sg13g2_o21ai_1 _4407_ (.B1(_1145_),
    .Y(_1146_),
    .A1(_1135_),
    .A2(_1142_));
 sg13g2_nand2_1 _4408_ (.Y(_1147_),
    .A(_1141_),
    .B(_1146_));
 sg13g2_xor2_1 _4409_ (.B(_1146_),
    .A(_1141_),
    .X(_1148_));
 sg13g2_nand2_2 _4410_ (.Y(_1149_),
    .A(\wirecube_top_inst.edge_function_inst.term3[5] ),
    .B(\wirecube_top_inst.edge_function_inst.term2[1] ));
 sg13g2_nor2_1 _4411_ (.A(_1142_),
    .B(_1149_),
    .Y(_1150_));
 sg13g2_or2_1 _4412_ (.X(_1151_),
    .B(_1149_),
    .A(_1142_));
 sg13g2_nand2_1 _4413_ (.Y(_1152_),
    .A(\wirecube_top_inst.edge_function_inst.term3[4] ),
    .B(net706));
 sg13g2_a22oi_1 _4414_ (.Y(_1153_),
    .B1(\wirecube_top_inst.edge_function_inst.term2[1] ),
    .B2(\wirecube_top_inst.edge_function_inst.term3[6] ),
    .A2(\wirecube_top_inst.edge_function_inst.term2[2] ),
    .A1(\wirecube_top_inst.edge_function_inst.term3[5] ));
 sg13g2_or2_1 _4415_ (.X(_1154_),
    .B(_1153_),
    .A(_1150_));
 sg13g2_o21ai_1 _4416_ (.B1(_1151_),
    .Y(_1155_),
    .A1(_1152_),
    .A2(_1154_));
 sg13g2_xnor2_1 _4417_ (.Y(_1156_),
    .A(_1143_),
    .B(_1144_));
 sg13g2_nand2_1 _4418_ (.Y(_1157_),
    .A(_1155_),
    .B(_1156_));
 sg13g2_nand2_2 _4419_ (.Y(_1158_),
    .A(\wirecube_top_inst.edge_function_inst.term2[6] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[2] ));
 sg13g2_xnor2_1 _4420_ (.Y(_1159_),
    .A(_1155_),
    .B(_1156_));
 sg13g2_o21ai_1 _4421_ (.B1(_1157_),
    .Y(_1160_),
    .A1(_1158_),
    .A2(_1159_));
 sg13g2_nand2_1 _4422_ (.Y(_1161_),
    .A(_1148_),
    .B(_1160_));
 sg13g2_xor2_1 _4423_ (.B(_1160_),
    .A(_1148_),
    .X(_1162_));
 sg13g2_nand2_1 _4424_ (.Y(_1163_),
    .A(\wirecube_top_inst.edge_function_inst.term2[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[6] ));
 sg13g2_nand2_1 _4425_ (.Y(_1164_),
    .A(\wirecube_top_inst.edge_function_inst.term3[4] ),
    .B(\wirecube_top_inst.edge_function_inst.term2[2] ));
 sg13g2_xor2_1 _4426_ (.B(_1163_),
    .A(_1149_),
    .X(_1165_));
 sg13g2_nand2b_1 _4427_ (.Y(_1166_),
    .B(_1165_),
    .A_N(_1164_));
 sg13g2_o21ai_1 _4428_ (.B1(_1166_),
    .Y(_1167_),
    .A1(_1149_),
    .A2(_1163_));
 sg13g2_xor2_1 _4429_ (.B(_1154_),
    .A(_1152_),
    .X(_1168_));
 sg13g2_nand2_1 _4430_ (.Y(_1169_),
    .A(_1167_),
    .B(_1168_));
 sg13g2_a22oi_1 _4431_ (.Y(_1170_),
    .B1(\wirecube_top_inst.edge_function_inst.term3[1] ),
    .B2(\wirecube_top_inst.edge_function_inst.term2[6] ),
    .A2(\wirecube_top_inst.edge_function_inst.term3[2] ),
    .A1(\wirecube_top_inst.edge_function_inst.term2[5] ));
 sg13g2_nand2_1 _4432_ (.Y(_1171_),
    .A(\wirecube_top_inst.edge_function_inst.term2[5] ),
    .B(net705));
 sg13g2_or2_1 _4433_ (.X(_1172_),
    .B(_1171_),
    .A(_1158_));
 sg13g2_nand2b_1 _4434_ (.Y(_1173_),
    .B(_1172_),
    .A_N(_1170_));
 sg13g2_xnor2_1 _4435_ (.Y(_1174_),
    .A(_1167_),
    .B(_1168_));
 sg13g2_o21ai_1 _4436_ (.B1(_1169_),
    .Y(_1175_),
    .A1(_1173_),
    .A2(_1174_));
 sg13g2_xor2_1 _4437_ (.B(_1159_),
    .A(_1158_),
    .X(_1176_));
 sg13g2_nand2_1 _4438_ (.Y(_1177_),
    .A(_1175_),
    .B(_1176_));
 sg13g2_xnor2_1 _4439_ (.Y(_1178_),
    .A(_1175_),
    .B(_1176_));
 sg13g2_o21ai_1 _4440_ (.B1(_1177_),
    .Y(_1179_),
    .A1(_1172_),
    .A2(_1178_));
 sg13g2_nand2_1 _4441_ (.Y(_1180_),
    .A(_1162_),
    .B(_1179_));
 sg13g2_nand2_1 _4442_ (.Y(_1181_),
    .A(\wirecube_top_inst.edge_function_inst.term2[6] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[3] ));
 sg13g2_nor2_1 _4443_ (.A(_1162_),
    .B(_1179_),
    .Y(_1182_));
 sg13g2_xor2_1 _4444_ (.B(_1179_),
    .A(_1162_),
    .X(_1183_));
 sg13g2_o21ai_1 _4445_ (.B1(_1180_),
    .Y(_1184_),
    .A1(_1181_),
    .A2(_1182_));
 sg13g2_nand2_1 _4446_ (.Y(_1185_),
    .A(\wirecube_top_inst.edge_function_inst.term2[6] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[4] ));
 sg13g2_nand2_2 _4447_ (.Y(_1186_),
    .A(\wirecube_top_inst.edge_function_inst.term2[5] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[5] ));
 sg13g2_xor2_1 _4448_ (.B(_1186_),
    .A(_1134_),
    .X(_1187_));
 sg13g2_nand2b_1 _4449_ (.Y(_1188_),
    .B(_1187_),
    .A_N(_1185_));
 sg13g2_xnor2_1 _4450_ (.Y(_1189_),
    .A(_1185_),
    .B(_1187_));
 sg13g2_and2_1 _4451_ (.A(_1138_),
    .B(_1140_),
    .X(_1190_));
 sg13g2_nand2b_1 _4452_ (.Y(_1191_),
    .B(_1189_),
    .A_N(_1190_));
 sg13g2_xnor2_1 _4453_ (.Y(_1192_),
    .A(_1189_),
    .B(_1190_));
 sg13g2_nand2_1 _4454_ (.Y(_1193_),
    .A(_1147_),
    .B(_1161_));
 sg13g2_nand2b_1 _4455_ (.Y(_1194_),
    .B(_1192_),
    .A_N(_1147_));
 sg13g2_nand3_1 _4456_ (.B(_1160_),
    .C(_1192_),
    .A(_1148_),
    .Y(_1195_));
 sg13g2_xor2_1 _4457_ (.B(_1193_),
    .A(_1192_),
    .X(_1196_));
 sg13g2_and2_1 _4458_ (.A(_1184_),
    .B(_1196_),
    .X(_1197_));
 sg13g2_nand2_1 _4459_ (.Y(_1198_),
    .A(\wirecube_top_inst.edge_function_inst.term2[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[4] ));
 sg13g2_nor2_1 _4460_ (.A(_1149_),
    .B(_1198_),
    .Y(_1199_));
 sg13g2_xnor2_1 _4461_ (.Y(_1200_),
    .A(_1164_),
    .B(_1165_));
 sg13g2_and2_1 _4462_ (.A(_1199_),
    .B(_1200_),
    .X(_1201_));
 sg13g2_xor2_1 _4463_ (.B(_1200_),
    .A(_1199_),
    .X(_1202_));
 sg13g2_nand2_1 _4464_ (.Y(_1203_),
    .A(\wirecube_top_inst.edge_function_inst.term2[4] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[2] ));
 sg13g2_nand2_1 _4465_ (.Y(_1204_),
    .A(\wirecube_top_inst.edge_function_inst.term3[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term2[5] ));
 sg13g2_nand2_1 _4466_ (.Y(_1205_),
    .A(\wirecube_top_inst.edge_function_inst.term3[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term2[6] ));
 sg13g2_xor2_1 _4467_ (.B(_1205_),
    .A(_1171_),
    .X(_1206_));
 sg13g2_nand2b_1 _4468_ (.Y(_1207_),
    .B(_1206_),
    .A_N(_1203_));
 sg13g2_xnor2_1 _4469_ (.Y(_1208_),
    .A(_1203_),
    .B(_1206_));
 sg13g2_a21o_1 _4470_ (.A2(_1208_),
    .A1(_1202_),
    .B1(_1201_),
    .X(_1209_));
 sg13g2_xor2_1 _4471_ (.B(_1174_),
    .A(_1173_),
    .X(_1210_));
 sg13g2_nand2_1 _4472_ (.Y(_1211_),
    .A(_1209_),
    .B(_1210_));
 sg13g2_o21ai_1 _4473_ (.B1(_1207_),
    .Y(_1212_),
    .A1(_1171_),
    .A2(_1205_));
 sg13g2_inv_1 _4474_ (.Y(_1213_),
    .A(_1212_));
 sg13g2_xnor2_1 _4475_ (.Y(_1214_),
    .A(_1209_),
    .B(_1210_));
 sg13g2_o21ai_1 _4476_ (.B1(_1211_),
    .Y(_1215_),
    .A1(_1213_),
    .A2(_1214_));
 sg13g2_xor2_1 _4477_ (.B(_1178_),
    .A(_1172_),
    .X(_1216_));
 sg13g2_nand2_1 _4478_ (.Y(_1217_),
    .A(_1215_),
    .B(_1216_));
 sg13g2_nand2_1 _4479_ (.Y(_1218_),
    .A(\wirecube_top_inst.edge_function_inst.term2[5] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[3] ));
 sg13g2_xnor2_1 _4480_ (.Y(_1219_),
    .A(_1215_),
    .B(_1216_));
 sg13g2_o21ai_1 _4481_ (.B1(_1217_),
    .Y(_1220_),
    .A1(_1218_),
    .A2(_1219_));
 sg13g2_xnor2_1 _4482_ (.Y(_1221_),
    .A(_1181_),
    .B(_1183_));
 sg13g2_nand2_1 _4483_ (.Y(_1222_),
    .A(net706),
    .B(\wirecube_top_inst.edge_function_inst.term3[2] ));
 sg13g2_nand2_1 _4484_ (.Y(_1223_),
    .A(\wirecube_top_inst.edge_function_inst.term2[4] ),
    .B(net705));
 sg13g2_or2_1 _4485_ (.X(_1224_),
    .B(_1223_),
    .A(_1204_));
 sg13g2_xor2_1 _4486_ (.B(_1223_),
    .A(_1204_),
    .X(_1225_));
 sg13g2_nand2b_1 _4487_ (.Y(_1226_),
    .B(_1225_),
    .A_N(_1222_));
 sg13g2_xnor2_1 _4488_ (.Y(_1227_),
    .A(_1222_),
    .B(_1225_));
 sg13g2_a22oi_1 _4489_ (.Y(_1228_),
    .B1(\wirecube_top_inst.edge_function_inst.term3[4] ),
    .B2(\wirecube_top_inst.edge_function_inst.term2[1] ),
    .A2(\wirecube_top_inst.edge_function_inst.term3[5] ),
    .A1(\wirecube_top_inst.edge_function_inst.term2[0] ));
 sg13g2_nor2_1 _4490_ (.A(_1199_),
    .B(_1228_),
    .Y(_1229_));
 sg13g2_nand2_1 _4491_ (.Y(_1230_),
    .A(_1227_),
    .B(_1229_));
 sg13g2_xnor2_1 _4492_ (.Y(_1231_),
    .A(_1202_),
    .B(_1208_));
 sg13g2_nor2_1 _4493_ (.A(_1230_),
    .B(_1231_),
    .Y(_1232_));
 sg13g2_and2_1 _4494_ (.A(_1224_),
    .B(_1226_),
    .X(_1233_));
 sg13g2_inv_1 _4495_ (.Y(_1234_),
    .A(_1233_));
 sg13g2_xor2_1 _4496_ (.B(_1231_),
    .A(_1230_),
    .X(_1235_));
 sg13g2_a21oi_1 _4497_ (.A1(_1234_),
    .A2(_1235_),
    .Y(_1236_),
    .B1(_1232_));
 sg13g2_xnor2_1 _4498_ (.Y(_1237_),
    .A(_1213_),
    .B(_1214_));
 sg13g2_nand2_1 _4499_ (.Y(_1238_),
    .A(\wirecube_top_inst.edge_function_inst.term2[4] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[3] ));
 sg13g2_xor2_1 _4500_ (.B(_1237_),
    .A(_1236_),
    .X(_1239_));
 sg13g2_nand2b_1 _4501_ (.Y(_1240_),
    .B(_1239_),
    .A_N(_1238_));
 sg13g2_o21ai_1 _4502_ (.B1(_1240_),
    .Y(_1241_),
    .A1(_1236_),
    .A2(_1237_));
 sg13g2_xor2_1 _4503_ (.B(_1219_),
    .A(_1218_),
    .X(_1242_));
 sg13g2_nand2_1 _4504_ (.Y(_1243_),
    .A(_1241_),
    .B(_1242_));
 sg13g2_xor2_1 _4505_ (.B(_1229_),
    .A(_1227_),
    .X(_1244_));
 sg13g2_and2_1 _4506_ (.A(\wirecube_top_inst.edge_function_inst.term2[2] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[2] ),
    .X(_1245_));
 sg13g2_nand2_1 _4507_ (.Y(_1246_),
    .A(\wirecube_top_inst.edge_function_inst.term2[3] ),
    .B(net705));
 sg13g2_nand4_1 _4508_ (.B(\wirecube_top_inst.edge_function_inst.term2[4] ),
    .C(\wirecube_top_inst.edge_function_inst.term2[3] ),
    .A(\wirecube_top_inst.edge_function_inst.term3[0] ),
    .Y(_1247_),
    .D(net705));
 sg13g2_inv_1 _4509_ (.Y(_1248_),
    .A(_1247_));
 sg13g2_a22oi_1 _4510_ (.Y(_1249_),
    .B1(net706),
    .B2(net705),
    .A2(\wirecube_top_inst.edge_function_inst.term2[4] ),
    .A1(\wirecube_top_inst.edge_function_inst.term3[0] ));
 sg13g2_nor2_1 _4511_ (.A(_1248_),
    .B(_1249_),
    .Y(_1250_));
 sg13g2_xor2_1 _4512_ (.B(_1250_),
    .A(_1245_),
    .X(_1251_));
 sg13g2_nand2b_1 _4513_ (.Y(_1252_),
    .B(_1251_),
    .A_N(_1198_));
 sg13g2_inv_1 _4514_ (.Y(_1253_),
    .A(_1252_));
 sg13g2_a21oi_1 _4515_ (.A1(_1245_),
    .A2(_1250_),
    .Y(_1254_),
    .B1(_1248_));
 sg13g2_xor2_1 _4516_ (.B(_1252_),
    .A(_1244_),
    .X(_1255_));
 sg13g2_nor2_1 _4517_ (.A(_1254_),
    .B(_1255_),
    .Y(_1256_));
 sg13g2_a21oi_1 _4518_ (.A1(_1244_),
    .A2(_1253_),
    .Y(_1257_),
    .B1(_1256_));
 sg13g2_xnor2_1 _4519_ (.Y(_1258_),
    .A(_1233_),
    .B(_1235_));
 sg13g2_nor2b_1 _4520_ (.A(_1257_),
    .B_N(_1258_),
    .Y(_1259_));
 sg13g2_and2_1 _4521_ (.A(net706),
    .B(\wirecube_top_inst.edge_function_inst.term3[3] ),
    .X(_1260_));
 sg13g2_nand2_1 _4522_ (.Y(_1261_),
    .A(net706),
    .B(\wirecube_top_inst.edge_function_inst.term3[3] ));
 sg13g2_xnor2_1 _4523_ (.Y(_1262_),
    .A(_1257_),
    .B(_1258_));
 sg13g2_a21oi_1 _4524_ (.A1(_1260_),
    .A2(_1262_),
    .Y(_1263_),
    .B1(_1259_));
 sg13g2_xnor2_1 _4525_ (.Y(_1264_),
    .A(_1238_),
    .B(_1239_));
 sg13g2_nor2b_1 _4526_ (.A(_1263_),
    .B_N(_1264_),
    .Y(_1265_));
 sg13g2_nand2_1 _4527_ (.Y(_1266_),
    .A(\wirecube_top_inst.edge_function_inst.term3[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term2[2] ));
 sg13g2_nor2_1 _4528_ (.A(_1246_),
    .B(_1266_),
    .Y(_1267_));
 sg13g2_or2_1 _4529_ (.X(_1268_),
    .B(_1266_),
    .A(_1246_));
 sg13g2_nand2_1 _4530_ (.Y(_1269_),
    .A(\wirecube_top_inst.edge_function_inst.term2[1] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[2] ));
 sg13g2_a22oi_1 _4531_ (.Y(_1270_),
    .B1(\wirecube_top_inst.edge_function_inst.term2[2] ),
    .B2(net705),
    .A2(net706),
    .A1(\wirecube_top_inst.edge_function_inst.term3[0] ));
 sg13g2_nor2_1 _4532_ (.A(_1267_),
    .B(_1270_),
    .Y(_1271_));
 sg13g2_o21ai_1 _4533_ (.B1(_1268_),
    .Y(_1272_),
    .A1(_1269_),
    .A2(_1270_));
 sg13g2_xnor2_1 _4534_ (.Y(_1273_),
    .A(_1198_),
    .B(_1251_));
 sg13g2_and2_1 _4535_ (.A(_1272_),
    .B(_1273_),
    .X(_1274_));
 sg13g2_xor2_1 _4536_ (.B(_1255_),
    .A(_1254_),
    .X(_1275_));
 sg13g2_nand2_1 _4537_ (.Y(_1276_),
    .A(_1274_),
    .B(_1275_));
 sg13g2_nand2_1 _4538_ (.Y(_1277_),
    .A(\wirecube_top_inst.edge_function_inst.term2[2] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[3] ));
 sg13g2_xnor2_1 _4539_ (.Y(_1278_),
    .A(_1274_),
    .B(_1275_));
 sg13g2_o21ai_1 _4540_ (.B1(_1276_),
    .Y(_1279_),
    .A1(_1277_),
    .A2(_1278_));
 sg13g2_xnor2_1 _4541_ (.Y(_1280_),
    .A(_1261_),
    .B(_1262_));
 sg13g2_xnor2_1 _4542_ (.Y(_1281_),
    .A(_1272_),
    .B(_1273_));
 sg13g2_or2_1 _4543_ (.X(_1282_),
    .B(_1266_),
    .A(_0903_));
 sg13g2_nand2_1 _4544_ (.Y(_1283_),
    .A(\wirecube_top_inst.edge_function_inst.term2[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[2] ));
 sg13g2_xor2_1 _4545_ (.B(_1266_),
    .A(_0903_),
    .X(_1284_));
 sg13g2_nand2b_1 _4546_ (.Y(_1285_),
    .B(_1284_),
    .A_N(_1283_));
 sg13g2_and2_1 _4547_ (.A(_1282_),
    .B(_1285_),
    .X(_1286_));
 sg13g2_xnor2_1 _4548_ (.Y(_1287_),
    .A(_1269_),
    .B(_1271_));
 sg13g2_nand2b_1 _4549_ (.Y(_1288_),
    .B(_1287_),
    .A_N(_1286_));
 sg13g2_nand2_1 _4550_ (.Y(_1289_),
    .A(\wirecube_top_inst.edge_function_inst.term2[1] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[3] ));
 sg13g2_xor2_1 _4551_ (.B(_1288_),
    .A(_1281_),
    .X(_1290_));
 sg13g2_nand2b_1 _4552_ (.Y(_1291_),
    .B(_1290_),
    .A_N(_1289_));
 sg13g2_o21ai_1 _4553_ (.B1(_1291_),
    .Y(_1292_),
    .A1(_1281_),
    .A2(_1288_));
 sg13g2_xor2_1 _4554_ (.B(_1278_),
    .A(_1277_),
    .X(_1293_));
 sg13g2_nand2_1 _4555_ (.Y(_1294_),
    .A(_1292_),
    .B(_1293_));
 sg13g2_xor2_1 _4556_ (.B(_1290_),
    .A(_1289_),
    .X(_1295_));
 sg13g2_xnor2_1 _4557_ (.Y(_1296_),
    .A(_1286_),
    .B(_1287_));
 sg13g2_xnor2_1 _4558_ (.Y(_1297_),
    .A(_1283_),
    .B(_1284_));
 sg13g2_nand2_1 _4559_ (.Y(_1298_),
    .A(_0904_),
    .B(_1297_));
 sg13g2_inv_1 _4560_ (.Y(_1299_),
    .A(_1298_));
 sg13g2_nand2_1 _4561_ (.Y(_1300_),
    .A(_1296_),
    .B(_1299_));
 sg13g2_nand2_1 _4562_ (.Y(_1301_),
    .A(\wirecube_top_inst.edge_function_inst.term2[0] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[3] ));
 sg13g2_xnor2_1 _4563_ (.Y(_1302_),
    .A(_1296_),
    .B(_1299_));
 sg13g2_or2_1 _4564_ (.X(_1303_),
    .B(_1302_),
    .A(_1301_));
 sg13g2_a21o_2 _4565_ (.A2(_1303_),
    .A1(_1300_),
    .B1(_1295_),
    .X(_1304_));
 sg13g2_xnor2_1 _4566_ (.Y(_1305_),
    .A(_1292_),
    .B(_1293_));
 sg13g2_o21ai_1 _4567_ (.B1(_1294_),
    .Y(_1306_),
    .A1(_1304_),
    .A2(_1305_));
 sg13g2_xnor2_1 _4568_ (.Y(_1307_),
    .A(_1279_),
    .B(_1280_));
 sg13g2_nor2b_1 _4569_ (.A(_1307_),
    .B_N(_1306_),
    .Y(_1308_));
 sg13g2_a21oi_1 _4570_ (.A1(_1279_),
    .A2(_1280_),
    .Y(_1309_),
    .B1(_1308_));
 sg13g2_xnor2_1 _4571_ (.Y(_1310_),
    .A(_1263_),
    .B(_1264_));
 sg13g2_nor2b_1 _4572_ (.A(_1309_),
    .B_N(_1310_),
    .Y(_1311_));
 sg13g2_nor2_1 _4573_ (.A(_1265_),
    .B(_1311_),
    .Y(_1312_));
 sg13g2_xnor2_1 _4574_ (.Y(_1313_),
    .A(_1241_),
    .B(_1242_));
 sg13g2_o21ai_1 _4575_ (.B1(_1243_),
    .Y(_1314_),
    .A1(_1312_),
    .A2(_1313_));
 sg13g2_xnor2_1 _4576_ (.Y(_1315_),
    .A(_1220_),
    .B(_1221_));
 sg13g2_nor2b_1 _4577_ (.A(_1315_),
    .B_N(_1314_),
    .Y(_1316_));
 sg13g2_a21o_1 _4578_ (.A2(_1221_),
    .A1(_1220_),
    .B1(_1316_),
    .X(_1317_));
 sg13g2_xor2_1 _4579_ (.B(_1196_),
    .A(_1184_),
    .X(_1318_));
 sg13g2_a21o_1 _4580_ (.A2(_1318_),
    .A1(_1317_),
    .B1(_1197_),
    .X(_1319_));
 sg13g2_nand2_1 _4581_ (.Y(_1320_),
    .A(\wirecube_top_inst.edge_function_inst.term2[6] ),
    .B(\wirecube_top_inst.edge_function_inst.term3[6] ));
 sg13g2_nor2_1 _4582_ (.A(_1186_),
    .B(_1320_),
    .Y(_1321_));
 sg13g2_a22oi_1 _4583_ (.Y(_1322_),
    .B1(\wirecube_top_inst.edge_function_inst.term3[5] ),
    .B2(\wirecube_top_inst.edge_function_inst.term2[6] ),
    .A2(\wirecube_top_inst.edge_function_inst.term2[5] ),
    .A1(\wirecube_top_inst.edge_function_inst.term3[6] ));
 sg13g2_nor2_1 _4584_ (.A(_1321_),
    .B(_1322_),
    .Y(_1323_));
 sg13g2_o21ai_1 _4585_ (.B1(_1188_),
    .Y(_1324_),
    .A1(_1134_),
    .A2(_1186_));
 sg13g2_nand2_1 _4586_ (.Y(_1325_),
    .A(_1323_),
    .B(_1324_));
 sg13g2_xnor2_1 _4587_ (.Y(_1326_),
    .A(_1323_),
    .B(_1324_));
 sg13g2_nand3_1 _4588_ (.B(_1194_),
    .C(_1195_),
    .A(_1191_),
    .Y(_1327_));
 sg13g2_xnor2_1 _4589_ (.Y(_1328_),
    .A(_1326_),
    .B(_1327_));
 sg13g2_nand2_1 _4590_ (.Y(_1329_),
    .A(_1319_),
    .B(_1328_));
 sg13g2_o21ai_1 _4591_ (.B1(_1329_),
    .Y(_1330_),
    .A1(_1195_),
    .A2(_1326_));
 sg13g2_nor2b_1 _4592_ (.A(_1320_),
    .B_N(_1186_),
    .Y(_1331_));
 sg13g2_o21ai_1 _4593_ (.B1(_1325_),
    .Y(_1332_),
    .A1(_1191_),
    .A2(_1326_));
 sg13g2_inv_1 _4594_ (.Y(_1333_),
    .A(_1332_));
 sg13g2_xnor2_1 _4595_ (.Y(_1334_),
    .A(_1331_),
    .B(_1332_));
 sg13g2_nor3_1 _4596_ (.A(_1194_),
    .B(_1326_),
    .C(_1334_),
    .Y(_1335_));
 sg13g2_o21ai_1 _4597_ (.B1(_1334_),
    .Y(_1336_),
    .A1(_1194_),
    .A2(_1326_));
 sg13g2_nand2b_1 _4598_ (.Y(_1337_),
    .B(_1336_),
    .A_N(_1335_));
 sg13g2_nor2b_1 _4599_ (.A(_1337_),
    .B_N(_1330_),
    .Y(_1338_));
 sg13g2_a21oi_1 _4600_ (.A1(_1186_),
    .A2(_1333_),
    .Y(_1339_),
    .B1(_1320_));
 sg13g2_nor3_2 _4601_ (.A(_1335_),
    .B(_1338_),
    .C(_1339_),
    .Y(_1340_));
 sg13g2_nor2b_1 _4602_ (.A(_1340_),
    .B_N(_1132_),
    .Y(_1341_));
 sg13g2_nand2b_1 _4603_ (.Y(_1342_),
    .B(_1340_),
    .A_N(_1132_));
 sg13g2_xor2_1 _4604_ (.B(_1337_),
    .A(_1330_),
    .X(_1343_));
 sg13g2_nand3_1 _4605_ (.B(_1123_),
    .C(_1129_),
    .A(_0977_),
    .Y(_1344_));
 sg13g2_nor2b_1 _4606_ (.A(_1130_),
    .B_N(_1344_),
    .Y(_1345_));
 sg13g2_nor2_1 _4607_ (.A(_1343_),
    .B(_1345_),
    .Y(_1346_));
 sg13g2_nand2_1 _4608_ (.Y(_1347_),
    .A(_1343_),
    .B(_1345_));
 sg13g2_or3_1 _4609_ (.A(_1003_),
    .B(_1121_),
    .C(_1122_),
    .X(_1348_));
 sg13g2_nand2_1 _4610_ (.Y(_1349_),
    .A(_1123_),
    .B(_1348_));
 sg13g2_xor2_1 _4611_ (.B(_1328_),
    .A(_1319_),
    .X(_1350_));
 sg13g2_nand2_1 _4612_ (.Y(_1351_),
    .A(_1349_),
    .B(_1350_));
 sg13g2_inv_1 _4613_ (.Y(_1352_),
    .A(_1351_));
 sg13g2_or2_1 _4614_ (.X(_1353_),
    .B(_1350_),
    .A(_1349_));
 sg13g2_nand2_1 _4615_ (.Y(_1354_),
    .A(_1351_),
    .B(_1353_));
 sg13g2_nand3_1 _4616_ (.B(_1119_),
    .C(_1120_),
    .A(_1026_),
    .Y(_1355_));
 sg13g2_nor2b_1 _4617_ (.A(_1121_),
    .B_N(_1355_),
    .Y(_1356_));
 sg13g2_xnor2_1 _4618_ (.Y(_1357_),
    .A(_1317_),
    .B(_1318_));
 sg13g2_nor2_1 _4619_ (.A(_1356_),
    .B(_1357_),
    .Y(_1358_));
 sg13g2_and2_1 _4620_ (.A(_1356_),
    .B(_1357_),
    .X(_1359_));
 sg13g2_nor2_1 _4621_ (.A(_1358_),
    .B(_1359_),
    .Y(_1360_));
 sg13g2_nor2b_1 _4622_ (.A(_1354_),
    .B_N(_1360_),
    .Y(_1361_));
 sg13g2_or3_1 _4623_ (.A(_1046_),
    .B(_1117_),
    .C(_1118_),
    .X(_1362_));
 sg13g2_nand2_1 _4624_ (.Y(_1363_),
    .A(_1119_),
    .B(_1362_));
 sg13g2_xnor2_1 _4625_ (.Y(_1364_),
    .A(_1314_),
    .B(_1315_));
 sg13g2_nand2_1 _4626_ (.Y(_1365_),
    .A(_1363_),
    .B(_1364_));
 sg13g2_nor2_1 _4627_ (.A(_1363_),
    .B(_1364_),
    .Y(_1366_));
 sg13g2_inv_1 _4628_ (.Y(_1367_),
    .A(_1366_));
 sg13g2_nand2_1 _4629_ (.Y(_1368_),
    .A(_1365_),
    .B(_1367_));
 sg13g2_nand3_1 _4630_ (.B(_1115_),
    .C(_1116_),
    .A(_1066_),
    .Y(_1369_));
 sg13g2_nor2b_1 _4631_ (.A(_1117_),
    .B_N(_1369_),
    .Y(_1370_));
 sg13g2_xnor2_1 _4632_ (.Y(_1371_),
    .A(_1312_),
    .B(_1313_));
 sg13g2_nor2_1 _4633_ (.A(_1370_),
    .B(_1371_),
    .Y(_1372_));
 sg13g2_inv_1 _4634_ (.Y(_1373_),
    .A(_1372_));
 sg13g2_nand2_1 _4635_ (.Y(_1374_),
    .A(_1370_),
    .B(_1371_));
 sg13g2_nor2b_1 _4636_ (.A(_1372_),
    .B_N(_1374_),
    .Y(_1375_));
 sg13g2_nor2b_1 _4637_ (.A(_1368_),
    .B_N(_1375_),
    .Y(_1376_));
 sg13g2_nand3_1 _4638_ (.B(_1113_),
    .C(_1114_),
    .A(_1082_),
    .Y(_1377_));
 sg13g2_and2_1 _4639_ (.A(_1115_),
    .B(_1377_),
    .X(_1378_));
 sg13g2_xor2_1 _4640_ (.B(_1310_),
    .A(_1309_),
    .X(_1379_));
 sg13g2_nor2_1 _4641_ (.A(_1378_),
    .B(_1379_),
    .Y(_1380_));
 sg13g2_nand2_1 _4642_ (.Y(_1381_),
    .A(_1378_),
    .B(_1379_));
 sg13g2_nor2b_1 _4643_ (.A(_1380_),
    .B_N(_1381_),
    .Y(_1382_));
 sg13g2_or3_1 _4644_ (.A(_1092_),
    .B(_1110_),
    .C(_1112_),
    .X(_1383_));
 sg13g2_nand2_1 _4645_ (.Y(_1384_),
    .A(_1113_),
    .B(_1383_));
 sg13g2_xnor2_1 _4646_ (.Y(_1385_),
    .A(_1306_),
    .B(_1307_));
 sg13g2_and2_1 _4647_ (.A(_1384_),
    .B(_1385_),
    .X(_1386_));
 sg13g2_nand2_1 _4648_ (.Y(_1387_),
    .A(_1384_),
    .B(_1385_));
 sg13g2_nor2_1 _4649_ (.A(_1384_),
    .B(_1385_),
    .Y(_1388_));
 sg13g2_inv_1 _4650_ (.Y(_1389_),
    .A(_1388_));
 sg13g2_nor2_1 _4651_ (.A(_1386_),
    .B(_1388_),
    .Y(_1390_));
 sg13g2_and2_1 _4652_ (.A(_1382_),
    .B(_1390_),
    .X(_1391_));
 sg13g2_xor2_1 _4653_ (.B(_1109_),
    .A(_1108_),
    .X(_1392_));
 sg13g2_xnor2_1 _4654_ (.Y(_1393_),
    .A(_1304_),
    .B(_1305_));
 sg13g2_or2_1 _4655_ (.X(_1394_),
    .B(_1393_),
    .A(_1392_));
 sg13g2_nand2_1 _4656_ (.Y(_1395_),
    .A(_1392_),
    .B(_1393_));
 sg13g2_nand2_1 _4657_ (.Y(_1396_),
    .A(_1394_),
    .B(_1395_));
 sg13g2_nand3_1 _4658_ (.B(_1300_),
    .C(_1303_),
    .A(_1295_),
    .Y(_1397_));
 sg13g2_xor2_1 _4659_ (.B(_1106_),
    .A(_1105_),
    .X(_1398_));
 sg13g2_nand3_1 _4660_ (.B(_1397_),
    .C(_1398_),
    .A(_1304_),
    .Y(_1399_));
 sg13g2_a21oi_2 _4661_ (.B1(_1398_),
    .Y(_1400_),
    .A2(_1397_),
    .A1(_1304_));
 sg13g2_inv_1 _4662_ (.Y(_1401_),
    .A(_1400_));
 sg13g2_nand2_1 _4663_ (.Y(_1402_),
    .A(_1399_),
    .B(_1401_));
 sg13g2_nor2_1 _4664_ (.A(_1396_),
    .B(_1402_),
    .Y(_1403_));
 sg13g2_xor2_1 _4665_ (.B(_1104_),
    .A(_1103_),
    .X(_1404_));
 sg13g2_xor2_1 _4666_ (.B(_1302_),
    .A(_1301_),
    .X(_1405_));
 sg13g2_nor2b_1 _4667_ (.A(_1405_),
    .B_N(_1404_),
    .Y(_1406_));
 sg13g2_inv_1 _4668_ (.Y(_1407_),
    .A(_1406_));
 sg13g2_nor2b_1 _4669_ (.A(_1404_),
    .B_N(_1405_),
    .Y(_1408_));
 sg13g2_xor2_1 _4670_ (.B(_1297_),
    .A(_0904_),
    .X(_1409_));
 sg13g2_xor2_1 _4671_ (.B(_1102_),
    .A(_0908_),
    .X(_1410_));
 sg13g2_nand2b_1 _4672_ (.Y(_1411_),
    .B(_1410_),
    .A_N(_1409_));
 sg13g2_nor2b_1 _4673_ (.A(_1410_),
    .B_N(_1409_),
    .Y(_1412_));
 sg13g2_o21ai_1 _4674_ (.B1(_0914_),
    .Y(_1413_),
    .A1(_0901_),
    .A2(_0911_));
 sg13g2_a21o_1 _4675_ (.A2(_1413_),
    .A1(_1411_),
    .B1(_1412_),
    .X(_1414_));
 sg13g2_xnor2_1 _4676_ (.Y(_1415_),
    .A(_1409_),
    .B(_1410_));
 sg13g2_o21ai_1 _4677_ (.B1(_0912_),
    .Y(_1416_),
    .A1(_0902_),
    .A2(_0913_));
 sg13g2_nand2b_1 _4678_ (.Y(_1417_),
    .B(_1415_),
    .A_N(_1416_));
 sg13g2_o21ai_1 _4679_ (.B1(_1407_),
    .Y(_1418_),
    .A1(_1408_),
    .A2(_1414_));
 sg13g2_o21ai_1 _4680_ (.B1(_1418_),
    .Y(_1419_),
    .A1(_1406_),
    .A2(_1417_));
 sg13g2_inv_1 _4681_ (.Y(_1420_),
    .A(_1419_));
 sg13g2_nand2_1 _4682_ (.Y(_1421_),
    .A(_1403_),
    .B(_1419_));
 sg13g2_nand2b_1 _4683_ (.Y(_1422_),
    .B(_1395_),
    .A_N(_1399_));
 sg13g2_nand3_1 _4684_ (.B(_1421_),
    .C(_1422_),
    .A(_1394_),
    .Y(_1423_));
 sg13g2_a221oi_1 _4685_ (.B2(_1423_),
    .C1(_1380_),
    .B1(_1391_),
    .A1(_1381_),
    .Y(_1424_),
    .A2(_1386_));
 sg13g2_inv_1 _4686_ (.Y(_1425_),
    .A(_1424_));
 sg13g2_o21ai_1 _4687_ (.B1(_1365_),
    .Y(_1426_),
    .A1(_1366_),
    .A2(_1373_));
 sg13g2_a21oi_1 _4688_ (.A1(_1376_),
    .A2(_1425_),
    .Y(_1427_),
    .B1(_1426_));
 sg13g2_inv_1 _4689_ (.Y(_1428_),
    .A(_1427_));
 sg13g2_a221oi_1 _4690_ (.B2(_1428_),
    .C1(_1352_),
    .B1(_1361_),
    .A1(_1353_),
    .Y(_1429_),
    .A2(_1358_));
 sg13g2_nand2b_1 _4691_ (.Y(_1430_),
    .B(_1429_),
    .A_N(_1346_));
 sg13g2_and2_1 _4692_ (.A(_1347_),
    .B(_1430_),
    .X(_1431_));
 sg13g2_o21ai_1 _4693_ (.B1(_1342_),
    .Y(_1432_),
    .A1(_1341_),
    .A2(_1431_));
 sg13g2_mux2_1 _4694_ (.A0(_0902_),
    .A1(_0901_),
    .S(net532),
    .X(_1433_));
 sg13g2_xor2_1 _4695_ (.B(_1433_),
    .A(_0915_),
    .X(_0019_));
 sg13g2_mux2_1 _4696_ (.A0(_1416_),
    .A1(_1413_),
    .S(net532),
    .X(_1434_));
 sg13g2_xnor2_1 _4697_ (.Y(_0020_),
    .A(_1415_),
    .B(_1434_));
 sg13g2_nor2_1 _4698_ (.A(_1406_),
    .B(_1408_),
    .Y(_1435_));
 sg13g2_nor2b_1 _4699_ (.A(_1412_),
    .B_N(_1417_),
    .Y(_1436_));
 sg13g2_mux2_1 _4700_ (.A0(_1436_),
    .A1(_1414_),
    .S(net532),
    .X(_1437_));
 sg13g2_xnor2_1 _4701_ (.Y(_0021_),
    .A(_1435_),
    .B(_1437_));
 sg13g2_nand2_1 _4702_ (.Y(_1438_),
    .A(_1418_),
    .B(_1432_));
 sg13g2_o21ai_1 _4703_ (.B1(_1438_),
    .Y(_1439_),
    .A1(_1420_),
    .A2(net532));
 sg13g2_xnor2_1 _4704_ (.Y(_0022_),
    .A(_1402_),
    .B(_1439_));
 sg13g2_o21ai_1 _4705_ (.B1(_1399_),
    .Y(_1440_),
    .A1(_1400_),
    .A2(_1420_));
 sg13g2_nor2_1 _4706_ (.A(_1432_),
    .B(_1440_),
    .Y(_1441_));
 sg13g2_a21oi_1 _4707_ (.A1(_1399_),
    .A2(_1418_),
    .Y(_1442_),
    .B1(_1400_));
 sg13g2_a21oi_1 _4708_ (.A1(_1432_),
    .A2(_1442_),
    .Y(_1443_),
    .B1(_1441_));
 sg13g2_xnor2_1 _4709_ (.Y(_0023_),
    .A(_1396_),
    .B(_1443_));
 sg13g2_a22oi_1 _4710_ (.Y(_1444_),
    .B1(_1403_),
    .B2(_1418_),
    .A2(_1400_),
    .A1(_1394_));
 sg13g2_nand2_1 _4711_ (.Y(_1445_),
    .A(_1395_),
    .B(_1444_));
 sg13g2_mux2_1 _4712_ (.A0(_1423_),
    .A1(_1445_),
    .S(net532),
    .X(_1446_));
 sg13g2_xor2_1 _4713_ (.B(_1446_),
    .A(_1390_),
    .X(_0024_));
 sg13g2_o21ai_1 _4714_ (.B1(_1387_),
    .Y(_1447_),
    .A1(_1388_),
    .A2(_1445_));
 sg13g2_o21ai_1 _4715_ (.B1(_1389_),
    .Y(_1448_),
    .A1(_1386_),
    .A2(_1423_));
 sg13g2_mux2_1 _4716_ (.A0(_1448_),
    .A1(_1447_),
    .S(net532),
    .X(_1449_));
 sg13g2_xnor2_1 _4717_ (.Y(_0025_),
    .A(_1382_),
    .B(_1449_));
 sg13g2_o21ai_1 _4718_ (.B1(_1381_),
    .Y(_1450_),
    .A1(_1380_),
    .A2(_1389_));
 sg13g2_a21oi_1 _4719_ (.A1(_1391_),
    .A2(_1445_),
    .Y(_1451_),
    .B1(_1450_));
 sg13g2_inv_1 _4720_ (.Y(_1452_),
    .A(_1451_));
 sg13g2_nor2_1 _4721_ (.A(_1424_),
    .B(net532),
    .Y(_1453_));
 sg13g2_a21oi_1 _4722_ (.A1(net531),
    .A2(_1452_),
    .Y(_1454_),
    .B1(_1453_));
 sg13g2_xnor2_1 _4723_ (.Y(_0026_),
    .A(_1375_),
    .B(_1454_));
 sg13g2_o21ai_1 _4724_ (.B1(_1374_),
    .Y(_1455_),
    .A1(_1372_),
    .A2(_1425_));
 sg13g2_o21ai_1 _4725_ (.B1(_1374_),
    .Y(_1456_),
    .A1(_1372_),
    .A2(_1451_));
 sg13g2_nand2_1 _4726_ (.Y(_1457_),
    .A(net531),
    .B(_1456_));
 sg13g2_o21ai_1 _4727_ (.B1(_1457_),
    .Y(_1458_),
    .A1(net531),
    .A2(_1455_));
 sg13g2_xnor2_1 _4728_ (.Y(_0027_),
    .A(_1368_),
    .B(_1458_));
 sg13g2_nand2_1 _4729_ (.Y(_1459_),
    .A(_1367_),
    .B(_1374_));
 sg13g2_a22oi_1 _4730_ (.Y(_1460_),
    .B1(_1459_),
    .B2(_1365_),
    .A2(_1452_),
    .A1(_1376_));
 sg13g2_nand2_1 _4731_ (.Y(_1461_),
    .A(net531),
    .B(_1460_));
 sg13g2_o21ai_1 _4732_ (.B1(_1461_),
    .Y(_1462_),
    .A1(_1428_),
    .A2(net531));
 sg13g2_xnor2_1 _4733_ (.Y(_0015_),
    .A(_1360_),
    .B(_1462_));
 sg13g2_nor2_1 _4734_ (.A(_1358_),
    .B(_1460_),
    .Y(_1463_));
 sg13g2_nor2_1 _4735_ (.A(_1358_),
    .B(_1428_),
    .Y(_1464_));
 sg13g2_nor3_1 _4736_ (.A(_1359_),
    .B(net531),
    .C(_1464_),
    .Y(_1465_));
 sg13g2_o21ai_1 _4737_ (.B1(net531),
    .Y(_1466_),
    .A1(_1359_),
    .A2(_1463_));
 sg13g2_nand2b_1 _4738_ (.Y(_1467_),
    .B(_1466_),
    .A_N(_1465_));
 sg13g2_xnor2_1 _4739_ (.Y(_0016_),
    .A(_1354_),
    .B(_1467_));
 sg13g2_nor2b_1 _4740_ (.A(_1346_),
    .B_N(_1347_),
    .Y(_1468_));
 sg13g2_nor2b_1 _4741_ (.A(_1460_),
    .B_N(_1361_),
    .Y(_1469_));
 sg13g2_a21oi_1 _4742_ (.A1(_1351_),
    .A2(_1359_),
    .Y(_1470_),
    .B1(_1469_));
 sg13g2_and2_1 _4743_ (.A(_1353_),
    .B(_1470_),
    .X(_1471_));
 sg13g2_mux2_1 _4744_ (.A0(_1429_),
    .A1(_1471_),
    .S(net531),
    .X(_1472_));
 sg13g2_xnor2_1 _4745_ (.Y(_0017_),
    .A(_1468_),
    .B(_1472_));
 sg13g2_nand2_1 _4746_ (.Y(_1473_),
    .A(_1347_),
    .B(_1471_));
 sg13g2_nor2_1 _4747_ (.A(_1342_),
    .B(_1346_),
    .Y(_1474_));
 sg13g2_a22oi_1 _4748_ (.Y(_1475_),
    .B1(_1473_),
    .B2(_1474_),
    .A2(_1431_),
    .A1(_1341_));
 sg13g2_inv_1 _4749_ (.Y(_0018_),
    .A(_1475_));
 sg13g2_mux2_1 _4750_ (.A0(_0255_),
    .A1(_0257_),
    .S(_0556_),
    .X(_1476_));
 sg13g2_xnor2_1 _4751_ (.Y(_0036_),
    .A(_0520_),
    .B(_1476_));
 sg13g2_nand2_1 _4752_ (.Y(_1477_),
    .A(_1850_),
    .B(_0516_));
 sg13g2_o21ai_1 _4753_ (.B1(_1477_),
    .Y(_1478_),
    .A1(_0256_),
    .A2(_0520_));
 sg13g2_mux2_1 _4754_ (.A0(_0524_),
    .A1(_1478_),
    .S(_0556_),
    .X(_1479_));
 sg13g2_xor2_1 _4755_ (.B(_1479_),
    .A(_0527_),
    .X(_0037_));
 sg13g2_nor2_1 _4756_ (.A(net681),
    .B(_0513_),
    .Y(_1480_));
 sg13g2_a21oi_1 _4757_ (.A1(_0527_),
    .A2(_1478_),
    .Y(_1481_),
    .B1(_1480_));
 sg13g2_mux2_1 _4758_ (.A0(_0528_),
    .A1(_1481_),
    .S(_0556_),
    .X(_1482_));
 sg13g2_xnor2_1 _4759_ (.Y(_0038_),
    .A(_0530_),
    .B(_1482_));
 sg13g2_a21oi_1 _4760_ (.A1(_0510_),
    .A2(_1481_),
    .Y(_1483_),
    .B1(_0508_));
 sg13g2_mux2_1 _4761_ (.A0(_0533_),
    .A1(_1483_),
    .S(_0556_),
    .X(_1484_));
 sg13g2_xnor2_1 _4762_ (.Y(_0039_),
    .A(_0500_),
    .B(_1484_));
 sg13g2_nor2_1 _4763_ (.A(\wirecube_top_inst.edge_function_inst.pixel_x_i[4] ),
    .B(_0499_),
    .Y(_1485_));
 sg13g2_a21o_1 _4764_ (.A2(_1483_),
    .A1(_0501_),
    .B1(_1485_),
    .X(_1486_));
 sg13g2_a21o_1 _4765_ (.A2(_0533_),
    .A1(_0501_),
    .B1(_0534_),
    .X(_1487_));
 sg13g2_mux2_1 _4766_ (.A0(_1486_),
    .A1(_1487_),
    .S(_0555_),
    .X(_1488_));
 sg13g2_xnor2_1 _4767_ (.Y(_0040_),
    .A(_0497_),
    .B(_1488_));
 sg13g2_a21oi_1 _4768_ (.A1(_0495_),
    .A2(_1486_),
    .Y(_1489_),
    .B1(_0496_));
 sg13g2_mux2_1 _4769_ (.A0(_0537_),
    .A1(_1489_),
    .S(_0556_),
    .X(_1490_));
 sg13g2_xnor2_1 _4770_ (.Y(_0041_),
    .A(_0558_),
    .B(_1490_));
 sg13g2_mux2_1 _4771_ (.A0(_0252_),
    .A1(_0253_),
    .S(_0555_),
    .X(_1491_));
 sg13g2_xnor2_1 _4772_ (.Y(_0029_),
    .A(_0460_),
    .B(_1491_));
 sg13g2_nor2_1 _4773_ (.A(\wirecube_top_inst.edge_function_inst.pixel_x_i[1] ),
    .B(_0457_),
    .Y(_1492_));
 sg13g2_a21o_1 _4774_ (.A2(_0459_),
    .A1(_0253_),
    .B1(_1492_),
    .X(_1493_));
 sg13g2_mux2_1 _4775_ (.A0(_0461_),
    .A1(_1493_),
    .S(_0555_),
    .X(_1494_));
 sg13g2_xor2_1 _4776_ (.B(_1494_),
    .A(_0462_),
    .X(_0030_));
 sg13g2_a22oi_1 _4777_ (.Y(_1495_),
    .B1(_0462_),
    .B2(_1493_),
    .A2(_0418_),
    .A1(_1849_));
 sg13g2_mux2_1 _4778_ (.A0(_0463_),
    .A1(_1495_),
    .S(_0555_),
    .X(_1496_));
 sg13g2_xor2_1 _4779_ (.B(_1496_),
    .A(_0484_),
    .X(_0031_));
 sg13g2_a21oi_1 _4780_ (.A1(_0409_),
    .A2(_1495_),
    .Y(_1497_),
    .B1(_0408_));
 sg13g2_mux2_1 _4781_ (.A0(_0465_),
    .A1(_1497_),
    .S(_0555_),
    .X(_1498_));
 sg13g2_xnor2_1 _4782_ (.Y(_0032_),
    .A(_0472_),
    .B(_1498_));
 sg13g2_a21oi_1 _4783_ (.A1(_0465_),
    .A2(_0473_),
    .Y(_1499_),
    .B1(_0474_));
 sg13g2_a22oi_1 _4784_ (.Y(_1500_),
    .B1(_0473_),
    .B2(_1497_),
    .A2(_0471_),
    .A1(_1847_));
 sg13g2_mux2_1 _4785_ (.A0(_1499_),
    .A1(_1500_),
    .S(_0555_),
    .X(_1501_));
 sg13g2_xor2_1 _4786_ (.B(_1501_),
    .A(_0478_),
    .X(_0033_));
 sg13g2_a21oi_1 _4787_ (.A1(_0399_),
    .A2(_1500_),
    .Y(_1502_),
    .B1(_0475_));
 sg13g2_mux2_1 _4788_ (.A0(_0481_),
    .A1(_1502_),
    .S(_0555_),
    .X(_1503_));
 sg13g2_xnor2_1 _4789_ (.Y(_0034_),
    .A(_0485_),
    .B(_1503_));
 sg13g2_nor2_1 _4790_ (.A(net113),
    .B(net628),
    .Y(_0043_));
 sg13g2_nor2_1 _4791_ (.A(net159),
    .B(net113),
    .Y(_1504_));
 sg13g2_nor3_1 _4792_ (.A(_1854_),
    .B(net628),
    .C(_1504_),
    .Y(_0044_));
 sg13g2_xnor2_1 _4793_ (.Y(_1505_),
    .A(net167),
    .B(_1854_));
 sg13g2_nor2_1 _4794_ (.A(net627),
    .B(_1505_),
    .Y(_0045_));
 sg13g2_a21oi_1 _4795_ (.A1(\wirecube_top_inst.counter_h[2] ),
    .A2(_1854_),
    .Y(_1506_),
    .B1(net151));
 sg13g2_nor3_1 _4796_ (.A(_1856_),
    .B(net628),
    .C(net152),
    .Y(_0046_));
 sg13g2_nor2_1 _4797_ (.A(net143),
    .B(_1856_),
    .Y(_1507_));
 sg13g2_nor3_1 _4798_ (.A(_1857_),
    .B(net627),
    .C(_1507_),
    .Y(_0047_));
 sg13g2_xor2_1 _4799_ (.B(_1857_),
    .A(net111),
    .X(_1508_));
 sg13g2_nor2_1 _4800_ (.A(net627),
    .B(net112),
    .Y(_0048_));
 sg13g2_nor3_1 _4801_ (.A(_1853_),
    .B(net120),
    .C(_1866_),
    .Y(_0049_));
 sg13g2_nand4_1 _4802_ (.B(\wirecube_top_inst.counter_h[5] ),
    .C(\wirecube_top_inst.counter_h[4] ),
    .A(\wirecube_top_inst.counter_h[6] ),
    .Y(_1509_),
    .D(_1863_));
 sg13g2_nand2b_1 _4803_ (.Y(_1510_),
    .B(net113),
    .A_N(\wirecube_top_inst.counter_h[1] ));
 sg13g2_nor4_2 _4804_ (.A(\wirecube_top_inst.counter_h[3] ),
    .B(\wirecube_top_inst.counter_h[2] ),
    .C(_1509_),
    .Y(_1511_),
    .D(_1510_));
 sg13g2_nor2_1 _4805_ (.A(net147),
    .B(_1511_),
    .Y(_0010_));
 sg13g2_nor3_1 _4806_ (.A(_2068_),
    .B(_2123_),
    .C(_1511_),
    .Y(_0011_));
 sg13g2_a21oi_1 _4807_ (.A1(net679),
    .A2(_2124_),
    .Y(_1512_),
    .B1(_2125_));
 sg13g2_nor2_2 _4808_ (.A(net655),
    .B(net646),
    .Y(_1513_));
 sg13g2_nor2_1 _4809_ (.A(net646),
    .B(_1512_),
    .Y(_0012_));
 sg13g2_nand2_1 _4810_ (.Y(_1514_),
    .A(net114),
    .B(_2124_));
 sg13g2_a21oi_1 _4811_ (.A1(net658),
    .A2(_1514_),
    .Y(_0013_),
    .B1(net646));
 sg13g2_nor4_2 _4812_ (.A(\wirecube_top_inst.counter_h[3] ),
    .B(\wirecube_top_inst.counter_h[2] ),
    .C(_1855_),
    .Y(_1515_),
    .D(_1509_));
 sg13g2_nor2_1 _4813_ (.A(net95),
    .B(_1515_),
    .Y(_0000_));
 sg13g2_and2_1 _4814_ (.A(net124),
    .B(net95),
    .X(_1516_));
 sg13g2_nand2_1 _4815_ (.Y(_1517_),
    .A(net124),
    .B(net95));
 sg13g2_nor2_1 _4816_ (.A(net124),
    .B(net95),
    .Y(_1518_));
 sg13g2_nor3_1 _4817_ (.A(_1515_),
    .B(_1516_),
    .C(_1518_),
    .Y(_0001_));
 sg13g2_nor3_1 _4818_ (.A(net126),
    .B(net145),
    .C(_1517_),
    .Y(_1519_));
 sg13g2_a21oi_1 _4819_ (.A1(net145),
    .A2(_1517_),
    .Y(_1520_),
    .B1(_1519_));
 sg13g2_nor2_1 _4820_ (.A(_1515_),
    .B(_1520_),
    .Y(_0002_));
 sg13g2_nor2_1 _4821_ (.A(net126),
    .B(_1516_),
    .Y(_1521_));
 sg13g2_nand2_2 _4822_ (.Y(_1522_),
    .A(net126),
    .B(_1516_));
 sg13g2_o21ai_1 _4823_ (.B1(_1522_),
    .Y(_1523_),
    .A1(net126),
    .A2(\wirecube_top_inst.linecounter_h[2] ));
 sg13g2_nor3_1 _4824_ (.A(_1515_),
    .B(_1521_),
    .C(_1523_),
    .Y(_0003_));
 sg13g2_o21ai_1 _4825_ (.B1(net116),
    .Y(_1524_),
    .A1(_1839_),
    .A2(_0628_));
 sg13g2_nand4_1 _4826_ (.B(net701),
    .C(\wirecube_top_inst.counter_v[7] ),
    .A(_1838_),
    .Y(_1525_),
    .D(net699));
 sg13g2_nand2b_1 _4827_ (.Y(_1526_),
    .B(_1525_),
    .A_N(net704));
 sg13g2_xor2_1 _4828_ (.B(net704),
    .A(\wirecube_top_inst.counter_v[0] ),
    .X(_1527_));
 sg13g2_nand2_1 _4829_ (.Y(_1528_),
    .A(net702),
    .B(net703));
 sg13g2_nor4_1 _4830_ (.A(net700),
    .B(_1840_),
    .C(_0631_),
    .D(_1528_),
    .Y(_1529_));
 sg13g2_nand4_1 _4831_ (.B(_1526_),
    .C(_1527_),
    .A(net117),
    .Y(\wirecube_top_inst.delay_inst_vsync.in_i ),
    .D(_1529_));
 sg13g2_nor3_1 _4832_ (.A(\wirecube_top_inst.counter_h[4] ),
    .B(\wirecube_top_inst.counter_h[3] ),
    .C(\wirecube_top_inst.counter_h[2] ),
    .Y(_1530_));
 sg13g2_nand3_1 _4833_ (.B(_1504_),
    .C(_1530_),
    .A(\wirecube_top_inst.counter_h[5] ),
    .Y(_1531_));
 sg13g2_nand3b_1 _4834_ (.B(net111),
    .C(_1531_),
    .Y(_1532_),
    .A_N(\wirecube_top_inst.counter_h[6] ));
 sg13g2_nand3_1 _4835_ (.B(_1863_),
    .C(_1532_),
    .A(net125),
    .Y(_1533_));
 sg13g2_nand3b_1 _4836_ (.B(net111),
    .C(_1531_),
    .Y(_1534_),
    .A_N(net119));
 sg13g2_nand3_1 _4837_ (.B(_1533_),
    .C(_1534_),
    .A(_0623_),
    .Y(\wirecube_top_inst.delay_inst_hsync.in_i ));
 sg13g2_xor2_1 _4838_ (.B(_0603_),
    .A(_2546_),
    .X(_0075_));
 sg13g2_o21ai_1 _4839_ (.B1(_0594_),
    .Y(_1535_),
    .A1(_0602_),
    .A2(_0604_));
 sg13g2_or3_1 _4840_ (.A(_0594_),
    .B(_0602_),
    .C(_0604_),
    .X(_1536_));
 sg13g2_and2_1 _4841_ (.A(_1535_),
    .B(_1536_),
    .X(_0076_));
 sg13g2_o21ai_1 _4842_ (.B1(_1535_),
    .Y(_1537_),
    .A1(\wirecube_top_inst.edge_function_inst.pixel_y_i[2] ),
    .A2(_0593_));
 sg13g2_xnor2_1 _4843_ (.Y(_0077_),
    .A(_0612_),
    .B(_1537_));
 sg13g2_o21ai_1 _4844_ (.B1(_0591_),
    .Y(_1538_),
    .A1(_0605_),
    .A2(_1537_));
 sg13g2_xor2_1 _4845_ (.B(_1538_),
    .A(_0609_),
    .X(_0078_));
 sg13g2_or2_1 _4846_ (.X(_1539_),
    .B(_0608_),
    .A(\wirecube_top_inst.edge_function_inst.pixel_y_i[4] ));
 sg13g2_o21ai_1 _4847_ (.B1(_1539_),
    .Y(_1540_),
    .A1(_0609_),
    .A2(_1538_));
 sg13g2_xor2_1 _4848_ (.B(_1540_),
    .A(_0599_),
    .X(_0079_));
 sg13g2_a21oi_1 _4849_ (.A1(_0597_),
    .A2(_1540_),
    .Y(_1541_),
    .B1(_0598_));
 sg13g2_xnor2_1 _4850_ (.Y(_0080_),
    .A(_0589_),
    .B(_1541_));
 sg13g2_xnor2_1 _4851_ (.Y(_0082_),
    .A(_0155_),
    .B(_0575_));
 sg13g2_xor2_1 _4852_ (.B(_0577_),
    .A(_0576_),
    .X(_0083_));
 sg13g2_xor2_1 _4853_ (.B(_0579_),
    .A(_0578_),
    .X(_0084_));
 sg13g2_xor2_1 _4854_ (.B(_0581_),
    .A(_0580_),
    .X(_0085_));
 sg13g2_xor2_1 _4855_ (.B(_0583_),
    .A(_0582_),
    .X(_0086_));
 sg13g2_xor2_1 _4856_ (.B(_0585_),
    .A(_0584_),
    .X(_0087_));
 sg13g2_nor2_1 _4857_ (.A(_1841_),
    .B(net109),
    .Y(_1542_));
 sg13g2_nor4_2 _4858_ (.A(_1841_),
    .B(net109),
    .C(net179),
    .Y(_1543_),
    .D(net626));
 sg13g2_nor4_1 _4859_ (.A(\wirecube_top_inst.counter_v[0] ),
    .B(net704),
    .C(\wirecube_top_inst.counter_v[10] ),
    .D(\wirecube_top_inst.counter_v[9] ),
    .Y(_1544_));
 sg13g2_nand3_1 _4860_ (.B(_0630_),
    .C(_1544_),
    .A(_0625_),
    .Y(_1545_));
 sg13g2_nor4_2 _4861_ (.A(\wirecube_top_inst.counter_v[7] ),
    .B(net155),
    .C(\wirecube_top_inst.counter_v[8] ),
    .Y(_1546_),
    .D(_1545_));
 sg13g2_nand2_1 _4862_ (.Y(_1547_),
    .A(net130),
    .B(_1543_));
 sg13g2_xnor2_1 _4863_ (.Y(_1548_),
    .A(net130),
    .B(_1543_));
 sg13g2_nor2_1 _4864_ (.A(_1546_),
    .B(net131),
    .Y(_0108_));
 sg13g2_xnor2_1 _4865_ (.Y(_1549_),
    .A(_1845_),
    .B(_1547_));
 sg13g2_nor2_1 _4866_ (.A(net156),
    .B(_1549_),
    .Y(_0109_));
 sg13g2_nor2_2 _4867_ (.A(_1543_),
    .B(_1546_),
    .Y(_1550_));
 sg13g2_nor2b_2 _4868_ (.A(_1546_),
    .B_N(_1543_),
    .Y(_1551_));
 sg13g2_nand2_2 _4869_ (.Y(_1552_),
    .A(net130),
    .B(\wirecube_top_inst.edge_function_inst.pixel_y_i[1] ));
 sg13g2_xor2_1 _4870_ (.B(_1552_),
    .A(_0053_),
    .X(_1553_));
 sg13g2_a22oi_1 _4871_ (.Y(_1554_),
    .B1(_1551_),
    .B2(_1553_),
    .A2(_1550_),
    .A1(net149));
 sg13g2_inv_1 _4872_ (.Y(_0110_),
    .A(net150));
 sg13g2_or3_1 _4873_ (.A(_1844_),
    .B(_1550_),
    .C(_1552_),
    .X(_1555_));
 sg13g2_nor3_2 _4874_ (.A(_1843_),
    .B(_1844_),
    .C(_1552_),
    .Y(_1556_));
 sg13g2_a221oi_1 _4875_ (.B2(_1543_),
    .C1(net156),
    .B1(_1556_),
    .A1(_1843_),
    .Y(_0111_),
    .A2(_1555_));
 sg13g2_nor2b_1 _4876_ (.A(_0052_),
    .B_N(_1556_),
    .Y(_1557_));
 sg13g2_xnor2_1 _4877_ (.Y(_1558_),
    .A(_0052_),
    .B(_1556_));
 sg13g2_a22oi_1 _4878_ (.Y(_1559_),
    .B1(_1551_),
    .B2(_1558_),
    .A2(_1550_),
    .A1(net153));
 sg13g2_inv_1 _4879_ (.Y(_0112_),
    .A(net154));
 sg13g2_xnor2_1 _4880_ (.Y(_1560_),
    .A(_0054_),
    .B(_1557_));
 sg13g2_a22oi_1 _4881_ (.Y(_1561_),
    .B1(_1551_),
    .B2(_1560_),
    .A2(_1550_),
    .A1(net122));
 sg13g2_inv_1 _4882_ (.Y(_0113_),
    .A(net123));
 sg13g2_nand3_1 _4883_ (.B(\wirecube_top_inst.edge_function_inst.pixel_y_i[4] ),
    .C(_1556_),
    .A(\wirecube_top_inst.edge_function_inst.pixel_y_i[5] ),
    .Y(_1562_));
 sg13g2_xor2_1 _4884_ (.B(_1562_),
    .A(_0051_),
    .X(_1563_));
 sg13g2_a22oi_1 _4885_ (.Y(_1564_),
    .B1(_1551_),
    .B2(_1563_),
    .A2(_1550_),
    .A1(net107));
 sg13g2_inv_1 _4886_ (.Y(_0114_),
    .A(net108));
 sg13g2_nand3_1 _4887_ (.B(net703),
    .C(_0626_),
    .A(net702),
    .Y(_1565_));
 sg13g2_nor2_1 _4888_ (.A(_1839_),
    .B(_1565_),
    .Y(_1566_));
 sg13g2_nor3_2 _4889_ (.A(_1838_),
    .B(_1839_),
    .C(_1565_),
    .Y(_1567_));
 sg13g2_nand2_1 _4890_ (.Y(_1568_),
    .A(net700),
    .B(_1566_));
 sg13g2_nor2_2 _4891_ (.A(_0628_),
    .B(_1568_),
    .Y(_1569_));
 sg13g2_nand2b_2 _4892_ (.Y(_1570_),
    .B(_1569_),
    .A_N(_0631_));
 sg13g2_and2_1 _4893_ (.A(net626),
    .B(_1570_),
    .X(_1571_));
 sg13g2_nand2_1 _4894_ (.Y(_1572_),
    .A(net115),
    .B(_1571_));
 sg13g2_nand2_1 _4895_ (.Y(_1573_),
    .A(net627),
    .B(_1570_));
 sg13g2_o21ai_1 _4896_ (.B1(_1572_),
    .Y(_0115_),
    .A1(net115),
    .A2(_1573_));
 sg13g2_nand2_1 _4897_ (.Y(_1574_),
    .A(net109),
    .B(_1571_));
 sg13g2_nor2b_1 _4898_ (.A(\wirecube_top_inst.subcounter_v[0] ),
    .B_N(net109),
    .Y(_1575_));
 sg13g2_a21oi_1 _4899_ (.A1(_0050_),
    .A2(_1542_),
    .Y(_1576_),
    .B1(_1575_));
 sg13g2_o21ai_1 _4900_ (.B1(_1574_),
    .Y(_0116_),
    .A1(_1573_),
    .A2(_1576_));
 sg13g2_xor2_1 _4901_ (.B(_0050_),
    .A(\wirecube_top_inst.subcounter_v[0] ),
    .X(_1577_));
 sg13g2_nor3_1 _4902_ (.A(_1542_),
    .B(_1573_),
    .C(_1577_),
    .Y(_1578_));
 sg13g2_a21o_1 _4903_ (.A2(_1571_),
    .A1(net97),
    .B1(_1578_),
    .X(_0117_));
 sg13g2_a21oi_1 _4904_ (.A1(net700),
    .A2(_0629_),
    .Y(_1579_),
    .B1(\wirecube_top_inst.counter_v[9] ));
 sg13g2_nor2_1 _4905_ (.A(\wirecube_top_inst.counter_v[10] ),
    .B(_1579_),
    .Y(_1580_));
 sg13g2_nor4_1 _4906_ (.A(\wirecube_top_inst.counter_v[10] ),
    .B(\wirecube_top_inst.counter_v[9] ),
    .C(_0624_),
    .D(_1565_),
    .Y(_1581_));
 sg13g2_a21oi_2 _4907_ (.B1(_1580_),
    .Y(_1582_),
    .A2(_1581_),
    .A1(_0629_));
 sg13g2_nand2_2 _4908_ (.Y(_1583_),
    .A(net628),
    .B(_1582_));
 sg13g2_inv_1 _4909_ (.Y(_1584_),
    .A(_1583_));
 sg13g2_a22oi_1 _4910_ (.Y(_1585_),
    .B1(_1584_),
    .B2(\wirecube_top_inst.counter_v[0] ),
    .A2(net625),
    .A1(net89));
 sg13g2_inv_1 _4911_ (.Y(_0118_),
    .A(net90));
 sg13g2_nand2_1 _4912_ (.Y(_1586_),
    .A(net81),
    .B(net625));
 sg13g2_o21ai_1 _4913_ (.B1(_1586_),
    .Y(_0119_),
    .A1(_1527_),
    .A2(_1583_));
 sg13g2_and3_1 _4914_ (.X(_1587_),
    .A(net703),
    .B(net628),
    .C(_0626_));
 sg13g2_nor2_2 _4915_ (.A(net626),
    .B(_1582_),
    .Y(_1588_));
 sg13g2_a21oi_1 _4916_ (.A1(net628),
    .A2(_0626_),
    .Y(_1589_),
    .B1(net703));
 sg13g2_nor3_1 _4917_ (.A(_1587_),
    .B(_1588_),
    .C(_1589_),
    .Y(_0120_));
 sg13g2_nor2_1 _4918_ (.A(net702),
    .B(_1587_),
    .Y(_1590_));
 sg13g2_nor2_1 _4919_ (.A(net625),
    .B(_1565_),
    .Y(_1591_));
 sg13g2_nor3_1 _4920_ (.A(_1588_),
    .B(_1590_),
    .C(_1591_),
    .Y(_0121_));
 sg13g2_nand2_1 _4921_ (.Y(_1592_),
    .A(net87),
    .B(net626));
 sg13g2_xnor2_1 _4922_ (.Y(_1593_),
    .A(net701),
    .B(_1565_));
 sg13g2_o21ai_1 _4923_ (.B1(_1592_),
    .Y(_0122_),
    .A1(_1583_),
    .A2(_1593_));
 sg13g2_nor2_1 _4924_ (.A(net625),
    .B(_1568_),
    .Y(_1594_));
 sg13g2_a21oi_1 _4925_ (.A1(net628),
    .A2(_1566_),
    .Y(_1595_),
    .B1(net700));
 sg13g2_nor3_1 _4926_ (.A(_1588_),
    .B(_1594_),
    .C(net176),
    .Y(_0123_));
 sg13g2_nand2_1 _4927_ (.Y(_1596_),
    .A(net85),
    .B(net625));
 sg13g2_xor2_1 _4928_ (.B(_1567_),
    .A(net699),
    .X(_1597_));
 sg13g2_o21ai_1 _4929_ (.B1(_1596_),
    .Y(_0124_),
    .A1(_1583_),
    .A2(_1597_));
 sg13g2_nand2_1 _4930_ (.Y(_1598_),
    .A(net93),
    .B(net625));
 sg13g2_nand3_1 _4931_ (.B(net699),
    .C(_1567_),
    .A(\wirecube_top_inst.counter_v[7] ),
    .Y(_1599_));
 sg13g2_a21o_1 _4932_ (.A2(_1567_),
    .A1(net699),
    .B1(\wirecube_top_inst.counter_v[7] ),
    .X(_1600_));
 sg13g2_and2_1 _4933_ (.A(_1599_),
    .B(_1600_),
    .X(_1601_));
 sg13g2_o21ai_1 _4934_ (.B1(_1598_),
    .Y(_0125_),
    .A1(_1583_),
    .A2(_1601_));
 sg13g2_nand2_1 _4935_ (.Y(_1602_),
    .A(net83),
    .B(net626));
 sg13g2_a21oi_1 _4936_ (.A1(_1840_),
    .A2(_1599_),
    .Y(_1603_),
    .B1(_1569_));
 sg13g2_o21ai_1 _4937_ (.B1(_1602_),
    .Y(_0126_),
    .A1(_1583_),
    .A2(_1603_));
 sg13g2_nand2_1 _4938_ (.Y(_1604_),
    .A(net79),
    .B(net625));
 sg13g2_xor2_1 _4939_ (.B(_1569_),
    .A(\wirecube_top_inst.counter_v[9] ),
    .X(_1605_));
 sg13g2_o21ai_1 _4940_ (.B1(_1604_),
    .Y(_0127_),
    .A1(_1583_),
    .A2(_1605_));
 sg13g2_a21o_1 _4941_ (.A2(_1569_),
    .A1(\wirecube_top_inst.counter_v[9] ),
    .B1(\wirecube_top_inst.counter_v[10] ),
    .X(_1606_));
 sg13g2_a21oi_1 _4942_ (.A1(_1570_),
    .A2(_1606_),
    .Y(_1607_),
    .B1(_1583_));
 sg13g2_a21o_1 _4943_ (.A2(net625),
    .A1(net99),
    .B1(_1607_),
    .X(_0128_));
 sg13g2_mux2_1 _4944_ (.A0(\wirecube_top_inst.frame_cnt[0] ),
    .A1(net77),
    .S(_1588_),
    .X(_0129_));
 sg13g2_and3_2 _4945_ (.X(_1608_),
    .A(net136),
    .B(net698),
    .C(_1588_));
 sg13g2_a21oi_1 _4946_ (.A1(net136),
    .A2(_1588_),
    .Y(_1609_),
    .B1(net698));
 sg13g2_nor2_1 _4947_ (.A(_1608_),
    .B(net137),
    .Y(_0130_));
 sg13g2_xor2_1 _4948_ (.B(_1608_),
    .A(net697),
    .X(_0131_));
 sg13g2_nand2_1 _4949_ (.Y(_1610_),
    .A(_1837_),
    .B(_1608_));
 sg13g2_xnor2_1 _4950_ (.Y(_0132_),
    .A(net696),
    .B(_1610_));
 sg13g2_nand3_1 _4951_ (.B(net697),
    .C(_1608_),
    .A(net696),
    .Y(_1611_));
 sg13g2_inv_1 _4952_ (.Y(_1612_),
    .A(_1611_));
 sg13g2_xnor2_1 _4953_ (.Y(_0133_),
    .A(net695),
    .B(_1611_));
 sg13g2_nor2_1 _4954_ (.A(net157),
    .B(_1611_),
    .Y(_1613_));
 sg13g2_xor2_1 _4955_ (.B(_1613_),
    .A(net694),
    .X(_0134_));
 sg13g2_and3_2 _4956_ (.X(_1614_),
    .A(net694),
    .B(net695),
    .C(_1612_));
 sg13g2_and2_1 _4957_ (.A(net692),
    .B(_1614_),
    .X(_1615_));
 sg13g2_xnor2_1 _4958_ (.Y(_0135_),
    .A(_1804_),
    .B(_1614_));
 sg13g2_nor2b_2 _4959_ (.A(net190),
    .B_N(_1614_),
    .Y(_1616_));
 sg13g2_xnor2_1 _4960_ (.Y(_0136_),
    .A(_1793_),
    .B(_1616_));
 sg13g2_nand2_1 _4961_ (.Y(_1617_),
    .A(net689),
    .B(_1615_));
 sg13g2_nand3_1 _4962_ (.B(_1922_),
    .C(_1614_),
    .A(net687),
    .Y(_1618_));
 sg13g2_xnor2_1 _4963_ (.Y(_0137_),
    .A(net687),
    .B(_1617_));
 sg13g2_a22oi_1 _4964_ (.Y(_0138_),
    .B1(_1618_),
    .B2(_1813_),
    .A2(_1615_),
    .A1(_1941_));
 sg13g2_nor2_2 _4965_ (.A(_1879_),
    .B(_1617_),
    .Y(_1619_));
 sg13g2_inv_1 _4966_ (.Y(_1620_),
    .A(_1619_));
 sg13g2_xnor2_1 _4967_ (.Y(_0139_),
    .A(_1821_),
    .B(_1619_));
 sg13g2_o21ai_1 _4968_ (.B1(net683),
    .Y(_1621_),
    .A1(_1821_),
    .A2(_1620_));
 sg13g2_o21ai_1 _4969_ (.B1(_1621_),
    .Y(_0140_),
    .A1(_1896_),
    .A2(_1620_));
 sg13g2_nand2b_1 _4970_ (.Y(_1622_),
    .B(_1619_),
    .A_N(_1890_));
 sg13g2_xnor2_1 _4971_ (.Y(_0141_),
    .A(net101),
    .B(_1622_));
 sg13g2_nor2_1 _4972_ (.A(\wirecube_top_inst.linecounter_h[2] ),
    .B(_1522_),
    .Y(_1623_));
 sg13g2_nand2_1 _4973_ (.Y(_1624_),
    .A(net674),
    .B(_1623_));
 sg13g2_nor2_1 _4974_ (.A(net102),
    .B(_1624_),
    .Y(_1625_));
 sg13g2_nand2_2 _4975_ (.Y(_1626_),
    .A(_2062_),
    .B(_2152_));
 sg13g2_nor2_1 _4976_ (.A(_2087_),
    .B(_2141_),
    .Y(_1627_));
 sg13g2_nand4_1 _4977_ (.B(_2372_),
    .C(_2383_),
    .A(_2300_),
    .Y(_1628_),
    .D(_1627_));
 sg13g2_and2_1 _4978_ (.A(net662),
    .B(_2127_),
    .X(_1629_));
 sg13g2_nand2_1 _4979_ (.Y(_1630_),
    .A(net662),
    .B(net658));
 sg13g2_nor2_1 _4980_ (.A(_2064_),
    .B(_2128_),
    .Y(_1631_));
 sg13g2_nand2_1 _4981_ (.Y(_1632_),
    .A(_2065_),
    .B(_2129_));
 sg13g2_a21oi_1 _4982_ (.A1(_1629_),
    .A2(_1631_),
    .Y(_1633_),
    .B1(_0161_));
 sg13g2_a21oi_1 _4983_ (.A1(_1626_),
    .A2(_1628_),
    .Y(_1634_),
    .B1(_1633_));
 sg13g2_nor3_1 _4984_ (.A(net566),
    .B(_2187_),
    .C(net540),
    .Y(_1635_));
 sg13g2_nand4_1 _4985_ (.B(_2320_),
    .C(_0164_),
    .A(_2078_),
    .Y(_1636_),
    .D(_1635_));
 sg13g2_o21ai_1 _4986_ (.B1(net677),
    .Y(_1637_),
    .A1(_2044_),
    .A2(_1636_));
 sg13g2_o21ai_1 _4987_ (.B1(_2067_),
    .Y(_1638_),
    .A1(net679),
    .A2(_2124_));
 sg13g2_o21ai_1 _4988_ (.B1(_2182_),
    .Y(_1639_),
    .A1(_2102_),
    .A2(_1638_));
 sg13g2_nand3_1 _4989_ (.B(_1637_),
    .C(_1639_),
    .A(_1634_),
    .Y(_1640_));
 sg13g2_and2_2 _4990_ (.A(net636),
    .B(_1640_),
    .X(_1641_));
 sg13g2_inv_1 _4991_ (.Y(_1642_),
    .A(_1641_));
 sg13g2_a21oi_1 _4992_ (.A1(\wirecube_top_inst.edge_function_inst.absolute[6] ),
    .A2(_1642_),
    .Y(_1643_),
    .B1(\wirecube_top_inst.edge_function_inst.absolute[7] ));
 sg13g2_a21o_2 _4993_ (.A2(_2151_),
    .A1(_2104_),
    .B1(net546),
    .X(_1644_));
 sg13g2_nor2_1 _4994_ (.A(_2126_),
    .B(net546),
    .Y(_1645_));
 sg13g2_a21o_1 _4995_ (.A2(_2149_),
    .A1(_2067_),
    .B1(net547),
    .X(_1646_));
 sg13g2_nor2b_2 _4996_ (.A(_1645_),
    .B_N(_1646_),
    .Y(_1647_));
 sg13g2_a22oi_1 _4997_ (.Y(_1648_),
    .B1(_1644_),
    .B2(_1647_),
    .A2(_2181_),
    .A1(_2043_));
 sg13g2_nand2_1 _4998_ (.Y(_1649_),
    .A(_2359_),
    .B(_1632_));
 sg13g2_nand3_1 _4999_ (.B(_2054_),
    .C(_2081_),
    .A(_2026_),
    .Y(_1650_));
 sg13g2_nor3_1 _5000_ (.A(_2173_),
    .B(_2214_),
    .C(_2256_),
    .Y(_1651_));
 sg13g2_nand2b_1 _5001_ (.Y(_1652_),
    .B(_1651_),
    .A_N(_1650_));
 sg13g2_nor3_1 _5002_ (.A(_2162_),
    .B(_2283_),
    .C(_2301_),
    .Y(_1653_));
 sg13g2_nand3b_1 _5003_ (.B(_1653_),
    .C(_2113_),
    .Y(_1654_),
    .A_N(_1652_));
 sg13g2_nor3_2 _5004_ (.A(_2048_),
    .B(_2087_),
    .C(_2206_),
    .Y(_1655_));
 sg13g2_nor4_1 _5005_ (.A(net575),
    .B(_2006_),
    .C(_2146_),
    .D(_1654_),
    .Y(_1656_));
 sg13g2_nand3_1 _5006_ (.B(_1655_),
    .C(_1656_),
    .A(_2296_),
    .Y(_1657_));
 sg13g2_nand2_1 _5007_ (.Y(_1658_),
    .A(_1630_),
    .B(_1657_));
 sg13g2_a221oi_1 _5008_ (.B2(_1658_),
    .C1(net588),
    .B1(_1649_),
    .A1(_2009_),
    .Y(_1659_),
    .A2(_2030_));
 sg13g2_nor2_1 _5009_ (.A(net555),
    .B(_2314_),
    .Y(_1660_));
 sg13g2_a21oi_1 _5010_ (.A1(_2080_),
    .A2(net677),
    .Y(_1661_),
    .B1(net547));
 sg13g2_and4_1 _5011_ (.A(_2372_),
    .B(_0258_),
    .C(_0341_),
    .D(_1661_),
    .X(_1662_));
 sg13g2_nor2_1 _5012_ (.A(net677),
    .B(_1626_),
    .Y(_1663_));
 sg13g2_nor2_1 _5013_ (.A(_2080_),
    .B(net547),
    .Y(_1664_));
 sg13g2_a21oi_1 _5014_ (.A1(_1660_),
    .A2(_1662_),
    .Y(_1665_),
    .B1(_1663_));
 sg13g2_nor3_2 _5015_ (.A(_1648_),
    .B(_1659_),
    .C(_1665_),
    .Y(_1666_));
 sg13g2_nor2_1 _5016_ (.A(net642),
    .B(_1666_),
    .Y(_1667_));
 sg13g2_and2_1 _5017_ (.A(_0063_),
    .B(_1667_),
    .X(_1668_));
 sg13g2_xor2_1 _5018_ (.B(_1667_),
    .A(\wirecube_top_inst.edge_function_inst.absolute[5] ),
    .X(_1669_));
 sg13g2_nand3_1 _5019_ (.B(_2081_),
    .C(_2084_),
    .A(_2019_),
    .Y(_1670_));
 sg13g2_nor3_1 _5020_ (.A(net566),
    .B(_2138_),
    .C(_1670_),
    .Y(_1671_));
 sg13g2_a21oi_2 _5021_ (.B1(_1644_),
    .Y(_1672_),
    .A2(_1671_),
    .A1(_2165_));
 sg13g2_nor4_1 _5022_ (.A(_2008_),
    .B(_2087_),
    .C(_2485_),
    .D(_1654_),
    .Y(_1673_));
 sg13g2_a21oi_1 _5023_ (.A1(_1657_),
    .A2(_1673_),
    .Y(_1674_),
    .B1(_1629_));
 sg13g2_nor4_2 _5024_ (.A(_2028_),
    .B(_2038_),
    .C(_2170_),
    .Y(_1675_),
    .D(_2256_));
 sg13g2_and2_1 _5025_ (.A(_2282_),
    .B(_1675_),
    .X(_1676_));
 sg13g2_nand4_1 _5026_ (.B(net560),
    .C(_2176_),
    .A(_2009_),
    .Y(_1677_),
    .D(_2265_));
 sg13g2_nor2_1 _5027_ (.A(_2485_),
    .B(_1677_),
    .Y(_1678_));
 sg13g2_nand3_1 _5028_ (.B(_1676_),
    .C(_1678_),
    .A(_2359_),
    .Y(_1679_));
 sg13g2_and4_1 _5029_ (.A(_2021_),
    .B(net556),
    .C(_2313_),
    .D(_0175_),
    .X(_1680_));
 sg13g2_nor4_2 _5030_ (.A(_2087_),
    .B(_2141_),
    .C(_2354_),
    .Y(_1681_),
    .D(_2498_));
 sg13g2_nand4_1 _5031_ (.B(_2331_),
    .C(_1680_),
    .A(_2207_),
    .Y(_1682_),
    .D(_1681_));
 sg13g2_o21ai_1 _5032_ (.B1(_1626_),
    .Y(_1683_),
    .A1(net546),
    .A2(_1682_));
 sg13g2_nand4_1 _5033_ (.B(_2313_),
    .C(_0271_),
    .A(_2282_),
    .Y(_1684_),
    .D(_1664_));
 sg13g2_nand4_1 _5034_ (.B(_2078_),
    .C(_2117_),
    .A(_1996_),
    .Y(_1685_),
    .D(net551));
 sg13g2_or4_1 _5035_ (.A(_2008_),
    .B(_2087_),
    .C(_1684_),
    .D(_1685_),
    .X(_1686_));
 sg13g2_nand2_1 _5036_ (.Y(_1687_),
    .A(_2079_),
    .B(_2136_));
 sg13g2_nor4_1 _5037_ (.A(_2018_),
    .B(_0161_),
    .C(_0225_),
    .D(_1687_),
    .Y(_1688_));
 sg13g2_nand4_1 _5038_ (.B(net557),
    .C(_0264_),
    .A(_2003_),
    .Y(_1689_),
    .D(_1688_));
 sg13g2_nand2b_1 _5039_ (.Y(_1690_),
    .B(_1689_),
    .A_N(_1647_));
 sg13g2_a22oi_1 _5040_ (.Y(_1691_),
    .B1(_1686_),
    .B2(net677),
    .A2(_1679_),
    .A1(_1632_));
 sg13g2_nand3_1 _5041_ (.B(_1690_),
    .C(_1691_),
    .A(_1683_),
    .Y(_1692_));
 sg13g2_nor3_2 _5042_ (.A(_1672_),
    .B(_1674_),
    .C(_1692_),
    .Y(_1693_));
 sg13g2_nor2_1 _5043_ (.A(net642),
    .B(_1693_),
    .Y(_1694_));
 sg13g2_a21oi_2 _5044_ (.B1(_1694_),
    .Y(_1695_),
    .A2(_1640_),
    .A1(net642));
 sg13g2_nand2b_1 _5045_ (.Y(_1696_),
    .B(_0064_),
    .A_N(_1695_));
 sg13g2_nand3_1 _5046_ (.B(_2196_),
    .C(_0258_),
    .A(_2022_),
    .Y(_1697_));
 sg13g2_nor4_1 _5047_ (.A(net559),
    .B(_2164_),
    .C(_2174_),
    .D(_1697_),
    .Y(_1698_));
 sg13g2_nand3_1 _5048_ (.B(net561),
    .C(_2145_),
    .A(_2003_),
    .Y(_1699_));
 sg13g2_nor3_1 _5049_ (.A(_2259_),
    .B(_1652_),
    .C(_1699_),
    .Y(_1700_));
 sg13g2_a21oi_1 _5050_ (.A1(_1657_),
    .A2(_1700_),
    .Y(_1701_),
    .B1(_1629_));
 sg13g2_nand4_1 _5051_ (.B(net560),
    .C(_2113_),
    .A(net561),
    .Y(_1702_),
    .D(_2265_));
 sg13g2_nor3_1 _5052_ (.A(_2075_),
    .B(net548),
    .C(_2259_),
    .Y(_1703_));
 sg13g2_nor3_1 _5053_ (.A(_2146_),
    .B(_2206_),
    .C(_1702_),
    .Y(_1704_));
 sg13g2_nand3_1 _5054_ (.B(_1703_),
    .C(_1704_),
    .A(_1675_),
    .Y(_1705_));
 sg13g2_nand2b_1 _5055_ (.Y(_1706_),
    .B(_1705_),
    .A_N(_1649_));
 sg13g2_and2_1 _5056_ (.A(net543),
    .B(_1626_),
    .X(_1707_));
 sg13g2_nor4_2 _5057_ (.A(net575),
    .B(_2010_),
    .C(_2044_),
    .Y(_1708_),
    .D(_2493_));
 sg13g2_nand3_1 _5058_ (.B(_2313_),
    .C(_1708_),
    .A(net556),
    .Y(_1709_));
 sg13g2_nor4_1 _5059_ (.A(_2042_),
    .B(net553),
    .C(net549),
    .D(_2187_),
    .Y(_1710_));
 sg13g2_nand4_1 _5060_ (.B(_1660_),
    .C(_1708_),
    .A(_2218_),
    .Y(_1711_),
    .D(_1710_));
 sg13g2_nand2_1 _5061_ (.Y(_1712_),
    .A(_1707_),
    .B(_1711_));
 sg13g2_nand4_1 _5062_ (.B(_2021_),
    .C(_2022_),
    .A(_2001_),
    .Y(_1713_),
    .D(_2079_));
 sg13g2_nor4_1 _5063_ (.A(_2010_),
    .B(_2310_),
    .C(_0210_),
    .D(_1713_),
    .Y(_1714_));
 sg13g2_nor2_1 _5064_ (.A(_2044_),
    .B(_2259_),
    .Y(_1715_));
 sg13g2_nand4_1 _5065_ (.B(_1660_),
    .C(_1710_),
    .A(_2081_),
    .Y(_1716_),
    .D(_1715_));
 sg13g2_and2_1 _5066_ (.A(net677),
    .B(_1716_),
    .X(_1717_));
 sg13g2_o21ai_1 _5067_ (.B1(_1712_),
    .Y(_1718_),
    .A1(_1644_),
    .A2(_1698_));
 sg13g2_o21ai_1 _5068_ (.B1(_1706_),
    .Y(_1719_),
    .A1(_1647_),
    .A2(_1714_));
 sg13g2_nor4_2 _5069_ (.A(_1701_),
    .B(_1717_),
    .C(_1718_),
    .Y(_1720_),
    .D(_1719_));
 sg13g2_mux2_2 _5070_ (.A0(_1666_),
    .A1(_1720_),
    .S(net636),
    .X(_1721_));
 sg13g2_a22oi_1 _5071_ (.Y(_1722_),
    .B1(_1721_),
    .B2(\wirecube_top_inst.edge_function_inst.absolute[3] ),
    .A2(_1695_),
    .A1(_1851_));
 sg13g2_nand3_1 _5072_ (.B(_2030_),
    .C(_2281_),
    .A(_2001_),
    .Y(_1723_));
 sg13g2_nor3_1 _5073_ (.A(_2174_),
    .B(_0225_),
    .C(_1723_),
    .Y(_1724_));
 sg13g2_or2_1 _5074_ (.X(_1725_),
    .B(_1724_),
    .A(_1644_));
 sg13g2_nor3_1 _5075_ (.A(_1995_),
    .B(_0161_),
    .C(_1650_),
    .Y(_1726_));
 sg13g2_nand3_1 _5076_ (.B(_1655_),
    .C(_1726_),
    .A(_1653_),
    .Y(_1727_));
 sg13g2_nor4_1 _5077_ (.A(_1995_),
    .B(_2143_),
    .C(_2283_),
    .D(_1702_),
    .Y(_1728_));
 sg13g2_a21oi_1 _5078_ (.A1(_2359_),
    .A2(_1728_),
    .Y(_1729_),
    .B1(_1631_));
 sg13g2_nand3_1 _5079_ (.B(net569),
    .C(_2076_),
    .A(_2021_),
    .Y(_1730_));
 sg13g2_nor3_1 _5080_ (.A(_2162_),
    .B(_0210_),
    .C(_1730_),
    .Y(_1731_));
 sg13g2_nor2_1 _5081_ (.A(_1647_),
    .B(_1731_),
    .Y(_1732_));
 sg13g2_a21oi_1 _5082_ (.A1(net658),
    .A2(_1646_),
    .Y(_1733_),
    .B1(_2296_));
 sg13g2_nor4_1 _5083_ (.A(net641),
    .B(_1729_),
    .C(_1732_),
    .D(_1733_),
    .Y(_1734_));
 sg13g2_nand3_1 _5084_ (.B(_1680_),
    .C(_1708_),
    .A(_0341_),
    .Y(_1735_));
 sg13g2_o21ai_1 _5085_ (.B1(_1626_),
    .Y(_1736_),
    .A1(net546),
    .A2(_1735_));
 sg13g2_nand3_1 _5086_ (.B(_2280_),
    .C(_1715_),
    .A(_2026_),
    .Y(_1737_));
 sg13g2_o21ai_1 _5087_ (.B1(net677),
    .Y(_1738_),
    .A1(_1684_),
    .A2(_1737_));
 sg13g2_nand3_1 _5088_ (.B(_1736_),
    .C(_1738_),
    .A(_1734_),
    .Y(_1739_));
 sg13g2_a21oi_1 _5089_ (.A1(_1630_),
    .A2(_1727_),
    .Y(_1740_),
    .B1(_1739_));
 sg13g2_a22oi_1 _5090_ (.Y(_1741_),
    .B1(_1725_),
    .B2(_1740_),
    .A2(_1693_),
    .A1(net641));
 sg13g2_xnor2_1 _5091_ (.Y(_1742_),
    .A(_0065_),
    .B(_1741_));
 sg13g2_nand2_1 _5092_ (.Y(_1743_),
    .A(net641),
    .B(_1720_));
 sg13g2_nand2b_1 _5093_ (.Y(_1744_),
    .B(_2491_),
    .A_N(_2352_));
 sg13g2_nand2_1 _5094_ (.Y(_1745_),
    .A(_2024_),
    .B(_0258_));
 sg13g2_nor4_1 _5095_ (.A(_2178_),
    .B(_2185_),
    .C(_2210_),
    .D(_0210_),
    .Y(_1746_));
 sg13g2_nor4_2 _5096_ (.A(net563),
    .B(_2217_),
    .C(_1744_),
    .Y(_1747_),
    .D(_1745_));
 sg13g2_a21oi_2 _5097_ (.B1(_1644_),
    .Y(_1748_),
    .A2(_1747_),
    .A1(_1746_));
 sg13g2_or2_1 _5098_ (.X(_1749_),
    .B(_1655_),
    .A(net658));
 sg13g2_nand3_1 _5099_ (.B(_1651_),
    .C(_1749_),
    .A(_0427_),
    .Y(_1750_));
 sg13g2_nand3_1 _5100_ (.B(_1657_),
    .C(_1750_),
    .A(_1630_),
    .Y(_1751_));
 sg13g2_a21oi_1 _5101_ (.A1(_2296_),
    .A2(_1655_),
    .Y(_1752_),
    .B1(net662));
 sg13g2_nor4_1 _5102_ (.A(net562),
    .B(_2141_),
    .C(net549),
    .D(_2314_),
    .Y(_1753_));
 sg13g2_nand3_1 _5103_ (.B(_0164_),
    .C(_1753_),
    .A(_2394_),
    .Y(_1754_));
 sg13g2_o21ai_1 _5104_ (.B1(net677),
    .Y(_1755_),
    .A1(_2492_),
    .A2(_1754_));
 sg13g2_nor3_1 _5105_ (.A(_2029_),
    .B(_2112_),
    .C(_2163_),
    .Y(_1756_));
 sg13g2_a21oi_1 _5106_ (.A1(_1676_),
    .A2(_1756_),
    .Y(_1757_),
    .B1(_1649_));
 sg13g2_or4_1 _5107_ (.A(_2206_),
    .B(_2332_),
    .C(_1709_),
    .D(_1745_),
    .X(_1758_));
 sg13g2_nor3_1 _5108_ (.A(net641),
    .B(_1752_),
    .C(_1757_),
    .Y(_1759_));
 sg13g2_nor4_1 _5109_ (.A(_2046_),
    .B(net562),
    .C(_0210_),
    .D(_1687_),
    .Y(_1760_));
 sg13g2_and4_1 _5110_ (.A(_2247_),
    .B(_2309_),
    .C(_0160_),
    .D(_1760_),
    .X(_1761_));
 sg13g2_a21oi_1 _5111_ (.A1(_2083_),
    .A2(_1761_),
    .Y(_1762_),
    .B1(_1646_));
 sg13g2_nor4_1 _5112_ (.A(net558),
    .B(net552),
    .C(net549),
    .D(_2493_),
    .Y(_1763_));
 sg13g2_nand4_1 _5113_ (.B(_1635_),
    .C(_1760_),
    .A(_2313_),
    .Y(_1764_),
    .D(_1763_));
 sg13g2_a221oi_1 _5114_ (.B2(_1645_),
    .C1(_1762_),
    .B1(_1764_),
    .A1(_1707_),
    .Y(_1765_),
    .A2(_1758_));
 sg13g2_nand4_1 _5115_ (.B(_1755_),
    .C(_1759_),
    .A(_1751_),
    .Y(_1766_),
    .D(_1765_));
 sg13g2_o21ai_1 _5116_ (.B1(_1743_),
    .Y(_1767_),
    .A1(_1748_),
    .A2(_1766_));
 sg13g2_nor3_1 _5117_ (.A(\wirecube_top_inst.edge_function_inst.absolute[1] ),
    .B(_1742_),
    .C(_1767_),
    .Y(_1768_));
 sg13g2_or2_1 _5118_ (.X(_1769_),
    .B(_1721_),
    .A(\wirecube_top_inst.edge_function_inst.absolute[3] ));
 sg13g2_nand2b_1 _5119_ (.Y(_1770_),
    .B(_1741_),
    .A_N(\wirecube_top_inst.edge_function_inst.absolute[2] ));
 sg13g2_nand2_1 _5120_ (.Y(_1771_),
    .A(_1769_),
    .B(_1770_));
 sg13g2_o21ai_1 _5121_ (.B1(_1722_),
    .Y(_1772_),
    .A1(_1768_),
    .A2(_1771_));
 sg13g2_a21oi_1 _5122_ (.A1(_1696_),
    .A2(_1772_),
    .Y(_1773_),
    .B1(_1669_));
 sg13g2_o21ai_1 _5123_ (.B1(_1643_),
    .Y(_1774_),
    .A1(_1668_),
    .A2(_1773_));
 sg13g2_nand2b_1 _5124_ (.Y(_1775_),
    .B(_1641_),
    .A_N(\wirecube_top_inst.edge_function_inst.absolute[6] ));
 sg13g2_o21ai_1 _5125_ (.B1(_1774_),
    .Y(_1776_),
    .A1(\wirecube_top_inst.edge_function_inst.absolute[7] ),
    .A2(_1775_));
 sg13g2_or4_1 _5126_ (.A(\wirecube_top_inst.edge_function_inst.absolute[11] ),
    .B(\wirecube_top_inst.edge_function_inst.absolute[10] ),
    .C(\wirecube_top_inst.edge_function_inst.absolute[9] ),
    .D(\wirecube_top_inst.edge_function_inst.absolute[8] ),
    .X(_1777_));
 sg13g2_nor3_2 _5127_ (.A(\wirecube_top_inst.edge_function_inst.absolute[12] ),
    .B(\wirecube_top_inst.edge_function_inst.absolute[13] ),
    .C(_1777_),
    .Y(_1778_));
 sg13g2_and2_1 _5128_ (.A(\wirecube_top_inst.edge_function_inst.visible_2 ),
    .B(_1778_),
    .X(_1779_));
 sg13g2_xnor2_1 _5129_ (.Y(_1780_),
    .A(_0067_),
    .B(_1767_));
 sg13g2_nand4_1 _5130_ (.B(_1643_),
    .C(_1696_),
    .A(_0066_),
    .Y(_1781_),
    .D(_1775_));
 sg13g2_nor3_1 _5131_ (.A(_1669_),
    .B(_1742_),
    .C(_1781_),
    .Y(_1782_));
 sg13g2_nand4_1 _5132_ (.B(_1769_),
    .C(_1780_),
    .A(_1722_),
    .Y(_1783_),
    .D(_1782_));
 sg13g2_nand3_1 _5133_ (.B(_1779_),
    .C(_1783_),
    .A(_1776_),
    .Y(_1784_));
 sg13g2_a22oi_1 _5134_ (.Y(_0142_),
    .B1(_1625_),
    .B2(_1784_),
    .A2(_1624_),
    .A1(_1852_));
 sg13g2_nor2_1 _5135_ (.A(net138),
    .B(_1623_),
    .Y(_1785_));
 sg13g2_nor3_1 _5136_ (.A(\wirecube_top_inst.linecounter_h[2] ),
    .B(net91),
    .C(_1522_),
    .Y(_1786_));
 sg13g2_and2_1 _5137_ (.A(\wirecube_top_inst.edge_function_inst.absolute[3] ),
    .B(_1695_),
    .X(_1787_));
 sg13g2_nor3_2 _5138_ (.A(\wirecube_top_inst.edge_function_inst.absolute[4] ),
    .B(net642),
    .C(_1666_),
    .Y(_1788_));
 sg13g2_xor2_1 _5139_ (.B(_1641_),
    .A(\wirecube_top_inst.edge_function_inst.absolute[5] ),
    .X(_1789_));
 sg13g2_inv_1 _5140_ (.Y(_1790_),
    .A(_1789_));
 sg13g2_nor2b_1 _5141_ (.A(_1667_),
    .B_N(\wirecube_top_inst.edge_function_inst.absolute[4] ),
    .Y(_1791_));
 sg13g2_nor4_1 _5142_ (.A(_1787_),
    .B(_1788_),
    .C(_1789_),
    .D(_1791_),
    .Y(_1792_));
 sg13g2_or4_1 _5143_ (.A(_1787_),
    .B(_1788_),
    .C(_1789_),
    .D(_1791_),
    .X(_1794_));
 sg13g2_xor2_1 _5144_ (.B(_1721_),
    .A(_0065_),
    .X(_1795_));
 sg13g2_xnor2_1 _5145_ (.Y(_1796_),
    .A(_0067_),
    .B(_1741_));
 sg13g2_a21o_1 _5146_ (.A2(_1767_),
    .A1(\wirecube_top_inst.edge_function_inst.absolute[0] ),
    .B1(_1796_),
    .X(_1797_));
 sg13g2_nand2b_1 _5147_ (.Y(_1798_),
    .B(_1741_),
    .A_N(\wirecube_top_inst.edge_function_inst.absolute[1] ));
 sg13g2_a21oi_1 _5148_ (.A1(_1797_),
    .A2(_1798_),
    .Y(_1799_),
    .B1(_1795_));
 sg13g2_or2_1 _5149_ (.X(_1800_),
    .B(_1695_),
    .A(\wirecube_top_inst.edge_function_inst.absolute[3] ));
 sg13g2_o21ai_1 _5150_ (.B1(_1800_),
    .Y(_1801_),
    .A1(\wirecube_top_inst.edge_function_inst.absolute[2] ),
    .A2(_1721_));
 sg13g2_o21ai_1 _5151_ (.B1(_1792_),
    .Y(_1802_),
    .A1(_1799_),
    .A2(_1801_));
 sg13g2_a22oi_1 _5152_ (.Y(_1803_),
    .B1(_1788_),
    .B2(_1790_),
    .A2(_1641_),
    .A1(_0063_));
 sg13g2_nand2_1 _5153_ (.Y(_1805_),
    .A(_1802_),
    .B(_1803_));
 sg13g2_xnor2_1 _5154_ (.Y(_1806_),
    .A(_0066_),
    .B(_1767_));
 sg13g2_nand3_1 _5155_ (.B(_1800_),
    .C(_1806_),
    .A(_1778_),
    .Y(_1807_));
 sg13g2_nor4_1 _5156_ (.A(_1794_),
    .B(_1795_),
    .C(_1796_),
    .D(_1807_),
    .Y(_1808_));
 sg13g2_nor3_1 _5157_ (.A(\wirecube_top_inst.edge_function_inst.absolute[6] ),
    .B(\wirecube_top_inst.edge_function_inst.absolute[7] ),
    .C(_1808_),
    .Y(_1809_));
 sg13g2_nand3_1 _5158_ (.B(_1805_),
    .C(_1809_),
    .A(_1779_),
    .Y(_1810_));
 sg13g2_a21oi_1 _5159_ (.A1(_1786_),
    .A2(_1810_),
    .Y(_0143_),
    .B1(net139));
 sg13g2_o21ai_1 _5160_ (.B1(\wirecube_top_inst.edge_function_inst.pixel_x_i[0] ),
    .Y(_1811_),
    .A1(net655),
    .A2(net646));
 sg13g2_nor2_2 _5161_ (.A(_2151_),
    .B(net646),
    .Y(_1812_));
 sg13g2_mux2_1 _5162_ (.A0(_1812_),
    .A1(_1513_),
    .S(net186),
    .X(_0144_));
 sg13g2_and2_1 _5163_ (.A(\wirecube_top_inst.edge_function_inst.pixel_x_i[1] ),
    .B(\wirecube_top_inst.edge_function_inst.pixel_x_i[0] ),
    .X(_1814_));
 sg13g2_a221oi_1 _5164_ (.B2(net655),
    .C1(net646),
    .B1(_1814_),
    .A1(_1850_),
    .Y(_0145_),
    .A2(_1811_));
 sg13g2_xnor2_1 _5165_ (.Y(_1815_),
    .A(net181),
    .B(_1814_));
 sg13g2_a22oi_1 _5166_ (.Y(_1816_),
    .B1(_1812_),
    .B2(_1815_),
    .A2(_1513_),
    .A1(net681));
 sg13g2_inv_1 _5167_ (.Y(_0146_),
    .A(_1816_));
 sg13g2_and2_1 _5168_ (.A(net681),
    .B(_1814_),
    .X(_1817_));
 sg13g2_a21oi_1 _5169_ (.A1(net655),
    .A2(_1817_),
    .Y(_1818_),
    .B1(net194));
 sg13g2_nand2_1 _5170_ (.Y(_1819_),
    .A(\wirecube_top_inst.edge_function_inst.pixel_x_i[3] ),
    .B(_1817_));
 sg13g2_nor2_1 _5171_ (.A(_2151_),
    .B(_1819_),
    .Y(_1820_));
 sg13g2_nor3_1 _5172_ (.A(net646),
    .B(_1818_),
    .C(_1820_),
    .Y(_0147_));
 sg13g2_xor2_1 _5173_ (.B(_1819_),
    .A(net183),
    .X(_1822_));
 sg13g2_a22oi_1 _5174_ (.Y(_1823_),
    .B1(_1812_),
    .B2(_1822_),
    .A2(_1513_),
    .A1(\wirecube_top_inst.edge_function_inst.pixel_x_i[4] ));
 sg13g2_inv_1 _5175_ (.Y(_0148_),
    .A(net184));
 sg13g2_a21oi_1 _5176_ (.A1(\wirecube_top_inst.edge_function_inst.pixel_x_i[4] ),
    .A2(_1820_),
    .Y(_1824_),
    .B1(net187));
 sg13g2_nand4_1 _5177_ (.B(\wirecube_top_inst.edge_function_inst.pixel_x_i[4] ),
    .C(\wirecube_top_inst.edge_function_inst.pixel_x_i[3] ),
    .A(\wirecube_top_inst.edge_function_inst.pixel_x_i[5] ),
    .Y(_1825_),
    .D(_1817_));
 sg13g2_nor2_1 _5178_ (.A(_2151_),
    .B(_1825_),
    .Y(_1826_));
 sg13g2_nor3_1 _5179_ (.A(net646),
    .B(net188),
    .C(_1826_),
    .Y(_0149_));
 sg13g2_xor2_1 _5180_ (.B(_1825_),
    .A(_0061_),
    .X(_1827_));
 sg13g2_a22oi_1 _5181_ (.Y(_1828_),
    .B1(_1812_),
    .B2(_1827_),
    .A2(_1513_),
    .A1(net133));
 sg13g2_inv_1 _5182_ (.Y(_0150_),
    .A(net134));
 sg13g2_or4_1 _5183_ (.A(\wirecube_top_inst.linecounter_h[1] ),
    .B(\wirecube_top_inst.linecounter_h[0] ),
    .C(\wirecube_top_inst.linecounter_h[3] ),
    .D(\wirecube_top_inst.linecounter_h[2] ),
    .X(_1830_));
 sg13g2_o21ai_1 _5184_ (.B1(net674),
    .Y(_1831_),
    .A1(\wirecube_top_inst.linecounter_h[2] ),
    .A2(_1522_));
 sg13g2_o21ai_1 _5185_ (.B1(net102),
    .Y(_1832_),
    .A1(_1830_),
    .A2(_1831_));
 sg13g2_o21ai_1 _5186_ (.B1(net103),
    .Y(_0151_),
    .A1(_1784_),
    .A2(_1831_));
 sg13g2_nand2_1 _5187_ (.Y(_1833_),
    .A(net91),
    .B(_1830_));
 sg13g2_o21ai_1 _5188_ (.B1(_1833_),
    .Y(_0152_),
    .A1(_1623_),
    .A2(_1810_));
 sg13g2_dfrbp_1 _5189_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net664),
    .D(net132),
    .Q_N(_0059_),
    .Q(\wirecube_top_inst.edge_function_inst.pixel_y_i[0] ));
 sg13g2_dfrbp_1 _5190_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net664),
    .D(_0109_),
    .Q_N(_2568_),
    .Q(\wirecube_top_inst.edge_function_inst.pixel_y_i[1] ));
 sg13g2_dfrbp_1 _5191_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net664),
    .D(_0110_),
    .Q_N(_0053_),
    .Q(\wirecube_top_inst.edge_function_inst.pixel_y_i[2] ));
 sg13g2_dfrbp_1 _5192_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net674),
    .D(net180),
    .Q_N(_2567_),
    .Q(\wirecube_top_inst.edge_function_inst.pixel_y_i[3] ));
 sg13g2_dfrbp_1 _5193_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net674),
    .D(_0112_),
    .Q_N(_0052_),
    .Q(\wirecube_top_inst.edge_function_inst.pixel_y_i[4] ));
 sg13g2_dfrbp_1 _5194_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net674),
    .D(_0113_),
    .Q_N(_0054_),
    .Q(\wirecube_top_inst.edge_function_inst.pixel_y_i[5] ));
 sg13g2_dfrbp_1 _5195_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net676),
    .D(_0114_),
    .Q_N(_0051_),
    .Q(\wirecube_top_inst.edge_function_inst.pixel_y_i[6] ));
 sg13g2_dfrbp_1 _5196_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net672),
    .D(net96),
    .Q_N(_2569_),
    .Q(\wirecube_top_inst.linecounter_h[0] ));
 sg13g2_dfrbp_1 _5197_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net672),
    .D(_0001_),
    .Q_N(_2570_),
    .Q(\wirecube_top_inst.linecounter_h[1] ));
 sg13g2_dfrbp_1 _5198_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net672),
    .D(net146),
    .Q_N(_2571_),
    .Q(\wirecube_top_inst.linecounter_h[2] ));
 sg13g2_dfrbp_1 _5199_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net672),
    .D(net127),
    .Q_N(_2566_),
    .Q(\wirecube_top_inst.linecounter_h[3] ));
 sg13g2_dfrbp_1 _5200_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net666),
    .D(_0115_),
    .Q_N(_2565_),
    .Q(\wirecube_top_inst.subcounter_v[0] ));
 sg13g2_dfrbp_1 _5201_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net666),
    .D(net110),
    .Q_N(_2564_),
    .Q(\wirecube_top_inst.subcounter_v[1] ));
 sg13g2_dfrbp_1 _5202_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net666),
    .D(net98),
    .Q_N(_0050_),
    .Q(\wirecube_top_inst.subcounter_v[2] ));
 sg13g2_dfrbp_1 _5203_ (.CLK(net73),
    .RESET_B(net25),
    .D(net1),
    .Q_N(_2572_),
    .Q(rst_n_sync));
 sg13g2_dfrbp_1 _5204_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net670),
    .D(net118),
    .Q_N(_2573_),
    .Q(\wirecube_top_inst.delay_inst_vsync.pipe[0] ));
 sg13g2_dfrbp_1 _5205_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net671),
    .D(net76),
    .Q_N(_2574_),
    .Q(vsync));
 sg13g2_dfrbp_1 _5206_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net667),
    .D(net142),
    .Q_N(_2575_),
    .Q(\wirecube_top_inst.delay_inst_hsync.pipe[0] ));
 sg13g2_dfrbp_1 _5207_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net668),
    .D(net74),
    .Q_N(_2576_),
    .Q(hsync));
 sg13g2_dfrbp_1 _5208_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net26),
    .D(_0042_),
    .Q_N(_2577_),
    .Q(\wirecube_top_inst.edge_function_inst.visible ));
 sg13g2_dfrbp_1 _5209_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net27),
    .D(_0014_),
    .Q_N(_0066_),
    .Q(\wirecube_top_inst.edge_function_inst.absolute[0] ));
 sg13g2_dfrbp_1 _5210_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net28),
    .D(_0019_),
    .Q_N(_0067_),
    .Q(\wirecube_top_inst.edge_function_inst.absolute[1] ));
 sg13g2_dfrbp_1 _5211_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net29),
    .D(_0020_),
    .Q_N(_0065_),
    .Q(\wirecube_top_inst.edge_function_inst.absolute[2] ));
 sg13g2_dfrbp_1 _5212_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net30),
    .D(_0021_),
    .Q_N(_2578_),
    .Q(\wirecube_top_inst.edge_function_inst.absolute[3] ));
 sg13g2_dfrbp_1 _5213_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net31),
    .D(_0022_),
    .Q_N(_0064_),
    .Q(\wirecube_top_inst.edge_function_inst.absolute[4] ));
 sg13g2_dfrbp_1 _5214_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net32),
    .D(_0023_),
    .Q_N(_0063_),
    .Q(\wirecube_top_inst.edge_function_inst.absolute[5] ));
 sg13g2_dfrbp_1 _5215_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net33),
    .D(_0024_),
    .Q_N(_2579_),
    .Q(\wirecube_top_inst.edge_function_inst.absolute[6] ));
 sg13g2_dfrbp_1 _5216_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net34),
    .D(_0025_),
    .Q_N(_2580_),
    .Q(\wirecube_top_inst.edge_function_inst.absolute[7] ));
 sg13g2_dfrbp_1 _5217_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net35),
    .D(_0026_),
    .Q_N(_2581_),
    .Q(\wirecube_top_inst.edge_function_inst.absolute[8] ));
 sg13g2_dfrbp_1 _5218_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net36),
    .D(_0027_),
    .Q_N(_2582_),
    .Q(\wirecube_top_inst.edge_function_inst.absolute[9] ));
 sg13g2_dfrbp_1 _5219_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net37),
    .D(_0015_),
    .Q_N(_2583_),
    .Q(\wirecube_top_inst.edge_function_inst.absolute[10] ));
 sg13g2_dfrbp_1 _5220_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net38),
    .D(_0016_),
    .Q_N(_2584_),
    .Q(\wirecube_top_inst.edge_function_inst.absolute[11] ));
 sg13g2_dfrbp_1 _5221_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net39),
    .D(_0017_),
    .Q_N(_2585_),
    .Q(\wirecube_top_inst.edge_function_inst.absolute[12] ));
 sg13g2_dfrbp_1 _5222_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net40),
    .D(_0018_),
    .Q_N(_2586_),
    .Q(\wirecube_top_inst.edge_function_inst.absolute[13] ));
 sg13g2_dfrbp_1 _5223_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net41),
    .D(net75),
    .Q_N(_2587_),
    .Q(\wirecube_top_inst.edge_function_inst.visible_2 ));
 sg13g2_dfrbp_1 _5224_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net42),
    .D(_0028_),
    .Q_N(_2588_),
    .Q(\wirecube_top_inst.edge_function_inst.term0[0] ));
 sg13g2_dfrbp_1 _5225_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net43),
    .D(_0029_),
    .Q_N(_2589_),
    .Q(\wirecube_top_inst.edge_function_inst.term0[1] ));
 sg13g2_dfrbp_1 _5226_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net44),
    .D(_0030_),
    .Q_N(_2590_),
    .Q(\wirecube_top_inst.edge_function_inst.term0[2] ));
 sg13g2_dfrbp_1 _5227_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net45),
    .D(_0031_),
    .Q_N(_2591_),
    .Q(\wirecube_top_inst.edge_function_inst.term0[3] ));
 sg13g2_dfrbp_1 _5228_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net46),
    .D(_0032_),
    .Q_N(_2592_),
    .Q(\wirecube_top_inst.edge_function_inst.term0[4] ));
 sg13g2_dfrbp_1 _5229_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net47),
    .D(_0033_),
    .Q_N(_2593_),
    .Q(\wirecube_top_inst.edge_function_inst.term0[5] ));
 sg13g2_dfrbp_1 _5230_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net48),
    .D(_0034_),
    .Q_N(_2594_),
    .Q(\wirecube_top_inst.edge_function_inst.term0[6] ));
 sg13g2_dfrbp_1 _5231_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net49),
    .D(_0074_),
    .Q_N(_2595_),
    .Q(\wirecube_top_inst.edge_function_inst.term1[0] ));
 sg13g2_dfrbp_1 _5232_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net50),
    .D(_0075_),
    .Q_N(_2596_),
    .Q(\wirecube_top_inst.edge_function_inst.term1[1] ));
 sg13g2_dfrbp_1 _5233_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net51),
    .D(_0076_),
    .Q_N(_2597_),
    .Q(\wirecube_top_inst.edge_function_inst.term1[2] ));
 sg13g2_dfrbp_1 _5234_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net52),
    .D(_0077_),
    .Q_N(_2598_),
    .Q(\wirecube_top_inst.edge_function_inst.term1[3] ));
 sg13g2_dfrbp_1 _5235_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net53),
    .D(_0078_),
    .Q_N(_2599_),
    .Q(\wirecube_top_inst.edge_function_inst.term1[4] ));
 sg13g2_dfrbp_1 _5236_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net54),
    .D(_0079_),
    .Q_N(_2600_),
    .Q(\wirecube_top_inst.edge_function_inst.term1[5] ));
 sg13g2_dfrbp_1 _5237_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net55),
    .D(_0080_),
    .Q_N(_2601_),
    .Q(\wirecube_top_inst.edge_function_inst.term1[6] ));
 sg13g2_dfrbp_1 _5238_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net56),
    .D(_0035_),
    .Q_N(_2602_),
    .Q(\wirecube_top_inst.edge_function_inst.term2[0] ));
 sg13g2_dfrbp_1 _5239_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net57),
    .D(_0036_),
    .Q_N(_2603_),
    .Q(\wirecube_top_inst.edge_function_inst.term2[1] ));
 sg13g2_dfrbp_1 _5240_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net58),
    .D(_0037_),
    .Q_N(_2604_),
    .Q(\wirecube_top_inst.edge_function_inst.term2[2] ));
 sg13g2_dfrbp_1 _5241_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net59),
    .D(_0038_),
    .Q_N(_2605_),
    .Q(\wirecube_top_inst.edge_function_inst.term2[3] ));
 sg13g2_dfrbp_1 _5242_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net60),
    .D(_0039_),
    .Q_N(_2606_),
    .Q(\wirecube_top_inst.edge_function_inst.term2[4] ));
 sg13g2_dfrbp_1 _5243_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net61),
    .D(_0040_),
    .Q_N(_2607_),
    .Q(\wirecube_top_inst.edge_function_inst.term2[5] ));
 sg13g2_dfrbp_1 _5244_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net62),
    .D(_0041_),
    .Q_N(_2608_),
    .Q(\wirecube_top_inst.edge_function_inst.term2[6] ));
 sg13g2_dfrbp_1 _5245_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net63),
    .D(_0081_),
    .Q_N(_2609_),
    .Q(\wirecube_top_inst.edge_function_inst.term3[0] ));
 sg13g2_dfrbp_1 _5246_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net64),
    .D(_0082_),
    .Q_N(_2610_),
    .Q(\wirecube_top_inst.edge_function_inst.term3[1] ));
 sg13g2_dfrbp_1 _5247_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net65),
    .D(_0083_),
    .Q_N(_2611_),
    .Q(\wirecube_top_inst.edge_function_inst.term3[2] ));
 sg13g2_dfrbp_1 _5248_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net66),
    .D(_0084_),
    .Q_N(_2612_),
    .Q(\wirecube_top_inst.edge_function_inst.term3[3] ));
 sg13g2_dfrbp_1 _5249_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net67),
    .D(_0085_),
    .Q_N(_2613_),
    .Q(\wirecube_top_inst.edge_function_inst.term3[4] ));
 sg13g2_dfrbp_1 _5250_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net70),
    .D(_0086_),
    .Q_N(_2614_),
    .Q(\wirecube_top_inst.edge_function_inst.term3[5] ));
 sg13g2_dfrbp_1 _5251_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net71),
    .D(_0087_),
    .Q_N(_2563_),
    .Q(\wirecube_top_inst.edge_function_inst.term3[6] ));
 sg13g2_dfrbp_1 _5252_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net670),
    .D(_0118_),
    .Q_N(\wirecube_top_inst.counter_v[0] ),
    .Q(_0089_));
 sg13g2_dfrbp_1 _5253_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net670),
    .D(net82),
    .Q_N(\wirecube_top_inst.counter_v[1] ),
    .Q(_0090_));
 sg13g2_dfrbp_1 _5254_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net670),
    .D(_0120_),
    .Q_N(_2562_),
    .Q(\wirecube_top_inst.counter_v[2] ));
 sg13g2_dfrbp_1 _5255_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net670),
    .D(_0121_),
    .Q_N(_2561_),
    .Q(\wirecube_top_inst.counter_v[3] ));
 sg13g2_dfrbp_1 _5256_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net666),
    .D(net88),
    .Q_N(\wirecube_top_inst.counter_v[4] ),
    .Q(_0091_));
 sg13g2_dfrbp_1 _5257_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net670),
    .D(_0123_),
    .Q_N(_2560_),
    .Q(\wirecube_top_inst.counter_v[5] ));
 sg13g2_dfrbp_1 _5258_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net667),
    .D(net86),
    .Q_N(\wirecube_top_inst.counter_v[6] ),
    .Q(_0092_));
 sg13g2_dfrbp_1 _5259_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net668),
    .D(net94),
    .Q_N(\wirecube_top_inst.counter_v[7] ),
    .Q(_0093_));
 sg13g2_dfrbp_1 _5260_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net668),
    .D(net84),
    .Q_N(\wirecube_top_inst.counter_v[8] ),
    .Q(_0094_));
 sg13g2_dfrbp_1 _5261_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net667),
    .D(net80),
    .Q_N(\wirecube_top_inst.counter_v[9] ),
    .Q(_0095_));
 sg13g2_dfrbp_1 _5262_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net668),
    .D(net100),
    .Q_N(\wirecube_top_inst.counter_v[10] ),
    .Q(_0096_));
 sg13g2_dfrbp_1 _5263_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net670),
    .D(net78),
    .Q_N(_0088_),
    .Q(\wirecube_top_inst.frame_cnt[0] ));
 sg13g2_dfrbp_1 _5264_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net671),
    .D(_0130_),
    .Q_N(_2559_),
    .Q(\wirecube_top_inst.frame_cnt[1] ));
 sg13g2_dfrbp_1 _5265_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net665),
    .D(_0131_),
    .Q_N(_0073_),
    .Q(\wirecube_top_inst.frame_cnt[2] ));
 sg13g2_dfrbp_1 _5266_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net664),
    .D(net161),
    .Q_N(_0070_),
    .Q(\wirecube_top_inst.frame_cnt[3] ));
 sg13g2_dfrbp_1 _5267_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net664),
    .D(net178),
    .Q_N(_0072_),
    .Q(\wirecube_top_inst.frame_cnt[4] ));
 sg13g2_dfrbp_1 _5268_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net665),
    .D(net158),
    .Q_N(_0069_),
    .Q(\wirecube_top_inst.frame_cnt[5] ));
 sg13g2_dfrbp_1 _5269_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net674),
    .D(_0135_),
    .Q_N(_0071_),
    .Q(\wirecube_top_inst.frame_cnt[6] ));
 sg13g2_dfrbp_1 _5270_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net673),
    .D(_0136_),
    .Q_N(_0060_),
    .Q(\wirecube_top_inst.frame_cnt[7] ));
 sg13g2_dfrbp_1 _5271_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net672),
    .D(_0137_),
    .Q_N(_2558_),
    .Q(\wirecube_top_inst.cur_state_background[0] ));
 sg13g2_dfrbp_1 _5272_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net672),
    .D(_0138_),
    .Q_N(_2557_),
    .Q(\wirecube_top_inst.cur_state_background[1] ));
 sg13g2_dfrbp_1 _5273_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net673),
    .D(_0139_),
    .Q_N(_2556_),
    .Q(\wirecube_top_inst.cur_state_background[2] ));
 sg13g2_dfrbp_1 _5274_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net672),
    .D(net198),
    .Q_N(_2555_),
    .Q(\wirecube_top_inst.cur_state_background[3] ));
 sg13g2_dfrbp_1 _5275_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net672),
    .D(_0141_),
    .Q_N(_0062_),
    .Q(\wirecube_top_inst.frame_cnt[12] ));
 sg13g2_dfrbp_1 _5276_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net671),
    .D(_0043_),
    .Q_N(_2615_),
    .Q(\wirecube_top_inst.counter_h[0] ));
 sg13g2_dfrbp_1 _5277_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net669),
    .D(_0044_),
    .Q_N(_2616_),
    .Q(\wirecube_top_inst.counter_h[1] ));
 sg13g2_dfrbp_1 _5278_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net669),
    .D(_0045_),
    .Q_N(_2617_),
    .Q(\wirecube_top_inst.counter_h[2] ));
 sg13g2_dfrbp_1 _5279_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net666),
    .D(_0046_),
    .Q_N(_2618_),
    .Q(\wirecube_top_inst.counter_h[3] ));
 sg13g2_dfrbp_1 _5280_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net666),
    .D(_0047_),
    .Q_N(_2619_),
    .Q(\wirecube_top_inst.counter_h[4] ));
 sg13g2_dfrbp_1 _5281_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net666),
    .D(_0048_),
    .Q_N(_0068_),
    .Q(\wirecube_top_inst.counter_h[5] ));
 sg13g2_dfrbp_1 _5282_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net666),
    .D(_0103_),
    .Q_N(\wirecube_top_inst.counter_h[6] ),
    .Q(_0097_));
 sg13g2_dfrbp_1 _5283_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net667),
    .D(_0104_),
    .Q_N(\wirecube_top_inst.counter_h[7] ),
    .Q(_0098_));
 sg13g2_dfrbp_1 _5284_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net667),
    .D(net121),
    .Q_N(_2554_),
    .Q(\wirecube_top_inst.counter_h[8] ));
 sg13g2_dfrbp_1 _5285_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net667),
    .D(_0105_),
    .Q_N(\wirecube_top_inst.counter_h[9] ),
    .Q(_0099_));
 sg13g2_dfrbp_1 _5286_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net667),
    .D(_0106_),
    .Q_N(\wirecube_top_inst.counter_h[10] ),
    .Q(_0100_));
 sg13g2_dfrbp_1 _5287_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net667),
    .D(_0107_),
    .Q_N(\wirecube_top_inst.timing_hor.counter[11] ),
    .Q(_0101_));
 sg13g2_dfrbp_1 _5288_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net68),
    .D(net106),
    .Q_N(_2553_),
    .Q(\wirecube_top_inst.final_pixel2 ));
 sg13g2_dfrbp_1 _5289_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net674),
    .D(net140),
    .Q_N(_2552_),
    .Q(\wirecube_top_inst.final_pixel ));
 sg13g2_dfrbp_1 _5290_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net676),
    .D(_0144_),
    .Q_N(_0058_),
    .Q(\wirecube_top_inst.edge_function_inst.pixel_x_i[0] ));
 sg13g2_dfrbp_1 _5291_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net676),
    .D(net169),
    .Q_N(_0057_),
    .Q(\wirecube_top_inst.edge_function_inst.pixel_x_i[1] ));
 sg13g2_dfrbp_1 _5292_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net676),
    .D(_0146_),
    .Q_N(_0056_),
    .Q(\wirecube_top_inst.edge_function_inst.pixel_x_i[2] ));
 sg13g2_dfrbp_1 _5293_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net676),
    .D(_0147_),
    .Q_N(_2551_),
    .Q(\wirecube_top_inst.edge_function_inst.pixel_x_i[3] ));
 sg13g2_dfrbp_1 _5294_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net676),
    .D(_0148_),
    .Q_N(_0055_),
    .Q(\wirecube_top_inst.edge_function_inst.pixel_x_i[4] ));
 sg13g2_dfrbp_1 _5295_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net676),
    .D(_0149_),
    .Q_N(_2550_),
    .Q(\wirecube_top_inst.edge_function_inst.pixel_x_i[5] ));
 sg13g2_dfrbp_1 _5296_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net676),
    .D(_0150_),
    .Q_N(_0061_),
    .Q(\wirecube_top_inst.edge_function_inst.pixel_x_i[6] ));
 sg13g2_dfrbp_1 _5297_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net69),
    .D(net104),
    .Q_N(_2549_),
    .Q(\wirecube_top_inst.any_line_set2 ));
 sg13g2_dfrbp_1 _5298_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net674),
    .D(net92),
    .Q_N(_2620_),
    .Q(\wirecube_top_inst.any_line_set ));
 sg13g2_dfrbp_1 _5299_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net664),
    .D(net148),
    .Q_N(_2621_),
    .Q(\wirecube_top_inst.line_rom_inst.line_i[0] ));
 sg13g2_dfrbp_1 _5300_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net664),
    .D(_0011_),
    .Q_N(_2622_),
    .Q(\wirecube_top_inst.line_rom_inst.line_i[1] ));
 sg13g2_dfrbp_1 _5301_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net664),
    .D(_0012_),
    .Q_N(_2623_),
    .Q(\wirecube_top_inst.line_rom_inst.line_i[2] ));
 sg13g2_dfrbp_1 _5302_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net665),
    .D(_0013_),
    .Q_N(_2624_),
    .Q(\wirecube_top_inst.line_rom_inst.line_i[3] ));
 sg13g2_dfrbp_1 _5303_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net673),
    .D(_0004_),
    .Q_N(_2625_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _5304_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net671),
    .D(_0005_),
    .Q_N(_2626_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _5305_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net673),
    .D(_0006_),
    .Q_N(_2627_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _5306_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net673),
    .D(_0007_),
    .Q_N(_2628_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _5307_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net673),
    .D(_0008_),
    .Q_N(_2629_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _5308_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net670),
    .D(_0009_),
    .Q_N(_2548_),
    .Q(uo_out[0]));
 sg13g2_tiehi _5208__26 (.L_HI(net26));
 sg13g2_tiehi _5209__27 (.L_HI(net27));
 sg13g2_tiehi _5210__28 (.L_HI(net28));
 sg13g2_tiehi _5211__29 (.L_HI(net29));
 sg13g2_tiehi _5212__30 (.L_HI(net30));
 sg13g2_tiehi _5213__31 (.L_HI(net31));
 sg13g2_tiehi _5214__32 (.L_HI(net32));
 sg13g2_tiehi _5215__33 (.L_HI(net33));
 sg13g2_tiehi _5216__34 (.L_HI(net34));
 sg13g2_tiehi _5217__35 (.L_HI(net35));
 sg13g2_tiehi _5218__36 (.L_HI(net36));
 sg13g2_tiehi _5219__37 (.L_HI(net37));
 sg13g2_tiehi _5220__38 (.L_HI(net38));
 sg13g2_tiehi _5221__39 (.L_HI(net39));
 sg13g2_tiehi _5222__40 (.L_HI(net40));
 sg13g2_tiehi _5223__41 (.L_HI(net41));
 sg13g2_tiehi _5224__42 (.L_HI(net42));
 sg13g2_tiehi _5225__43 (.L_HI(net43));
 sg13g2_tiehi _5226__44 (.L_HI(net44));
 sg13g2_tiehi _5227__45 (.L_HI(net45));
 sg13g2_tiehi _5228__46 (.L_HI(net46));
 sg13g2_tiehi _5229__47 (.L_HI(net47));
 sg13g2_tiehi _5230__48 (.L_HI(net48));
 sg13g2_tiehi _5231__49 (.L_HI(net49));
 sg13g2_tiehi _5232__50 (.L_HI(net50));
 sg13g2_tiehi _5233__51 (.L_HI(net51));
 sg13g2_tiehi _5234__52 (.L_HI(net52));
 sg13g2_tiehi _5235__53 (.L_HI(net53));
 sg13g2_tiehi _5236__54 (.L_HI(net54));
 sg13g2_tiehi _5237__55 (.L_HI(net55));
 sg13g2_tiehi _5238__56 (.L_HI(net56));
 sg13g2_tiehi _5239__57 (.L_HI(net57));
 sg13g2_tiehi _5240__58 (.L_HI(net58));
 sg13g2_tiehi _5241__59 (.L_HI(net59));
 sg13g2_tiehi _5242__60 (.L_HI(net60));
 sg13g2_tiehi _5243__61 (.L_HI(net61));
 sg13g2_tiehi _5244__62 (.L_HI(net62));
 sg13g2_tiehi _5245__63 (.L_HI(net63));
 sg13g2_tiehi _5246__64 (.L_HI(net64));
 sg13g2_tiehi _5247__65 (.L_HI(net65));
 sg13g2_tiehi _5248__66 (.L_HI(net66));
 sg13g2_tiehi _5249__67 (.L_HI(net67));
 sg13g2_tiehi _5288__68 (.L_HI(net68));
 sg13g2_tiehi _5297__69 (.L_HI(net69));
 sg13g2_tiehi _5250__70 (.L_HI(net70));
 sg13g2_tiehi _5251__71 (.L_HI(net71));
 sg13g2_tiehi tt_um_tt08_wirecube_72 (.L_HI(net72));
 sg13g2_inv_1 _2701__1 (.Y(net73),
    .A(clknet_1_0__leaf_clk));
 sg13g2_tielo tt_um_tt08_wirecube_11 (.L_LO(net11));
 sg13g2_tielo tt_um_tt08_wirecube_12 (.L_LO(net12));
 sg13g2_tielo tt_um_tt08_wirecube_13 (.L_LO(net13));
 sg13g2_tielo tt_um_tt08_wirecube_14 (.L_LO(net14));
 sg13g2_tielo tt_um_tt08_wirecube_15 (.L_LO(net15));
 sg13g2_tielo tt_um_tt08_wirecube_16 (.L_LO(net16));
 sg13g2_tielo tt_um_tt08_wirecube_17 (.L_LO(net17));
 sg13g2_tielo tt_um_tt08_wirecube_18 (.L_LO(net18));
 sg13g2_tielo tt_um_tt08_wirecube_19 (.L_LO(net19));
 sg13g2_tielo tt_um_tt08_wirecube_20 (.L_LO(net20));
 sg13g2_tielo tt_um_tt08_wirecube_21 (.L_LO(net21));
 sg13g2_tielo tt_um_tt08_wirecube_22 (.L_LO(net22));
 sg13g2_tielo tt_um_tt08_wirecube_23 (.L_LO(net23));
 sg13g2_tielo tt_um_tt08_wirecube_24 (.L_LO(net24));
 sg13g2_tiehi _5203__25 (.L_HI(net25));
 sg13g2_buf_1 _5372_ (.A(vsync),
    .X(uo_out[3]));
 sg13g2_buf_1 _5373_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout531 (.A(net532),
    .X(net531));
 sg13g2_buf_4 fanout532 (.X(net532),
    .A(_1432_));
 sg13g2_buf_2 fanout533 (.A(net534),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(net537),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(net536),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(net537),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_2543_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(_2538_),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(_2542_),
    .X(net539));
 sg13g2_buf_4 fanout540 (.X(net540),
    .A(_2295_));
 sg13g2_buf_2 fanout541 (.A(net542),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(net543),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(_2184_),
    .X(net543));
 sg13g2_buf_4 fanout544 (.X(net544),
    .A(net545));
 sg13g2_buf_2 fanout545 (.A(_2183_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_2183_),
    .X(net546));
 sg13g2_buf_1 fanout547 (.A(_2183_),
    .X(net547));
 sg13g2_buf_4 fanout548 (.X(net548),
    .A(_2175_));
 sg13g2_buf_2 fanout549 (.A(_2175_),
    .X(net549));
 sg13g2_buf_4 fanout550 (.X(net550),
    .A(net551));
 sg13g2_buf_2 fanout551 (.A(_2121_),
    .X(net551));
 sg13g2_buf_4 fanout552 (.X(net552),
    .A(_2120_));
 sg13g2_buf_4 fanout553 (.X(net553),
    .A(_2109_));
 sg13g2_buf_2 fanout554 (.A(_2109_),
    .X(net554));
 sg13g2_buf_4 fanout555 (.X(net555),
    .A(_2092_));
 sg13g2_buf_4 fanout556 (.X(net556),
    .A(_2090_));
 sg13g2_buf_4 fanout557 (.X(net557),
    .A(_2083_));
 sg13g2_buf_4 fanout558 (.X(net558),
    .A(_2082_));
 sg13g2_buf_1 fanout559 (.A(_2082_),
    .X(net559));
 sg13g2_buf_4 fanout560 (.X(net560),
    .A(_2054_));
 sg13g2_buf_4 fanout561 (.X(net561),
    .A(_2050_));
 sg13g2_buf_4 fanout562 (.X(net562),
    .A(_2049_));
 sg13g2_buf_2 fanout563 (.A(_2049_),
    .X(net563));
 sg13g2_buf_4 fanout564 (.X(net564),
    .A(_2039_));
 sg13g2_buf_4 fanout565 (.X(net565),
    .A(_2037_));
 sg13g2_buf_4 fanout566 (.X(net566),
    .A(_2036_));
 sg13g2_buf_2 fanout567 (.A(_2036_),
    .X(net567));
 sg13g2_buf_4 fanout568 (.X(net568),
    .A(_2034_));
 sg13g2_buf_4 fanout569 (.X(net569),
    .A(_2030_));
 sg13g2_buf_4 fanout570 (.X(net570),
    .A(_2025_));
 sg13g2_buf_1 fanout571 (.A(_2025_),
    .X(net571));
 sg13g2_buf_4 fanout572 (.X(net572),
    .A(_2007_));
 sg13g2_buf_4 fanout573 (.X(net573),
    .A(_2006_));
 sg13g2_buf_4 fanout574 (.X(net574),
    .A(_2003_));
 sg13g2_buf_4 fanout575 (.X(net575),
    .A(_2002_));
 sg13g2_buf_2 fanout576 (.A(net580),
    .X(net576));
 sg13g2_buf_1 fanout577 (.A(net580),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(net580),
    .X(net578));
 sg13g2_buf_1 fanout579 (.A(net580),
    .X(net579));
 sg13g2_buf_4 fanout580 (.X(net580),
    .A(_2020_));
 sg13g2_buf_2 fanout581 (.A(net582),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(net584),
    .X(net582));
 sg13g2_buf_4 fanout583 (.X(net583),
    .A(net584));
 sg13g2_buf_2 fanout584 (.A(_2014_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(net586),
    .X(net585));
 sg13g2_buf_4 fanout586 (.X(net586),
    .A(_2013_));
 sg13g2_buf_2 fanout587 (.A(_2013_),
    .X(net587));
 sg13g2_buf_1 fanout588 (.A(_2013_),
    .X(net588));
 sg13g2_buf_4 fanout589 (.X(net589),
    .A(_2005_));
 sg13g2_buf_2 fanout590 (.A(_2005_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(net592),
    .X(net591));
 sg13g2_buf_4 fanout592 (.X(net592),
    .A(_2004_));
 sg13g2_buf_2 fanout593 (.A(net594),
    .X(net593));
 sg13g2_buf_1 fanout594 (.A(net595),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(_1998_),
    .X(net595));
 sg13g2_buf_4 fanout596 (.X(net596),
    .A(_1998_));
 sg13g2_buf_2 fanout597 (.A(net598),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(net599),
    .X(net598));
 sg13g2_buf_4 fanout599 (.X(net599),
    .A(_1997_));
 sg13g2_buf_2 fanout600 (.A(net602),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(net602),
    .X(net601));
 sg13g2_buf_4 fanout602 (.X(net602),
    .A(_1994_));
 sg13g2_buf_4 fanout603 (.X(net603),
    .A(_1985_));
 sg13g2_buf_4 fanout604 (.X(net604),
    .A(_1984_));
 sg13g2_buf_1 fanout605 (.A(net606),
    .X(net605));
 sg13g2_buf_4 fanout606 (.X(net606),
    .A(_1984_));
 sg13g2_buf_2 fanout607 (.A(net608),
    .X(net607));
 sg13g2_buf_4 fanout608 (.X(net608),
    .A(_1977_));
 sg13g2_buf_2 fanout609 (.A(net610),
    .X(net609));
 sg13g2_buf_1 fanout610 (.A(_1977_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(net612),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(net617),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(net614),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(net615),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(net616),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(net617),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_1963_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(net620),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(net620),
    .X(net619));
 sg13g2_buf_4 fanout620 (.X(net620),
    .A(_1962_));
 sg13g2_buf_2 fanout621 (.A(net622),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(net623),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(net624),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_1962_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(net626),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_1862_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_1861_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_1861_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_1956_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_1940_),
    .X(net630));
 sg13g2_buf_1 fanout631 (.A(_1940_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(net633),
    .X(net632));
 sg13g2_buf_1 fanout633 (.A(net634),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(_1918_),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(net636),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(_1918_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(net638),
    .X(net637));
 sg13g2_buf_4 fanout638 (.X(net638),
    .A(_1917_));
 sg13g2_buf_2 fanout639 (.A(net640),
    .X(net639));
 sg13g2_buf_1 fanout640 (.A(net641),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(net642),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(_1917_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_1938_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(net645),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_1937_),
    .X(net645));
 sg13g2_buf_4 fanout646 (.X(net646),
    .A(_1511_));
 sg13g2_buf_4 fanout647 (.X(net647),
    .A(_2148_));
 sg13g2_buf_4 fanout648 (.X(net648),
    .A(_2131_));
 sg13g2_buf_4 fanout649 (.X(net649),
    .A(_2073_));
 sg13g2_buf_4 fanout650 (.X(net650),
    .A(_2072_));
 sg13g2_buf_2 fanout651 (.A(_2072_),
    .X(net651));
 sg13g2_buf_4 fanout652 (.X(net652),
    .A(_2071_));
 sg13g2_buf_4 fanout653 (.X(net653),
    .A(net654));
 sg13g2_buf_4 fanout654 (.X(net654),
    .A(_2066_));
 sg13g2_buf_4 fanout655 (.X(net655),
    .A(net656));
 sg13g2_buf_4 fanout656 (.X(net656),
    .A(_2150_));
 sg13g2_buf_2 fanout657 (.A(_2128_),
    .X(net657));
 sg13g2_buf_4 fanout658 (.X(net658),
    .A(_2127_));
 sg13g2_buf_4 fanout659 (.X(net659),
    .A(_2125_));
 sg13g2_buf_4 fanout660 (.X(net660),
    .A(_2103_));
 sg13g2_buf_4 fanout661 (.X(net661),
    .A(net662));
 sg13g2_buf_2 fanout662 (.A(_2100_),
    .X(net662));
 sg13g2_buf_4 fanout663 (.X(net663),
    .A(_2097_));
 sg13g2_buf_4 fanout664 (.X(net664),
    .A(net665));
 sg13g2_buf_2 fanout665 (.A(net675),
    .X(net665));
 sg13g2_buf_4 fanout666 (.X(net666),
    .A(net669));
 sg13g2_buf_4 fanout667 (.X(net667),
    .A(net669));
 sg13g2_buf_2 fanout668 (.A(net669),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(net675),
    .X(net669));
 sg13g2_buf_4 fanout670 (.X(net670),
    .A(net671));
 sg13g2_buf_2 fanout671 (.A(net675),
    .X(net671));
 sg13g2_buf_4 fanout672 (.X(net672),
    .A(net673));
 sg13g2_buf_4 fanout673 (.X(net673),
    .A(net675));
 sg13g2_buf_4 fanout674 (.X(net674),
    .A(net675));
 sg13g2_buf_4 fanout675 (.X(net675),
    .A(rst_n_sync));
 sg13g2_buf_8 fanout676 (.A(rst_n_sync),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(_2096_),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(\wirecube_top_inst.line_rom_inst.line_i[3] ),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(net680),
    .X(net679));
 sg13g2_buf_1 fanout680 (.A(\wirecube_top_inst.line_rom_inst.line_i[2] ),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(\wirecube_top_inst.edge_function_inst.pixel_x_i[2] ),
    .X(net681));
 sg13g2_buf_4 fanout682 (.X(net682),
    .A(\wirecube_top_inst.frame_cnt[12] ));
 sg13g2_buf_2 fanout683 (.A(net197),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(net200),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(net686),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(\wirecube_top_inst.cur_state_background[1] ),
    .X(net686));
 sg13g2_buf_4 fanout687 (.X(net687),
    .A(net162));
 sg13g2_buf_2 fanout688 (.A(\wirecube_top_inst.cur_state_background[0] ),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(net690),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(net691),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(net164),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(\wirecube_top_inst.frame_cnt[6] ),
    .X(net693));
 sg13g2_buf_4 fanout694 (.X(net694),
    .A(\wirecube_top_inst.frame_cnt[5] ));
 sg13g2_buf_4 fanout695 (.X(net695),
    .A(net177));
 sg13g2_buf_4 fanout696 (.X(net696),
    .A(\wirecube_top_inst.frame_cnt[3] ));
 sg13g2_buf_4 fanout697 (.X(net697),
    .A(net192));
 sg13g2_buf_2 fanout698 (.A(\wirecube_top_inst.frame_cnt[1] ),
    .X(net698));
 sg13g2_buf_4 fanout699 (.X(net699),
    .A(\wirecube_top_inst.counter_v[6] ));
 sg13g2_buf_2 fanout700 (.A(\wirecube_top_inst.counter_v[5] ),
    .X(net700));
 sg13g2_buf_4 fanout701 (.X(net701),
    .A(\wirecube_top_inst.counter_v[4] ));
 sg13g2_buf_2 fanout702 (.A(net199),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(net170),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(\wirecube_top_inst.counter_v[1] ),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(\wirecube_top_inst.edge_function_inst.term3[1] ),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(\wirecube_top_inst.edge_function_inst.term2[3] ),
    .X(net706));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_tielo tt_um_tt08_wirecube_10 (.L_LO(net10));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_2 clkbuf_5_0__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_1__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_2__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_3__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_4__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_5__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_6__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_7__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_8__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_9__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_10__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_11__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_12__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_13__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_14__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_15__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_16__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_17__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_18__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_19__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_20__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_21__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_22__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_23__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_24__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_25__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_26__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_27__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_28__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_29__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_30__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_31__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_5_7__leaf_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_5_11__leaf_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_5_15__leaf_clk_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_5_19__leaf_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_5_23__leaf_clk_regs));
 sg13g2_inv_1 clkload6 (.A(clknet_5_27__leaf_clk_regs));
 sg13g2_inv_1 clkload7 (.A(clknet_5_29__leaf_clk_regs));
 sg13g2_inv_1 clkload8 (.A(clknet_5_31__leaf_clk_regs));
 sg13g2_buf_2 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\wirecube_top_inst.delay_inst_hsync.pipe[0] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold2 (.A(\wirecube_top_inst.edge_function_inst.visible ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold3 (.A(\wirecube_top_inst.delay_inst_vsync.pipe[0] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0088_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0129_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0095_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0127_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0090_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0119_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0094_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0126_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0092_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0124_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0091_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0122_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0089_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold17 (.A(_1585_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold18 (.A(\wirecube_top_inst.any_line_set ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0152_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0093_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0125_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold22 (.A(\wirecube_top_inst.linecounter_h[0] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0000_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold24 (.A(\wirecube_top_inst.subcounter_v[2] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0117_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0096_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0128_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold28 (.A(\wirecube_top_inst.frame_cnt[12] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold29 (.A(\wirecube_top_inst.any_line_set2 ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold30 (.A(_1832_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0151_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold32 (.A(\wirecube_top_inst.final_pixel2 ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0142_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold34 (.A(\wirecube_top_inst.edge_function_inst.pixel_y_i[6] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold35 (.A(_1564_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold36 (.A(\wirecube_top_inst.subcounter_v[1] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0116_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0068_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold39 (.A(_1508_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold40 (.A(\wirecube_top_inst.counter_h[0] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold41 (.A(\wirecube_top_inst.line_rom_inst.line_i[3] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold42 (.A(\wirecube_top_inst.subcounter_v[0] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold43 (.A(\wirecube_top_inst.counter_v[1] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold44 (.A(_1524_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold45 (.A(\wirecube_top_inst.delay_inst_vsync.in_i ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold46 (.A(\wirecube_top_inst.counter_h[8] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold47 (.A(_1859_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0049_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold49 (.A(\wirecube_top_inst.edge_function_inst.pixel_y_i[5] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold50 (.A(_1561_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold51 (.A(\wirecube_top_inst.linecounter_h[1] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold52 (.A(\wirecube_top_inst.timing_hor.counter[11] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold53 (.A(\wirecube_top_inst.linecounter_h[3] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0003_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold55 (.A(\wirecube_top_inst.counter_h[10] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold56 (.A(_1867_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold57 (.A(\wirecube_top_inst.edge_function_inst.pixel_y_i[0] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold58 (.A(_1548_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0108_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold60 (.A(\wirecube_top_inst.edge_function_inst.pixel_x_i[6] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold61 (.A(_1828_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold62 (.A(\wirecube_top_inst.counter_h[9] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold63 (.A(\wirecube_top_inst.frame_cnt[0] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold64 (.A(_1609_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold65 (.A(\wirecube_top_inst.final_pixel ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold66 (.A(_1785_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0143_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold68 (.A(\wirecube_top_inst.counter_h[9] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold69 (.A(\wirecube_top_inst.delay_inst_hsync.in_i ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold70 (.A(\wirecube_top_inst.counter_h[4] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0059_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold72 (.A(\wirecube_top_inst.linecounter_h[2] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0002_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold74 (.A(\wirecube_top_inst.line_rom_inst.line_i[0] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0010_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold76 (.A(\wirecube_top_inst.edge_function_inst.pixel_y_i[2] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold77 (.A(_1554_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold78 (.A(\wirecube_top_inst.counter_h[3] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold79 (.A(_1506_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold80 (.A(\wirecube_top_inst.edge_function_inst.pixel_y_i[4] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold81 (.A(_1559_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold82 (.A(\wirecube_top_inst.counter_v[6] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold83 (.A(_1546_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0072_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0134_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold86 (.A(\wirecube_top_inst.counter_h[1] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0073_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0132_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold89 (.A(\wirecube_top_inst.cur_state_background[0] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold90 (.A(\wirecube_top_inst.counter_h[7] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold91 (.A(\wirecube_top_inst.frame_cnt[7] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0059_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0054_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold94 (.A(\wirecube_top_inst.counter_h[2] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold95 (.A(\wirecube_top_inst.edge_function_inst.pixel_x_i[1] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0145_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold97 (.A(\wirecube_top_inst.counter_v[2] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold98 (.A(\wirecube_top_inst.final_pixel ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold99 (.A(\wirecube_top_inst.counter_h[7] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold100 (.A(\wirecube_top_inst.counter_h[6] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold101 (.A(_1870_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold102 (.A(\wirecube_top_inst.counter_v[4] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold103 (.A(_1595_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold104 (.A(\wirecube_top_inst.frame_cnt[4] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0133_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0050_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0111_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0056_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0058_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0055_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold111 (.A(_1823_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0058_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold113 (.A(\wirecube_top_inst.edge_function_inst.pixel_x_i[0] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold114 (.A(\wirecube_top_inst.edge_function_inst.pixel_x_i[5] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold115 (.A(_1824_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0061_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0071_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0051_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold119 (.A(\wirecube_top_inst.frame_cnt[2] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0053_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold121 (.A(\wirecube_top_inst.edge_function_inst.pixel_x_i[3] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0052_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0057_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold124 (.A(\wirecube_top_inst.cur_state_background[3] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0140_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold126 (.A(\wirecube_top_inst.counter_v[3] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold127 (.A(\wirecube_top_inst.cur_state_background[2] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold128 (.A(\wirecube_top_inst.line_rom_inst.line_i[1] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold129 (.A(\wirecube_top_inst.counter_h[1] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0055_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold131 (.A(\wirecube_top_inst.edge_function_inst.pixel_y_i[2] ),
    .X(net204));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_fill_1 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_263 ();
 sg13g2_decap_8 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_277 ();
 sg13g2_decap_8 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_decap_4 FILLER_3_326 ();
 sg13g2_fill_2 FILLER_3_330 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_fill_2 FILLER_4_252 ();
 sg13g2_fill_1 FILLER_4_254 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_fill_2 FILLER_4_315 ();
 sg13g2_fill_2 FILLER_4_321 ();
 sg13g2_fill_1 FILLER_4_323 ();
 sg13g2_fill_1 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_354 ();
 sg13g2_decap_8 FILLER_4_361 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_4 FILLER_4_403 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_fill_2 FILLER_5_283 ();
 sg13g2_decap_8 FILLER_5_360 ();
 sg13g2_decap_8 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_374 ();
 sg13g2_decap_8 FILLER_5_381 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_fill_1 FILLER_6_203 ();
 sg13g2_fill_2 FILLER_6_230 ();
 sg13g2_fill_1 FILLER_6_356 ();
 sg13g2_decap_8 FILLER_6_365 ();
 sg13g2_decap_8 FILLER_6_372 ();
 sg13g2_decap_8 FILLER_6_379 ();
 sg13g2_decap_8 FILLER_6_386 ();
 sg13g2_decap_8 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_400 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_4 FILLER_7_196 ();
 sg13g2_fill_1 FILLER_7_200 ();
 sg13g2_decap_4 FILLER_7_233 ();
 sg13g2_fill_2 FILLER_7_237 ();
 sg13g2_fill_2 FILLER_7_257 ();
 sg13g2_fill_1 FILLER_7_307 ();
 sg13g2_fill_2 FILLER_7_336 ();
 sg13g2_fill_1 FILLER_7_338 ();
 sg13g2_fill_2 FILLER_7_344 ();
 sg13g2_fill_2 FILLER_7_359 ();
 sg13g2_fill_1 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_376 ();
 sg13g2_decap_8 FILLER_7_383 ();
 sg13g2_decap_8 FILLER_7_390 ();
 sg13g2_decap_8 FILLER_7_397 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_4 FILLER_8_196 ();
 sg13g2_fill_1 FILLER_8_200 ();
 sg13g2_decap_8 FILLER_8_281 ();
 sg13g2_decap_8 FILLER_8_288 ();
 sg13g2_decap_8 FILLER_8_299 ();
 sg13g2_fill_2 FILLER_8_306 ();
 sg13g2_fill_1 FILLER_8_308 ();
 sg13g2_fill_2 FILLER_8_322 ();
 sg13g2_fill_1 FILLER_8_324 ();
 sg13g2_fill_2 FILLER_8_345 ();
 sg13g2_decap_8 FILLER_8_352 ();
 sg13g2_fill_2 FILLER_8_359 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_fill_2 FILLER_9_196 ();
 sg13g2_fill_1 FILLER_9_198 ();
 sg13g2_fill_1 FILLER_9_214 ();
 sg13g2_fill_1 FILLER_9_239 ();
 sg13g2_fill_2 FILLER_9_254 ();
 sg13g2_fill_1 FILLER_9_278 ();
 sg13g2_fill_1 FILLER_9_305 ();
 sg13g2_decap_4 FILLER_9_327 ();
 sg13g2_fill_2 FILLER_9_331 ();
 sg13g2_fill_1 FILLER_9_358 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_4 FILLER_10_182 ();
 sg13g2_fill_2 FILLER_10_186 ();
 sg13g2_fill_2 FILLER_10_254 ();
 sg13g2_fill_2 FILLER_10_266 ();
 sg13g2_decap_4 FILLER_10_287 ();
 sg13g2_fill_1 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_fill_2 FILLER_10_308 ();
 sg13g2_fill_1 FILLER_10_334 ();
 sg13g2_fill_2 FILLER_10_348 ();
 sg13g2_fill_1 FILLER_10_350 ();
 sg13g2_decap_4 FILLER_10_359 ();
 sg13g2_fill_1 FILLER_10_363 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_8 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_fill_2 FILLER_11_196 ();
 sg13g2_fill_1 FILLER_11_198 ();
 sg13g2_decap_4 FILLER_11_284 ();
 sg13g2_fill_1 FILLER_11_288 ();
 sg13g2_decap_8 FILLER_11_293 ();
 sg13g2_fill_2 FILLER_11_300 ();
 sg13g2_fill_1 FILLER_11_324 ();
 sg13g2_fill_1 FILLER_11_343 ();
 sg13g2_decap_4 FILLER_11_352 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_123 ();
 sg13g2_fill_2 FILLER_12_130 ();
 sg13g2_decap_4 FILLER_12_136 ();
 sg13g2_fill_1 FILLER_12_140 ();
 sg13g2_fill_2 FILLER_12_145 ();
 sg13g2_decap_8 FILLER_12_155 ();
 sg13g2_decap_8 FILLER_12_162 ();
 sg13g2_decap_8 FILLER_12_169 ();
 sg13g2_decap_8 FILLER_12_176 ();
 sg13g2_decap_8 FILLER_12_183 ();
 sg13g2_decap_8 FILLER_12_190 ();
 sg13g2_fill_2 FILLER_12_214 ();
 sg13g2_fill_1 FILLER_12_225 ();
 sg13g2_fill_2 FILLER_12_263 ();
 sg13g2_fill_1 FILLER_12_265 ();
 sg13g2_decap_4 FILLER_12_274 ();
 sg13g2_fill_2 FILLER_12_304 ();
 sg13g2_fill_1 FILLER_12_306 ();
 sg13g2_fill_1 FILLER_12_311 ();
 sg13g2_fill_2 FILLER_12_330 ();
 sg13g2_decap_8 FILLER_12_337 ();
 sg13g2_decap_8 FILLER_12_344 ();
 sg13g2_fill_2 FILLER_12_351 ();
 sg13g2_decap_4 FILLER_12_357 ();
 sg13g2_fill_1 FILLER_12_365 ();
 sg13g2_decap_4 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_fill_2 FILLER_13_91 ();
 sg13g2_fill_1 FILLER_13_93 ();
 sg13g2_decap_8 FILLER_13_99 ();
 sg13g2_fill_2 FILLER_13_106 ();
 sg13g2_decap_8 FILLER_13_114 ();
 sg13g2_fill_2 FILLER_13_137 ();
 sg13g2_fill_1 FILLER_13_139 ();
 sg13g2_fill_1 FILLER_13_148 ();
 sg13g2_decap_8 FILLER_13_183 ();
 sg13g2_fill_2 FILLER_13_190 ();
 sg13g2_fill_1 FILLER_13_192 ();
 sg13g2_decap_4 FILLER_13_201 ();
 sg13g2_fill_1 FILLER_13_205 ();
 sg13g2_fill_2 FILLER_13_254 ();
 sg13g2_fill_2 FILLER_13_266 ();
 sg13g2_fill_1 FILLER_13_276 ();
 sg13g2_decap_8 FILLER_13_313 ();
 sg13g2_fill_2 FILLER_13_324 ();
 sg13g2_fill_1 FILLER_13_326 ();
 sg13g2_fill_2 FILLER_13_335 ();
 sg13g2_decap_8 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_4 FILLER_14_88 ();
 sg13g2_fill_1 FILLER_14_92 ();
 sg13g2_fill_2 FILLER_14_97 ();
 sg13g2_fill_2 FILLER_14_108 ();
 sg13g2_fill_1 FILLER_14_110 ();
 sg13g2_fill_2 FILLER_14_133 ();
 sg13g2_fill_2 FILLER_14_161 ();
 sg13g2_fill_1 FILLER_14_163 ();
 sg13g2_decap_8 FILLER_14_194 ();
 sg13g2_decap_8 FILLER_14_201 ();
 sg13g2_fill_1 FILLER_14_208 ();
 sg13g2_fill_2 FILLER_14_226 ();
 sg13g2_fill_1 FILLER_14_228 ();
 sg13g2_decap_8 FILLER_14_300 ();
 sg13g2_fill_1 FILLER_14_307 ();
 sg13g2_fill_1 FILLER_14_312 ();
 sg13g2_fill_2 FILLER_14_342 ();
 sg13g2_fill_2 FILLER_14_357 ();
 sg13g2_fill_1 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_fill_1 FILLER_15_104 ();
 sg13g2_fill_2 FILLER_15_111 ();
 sg13g2_fill_2 FILLER_15_137 ();
 sg13g2_fill_1 FILLER_15_148 ();
 sg13g2_fill_2 FILLER_15_160 ();
 sg13g2_decap_8 FILLER_15_199 ();
 sg13g2_decap_8 FILLER_15_206 ();
 sg13g2_fill_2 FILLER_15_213 ();
 sg13g2_fill_1 FILLER_15_215 ();
 sg13g2_decap_4 FILLER_15_290 ();
 sg13g2_fill_2 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_fill_2 FILLER_16_89 ();
 sg13g2_decap_8 FILLER_16_114 ();
 sg13g2_fill_2 FILLER_16_121 ();
 sg13g2_decap_4 FILLER_16_128 ();
 sg13g2_decap_8 FILLER_16_137 ();
 sg13g2_fill_2 FILLER_16_144 ();
 sg13g2_fill_1 FILLER_16_153 ();
 sg13g2_fill_2 FILLER_16_166 ();
 sg13g2_decap_8 FILLER_16_190 ();
 sg13g2_decap_8 FILLER_16_214 ();
 sg13g2_fill_2 FILLER_16_221 ();
 sg13g2_fill_1 FILLER_16_223 ();
 sg13g2_fill_1 FILLER_16_247 ();
 sg13g2_fill_2 FILLER_16_252 ();
 sg13g2_fill_1 FILLER_16_254 ();
 sg13g2_decap_4 FILLER_16_259 ();
 sg13g2_fill_2 FILLER_16_277 ();
 sg13g2_fill_1 FILLER_16_279 ();
 sg13g2_fill_2 FILLER_16_306 ();
 sg13g2_fill_1 FILLER_16_308 ();
 sg13g2_fill_2 FILLER_16_315 ();
 sg13g2_fill_1 FILLER_16_317 ();
 sg13g2_decap_4 FILLER_16_330 ();
 sg13g2_fill_1 FILLER_16_334 ();
 sg13g2_decap_4 FILLER_16_348 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_fill_2 FILLER_16_391 ();
 sg13g2_fill_1 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_fill_2 FILLER_17_63 ();
 sg13g2_fill_1 FILLER_17_65 ();
 sg13g2_decap_4 FILLER_17_87 ();
 sg13g2_fill_2 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_4 FILLER_17_112 ();
 sg13g2_fill_2 FILLER_17_116 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_fill_1 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_164 ();
 sg13g2_fill_2 FILLER_17_171 ();
 sg13g2_fill_2 FILLER_17_187 ();
 sg13g2_decap_8 FILLER_17_235 ();
 sg13g2_decap_4 FILLER_17_242 ();
 sg13g2_fill_2 FILLER_17_246 ();
 sg13g2_fill_2 FILLER_17_278 ();
 sg13g2_fill_2 FILLER_17_316 ();
 sg13g2_fill_1 FILLER_17_318 ();
 sg13g2_fill_2 FILLER_17_324 ();
 sg13g2_fill_2 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_fill_2 FILLER_17_363 ();
 sg13g2_fill_1 FILLER_17_365 ();
 sg13g2_decap_4 FILLER_17_369 ();
 sg13g2_fill_1 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_4 FILLER_18_56 ();
 sg13g2_decap_4 FILLER_18_71 ();
 sg13g2_fill_1 FILLER_18_75 ();
 sg13g2_decap_4 FILLER_18_88 ();
 sg13g2_fill_2 FILLER_18_92 ();
 sg13g2_decap_4 FILLER_18_111 ();
 sg13g2_fill_1 FILLER_18_115 ();
 sg13g2_decap_8 FILLER_18_135 ();
 sg13g2_fill_1 FILLER_18_167 ();
 sg13g2_fill_2 FILLER_18_196 ();
 sg13g2_fill_2 FILLER_18_221 ();
 sg13g2_fill_2 FILLER_18_238 ();
 sg13g2_fill_2 FILLER_18_289 ();
 sg13g2_decap_8 FILLER_18_299 ();
 sg13g2_fill_2 FILLER_18_306 ();
 sg13g2_fill_2 FILLER_18_325 ();
 sg13g2_fill_2 FILLER_18_338 ();
 sg13g2_fill_1 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_349 ();
 sg13g2_decap_8 FILLER_18_356 ();
 sg13g2_fill_2 FILLER_18_363 ();
 sg13g2_fill_1 FILLER_18_365 ();
 sg13g2_fill_2 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_4 FILLER_19_56 ();
 sg13g2_fill_2 FILLER_19_60 ();
 sg13g2_fill_1 FILLER_19_74 ();
 sg13g2_decap_8 FILLER_19_95 ();
 sg13g2_decap_4 FILLER_19_102 ();
 sg13g2_fill_2 FILLER_19_106 ();
 sg13g2_fill_2 FILLER_19_146 ();
 sg13g2_fill_1 FILLER_19_148 ();
 sg13g2_fill_2 FILLER_19_165 ();
 sg13g2_fill_1 FILLER_19_167 ();
 sg13g2_fill_2 FILLER_19_197 ();
 sg13g2_fill_1 FILLER_19_218 ();
 sg13g2_fill_2 FILLER_19_250 ();
 sg13g2_fill_1 FILLER_19_260 ();
 sg13g2_decap_8 FILLER_19_296 ();
 sg13g2_fill_1 FILLER_19_307 ();
 sg13g2_fill_2 FILLER_19_312 ();
 sg13g2_fill_2 FILLER_19_335 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_fill_1 FILLER_20_63 ();
 sg13g2_fill_1 FILLER_20_76 ();
 sg13g2_fill_1 FILLER_20_83 ();
 sg13g2_fill_2 FILLER_20_94 ();
 sg13g2_fill_2 FILLER_20_108 ();
 sg13g2_fill_1 FILLER_20_110 ();
 sg13g2_decap_4 FILLER_20_137 ();
 sg13g2_fill_2 FILLER_20_141 ();
 sg13g2_fill_2 FILLER_20_160 ();
 sg13g2_fill_1 FILLER_20_162 ();
 sg13g2_decap_4 FILLER_20_171 ();
 sg13g2_fill_2 FILLER_20_175 ();
 sg13g2_fill_1 FILLER_20_185 ();
 sg13g2_decap_8 FILLER_20_191 ();
 sg13g2_decap_4 FILLER_20_198 ();
 sg13g2_fill_1 FILLER_20_202 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_fill_2 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_244 ();
 sg13g2_fill_2 FILLER_20_279 ();
 sg13g2_fill_1 FILLER_20_281 ();
 sg13g2_fill_1 FILLER_20_343 ();
 sg13g2_fill_1 FILLER_20_360 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_fill_2 FILLER_21_49 ();
 sg13g2_fill_2 FILLER_21_105 ();
 sg13g2_fill_1 FILLER_21_107 ();
 sg13g2_fill_2 FILLER_21_126 ();
 sg13g2_fill_1 FILLER_21_128 ();
 sg13g2_decap_4 FILLER_21_140 ();
 sg13g2_fill_1 FILLER_21_144 ();
 sg13g2_fill_2 FILLER_21_160 ();
 sg13g2_fill_2 FILLER_21_174 ();
 sg13g2_fill_1 FILLER_21_176 ();
 sg13g2_fill_1 FILLER_21_181 ();
 sg13g2_decap_8 FILLER_21_187 ();
 sg13g2_fill_2 FILLER_21_194 ();
 sg13g2_fill_2 FILLER_21_201 ();
 sg13g2_fill_1 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_208 ();
 sg13g2_decap_8 FILLER_21_215 ();
 sg13g2_fill_1 FILLER_21_222 ();
 sg13g2_fill_2 FILLER_21_238 ();
 sg13g2_fill_1 FILLER_21_240 ();
 sg13g2_fill_1 FILLER_21_246 ();
 sg13g2_fill_2 FILLER_21_262 ();
 sg13g2_fill_1 FILLER_21_264 ();
 sg13g2_decap_8 FILLER_21_284 ();
 sg13g2_fill_2 FILLER_21_291 ();
 sg13g2_decap_8 FILLER_21_297 ();
 sg13g2_fill_1 FILLER_21_304 ();
 sg13g2_fill_2 FILLER_21_309 ();
 sg13g2_fill_1 FILLER_21_311 ();
 sg13g2_fill_1 FILLER_21_331 ();
 sg13g2_decap_8 FILLER_21_345 ();
 sg13g2_fill_1 FILLER_21_352 ();
 sg13g2_decap_4 FILLER_21_388 ();
 sg13g2_fill_2 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_fill_2 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_71 ();
 sg13g2_fill_2 FILLER_22_78 ();
 sg13g2_fill_2 FILLER_22_124 ();
 sg13g2_fill_1 FILLER_22_126 ();
 sg13g2_decap_4 FILLER_22_140 ();
 sg13g2_fill_2 FILLER_22_144 ();
 sg13g2_fill_2 FILLER_22_186 ();
 sg13g2_fill_2 FILLER_22_194 ();
 sg13g2_decap_8 FILLER_22_216 ();
 sg13g2_fill_2 FILLER_22_223 ();
 sg13g2_fill_2 FILLER_22_258 ();
 sg13g2_fill_2 FILLER_22_269 ();
 sg13g2_fill_1 FILLER_22_271 ();
 sg13g2_decap_4 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_316 ();
 sg13g2_fill_2 FILLER_22_323 ();
 sg13g2_fill_1 FILLER_22_325 ();
 sg13g2_fill_1 FILLER_22_334 ();
 sg13g2_fill_2 FILLER_22_343 ();
 sg13g2_fill_1 FILLER_22_345 ();
 sg13g2_decap_8 FILLER_22_359 ();
 sg13g2_decap_8 FILLER_22_366 ();
 sg13g2_fill_1 FILLER_22_373 ();
 sg13g2_fill_2 FILLER_22_381 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_fill_2 FILLER_23_49 ();
 sg13g2_fill_1 FILLER_23_51 ();
 sg13g2_decap_4 FILLER_23_66 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_decap_4 FILLER_23_128 ();
 sg13g2_fill_2 FILLER_23_147 ();
 sg13g2_fill_2 FILLER_23_160 ();
 sg13g2_fill_1 FILLER_23_194 ();
 sg13g2_fill_2 FILLER_23_210 ();
 sg13g2_fill_2 FILLER_23_226 ();
 sg13g2_decap_8 FILLER_23_233 ();
 sg13g2_fill_2 FILLER_23_240 ();
 sg13g2_fill_1 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_fill_1 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_286 ();
 sg13g2_fill_2 FILLER_23_293 ();
 sg13g2_decap_8 FILLER_23_299 ();
 sg13g2_fill_2 FILLER_23_306 ();
 sg13g2_fill_1 FILLER_23_323 ();
 sg13g2_fill_2 FILLER_23_337 ();
 sg13g2_decap_8 FILLER_23_352 ();
 sg13g2_fill_2 FILLER_23_359 ();
 sg13g2_fill_1 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_fill_2 FILLER_24_42 ();
 sg13g2_fill_1 FILLER_24_44 ();
 sg13g2_decap_4 FILLER_24_78 ();
 sg13g2_fill_1 FILLER_24_82 ();
 sg13g2_decap_4 FILLER_24_99 ();
 sg13g2_fill_1 FILLER_24_120 ();
 sg13g2_fill_2 FILLER_24_127 ();
 sg13g2_fill_1 FILLER_24_129 ();
 sg13g2_fill_2 FILLER_24_135 ();
 sg13g2_decap_8 FILLER_24_142 ();
 sg13g2_decap_8 FILLER_24_149 ();
 sg13g2_fill_1 FILLER_24_156 ();
 sg13g2_fill_2 FILLER_24_165 ();
 sg13g2_fill_2 FILLER_24_181 ();
 sg13g2_fill_1 FILLER_24_193 ();
 sg13g2_fill_2 FILLER_24_226 ();
 sg13g2_fill_1 FILLER_24_228 ();
 sg13g2_fill_2 FILLER_24_244 ();
 sg13g2_fill_1 FILLER_24_246 ();
 sg13g2_fill_1 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_285 ();
 sg13g2_decap_8 FILLER_24_292 ();
 sg13g2_fill_2 FILLER_24_299 ();
 sg13g2_fill_2 FILLER_24_346 ();
 sg13g2_fill_1 FILLER_24_348 ();
 sg13g2_fill_2 FILLER_24_356 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_4 FILLER_25_42 ();
 sg13g2_fill_1 FILLER_25_46 ();
 sg13g2_fill_2 FILLER_25_55 ();
 sg13g2_fill_1 FILLER_25_57 ();
 sg13g2_fill_1 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_76 ();
 sg13g2_decap_8 FILLER_25_83 ();
 sg13g2_decap_8 FILLER_25_90 ();
 sg13g2_decap_8 FILLER_25_97 ();
 sg13g2_fill_2 FILLER_25_104 ();
 sg13g2_fill_1 FILLER_25_122 ();
 sg13g2_decap_4 FILLER_25_144 ();
 sg13g2_fill_1 FILLER_25_148 ();
 sg13g2_decap_8 FILLER_25_166 ();
 sg13g2_fill_1 FILLER_25_177 ();
 sg13g2_decap_8 FILLER_25_186 ();
 sg13g2_decap_4 FILLER_25_193 ();
 sg13g2_fill_2 FILLER_25_197 ();
 sg13g2_fill_1 FILLER_25_203 ();
 sg13g2_decap_4 FILLER_25_238 ();
 sg13g2_decap_4 FILLER_25_248 ();
 sg13g2_decap_8 FILLER_25_270 ();
 sg13g2_decap_4 FILLER_25_303 ();
 sg13g2_fill_2 FILLER_25_307 ();
 sg13g2_decap_4 FILLER_25_318 ();
 sg13g2_fill_2 FILLER_25_339 ();
 sg13g2_fill_1 FILLER_25_341 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_4 FILLER_26_35 ();
 sg13g2_fill_1 FILLER_26_39 ();
 sg13g2_fill_1 FILLER_26_99 ();
 sg13g2_decap_4 FILLER_26_106 ();
 sg13g2_fill_1 FILLER_26_110 ();
 sg13g2_decap_4 FILLER_26_121 ();
 sg13g2_fill_1 FILLER_26_141 ();
 sg13g2_fill_1 FILLER_26_157 ();
 sg13g2_fill_1 FILLER_26_178 ();
 sg13g2_decap_8 FILLER_26_200 ();
 sg13g2_fill_1 FILLER_26_213 ();
 sg13g2_fill_2 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_fill_1 FILLER_26_323 ();
 sg13g2_decap_4 FILLER_26_329 ();
 sg13g2_fill_1 FILLER_26_333 ();
 sg13g2_decap_8 FILLER_26_342 ();
 sg13g2_fill_1 FILLER_26_349 ();
 sg13g2_decap_4 FILLER_26_355 ();
 sg13g2_fill_1 FILLER_26_359 ();
 sg13g2_fill_2 FILLER_26_367 ();
 sg13g2_decap_8 FILLER_26_379 ();
 sg13g2_fill_1 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_fill_2 FILLER_27_61 ();
 sg13g2_fill_2 FILLER_27_69 ();
 sg13g2_fill_2 FILLER_27_87 ();
 sg13g2_fill_1 FILLER_27_113 ();
 sg13g2_decap_8 FILLER_27_120 ();
 sg13g2_decap_8 FILLER_27_206 ();
 sg13g2_decap_8 FILLER_27_213 ();
 sg13g2_fill_2 FILLER_27_220 ();
 sg13g2_fill_1 FILLER_27_222 ();
 sg13g2_fill_1 FILLER_27_238 ();
 sg13g2_fill_2 FILLER_27_244 ();
 sg13g2_fill_2 FILLER_27_302 ();
 sg13g2_fill_1 FILLER_27_330 ();
 sg13g2_fill_1 FILLER_27_340 ();
 sg13g2_fill_2 FILLER_27_346 ();
 sg13g2_decap_8 FILLER_27_351 ();
 sg13g2_decap_8 FILLER_27_358 ();
 sg13g2_decap_4 FILLER_27_365 ();
 sg13g2_decap_8 FILLER_27_373 ();
 sg13g2_fill_1 FILLER_27_380 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_67 ();
 sg13g2_fill_2 FILLER_28_74 ();
 sg13g2_fill_1 FILLER_28_76 ();
 sg13g2_decap_4 FILLER_28_81 ();
 sg13g2_decap_4 FILLER_28_97 ();
 sg13g2_fill_2 FILLER_28_101 ();
 sg13g2_fill_2 FILLER_28_109 ();
 sg13g2_fill_1 FILLER_28_111 ();
 sg13g2_fill_1 FILLER_28_127 ();
 sg13g2_fill_2 FILLER_28_144 ();
 sg13g2_fill_1 FILLER_28_146 ();
 sg13g2_fill_2 FILLER_28_170 ();
 sg13g2_decap_8 FILLER_28_211 ();
 sg13g2_decap_8 FILLER_28_218 ();
 sg13g2_fill_1 FILLER_28_225 ();
 sg13g2_decap_4 FILLER_28_231 ();
 sg13g2_fill_1 FILLER_28_247 ();
 sg13g2_fill_2 FILLER_28_254 ();
 sg13g2_fill_1 FILLER_28_309 ();
 sg13g2_fill_1 FILLER_28_322 ();
 sg13g2_fill_2 FILLER_28_336 ();
 sg13g2_fill_2 FILLER_28_358 ();
 sg13g2_decap_8 FILLER_28_368 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_4 FILLER_29_49 ();
 sg13g2_fill_1 FILLER_29_53 ();
 sg13g2_decap_8 FILLER_29_69 ();
 sg13g2_decap_4 FILLER_29_76 ();
 sg13g2_decap_4 FILLER_29_92 ();
 sg13g2_fill_2 FILLER_29_121 ();
 sg13g2_fill_1 FILLER_29_123 ();
 sg13g2_fill_2 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_163 ();
 sg13g2_fill_2 FILLER_29_170 ();
 sg13g2_decap_4 FILLER_29_190 ();
 sg13g2_decap_8 FILLER_29_198 ();
 sg13g2_decap_4 FILLER_29_205 ();
 sg13g2_fill_1 FILLER_29_209 ();
 sg13g2_fill_2 FILLER_29_224 ();
 sg13g2_fill_2 FILLER_29_240 ();
 sg13g2_fill_1 FILLER_29_242 ();
 sg13g2_fill_2 FILLER_29_247 ();
 sg13g2_fill_1 FILLER_29_249 ();
 sg13g2_fill_1 FILLER_29_255 ();
 sg13g2_fill_2 FILLER_29_266 ();
 sg13g2_fill_1 FILLER_29_286 ();
 sg13g2_fill_2 FILLER_29_313 ();
 sg13g2_fill_1 FILLER_29_315 ();
 sg13g2_fill_1 FILLER_29_329 ();
 sg13g2_decap_4 FILLER_29_338 ();
 sg13g2_fill_2 FILLER_29_374 ();
 sg13g2_fill_1 FILLER_29_376 ();
 sg13g2_fill_2 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_4 FILLER_30_35 ();
 sg13g2_fill_2 FILLER_30_39 ();
 sg13g2_fill_2 FILLER_30_59 ();
 sg13g2_fill_1 FILLER_30_76 ();
 sg13g2_fill_2 FILLER_30_88 ();
 sg13g2_fill_1 FILLER_30_90 ();
 sg13g2_fill_2 FILLER_30_109 ();
 sg13g2_fill_2 FILLER_30_117 ();
 sg13g2_fill_2 FILLER_30_147 ();
 sg13g2_fill_1 FILLER_30_149 ();
 sg13g2_decap_8 FILLER_30_155 ();
 sg13g2_decap_8 FILLER_30_162 ();
 sg13g2_decap_8 FILLER_30_169 ();
 sg13g2_fill_2 FILLER_30_176 ();
 sg13g2_fill_1 FILLER_30_190 ();
 sg13g2_decap_8 FILLER_30_199 ();
 sg13g2_fill_2 FILLER_30_206 ();
 sg13g2_decap_4 FILLER_30_216 ();
 sg13g2_fill_2 FILLER_30_225 ();
 sg13g2_fill_1 FILLER_30_227 ();
 sg13g2_decap_4 FILLER_30_245 ();
 sg13g2_fill_1 FILLER_30_253 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_decap_4 FILLER_30_265 ();
 sg13g2_fill_1 FILLER_30_274 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_4 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_302 ();
 sg13g2_fill_1 FILLER_30_309 ();
 sg13g2_decap_8 FILLER_30_314 ();
 sg13g2_fill_2 FILLER_30_321 ();
 sg13g2_fill_1 FILLER_30_323 ();
 sg13g2_fill_2 FILLER_30_329 ();
 sg13g2_fill_2 FILLER_30_339 ();
 sg13g2_fill_2 FILLER_30_376 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_4 FILLER_31_35 ();
 sg13g2_fill_2 FILLER_31_62 ();
 sg13g2_fill_1 FILLER_31_64 ();
 sg13g2_decap_4 FILLER_31_93 ();
 sg13g2_decap_4 FILLER_31_124 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_decap_4 FILLER_31_135 ();
 sg13g2_decap_4 FILLER_31_148 ();
 sg13g2_fill_2 FILLER_31_152 ();
 sg13g2_decap_8 FILLER_31_159 ();
 sg13g2_fill_1 FILLER_31_170 ();
 sg13g2_fill_2 FILLER_31_185 ();
 sg13g2_decap_8 FILLER_31_209 ();
 sg13g2_fill_1 FILLER_31_216 ();
 sg13g2_fill_1 FILLER_31_227 ();
 sg13g2_decap_8 FILLER_31_248 ();
 sg13g2_decap_8 FILLER_31_255 ();
 sg13g2_decap_8 FILLER_31_262 ();
 sg13g2_decap_4 FILLER_31_269 ();
 sg13g2_fill_2 FILLER_31_273 ();
 sg13g2_fill_2 FILLER_31_301 ();
 sg13g2_fill_1 FILLER_31_303 ();
 sg13g2_fill_1 FILLER_31_318 ();
 sg13g2_decap_4 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_31_341 ();
 sg13g2_fill_2 FILLER_31_348 ();
 sg13g2_fill_1 FILLER_31_350 ();
 sg13g2_fill_2 FILLER_31_364 ();
 sg13g2_decap_4 FILLER_31_374 ();
 sg13g2_fill_2 FILLER_31_378 ();
 sg13g2_fill_2 FILLER_31_393 ();
 sg13g2_fill_1 FILLER_31_395 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_fill_2 FILLER_32_42 ();
 sg13g2_fill_2 FILLER_32_54 ();
 sg13g2_fill_1 FILLER_32_56 ();
 sg13g2_fill_1 FILLER_32_62 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_110 ();
 sg13g2_decap_8 FILLER_32_117 ();
 sg13g2_decap_4 FILLER_32_132 ();
 sg13g2_fill_1 FILLER_32_136 ();
 sg13g2_fill_2 FILLER_32_149 ();
 sg13g2_fill_2 FILLER_32_181 ();
 sg13g2_fill_2 FILLER_32_213 ();
 sg13g2_fill_1 FILLER_32_215 ();
 sg13g2_decap_4 FILLER_32_220 ();
 sg13g2_fill_1 FILLER_32_224 ();
 sg13g2_decap_4 FILLER_32_238 ();
 sg13g2_decap_4 FILLER_32_270 ();
 sg13g2_fill_2 FILLER_32_274 ();
 sg13g2_fill_1 FILLER_32_330 ();
 sg13g2_decap_8 FILLER_32_339 ();
 sg13g2_decap_4 FILLER_32_346 ();
 sg13g2_decap_8 FILLER_32_354 ();
 sg13g2_decap_8 FILLER_32_365 ();
 sg13g2_decap_8 FILLER_32_372 ();
 sg13g2_decap_4 FILLER_32_379 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_4 FILLER_33_42 ();
 sg13g2_fill_2 FILLER_33_46 ();
 sg13g2_fill_2 FILLER_33_52 ();
 sg13g2_fill_2 FILLER_33_72 ();
 sg13g2_fill_1 FILLER_33_74 ();
 sg13g2_fill_2 FILLER_33_81 ();
 sg13g2_fill_2 FILLER_33_111 ();
 sg13g2_fill_1 FILLER_33_132 ();
 sg13g2_decap_4 FILLER_33_147 ();
 sg13g2_fill_2 FILLER_33_160 ();
 sg13g2_fill_1 FILLER_33_162 ();
 sg13g2_fill_1 FILLER_33_190 ();
 sg13g2_fill_2 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_230 ();
 sg13g2_fill_2 FILLER_33_247 ();
 sg13g2_decap_4 FILLER_33_277 ();
 sg13g2_decap_8 FILLER_33_330 ();
 sg13g2_fill_2 FILLER_33_337 ();
 sg13g2_fill_1 FILLER_33_346 ();
 sg13g2_fill_1 FILLER_33_387 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_4 FILLER_34_35 ();
 sg13g2_fill_2 FILLER_34_64 ();
 sg13g2_decap_4 FILLER_34_79 ();
 sg13g2_fill_1 FILLER_34_83 ();
 sg13g2_fill_2 FILLER_34_122 ();
 sg13g2_fill_1 FILLER_34_124 ();
 sg13g2_fill_1 FILLER_34_129 ();
 sg13g2_fill_2 FILLER_34_135 ();
 sg13g2_decap_4 FILLER_34_142 ();
 sg13g2_fill_1 FILLER_34_160 ();
 sg13g2_fill_1 FILLER_34_215 ();
 sg13g2_fill_1 FILLER_34_246 ();
 sg13g2_decap_8 FILLER_34_275 ();
 sg13g2_decap_4 FILLER_34_282 ();
 sg13g2_fill_1 FILLER_34_286 ();
 sg13g2_fill_1 FILLER_34_291 ();
 sg13g2_decap_8 FILLER_34_296 ();
 sg13g2_fill_2 FILLER_34_303 ();
 sg13g2_fill_1 FILLER_34_305 ();
 sg13g2_fill_2 FILLER_34_328 ();
 sg13g2_fill_1 FILLER_34_330 ();
 sg13g2_fill_1 FILLER_34_343 ();
 sg13g2_fill_1 FILLER_34_369 ();
 sg13g2_fill_2 FILLER_34_393 ();
 sg13g2_fill_1 FILLER_34_395 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_fill_2 FILLER_35_47 ();
 sg13g2_fill_1 FILLER_35_49 ();
 sg13g2_fill_2 FILLER_35_55 ();
 sg13g2_fill_1 FILLER_35_73 ();
 sg13g2_fill_1 FILLER_35_79 ();
 sg13g2_decap_8 FILLER_35_101 ();
 sg13g2_fill_1 FILLER_35_108 ();
 sg13g2_decap_4 FILLER_35_125 ();
 sg13g2_fill_1 FILLER_35_129 ();
 sg13g2_decap_4 FILLER_35_148 ();
 sg13g2_decap_4 FILLER_35_174 ();
 sg13g2_decap_4 FILLER_35_189 ();
 sg13g2_fill_1 FILLER_35_193 ();
 sg13g2_decap_8 FILLER_35_198 ();
 sg13g2_decap_8 FILLER_35_205 ();
 sg13g2_decap_8 FILLER_35_212 ();
 sg13g2_fill_2 FILLER_35_219 ();
 sg13g2_decap_8 FILLER_35_236 ();
 sg13g2_decap_8 FILLER_35_243 ();
 sg13g2_decap_4 FILLER_35_250 ();
 sg13g2_fill_2 FILLER_35_258 ();
 sg13g2_decap_8 FILLER_35_265 ();
 sg13g2_decap_8 FILLER_35_272 ();
 sg13g2_decap_8 FILLER_35_279 ();
 sg13g2_fill_2 FILLER_35_286 ();
 sg13g2_fill_1 FILLER_35_288 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_fill_2 FILLER_35_322 ();
 sg13g2_fill_2 FILLER_35_327 ();
 sg13g2_fill_2 FILLER_35_365 ();
 sg13g2_fill_1 FILLER_35_384 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_4 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_46 ();
 sg13g2_decap_8 FILLER_36_57 ();
 sg13g2_fill_2 FILLER_36_79 ();
 sg13g2_fill_1 FILLER_36_86 ();
 sg13g2_decap_8 FILLER_36_92 ();
 sg13g2_decap_8 FILLER_36_99 ();
 sg13g2_fill_2 FILLER_36_106 ();
 sg13g2_decap_8 FILLER_36_114 ();
 sg13g2_fill_2 FILLER_36_121 ();
 sg13g2_decap_8 FILLER_36_128 ();
 sg13g2_decap_4 FILLER_36_135 ();
 sg13g2_fill_1 FILLER_36_139 ();
 sg13g2_decap_8 FILLER_36_145 ();
 sg13g2_decap_4 FILLER_36_152 ();
 sg13g2_fill_1 FILLER_36_156 ();
 sg13g2_decap_8 FILLER_36_170 ();
 sg13g2_fill_2 FILLER_36_177 ();
 sg13g2_fill_1 FILLER_36_179 ();
 sg13g2_decap_4 FILLER_36_185 ();
 sg13g2_decap_8 FILLER_36_206 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_fill_1 FILLER_36_220 ();
 sg13g2_fill_2 FILLER_36_228 ();
 sg13g2_fill_1 FILLER_36_234 ();
 sg13g2_fill_1 FILLER_36_240 ();
 sg13g2_fill_2 FILLER_36_249 ();
 sg13g2_fill_1 FILLER_36_251 ();
 sg13g2_fill_1 FILLER_36_275 ();
 sg13g2_decap_4 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_318 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_fill_2 FILLER_36_354 ();
 sg13g2_fill_1 FILLER_36_385 ();
 sg13g2_fill_2 FILLER_36_390 ();
 sg13g2_fill_1 FILLER_36_392 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_fill_1 FILLER_37_49 ();
 sg13g2_decap_4 FILLER_37_67 ();
 sg13g2_fill_2 FILLER_37_71 ();
 sg13g2_fill_2 FILLER_37_83 ();
 sg13g2_decap_4 FILLER_37_95 ();
 sg13g2_fill_2 FILLER_37_105 ();
 sg13g2_fill_1 FILLER_37_107 ();
 sg13g2_fill_1 FILLER_37_114 ();
 sg13g2_fill_1 FILLER_37_121 ();
 sg13g2_fill_1 FILLER_37_146 ();
 sg13g2_fill_1 FILLER_37_157 ();
 sg13g2_fill_1 FILLER_37_165 ();
 sg13g2_fill_2 FILLER_37_174 ();
 sg13g2_fill_1 FILLER_37_176 ();
 sg13g2_fill_2 FILLER_37_184 ();
 sg13g2_fill_1 FILLER_37_186 ();
 sg13g2_fill_2 FILLER_37_216 ();
 sg13g2_fill_2 FILLER_37_239 ();
 sg13g2_decap_4 FILLER_37_249 ();
 sg13g2_fill_2 FILLER_37_273 ();
 sg13g2_fill_1 FILLER_37_291 ();
 sg13g2_fill_2 FILLER_37_297 ();
 sg13g2_decap_8 FILLER_37_307 ();
 sg13g2_fill_1 FILLER_37_314 ();
 sg13g2_fill_2 FILLER_37_324 ();
 sg13g2_fill_1 FILLER_37_326 ();
 sg13g2_decap_4 FILLER_37_331 ();
 sg13g2_fill_2 FILLER_37_335 ();
 sg13g2_fill_2 FILLER_37_342 ();
 sg13g2_fill_1 FILLER_37_344 ();
 sg13g2_decap_8 FILLER_37_353 ();
 sg13g2_decap_4 FILLER_37_360 ();
 sg13g2_fill_2 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_376 ();
 sg13g2_decap_4 FILLER_37_383 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_fill_2 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_44 ();
 sg13g2_fill_2 FILLER_38_52 ();
 sg13g2_fill_2 FILLER_38_74 ();
 sg13g2_fill_2 FILLER_38_94 ();
 sg13g2_fill_1 FILLER_38_96 ();
 sg13g2_decap_8 FILLER_38_106 ();
 sg13g2_decap_4 FILLER_38_113 ();
 sg13g2_fill_2 FILLER_38_123 ();
 sg13g2_fill_1 FILLER_38_125 ();
 sg13g2_fill_2 FILLER_38_140 ();
 sg13g2_fill_2 FILLER_38_150 ();
 sg13g2_fill_1 FILLER_38_152 ();
 sg13g2_fill_1 FILLER_38_169 ();
 sg13g2_fill_2 FILLER_38_198 ();
 sg13g2_decap_4 FILLER_38_225 ();
 sg13g2_fill_2 FILLER_38_229 ();
 sg13g2_fill_1 FILLER_38_265 ();
 sg13g2_decap_4 FILLER_38_304 ();
 sg13g2_fill_2 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_338 ();
 sg13g2_fill_2 FILLER_38_345 ();
 sg13g2_fill_1 FILLER_38_347 ();
 sg13g2_decap_8 FILLER_38_353 ();
 sg13g2_decap_4 FILLER_38_360 ();
 sg13g2_fill_2 FILLER_38_383 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_4 FILLER_39_42 ();
 sg13g2_fill_2 FILLER_39_46 ();
 sg13g2_fill_2 FILLER_39_54 ();
 sg13g2_fill_1 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_62 ();
 sg13g2_fill_2 FILLER_39_69 ();
 sg13g2_fill_2 FILLER_39_76 ();
 sg13g2_fill_2 FILLER_39_90 ();
 sg13g2_fill_1 FILLER_39_108 ();
 sg13g2_decap_4 FILLER_39_125 ();
 sg13g2_fill_2 FILLER_39_139 ();
 sg13g2_fill_1 FILLER_39_183 ();
 sg13g2_decap_4 FILLER_39_214 ();
 sg13g2_fill_2 FILLER_39_226 ();
 sg13g2_decap_8 FILLER_39_244 ();
 sg13g2_fill_2 FILLER_39_287 ();
 sg13g2_fill_2 FILLER_39_315 ();
 sg13g2_fill_2 FILLER_39_324 ();
 sg13g2_fill_2 FILLER_39_334 ();
 sg13g2_fill_1 FILLER_39_336 ();
 sg13g2_decap_4 FILLER_39_350 ();
 sg13g2_fill_2 FILLER_39_362 ();
 sg13g2_fill_2 FILLER_39_376 ();
 sg13g2_fill_1 FILLER_39_378 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_4 FILLER_40_49 ();
 sg13g2_fill_1 FILLER_40_53 ();
 sg13g2_fill_1 FILLER_40_59 ();
 sg13g2_fill_2 FILLER_40_80 ();
 sg13g2_fill_2 FILLER_40_98 ();
 sg13g2_fill_2 FILLER_40_106 ();
 sg13g2_fill_2 FILLER_40_120 ();
 sg13g2_fill_2 FILLER_40_131 ();
 sg13g2_fill_1 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_138 ();
 sg13g2_decap_4 FILLER_40_145 ();
 sg13g2_fill_2 FILLER_40_149 ();
 sg13g2_fill_2 FILLER_40_172 ();
 sg13g2_fill_1 FILLER_40_196 ();
 sg13g2_decap_8 FILLER_40_204 ();
 sg13g2_decap_8 FILLER_40_211 ();
 sg13g2_fill_2 FILLER_40_218 ();
 sg13g2_fill_1 FILLER_40_220 ();
 sg13g2_fill_1 FILLER_40_240 ();
 sg13g2_decap_8 FILLER_40_249 ();
 sg13g2_decap_4 FILLER_40_256 ();
 sg13g2_fill_2 FILLER_40_260 ();
 sg13g2_fill_1 FILLER_40_291 ();
 sg13g2_decap_4 FILLER_40_297 ();
 sg13g2_fill_1 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_306 ();
 sg13g2_fill_1 FILLER_40_313 ();
 sg13g2_fill_1 FILLER_40_327 ();
 sg13g2_fill_2 FILLER_40_336 ();
 sg13g2_fill_1 FILLER_40_338 ();
 sg13g2_fill_2 FILLER_40_355 ();
 sg13g2_fill_1 FILLER_40_357 ();
 sg13g2_fill_2 FILLER_40_382 ();
 sg13g2_fill_1 FILLER_40_384 ();
 sg13g2_fill_2 FILLER_40_406 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_fill_2 FILLER_41_35 ();
 sg13g2_fill_1 FILLER_41_37 ();
 sg13g2_decap_4 FILLER_41_65 ();
 sg13g2_fill_1 FILLER_41_94 ();
 sg13g2_fill_2 FILLER_41_109 ();
 sg13g2_fill_1 FILLER_41_134 ();
 sg13g2_fill_2 FILLER_41_145 ();
 sg13g2_fill_1 FILLER_41_147 ();
 sg13g2_decap_4 FILLER_41_165 ();
 sg13g2_fill_2 FILLER_41_181 ();
 sg13g2_fill_2 FILLER_41_191 ();
 sg13g2_fill_1 FILLER_41_193 ();
 sg13g2_decap_4 FILLER_41_207 ();
 sg13g2_fill_2 FILLER_41_228 ();
 sg13g2_fill_2 FILLER_41_236 ();
 sg13g2_fill_1 FILLER_41_238 ();
 sg13g2_fill_1 FILLER_41_246 ();
 sg13g2_fill_2 FILLER_41_255 ();
 sg13g2_fill_1 FILLER_41_257 ();
 sg13g2_fill_1 FILLER_41_271 ();
 sg13g2_fill_2 FILLER_41_276 ();
 sg13g2_fill_1 FILLER_41_278 ();
 sg13g2_fill_1 FILLER_41_291 ();
 sg13g2_decap_8 FILLER_41_318 ();
 sg13g2_decap_4 FILLER_41_328 ();
 sg13g2_fill_2 FILLER_41_332 ();
 sg13g2_fill_1 FILLER_41_360 ();
 sg13g2_fill_2 FILLER_41_376 ();
 sg13g2_decap_8 FILLER_41_382 ();
 sg13g2_decap_4 FILLER_41_389 ();
 sg13g2_fill_2 FILLER_41_393 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_fill_2 FILLER_42_35 ();
 sg13g2_fill_1 FILLER_42_37 ();
 sg13g2_decap_4 FILLER_42_54 ();
 sg13g2_decap_8 FILLER_42_99 ();
 sg13g2_decap_4 FILLER_42_106 ();
 sg13g2_fill_1 FILLER_42_110 ();
 sg13g2_decap_4 FILLER_42_117 ();
 sg13g2_fill_1 FILLER_42_121 ();
 sg13g2_fill_2 FILLER_42_128 ();
 sg13g2_fill_2 FILLER_42_144 ();
 sg13g2_fill_1 FILLER_42_146 ();
 sg13g2_fill_2 FILLER_42_168 ();
 sg13g2_fill_1 FILLER_42_170 ();
 sg13g2_fill_2 FILLER_42_201 ();
 sg13g2_decap_8 FILLER_42_281 ();
 sg13g2_fill_2 FILLER_42_288 ();
 sg13g2_decap_8 FILLER_42_306 ();
 sg13g2_fill_2 FILLER_42_313 ();
 sg13g2_decap_8 FILLER_42_327 ();
 sg13g2_decap_8 FILLER_42_334 ();
 sg13g2_fill_2 FILLER_42_362 ();
 sg13g2_fill_1 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_373 ();
 sg13g2_decap_4 FILLER_42_380 ();
 sg13g2_fill_2 FILLER_42_384 ();
 sg13g2_fill_1 FILLER_42_390 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_4 FILLER_43_42 ();
 sg13g2_decap_4 FILLER_43_67 ();
 sg13g2_fill_1 FILLER_43_71 ();
 sg13g2_decap_8 FILLER_43_78 ();
 sg13g2_decap_8 FILLER_43_85 ();
 sg13g2_decap_4 FILLER_43_92 ();
 sg13g2_fill_2 FILLER_43_105 ();
 sg13g2_fill_1 FILLER_43_107 ();
 sg13g2_decap_4 FILLER_43_118 ();
 sg13g2_fill_1 FILLER_43_122 ();
 sg13g2_decap_4 FILLER_43_127 ();
 sg13g2_fill_2 FILLER_43_131 ();
 sg13g2_fill_2 FILLER_43_145 ();
 sg13g2_fill_2 FILLER_43_163 ();
 sg13g2_fill_1 FILLER_43_165 ();
 sg13g2_decap_4 FILLER_43_190 ();
 sg13g2_fill_2 FILLER_43_247 ();
 sg13g2_fill_2 FILLER_43_269 ();
 sg13g2_fill_1 FILLER_43_276 ();
 sg13g2_fill_2 FILLER_43_282 ();
 sg13g2_fill_1 FILLER_43_310 ();
 sg13g2_fill_2 FILLER_43_328 ();
 sg13g2_fill_1 FILLER_43_330 ();
 sg13g2_decap_4 FILLER_43_344 ();
 sg13g2_fill_2 FILLER_43_348 ();
 sg13g2_decap_8 FILLER_43_362 ();
 sg13g2_fill_2 FILLER_43_369 ();
 sg13g2_fill_1 FILLER_43_371 ();
 sg13g2_fill_2 FILLER_43_377 ();
 sg13g2_fill_1 FILLER_43_379 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_4 FILLER_44_42 ();
 sg13g2_fill_1 FILLER_44_46 ();
 sg13g2_decap_8 FILLER_44_55 ();
 sg13g2_decap_4 FILLER_44_62 ();
 sg13g2_fill_2 FILLER_44_66 ();
 sg13g2_fill_2 FILLER_44_74 ();
 sg13g2_fill_2 FILLER_44_101 ();
 sg13g2_fill_2 FILLER_44_111 ();
 sg13g2_fill_2 FILLER_44_124 ();
 sg13g2_fill_1 FILLER_44_134 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_158 ();
 sg13g2_decap_4 FILLER_44_165 ();
 sg13g2_fill_2 FILLER_44_169 ();
 sg13g2_fill_2 FILLER_44_183 ();
 sg13g2_fill_1 FILLER_44_185 ();
 sg13g2_decap_8 FILLER_44_192 ();
 sg13g2_decap_4 FILLER_44_199 ();
 sg13g2_fill_2 FILLER_44_203 ();
 sg13g2_fill_2 FILLER_44_238 ();
 sg13g2_fill_1 FILLER_44_240 ();
 sg13g2_fill_2 FILLER_44_273 ();
 sg13g2_fill_2 FILLER_44_283 ();
 sg13g2_fill_2 FILLER_44_316 ();
 sg13g2_fill_1 FILLER_44_341 ();
 sg13g2_fill_2 FILLER_44_360 ();
 sg13g2_fill_1 FILLER_44_381 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_fill_1 FILLER_45_62 ();
 sg13g2_decap_8 FILLER_45_89 ();
 sg13g2_fill_2 FILLER_45_104 ();
 sg13g2_fill_1 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_fill_1 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_170 ();
 sg13g2_decap_4 FILLER_45_177 ();
 sg13g2_fill_1 FILLER_45_181 ();
 sg13g2_decap_4 FILLER_45_192 ();
 sg13g2_decap_8 FILLER_45_202 ();
 sg13g2_decap_4 FILLER_45_209 ();
 sg13g2_fill_2 FILLER_45_213 ();
 sg13g2_decap_4 FILLER_45_238 ();
 sg13g2_fill_2 FILLER_45_242 ();
 sg13g2_fill_1 FILLER_45_315 ();
 sg13g2_fill_2 FILLER_45_359 ();
 sg13g2_fill_1 FILLER_45_361 ();
 sg13g2_decap_4 FILLER_45_404 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_fill_1 FILLER_46_35 ();
 sg13g2_fill_2 FILLER_46_83 ();
 sg13g2_fill_1 FILLER_46_85 ();
 sg13g2_fill_2 FILLER_46_92 ();
 sg13g2_fill_2 FILLER_46_118 ();
 sg13g2_fill_1 FILLER_46_120 ();
 sg13g2_fill_1 FILLER_46_127 ();
 sg13g2_fill_1 FILLER_46_150 ();
 sg13g2_fill_2 FILLER_46_160 ();
 sg13g2_fill_1 FILLER_46_162 ();
 sg13g2_decap_4 FILLER_46_169 ();
 sg13g2_fill_2 FILLER_46_173 ();
 sg13g2_fill_2 FILLER_46_181 ();
 sg13g2_fill_1 FILLER_46_183 ();
 sg13g2_fill_1 FILLER_46_193 ();
 sg13g2_decap_8 FILLER_46_207 ();
 sg13g2_decap_8 FILLER_46_214 ();
 sg13g2_fill_2 FILLER_46_221 ();
 sg13g2_decap_4 FILLER_46_231 ();
 sg13g2_fill_2 FILLER_46_247 ();
 sg13g2_decap_4 FILLER_46_311 ();
 sg13g2_fill_2 FILLER_46_333 ();
 sg13g2_fill_1 FILLER_46_335 ();
 sg13g2_fill_1 FILLER_46_347 ();
 sg13g2_decap_4 FILLER_46_360 ();
 sg13g2_fill_1 FILLER_46_368 ();
 sg13g2_decap_4 FILLER_46_373 ();
 sg13g2_fill_2 FILLER_46_381 ();
 sg13g2_fill_1 FILLER_46_387 ();
 sg13g2_decap_4 FILLER_46_393 ();
 sg13g2_decap_4 FILLER_46_404 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_fill_2 FILLER_47_42 ();
 sg13g2_fill_1 FILLER_47_65 ();
 sg13g2_decap_8 FILLER_47_82 ();
 sg13g2_fill_2 FILLER_47_89 ();
 sg13g2_fill_2 FILLER_47_105 ();
 sg13g2_fill_1 FILLER_47_107 ();
 sg13g2_fill_2 FILLER_47_132 ();
 sg13g2_fill_1 FILLER_47_164 ();
 sg13g2_fill_2 FILLER_47_212 ();
 sg13g2_fill_1 FILLER_47_214 ();
 sg13g2_decap_8 FILLER_47_219 ();
 sg13g2_decap_4 FILLER_47_226 ();
 sg13g2_fill_1 FILLER_47_279 ();
 sg13g2_fill_2 FILLER_47_315 ();
 sg13g2_decap_4 FILLER_47_325 ();
 sg13g2_fill_2 FILLER_47_333 ();
 sg13g2_fill_2 FILLER_47_366 ();
 sg13g2_fill_2 FILLER_47_376 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_fill_2 FILLER_48_49 ();
 sg13g2_fill_1 FILLER_48_61 ();
 sg13g2_fill_2 FILLER_48_69 ();
 sg13g2_fill_1 FILLER_48_71 ();
 sg13g2_fill_2 FILLER_48_95 ();
 sg13g2_fill_1 FILLER_48_122 ();
 sg13g2_fill_1 FILLER_48_129 ();
 sg13g2_fill_1 FILLER_48_135 ();
 sg13g2_fill_2 FILLER_48_150 ();
 sg13g2_fill_2 FILLER_48_161 ();
 sg13g2_fill_1 FILLER_48_163 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_fill_1 FILLER_48_200 ();
 sg13g2_fill_2 FILLER_48_307 ();
 sg13g2_decap_8 FILLER_48_333 ();
 sg13g2_fill_2 FILLER_48_343 ();
 sg13g2_fill_1 FILLER_48_350 ();
 sg13g2_fill_2 FILLER_48_366 ();
 sg13g2_fill_1 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_fill_2 FILLER_49_42 ();
 sg13g2_fill_1 FILLER_49_44 ();
 sg13g2_fill_2 FILLER_49_57 ();
 sg13g2_fill_2 FILLER_49_76 ();
 sg13g2_fill_1 FILLER_49_78 ();
 sg13g2_decap_4 FILLER_49_87 ();
 sg13g2_fill_2 FILLER_49_91 ();
 sg13g2_fill_2 FILLER_49_111 ();
 sg13g2_fill_1 FILLER_49_113 ();
 sg13g2_fill_2 FILLER_49_120 ();
 sg13g2_fill_1 FILLER_49_122 ();
 sg13g2_fill_2 FILLER_49_129 ();
 sg13g2_fill_1 FILLER_49_131 ();
 sg13g2_decap_8 FILLER_49_141 ();
 sg13g2_fill_1 FILLER_49_148 ();
 sg13g2_decap_8 FILLER_49_156 ();
 sg13g2_decap_8 FILLER_49_163 ();
 sg13g2_fill_2 FILLER_49_170 ();
 sg13g2_decap_4 FILLER_49_178 ();
 sg13g2_fill_2 FILLER_49_192 ();
 sg13g2_fill_1 FILLER_49_194 ();
 sg13g2_fill_1 FILLER_49_200 ();
 sg13g2_decap_8 FILLER_49_213 ();
 sg13g2_fill_2 FILLER_49_260 ();
 sg13g2_fill_1 FILLER_49_270 ();
 sg13g2_decap_8 FILLER_49_347 ();
 sg13g2_fill_2 FILLER_49_354 ();
 sg13g2_fill_1 FILLER_49_365 ();
 sg13g2_fill_2 FILLER_49_392 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_4 FILLER_50_64 ();
 sg13g2_fill_2 FILLER_50_68 ();
 sg13g2_decap_8 FILLER_50_85 ();
 sg13g2_fill_2 FILLER_50_92 ();
 sg13g2_fill_1 FILLER_50_94 ();
 sg13g2_fill_2 FILLER_50_109 ();
 sg13g2_fill_1 FILLER_50_111 ();
 sg13g2_fill_2 FILLER_50_123 ();
 sg13g2_fill_2 FILLER_50_133 ();
 sg13g2_fill_2 FILLER_50_151 ();
 sg13g2_decap_4 FILLER_50_158 ();
 sg13g2_fill_1 FILLER_50_166 ();
 sg13g2_fill_2 FILLER_50_178 ();
 sg13g2_fill_1 FILLER_50_180 ();
 sg13g2_fill_2 FILLER_50_200 ();
 sg13g2_fill_1 FILLER_50_286 ();
 sg13g2_fill_2 FILLER_50_313 ();
 sg13g2_fill_1 FILLER_50_325 ();
 sg13g2_fill_2 FILLER_50_352 ();
 sg13g2_fill_1 FILLER_50_354 ();
 sg13g2_fill_1 FILLER_50_385 ();
 sg13g2_fill_1 FILLER_50_390 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_fill_2 FILLER_51_70 ();
 sg13g2_fill_2 FILLER_51_119 ();
 sg13g2_fill_1 FILLER_51_121 ();
 sg13g2_fill_1 FILLER_51_134 ();
 sg13g2_fill_1 FILLER_51_145 ();
 sg13g2_fill_1 FILLER_51_167 ();
 sg13g2_fill_2 FILLER_51_327 ();
 sg13g2_decap_8 FILLER_51_355 ();
 sg13g2_fill_2 FILLER_51_362 ();
 sg13g2_fill_1 FILLER_51_364 ();
 sg13g2_fill_2 FILLER_51_383 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_4 FILLER_52_49 ();
 sg13g2_fill_1 FILLER_52_53 ();
 sg13g2_fill_2 FILLER_52_59 ();
 sg13g2_fill_1 FILLER_52_68 ();
 sg13g2_fill_1 FILLER_52_83 ();
 sg13g2_fill_2 FILLER_52_105 ();
 sg13g2_fill_1 FILLER_52_107 ();
 sg13g2_fill_2 FILLER_52_144 ();
 sg13g2_decap_8 FILLER_52_154 ();
 sg13g2_decap_8 FILLER_52_161 ();
 sg13g2_fill_2 FILLER_52_176 ();
 sg13g2_fill_2 FILLER_52_185 ();
 sg13g2_fill_1 FILLER_52_187 ();
 sg13g2_fill_1 FILLER_52_280 ();
 sg13g2_decap_8 FILLER_52_319 ();
 sg13g2_decap_8 FILLER_52_326 ();
 sg13g2_decap_4 FILLER_52_333 ();
 sg13g2_fill_2 FILLER_52_337 ();
 sg13g2_fill_2 FILLER_52_347 ();
 sg13g2_fill_1 FILLER_52_349 ();
 sg13g2_decap_8 FILLER_52_357 ();
 sg13g2_decap_8 FILLER_52_364 ();
 sg13g2_decap_8 FILLER_52_371 ();
 sg13g2_decap_8 FILLER_52_378 ();
 sg13g2_fill_1 FILLER_52_385 ();
 sg13g2_fill_2 FILLER_52_407 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_4 FILLER_53_42 ();
 sg13g2_fill_1 FILLER_53_46 ();
 sg13g2_decap_4 FILLER_53_78 ();
 sg13g2_fill_1 FILLER_53_103 ();
 sg13g2_fill_1 FILLER_53_109 ();
 sg13g2_fill_1 FILLER_53_124 ();
 sg13g2_decap_8 FILLER_53_130 ();
 sg13g2_decap_4 FILLER_53_137 ();
 sg13g2_fill_1 FILLER_53_146 ();
 sg13g2_fill_2 FILLER_53_235 ();
 sg13g2_fill_1 FILLER_53_237 ();
 sg13g2_fill_1 FILLER_53_247 ();
 sg13g2_fill_2 FILLER_53_265 ();
 sg13g2_decap_8 FILLER_53_309 ();
 sg13g2_decap_4 FILLER_53_342 ();
 sg13g2_decap_8 FILLER_53_367 ();
 sg13g2_decap_8 FILLER_53_374 ();
 sg13g2_decap_8 FILLER_53_381 ();
 sg13g2_decap_8 FILLER_53_388 ();
 sg13g2_decap_8 FILLER_53_395 ();
 sg13g2_decap_8 FILLER_53_402 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_fill_2 FILLER_54_35 ();
 sg13g2_fill_1 FILLER_54_37 ();
 sg13g2_fill_2 FILLER_54_89 ();
 sg13g2_fill_1 FILLER_54_91 ();
 sg13g2_fill_2 FILLER_54_97 ();
 sg13g2_decap_4 FILLER_54_104 ();
 sg13g2_fill_1 FILLER_54_108 ();
 sg13g2_decap_4 FILLER_54_124 ();
 sg13g2_fill_1 FILLER_54_133 ();
 sg13g2_fill_1 FILLER_54_159 ();
 sg13g2_fill_2 FILLER_54_184 ();
 sg13g2_decap_4 FILLER_54_218 ();
 sg13g2_fill_1 FILLER_54_230 ();
 sg13g2_decap_4 FILLER_54_252 ();
 sg13g2_fill_2 FILLER_54_256 ();
 sg13g2_decap_8 FILLER_54_261 ();
 sg13g2_fill_2 FILLER_54_268 ();
 sg13g2_fill_1 FILLER_54_270 ();
 sg13g2_decap_4 FILLER_54_285 ();
 sg13g2_fill_2 FILLER_54_334 ();
 sg13g2_fill_1 FILLER_54_336 ();
 sg13g2_fill_2 FILLER_54_375 ();
 sg13g2_fill_1 FILLER_54_377 ();
 sg13g2_decap_4 FILLER_54_404 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_fill_2 FILLER_55_42 ();
 sg13g2_fill_1 FILLER_55_66 ();
 sg13g2_fill_1 FILLER_55_74 ();
 sg13g2_decap_8 FILLER_55_87 ();
 sg13g2_decap_4 FILLER_55_94 ();
 sg13g2_fill_1 FILLER_55_104 ();
 sg13g2_fill_1 FILLER_55_128 ();
 sg13g2_decap_4 FILLER_55_144 ();
 sg13g2_decap_8 FILLER_55_172 ();
 sg13g2_decap_8 FILLER_55_179 ();
 sg13g2_fill_2 FILLER_55_186 ();
 sg13g2_fill_1 FILLER_55_188 ();
 sg13g2_decap_8 FILLER_55_202 ();
 sg13g2_fill_1 FILLER_55_209 ();
 sg13g2_decap_4 FILLER_55_218 ();
 sg13g2_fill_2 FILLER_55_222 ();
 sg13g2_fill_2 FILLER_55_229 ();
 sg13g2_decap_8 FILLER_55_244 ();
 sg13g2_decap_8 FILLER_55_256 ();
 sg13g2_decap_4 FILLER_55_268 ();
 sg13g2_decap_8 FILLER_55_284 ();
 sg13g2_fill_2 FILLER_55_299 ();
 sg13g2_fill_1 FILLER_55_301 ();
 sg13g2_fill_2 FILLER_55_337 ();
 sg13g2_fill_2 FILLER_55_354 ();
 sg13g2_fill_1 FILLER_55_356 ();
 sg13g2_fill_2 FILLER_55_379 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_4 FILLER_56_49 ();
 sg13g2_decap_4 FILLER_56_73 ();
 sg13g2_fill_1 FILLER_56_94 ();
 sg13g2_fill_2 FILLER_56_123 ();
 sg13g2_fill_2 FILLER_56_163 ();
 sg13g2_decap_8 FILLER_56_170 ();
 sg13g2_decap_4 FILLER_56_177 ();
 sg13g2_decap_4 FILLER_56_215 ();
 sg13g2_fill_1 FILLER_56_219 ();
 sg13g2_fill_2 FILLER_56_311 ();
 sg13g2_fill_1 FILLER_56_313 ();
 sg13g2_decap_4 FILLER_56_318 ();
 sg13g2_decap_8 FILLER_56_326 ();
 sg13g2_fill_2 FILLER_56_362 ();
 sg13g2_fill_1 FILLER_56_364 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_fill_1 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_58 ();
 sg13g2_fill_1 FILLER_57_65 ();
 sg13g2_fill_2 FILLER_57_70 ();
 sg13g2_fill_1 FILLER_57_72 ();
 sg13g2_decap_8 FILLER_57_89 ();
 sg13g2_fill_1 FILLER_57_96 ();
 sg13g2_decap_8 FILLER_57_126 ();
 sg13g2_decap_8 FILLER_57_151 ();
 sg13g2_decap_4 FILLER_57_158 ();
 sg13g2_fill_1 FILLER_57_177 ();
 sg13g2_decap_8 FILLER_57_181 ();
 sg13g2_fill_2 FILLER_57_188 ();
 sg13g2_decap_8 FILLER_57_283 ();
 sg13g2_decap_8 FILLER_57_290 ();
 sg13g2_fill_2 FILLER_57_297 ();
 sg13g2_fill_1 FILLER_57_299 ();
 sg13g2_decap_8 FILLER_57_304 ();
 sg13g2_fill_2 FILLER_57_311 ();
 sg13g2_fill_1 FILLER_57_313 ();
 sg13g2_fill_1 FILLER_57_349 ();
 sg13g2_fill_2 FILLER_57_406 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_4 FILLER_58_49 ();
 sg13g2_fill_1 FILLER_58_53 ();
 sg13g2_fill_2 FILLER_58_66 ();
 sg13g2_fill_1 FILLER_58_68 ();
 sg13g2_decap_4 FILLER_58_101 ();
 sg13g2_fill_2 FILLER_58_105 ();
 sg13g2_decap_4 FILLER_58_120 ();
 sg13g2_fill_1 FILLER_58_124 ();
 sg13g2_decap_4 FILLER_58_131 ();
 sg13g2_fill_1 FILLER_58_135 ();
 sg13g2_decap_8 FILLER_58_141 ();
 sg13g2_fill_1 FILLER_58_148 ();
 sg13g2_fill_2 FILLER_58_155 ();
 sg13g2_fill_1 FILLER_58_157 ();
 sg13g2_fill_1 FILLER_58_171 ();
 sg13g2_fill_1 FILLER_58_188 ();
 sg13g2_fill_2 FILLER_58_217 ();
 sg13g2_fill_2 FILLER_58_241 ();
 sg13g2_decap_8 FILLER_58_280 ();
 sg13g2_decap_4 FILLER_58_287 ();
 sg13g2_decap_8 FILLER_58_313 ();
 sg13g2_decap_4 FILLER_58_320 ();
 sg13g2_fill_1 FILLER_58_324 ();
 sg13g2_decap_4 FILLER_58_329 ();
 sg13g2_decap_8 FILLER_58_337 ();
 sg13g2_fill_2 FILLER_58_354 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_4 FILLER_59_42 ();
 sg13g2_fill_2 FILLER_59_125 ();
 sg13g2_fill_1 FILLER_59_127 ();
 sg13g2_fill_2 FILLER_59_141 ();
 sg13g2_fill_1 FILLER_59_143 ();
 sg13g2_fill_2 FILLER_59_152 ();
 sg13g2_fill_1 FILLER_59_162 ();
 sg13g2_fill_1 FILLER_59_219 ();
 sg13g2_fill_1 FILLER_59_233 ();
 sg13g2_fill_1 FILLER_59_255 ();
 sg13g2_fill_2 FILLER_59_263 ();
 sg13g2_decap_8 FILLER_59_339 ();
 sg13g2_decap_4 FILLER_59_346 ();
 sg13g2_fill_2 FILLER_59_350 ();
 sg13g2_fill_2 FILLER_59_378 ();
 sg13g2_fill_1 FILLER_59_380 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_fill_1 FILLER_60_56 ();
 sg13g2_fill_2 FILLER_60_103 ();
 sg13g2_fill_2 FILLER_60_120 ();
 sg13g2_fill_1 FILLER_60_134 ();
 sg13g2_fill_1 FILLER_60_178 ();
 sg13g2_fill_2 FILLER_60_218 ();
 sg13g2_decap_8 FILLER_60_239 ();
 sg13g2_fill_1 FILLER_60_246 ();
 sg13g2_decap_8 FILLER_60_250 ();
 sg13g2_fill_1 FILLER_60_294 ();
 sg13g2_decap_4 FILLER_60_318 ();
 sg13g2_fill_1 FILLER_60_322 ();
 sg13g2_fill_1 FILLER_60_337 ();
 sg13g2_decap_8 FILLER_60_351 ();
 sg13g2_fill_1 FILLER_60_358 ();
 sg13g2_fill_2 FILLER_60_367 ();
 sg13g2_fill_1 FILLER_60_369 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_fill_1 FILLER_61_77 ();
 sg13g2_fill_2 FILLER_61_95 ();
 sg13g2_fill_1 FILLER_61_97 ();
 sg13g2_fill_2 FILLER_61_106 ();
 sg13g2_decap_4 FILLER_61_128 ();
 sg13g2_fill_1 FILLER_61_132 ();
 sg13g2_fill_2 FILLER_61_138 ();
 sg13g2_fill_1 FILLER_61_140 ();
 sg13g2_fill_2 FILLER_61_167 ();
 sg13g2_decap_4 FILLER_61_200 ();
 sg13g2_fill_2 FILLER_61_224 ();
 sg13g2_fill_1 FILLER_61_240 ();
 sg13g2_decap_8 FILLER_61_248 ();
 sg13g2_decap_8 FILLER_61_255 ();
 sg13g2_fill_2 FILLER_61_262 ();
 sg13g2_fill_2 FILLER_61_301 ();
 sg13g2_fill_1 FILLER_61_339 ();
 sg13g2_fill_1 FILLER_61_359 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_fill_2 FILLER_62_109 ();
 sg13g2_fill_1 FILLER_62_111 ();
 sg13g2_decap_8 FILLER_62_117 ();
 sg13g2_decap_8 FILLER_62_124 ();
 sg13g2_decap_8 FILLER_62_131 ();
 sg13g2_decap_8 FILLER_62_149 ();
 sg13g2_fill_2 FILLER_62_156 ();
 sg13g2_decap_8 FILLER_62_175 ();
 sg13g2_decap_4 FILLER_62_182 ();
 sg13g2_fill_2 FILLER_62_211 ();
 sg13g2_fill_2 FILLER_62_218 ();
 sg13g2_fill_1 FILLER_62_235 ();
 sg13g2_fill_1 FILLER_62_244 ();
 sg13g2_decap_4 FILLER_62_258 ();
 sg13g2_fill_1 FILLER_62_262 ();
 sg13g2_fill_2 FILLER_62_267 ();
 sg13g2_decap_8 FILLER_62_273 ();
 sg13g2_fill_1 FILLER_62_280 ();
 sg13g2_fill_1 FILLER_62_291 ();
 sg13g2_decap_8 FILLER_62_314 ();
 sg13g2_decap_8 FILLER_62_321 ();
 sg13g2_fill_2 FILLER_62_337 ();
 sg13g2_fill_2 FILLER_62_344 ();
 sg13g2_fill_1 FILLER_62_346 ();
 sg13g2_fill_2 FILLER_62_363 ();
 sg13g2_fill_1 FILLER_62_365 ();
 sg13g2_fill_1 FILLER_62_392 ();
 sg13g2_fill_2 FILLER_62_407 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_fill_2 FILLER_63_126 ();
 sg13g2_fill_1 FILLER_63_128 ();
 sg13g2_fill_2 FILLER_63_138 ();
 sg13g2_fill_1 FILLER_63_140 ();
 sg13g2_decap_4 FILLER_63_177 ();
 sg13g2_fill_1 FILLER_63_181 ();
 sg13g2_decap_8 FILLER_63_187 ();
 sg13g2_decap_8 FILLER_63_194 ();
 sg13g2_fill_2 FILLER_63_201 ();
 sg13g2_fill_1 FILLER_63_203 ();
 sg13g2_fill_2 FILLER_63_283 ();
 sg13g2_decap_8 FILLER_63_305 ();
 sg13g2_decap_8 FILLER_63_312 ();
 sg13g2_fill_2 FILLER_63_319 ();
 sg13g2_fill_1 FILLER_63_321 ();
 sg13g2_fill_2 FILLER_63_326 ();
 sg13g2_fill_2 FILLER_63_342 ();
 sg13g2_fill_1 FILLER_63_344 ();
 sg13g2_fill_2 FILLER_63_406 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_fill_2 FILLER_64_112 ();
 sg13g2_decap_4 FILLER_64_197 ();
 sg13g2_fill_1 FILLER_64_221 ();
 sg13g2_fill_2 FILLER_64_259 ();
 sg13g2_fill_2 FILLER_64_298 ();
 sg13g2_decap_8 FILLER_64_305 ();
 sg13g2_fill_2 FILLER_64_316 ();
 sg13g2_fill_1 FILLER_64_318 ();
 sg13g2_fill_2 FILLER_64_324 ();
 sg13g2_fill_1 FILLER_64_326 ();
 sg13g2_fill_2 FILLER_64_343 ();
 sg13g2_fill_1 FILLER_64_345 ();
 sg13g2_fill_1 FILLER_64_365 ();
 sg13g2_fill_2 FILLER_64_374 ();
 sg13g2_fill_1 FILLER_64_376 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_fill_2 FILLER_65_105 ();
 sg13g2_decap_4 FILLER_65_244 ();
 sg13g2_decap_8 FILLER_65_255 ();
 sg13g2_fill_2 FILLER_65_290 ();
 sg13g2_fill_2 FILLER_65_310 ();
 sg13g2_fill_1 FILLER_65_312 ();
 sg13g2_fill_2 FILLER_65_327 ();
 sg13g2_fill_1 FILLER_65_329 ();
 sg13g2_fill_1 FILLER_65_359 ();
 sg13g2_fill_1 FILLER_65_382 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_fill_2 FILLER_66_98 ();
 sg13g2_fill_1 FILLER_66_100 ();
 sg13g2_fill_1 FILLER_66_146 ();
 sg13g2_fill_2 FILLER_66_199 ();
 sg13g2_decap_8 FILLER_66_217 ();
 sg13g2_fill_1 FILLER_66_229 ();
 sg13g2_decap_4 FILLER_66_235 ();
 sg13g2_fill_1 FILLER_66_239 ();
 sg13g2_decap_4 FILLER_66_261 ();
 sg13g2_decap_8 FILLER_66_305 ();
 sg13g2_fill_1 FILLER_66_347 ();
 sg13g2_fill_2 FILLER_66_379 ();
 sg13g2_fill_1 FILLER_66_381 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_fill_1 FILLER_67_112 ();
 sg13g2_fill_2 FILLER_67_148 ();
 sg13g2_decap_4 FILLER_67_181 ();
 sg13g2_fill_2 FILLER_67_207 ();
 sg13g2_fill_2 FILLER_67_248 ();
 sg13g2_decap_8 FILLER_67_259 ();
 sg13g2_fill_2 FILLER_67_266 ();
 sg13g2_fill_1 FILLER_67_286 ();
 sg13g2_decap_8 FILLER_67_299 ();
 sg13g2_decap_8 FILLER_67_306 ();
 sg13g2_fill_2 FILLER_67_313 ();
 sg13g2_fill_1 FILLER_67_335 ();
 sg13g2_fill_1 FILLER_67_345 ();
 sg13g2_fill_2 FILLER_67_372 ();
 sg13g2_fill_1 FILLER_67_379 ();
 sg13g2_fill_1 FILLER_67_395 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_4 FILLER_68_112 ();
 sg13g2_fill_1 FILLER_68_116 ();
 sg13g2_fill_2 FILLER_68_144 ();
 sg13g2_fill_2 FILLER_68_203 ();
 sg13g2_fill_2 FILLER_68_222 ();
 sg13g2_fill_2 FILLER_68_244 ();
 sg13g2_fill_1 FILLER_68_246 ();
 sg13g2_fill_1 FILLER_68_263 ();
 sg13g2_fill_1 FILLER_68_294 ();
 sg13g2_decap_8 FILLER_68_311 ();
 sg13g2_fill_2 FILLER_68_327 ();
 sg13g2_fill_1 FILLER_68_329 ();
 sg13g2_fill_2 FILLER_68_348 ();
 sg13g2_fill_2 FILLER_68_375 ();
 sg13g2_fill_1 FILLER_68_391 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_fill_2 FILLER_69_119 ();
 sg13g2_fill_1 FILLER_69_121 ();
 sg13g2_fill_1 FILLER_69_133 ();
 sg13g2_fill_2 FILLER_69_196 ();
 sg13g2_fill_1 FILLER_69_198 ();
 sg13g2_fill_2 FILLER_69_208 ();
 sg13g2_fill_1 FILLER_69_210 ();
 sg13g2_fill_1 FILLER_69_223 ();
 sg13g2_fill_2 FILLER_69_234 ();
 sg13g2_fill_1 FILLER_69_252 ();
 sg13g2_fill_1 FILLER_69_274 ();
 sg13g2_fill_1 FILLER_69_285 ();
 sg13g2_fill_1 FILLER_69_343 ();
 sg13g2_fill_2 FILLER_69_380 ();
 sg13g2_fill_1 FILLER_69_382 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_4 FILLER_70_119 ();
 sg13g2_fill_1 FILLER_70_123 ();
 sg13g2_fill_2 FILLER_70_155 ();
 sg13g2_fill_1 FILLER_70_157 ();
 sg13g2_fill_2 FILLER_70_286 ();
 sg13g2_fill_2 FILLER_70_293 ();
 sg13g2_fill_1 FILLER_70_310 ();
 sg13g2_fill_2 FILLER_70_316 ();
 sg13g2_fill_2 FILLER_70_358 ();
 sg13g2_fill_1 FILLER_70_370 ();
 sg13g2_fill_2 FILLER_70_376 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_4 FILLER_71_119 ();
 sg13g2_fill_1 FILLER_71_123 ();
 sg13g2_fill_2 FILLER_71_138 ();
 sg13g2_fill_2 FILLER_71_176 ();
 sg13g2_fill_1 FILLER_71_183 ();
 sg13g2_fill_2 FILLER_71_203 ();
 sg13g2_fill_1 FILLER_71_205 ();
 sg13g2_decap_4 FILLER_71_275 ();
 sg13g2_fill_1 FILLER_71_279 ();
 sg13g2_decap_4 FILLER_71_299 ();
 sg13g2_fill_2 FILLER_71_330 ();
 sg13g2_fill_1 FILLER_71_344 ();
 sg13g2_fill_1 FILLER_71_399 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_fill_1 FILLER_72_119 ();
 sg13g2_fill_2 FILLER_72_194 ();
 sg13g2_fill_1 FILLER_72_206 ();
 sg13g2_decap_8 FILLER_72_289 ();
 sg13g2_decap_8 FILLER_72_296 ();
 sg13g2_fill_1 FILLER_72_340 ();
 sg13g2_fill_2 FILLER_72_363 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_4 FILLER_73_112 ();
 sg13g2_fill_1 FILLER_73_175 ();
 sg13g2_decap_8 FILLER_73_302 ();
 sg13g2_decap_4 FILLER_73_309 ();
 sg13g2_fill_1 FILLER_73_313 ();
 sg13g2_fill_1 FILLER_73_324 ();
 sg13g2_fill_2 FILLER_73_398 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_fill_1 FILLER_74_112 ();
 sg13g2_fill_2 FILLER_74_161 ();
 sg13g2_fill_1 FILLER_74_229 ();
 sg13g2_fill_2 FILLER_74_243 ();
 sg13g2_fill_2 FILLER_74_298 ();
 sg13g2_fill_1 FILLER_74_300 ();
 sg13g2_fill_1 FILLER_74_306 ();
 sg13g2_fill_2 FILLER_74_323 ();
 sg13g2_fill_1 FILLER_74_330 ();
 sg13g2_fill_2 FILLER_74_346 ();
 sg13g2_fill_1 FILLER_74_348 ();
 sg13g2_fill_1 FILLER_74_362 ();
 sg13g2_fill_2 FILLER_74_391 ();
 sg13g2_fill_1 FILLER_74_393 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_4 FILLER_75_105 ();
 sg13g2_fill_2 FILLER_75_109 ();
 sg13g2_fill_1 FILLER_75_164 ();
 sg13g2_fill_2 FILLER_75_184 ();
 sg13g2_fill_2 FILLER_75_202 ();
 sg13g2_fill_2 FILLER_75_272 ();
 sg13g2_fill_2 FILLER_75_283 ();
 sg13g2_fill_2 FILLER_75_311 ();
 sg13g2_fill_2 FILLER_75_356 ();
 sg13g2_fill_1 FILLER_75_358 ();
 sg13g2_fill_2 FILLER_75_388 ();
 sg13g2_fill_1 FILLER_75_390 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_fill_1 FILLER_76_119 ();
 sg13g2_fill_2 FILLER_76_160 ();
 sg13g2_fill_2 FILLER_76_195 ();
 sg13g2_fill_2 FILLER_76_243 ();
 sg13g2_fill_1 FILLER_76_298 ();
 sg13g2_fill_1 FILLER_76_344 ();
 sg13g2_fill_2 FILLER_76_351 ();
 sg13g2_fill_1 FILLER_76_353 ();
 sg13g2_fill_1 FILLER_76_361 ();
 sg13g2_decap_8 FILLER_76_393 ();
 sg13g2_decap_8 FILLER_76_400 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_fill_1 FILLER_77_112 ();
 sg13g2_fill_1 FILLER_77_198 ();
 sg13g2_decap_8 FILLER_77_325 ();
 sg13g2_fill_2 FILLER_77_332 ();
 sg13g2_fill_1 FILLER_77_334 ();
 sg13g2_fill_2 FILLER_77_342 ();
 sg13g2_decap_8 FILLER_77_397 ();
 sg13g2_decap_4 FILLER_77_404 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_4 FILLER_78_112 ();
 sg13g2_fill_1 FILLER_78_116 ();
 sg13g2_fill_2 FILLER_78_218 ();
 sg13g2_fill_1 FILLER_78_237 ();
 sg13g2_decap_8 FILLER_78_316 ();
 sg13g2_fill_2 FILLER_78_323 ();
 sg13g2_fill_2 FILLER_78_339 ();
 sg13g2_fill_1 FILLER_78_341 ();
 sg13g2_fill_1 FILLER_78_350 ();
 sg13g2_fill_1 FILLER_78_368 ();
 sg13g2_decap_8 FILLER_78_395 ();
 sg13g2_decap_8 FILLER_78_402 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_4 FILLER_79_119 ();
 sg13g2_fill_1 FILLER_79_123 ();
 sg13g2_fill_1 FILLER_79_168 ();
 sg13g2_fill_1 FILLER_79_221 ();
 sg13g2_fill_1 FILLER_79_275 ();
 sg13g2_decap_8 FILLER_79_394 ();
 sg13g2_decap_8 FILLER_79_401 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_fill_2 FILLER_80_132 ();
 sg13g2_fill_1 FILLER_80_134 ();
 sg13g2_fill_1 FILLER_80_224 ();
 sg13g2_fill_1 FILLER_80_264 ();
 sg13g2_fill_1 FILLER_80_306 ();
 sg13g2_decap_4 FILLER_80_332 ();
 sg13g2_decap_4 FILLER_80_340 ();
 sg13g2_fill_2 FILLER_80_348 ();
 sg13g2_decap_8 FILLER_80_392 ();
 sg13g2_decap_8 FILLER_80_399 ();
 sg13g2_fill_2 FILLER_80_406 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net10;
 assign uio_oe[1] = net11;
 assign uio_oe[2] = net72;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule

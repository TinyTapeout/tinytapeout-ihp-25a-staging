module tt_um_wokwi_414120248222232577 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire clknet_0_clk;
 wire \boxcar_filter[0] ;
 wire \boxcar_filter[1] ;
 wire \boxcar_filter[2] ;
 wire \boxcar_filter[3] ;
 wire \boxcar_filter[4] ;
 wire \boxcar_filter[5] ;
 wire \boxcar_filter[6] ;
 wire \boxcar_filter[7] ;
 wire \boxcar_filter[8] ;
 wire \boxcar_filter[9] ;
 wire \boxcar_storage[1][0] ;
 wire \boxcar_storage[1][1] ;
 wire \boxcar_storage[1][2] ;
 wire \boxcar_storage[1][3] ;
 wire \boxcar_storage[1][4] ;
 wire \boxcar_storage[1][5] ;
 wire \boxcar_storage[1][6] ;
 wire \boxcar_storage[1][7] ;
 wire \boxcar_storage[2][0] ;
 wire \boxcar_storage[2][1] ;
 wire \boxcar_storage[2][2] ;
 wire \boxcar_storage[2][3] ;
 wire \boxcar_storage[2][4] ;
 wire \boxcar_storage[2][5] ;
 wire \boxcar_storage[2][6] ;
 wire \boxcar_storage[2][7] ;
 wire \boxcar_storage[3][0] ;
 wire \boxcar_storage[3][1] ;
 wire \boxcar_storage[3][2] ;
 wire \boxcar_storage[3][3] ;
 wire \boxcar_storage[3][4] ;
 wire \boxcar_storage[3][5] ;
 wire \boxcar_storage[3][6] ;
 wire \boxcar_storage[3][7] ;
 wire \boxcar_storage[4][0] ;
 wire \boxcar_storage[4][1] ;
 wire \boxcar_storage[4][2] ;
 wire \boxcar_storage[4][3] ;
 wire \boxcar_storage[4][4] ;
 wire \boxcar_storage[4][5] ;
 wire \boxcar_storage[4][6] ;
 wire \boxcar_storage[4][7] ;
 wire bypass_B;
 wire filter_on;
 wire \inst_sine_A.phase[0] ;
 wire \inst_sine_A.phase[1] ;
 wire \inst_sine_A.phase[2] ;
 wire \inst_sine_A.phase[3] ;
 wire \inst_sine_A.phase[4] ;
 wire \inst_sine_A.phase[5] ;
 wire \inst_sine_A.phase[6] ;
 wire \inst_sine_A.phase[7] ;
 wire \inst_sine_A.sample[0] ;
 wire \inst_sine_A.sample[1] ;
 wire \inst_sine_A.sample[2] ;
 wire \inst_sine_A.sample[3] ;
 wire \inst_sine_A.sample[4] ;
 wire \inst_sine_A.sample[5] ;
 wire \inst_sine_A.sample[6] ;
 wire \inst_sine_B.phase[0] ;
 wire \inst_sine_B.phase[1] ;
 wire \inst_sine_B.phase[2] ;
 wire \inst_sine_B.phase[3] ;
 wire \inst_sine_B.phase[4] ;
 wire \inst_sine_B.phase[5] ;
 wire \inst_sine_B.phase[6] ;
 wire \inst_sine_B.phase[7] ;
 wire lowamp_B;
 wire \mixer_out[0] ;
 wire \mixer_out[1] ;
 wire \mixer_out[2] ;
 wire \mixer_out[3] ;
 wire \mixer_out[4] ;
 wire \mixer_out[5] ;
 wire \mixer_out[6] ;
 wire \mixer_out[7] ;
 wire \phase_incr_A[0] ;
 wire \phase_incr_A[1] ;
 wire \phase_incr_A[2] ;
 wire \phase_incr_A[3] ;
 wire \phase_incr_A[4] ;
 wire \phase_incr_A[5] ;
 wire \phase_incr_A[6] ;
 wire \phase_incr_B[0] ;
 wire \phase_incr_B[1] ;
 wire \phase_incr_B[2] ;
 wire \phase_incr_B[3] ;
 wire \phase_incr_B[4] ;
 wire \phase_incr_B[5] ;
 wire \product[10] ;
 wire \product[11] ;
 wire \product[12] ;
 wire \product[13] ;
 wire \product[14] ;
 wire \product[7] ;
 wire \product[8] ;
 wire \product[9] ;
 wire \sine_Areg[0] ;
 wire \sine_Areg[1] ;
 wire \sine_Areg[2] ;
 wire \sine_Areg[3] ;
 wire \sine_Areg[4] ;
 wire \sine_Areg[5] ;
 wire \sine_Areg[6] ;
 wire \sine_Areg[7] ;
 wire \sine_Breg[0] ;
 wire \sine_Breg[1] ;
 wire \sine_Breg[2] ;
 wire \sine_Breg[3] ;
 wire \sine_Breg[4] ;
 wire \sine_Breg[5] ;
 wire \sine_Breg[6] ;
 wire \sine_Breg[7] ;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net148;
 wire net149;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;

 sg13g2_inv_1 _0990_ (.Y(_0099_),
    .A(net259));
 sg13g2_inv_1 _0991_ (.Y(_0100_),
    .A(net251));
 sg13g2_inv_1 _0992_ (.Y(_0101_),
    .A(net189));
 sg13g2_inv_1 _0993_ (.Y(_0102_),
    .A(net161));
 sg13g2_inv_1 _0994_ (.Y(_0103_),
    .A(net179));
 sg13g2_inv_1 _0995_ (.Y(_0104_),
    .A(net164));
 sg13g2_inv_1 _0996_ (.Y(_0105_),
    .A(net201));
 sg13g2_xor2_1 _0997_ (.B(net157),
    .A(\inst_sine_A.phase[5] ),
    .X(_0106_));
 sg13g2_xnor2_1 _0998_ (.Y(_0107_),
    .A(\inst_sine_A.phase[5] ),
    .B(net157));
 sg13g2_xor2_1 _0999_ (.B(\inst_sine_A.phase[4] ),
    .A(net157),
    .X(_0108_));
 sg13g2_xnor2_1 _1000_ (.Y(_0109_),
    .A(net157),
    .B(\inst_sine_A.phase[4] ));
 sg13g2_xor2_1 _1001_ (.B(\inst_sine_A.phase[3] ),
    .A(net158),
    .X(_0110_));
 sg13g2_xnor2_1 _1002_ (.Y(_0111_),
    .A(net157),
    .B(\inst_sine_A.phase[3] ));
 sg13g2_xor2_1 _1003_ (.B(\inst_sine_A.phase[0] ),
    .A(net158),
    .X(_0112_));
 sg13g2_xnor2_1 _1004_ (.Y(_0113_),
    .A(net158),
    .B(\inst_sine_A.phase[0] ));
 sg13g2_xor2_1 _1005_ (.B(\inst_sine_A.phase[1] ),
    .A(net158),
    .X(_0114_));
 sg13g2_xnor2_1 _1006_ (.Y(_0115_),
    .A(net158),
    .B(\inst_sine_A.phase[1] ));
 sg13g2_nand2_2 _1007_ (.Y(_0116_),
    .A(_0112_),
    .B(_0114_));
 sg13g2_xor2_1 _1008_ (.B(\inst_sine_A.phase[2] ),
    .A(net157),
    .X(_0117_));
 sg13g2_xnor2_1 _1009_ (.Y(_0118_),
    .A(net158),
    .B(\inst_sine_A.phase[2] ));
 sg13g2_o21ai_1 _1010_ (.B1(_0116_),
    .Y(_0119_),
    .A1(_0112_),
    .A2(_0118_));
 sg13g2_nor2_1 _1011_ (.A(_0111_),
    .B(_0119_),
    .Y(_0120_));
 sg13g2_nand2_1 _1012_ (.Y(_0121_),
    .A(_0109_),
    .B(_0120_));
 sg13g2_nand2_1 _1013_ (.Y(_0122_),
    .A(_0114_),
    .B(_0117_));
 sg13g2_a21oi_2 _1014_ (.B1(net155),
    .Y(_0123_),
    .A2(_0117_),
    .A1(_0114_));
 sg13g2_nand2_1 _1015_ (.Y(_0124_),
    .A(net154),
    .B(_0112_));
 sg13g2_nand2_1 _1016_ (.Y(_0125_),
    .A(_0112_),
    .B(_0123_));
 sg13g2_o21ai_1 _1017_ (.B1(net155),
    .Y(_0126_),
    .A1(_0115_),
    .A2(net153));
 sg13g2_nand3_1 _1018_ (.B(_0125_),
    .C(_0126_),
    .A(_0108_),
    .Y(_0127_));
 sg13g2_a21oi_1 _1019_ (.A1(_0121_),
    .A2(_0127_),
    .Y(_0128_),
    .B1(_0107_));
 sg13g2_nand2_1 _1020_ (.Y(_0129_),
    .A(_0113_),
    .B(_0115_));
 sg13g2_o21ai_1 _1021_ (.B1(_0129_),
    .Y(_0130_),
    .A1(_0115_),
    .A2(net153));
 sg13g2_nand2_1 _1022_ (.Y(_0131_),
    .A(_0124_),
    .B(_0130_));
 sg13g2_nor2_1 _1023_ (.A(_0106_),
    .B(net156),
    .Y(_0132_));
 sg13g2_nand2_1 _1024_ (.Y(_0133_),
    .A(_0107_),
    .B(_0108_));
 sg13g2_nor2_1 _1025_ (.A(_0118_),
    .B(_0124_),
    .Y(_0134_));
 sg13g2_nor2_1 _1026_ (.A(_0133_),
    .B(_0134_),
    .Y(_0135_));
 sg13g2_o21ai_1 _1027_ (.B1(_0125_),
    .Y(_0136_),
    .A1(_0111_),
    .A2(_0112_));
 sg13g2_nand2_1 _1028_ (.Y(_0137_),
    .A(_0107_),
    .B(net156));
 sg13g2_inv_1 _1029_ (.Y(_0138_),
    .A(_0137_));
 sg13g2_a221oi_1 _1030_ (.B2(_0138_),
    .C1(_0128_),
    .B1(_0136_),
    .A1(_0131_),
    .Y(\inst_sine_A.sample[0] ),
    .A2(_0135_));
 sg13g2_mux2_1 _1031_ (.A0(net245),
    .A1(net275),
    .S(filter_on),
    .X(_0000_));
 sg13g2_mux2_1 _1032_ (.A0(net240),
    .A1(net270),
    .S(filter_on),
    .X(_0001_));
 sg13g2_mux2_1 _1033_ (.A0(net241),
    .A1(net264),
    .S(filter_on),
    .X(_0002_));
 sg13g2_mux2_1 _1034_ (.A0(net246),
    .A1(net278),
    .S(filter_on),
    .X(_0003_));
 sg13g2_mux2_1 _1035_ (.A0(\mixer_out[4] ),
    .A1(net266),
    .S(filter_on),
    .X(_0004_));
 sg13g2_mux2_1 _1036_ (.A0(\mixer_out[5] ),
    .A1(net260),
    .S(filter_on),
    .X(_0005_));
 sg13g2_mux2_1 _1037_ (.A0(net258),
    .A1(net287),
    .S(filter_on),
    .X(_0006_));
 sg13g2_mux2_1 _1038_ (.A0(\mixer_out[7] ),
    .A1(net249),
    .S(filter_on),
    .X(_0007_));
 sg13g2_nor2b_2 _1039_ (.A(net255),
    .B_N(net257),
    .Y(_0139_));
 sg13g2_nand2b_1 _1040_ (.Y(_0140_),
    .B(net257),
    .A_N(net255));
 sg13g2_xor2_1 _1041_ (.B(\inst_sine_B.phase[1] ),
    .A(net188),
    .X(_0141_));
 sg13g2_xnor2_1 _1042_ (.Y(_0142_),
    .A(net188),
    .B(\inst_sine_B.phase[1] ));
 sg13g2_xor2_1 _1043_ (.B(\inst_sine_B.phase[2] ),
    .A(net188),
    .X(_0143_));
 sg13g2_xnor2_1 _1044_ (.Y(_0144_),
    .A(net188),
    .B(\inst_sine_B.phase[2] ));
 sg13g2_nor2_1 _1045_ (.A(_0141_),
    .B(net152),
    .Y(_0145_));
 sg13g2_nand2_2 _1046_ (.Y(_0146_),
    .A(_0142_),
    .B(_0144_));
 sg13g2_xor2_1 _1047_ (.B(\inst_sine_B.phase[0] ),
    .A(net187),
    .X(_0147_));
 sg13g2_xnor2_1 _1048_ (.Y(_0148_),
    .A(net187),
    .B(\inst_sine_B.phase[0] ));
 sg13g2_nor2_1 _1049_ (.A(_0141_),
    .B(_0148_),
    .Y(_0149_));
 sg13g2_xnor2_1 _1050_ (.Y(_0150_),
    .A(\inst_sine_B.phase[1] ),
    .B(\inst_sine_B.phase[0] ));
 sg13g2_xor2_1 _1051_ (.B(\inst_sine_B.phase[0] ),
    .A(\inst_sine_B.phase[1] ),
    .X(_0151_));
 sg13g2_o21ai_1 _1052_ (.B1(_0146_),
    .Y(_0152_),
    .A1(_0144_),
    .A2(_0151_));
 sg13g2_nand2_1 _1053_ (.Y(_0153_),
    .A(_0144_),
    .B(_0148_));
 sg13g2_xor2_1 _1054_ (.B(\inst_sine_B.phase[3] ),
    .A(net188),
    .X(_0154_));
 sg13g2_xnor2_1 _1055_ (.Y(_0155_),
    .A(net188),
    .B(\inst_sine_B.phase[3] ));
 sg13g2_nand3_1 _1056_ (.B(_0153_),
    .C(net151),
    .A(_0152_),
    .Y(_0156_));
 sg13g2_xor2_1 _1057_ (.B(\inst_sine_B.phase[4] ),
    .A(net187),
    .X(_0157_));
 sg13g2_xnor2_1 _1058_ (.Y(_0158_),
    .A(net187),
    .B(\inst_sine_B.phase[4] ));
 sg13g2_nor2_2 _1059_ (.A(_0148_),
    .B(net151),
    .Y(_0159_));
 sg13g2_nor2_1 _1060_ (.A(_0157_),
    .B(_0159_),
    .Y(_0160_));
 sg13g2_xor2_1 _1061_ (.B(\inst_sine_B.phase[5] ),
    .A(net187),
    .X(_0161_));
 sg13g2_xnor2_1 _1062_ (.Y(_0162_),
    .A(net187),
    .B(\inst_sine_B.phase[5] ));
 sg13g2_nor2_1 _1063_ (.A(_0146_),
    .B(_0155_),
    .Y(_0163_));
 sg13g2_nand2_1 _1064_ (.Y(_0164_),
    .A(_0141_),
    .B(_0155_));
 sg13g2_nor2_1 _1065_ (.A(_0158_),
    .B(_0163_),
    .Y(_0165_));
 sg13g2_a221oi_1 _1066_ (.B2(_0165_),
    .C1(_0162_),
    .B1(_0164_),
    .A1(_0156_),
    .Y(_0166_),
    .A2(_0160_));
 sg13g2_nor2b_1 _1067_ (.A(_0149_),
    .B_N(_0153_),
    .Y(_0167_));
 sg13g2_nor2_1 _1068_ (.A(_0155_),
    .B(_0167_),
    .Y(_0168_));
 sg13g2_or2_1 _1069_ (.X(_0169_),
    .B(_0168_),
    .A(_0152_));
 sg13g2_nand2_1 _1070_ (.Y(_0170_),
    .A(_0157_),
    .B(_0162_));
 sg13g2_nor2_1 _1071_ (.A(_0163_),
    .B(_0170_),
    .Y(_0171_));
 sg13g2_nand2_2 _1072_ (.Y(_0172_),
    .A(_0158_),
    .B(_0162_));
 sg13g2_a21oi_1 _1073_ (.A1(_0150_),
    .A2(net151),
    .Y(_0173_),
    .B1(_0172_));
 sg13g2_a221oi_1 _1074_ (.B2(_0164_),
    .C1(_0166_),
    .B1(_0173_),
    .A1(_0169_),
    .Y(_0174_),
    .A2(_0171_));
 sg13g2_nand2_1 _1075_ (.Y(_0175_),
    .A(_0158_),
    .B(_0168_));
 sg13g2_o21ai_1 _1076_ (.B1(net150),
    .Y(_0176_),
    .A1(_0142_),
    .A2(net152));
 sg13g2_nand2_1 _1077_ (.Y(_0177_),
    .A(_0141_),
    .B(_0143_));
 sg13g2_a21oi_2 _1078_ (.B1(net150),
    .Y(_0178_),
    .A2(net152),
    .A1(_0141_));
 sg13g2_nand2_1 _1079_ (.Y(_0179_),
    .A(_0147_),
    .B(_0178_));
 sg13g2_nand3_1 _1080_ (.B(_0176_),
    .C(_0179_),
    .A(_0157_),
    .Y(_0180_));
 sg13g2_a21oi_1 _1081_ (.A1(_0175_),
    .A2(_0180_),
    .Y(_0181_),
    .B1(_0162_));
 sg13g2_nand2_1 _1082_ (.Y(_0182_),
    .A(_0142_),
    .B(_0148_));
 sg13g2_nor2_1 _1083_ (.A(_0149_),
    .B(_0159_),
    .Y(_0183_));
 sg13g2_nor2_1 _1084_ (.A(_0144_),
    .B(net151),
    .Y(_0184_));
 sg13g2_a221oi_1 _1085_ (.B2(_0183_),
    .C1(_0170_),
    .B1(_0177_),
    .A1(net152),
    .Y(_0185_),
    .A2(_0159_));
 sg13g2_nand2_1 _1086_ (.Y(_0186_),
    .A(_0148_),
    .B(net150));
 sg13g2_a21oi_1 _1087_ (.A1(_0179_),
    .A2(_0186_),
    .Y(_0187_),
    .B1(_0172_));
 sg13g2_nor3_2 _1088_ (.A(_0181_),
    .B(_0185_),
    .C(_0187_),
    .Y(_0188_));
 sg13g2_nand2_1 _1089_ (.Y(_0189_),
    .A(net268),
    .B(_0188_));
 sg13g2_xnor2_1 _1090_ (.Y(_0190_),
    .A(_0174_),
    .B(_0189_));
 sg13g2_nand2_1 _1091_ (.Y(_0191_),
    .A(net255),
    .B(net252));
 sg13g2_nor2_2 _1092_ (.A(net257),
    .B(net255),
    .Y(_0192_));
 sg13g2_or2_1 _1093_ (.X(_0193_),
    .B(net255),
    .A(net257));
 sg13g2_a22oi_1 _1094_ (.Y(_0194_),
    .B1(_0192_),
    .B2(_0188_),
    .A2(_0190_),
    .A1(_0139_));
 sg13g2_nand2_1 _1095_ (.Y(_0008_),
    .A(_0191_),
    .B(_0194_));
 sg13g2_nand3_1 _1096_ (.B(_0157_),
    .C(_0178_),
    .A(_0146_),
    .Y(_0195_));
 sg13g2_nand2_1 _1097_ (.Y(_0196_),
    .A(_0141_),
    .B(_0147_));
 sg13g2_nand2_1 _1098_ (.Y(_0197_),
    .A(net152),
    .B(_0196_));
 sg13g2_a21oi_1 _1099_ (.A1(_0182_),
    .A2(_0197_),
    .Y(_0198_),
    .B1(_0155_));
 sg13g2_a21oi_1 _1100_ (.A1(_0150_),
    .A2(_0155_),
    .Y(_0199_),
    .B1(_0198_));
 sg13g2_o21ai_1 _1101_ (.B1(_0195_),
    .Y(_0200_),
    .A1(_0157_),
    .A2(_0199_));
 sg13g2_nor2_1 _1102_ (.A(_0147_),
    .B(_0164_),
    .Y(_0201_));
 sg13g2_nor2_1 _1103_ (.A(_0149_),
    .B(_0201_),
    .Y(_0202_));
 sg13g2_xnor2_1 _1104_ (.Y(_0203_),
    .A(net152),
    .B(_0202_));
 sg13g2_a21oi_1 _1105_ (.A1(_0158_),
    .A2(_0203_),
    .Y(_0204_),
    .B1(_0161_));
 sg13g2_nor2_1 _1106_ (.A(net152),
    .B(net150),
    .Y(_0205_));
 sg13g2_nand2_1 _1107_ (.Y(_0206_),
    .A(_0144_),
    .B(_0151_));
 sg13g2_o21ai_1 _1108_ (.B1(_0206_),
    .Y(_0207_),
    .A1(_0201_),
    .A2(_0205_));
 sg13g2_nand3_1 _1109_ (.B(_0157_),
    .C(_0207_),
    .A(_0156_),
    .Y(_0208_));
 sg13g2_a22oi_1 _1110_ (.Y(_0209_),
    .B1(_0204_),
    .B2(_0208_),
    .A2(_0200_),
    .A1(_0161_));
 sg13g2_or2_1 _1111_ (.X(_0210_),
    .B(_0188_),
    .A(_0174_));
 sg13g2_nand2_1 _1112_ (.Y(_0211_),
    .A(net268),
    .B(_0210_));
 sg13g2_xnor2_1 _1113_ (.Y(_0212_),
    .A(_0209_),
    .B(_0211_));
 sg13g2_a22oi_1 _1114_ (.Y(_0213_),
    .B1(_0212_),
    .B2(_0139_),
    .A2(_0192_),
    .A1(_0190_));
 sg13g2_nand2_1 _1115_ (.Y(_0009_),
    .A(_0191_),
    .B(_0213_));
 sg13g2_nor2_1 _1116_ (.A(_0145_),
    .B(_0157_),
    .Y(_0214_));
 sg13g2_o21ai_1 _1117_ (.B1(_0179_),
    .Y(_0215_),
    .A1(_0144_),
    .A2(_0159_));
 sg13g2_nor3_1 _1118_ (.A(_0146_),
    .B(net150),
    .C(_0158_),
    .Y(_0216_));
 sg13g2_a21o_1 _1119_ (.A2(_0215_),
    .A1(_0214_),
    .B1(_0216_),
    .X(_0217_));
 sg13g2_nand2_1 _1120_ (.Y(_0218_),
    .A(_0196_),
    .B(_0205_));
 sg13g2_a21oi_1 _1121_ (.A1(_0141_),
    .A2(_0184_),
    .Y(_0219_),
    .B1(_0198_));
 sg13g2_a21oi_1 _1122_ (.A1(_0218_),
    .A2(_0219_),
    .Y(_0220_),
    .B1(_0170_));
 sg13g2_a21o_1 _1123_ (.A2(_0177_),
    .A1(_0167_),
    .B1(_0176_),
    .X(_0221_));
 sg13g2_a21oi_1 _1124_ (.A1(_0167_),
    .A2(_0178_),
    .Y(_0222_),
    .B1(_0172_));
 sg13g2_a221oi_1 _1125_ (.B2(_0222_),
    .C1(_0220_),
    .B1(_0221_),
    .A1(_0161_),
    .Y(_0223_),
    .A2(_0217_));
 sg13g2_or2_1 _1126_ (.X(_0224_),
    .B(_0210_),
    .A(_0209_));
 sg13g2_nand2_1 _1127_ (.Y(_0225_),
    .A(net268),
    .B(_0224_));
 sg13g2_xor2_1 _1128_ (.B(_0225_),
    .A(_0223_),
    .X(_0226_));
 sg13g2_a22oi_1 _1129_ (.Y(_0227_),
    .B1(_0192_),
    .B2(_0212_),
    .A2(net252),
    .A1(bypass_B));
 sg13g2_o21ai_1 _1130_ (.B1(net253),
    .Y(_0010_),
    .A1(_0140_),
    .A2(_0226_));
 sg13g2_o21ai_1 _1131_ (.B1(_0162_),
    .Y(_0228_),
    .A1(_0158_),
    .A2(_0178_));
 sg13g2_o21ai_1 _1132_ (.B1(_0218_),
    .Y(_0229_),
    .A1(_0158_),
    .A2(_0162_));
 sg13g2_a21oi_1 _1133_ (.A1(net152),
    .A2(net150),
    .Y(_0230_),
    .B1(_0229_));
 sg13g2_a221oi_1 _1134_ (.B2(_0184_),
    .C1(_0172_),
    .B1(_0182_),
    .A1(_0145_),
    .Y(_0231_),
    .A2(net150));
 sg13g2_a21oi_1 _1135_ (.A1(_0228_),
    .A2(_0230_),
    .Y(_0232_),
    .B1(_0231_));
 sg13g2_nor2_1 _1136_ (.A(_0223_),
    .B(_0224_),
    .Y(_0233_));
 sg13g2_nor2_1 _1137_ (.A(_0099_),
    .B(_0233_),
    .Y(_0234_));
 sg13g2_xor2_1 _1138_ (.B(_0234_),
    .A(_0232_),
    .X(_0235_));
 sg13g2_a22oi_1 _1139_ (.Y(_0236_),
    .B1(_0139_),
    .B2(_0235_),
    .A2(net252),
    .A1(net255));
 sg13g2_o21ai_1 _1140_ (.B1(_0236_),
    .Y(_0011_),
    .A1(_0193_),
    .A2(_0226_));
 sg13g2_a22oi_1 _1141_ (.Y(_0237_),
    .B1(_0214_),
    .B2(net150),
    .A2(_0178_),
    .A1(_0157_));
 sg13g2_nand2_1 _1142_ (.Y(_0238_),
    .A(_0161_),
    .B(_0218_));
 sg13g2_a21oi_1 _1143_ (.A1(_0237_),
    .A2(_0238_),
    .Y(_0239_),
    .B1(_0233_));
 sg13g2_and2_1 _1144_ (.A(_0099_),
    .B(_0237_),
    .X(_0240_));
 sg13g2_mux2_1 _1145_ (.A0(_0240_),
    .A1(net259),
    .S(_0239_),
    .X(_0241_));
 sg13g2_a22oi_1 _1146_ (.Y(_0242_),
    .B1(_0192_),
    .B2(_0235_),
    .A2(net252),
    .A1(net255));
 sg13g2_o21ai_1 _1147_ (.B1(_0242_),
    .Y(_0012_),
    .A1(_0140_),
    .A2(_0241_));
 sg13g2_xnor2_1 _1148_ (.Y(_0243_),
    .A(net259),
    .B(_0228_));
 sg13g2_nor2_1 _1149_ (.A(_0140_),
    .B(_0243_),
    .Y(_0244_));
 sg13g2_o21ai_1 _1150_ (.B1(_0191_),
    .Y(_0245_),
    .A1(_0193_),
    .A2(_0241_));
 sg13g2_or2_1 _1151_ (.X(_0013_),
    .B(_0245_),
    .A(_0244_));
 sg13g2_nand2_1 _1152_ (.Y(_0246_),
    .A(net251),
    .B(\inst_sine_A.sample[0] ));
 sg13g2_nor2_1 _1153_ (.A(_0114_),
    .B(net153),
    .Y(_0247_));
 sg13g2_nand2_2 _1154_ (.Y(_0248_),
    .A(_0115_),
    .B(_0118_));
 sg13g2_nor2_1 _1155_ (.A(net154),
    .B(_0248_),
    .Y(_0249_));
 sg13g2_nor2_2 _1156_ (.A(_0110_),
    .B(_0115_),
    .Y(_0250_));
 sg13g2_and2_1 _1157_ (.A(_0116_),
    .B(_0129_),
    .X(_0251_));
 sg13g2_nor2_1 _1158_ (.A(_0118_),
    .B(_0251_),
    .Y(_0252_));
 sg13g2_nor2_1 _1159_ (.A(_0113_),
    .B(_0248_),
    .Y(_0253_));
 sg13g2_o21ai_1 _1160_ (.B1(net155),
    .Y(_0254_),
    .A1(_0252_),
    .A2(_0253_));
 sg13g2_o21ai_1 _1161_ (.B1(_0108_),
    .Y(_0255_),
    .A1(_0249_),
    .A2(_0250_));
 sg13g2_a21o_1 _1162_ (.A2(_0254_),
    .A1(_0124_),
    .B1(_0108_),
    .X(_0256_));
 sg13g2_nand3_1 _1163_ (.B(_0255_),
    .C(_0256_),
    .A(_0106_),
    .Y(_0257_));
 sg13g2_nor3_1 _1164_ (.A(_0120_),
    .B(_0247_),
    .C(_0252_),
    .Y(_0258_));
 sg13g2_o21ai_1 _1165_ (.B1(_0132_),
    .Y(_0259_),
    .A1(_0249_),
    .A2(_0258_));
 sg13g2_nor2_1 _1166_ (.A(_0111_),
    .B(_0251_),
    .Y(_0260_));
 sg13g2_o21ai_1 _1167_ (.B1(_0138_),
    .Y(_0261_),
    .A1(_0250_),
    .A2(_0260_));
 sg13g2_nand3_1 _1168_ (.B(_0259_),
    .C(_0261_),
    .A(_0257_),
    .Y(_0262_));
 sg13g2_xnor2_1 _1169_ (.Y(\inst_sine_A.sample[1] ),
    .A(_0246_),
    .B(_0262_));
 sg13g2_nor2_1 _1170_ (.A(net156),
    .B(net155),
    .Y(_0263_));
 sg13g2_nand3_1 _1171_ (.B(_0123_),
    .C(_0248_),
    .A(_0108_),
    .Y(_0264_));
 sg13g2_nor2_1 _1172_ (.A(net155),
    .B(_0251_),
    .Y(_0265_));
 sg13g2_nand2_1 _1173_ (.Y(_0266_),
    .A(_0116_),
    .B(net153));
 sg13g2_a21oi_1 _1174_ (.A1(_0129_),
    .A2(_0266_),
    .Y(_0267_),
    .B1(net154));
 sg13g2_o21ai_1 _1175_ (.B1(net156),
    .Y(_0268_),
    .A1(_0265_),
    .A2(_0267_));
 sg13g2_a21oi_1 _1176_ (.A1(_0264_),
    .A2(_0268_),
    .Y(_0269_),
    .B1(_0107_));
 sg13g2_nor2_1 _1177_ (.A(net155),
    .B(_0122_),
    .Y(_0270_));
 sg13g2_a221oi_1 _1178_ (.B2(_0113_),
    .C1(net156),
    .B1(_0270_),
    .A1(_0118_),
    .Y(_0271_),
    .A2(_0265_));
 sg13g2_xnor2_1 _1179_ (.Y(_0272_),
    .A(_0116_),
    .B(net153));
 sg13g2_o21ai_1 _1180_ (.B1(_0272_),
    .Y(_0273_),
    .A1(_0112_),
    .A2(_0250_));
 sg13g2_nor3_1 _1181_ (.A(_0112_),
    .B(net153),
    .C(_0250_),
    .Y(_0274_));
 sg13g2_nor2_1 _1182_ (.A(_0108_),
    .B(_0274_),
    .Y(_0275_));
 sg13g2_a221oi_1 _1183_ (.B2(_0275_),
    .C1(_0106_),
    .B1(_0273_),
    .A1(_0254_),
    .Y(_0276_),
    .A2(_0271_));
 sg13g2_nor2_1 _1184_ (.A(_0269_),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_or2_1 _1185_ (.X(_0278_),
    .B(_0262_),
    .A(\inst_sine_A.sample[0] ));
 sg13g2_nand2_1 _1186_ (.Y(_0279_),
    .A(net251),
    .B(_0278_));
 sg13g2_xnor2_1 _1187_ (.Y(\inst_sine_A.sample[2] ),
    .A(_0277_),
    .B(_0279_));
 sg13g2_nor2_1 _1188_ (.A(_0277_),
    .B(_0278_),
    .Y(_0280_));
 sg13g2_nor2_1 _1189_ (.A(_0100_),
    .B(_0280_),
    .Y(_0281_));
 sg13g2_nand2_1 _1190_ (.Y(_0282_),
    .A(net154),
    .B(_0272_));
 sg13g2_o21ai_1 _1191_ (.B1(_0282_),
    .Y(_0283_),
    .A1(net154),
    .A2(_0118_));
 sg13g2_a22oi_1 _1192_ (.Y(_0284_),
    .B1(_0283_),
    .B2(net156),
    .A2(_0263_),
    .A1(_0247_));
 sg13g2_nand2_1 _1193_ (.Y(_0285_),
    .A(_0119_),
    .B(_0122_));
 sg13g2_nand3_1 _1194_ (.B(_0119_),
    .C(_0122_),
    .A(net155),
    .Y(_0286_));
 sg13g2_a21oi_1 _1195_ (.A1(_0126_),
    .A2(_0285_),
    .Y(_0287_),
    .B1(_0137_));
 sg13g2_nand3_1 _1196_ (.B(_0116_),
    .C(_0118_),
    .A(net154),
    .Y(_0288_));
 sg13g2_inv_1 _1197_ (.Y(_0289_),
    .A(_0288_));
 sg13g2_nor4_1 _1198_ (.A(_0133_),
    .B(_0267_),
    .C(_0270_),
    .D(_0289_),
    .Y(_0290_));
 sg13g2_a221oi_1 _1199_ (.B2(_0287_),
    .C1(_0290_),
    .B1(_0286_),
    .A1(_0106_),
    .Y(_0291_),
    .A2(_0284_));
 sg13g2_xnor2_1 _1200_ (.Y(\inst_sine_A.sample[3] ),
    .A(_0281_),
    .B(_0291_));
 sg13g2_o21ai_1 _1201_ (.B1(_0107_),
    .Y(_0292_),
    .A1(net156),
    .A2(_0123_));
 sg13g2_nand2_1 _1202_ (.Y(_0293_),
    .A(net156),
    .B(_0288_));
 sg13g2_a22oi_1 _1203_ (.Y(_0294_),
    .B1(_0293_),
    .B2(_0106_),
    .A2(net153),
    .A1(net155));
 sg13g2_nand3_1 _1204_ (.B(net153),
    .C(_0129_),
    .A(net154),
    .Y(_0295_));
 sg13g2_nor2_1 _1205_ (.A(_0137_),
    .B(_0249_),
    .Y(_0296_));
 sg13g2_a22oi_1 _1206_ (.Y(_0297_),
    .B1(_0295_),
    .B2(_0296_),
    .A2(_0294_),
    .A1(_0292_));
 sg13g2_a21oi_1 _1207_ (.A1(_0280_),
    .A2(_0291_),
    .Y(_0298_),
    .B1(_0100_));
 sg13g2_xor2_1 _1208_ (.B(_0298_),
    .A(_0297_),
    .X(\inst_sine_A.sample[4] ));
 sg13g2_nand2_1 _1209_ (.Y(_0299_),
    .A(_0106_),
    .B(_0288_));
 sg13g2_nor2_1 _1210_ (.A(_0108_),
    .B(net154),
    .Y(_0300_));
 sg13g2_a22oi_1 _1211_ (.Y(_0301_),
    .B1(_0248_),
    .B2(_0300_),
    .A2(_0123_),
    .A1(_0108_));
 sg13g2_a22oi_1 _1212_ (.Y(_0302_),
    .B1(_0299_),
    .B2(_0301_),
    .A2(_0291_),
    .A1(_0280_));
 sg13g2_a21oi_1 _1213_ (.A1(_0100_),
    .A2(_0301_),
    .Y(_0303_),
    .B1(_0302_));
 sg13g2_a21o_1 _1214_ (.A2(_0302_),
    .A1(_0100_),
    .B1(_0303_),
    .X(\inst_sine_A.sample[5] ));
 sg13g2_xnor2_1 _1215_ (.Y(\inst_sine_A.sample[6] ),
    .A(_0100_),
    .B(_0292_));
 sg13g2_xnor2_1 _1216_ (.Y(_0023_),
    .A(\product[7] ),
    .B(net238));
 sg13g2_nor3_2 _1217_ (.A(\product[7] ),
    .B(net238),
    .C(net242),
    .Y(_0304_));
 sg13g2_o21ai_1 _1218_ (.B1(net242),
    .Y(_0305_),
    .A1(\product[7] ),
    .A2(net238));
 sg13g2_nand2b_1 _1219_ (.Y(_0024_),
    .B(net243),
    .A_N(_0304_));
 sg13g2_nor2b_1 _1220_ (.A(\product[10] ),
    .B_N(_0304_),
    .Y(_0306_));
 sg13g2_xor2_1 _1221_ (.B(_0304_),
    .A(net236),
    .X(_0025_));
 sg13g2_nor2b_1 _1222_ (.A(net230),
    .B_N(_0306_),
    .Y(_0307_));
 sg13g2_xor2_1 _1223_ (.B(_0306_),
    .A(net230),
    .X(_0026_));
 sg13g2_nor2b_1 _1224_ (.A(\product[12] ),
    .B_N(_0307_),
    .Y(_0308_));
 sg13g2_xor2_1 _1225_ (.B(_0307_),
    .A(net234),
    .X(_0027_));
 sg13g2_nor2b_1 _1226_ (.A(\product[13] ),
    .B_N(_0308_),
    .Y(_0309_));
 sg13g2_xor2_1 _1227_ (.B(_0308_),
    .A(net232),
    .X(_0028_));
 sg13g2_xnor2_1 _1228_ (.Y(_0029_),
    .A(net228),
    .B(_0309_));
 sg13g2_nand2_1 _1229_ (.Y(_0310_),
    .A(net174),
    .B(net170));
 sg13g2_nand2_1 _1230_ (.Y(_0311_),
    .A(net176),
    .B(net168));
 sg13g2_nand2_1 _1231_ (.Y(_0312_),
    .A(\sine_Breg[5] ),
    .B(\sine_Areg[0] ));
 sg13g2_xor2_1 _1232_ (.B(_0311_),
    .A(_0310_),
    .X(_0313_));
 sg13g2_nand2b_1 _1233_ (.Y(_0314_),
    .B(_0313_),
    .A_N(_0312_));
 sg13g2_o21ai_1 _1234_ (.B1(_0314_),
    .Y(_0315_),
    .A1(_0310_),
    .A2(_0311_));
 sg13g2_nand2_1 _1235_ (.Y(_0316_),
    .A(net192),
    .B(\sine_Areg[0] ));
 sg13g2_nor2b_1 _1236_ (.A(_0316_),
    .B_N(_0315_),
    .Y(_0317_));
 sg13g2_nand2b_1 _1237_ (.Y(_0318_),
    .B(_0315_),
    .A_N(_0316_));
 sg13g2_and4_1 _1238_ (.A(net185),
    .B(net181),
    .C(net165),
    .D(net167),
    .X(_0319_));
 sg13g2_nand4_1 _1239_ (.B(net181),
    .C(net165),
    .A(net185),
    .Y(_0320_),
    .D(net167));
 sg13g2_nand2_1 _1240_ (.Y(_0321_),
    .A(net179),
    .B(net169));
 sg13g2_a22oi_1 _1241_ (.Y(_0322_),
    .B1(net167),
    .B2(net181),
    .A2(net165),
    .A1(net185));
 sg13g2_or3_1 _1242_ (.A(_0319_),
    .B(_0321_),
    .C(_0322_),
    .X(_0323_));
 sg13g2_o21ai_1 _1243_ (.B1(_0320_),
    .Y(_0324_),
    .A1(_0321_),
    .A2(_0322_));
 sg13g2_nand2_1 _1244_ (.Y(_0325_),
    .A(net179),
    .B(net167));
 sg13g2_and4_1 _1245_ (.A(net185),
    .B(net181),
    .C(net163),
    .D(net165),
    .X(_0326_));
 sg13g2_nand4_1 _1246_ (.B(net181),
    .C(net163),
    .A(net185),
    .Y(_0327_),
    .D(net165));
 sg13g2_a22oi_1 _1247_ (.Y(_0328_),
    .B1(net165),
    .B2(net181),
    .A2(net163),
    .A1(net185));
 sg13g2_or3_1 _1248_ (.A(_0325_),
    .B(_0326_),
    .C(_0328_),
    .X(_0329_));
 sg13g2_o21ai_1 _1249_ (.B1(_0325_),
    .Y(_0330_),
    .A1(_0326_),
    .A2(_0328_));
 sg13g2_and3_1 _1250_ (.X(_0331_),
    .A(_0324_),
    .B(_0329_),
    .C(_0330_));
 sg13g2_nand3_1 _1251_ (.B(_0329_),
    .C(_0330_),
    .A(_0324_),
    .Y(_0332_));
 sg13g2_a21o_1 _1252_ (.A2(_0330_),
    .A1(_0329_),
    .B1(_0324_),
    .X(_0333_));
 sg13g2_xnor2_1 _1253_ (.Y(_0334_),
    .A(_0312_),
    .B(_0313_));
 sg13g2_and3_1 _1254_ (.X(_0335_),
    .A(_0332_),
    .B(_0333_),
    .C(_0334_));
 sg13g2_a21o_1 _1255_ (.A2(_0334_),
    .A1(_0333_),
    .B1(_0331_),
    .X(_0336_));
 sg13g2_o21ai_1 _1256_ (.B1(_0327_),
    .Y(_0337_),
    .A1(_0325_),
    .A2(_0328_));
 sg13g2_nand2_1 _1257_ (.Y(_0338_),
    .A(net178),
    .B(net165));
 sg13g2_nand2_1 _1258_ (.Y(_0339_),
    .A(net180),
    .B(net160));
 sg13g2_and4_1 _1259_ (.A(net184),
    .B(net180),
    .C(net160),
    .D(net163),
    .X(_0340_));
 sg13g2_nand4_1 _1260_ (.B(net180),
    .C(net160),
    .A(net184),
    .Y(_0341_),
    .D(net163));
 sg13g2_a22oi_1 _1261_ (.Y(_0342_),
    .B1(net163),
    .B2(net181),
    .A2(net160),
    .A1(net183));
 sg13g2_or3_1 _1262_ (.A(_0338_),
    .B(_0340_),
    .C(_0342_),
    .X(_0343_));
 sg13g2_o21ai_1 _1263_ (.B1(_0338_),
    .Y(_0344_),
    .A1(_0340_),
    .A2(_0342_));
 sg13g2_and3_1 _1264_ (.X(_0345_),
    .A(_0337_),
    .B(_0343_),
    .C(_0344_));
 sg13g2_nand3_1 _1265_ (.B(_0343_),
    .C(_0344_),
    .A(_0337_),
    .Y(_0346_));
 sg13g2_a21oi_1 _1266_ (.A1(_0343_),
    .A2(_0344_),
    .Y(_0347_),
    .B1(_0337_));
 sg13g2_nand2_1 _1267_ (.Y(_0348_),
    .A(\sine_Breg[5] ),
    .B(net170));
 sg13g2_nand2_1 _1268_ (.Y(_0349_),
    .A(net173),
    .B(net166));
 sg13g2_and4_1 _1269_ (.A(net176),
    .B(net174),
    .C(net166),
    .D(net168),
    .X(_0350_));
 sg13g2_a22oi_1 _1270_ (.Y(_0351_),
    .B1(net168),
    .B2(net174),
    .A2(net166),
    .A1(net176));
 sg13g2_nor3_1 _1271_ (.A(_0348_),
    .B(_0350_),
    .C(_0351_),
    .Y(_0352_));
 sg13g2_o21ai_1 _1272_ (.B1(_0348_),
    .Y(_0353_),
    .A1(_0350_),
    .A2(_0351_));
 sg13g2_nand2b_1 _1273_ (.Y(_0354_),
    .B(_0353_),
    .A_N(_0352_));
 sg13g2_or3_1 _1274_ (.A(_0345_),
    .B(_0347_),
    .C(_0354_),
    .X(_0355_));
 sg13g2_o21ai_1 _1275_ (.B1(_0354_),
    .Y(_0356_),
    .A1(_0345_),
    .A2(_0347_));
 sg13g2_nand3_1 _1276_ (.B(_0355_),
    .C(_0356_),
    .A(_0336_),
    .Y(_0357_));
 sg13g2_xor2_1 _1277_ (.B(_0316_),
    .A(_0315_),
    .X(_0358_));
 sg13g2_a21oi_1 _1278_ (.A1(_0355_),
    .A2(_0356_),
    .Y(_0359_),
    .B1(_0336_));
 sg13g2_a21o_1 _1279_ (.A2(_0356_),
    .A1(_0355_),
    .B1(_0336_),
    .X(_0360_));
 sg13g2_o21ai_1 _1280_ (.B1(_0357_),
    .Y(_0361_),
    .A1(_0358_),
    .A2(_0359_));
 sg13g2_or2_1 _1281_ (.X(_0362_),
    .B(_0352_),
    .A(_0350_));
 sg13g2_nor2b_1 _1282_ (.A(\sine_Areg[0] ),
    .B_N(net172),
    .Y(_0363_));
 sg13g2_nand2_1 _1283_ (.Y(_0364_),
    .A(net168),
    .B(net192));
 sg13g2_nor2_1 _1284_ (.A(_0348_),
    .B(_0364_),
    .Y(_0365_));
 sg13g2_a22oi_1 _1285_ (.Y(_0366_),
    .B1(net170),
    .B2(net192),
    .A2(\sine_Breg[5] ),
    .A1(net168));
 sg13g2_nor2_1 _1286_ (.A(_0365_),
    .B(_0366_),
    .Y(_0367_));
 sg13g2_xor2_1 _1287_ (.B(_0367_),
    .A(_0363_),
    .X(_0368_));
 sg13g2_xnor2_1 _1288_ (.Y(_0369_),
    .A(_0362_),
    .B(_0368_));
 sg13g2_o21ai_1 _1289_ (.B1(_0346_),
    .Y(_0370_),
    .A1(_0347_),
    .A2(_0354_));
 sg13g2_and4_1 _1290_ (.A(net162),
    .B(net178),
    .C(net164),
    .D(net175),
    .X(_0371_));
 sg13g2_a22oi_1 _1291_ (.Y(_0372_),
    .B1(net164),
    .B2(net176),
    .A2(net178),
    .A1(net162));
 sg13g2_nor3_1 _1292_ (.A(_0349_),
    .B(_0371_),
    .C(_0372_),
    .Y(_0373_));
 sg13g2_o21ai_1 _1293_ (.B1(_0349_),
    .Y(_0374_),
    .A1(_0371_),
    .A2(_0372_));
 sg13g2_nand2b_1 _1294_ (.Y(_0375_),
    .B(_0374_),
    .A_N(_0373_));
 sg13g2_o21ai_1 _1295_ (.B1(_0341_),
    .Y(_0376_),
    .A1(_0338_),
    .A2(_0342_));
 sg13g2_a21oi_1 _1296_ (.A1(net183),
    .A2(net189),
    .Y(_0377_),
    .B1(net172));
 sg13g2_and3_1 _1297_ (.X(_0378_),
    .A(net183),
    .B(\sine_Areg[7] ),
    .C(net171));
 sg13g2_nand3_1 _1298_ (.B(net189),
    .C(net171),
    .A(net183),
    .Y(_0379_));
 sg13g2_or3_1 _1299_ (.A(_0339_),
    .B(_0377_),
    .C(_0378_),
    .X(_0380_));
 sg13g2_o21ai_1 _1300_ (.B1(_0339_),
    .Y(_0381_),
    .A1(_0377_),
    .A2(_0378_));
 sg13g2_and3_1 _1301_ (.X(_0382_),
    .A(_0376_),
    .B(_0380_),
    .C(_0381_));
 sg13g2_nand3_1 _1302_ (.B(_0380_),
    .C(_0381_),
    .A(_0376_),
    .Y(_0383_));
 sg13g2_a21oi_1 _1303_ (.A1(_0380_),
    .A2(_0381_),
    .Y(_0384_),
    .B1(_0376_));
 sg13g2_or3_1 _1304_ (.A(_0375_),
    .B(_0382_),
    .C(_0384_),
    .X(_0385_));
 sg13g2_o21ai_1 _1305_ (.B1(_0375_),
    .Y(_0386_),
    .A1(_0382_),
    .A2(_0384_));
 sg13g2_and3_1 _1306_ (.X(_0387_),
    .A(_0370_),
    .B(_0385_),
    .C(_0386_));
 sg13g2_nand3_1 _1307_ (.B(_0385_),
    .C(_0386_),
    .A(_0370_),
    .Y(_0388_));
 sg13g2_a21oi_1 _1308_ (.A1(_0385_),
    .A2(_0386_),
    .Y(_0389_),
    .B1(_0370_));
 sg13g2_or3_1 _1309_ (.A(_0369_),
    .B(_0387_),
    .C(_0389_),
    .X(_0390_));
 sg13g2_o21ai_1 _1310_ (.B1(_0369_),
    .Y(_0391_),
    .A1(_0387_),
    .A2(_0389_));
 sg13g2_and3_1 _1311_ (.X(_0392_),
    .A(_0361_),
    .B(_0390_),
    .C(_0391_));
 sg13g2_nand3_1 _1312_ (.B(_0390_),
    .C(_0391_),
    .A(_0361_),
    .Y(_0393_));
 sg13g2_a21o_1 _1313_ (.A2(_0391_),
    .A1(_0390_),
    .B1(_0361_),
    .X(_0394_));
 sg13g2_nand3_1 _1314_ (.B(_0393_),
    .C(_0394_),
    .A(_0318_),
    .Y(_0395_));
 sg13g2_a21o_1 _1315_ (.A2(_0394_),
    .A1(_0393_),
    .B1(_0318_),
    .X(_0396_));
 sg13g2_nand2_1 _1316_ (.Y(_0397_),
    .A(_0395_),
    .B(_0396_));
 sg13g2_and4_1 _1317_ (.A(net186),
    .B(net182),
    .C(net166),
    .D(net169),
    .X(_0398_));
 sg13g2_nand4_1 _1318_ (.B(net182),
    .C(net167),
    .A(net186),
    .Y(_0399_),
    .D(net169));
 sg13g2_nand2_1 _1319_ (.Y(_0400_),
    .A(net179),
    .B(\sine_Areg[1] ));
 sg13g2_a22oi_1 _1320_ (.Y(_0401_),
    .B1(net169),
    .B2(net182),
    .A2(net167),
    .A1(net186));
 sg13g2_nor3_1 _1321_ (.A(_0398_),
    .B(_0400_),
    .C(_0401_),
    .Y(_0402_));
 sg13g2_o21ai_1 _1322_ (.B1(_0399_),
    .Y(_0403_),
    .A1(_0400_),
    .A2(_0401_));
 sg13g2_o21ai_1 _1323_ (.B1(_0321_),
    .Y(_0404_),
    .A1(_0319_),
    .A2(_0322_));
 sg13g2_and3_1 _1324_ (.X(_0405_),
    .A(_0323_),
    .B(_0403_),
    .C(_0404_));
 sg13g2_and4_1 _1325_ (.A(net177),
    .B(net174),
    .C(\sine_Areg[1] ),
    .D(\sine_Areg[0] ),
    .X(_0406_));
 sg13g2_a22oi_1 _1326_ (.Y(_0407_),
    .B1(\sine_Areg[0] ),
    .B2(net174),
    .A2(net170),
    .A1(net177));
 sg13g2_nor2_1 _1327_ (.A(_0406_),
    .B(_0407_),
    .Y(_0408_));
 sg13g2_a21o_1 _1328_ (.A2(_0404_),
    .A1(_0323_),
    .B1(_0403_),
    .X(_0409_));
 sg13g2_nor2b_1 _1329_ (.A(_0405_),
    .B_N(_0409_),
    .Y(_0410_));
 sg13g2_a21oi_1 _1330_ (.A1(_0408_),
    .A2(_0409_),
    .Y(_0411_),
    .B1(_0405_));
 sg13g2_a21oi_1 _1331_ (.A1(_0332_),
    .A2(_0333_),
    .Y(_0412_),
    .B1(_0334_));
 sg13g2_nor3_1 _1332_ (.A(_0335_),
    .B(_0411_),
    .C(_0412_),
    .Y(_0413_));
 sg13g2_o21ai_1 _1333_ (.B1(_0411_),
    .Y(_0414_),
    .A1(_0335_),
    .A2(_0412_));
 sg13g2_nand2b_1 _1334_ (.Y(_0415_),
    .B(_0414_),
    .A_N(_0413_));
 sg13g2_a21oi_1 _1335_ (.A1(_0406_),
    .A2(_0414_),
    .Y(_0416_),
    .B1(_0413_));
 sg13g2_a21o_1 _1336_ (.A2(_0360_),
    .A1(_0357_),
    .B1(_0358_),
    .X(_0417_));
 sg13g2_nand3_1 _1337_ (.B(_0358_),
    .C(_0360_),
    .A(_0357_),
    .Y(_0418_));
 sg13g2_a21o_1 _1338_ (.A2(_0418_),
    .A1(_0417_),
    .B1(_0416_),
    .X(_0419_));
 sg13g2_nand3_1 _1339_ (.B(_0417_),
    .C(_0418_),
    .A(_0416_),
    .Y(_0420_));
 sg13g2_xnor2_1 _1340_ (.Y(_0421_),
    .A(_0408_),
    .B(_0410_));
 sg13g2_nand4_1 _1341_ (.B(net182),
    .C(net169),
    .A(net186),
    .Y(_0422_),
    .D(net170));
 sg13g2_a22oi_1 _1342_ (.Y(_0423_),
    .B1(net170),
    .B2(net182),
    .A2(net168),
    .A1(net186));
 sg13g2_nand2_1 _1343_ (.Y(_0424_),
    .A(net179),
    .B(\sine_Areg[0] ));
 sg13g2_nor2_1 _1344_ (.A(_0423_),
    .B(_0424_),
    .Y(_0425_));
 sg13g2_nand4_1 _1345_ (.B(net182),
    .C(net170),
    .A(net186),
    .Y(_0426_),
    .D(\sine_Areg[0] ));
 sg13g2_a221oi_1 _1346_ (.B2(_0425_),
    .C1(_0426_),
    .B1(_0422_),
    .A1(_0103_),
    .Y(_0427_),
    .A2(net168));
 sg13g2_a21oi_1 _1347_ (.A1(net177),
    .A2(\sine_Areg[0] ),
    .Y(_0428_),
    .B1(_0427_));
 sg13g2_o21ai_1 _1348_ (.B1(_0422_),
    .Y(_0429_),
    .A1(_0423_),
    .A2(_0424_));
 sg13g2_o21ai_1 _1349_ (.B1(_0400_),
    .Y(_0430_),
    .A1(_0398_),
    .A2(_0401_));
 sg13g2_nor2b_1 _1350_ (.A(_0402_),
    .B_N(_0430_),
    .Y(_0431_));
 sg13g2_nand2_1 _1351_ (.Y(_0432_),
    .A(_0429_),
    .B(_0431_));
 sg13g2_o21ai_1 _1352_ (.B1(_0432_),
    .Y(_0433_),
    .A1(_0421_),
    .A2(_0428_));
 sg13g2_nand2_1 _1353_ (.Y(_0434_),
    .A(net177),
    .B(_0427_));
 sg13g2_nor2_1 _1354_ (.A(_0429_),
    .B(_0431_),
    .Y(_0435_));
 sg13g2_o21ai_1 _1355_ (.B1(_0434_),
    .Y(_0436_),
    .A1(_0421_),
    .A2(_0435_));
 sg13g2_xnor2_1 _1356_ (.Y(_0437_),
    .A(_0406_),
    .B(_0415_));
 sg13g2_nand4_1 _1357_ (.B(_0433_),
    .C(_0436_),
    .A(_0420_),
    .Y(_0438_),
    .D(_0437_));
 sg13g2_nand2_1 _1358_ (.Y(_0439_),
    .A(_0419_),
    .B(_0438_));
 sg13g2_a22oi_1 _1359_ (.Y(_0440_),
    .B1(_0419_),
    .B2(_0438_),
    .A2(_0396_),
    .A1(_0395_));
 sg13g2_xor2_1 _1360_ (.B(_0439_),
    .A(_0397_),
    .X(_0035_));
 sg13g2_o21ai_1 _1361_ (.B1(_0388_),
    .Y(_0441_),
    .A1(_0369_),
    .A2(_0389_));
 sg13g2_a21oi_1 _1362_ (.A1(_0363_),
    .A2(_0367_),
    .Y(_0442_),
    .B1(_0365_));
 sg13g2_or2_1 _1363_ (.X(_0443_),
    .B(_0373_),
    .A(_0371_));
 sg13g2_nor2b_1 _1364_ (.A(net170),
    .B_N(net172),
    .Y(_0444_));
 sg13g2_nor2b_1 _1365_ (.A(_0364_),
    .B_N(_0444_),
    .Y(_0445_));
 sg13g2_xnor2_1 _1366_ (.Y(_0446_),
    .A(_0364_),
    .B(_0444_));
 sg13g2_nand2_1 _1367_ (.Y(_0447_),
    .A(_0443_),
    .B(_0446_));
 sg13g2_xnor2_1 _1368_ (.Y(_0448_),
    .A(_0443_),
    .B(_0446_));
 sg13g2_xor2_1 _1369_ (.B(_0448_),
    .A(_0442_),
    .X(_0449_));
 sg13g2_o21ai_1 _1370_ (.B1(_0383_),
    .Y(_0450_),
    .A1(_0375_),
    .A2(_0384_));
 sg13g2_nand2_1 _1371_ (.Y(_0451_),
    .A(net166),
    .B(\sine_Breg[5] ));
 sg13g2_and4_1 _1372_ (.A(net161),
    .B(net164),
    .C(net175),
    .D(net173),
    .X(_0452_));
 sg13g2_a22oi_1 _1373_ (.Y(_0453_),
    .B1(net173),
    .B2(net164),
    .A2(net175),
    .A1(net161));
 sg13g2_nor3_1 _1374_ (.A(_0451_),
    .B(_0452_),
    .C(_0453_),
    .Y(_0454_));
 sg13g2_o21ai_1 _1375_ (.B1(_0451_),
    .Y(_0455_),
    .A1(_0452_),
    .A2(_0453_));
 sg13g2_nor2b_1 _1376_ (.A(_0454_),
    .B_N(_0455_),
    .Y(_0456_));
 sg13g2_o21ai_1 _1377_ (.B1(_0379_),
    .Y(_0457_),
    .A1(_0339_),
    .A2(_0377_));
 sg13g2_and3_1 _1378_ (.X(_0458_),
    .A(net184),
    .B(net189),
    .C(net180));
 sg13g2_nand3_1 _1379_ (.B(net189),
    .C(net180),
    .A(net183),
    .Y(_0459_));
 sg13g2_o21ai_1 _1380_ (.B1(net189),
    .Y(_0460_),
    .A1(net183),
    .A2(net180));
 sg13g2_nand2_1 _1381_ (.Y(_0461_),
    .A(net160),
    .B(net178));
 sg13g2_or3_1 _1382_ (.A(_0458_),
    .B(_0460_),
    .C(_0461_),
    .X(_0462_));
 sg13g2_o21ai_1 _1383_ (.B1(_0461_),
    .Y(_0463_),
    .A1(_0458_),
    .A2(_0460_));
 sg13g2_nand3_1 _1384_ (.B(_0462_),
    .C(_0463_),
    .A(_0457_),
    .Y(_0464_));
 sg13g2_a21o_1 _1385_ (.A2(_0463_),
    .A1(_0462_),
    .B1(_0457_),
    .X(_0465_));
 sg13g2_nand3_1 _1386_ (.B(_0464_),
    .C(_0465_),
    .A(_0456_),
    .Y(_0466_));
 sg13g2_a21o_1 _1387_ (.A2(_0465_),
    .A1(_0464_),
    .B1(_0456_),
    .X(_0467_));
 sg13g2_nand3_1 _1388_ (.B(_0466_),
    .C(_0467_),
    .A(_0450_),
    .Y(_0468_));
 sg13g2_a21o_1 _1389_ (.A2(_0467_),
    .A1(_0466_),
    .B1(_0450_),
    .X(_0469_));
 sg13g2_nand3_1 _1390_ (.B(_0468_),
    .C(_0469_),
    .A(_0449_),
    .Y(_0470_));
 sg13g2_a21o_1 _1391_ (.A2(_0469_),
    .A1(_0468_),
    .B1(_0449_),
    .X(_0471_));
 sg13g2_and2_1 _1392_ (.A(_0470_),
    .B(_0471_),
    .X(_0472_));
 sg13g2_nand3_1 _1393_ (.B(_0470_),
    .C(_0471_),
    .A(_0441_),
    .Y(_0473_));
 sg13g2_a21o_1 _1394_ (.A2(_0471_),
    .A1(_0470_),
    .B1(_0441_),
    .X(_0474_));
 sg13g2_and4_1 _1395_ (.A(_0362_),
    .B(_0368_),
    .C(_0473_),
    .D(_0474_),
    .X(_0475_));
 sg13g2_a22oi_1 _1396_ (.Y(_0476_),
    .B1(_0473_),
    .B2(_0474_),
    .A2(_0368_),
    .A1(_0362_));
 sg13g2_a21oi_1 _1397_ (.A1(_0317_),
    .A2(_0394_),
    .Y(_0477_),
    .B1(_0392_));
 sg13g2_nor3_1 _1398_ (.A(_0475_),
    .B(_0476_),
    .C(_0477_),
    .Y(_0478_));
 sg13g2_o21ai_1 _1399_ (.B1(_0477_),
    .Y(_0479_),
    .A1(_0475_),
    .A2(_0476_));
 sg13g2_nand2b_1 _1400_ (.Y(_0480_),
    .B(_0479_),
    .A_N(_0478_));
 sg13g2_xnor2_1 _1401_ (.Y(_0036_),
    .A(_0440_),
    .B(_0480_));
 sg13g2_a21o_1 _1402_ (.A2(_0472_),
    .A1(_0441_),
    .B1(_0475_),
    .X(_0481_));
 sg13g2_o21ai_1 _1403_ (.B1(_0447_),
    .Y(_0482_),
    .A1(_0442_),
    .A2(_0448_));
 sg13g2_inv_1 _1404_ (.Y(_0483_),
    .A(_0482_));
 sg13g2_nand2_1 _1405_ (.Y(_0484_),
    .A(_0468_),
    .B(_0470_));
 sg13g2_or2_1 _1406_ (.X(_0485_),
    .B(_0454_),
    .A(_0452_));
 sg13g2_nor2b_1 _1407_ (.A(net168),
    .B_N(net172),
    .Y(_0486_));
 sg13g2_nand2_1 _1408_ (.Y(_0487_),
    .A(net166),
    .B(net192));
 sg13g2_and3_1 _1409_ (.X(_0488_),
    .A(net166),
    .B(net191),
    .C(_0486_));
 sg13g2_xnor2_1 _1410_ (.Y(_0489_),
    .A(_0486_),
    .B(_0487_));
 sg13g2_and2_1 _1411_ (.A(_0485_),
    .B(_0489_),
    .X(_0490_));
 sg13g2_xor2_1 _1412_ (.B(_0489_),
    .A(_0485_),
    .X(_0491_));
 sg13g2_xnor2_1 _1413_ (.Y(_0492_),
    .A(_0445_),
    .B(_0491_));
 sg13g2_nand2_1 _1414_ (.Y(_0493_),
    .A(_0464_),
    .B(_0466_));
 sg13g2_nand2_1 _1415_ (.Y(_0494_),
    .A(net164),
    .B(\sine_Breg[5] ));
 sg13g2_and4_1 _1416_ (.A(net159),
    .B(net161),
    .C(net175),
    .D(net173),
    .X(_0495_));
 sg13g2_a22oi_1 _1417_ (.Y(_0496_),
    .B1(net173),
    .B2(net161),
    .A2(net175),
    .A1(net159));
 sg13g2_nor3_1 _1418_ (.A(_0494_),
    .B(_0495_),
    .C(_0496_),
    .Y(_0497_));
 sg13g2_o21ai_1 _1419_ (.B1(_0494_),
    .Y(_0498_),
    .A1(_0495_),
    .A2(_0496_));
 sg13g2_nand2b_1 _1420_ (.Y(_0499_),
    .B(_0498_),
    .A_N(_0497_));
 sg13g2_and2_1 _1421_ (.A(net189),
    .B(net178),
    .X(_0500_));
 sg13g2_nand2_1 _1422_ (.Y(_0501_),
    .A(net189),
    .B(net178));
 sg13g2_or3_1 _1423_ (.A(_0458_),
    .B(_0460_),
    .C(_0500_),
    .X(_0502_));
 sg13g2_o21ai_1 _1424_ (.B1(_0500_),
    .Y(_0503_),
    .A1(_0458_),
    .A2(_0460_));
 sg13g2_and4_2 _1425_ (.A(net183),
    .B(net190),
    .C(net180),
    .D(net178),
    .X(_0504_));
 sg13g2_nand4_1 _1426_ (.B(net190),
    .C(net180),
    .A(net183),
    .Y(_0505_),
    .D(net178));
 sg13g2_and4_1 _1427_ (.A(_0459_),
    .B(_0462_),
    .C(_0502_),
    .D(_0503_),
    .X(_0506_));
 sg13g2_nor2_1 _1428_ (.A(_0504_),
    .B(_0506_),
    .Y(_0507_));
 sg13g2_xnor2_1 _1429_ (.Y(_0508_),
    .A(_0499_),
    .B(_0507_));
 sg13g2_nand2_1 _1430_ (.Y(_0509_),
    .A(_0493_),
    .B(_0508_));
 sg13g2_xnor2_1 _1431_ (.Y(_0510_),
    .A(_0493_),
    .B(_0508_));
 sg13g2_xor2_1 _1432_ (.B(_0510_),
    .A(_0492_),
    .X(_0511_));
 sg13g2_nand2_1 _1433_ (.Y(_0512_),
    .A(_0484_),
    .B(_0511_));
 sg13g2_xnor2_1 _1434_ (.Y(_0513_),
    .A(_0484_),
    .B(_0511_));
 sg13g2_xnor2_1 _1435_ (.Y(_0514_),
    .A(_0482_),
    .B(_0513_));
 sg13g2_nor2_1 _1436_ (.A(_0481_),
    .B(_0514_),
    .Y(_0515_));
 sg13g2_xnor2_1 _1437_ (.Y(_0516_),
    .A(_0481_),
    .B(_0514_));
 sg13g2_a21oi_1 _1438_ (.A1(_0440_),
    .A2(_0479_),
    .Y(_0517_),
    .B1(_0478_));
 sg13g2_xor2_1 _1439_ (.B(_0517_),
    .A(_0516_),
    .X(_0037_));
 sg13g2_a21oi_1 _1440_ (.A1(_0445_),
    .A2(_0491_),
    .Y(_0518_),
    .B1(_0490_));
 sg13g2_o21ai_1 _1441_ (.B1(_0509_),
    .Y(_0519_),
    .A1(_0492_),
    .A2(_0510_));
 sg13g2_or2_1 _1442_ (.X(_0520_),
    .B(_0497_),
    .A(_0495_));
 sg13g2_nor2b_1 _1443_ (.A(net166),
    .B_N(net171),
    .Y(_0521_));
 sg13g2_nand2_1 _1444_ (.Y(_0522_),
    .A(net164),
    .B(net191));
 sg13g2_and3_1 _1445_ (.X(_0523_),
    .A(net164),
    .B(net191),
    .C(_0521_));
 sg13g2_xnor2_1 _1446_ (.Y(_0524_),
    .A(_0521_),
    .B(_0522_));
 sg13g2_and2_1 _1447_ (.A(_0520_),
    .B(_0524_),
    .X(_0525_));
 sg13g2_xor2_1 _1448_ (.B(_0524_),
    .A(_0520_),
    .X(_0526_));
 sg13g2_xnor2_1 _1449_ (.Y(_0527_),
    .A(_0488_),
    .B(_0526_));
 sg13g2_o21ai_1 _1450_ (.B1(_0505_),
    .Y(_0528_),
    .A1(_0499_),
    .A2(_0506_));
 sg13g2_and2_1 _1451_ (.A(net161),
    .B(\sine_Breg[5] ),
    .X(_0529_));
 sg13g2_and3_2 _1452_ (.X(_0530_),
    .A(net190),
    .B(net175),
    .C(net173));
 sg13g2_a22oi_1 _1453_ (.Y(_0531_),
    .B1(net173),
    .B2(net159),
    .A2(net175),
    .A1(net190));
 sg13g2_a21oi_1 _1454_ (.A1(net159),
    .A2(_0530_),
    .Y(_0532_),
    .B1(_0531_));
 sg13g2_xor2_1 _1455_ (.B(_0532_),
    .A(_0529_),
    .X(_0533_));
 sg13g2_a21oi_2 _1456_ (.B1(_0504_),
    .Y(_0534_),
    .A2(_0501_),
    .A1(_0460_));
 sg13g2_xnor2_1 _1457_ (.Y(_0535_),
    .A(_0533_),
    .B(_0534_));
 sg13g2_nand2b_1 _1458_ (.Y(_0536_),
    .B(_0528_),
    .A_N(_0535_));
 sg13g2_xor2_1 _1459_ (.B(_0535_),
    .A(_0528_),
    .X(_0537_));
 sg13g2_xor2_1 _1460_ (.B(_0537_),
    .A(_0527_),
    .X(_0538_));
 sg13g2_and2_1 _1461_ (.A(_0519_),
    .B(_0538_),
    .X(_0539_));
 sg13g2_xnor2_1 _1462_ (.Y(_0540_),
    .A(_0519_),
    .B(_0538_));
 sg13g2_nor2_1 _1463_ (.A(_0518_),
    .B(_0540_),
    .Y(_0541_));
 sg13g2_xor2_1 _1464_ (.B(_0540_),
    .A(_0518_),
    .X(_0542_));
 sg13g2_o21ai_1 _1465_ (.B1(_0512_),
    .Y(_0543_),
    .A1(_0483_),
    .A2(_0513_));
 sg13g2_nand2_1 _1466_ (.Y(_0544_),
    .A(_0542_),
    .B(_0543_));
 sg13g2_xnor2_1 _1467_ (.Y(_0545_),
    .A(_0542_),
    .B(_0543_));
 sg13g2_a221oi_1 _1468_ (.B2(_0514_),
    .C1(_0478_),
    .B1(_0481_),
    .A1(_0440_),
    .Y(_0546_),
    .A2(_0479_));
 sg13g2_or2_1 _1469_ (.X(_0547_),
    .B(_0546_),
    .A(_0515_));
 sg13g2_nor3_1 _1470_ (.A(_0515_),
    .B(_0545_),
    .C(_0546_),
    .Y(_0548_));
 sg13g2_xor2_1 _1471_ (.B(_0547_),
    .A(_0545_),
    .X(_0030_));
 sg13g2_a21oi_1 _1472_ (.A1(_0488_),
    .A2(_0526_),
    .Y(_0549_),
    .B1(_0525_));
 sg13g2_o21ai_1 _1473_ (.B1(_0536_),
    .Y(_0550_),
    .A1(_0527_),
    .A2(_0537_));
 sg13g2_a22oi_1 _1474_ (.Y(_0551_),
    .B1(_0532_),
    .B2(_0529_),
    .A2(_0530_),
    .A1(net159));
 sg13g2_a22oi_1 _1475_ (.Y(_0552_),
    .B1(net191),
    .B2(net161),
    .A2(_0104_),
    .A1(net171));
 sg13g2_and4_1 _1476_ (.A(net171),
    .B(net161),
    .C(_0104_),
    .D(net191),
    .X(_0553_));
 sg13g2_nor2_1 _1477_ (.A(_0552_),
    .B(_0553_),
    .Y(_0554_));
 sg13g2_nor2b_1 _1478_ (.A(_0551_),
    .B_N(_0554_),
    .Y(_0555_));
 sg13g2_xnor2_1 _1479_ (.Y(_0556_),
    .A(_0551_),
    .B(_0554_));
 sg13g2_xnor2_1 _1480_ (.Y(_0557_),
    .A(_0523_),
    .B(_0556_));
 sg13g2_a21o_1 _1481_ (.A2(_0534_),
    .A1(_0533_),
    .B1(_0504_),
    .X(_0558_));
 sg13g2_o21ai_1 _1482_ (.B1(net190),
    .Y(_0559_),
    .A1(net175),
    .A2(net173));
 sg13g2_or2_2 _1483_ (.X(_0560_),
    .B(_0559_),
    .A(_0530_));
 sg13g2_nand2_1 _1484_ (.Y(_0561_),
    .A(net159),
    .B(\sine_Breg[5] ));
 sg13g2_nor2_1 _1485_ (.A(_0560_),
    .B(_0561_),
    .Y(_0562_));
 sg13g2_xor2_1 _1486_ (.B(_0561_),
    .A(_0560_),
    .X(_0563_));
 sg13g2_nand2_1 _1487_ (.Y(_0564_),
    .A(_0534_),
    .B(_0563_));
 sg13g2_xnor2_1 _1488_ (.Y(_0565_),
    .A(_0534_),
    .B(_0563_));
 sg13g2_nand2b_1 _1489_ (.Y(_0566_),
    .B(_0558_),
    .A_N(_0565_));
 sg13g2_xor2_1 _1490_ (.B(_0565_),
    .A(_0558_),
    .X(_0567_));
 sg13g2_xor2_1 _1491_ (.B(_0567_),
    .A(_0557_),
    .X(_0568_));
 sg13g2_nand2_1 _1492_ (.Y(_0569_),
    .A(_0550_),
    .B(_0568_));
 sg13g2_xnor2_1 _1493_ (.Y(_0570_),
    .A(_0550_),
    .B(_0568_));
 sg13g2_xor2_1 _1494_ (.B(_0570_),
    .A(_0549_),
    .X(_0571_));
 sg13g2_or3_1 _1495_ (.A(_0539_),
    .B(_0541_),
    .C(_0571_),
    .X(_0572_));
 sg13g2_o21ai_1 _1496_ (.B1(_0571_),
    .Y(_0573_),
    .A1(_0539_),
    .A2(_0541_));
 sg13g2_and2_1 _1497_ (.A(_0572_),
    .B(_0573_),
    .X(_0574_));
 sg13g2_o21ai_1 _1498_ (.B1(_0544_),
    .Y(_0575_),
    .A1(_0545_),
    .A2(_0547_));
 sg13g2_xor2_1 _1499_ (.B(_0575_),
    .A(_0574_),
    .X(_0031_));
 sg13g2_a21o_1 _1500_ (.A2(_0556_),
    .A1(_0523_),
    .B1(_0555_),
    .X(_0576_));
 sg13g2_o21ai_1 _1501_ (.B1(_0566_),
    .Y(_0577_),
    .A1(_0557_),
    .A2(_0567_));
 sg13g2_nand2_1 _1502_ (.Y(_0578_),
    .A(net190),
    .B(\sine_Breg[5] ));
 sg13g2_nor2_1 _1503_ (.A(_0560_),
    .B(_0578_),
    .Y(_0579_));
 sg13g2_xor2_1 _1504_ (.B(_0578_),
    .A(_0560_),
    .X(_0580_));
 sg13g2_xnor2_1 _1505_ (.Y(_0581_),
    .A(_0534_),
    .B(_0580_));
 sg13g2_a21oi_1 _1506_ (.A1(_0505_),
    .A2(_0564_),
    .Y(_0582_),
    .B1(_0581_));
 sg13g2_nand3_1 _1507_ (.B(_0564_),
    .C(_0581_),
    .A(_0505_),
    .Y(_0583_));
 sg13g2_nand2b_1 _1508_ (.Y(_0584_),
    .B(_0583_),
    .A_N(_0582_));
 sg13g2_nor2_1 _1509_ (.A(_0530_),
    .B(_0562_),
    .Y(_0585_));
 sg13g2_a22oi_1 _1510_ (.Y(_0586_),
    .B1(net191),
    .B2(net159),
    .A2(_0102_),
    .A1(net171));
 sg13g2_nand3_1 _1511_ (.B(net159),
    .C(net191),
    .A(net171),
    .Y(_0587_));
 sg13g2_nor2_1 _1512_ (.A(net162),
    .B(_0587_),
    .Y(_0588_));
 sg13g2_nor2_1 _1513_ (.A(_0586_),
    .B(_0588_),
    .Y(_0589_));
 sg13g2_nor2b_1 _1514_ (.A(_0585_),
    .B_N(_0589_),
    .Y(_0590_));
 sg13g2_xnor2_1 _1515_ (.Y(_0591_),
    .A(_0585_),
    .B(_0589_));
 sg13g2_xor2_1 _1516_ (.B(_0591_),
    .A(_0553_),
    .X(_0592_));
 sg13g2_xnor2_1 _1517_ (.Y(_0593_),
    .A(_0584_),
    .B(_0592_));
 sg13g2_and2_1 _1518_ (.A(_0577_),
    .B(_0593_),
    .X(_0594_));
 sg13g2_xor2_1 _1519_ (.B(_0593_),
    .A(_0577_),
    .X(_0595_));
 sg13g2_and2_1 _1520_ (.A(_0576_),
    .B(_0595_),
    .X(_0596_));
 sg13g2_xor2_1 _1521_ (.B(_0595_),
    .A(_0576_),
    .X(_0597_));
 sg13g2_o21ai_1 _1522_ (.B1(_0569_),
    .Y(_0598_),
    .A1(_0549_),
    .A2(_0570_));
 sg13g2_nand2_1 _1523_ (.Y(_0599_),
    .A(_0597_),
    .B(_0598_));
 sg13g2_xnor2_1 _1524_ (.Y(_0600_),
    .A(_0597_),
    .B(_0598_));
 sg13g2_nand2_1 _1525_ (.Y(_0601_),
    .A(_0544_),
    .B(_0573_));
 sg13g2_a22oi_1 _1526_ (.Y(_0602_),
    .B1(_0601_),
    .B2(_0572_),
    .A2(_0574_),
    .A1(_0548_));
 sg13g2_xor2_1 _1527_ (.B(_0602_),
    .A(_0600_),
    .X(_0032_));
 sg13g2_a21oi_2 _1528_ (.B1(_0590_),
    .Y(_0603_),
    .A2(_0591_),
    .A1(_0553_));
 sg13g2_a21oi_1 _1529_ (.A1(_0583_),
    .A2(_0592_),
    .Y(_0604_),
    .B1(_0582_));
 sg13g2_or3_1 _1530_ (.A(_0504_),
    .B(_0534_),
    .C(_0580_),
    .X(_0605_));
 sg13g2_nand2_1 _1531_ (.Y(_0606_),
    .A(_0504_),
    .B(_0580_));
 sg13g2_nand2_1 _1532_ (.Y(_0607_),
    .A(_0605_),
    .B(_0606_));
 sg13g2_nor2_2 _1533_ (.A(_0530_),
    .B(_0579_),
    .Y(_0608_));
 sg13g2_nand2_1 _1534_ (.Y(_0609_),
    .A(net190),
    .B(net191));
 sg13g2_nor2b_1 _1535_ (.A(net160),
    .B_N(net172),
    .Y(_0610_));
 sg13g2_nor2_1 _1536_ (.A(_0609_),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_xnor2_1 _1537_ (.Y(_0612_),
    .A(_0609_),
    .B(_0610_));
 sg13g2_nor2b_1 _1538_ (.A(_0608_),
    .B_N(_0612_),
    .Y(_0613_));
 sg13g2_xor2_1 _1539_ (.B(_0612_),
    .A(_0608_),
    .X(_0614_));
 sg13g2_nor3_1 _1540_ (.A(net162),
    .B(_0587_),
    .C(_0614_),
    .Y(_0615_));
 sg13g2_xor2_1 _1541_ (.B(_0614_),
    .A(_0588_),
    .X(_0616_));
 sg13g2_xor2_1 _1542_ (.B(_0616_),
    .A(_0607_),
    .X(_0617_));
 sg13g2_nand2b_1 _1543_ (.Y(_0618_),
    .B(_0617_),
    .A_N(_0604_));
 sg13g2_xor2_1 _1544_ (.B(_0617_),
    .A(_0604_),
    .X(_0619_));
 sg13g2_xor2_1 _1545_ (.B(_0619_),
    .A(_0603_),
    .X(_0620_));
 sg13g2_nor3_1 _1546_ (.A(_0594_),
    .B(_0596_),
    .C(_0620_),
    .Y(_0621_));
 sg13g2_o21ai_1 _1547_ (.B1(_0620_),
    .Y(_0622_),
    .A1(_0594_),
    .A2(_0596_));
 sg13g2_nand2b_1 _1548_ (.Y(_0623_),
    .B(_0622_),
    .A_N(_0621_));
 sg13g2_o21ai_1 _1549_ (.B1(_0599_),
    .Y(_0624_),
    .A1(_0600_),
    .A2(_0602_));
 sg13g2_xnor2_1 _1550_ (.Y(_0033_),
    .A(_0623_),
    .B(_0624_));
 sg13g2_or2_1 _1551_ (.X(_0625_),
    .B(_0623_),
    .A(_0600_));
 sg13g2_a21o_1 _1552_ (.A2(_0622_),
    .A1(_0599_),
    .B1(_0621_),
    .X(_0626_));
 sg13g2_o21ai_1 _1553_ (.B1(_0626_),
    .Y(_0627_),
    .A1(_0602_),
    .A2(_0625_));
 sg13g2_o21ai_1 _1554_ (.B1(_0618_),
    .Y(_0628_),
    .A1(_0603_),
    .A2(_0619_));
 sg13g2_a22oi_1 _1555_ (.Y(_0629_),
    .B1(_0605_),
    .B2(_0616_),
    .A2(_0580_),
    .A1(_0504_));
 sg13g2_a21oi_1 _1556_ (.A1(_0101_),
    .A2(net171),
    .Y(_0630_),
    .B1(_0611_));
 sg13g2_nor2_1 _1557_ (.A(_0608_),
    .B(_0630_),
    .Y(_0631_));
 sg13g2_nor2_1 _1558_ (.A(_0613_),
    .B(_0615_),
    .Y(_0632_));
 sg13g2_nand2_1 _1559_ (.Y(_0633_),
    .A(_0608_),
    .B(_0630_));
 sg13g2_o21ai_1 _1560_ (.B1(_0633_),
    .Y(_0634_),
    .A1(_0631_),
    .A2(_0632_));
 sg13g2_xor2_1 _1561_ (.B(_0634_),
    .A(_0629_),
    .X(_0635_));
 sg13g2_xnor2_1 _1562_ (.Y(_0636_),
    .A(_0628_),
    .B(_0635_));
 sg13g2_xnor2_1 _1563_ (.Y(_0034_),
    .A(_0627_),
    .B(_0636_));
 sg13g2_a22oi_1 _1564_ (.Y(_0038_),
    .B1(_0192_),
    .B2(_0243_),
    .A2(_0139_),
    .A1(_0099_));
 sg13g2_nor2b_1 _1565_ (.A(\mixer_out[0] ),
    .B_N(net262),
    .Y(_0637_));
 sg13g2_xor2_1 _1566_ (.B(net262),
    .A(net245),
    .X(_0638_));
 sg13g2_nand2_1 _1567_ (.Y(_0639_),
    .A(net247),
    .B(_0638_));
 sg13g2_o21ai_1 _1568_ (.B1(net195),
    .Y(_0640_),
    .A1(net247),
    .A2(_0638_));
 sg13g2_nor2b_1 _1569_ (.A(net248),
    .B_N(_0639_),
    .Y(_0039_));
 sg13g2_and2_1 _1570_ (.A(\mixer_out[1] ),
    .B(\boxcar_filter[1] ),
    .X(_0641_));
 sg13g2_xor2_1 _1571_ (.B(\boxcar_filter[1] ),
    .A(\mixer_out[1] ),
    .X(_0642_));
 sg13g2_xnor2_1 _1572_ (.Y(_0643_),
    .A(_0016_),
    .B(_0642_));
 sg13g2_or2_1 _1573_ (.X(_0644_),
    .B(_0643_),
    .A(_0637_));
 sg13g2_xnor2_1 _1574_ (.Y(_0645_),
    .A(_0637_),
    .B(_0643_));
 sg13g2_or2_1 _1575_ (.X(_0646_),
    .B(_0645_),
    .A(_0639_));
 sg13g2_nand2_1 _1576_ (.Y(_0647_),
    .A(net198),
    .B(_0646_));
 sg13g2_a21oi_1 _1577_ (.A1(_0639_),
    .A2(_0645_),
    .Y(_0040_),
    .B1(_0647_));
 sg13g2_and2_1 _1578_ (.A(_0644_),
    .B(_0646_),
    .X(_0648_));
 sg13g2_o21ai_1 _1579_ (.B1(_0644_),
    .Y(_0649_),
    .A1(_0639_),
    .A2(_0645_));
 sg13g2_and2_1 _1580_ (.A(\boxcar_filter[2] ),
    .B(\mixer_out[2] ),
    .X(_0650_));
 sg13g2_xor2_1 _1581_ (.B(\mixer_out[2] ),
    .A(\boxcar_filter[2] ),
    .X(_0651_));
 sg13g2_xnor2_1 _1582_ (.Y(_0652_),
    .A(_0017_),
    .B(_0651_));
 sg13g2_a21oi_1 _1583_ (.A1(net324),
    .A2(_0642_),
    .Y(_0653_),
    .B1(_0641_));
 sg13g2_nor2_1 _1584_ (.A(_0652_),
    .B(_0653_),
    .Y(_0654_));
 sg13g2_xnor2_1 _1585_ (.Y(_0655_),
    .A(_0652_),
    .B(_0653_));
 sg13g2_inv_1 _1586_ (.Y(_0656_),
    .A(_0655_));
 sg13g2_o21ai_1 _1587_ (.B1(net198),
    .Y(_0657_),
    .A1(_0648_),
    .A2(_0655_));
 sg13g2_a21oi_1 _1588_ (.A1(_0648_),
    .A2(net325),
    .Y(_0041_),
    .B1(_0657_));
 sg13g2_a21oi_1 _1589_ (.A1(_0649_),
    .A2(_0656_),
    .Y(_0658_),
    .B1(_0654_));
 sg13g2_and2_1 _1590_ (.A(\boxcar_filter[3] ),
    .B(\mixer_out[3] ),
    .X(_0659_));
 sg13g2_xor2_1 _1591_ (.B(\mixer_out[3] ),
    .A(\boxcar_filter[3] ),
    .X(_0660_));
 sg13g2_xnor2_1 _1592_ (.Y(_0661_),
    .A(_0018_),
    .B(_0660_));
 sg13g2_a21oi_1 _1593_ (.A1(net319),
    .A2(_0651_),
    .Y(_0662_),
    .B1(_0650_));
 sg13g2_or2_1 _1594_ (.X(_0663_),
    .B(_0662_),
    .A(_0661_));
 sg13g2_xnor2_1 _1595_ (.Y(_0664_),
    .A(_0661_),
    .B(_0662_));
 sg13g2_or2_1 _1596_ (.X(_0665_),
    .B(_0664_),
    .A(_0658_));
 sg13g2_nand2_1 _1597_ (.Y(_0666_),
    .A(net198),
    .B(_0665_));
 sg13g2_a21oi_1 _1598_ (.A1(_0658_),
    .A2(net320),
    .Y(_0042_),
    .B1(_0666_));
 sg13g2_and2_1 _1599_ (.A(_0663_),
    .B(_0665_),
    .X(_0667_));
 sg13g2_o21ai_1 _1600_ (.B1(_0663_),
    .Y(_0668_),
    .A1(_0658_),
    .A2(_0664_));
 sg13g2_and2_1 _1601_ (.A(\boxcar_filter[4] ),
    .B(\mixer_out[4] ),
    .X(_0669_));
 sg13g2_xor2_1 _1602_ (.B(\mixer_out[4] ),
    .A(\boxcar_filter[4] ),
    .X(_0670_));
 sg13g2_xnor2_1 _1603_ (.Y(_0671_),
    .A(_0019_),
    .B(_0670_));
 sg13g2_a21oi_1 _1604_ (.A1(net322),
    .A2(_0660_),
    .Y(_0672_),
    .B1(_0659_));
 sg13g2_nor2_1 _1605_ (.A(_0671_),
    .B(_0672_),
    .Y(_0673_));
 sg13g2_xnor2_1 _1606_ (.Y(_0674_),
    .A(_0671_),
    .B(_0672_));
 sg13g2_inv_1 _1607_ (.Y(_0675_),
    .A(_0674_));
 sg13g2_o21ai_1 _1608_ (.B1(net198),
    .Y(_0676_),
    .A1(_0667_),
    .A2(_0674_));
 sg13g2_a21oi_1 _1609_ (.A1(_0667_),
    .A2(_0674_),
    .Y(_0043_),
    .B1(_0676_));
 sg13g2_a21o_1 _1610_ (.A2(_0675_),
    .A1(_0668_),
    .B1(_0673_),
    .X(_0677_));
 sg13g2_a21o_1 _1611_ (.A2(_0670_),
    .A1(_0019_),
    .B1(_0669_),
    .X(_0678_));
 sg13g2_and2_1 _1612_ (.A(\boxcar_filter[5] ),
    .B(\mixer_out[5] ),
    .X(_0679_));
 sg13g2_xor2_1 _1613_ (.B(\mixer_out[5] ),
    .A(\boxcar_filter[5] ),
    .X(_0680_));
 sg13g2_xnor2_1 _1614_ (.Y(_0681_),
    .A(net323),
    .B(_0680_));
 sg13g2_inv_1 _1615_ (.Y(_0682_),
    .A(_0681_));
 sg13g2_nor2_1 _1616_ (.A(_0678_),
    .B(_0682_),
    .Y(_0683_));
 sg13g2_xnor2_1 _1617_ (.Y(_0684_),
    .A(_0678_),
    .B(_0681_));
 sg13g2_o21ai_1 _1618_ (.B1(net197),
    .Y(_0685_),
    .A1(_0677_),
    .A2(_0684_));
 sg13g2_a21oi_1 _1619_ (.A1(_0677_),
    .A2(_0684_),
    .Y(_0044_),
    .B1(_0685_));
 sg13g2_and2_1 _1620_ (.A(\boxcar_filter[6] ),
    .B(\mixer_out[6] ),
    .X(_0686_));
 sg13g2_xor2_1 _1621_ (.B(\mixer_out[6] ),
    .A(\boxcar_filter[6] ),
    .X(_0687_));
 sg13g2_xnor2_1 _1622_ (.Y(_0688_),
    .A(_0021_),
    .B(_0687_));
 sg13g2_a21oi_1 _1623_ (.A1(net326),
    .A2(_0680_),
    .Y(_0689_),
    .B1(_0679_));
 sg13g2_nor2_1 _1624_ (.A(_0688_),
    .B(_0689_),
    .Y(_0690_));
 sg13g2_xnor2_1 _1625_ (.Y(_0691_),
    .A(_0688_),
    .B(_0689_));
 sg13g2_a221oi_1 _1626_ (.B2(_0682_),
    .C1(_0673_),
    .B1(_0678_),
    .A1(_0668_),
    .Y(_0692_),
    .A2(_0675_));
 sg13g2_o21ai_1 _1627_ (.B1(_0691_),
    .Y(_0693_),
    .A1(_0683_),
    .A2(_0692_));
 sg13g2_nor3_2 _1628_ (.A(_0683_),
    .B(_0691_),
    .C(_0692_),
    .Y(_0694_));
 sg13g2_nand2_1 _1629_ (.Y(_0695_),
    .A(net197),
    .B(_0693_));
 sg13g2_nor2_1 _1630_ (.A(_0694_),
    .B(_0695_),
    .Y(_0045_));
 sg13g2_and2_1 _1631_ (.A(\boxcar_filter[7] ),
    .B(\mixer_out[7] ),
    .X(_0696_));
 sg13g2_xor2_1 _1632_ (.B(\mixer_out[7] ),
    .A(\boxcar_filter[7] ),
    .X(_0697_));
 sg13g2_xnor2_1 _1633_ (.Y(_0698_),
    .A(_0022_),
    .B(_0697_));
 sg13g2_a21oi_1 _1634_ (.A1(_0021_),
    .A2(_0687_),
    .Y(_0699_),
    .B1(_0686_));
 sg13g2_nor2_1 _1635_ (.A(_0698_),
    .B(_0699_),
    .Y(_0700_));
 sg13g2_xnor2_1 _1636_ (.Y(_0701_),
    .A(_0698_),
    .B(_0699_));
 sg13g2_inv_1 _1637_ (.Y(_0702_),
    .A(_0701_));
 sg13g2_nor3_1 _1638_ (.A(_0690_),
    .B(_0694_),
    .C(_0702_),
    .Y(_0703_));
 sg13g2_o21ai_1 _1639_ (.B1(_0702_),
    .Y(_0704_),
    .A1(_0690_),
    .A2(_0694_));
 sg13g2_nand2_1 _1640_ (.Y(_0705_),
    .A(net197),
    .B(_0704_));
 sg13g2_nor2_1 _1641_ (.A(_0703_),
    .B(_0705_),
    .Y(_0046_));
 sg13g2_nor2b_1 _1642_ (.A(_0700_),
    .B_N(_0704_),
    .Y(_0706_));
 sg13g2_a21oi_1 _1643_ (.A1(net302),
    .A2(_0697_),
    .Y(_0707_),
    .B1(_0696_));
 sg13g2_nor2_1 _1644_ (.A(net287),
    .B(_0707_),
    .Y(_0708_));
 sg13g2_xnor2_1 _1645_ (.Y(_0709_),
    .A(net287),
    .B(_0707_));
 sg13g2_and2_1 _1646_ (.A(_0706_),
    .B(_0709_),
    .X(_0710_));
 sg13g2_nor2_1 _1647_ (.A(_0706_),
    .B(_0709_),
    .Y(_0711_));
 sg13g2_nor3_1 _1648_ (.A(net193),
    .B(_0710_),
    .C(_0711_),
    .Y(_0047_));
 sg13g2_nor2_1 _1649_ (.A(_0708_),
    .B(_0711_),
    .Y(_0712_));
 sg13g2_xor2_1 _1650_ (.B(net249),
    .A(net287),
    .X(_0713_));
 sg13g2_o21ai_1 _1651_ (.B1(net199),
    .Y(_0714_),
    .A1(_0712_),
    .A2(_0713_));
 sg13g2_a21oi_1 _1652_ (.A1(_0712_),
    .A2(_0713_),
    .Y(_0048_),
    .B1(_0714_));
 sg13g2_and2_1 _1653_ (.A(net245),
    .B(net194),
    .X(_0049_));
 sg13g2_and2_1 _1654_ (.A(net240),
    .B(net198),
    .X(_0050_));
 sg13g2_and2_1 _1655_ (.A(net241),
    .B(net199),
    .X(_0051_));
 sg13g2_and2_1 _1656_ (.A(net246),
    .B(net194),
    .X(_0052_));
 sg13g2_and2_1 _1657_ (.A(net269),
    .B(net194),
    .X(_0053_));
 sg13g2_and2_1 _1658_ (.A(net276),
    .B(net196),
    .X(_0054_));
 sg13g2_and2_1 _1659_ (.A(net258),
    .B(net196),
    .X(_0055_));
 sg13g2_and2_1 _1660_ (.A(net277),
    .B(net197),
    .X(_0056_));
 sg13g2_and2_1 _1661_ (.A(net194),
    .B(net209),
    .X(_0057_));
 sg13g2_and2_1 _1662_ (.A(net198),
    .B(net216),
    .X(_0058_));
 sg13g2_and2_1 _1663_ (.A(net199),
    .B(net224),
    .X(_0059_));
 sg13g2_and2_1 _1664_ (.A(net194),
    .B(net219),
    .X(_0060_));
 sg13g2_and2_1 _1665_ (.A(net195),
    .B(net215),
    .X(_0061_));
 sg13g2_and2_1 _1666_ (.A(net196),
    .B(net226),
    .X(_0062_));
 sg13g2_and2_1 _1667_ (.A(net196),
    .B(net227),
    .X(_0063_));
 sg13g2_and2_1 _1668_ (.A(net196),
    .B(net217),
    .X(_0064_));
 sg13g2_and2_1 _1669_ (.A(net194),
    .B(net208),
    .X(_0065_));
 sg13g2_and2_1 _1670_ (.A(net198),
    .B(net220),
    .X(_0066_));
 sg13g2_and2_1 _1671_ (.A(net199),
    .B(net149),
    .X(_0067_));
 sg13g2_and2_1 _1672_ (.A(net194),
    .B(net212),
    .X(_0068_));
 sg13g2_and2_1 _1673_ (.A(net194),
    .B(net222),
    .X(_0069_));
 sg13g2_and2_1 _1674_ (.A(net196),
    .B(net218),
    .X(_0070_));
 sg13g2_and2_1 _1675_ (.A(net196),
    .B(net213),
    .X(_0071_));
 sg13g2_and2_1 _1676_ (.A(net197),
    .B(net223),
    .X(_0072_));
 sg13g2_and2_1 _1677_ (.A(net195),
    .B(net205),
    .X(_0073_));
 sg13g2_and2_1 _1678_ (.A(net201),
    .B(net214),
    .X(_0074_));
 sg13g2_and2_1 _1679_ (.A(net198),
    .B(net225),
    .X(_0075_));
 sg13g2_and2_1 _1680_ (.A(net195),
    .B(net207),
    .X(_0076_));
 sg13g2_and2_1 _1681_ (.A(net195),
    .B(net211),
    .X(_0077_));
 sg13g2_and2_1 _1682_ (.A(net196),
    .B(net210),
    .X(_0078_));
 sg13g2_and2_1 _1683_ (.A(net197),
    .B(net221),
    .X(_0079_));
 sg13g2_and2_1 _1684_ (.A(net197),
    .B(net206),
    .X(_0080_));
 sg13g2_or2_1 _1685_ (.X(_0715_),
    .B(net289),
    .A(\inst_sine_B.phase[0] ));
 sg13g2_nand2_1 _1686_ (.Y(_0716_),
    .A(\inst_sine_B.phase[0] ),
    .B(net289));
 sg13g2_and3_1 _1687_ (.X(_0082_),
    .A(net1),
    .B(net290),
    .C(_0716_));
 sg13g2_xnor2_1 _1688_ (.Y(_0717_),
    .A(\inst_sine_B.phase[1] ),
    .B(net300));
 sg13g2_and2_1 _1689_ (.A(_0716_),
    .B(_0717_),
    .X(_0718_));
 sg13g2_nor2_1 _1690_ (.A(_0716_),
    .B(_0717_),
    .Y(_0719_));
 sg13g2_nor3_1 _1691_ (.A(net193),
    .B(_0718_),
    .C(_0719_),
    .Y(_0083_));
 sg13g2_xnor2_1 _1692_ (.Y(_0720_),
    .A(\inst_sine_B.phase[2] ),
    .B(net315));
 sg13g2_a21oi_1 _1693_ (.A1(\inst_sine_B.phase[1] ),
    .A2(net300),
    .Y(_0721_),
    .B1(_0719_));
 sg13g2_and2_1 _1694_ (.A(net316),
    .B(_0721_),
    .X(_0722_));
 sg13g2_nor2_1 _1695_ (.A(_0720_),
    .B(_0721_),
    .Y(_0723_));
 sg13g2_nor3_1 _1696_ (.A(net193),
    .B(_0722_),
    .C(_0723_),
    .Y(_0084_));
 sg13g2_nand2_1 _1697_ (.Y(_0724_),
    .A(\inst_sine_B.phase[3] ),
    .B(net280));
 sg13g2_xnor2_1 _1698_ (.Y(_0725_),
    .A(\inst_sine_B.phase[3] ),
    .B(net280));
 sg13g2_a21oi_1 _1699_ (.A1(\inst_sine_B.phase[2] ),
    .A2(\phase_incr_B[2] ),
    .Y(_0726_),
    .B1(_0723_));
 sg13g2_or2_1 _1700_ (.X(_0727_),
    .B(_0726_),
    .A(_0725_));
 sg13g2_nand2_1 _1701_ (.Y(_0728_),
    .A(net201),
    .B(_0727_));
 sg13g2_a21oi_1 _1702_ (.A1(net281),
    .A2(_0726_),
    .Y(_0085_),
    .B1(_0728_));
 sg13g2_xnor2_1 _1703_ (.Y(_0729_),
    .A(\inst_sine_B.phase[4] ),
    .B(net307));
 sg13g2_and2_1 _1704_ (.A(_0724_),
    .B(_0727_),
    .X(_0730_));
 sg13g2_and2_1 _1705_ (.A(net308),
    .B(_0730_),
    .X(_0731_));
 sg13g2_nor2_1 _1706_ (.A(net308),
    .B(_0730_),
    .Y(_0732_));
 sg13g2_nor3_1 _1707_ (.A(net193),
    .B(_0731_),
    .C(_0732_),
    .Y(_0086_));
 sg13g2_nand2_1 _1708_ (.Y(_0733_),
    .A(net309),
    .B(net283));
 sg13g2_xnor2_1 _1709_ (.Y(_0734_),
    .A(\inst_sine_B.phase[5] ),
    .B(net283));
 sg13g2_a21oi_1 _1710_ (.A1(\inst_sine_B.phase[4] ),
    .A2(\phase_incr_B[4] ),
    .Y(_0735_),
    .B1(_0732_));
 sg13g2_or2_1 _1711_ (.X(_0736_),
    .B(_0735_),
    .A(_0734_));
 sg13g2_nand2_1 _1712_ (.Y(_0737_),
    .A(net201),
    .B(_0736_));
 sg13g2_a21oi_1 _1713_ (.A1(net284),
    .A2(_0735_),
    .Y(_0087_),
    .B1(_0737_));
 sg13g2_nand2_1 _1714_ (.Y(_0738_),
    .A(_0733_),
    .B(_0736_));
 sg13g2_nor2_1 _1715_ (.A(net187),
    .B(_0738_),
    .Y(_0739_));
 sg13g2_and2_1 _1716_ (.A(net187),
    .B(_0738_),
    .X(_0740_));
 sg13g2_nor3_1 _1717_ (.A(net193),
    .B(_0739_),
    .C(_0740_),
    .Y(_0088_));
 sg13g2_xnor2_1 _1718_ (.Y(_0741_),
    .A(net259),
    .B(_0740_));
 sg13g2_nor2_1 _1719_ (.A(net193),
    .B(_0741_),
    .Y(_0089_));
 sg13g2_nor2_1 _1720_ (.A(_0099_),
    .B(_0193_),
    .Y(_0090_));
 sg13g2_or2_1 _1721_ (.X(_0742_),
    .B(net295),
    .A(\inst_sine_A.phase[0] ));
 sg13g2_nand2_1 _1722_ (.Y(_0743_),
    .A(\inst_sine_A.phase[0] ),
    .B(net295));
 sg13g2_and3_1 _1723_ (.X(_0091_),
    .A(net201),
    .B(net296),
    .C(_0743_));
 sg13g2_xnor2_1 _1724_ (.Y(_0744_),
    .A(\inst_sine_A.phase[1] ),
    .B(net303));
 sg13g2_and2_1 _1725_ (.A(_0743_),
    .B(net304),
    .X(_0745_));
 sg13g2_nor2_1 _1726_ (.A(_0743_),
    .B(_0744_),
    .Y(_0746_));
 sg13g2_nor3_1 _1727_ (.A(_0105_),
    .B(net305),
    .C(_0746_),
    .Y(_0092_));
 sg13g2_xnor2_1 _1728_ (.Y(_0747_),
    .A(\inst_sine_A.phase[2] ),
    .B(net310));
 sg13g2_a21oi_1 _1729_ (.A1(\inst_sine_A.phase[1] ),
    .A2(net303),
    .Y(_0748_),
    .B1(_0746_));
 sg13g2_and2_1 _1730_ (.A(net311),
    .B(_0748_),
    .X(_0749_));
 sg13g2_nor2_1 _1731_ (.A(_0747_),
    .B(_0748_),
    .Y(_0750_));
 sg13g2_nor3_1 _1732_ (.A(_0105_),
    .B(net312),
    .C(_0750_),
    .Y(_0093_));
 sg13g2_nand2_1 _1733_ (.Y(_0751_),
    .A(\inst_sine_A.phase[3] ),
    .B(net292));
 sg13g2_xnor2_1 _1734_ (.Y(_0752_),
    .A(\inst_sine_A.phase[3] ),
    .B(net292));
 sg13g2_a21oi_1 _1735_ (.A1(\inst_sine_A.phase[2] ),
    .A2(\phase_incr_A[2] ),
    .Y(_0753_),
    .B1(_0750_));
 sg13g2_or2_1 _1736_ (.X(_0754_),
    .B(_0753_),
    .A(_0752_));
 sg13g2_nand2_1 _1737_ (.Y(_0755_),
    .A(net201),
    .B(_0754_));
 sg13g2_a21oi_1 _1738_ (.A1(net293),
    .A2(_0753_),
    .Y(_0094_),
    .B1(_0755_));
 sg13g2_xnor2_1 _1739_ (.Y(_0756_),
    .A(net298),
    .B(net314));
 sg13g2_and2_1 _1740_ (.A(_0751_),
    .B(_0754_),
    .X(_0757_));
 sg13g2_and2_1 _1741_ (.A(_0756_),
    .B(_0757_),
    .X(_0758_));
 sg13g2_nor2_1 _1742_ (.A(_0756_),
    .B(_0757_),
    .Y(_0759_));
 sg13g2_nor3_1 _1743_ (.A(net193),
    .B(_0758_),
    .C(_0759_),
    .Y(_0095_));
 sg13g2_nand2_1 _1744_ (.Y(_0760_),
    .A(net286),
    .B(net272));
 sg13g2_xnor2_1 _1745_ (.Y(_0761_),
    .A(\inst_sine_A.phase[5] ),
    .B(net272));
 sg13g2_a21oi_1 _1746_ (.A1(\inst_sine_A.phase[4] ),
    .A2(\phase_incr_A[4] ),
    .Y(_0762_),
    .B1(_0759_));
 sg13g2_or2_1 _1747_ (.X(_0763_),
    .B(_0762_),
    .A(_0761_));
 sg13g2_nand2_1 _1748_ (.Y(_0764_),
    .A(net201),
    .B(_0763_));
 sg13g2_a21oi_1 _1749_ (.A1(net273),
    .A2(_0762_),
    .Y(_0096_),
    .B1(_0764_));
 sg13g2_nand2_1 _1750_ (.Y(_0765_),
    .A(net157),
    .B(\phase_incr_A[6] ));
 sg13g2_xnor2_1 _1751_ (.Y(_0766_),
    .A(net157),
    .B(net318));
 sg13g2_nand3_1 _1752_ (.B(_0763_),
    .C(_0766_),
    .A(_0760_),
    .Y(_0767_));
 sg13g2_a21o_1 _1753_ (.A2(_0763_),
    .A1(_0760_),
    .B1(_0766_),
    .X(_0768_));
 sg13g2_and3_1 _1754_ (.X(_0097_),
    .A(net201),
    .B(_0767_),
    .C(_0768_));
 sg13g2_and3_1 _1755_ (.X(_0769_),
    .A(net202),
    .B(_0765_),
    .C(_0768_));
 sg13g2_a21oi_1 _1756_ (.A1(_0765_),
    .A2(_0768_),
    .Y(_0770_),
    .B1(net202));
 sg13g2_nor3_1 _1757_ (.A(net193),
    .B(_0769_),
    .C(net203),
    .Y(_0098_));
 sg13g2_buf_1 _1758_ (.A(net251),
    .X(_0081_));
 sg13g2_dfrbp_1 _1759_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net36),
    .D(_0038_),
    .Q_N(_0826_),
    .Q(\sine_Breg[6] ));
 sg13g2_dfrbp_1 _1760_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net37),
    .D(_0000_),
    .Q_N(_0827_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _1761_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net38),
    .D(net271),
    .Q_N(_0828_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1762_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net39),
    .D(net265),
    .Q_N(_0829_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1763_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net40),
    .D(net279),
    .Q_N(_0830_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _1764_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net41),
    .D(net267),
    .Q_N(_0831_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _1765_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net42),
    .D(net261),
    .Q_N(_0832_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1766_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net85),
    .D(net288),
    .Q_N(_0833_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1767_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net35),
    .D(net250),
    .Q_N(_0825_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _1768_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net44),
    .D(_0039_),
    .Q_N(_0824_),
    .Q(\boxcar_filter[0] ));
 sg13g2_dfrbp_1 _1769_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net43),
    .D(net263),
    .Q_N(_0823_),
    .Q(\boxcar_filter[1] ));
 sg13g2_dfrbp_1 _1770_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net34),
    .D(_0041_),
    .Q_N(_0822_),
    .Q(\boxcar_filter[2] ));
 sg13g2_dfrbp_1 _1771_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net147),
    .D(net321),
    .Q_N(_0821_),
    .Q(\boxcar_filter[3] ));
 sg13g2_dfrbp_1 _1772_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net146),
    .D(_0043_),
    .Q_N(_0820_),
    .Q(\boxcar_filter[4] ));
 sg13g2_dfrbp_1 _1773_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net145),
    .D(_0044_),
    .Q_N(_0819_),
    .Q(\boxcar_filter[5] ));
 sg13g2_dfrbp_1 _1774_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net144),
    .D(_0045_),
    .Q_N(_0818_),
    .Q(\boxcar_filter[6] ));
 sg13g2_dfrbp_1 _1775_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net143),
    .D(_0046_),
    .Q_N(_0817_),
    .Q(\boxcar_filter[7] ));
 sg13g2_dfrbp_1 _1776_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net142),
    .D(_0047_),
    .Q_N(_0816_),
    .Q(\boxcar_filter[8] ));
 sg13g2_dfrbp_1 _1777_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net141),
    .D(_0048_),
    .Q_N(_0815_),
    .Q(\boxcar_filter[9] ));
 sg13g2_dfrbp_1 _1778_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net140),
    .D(_0049_),
    .Q_N(_0814_),
    .Q(\boxcar_storage[1][0] ));
 sg13g2_dfrbp_1 _1779_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net132),
    .D(_0050_),
    .Q_N(_0813_),
    .Q(\boxcar_storage[1][1] ));
 sg13g2_dfrbp_1 _1780_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net109),
    .D(_0051_),
    .Q_N(_0812_),
    .Q(\boxcar_storage[1][2] ));
 sg13g2_dfrbp_1 _1781_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net108),
    .D(_0052_),
    .Q_N(_0811_),
    .Q(\boxcar_storage[1][3] ));
 sg13g2_dfrbp_1 _1782_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net107),
    .D(_0053_),
    .Q_N(_0810_),
    .Q(\boxcar_storage[1][4] ));
 sg13g2_dfrbp_1 _1783_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net106),
    .D(_0054_),
    .Q_N(_0809_),
    .Q(\boxcar_storage[1][5] ));
 sg13g2_dfrbp_1 _1784_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net105),
    .D(_0055_),
    .Q_N(_0808_),
    .Q(\boxcar_storage[1][6] ));
 sg13g2_dfrbp_1 _1785_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net104),
    .D(_0056_),
    .Q_N(_0807_),
    .Q(\boxcar_storage[1][7] ));
 sg13g2_dfrbp_1 _1786_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net103),
    .D(_0057_),
    .Q_N(_0806_),
    .Q(\boxcar_storage[2][0] ));
 sg13g2_dfrbp_1 _1787_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net102),
    .D(_0058_),
    .Q_N(_0805_),
    .Q(\boxcar_storage[2][1] ));
 sg13g2_dfrbp_1 _1788_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net101),
    .D(_0059_),
    .Q_N(_0804_),
    .Q(\boxcar_storage[2][2] ));
 sg13g2_dfrbp_1 _1789_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net84),
    .D(_0060_),
    .Q_N(_0803_),
    .Q(\boxcar_storage[2][3] ));
 sg13g2_dfrbp_1 _1790_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net83),
    .D(_0061_),
    .Q_N(_0802_),
    .Q(\boxcar_storage[2][4] ));
 sg13g2_dfrbp_1 _1791_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net82),
    .D(_0062_),
    .Q_N(_0801_),
    .Q(\boxcar_storage[2][5] ));
 sg13g2_dfrbp_1 _1792_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net81),
    .D(_0063_),
    .Q_N(_0800_),
    .Q(\boxcar_storage[2][6] ));
 sg13g2_dfrbp_1 _1793_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net80),
    .D(_0064_),
    .Q_N(_0799_),
    .Q(\boxcar_storage[2][7] ));
 sg13g2_dfrbp_1 _1794_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net79),
    .D(_0065_),
    .Q_N(_0798_),
    .Q(\boxcar_storage[3][0] ));
 sg13g2_dfrbp_1 _1795_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net78),
    .D(_0066_),
    .Q_N(_0797_),
    .Q(\boxcar_storage[3][1] ));
 sg13g2_dfrbp_1 _1796_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net77),
    .D(_0067_),
    .Q_N(_0796_),
    .Q(\boxcar_storage[3][2] ));
 sg13g2_dfrbp_1 _1797_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net76),
    .D(_0068_),
    .Q_N(_0795_),
    .Q(\boxcar_storage[3][3] ));
 sg13g2_dfrbp_1 _1798_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net75),
    .D(_0069_),
    .Q_N(_0794_),
    .Q(\boxcar_storage[3][4] ));
 sg13g2_dfrbp_1 _1799_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net74),
    .D(_0070_),
    .Q_N(_0793_),
    .Q(\boxcar_storage[3][5] ));
 sg13g2_dfrbp_1 _1800_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net73),
    .D(_0071_),
    .Q_N(_0792_),
    .Q(\boxcar_storage[3][6] ));
 sg13g2_dfrbp_1 _1801_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net72),
    .D(_0072_),
    .Q_N(_0791_),
    .Q(\boxcar_storage[3][7] ));
 sg13g2_dfrbp_1 _1802_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net71),
    .D(_0073_),
    .Q_N(_0790_),
    .Q(\boxcar_storage[4][0] ));
 sg13g2_dfrbp_1 _1803_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net70),
    .D(_0074_),
    .Q_N(_0016_),
    .Q(\boxcar_storage[4][1] ));
 sg13g2_dfrbp_1 _1804_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net69),
    .D(_0075_),
    .Q_N(_0017_),
    .Q(\boxcar_storage[4][2] ));
 sg13g2_dfrbp_1 _1805_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net68),
    .D(_0076_),
    .Q_N(_0018_),
    .Q(\boxcar_storage[4][3] ));
 sg13g2_dfrbp_1 _1806_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net67),
    .D(_0077_),
    .Q_N(_0019_),
    .Q(\boxcar_storage[4][4] ));
 sg13g2_dfrbp_1 _1807_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net66),
    .D(_0078_),
    .Q_N(_0020_),
    .Q(\boxcar_storage[4][5] ));
 sg13g2_dfrbp_1 _1808_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net65),
    .D(_0079_),
    .Q_N(_0021_),
    .Q(\boxcar_storage[4][6] ));
 sg13g2_dfrbp_1 _1809_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net86),
    .D(_0080_),
    .Q_N(_0022_),
    .Q(\boxcar_storage[4][7] ));
 sg13g2_dfrbp_1 _1810_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net87),
    .D(_0035_),
    .Q_N(_0771_),
    .Q(\product[7] ));
 sg13g2_dfrbp_1 _1811_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net88),
    .D(_0036_),
    .Q_N(_0834_),
    .Q(\product[8] ));
 sg13g2_dfrbp_1 _1812_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net89),
    .D(_0037_),
    .Q_N(_0835_),
    .Q(\product[9] ));
 sg13g2_dfrbp_1 _1813_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net90),
    .D(_0030_),
    .Q_N(_0836_),
    .Q(\product[10] ));
 sg13g2_dfrbp_1 _1814_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net91),
    .D(_0031_),
    .Q_N(_0837_),
    .Q(\product[11] ));
 sg13g2_dfrbp_1 _1815_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net92),
    .D(_0032_),
    .Q_N(_0838_),
    .Q(\product[12] ));
 sg13g2_dfrbp_1 _1816_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net93),
    .D(_0033_),
    .Q_N(_0839_),
    .Q(\product[13] ));
 sg13g2_dfrbp_1 _1817_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net94),
    .D(_0034_),
    .Q_N(_0840_),
    .Q(\product[14] ));
 sg13g2_dfrbp_1 _1818_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net95),
    .D(net148),
    .Q_N(_0841_),
    .Q(\mixer_out[0] ));
 sg13g2_dfrbp_1 _1819_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net96),
    .D(net239),
    .Q_N(_0842_),
    .Q(\mixer_out[1] ));
 sg13g2_dfrbp_1 _1820_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net97),
    .D(net244),
    .Q_N(_0843_),
    .Q(\mixer_out[2] ));
 sg13g2_dfrbp_1 _1821_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net98),
    .D(net237),
    .Q_N(_0844_),
    .Q(\mixer_out[3] ));
 sg13g2_dfrbp_1 _1822_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net99),
    .D(net231),
    .Q_N(_0845_),
    .Q(\mixer_out[4] ));
 sg13g2_dfrbp_1 _1823_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net100),
    .D(net235),
    .Q_N(_0846_),
    .Q(\mixer_out[5] ));
 sg13g2_dfrbp_1 _1824_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net110),
    .D(net233),
    .Q_N(_0847_),
    .Q(\mixer_out[6] ));
 sg13g2_dfrbp_1 _1825_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net64),
    .D(net229),
    .Q_N(_0789_),
    .Q(\mixer_out[7] ));
 sg13g2_dfrbp_1 _1826_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net63),
    .D(_0081_),
    .Q_N(_0788_),
    .Q(\sine_Areg[7] ));
 sg13g2_dfrbp_1 _1827_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net62),
    .D(net291),
    .Q_N(_0787_),
    .Q(\inst_sine_B.phase[0] ));
 sg13g2_dfrbp_1 _1828_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net61),
    .D(net301),
    .Q_N(_0786_),
    .Q(\inst_sine_B.phase[1] ));
 sg13g2_dfrbp_1 _1829_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net60),
    .D(net317),
    .Q_N(_0785_),
    .Q(\inst_sine_B.phase[2] ));
 sg13g2_dfrbp_1 _1830_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net59),
    .D(net282),
    .Q_N(_0784_),
    .Q(\inst_sine_B.phase[3] ));
 sg13g2_dfrbp_1 _1831_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net58),
    .D(_0086_),
    .Q_N(_0783_),
    .Q(\inst_sine_B.phase[4] ));
 sg13g2_dfrbp_1 _1832_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net57),
    .D(net285),
    .Q_N(_0782_),
    .Q(\inst_sine_B.phase[5] ));
 sg13g2_dfrbp_1 _1833_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net56),
    .D(_0088_),
    .Q_N(_0781_),
    .Q(\inst_sine_B.phase[6] ));
 sg13g2_dfrbp_1 _1834_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net111),
    .D(_0089_),
    .Q_N(_0848_),
    .Q(\inst_sine_B.phase[7] ));
 sg13g2_dfrbp_1 _1835_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net112),
    .D(net9),
    .Q_N(_0849_),
    .Q(filter_on));
 sg13g2_dfrbp_1 _1836_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net113),
    .D(net2),
    .Q_N(_0850_),
    .Q(\phase_incr_A[0] ));
 sg13g2_dfrbp_1 _1837_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net114),
    .D(net3),
    .Q_N(_0851_),
    .Q(\phase_incr_A[1] ));
 sg13g2_dfrbp_1 _1838_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net115),
    .D(net4),
    .Q_N(_0852_),
    .Q(\phase_incr_A[2] ));
 sg13g2_dfrbp_1 _1839_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net116),
    .D(net5),
    .Q_N(_0853_),
    .Q(\phase_incr_A[3] ));
 sg13g2_dfrbp_1 _1840_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net117),
    .D(net6),
    .Q_N(_0854_),
    .Q(\phase_incr_A[4] ));
 sg13g2_dfrbp_1 _1841_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net118),
    .D(net7),
    .Q_N(_0855_),
    .Q(\phase_incr_A[5] ));
 sg13g2_dfrbp_1 _1842_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net119),
    .D(net8),
    .Q_N(_0856_),
    .Q(\phase_incr_A[6] ));
 sg13g2_dfrbp_1 _1843_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net120),
    .D(net17),
    .Q_N(_0857_),
    .Q(bypass_B));
 sg13g2_dfrbp_1 _1844_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net121),
    .D(net16),
    .Q_N(_0014_),
    .Q(lowamp_B));
 sg13g2_dfrbp_1 _1845_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net122),
    .D(net10),
    .Q_N(_0858_),
    .Q(\phase_incr_B[0] ));
 sg13g2_dfrbp_1 _1846_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net123),
    .D(net11),
    .Q_N(_0859_),
    .Q(\phase_incr_B[1] ));
 sg13g2_dfrbp_1 _1847_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net124),
    .D(net12),
    .Q_N(_0860_),
    .Q(\phase_incr_B[2] ));
 sg13g2_dfrbp_1 _1848_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net125),
    .D(net13),
    .Q_N(_0861_),
    .Q(\phase_incr_B[3] ));
 sg13g2_dfrbp_1 _1849_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net126),
    .D(net14),
    .Q_N(_0862_),
    .Q(\phase_incr_B[4] ));
 sg13g2_dfrbp_1 _1850_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net127),
    .D(net15),
    .Q_N(_0863_),
    .Q(\phase_incr_B[5] ));
 sg13g2_dfrbp_1 _1851_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net128),
    .D(net256),
    .Q_N(_0864_),
    .Q(\sine_Breg[0] ));
 sg13g2_dfrbp_1 _1852_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net129),
    .D(_0009_),
    .Q_N(_0865_),
    .Q(\sine_Breg[1] ));
 sg13g2_dfrbp_1 _1853_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net130),
    .D(net254),
    .Q_N(_0866_),
    .Q(\sine_Breg[2] ));
 sg13g2_dfrbp_1 _1854_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net131),
    .D(_0011_),
    .Q_N(_0867_),
    .Q(\sine_Breg[3] ));
 sg13g2_dfrbp_1 _1855_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net133),
    .D(_0012_),
    .Q_N(_0868_),
    .Q(\sine_Breg[4] ));
 sg13g2_dfrbp_1 _1856_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net55),
    .D(_0013_),
    .Q_N(_0780_),
    .Q(\sine_Breg[5] ));
 sg13g2_dfrbp_1 _1857_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net134),
    .D(_0090_),
    .Q_N(_0869_),
    .Q(\sine_Breg[7] ));
 sg13g2_dfrbp_1 _1858_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net135),
    .D(\inst_sine_A.sample[0] ),
    .Q_N(_0870_),
    .Q(\sine_Areg[0] ));
 sg13g2_dfrbp_1 _1859_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net136),
    .D(\inst_sine_A.sample[1] ),
    .Q_N(_0871_),
    .Q(\sine_Areg[1] ));
 sg13g2_dfrbp_1 _1860_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net137),
    .D(\inst_sine_A.sample[2] ),
    .Q_N(_0872_),
    .Q(\sine_Areg[2] ));
 sg13g2_dfrbp_1 _1861_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net138),
    .D(\inst_sine_A.sample[3] ),
    .Q_N(_0873_),
    .Q(\sine_Areg[3] ));
 sg13g2_dfrbp_1 _1862_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net139),
    .D(\inst_sine_A.sample[4] ),
    .Q_N(_0874_),
    .Q(\sine_Areg[4] ));
 sg13g2_dfrbp_1 _1863_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net45),
    .D(\inst_sine_A.sample[5] ),
    .Q_N(_0875_),
    .Q(\sine_Areg[5] ));
 sg13g2_dfrbp_1 _1864_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net54),
    .D(\inst_sine_A.sample[6] ),
    .Q_N(_0779_),
    .Q(\sine_Areg[6] ));
 sg13g2_dfrbp_1 _1865_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net53),
    .D(net297),
    .Q_N(_0778_),
    .Q(\inst_sine_A.phase[0] ));
 sg13g2_dfrbp_1 _1866_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net52),
    .D(net306),
    .Q_N(_0777_),
    .Q(\inst_sine_A.phase[1] ));
 sg13g2_dfrbp_1 _1867_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net51),
    .D(net313),
    .Q_N(_0776_),
    .Q(\inst_sine_A.phase[2] ));
 sg13g2_dfrbp_1 _1868_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net50),
    .D(net294),
    .Q_N(_0775_),
    .Q(\inst_sine_A.phase[3] ));
 sg13g2_dfrbp_1 _1869_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net49),
    .D(_0095_),
    .Q_N(_0774_),
    .Q(\inst_sine_A.phase[4] ));
 sg13g2_dfrbp_1 _1870_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net48),
    .D(net274),
    .Q_N(_0773_),
    .Q(\inst_sine_A.phase[5] ));
 sg13g2_dfrbp_1 _1871_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net47),
    .D(_0097_),
    .Q_N(_0772_),
    .Q(\inst_sine_A.phase[6] ));
 sg13g2_dfrbp_1 _1872_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net46),
    .D(net204),
    .Q_N(_0015_),
    .Q(\inst_sine_A.phase[7] ));
 sg13g2_tiehi _1767__35 (.L_HI(net35));
 sg13g2_tiehi _1759__36 (.L_HI(net36));
 sg13g2_tiehi _1760__37 (.L_HI(net37));
 sg13g2_tiehi _1761__38 (.L_HI(net38));
 sg13g2_tiehi _1762__39 (.L_HI(net39));
 sg13g2_tiehi _1763__40 (.L_HI(net40));
 sg13g2_tiehi _1764__41 (.L_HI(net41));
 sg13g2_tiehi _1765__42 (.L_HI(net42));
 sg13g2_tiehi _1769__43 (.L_HI(net43));
 sg13g2_tiehi _1768__44 (.L_HI(net44));
 sg13g2_tiehi _1863__45 (.L_HI(net45));
 sg13g2_tiehi _1872__46 (.L_HI(net46));
 sg13g2_tiehi _1871__47 (.L_HI(net47));
 sg13g2_tiehi _1870__48 (.L_HI(net48));
 sg13g2_tiehi _1869__49 (.L_HI(net49));
 sg13g2_tiehi _1868__50 (.L_HI(net50));
 sg13g2_tiehi _1867__51 (.L_HI(net51));
 sg13g2_tiehi _1866__52 (.L_HI(net52));
 sg13g2_tiehi _1865__53 (.L_HI(net53));
 sg13g2_tiehi _1864__54 (.L_HI(net54));
 sg13g2_tiehi _1856__55 (.L_HI(net55));
 sg13g2_tiehi _1833__56 (.L_HI(net56));
 sg13g2_tiehi _1832__57 (.L_HI(net57));
 sg13g2_tiehi _1831__58 (.L_HI(net58));
 sg13g2_tiehi _1830__59 (.L_HI(net59));
 sg13g2_tiehi _1829__60 (.L_HI(net60));
 sg13g2_tiehi _1828__61 (.L_HI(net61));
 sg13g2_tiehi _1827__62 (.L_HI(net62));
 sg13g2_tiehi _1826__63 (.L_HI(net63));
 sg13g2_tiehi _1825__64 (.L_HI(net64));
 sg13g2_tiehi _1808__65 (.L_HI(net65));
 sg13g2_tiehi _1807__66 (.L_HI(net66));
 sg13g2_tiehi _1806__67 (.L_HI(net67));
 sg13g2_tiehi _1805__68 (.L_HI(net68));
 sg13g2_tiehi _1804__69 (.L_HI(net69));
 sg13g2_tiehi _1803__70 (.L_HI(net70));
 sg13g2_tiehi _1802__71 (.L_HI(net71));
 sg13g2_tiehi _1801__72 (.L_HI(net72));
 sg13g2_tiehi _1800__73 (.L_HI(net73));
 sg13g2_tiehi _1799__74 (.L_HI(net74));
 sg13g2_tiehi _1798__75 (.L_HI(net75));
 sg13g2_tiehi _1797__76 (.L_HI(net76));
 sg13g2_tiehi _1796__77 (.L_HI(net77));
 sg13g2_tiehi _1795__78 (.L_HI(net78));
 sg13g2_tiehi _1794__79 (.L_HI(net79));
 sg13g2_tiehi _1793__80 (.L_HI(net80));
 sg13g2_tiehi _1792__81 (.L_HI(net81));
 sg13g2_tiehi _1791__82 (.L_HI(net82));
 sg13g2_tiehi _1790__83 (.L_HI(net83));
 sg13g2_tiehi _1789__84 (.L_HI(net84));
 sg13g2_tiehi _1766__85 (.L_HI(net85));
 sg13g2_tiehi _1809__86 (.L_HI(net86));
 sg13g2_tiehi _1810__87 (.L_HI(net87));
 sg13g2_tiehi _1811__88 (.L_HI(net88));
 sg13g2_tiehi _1812__89 (.L_HI(net89));
 sg13g2_tiehi _1813__90 (.L_HI(net90));
 sg13g2_tiehi _1814__91 (.L_HI(net91));
 sg13g2_tiehi _1815__92 (.L_HI(net92));
 sg13g2_tiehi _1816__93 (.L_HI(net93));
 sg13g2_tiehi _1817__94 (.L_HI(net94));
 sg13g2_tiehi _1818__95 (.L_HI(net95));
 sg13g2_tiehi _1819__96 (.L_HI(net96));
 sg13g2_tiehi _1820__97 (.L_HI(net97));
 sg13g2_tiehi _1821__98 (.L_HI(net98));
 sg13g2_tiehi _1822__99 (.L_HI(net99));
 sg13g2_tiehi _1823__100 (.L_HI(net100));
 sg13g2_tiehi _1788__101 (.L_HI(net101));
 sg13g2_tiehi _1787__102 (.L_HI(net102));
 sg13g2_tiehi _1786__103 (.L_HI(net103));
 sg13g2_tiehi _1785__104 (.L_HI(net104));
 sg13g2_tiehi _1784__105 (.L_HI(net105));
 sg13g2_tiehi _1783__106 (.L_HI(net106));
 sg13g2_tiehi _1782__107 (.L_HI(net107));
 sg13g2_tiehi _1781__108 (.L_HI(net108));
 sg13g2_tiehi _1780__109 (.L_HI(net109));
 sg13g2_tiehi _1824__110 (.L_HI(net110));
 sg13g2_tiehi _1834__111 (.L_HI(net111));
 sg13g2_tiehi _1835__112 (.L_HI(net112));
 sg13g2_tiehi _1836__113 (.L_HI(net113));
 sg13g2_tiehi _1837__114 (.L_HI(net114));
 sg13g2_tiehi _1838__115 (.L_HI(net115));
 sg13g2_tiehi _1839__116 (.L_HI(net116));
 sg13g2_tiehi _1840__117 (.L_HI(net117));
 sg13g2_tiehi _1841__118 (.L_HI(net118));
 sg13g2_tiehi _1842__119 (.L_HI(net119));
 sg13g2_tiehi _1843__120 (.L_HI(net120));
 sg13g2_tiehi _1844__121 (.L_HI(net121));
 sg13g2_tiehi _1845__122 (.L_HI(net122));
 sg13g2_tiehi _1846__123 (.L_HI(net123));
 sg13g2_tiehi _1847__124 (.L_HI(net124));
 sg13g2_tiehi _1848__125 (.L_HI(net125));
 sg13g2_tiehi _1849__126 (.L_HI(net126));
 sg13g2_tiehi _1850__127 (.L_HI(net127));
 sg13g2_tiehi _1851__128 (.L_HI(net128));
 sg13g2_tiehi _1852__129 (.L_HI(net129));
 sg13g2_tiehi _1853__130 (.L_HI(net130));
 sg13g2_tiehi _1854__131 (.L_HI(net131));
 sg13g2_tiehi _1779__132 (.L_HI(net132));
 sg13g2_tiehi _1855__133 (.L_HI(net133));
 sg13g2_tiehi _1857__134 (.L_HI(net134));
 sg13g2_tiehi _1858__135 (.L_HI(net135));
 sg13g2_tiehi _1859__136 (.L_HI(net136));
 sg13g2_tiehi _1860__137 (.L_HI(net137));
 sg13g2_tiehi _1861__138 (.L_HI(net138));
 sg13g2_tiehi _1862__139 (.L_HI(net139));
 sg13g2_tiehi _1778__140 (.L_HI(net140));
 sg13g2_tiehi _1777__141 (.L_HI(net141));
 sg13g2_tiehi _1776__142 (.L_HI(net142));
 sg13g2_tiehi _1775__143 (.L_HI(net143));
 sg13g2_tiehi _1774__144 (.L_HI(net144));
 sg13g2_tiehi _1773__145 (.L_HI(net145));
 sg13g2_tiehi _1772__146 (.L_HI(net146));
 sg13g2_tiehi _1771__147 (.L_HI(net147));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_wokwi_414120248222232577_19 (.L_LO(net19));
 sg13g2_tielo tt_um_wokwi_414120248222232577_20 (.L_LO(net20));
 sg13g2_tielo tt_um_wokwi_414120248222232577_21 (.L_LO(net21));
 sg13g2_tielo tt_um_wokwi_414120248222232577_22 (.L_LO(net22));
 sg13g2_tielo tt_um_wokwi_414120248222232577_23 (.L_LO(net23));
 sg13g2_tielo tt_um_wokwi_414120248222232577_24 (.L_LO(net24));
 sg13g2_tielo tt_um_wokwi_414120248222232577_25 (.L_LO(net25));
 sg13g2_tielo tt_um_wokwi_414120248222232577_26 (.L_LO(net26));
 sg13g2_tielo tt_um_wokwi_414120248222232577_27 (.L_LO(net27));
 sg13g2_tielo tt_um_wokwi_414120248222232577_28 (.L_LO(net28));
 sg13g2_tielo tt_um_wokwi_414120248222232577_29 (.L_LO(net29));
 sg13g2_tielo tt_um_wokwi_414120248222232577_30 (.L_LO(net30));
 sg13g2_tielo tt_um_wokwi_414120248222232577_31 (.L_LO(net31));
 sg13g2_tielo tt_um_wokwi_414120248222232577_32 (.L_LO(net32));
 sg13g2_tielo tt_um_wokwi_414120248222232577_33 (.L_LO(net33));
 sg13g2_tiehi _1770__34 (.L_HI(net34));
 sg13g2_buf_2 fanout150 (.A(_0154_),
    .X(net150));
 sg13g2_buf_1 fanout151 (.A(_0154_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_0143_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_0117_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_0111_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_0110_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_0109_),
    .X(net156));
 sg13g2_buf_4 fanout157 (.X(net157),
    .A(\inst_sine_A.phase[6] ));
 sg13g2_buf_2 fanout158 (.A(\inst_sine_A.phase[6] ),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(\sine_Areg[6] ),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(\sine_Areg[6] ),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(net163),
    .X(net161));
 sg13g2_buf_1 fanout162 (.A(net163),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(\sine_Areg[5] ),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(\sine_Areg[4] ),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(\sine_Areg[4] ),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(\sine_Areg[3] ),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(\sine_Areg[3] ),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(\sine_Areg[2] ),
    .X(net168));
 sg13g2_buf_1 fanout169 (.A(\sine_Areg[2] ),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(\sine_Areg[1] ),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(net172),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(\sine_Breg[7] ),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(net174),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(\sine_Breg[4] ),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(net176),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(net177),
    .X(net176));
 sg13g2_buf_1 fanout177 (.A(\sine_Breg[3] ),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(net179),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(\sine_Breg[2] ),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(net182),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(net182),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(\sine_Breg[1] ),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(net184),
    .X(net183));
 sg13g2_buf_1 fanout184 (.A(net185),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(net186),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(\sine_Breg[0] ),
    .X(net186));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(net299));
 sg13g2_buf_2 fanout188 (.A(\inst_sine_B.phase[6] ),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(net190),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(\sine_Areg[7] ),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(\sine_Breg[6] ),
    .X(net191));
 sg13g2_buf_1 fanout192 (.A(\sine_Breg[6] ),
    .X(net192));
 sg13g2_buf_4 fanout193 (.X(net193),
    .A(_0105_));
 sg13g2_buf_2 fanout194 (.A(net195),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(net200),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(net197),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(net200),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(net200),
    .X(net198));
 sg13g2_buf_1 fanout199 (.A(net200),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(net1),
    .X(net200));
 sg13g2_buf_4 fanout201 (.X(net201),
    .A(net1));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[1]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[2]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[3]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[4]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[5]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[6]),
    .X(net16));
 sg13g2_buf_1 input17 (.A(uio_in[7]),
    .X(net17));
 sg13g2_tielo tt_um_wokwi_414120248222232577_18 (.L_LO(net18));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0771_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold2 (.A(\boxcar_storage[2][2] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0015_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0770_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0098_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold6 (.A(\boxcar_storage[3][0] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold7 (.A(\boxcar_storage[3][7] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold8 (.A(\boxcar_storage[3][3] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold9 (.A(\boxcar_storage[2][0] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold10 (.A(\boxcar_storage[1][0] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold11 (.A(\boxcar_storage[3][5] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold12 (.A(\boxcar_storage[3][4] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold13 (.A(\boxcar_storage[2][3] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold14 (.A(\boxcar_storage[2][6] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold15 (.A(\boxcar_storage[3][1] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold16 (.A(\boxcar_storage[1][4] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold17 (.A(\boxcar_storage[1][1] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold18 (.A(\boxcar_storage[1][7] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold19 (.A(\boxcar_storage[2][5] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold20 (.A(\boxcar_storage[1][3] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold21 (.A(\boxcar_storage[2][1] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold22 (.A(\boxcar_storage[3][6] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold23 (.A(\boxcar_storage[2][4] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold24 (.A(\boxcar_storage[2][7] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold25 (.A(\boxcar_storage[1][2] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold26 (.A(\boxcar_storage[3][2] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold27 (.A(\boxcar_storage[1][5] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold28 (.A(\boxcar_storage[1][6] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold29 (.A(\product[14] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0029_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold31 (.A(\product[11] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0026_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold33 (.A(\product[13] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0028_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold35 (.A(\product[12] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0027_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold37 (.A(\product[10] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0025_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold39 (.A(\product[8] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0023_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold41 (.A(\mixer_out[1] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold42 (.A(\mixer_out[2] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold43 (.A(\product[9] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0305_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0024_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold46 (.A(\mixer_out[0] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold47 (.A(\mixer_out[3] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold48 (.A(\boxcar_filter[0] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0640_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold50 (.A(\boxcar_filter[9] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0007_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold52 (.A(\inst_sine_A.phase[7] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0014_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0227_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0010_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold56 (.A(bypass_B),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0008_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold58 (.A(lowamp_B),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold59 (.A(\mixer_out[6] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold60 (.A(\inst_sine_B.phase[7] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold61 (.A(\boxcar_filter[7] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0005_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold63 (.A(\boxcar_storage[4][0] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0040_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold65 (.A(\boxcar_filter[4] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0002_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold67 (.A(\boxcar_filter[6] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0004_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold69 (.A(\inst_sine_B.phase[7] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold70 (.A(\mixer_out[4] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold71 (.A(\boxcar_filter[3] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0001_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold73 (.A(\phase_incr_A[5] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0761_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0096_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold76 (.A(\boxcar_filter[2] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold77 (.A(\mixer_out[5] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold78 (.A(\mixer_out[7] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold79 (.A(\boxcar_filter[5] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0003_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold81 (.A(\phase_incr_B[3] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0725_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0085_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold84 (.A(\phase_incr_B[5] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0734_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0087_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold87 (.A(\inst_sine_A.phase[5] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold88 (.A(\boxcar_filter[8] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0006_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold90 (.A(\phase_incr_B[0] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0715_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0082_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold93 (.A(\phase_incr_A[3] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0752_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0094_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold96 (.A(\phase_incr_A[0] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0742_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0091_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold99 (.A(\inst_sine_A.phase[4] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold100 (.A(\inst_sine_B.phase[6] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold101 (.A(\phase_incr_B[1] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0083_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0022_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold104 (.A(\phase_incr_A[1] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0744_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0745_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0092_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold108 (.A(\phase_incr_B[4] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0729_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold110 (.A(\inst_sine_B.phase[5] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold111 (.A(\phase_incr_A[2] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0747_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0749_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0093_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold115 (.A(\phase_incr_A[4] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold116 (.A(\phase_incr_B[2] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0720_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0084_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold119 (.A(\phase_incr_A[6] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0017_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0664_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0042_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0018_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0020_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0016_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0655_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0020_),
    .X(net326));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_4 FILLER_7_98 ();
 sg13g2_fill_1 FILLER_7_102 ();
 sg13g2_decap_8 FILLER_7_116 ();
 sg13g2_fill_2 FILLER_7_128 ();
 sg13g2_fill_1 FILLER_7_130 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_162 ();
 sg13g2_decap_8 FILLER_7_169 ();
 sg13g2_decap_4 FILLER_7_184 ();
 sg13g2_fill_2 FILLER_7_188 ();
 sg13g2_decap_4 FILLER_7_198 ();
 sg13g2_fill_2 FILLER_7_202 ();
 sg13g2_decap_4 FILLER_7_208 ();
 sg13g2_fill_2 FILLER_7_212 ();
 sg13g2_decap_4 FILLER_7_218 ();
 sg13g2_decap_4 FILLER_7_226 ();
 sg13g2_fill_2 FILLER_7_230 ();
 sg13g2_decap_8 FILLER_7_242 ();
 sg13g2_decap_8 FILLER_7_249 ();
 sg13g2_decap_8 FILLER_7_256 ();
 sg13g2_decap_8 FILLER_7_263 ();
 sg13g2_decap_8 FILLER_7_270 ();
 sg13g2_decap_8 FILLER_7_277 ();
 sg13g2_decap_8 FILLER_7_284 ();
 sg13g2_decap_8 FILLER_7_291 ();
 sg13g2_decap_8 FILLER_7_298 ();
 sg13g2_decap_8 FILLER_7_305 ();
 sg13g2_decap_8 FILLER_7_312 ();
 sg13g2_decap_8 FILLER_7_319 ();
 sg13g2_decap_8 FILLER_7_326 ();
 sg13g2_decap_8 FILLER_7_333 ();
 sg13g2_decap_8 FILLER_7_340 ();
 sg13g2_decap_8 FILLER_7_347 ();
 sg13g2_decap_8 FILLER_7_354 ();
 sg13g2_decap_8 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_368 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_4 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_fill_2 FILLER_8_98 ();
 sg13g2_fill_2 FILLER_8_116 ();
 sg13g2_fill_2 FILLER_8_126 ();
 sg13g2_fill_1 FILLER_8_165 ();
 sg13g2_fill_2 FILLER_8_195 ();
 sg13g2_fill_2 FILLER_8_217 ();
 sg13g2_fill_1 FILLER_8_219 ();
 sg13g2_decap_8 FILLER_8_253 ();
 sg13g2_decap_8 FILLER_8_260 ();
 sg13g2_decap_8 FILLER_8_267 ();
 sg13g2_decap_8 FILLER_8_274 ();
 sg13g2_decap_8 FILLER_8_281 ();
 sg13g2_decap_8 FILLER_8_288 ();
 sg13g2_decap_8 FILLER_8_295 ();
 sg13g2_decap_8 FILLER_8_302 ();
 sg13g2_decap_8 FILLER_8_309 ();
 sg13g2_decap_8 FILLER_8_316 ();
 sg13g2_decap_8 FILLER_8_323 ();
 sg13g2_decap_8 FILLER_8_330 ();
 sg13g2_decap_8 FILLER_8_337 ();
 sg13g2_decap_8 FILLER_8_344 ();
 sg13g2_decap_8 FILLER_8_351 ();
 sg13g2_decap_8 FILLER_8_358 ();
 sg13g2_decap_8 FILLER_8_365 ();
 sg13g2_decap_8 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_8_379 ();
 sg13g2_decap_8 FILLER_8_386 ();
 sg13g2_decap_8 FILLER_8_393 ();
 sg13g2_decap_8 FILLER_8_400 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_fill_2 FILLER_9_105 ();
 sg13g2_fill_1 FILLER_9_107 ();
 sg13g2_decap_8 FILLER_9_113 ();
 sg13g2_fill_2 FILLER_9_120 ();
 sg13g2_fill_1 FILLER_9_127 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_fill_2 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_162 ();
 sg13g2_fill_1 FILLER_9_173 ();
 sg13g2_decap_8 FILLER_9_177 ();
 sg13g2_fill_1 FILLER_9_189 ();
 sg13g2_decap_4 FILLER_9_194 ();
 sg13g2_decap_4 FILLER_9_207 ();
 sg13g2_fill_2 FILLER_9_211 ();
 sg13g2_decap_4 FILLER_9_219 ();
 sg13g2_fill_1 FILLER_9_228 ();
 sg13g2_fill_2 FILLER_9_237 ();
 sg13g2_fill_1 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_261 ();
 sg13g2_fill_2 FILLER_9_268 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_4 FILLER_10_91 ();
 sg13g2_decap_4 FILLER_10_113 ();
 sg13g2_decap_4 FILLER_10_143 ();
 sg13g2_fill_2 FILLER_10_147 ();
 sg13g2_decap_4 FILLER_10_161 ();
 sg13g2_fill_1 FILLER_10_198 ();
 sg13g2_decap_8 FILLER_10_220 ();
 sg13g2_fill_2 FILLER_10_231 ();
 sg13g2_fill_1 FILLER_10_233 ();
 sg13g2_fill_2 FILLER_10_253 ();
 sg13g2_decap_4 FILLER_10_259 ();
 sg13g2_fill_2 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_290 ();
 sg13g2_decap_8 FILLER_10_297 ();
 sg13g2_decap_8 FILLER_10_304 ();
 sg13g2_decap_8 FILLER_10_311 ();
 sg13g2_decap_8 FILLER_10_318 ();
 sg13g2_decap_8 FILLER_10_325 ();
 sg13g2_decap_8 FILLER_10_332 ();
 sg13g2_decap_8 FILLER_10_339 ();
 sg13g2_decap_8 FILLER_10_346 ();
 sg13g2_decap_8 FILLER_10_353 ();
 sg13g2_decap_8 FILLER_10_360 ();
 sg13g2_decap_8 FILLER_10_367 ();
 sg13g2_decap_8 FILLER_10_374 ();
 sg13g2_decap_8 FILLER_10_381 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_395 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_4 FILLER_11_89 ();
 sg13g2_fill_2 FILLER_11_93 ();
 sg13g2_decap_4 FILLER_11_113 ();
 sg13g2_fill_1 FILLER_11_140 ();
 sg13g2_decap_4 FILLER_11_167 ();
 sg13g2_fill_2 FILLER_11_171 ();
 sg13g2_decap_4 FILLER_11_178 ();
 sg13g2_decap_4 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_214 ();
 sg13g2_fill_2 FILLER_11_221 ();
 sg13g2_fill_1 FILLER_11_223 ();
 sg13g2_decap_4 FILLER_11_229 ();
 sg13g2_fill_2 FILLER_11_233 ();
 sg13g2_decap_8 FILLER_11_240 ();
 sg13g2_fill_1 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_281 ();
 sg13g2_fill_1 FILLER_11_288 ();
 sg13g2_fill_1 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_305 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_4 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_60 ();
 sg13g2_decap_8 FILLER_12_113 ();
 sg13g2_decap_4 FILLER_12_120 ();
 sg13g2_decap_8 FILLER_12_136 ();
 sg13g2_fill_1 FILLER_12_143 ();
 sg13g2_fill_2 FILLER_12_149 ();
 sg13g2_fill_1 FILLER_12_164 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_fill_2 FILLER_12_196 ();
 sg13g2_fill_1 FILLER_12_198 ();
 sg13g2_decap_4 FILLER_12_213 ();
 sg13g2_fill_1 FILLER_12_239 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_fill_2 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_299 ();
 sg13g2_decap_8 FILLER_12_306 ();
 sg13g2_decap_8 FILLER_12_313 ();
 sg13g2_decap_8 FILLER_12_320 ();
 sg13g2_decap_4 FILLER_12_337 ();
 sg13g2_fill_1 FILLER_12_341 ();
 sg13g2_fill_2 FILLER_12_346 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_decap_4 FILLER_12_359 ();
 sg13g2_fill_1 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_fill_2 FILLER_13_63 ();
 sg13g2_fill_1 FILLER_13_93 ();
 sg13g2_fill_2 FILLER_13_119 ();
 sg13g2_fill_1 FILLER_13_121 ();
 sg13g2_decap_4 FILLER_13_135 ();
 sg13g2_fill_1 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_4 FILLER_13_168 ();
 sg13g2_fill_2 FILLER_13_172 ();
 sg13g2_decap_8 FILLER_13_181 ();
 sg13g2_fill_2 FILLER_13_188 ();
 sg13g2_decap_8 FILLER_13_214 ();
 sg13g2_fill_2 FILLER_13_221 ();
 sg13g2_fill_1 FILLER_13_223 ();
 sg13g2_decap_8 FILLER_13_230 ();
 sg13g2_decap_8 FILLER_13_237 ();
 sg13g2_fill_2 FILLER_13_244 ();
 sg13g2_fill_1 FILLER_13_258 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_fill_2 FILLER_13_273 ();
 sg13g2_fill_1 FILLER_13_275 ();
 sg13g2_fill_2 FILLER_13_293 ();
 sg13g2_decap_4 FILLER_13_316 ();
 sg13g2_fill_1 FILLER_13_336 ();
 sg13g2_fill_2 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_370 ();
 sg13g2_fill_1 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_decap_8 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_fill_2 FILLER_14_56 ();
 sg13g2_fill_1 FILLER_14_58 ();
 sg13g2_fill_2 FILLER_14_85 ();
 sg13g2_fill_2 FILLER_14_96 ();
 sg13g2_fill_1 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_fill_2 FILLER_14_126 ();
 sg13g2_fill_1 FILLER_14_128 ();
 sg13g2_decap_4 FILLER_14_142 ();
 sg13g2_fill_1 FILLER_14_146 ();
 sg13g2_decap_4 FILLER_14_164 ();
 sg13g2_fill_2 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_183 ();
 sg13g2_decap_4 FILLER_14_190 ();
 sg13g2_decap_4 FILLER_14_210 ();
 sg13g2_fill_2 FILLER_14_214 ();
 sg13g2_fill_1 FILLER_14_241 ();
 sg13g2_decap_8 FILLER_14_264 ();
 sg13g2_fill_2 FILLER_14_271 ();
 sg13g2_decap_8 FILLER_14_278 ();
 sg13g2_decap_4 FILLER_14_285 ();
 sg13g2_decap_4 FILLER_14_309 ();
 sg13g2_fill_1 FILLER_14_313 ();
 sg13g2_decap_8 FILLER_14_332 ();
 sg13g2_decap_8 FILLER_14_339 ();
 sg13g2_fill_2 FILLER_14_346 ();
 sg13g2_decap_8 FILLER_14_400 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_4 FILLER_15_42 ();
 sg13g2_fill_1 FILLER_15_46 ();
 sg13g2_decap_4 FILLER_15_113 ();
 sg13g2_decap_8 FILLER_15_141 ();
 sg13g2_fill_2 FILLER_15_148 ();
 sg13g2_decap_8 FILLER_15_158 ();
 sg13g2_fill_1 FILLER_15_165 ();
 sg13g2_fill_2 FILLER_15_191 ();
 sg13g2_fill_2 FILLER_15_205 ();
 sg13g2_decap_8 FILLER_15_212 ();
 sg13g2_fill_2 FILLER_15_219 ();
 sg13g2_fill_1 FILLER_15_225 ();
 sg13g2_decap_8 FILLER_15_236 ();
 sg13g2_fill_2 FILLER_15_243 ();
 sg13g2_fill_1 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_258 ();
 sg13g2_fill_2 FILLER_15_265 ();
 sg13g2_decap_8 FILLER_15_284 ();
 sg13g2_decap_4 FILLER_15_291 ();
 sg13g2_fill_1 FILLER_15_295 ();
 sg13g2_decap_8 FILLER_15_306 ();
 sg13g2_fill_1 FILLER_15_313 ();
 sg13g2_fill_2 FILLER_15_336 ();
 sg13g2_fill_1 FILLER_15_338 ();
 sg13g2_decap_4 FILLER_15_354 ();
 sg13g2_fill_1 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_4 FILLER_15_377 ();
 sg13g2_fill_2 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_4 FILLER_16_49 ();
 sg13g2_fill_2 FILLER_16_88 ();
 sg13g2_fill_2 FILLER_16_99 ();
 sg13g2_fill_1 FILLER_16_101 ();
 sg13g2_decap_8 FILLER_16_110 ();
 sg13g2_fill_2 FILLER_16_128 ();
 sg13g2_fill_2 FILLER_16_146 ();
 sg13g2_decap_4 FILLER_16_165 ();
 sg13g2_fill_1 FILLER_16_169 ();
 sg13g2_fill_2 FILLER_16_191 ();
 sg13g2_fill_1 FILLER_16_193 ();
 sg13g2_decap_4 FILLER_16_265 ();
 sg13g2_decap_8 FILLER_16_281 ();
 sg13g2_fill_2 FILLER_16_309 ();
 sg13g2_decap_8 FILLER_16_316 ();
 sg13g2_fill_2 FILLER_16_323 ();
 sg13g2_fill_1 FILLER_16_325 ();
 sg13g2_fill_1 FILLER_16_330 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_fill_1 FILLER_16_361 ();
 sg13g2_decap_4 FILLER_16_373 ();
 sg13g2_decap_4 FILLER_16_389 ();
 sg13g2_fill_1 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_4 FILLER_17_49 ();
 sg13g2_fill_1 FILLER_17_117 ();
 sg13g2_decap_8 FILLER_17_141 ();
 sg13g2_fill_1 FILLER_17_148 ();
 sg13g2_decap_8 FILLER_17_164 ();
 sg13g2_fill_2 FILLER_17_198 ();
 sg13g2_fill_1 FILLER_17_200 ();
 sg13g2_decap_8 FILLER_17_214 ();
 sg13g2_fill_2 FILLER_17_221 ();
 sg13g2_fill_1 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_237 ();
 sg13g2_fill_2 FILLER_17_244 ();
 sg13g2_decap_8 FILLER_17_258 ();
 sg13g2_decap_4 FILLER_17_287 ();
 sg13g2_fill_2 FILLER_17_313 ();
 sg13g2_fill_1 FILLER_17_315 ();
 sg13g2_fill_1 FILLER_17_330 ();
 sg13g2_decap_8 FILLER_17_359 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_fill_2 FILLER_18_42 ();
 sg13g2_fill_1 FILLER_18_44 ();
 sg13g2_fill_2 FILLER_18_97 ();
 sg13g2_fill_1 FILLER_18_99 ();
 sg13g2_decap_8 FILLER_18_109 ();
 sg13g2_decap_8 FILLER_18_116 ();
 sg13g2_fill_2 FILLER_18_123 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_4 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_167 ();
 sg13g2_decap_8 FILLER_18_190 ();
 sg13g2_fill_1 FILLER_18_197 ();
 sg13g2_fill_2 FILLER_18_221 ();
 sg13g2_decap_8 FILLER_18_227 ();
 sg13g2_decap_4 FILLER_18_234 ();
 sg13g2_fill_2 FILLER_18_238 ();
 sg13g2_decap_4 FILLER_18_264 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_fill_2 FILLER_18_287 ();
 sg13g2_fill_1 FILLER_18_289 ();
 sg13g2_fill_2 FILLER_18_305 ();
 sg13g2_fill_1 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_320 ();
 sg13g2_fill_1 FILLER_18_343 ();
 sg13g2_fill_2 FILLER_18_380 ();
 sg13g2_fill_1 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_4 FILLER_19_49 ();
 sg13g2_fill_2 FILLER_19_66 ();
 sg13g2_fill_1 FILLER_19_68 ();
 sg13g2_fill_2 FILLER_19_87 ();
 sg13g2_fill_2 FILLER_19_115 ();
 sg13g2_decap_4 FILLER_19_147 ();
 sg13g2_decap_4 FILLER_19_185 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_194 ();
 sg13g2_fill_2 FILLER_19_201 ();
 sg13g2_fill_1 FILLER_19_203 ();
 sg13g2_decap_4 FILLER_19_230 ();
 sg13g2_fill_1 FILLER_19_234 ();
 sg13g2_fill_2 FILLER_19_266 ();
 sg13g2_fill_1 FILLER_19_268 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_fill_2 FILLER_19_324 ();
 sg13g2_decap_4 FILLER_19_337 ();
 sg13g2_fill_2 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_fill_2 FILLER_19_371 ();
 sg13g2_fill_1 FILLER_19_373 ();
 sg13g2_decap_4 FILLER_19_390 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_11 ();
 sg13g2_decap_8 FILLER_20_16 ();
 sg13g2_fill_2 FILLER_20_23 ();
 sg13g2_fill_1 FILLER_20_25 ();
 sg13g2_fill_2 FILLER_20_31 ();
 sg13g2_fill_2 FILLER_20_42 ();
 sg13g2_fill_1 FILLER_20_44 ();
 sg13g2_fill_1 FILLER_20_93 ();
 sg13g2_fill_2 FILLER_20_120 ();
 sg13g2_fill_1 FILLER_20_122 ();
 sg13g2_fill_1 FILLER_20_132 ();
 sg13g2_fill_2 FILLER_20_164 ();
 sg13g2_decap_8 FILLER_20_205 ();
 sg13g2_fill_2 FILLER_20_212 ();
 sg13g2_fill_1 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_219 ();
 sg13g2_decap_4 FILLER_20_226 ();
 sg13g2_fill_2 FILLER_20_234 ();
 sg13g2_fill_2 FILLER_20_253 ();
 sg13g2_decap_4 FILLER_20_276 ();
 sg13g2_fill_2 FILLER_20_285 ();
 sg13g2_fill_1 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_298 ();
 sg13g2_fill_2 FILLER_20_305 ();
 sg13g2_decap_4 FILLER_20_316 ();
 sg13g2_fill_1 FILLER_20_320 ();
 sg13g2_decap_8 FILLER_20_339 ();
 sg13g2_fill_2 FILLER_20_346 ();
 sg13g2_decap_8 FILLER_20_352 ();
 sg13g2_decap_4 FILLER_20_359 ();
 sg13g2_fill_2 FILLER_20_363 ();
 sg13g2_fill_2 FILLER_20_380 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_12 ();
 sg13g2_fill_2 FILLER_21_80 ();
 sg13g2_fill_2 FILLER_21_108 ();
 sg13g2_fill_2 FILLER_21_145 ();
 sg13g2_decap_8 FILLER_21_195 ();
 sg13g2_fill_2 FILLER_21_202 ();
 sg13g2_fill_1 FILLER_21_204 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_247 ();
 sg13g2_decap_4 FILLER_21_254 ();
 sg13g2_fill_1 FILLER_21_258 ();
 sg13g2_decap_8 FILLER_21_272 ();
 sg13g2_decap_4 FILLER_21_279 ();
 sg13g2_fill_1 FILLER_21_283 ();
 sg13g2_fill_2 FILLER_21_289 ();
 sg13g2_fill_1 FILLER_21_291 ();
 sg13g2_decap_8 FILLER_21_296 ();
 sg13g2_fill_1 FILLER_21_303 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_fill_2 FILLER_21_315 ();
 sg13g2_fill_1 FILLER_21_317 ();
 sg13g2_decap_4 FILLER_21_334 ();
 sg13g2_fill_2 FILLER_21_338 ();
 sg13g2_fill_1 FILLER_21_360 ();
 sg13g2_fill_2 FILLER_21_385 ();
 sg13g2_fill_2 FILLER_22_26 ();
 sg13g2_fill_1 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_64 ();
 sg13g2_fill_2 FILLER_22_74 ();
 sg13g2_fill_2 FILLER_22_89 ();
 sg13g2_fill_1 FILLER_22_109 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_fill_2 FILLER_22_199 ();
 sg13g2_fill_2 FILLER_22_253 ();
 sg13g2_decap_4 FILLER_22_259 ();
 sg13g2_fill_2 FILLER_22_341 ();
 sg13g2_fill_1 FILLER_22_343 ();
 sg13g2_fill_2 FILLER_22_363 ();
 sg13g2_fill_1 FILLER_22_365 ();
 sg13g2_fill_2 FILLER_22_379 ();
 sg13g2_fill_2 FILLER_22_385 ();
 sg13g2_fill_1 FILLER_22_387 ();
 sg13g2_fill_2 FILLER_22_392 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_fill_1 FILLER_23_26 ();
 sg13g2_fill_2 FILLER_23_36 ();
 sg13g2_fill_1 FILLER_23_38 ();
 sg13g2_fill_2 FILLER_23_57 ();
 sg13g2_fill_1 FILLER_23_59 ();
 sg13g2_fill_2 FILLER_23_108 ();
 sg13g2_fill_1 FILLER_23_110 ();
 sg13g2_fill_1 FILLER_23_125 ();
 sg13g2_fill_2 FILLER_23_140 ();
 sg13g2_fill_1 FILLER_23_164 ();
 sg13g2_fill_2 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_221 ();
 sg13g2_decap_8 FILLER_23_228 ();
 sg13g2_fill_2 FILLER_23_270 ();
 sg13g2_decap_4 FILLER_23_281 ();
 sg13g2_fill_1 FILLER_23_285 ();
 sg13g2_decap_8 FILLER_23_295 ();
 sg13g2_decap_4 FILLER_23_302 ();
 sg13g2_decap_8 FILLER_23_311 ();
 sg13g2_decap_4 FILLER_23_318 ();
 sg13g2_fill_1 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_328 ();
 sg13g2_fill_1 FILLER_23_374 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_71 ();
 sg13g2_fill_1 FILLER_24_94 ();
 sg13g2_fill_2 FILLER_24_108 ();
 sg13g2_fill_2 FILLER_24_125 ();
 sg13g2_fill_1 FILLER_24_127 ();
 sg13g2_fill_1 FILLER_24_180 ();
 sg13g2_fill_2 FILLER_24_190 ();
 sg13g2_fill_2 FILLER_24_201 ();
 sg13g2_fill_1 FILLER_24_203 ();
 sg13g2_fill_1 FILLER_24_209 ();
 sg13g2_fill_2 FILLER_24_248 ();
 sg13g2_decap_4 FILLER_24_260 ();
 sg13g2_fill_1 FILLER_24_341 ();
 sg13g2_fill_2 FILLER_24_382 ();
 sg13g2_fill_2 FILLER_24_388 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_53 ();
 sg13g2_fill_1 FILLER_25_104 ();
 sg13g2_fill_1 FILLER_25_115 ();
 sg13g2_fill_2 FILLER_25_159 ();
 sg13g2_fill_2 FILLER_25_218 ();
 sg13g2_fill_1 FILLER_25_220 ();
 sg13g2_fill_2 FILLER_25_240 ();
 sg13g2_fill_2 FILLER_25_269 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_decap_8 FILLER_25_331 ();
 sg13g2_fill_2 FILLER_25_338 ();
 sg13g2_fill_2 FILLER_25_360 ();
 sg13g2_fill_1 FILLER_25_362 ();
 sg13g2_fill_2 FILLER_25_373 ();
 sg13g2_fill_2 FILLER_25_387 ();
 sg13g2_fill_1 FILLER_25_389 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_2 FILLER_26_83 ();
 sg13g2_fill_1 FILLER_26_134 ();
 sg13g2_fill_1 FILLER_26_139 ();
 sg13g2_decap_8 FILLER_26_211 ();
 sg13g2_fill_1 FILLER_26_218 ();
 sg13g2_fill_1 FILLER_26_297 ();
 sg13g2_fill_2 FILLER_26_302 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_fill_1 FILLER_26_367 ();
 sg13g2_fill_1 FILLER_26_378 ();
 sg13g2_fill_1 FILLER_26_383 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_15 ();
 sg13g2_fill_1 FILLER_27_17 ();
 sg13g2_fill_2 FILLER_27_53 ();
 sg13g2_fill_1 FILLER_27_55 ();
 sg13g2_fill_2 FILLER_27_65 ();
 sg13g2_fill_2 FILLER_27_80 ();
 sg13g2_fill_1 FILLER_27_82 ();
 sg13g2_fill_2 FILLER_27_121 ();
 sg13g2_fill_2 FILLER_27_149 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_fill_2 FILLER_27_187 ();
 sg13g2_fill_1 FILLER_27_189 ();
 sg13g2_fill_1 FILLER_27_216 ();
 sg13g2_fill_1 FILLER_27_225 ();
 sg13g2_decap_4 FILLER_27_230 ();
 sg13g2_fill_2 FILLER_27_234 ();
 sg13g2_fill_2 FILLER_27_307 ();
 sg13g2_fill_1 FILLER_27_309 ();
 sg13g2_fill_2 FILLER_27_336 ();
 sg13g2_fill_2 FILLER_27_388 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_29 ();
 sg13g2_fill_1 FILLER_28_31 ();
 sg13g2_fill_2 FILLER_28_45 ();
 sg13g2_fill_1 FILLER_28_47 ();
 sg13g2_fill_1 FILLER_28_52 ();
 sg13g2_fill_1 FILLER_28_58 ();
 sg13g2_fill_2 FILLER_28_79 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_fill_2 FILLER_28_140 ();
 sg13g2_fill_2 FILLER_28_186 ();
 sg13g2_fill_1 FILLER_28_188 ();
 sg13g2_fill_2 FILLER_28_198 ();
 sg13g2_fill_1 FILLER_28_200 ();
 sg13g2_decap_4 FILLER_28_205 ();
 sg13g2_fill_2 FILLER_28_209 ();
 sg13g2_decap_8 FILLER_28_241 ();
 sg13g2_fill_2 FILLER_28_248 ();
 sg13g2_fill_1 FILLER_28_281 ();
 sg13g2_decap_4 FILLER_28_287 ();
 sg13g2_fill_1 FILLER_28_296 ();
 sg13g2_fill_1 FILLER_28_302 ();
 sg13g2_decap_8 FILLER_28_307 ();
 sg13g2_fill_2 FILLER_28_314 ();
 sg13g2_fill_1 FILLER_28_324 ();
 sg13g2_fill_2 FILLER_28_389 ();
 sg13g2_fill_1 FILLER_28_391 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_32 ();
 sg13g2_fill_1 FILLER_29_73 ();
 sg13g2_decap_8 FILLER_29_167 ();
 sg13g2_fill_1 FILLER_29_209 ();
 sg13g2_decap_8 FILLER_29_214 ();
 sg13g2_decap_8 FILLER_29_221 ();
 sg13g2_decap_8 FILLER_29_228 ();
 sg13g2_decap_8 FILLER_29_235 ();
 sg13g2_decap_4 FILLER_29_242 ();
 sg13g2_fill_2 FILLER_29_246 ();
 sg13g2_fill_1 FILLER_29_253 ();
 sg13g2_fill_2 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_267 ();
 sg13g2_fill_2 FILLER_29_288 ();
 sg13g2_fill_1 FILLER_29_318 ();
 sg13g2_fill_1 FILLER_29_397 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_decap_4 FILLER_30_33 ();
 sg13g2_fill_2 FILLER_30_37 ();
 sg13g2_fill_1 FILLER_30_47 ();
 sg13g2_fill_2 FILLER_30_52 ();
 sg13g2_fill_2 FILLER_30_105 ();
 sg13g2_fill_1 FILLER_30_129 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_fill_1 FILLER_30_177 ();
 sg13g2_fill_2 FILLER_30_187 ();
 sg13g2_fill_1 FILLER_30_189 ();
 sg13g2_decap_4 FILLER_30_195 ();
 sg13g2_decap_4 FILLER_30_225 ();
 sg13g2_fill_2 FILLER_30_251 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_decap_4 FILLER_30_280 ();
 sg13g2_fill_1 FILLER_30_284 ();
 sg13g2_fill_2 FILLER_30_304 ();
 sg13g2_fill_1 FILLER_30_306 ();
 sg13g2_fill_1 FILLER_30_312 ();
 sg13g2_fill_2 FILLER_30_326 ();
 sg13g2_fill_2 FILLER_30_344 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_73 ();
 sg13g2_fill_1 FILLER_31_145 ();
 sg13g2_fill_2 FILLER_31_155 ();
 sg13g2_fill_1 FILLER_31_213 ();
 sg13g2_decap_4 FILLER_31_268 ();
 sg13g2_fill_1 FILLER_31_279 ();
 sg13g2_fill_2 FILLER_31_298 ();
 sg13g2_fill_2 FILLER_31_305 ();
 sg13g2_fill_2 FILLER_31_327 ();
 sg13g2_fill_1 FILLER_31_355 ();
 sg13g2_fill_1 FILLER_31_365 ();
 sg13g2_fill_1 FILLER_31_382 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_11 ();
 sg13g2_fill_1 FILLER_32_22 ();
 sg13g2_fill_1 FILLER_32_32 ();
 sg13g2_fill_2 FILLER_32_52 ();
 sg13g2_fill_2 FILLER_32_84 ();
 sg13g2_fill_1 FILLER_32_94 ();
 sg13g2_fill_2 FILLER_32_144 ();
 sg13g2_fill_2 FILLER_32_150 ();
 sg13g2_fill_2 FILLER_32_170 ();
 sg13g2_decap_8 FILLER_32_234 ();
 sg13g2_decap_4 FILLER_32_241 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_fill_2 FILLER_32_273 ();
 sg13g2_fill_1 FILLER_32_275 ();
 sg13g2_fill_2 FILLER_32_281 ();
 sg13g2_fill_2 FILLER_32_300 ();
 sg13g2_fill_1 FILLER_32_302 ();
 sg13g2_fill_2 FILLER_32_325 ();
 sg13g2_fill_1 FILLER_32_337 ();
 sg13g2_fill_2 FILLER_32_359 ();
 sg13g2_fill_1 FILLER_32_392 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_12 ();
 sg13g2_fill_2 FILLER_33_16 ();
 sg13g2_fill_1 FILLER_33_44 ();
 sg13g2_fill_2 FILLER_33_77 ();
 sg13g2_fill_2 FILLER_33_97 ();
 sg13g2_fill_2 FILLER_33_120 ();
 sg13g2_fill_1 FILLER_33_188 ();
 sg13g2_fill_2 FILLER_33_279 ();
 sg13g2_fill_1 FILLER_33_281 ();
 sg13g2_fill_1 FILLER_33_326 ();
 sg13g2_fill_1 FILLER_33_353 ();
 sg13g2_fill_2 FILLER_33_373 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_fill_2 FILLER_34_26 ();
 sg13g2_fill_2 FILLER_34_141 ();
 sg13g2_fill_1 FILLER_34_143 ();
 sg13g2_decap_4 FILLER_34_156 ();
 sg13g2_fill_1 FILLER_34_160 ();
 sg13g2_fill_2 FILLER_34_165 ();
 sg13g2_fill_1 FILLER_34_167 ();
 sg13g2_decap_4 FILLER_34_172 ();
 sg13g2_fill_1 FILLER_34_176 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_decap_4 FILLER_34_227 ();
 sg13g2_fill_1 FILLER_34_297 ();
 sg13g2_fill_2 FILLER_34_322 ();
 sg13g2_fill_1 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_355 ();
 sg13g2_fill_2 FILLER_34_371 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_68 ();
 sg13g2_fill_1 FILLER_35_70 ();
 sg13g2_fill_1 FILLER_35_126 ();
 sg13g2_fill_2 FILLER_35_196 ();
 sg13g2_fill_2 FILLER_35_235 ();
 sg13g2_fill_2 FILLER_35_242 ();
 sg13g2_fill_1 FILLER_35_244 ();
 sg13g2_fill_1 FILLER_35_302 ();
 sg13g2_fill_1 FILLER_35_340 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_fill_2 FILLER_36_52 ();
 sg13g2_fill_1 FILLER_36_54 ();
 sg13g2_fill_2 FILLER_36_81 ();
 sg13g2_fill_1 FILLER_36_83 ();
 sg13g2_fill_1 FILLER_36_133 ();
 sg13g2_fill_1 FILLER_36_159 ();
 sg13g2_fill_1 FILLER_36_177 ();
 sg13g2_fill_2 FILLER_36_196 ();
 sg13g2_fill_2 FILLER_36_264 ();
 sg13g2_fill_1 FILLER_36_266 ();
 sg13g2_fill_2 FILLER_36_326 ();
 sg13g2_fill_1 FILLER_36_363 ();
 sg13g2_fill_1 FILLER_36_377 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_4 FILLER_37_21 ();
 sg13g2_fill_2 FILLER_37_30 ();
 sg13g2_fill_2 FILLER_37_36 ();
 sg13g2_fill_2 FILLER_37_130 ();
 sg13g2_fill_2 FILLER_37_158 ();
 sg13g2_fill_1 FILLER_37_212 ();
 sg13g2_fill_1 FILLER_37_266 ();
 sg13g2_fill_1 FILLER_37_276 ();
 sg13g2_fill_2 FILLER_37_285 ();
 sg13g2_fill_1 FILLER_37_306 ();
 sg13g2_fill_1 FILLER_37_316 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_fill_1 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_105 ();
 sg13g2_fill_2 FILLER_38_137 ();
 sg13g2_fill_1 FILLER_38_139 ();
 sg13g2_fill_2 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_150 ();
 sg13g2_fill_2 FILLER_38_164 ();
 sg13g2_fill_1 FILLER_38_166 ();
 sg13g2_fill_1 FILLER_38_175 ();
 sg13g2_fill_2 FILLER_38_188 ();
 sg13g2_fill_1 FILLER_38_190 ();
 sg13g2_fill_2 FILLER_38_200 ();
 sg13g2_fill_2 FILLER_38_250 ();
 sg13g2_fill_2 FILLER_38_282 ();
 sg13g2_fill_1 FILLER_38_284 ();
 sg13g2_fill_2 FILLER_38_290 ();
 sg13g2_fill_1 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_342 ();
 assign uio_oe[0] = net18;
 assign uio_oe[1] = net19;
 assign uio_oe[2] = net20;
 assign uio_oe[3] = net21;
 assign uio_oe[4] = net22;
 assign uio_oe[5] = net23;
 assign uio_oe[6] = net24;
 assign uio_oe[7] = net25;
 assign uio_out[0] = net26;
 assign uio_out[1] = net27;
 assign uio_out[2] = net28;
 assign uio_out[3] = net29;
 assign uio_out[4] = net30;
 assign uio_out[5] = net31;
 assign uio_out[6] = net32;
 assign uio_out[7] = net33;
endmodule

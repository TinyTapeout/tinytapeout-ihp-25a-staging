module tt_um_top (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \LFSR[0] ;
 wire \LFSR[1] ;
 wire \LFSR[2] ;
 wire \LFSR[3] ;
 wire \LFSR[4] ;
 wire \LFSR[5] ;
 wire \VAL[0] ;
 wire \VAL[10] ;
 wire \VAL[11] ;
 wire \VAL[12] ;
 wire \VAL[13] ;
 wire \VAL[14] ;
 wire \VAL[15] ;
 wire \VAL[16] ;
 wire \VAL[17] ;
 wire \VAL[18] ;
 wire \VAL[19] ;
 wire \VAL[1] ;
 wire \VAL[20] ;
 wire \VAL[21] ;
 wire \VAL[22] ;
 wire \VAL[23] ;
 wire \VAL[2] ;
 wire \VAL[3] ;
 wire \VAL[4] ;
 wire \VAL[5] ;
 wire \VAL[6] ;
 wire \VAL[7] ;
 wire \VAL[8] ;
 wire \VAL[9] ;
 wire \Voice1.accumulator[0] ;
 wire \Voice1.accumulator[10] ;
 wire \Voice1.accumulator[11] ;
 wire \Voice1.accumulator[12] ;
 wire \Voice1.accumulator[13] ;
 wire \Voice1.accumulator[14] ;
 wire \Voice1.accumulator[15] ;
 wire \Voice1.accumulator[16] ;
 wire \Voice1.accumulator[17] ;
 wire \Voice1.accumulator[18] ;
 wire \Voice1.accumulator[19] ;
 wire \Voice1.accumulator[1] ;
 wire \Voice1.accumulator[20] ;
 wire \Voice1.accumulator[21] ;
 wire \Voice1.accumulator[22] ;
 wire \Voice1.accumulator[23] ;
 wire \Voice1.accumulator[2] ;
 wire \Voice1.accumulator[3] ;
 wire \Voice1.accumulator[4] ;
 wire \Voice1.accumulator[5] ;
 wire \Voice1.accumulator[6] ;
 wire \Voice1.accumulator[7] ;
 wire \Voice1.accumulator[8] ;
 wire \Voice1.accumulator[9] ;
 wire \Voice1.en ;
 wire \Voice1.pulse ;
 wire \Voice1.pulsewidth[0] ;
 wire \Voice1.pulsewidth[10] ;
 wire \Voice1.pulsewidth[1] ;
 wire \Voice1.pulsewidth[2] ;
 wire \Voice1.pulsewidth[3] ;
 wire \Voice1.pulsewidth[4] ;
 wire \Voice1.pulsewidth[5] ;
 wire \Voice1.pulsewidth[6] ;
 wire \Voice1.pulsewidth[7] ;
 wire \Voice1.pulsewidth[8] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \ctr_audio[0] ;
 wire \ctr_audio[19] ;
 wire \ctr_audio[1] ;
 wire \ctr_audio[20] ;
 wire \ctr_audio[21] ;
 wire \ctr_audio[22] ;
 wire \ctr_audio[2] ;
 wire \ctr_audio[3] ;
 wire \ctr_audio[4] ;
 wire \ctr_audio[5] ;
 wire \ctr_audio[6] ;
 wire \ctr_audio[7] ;
 wire \ctr_audio[8] ;
 wire \ctr_audio[9] ;
 wire \ctr_clkdiv25[0] ;
 wire \ctr_clkdiv25[1] ;
 wire \ctr_clkdiv25[2] ;
 wire \ctr_clkdiv25[3] ;
 wire \ctr_clkdiv25[4] ;
 wire \ctr_clkdiv25[5] ;
 wire \ctr_clkdiv25[6] ;
 wire \ctr_clkdiv25[7] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_0_clk;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire \xq[0] ;
 wire \xq[10] ;
 wire \xq[11] ;
 wire \xq[1] ;
 wire \xq[2] ;
 wire \xq[3] ;
 wire \xq[4] ;
 wire \xq[5] ;
 wire \xq[6] ;
 wire \xq[7] ;
 wire \xq[8] ;
 wire \xq[9] ;
 wire \xqo[0] ;
 wire \xqo[10] ;
 wire \xqo[11] ;
 wire \xqo[1] ;
 wire \xqo[2] ;
 wire \xqo[3] ;
 wire \xqo[4] ;
 wire \xqo[5] ;
 wire \xqo[6] ;
 wire \xqo[7] ;
 wire \xqo[8] ;
 wire \xqo[9] ;
 wire \yq[0] ;
 wire \yq[10] ;
 wire \yq[11] ;
 wire \yq[12] ;
 wire \yq[1] ;
 wire \yq[2] ;
 wire \yq[3] ;
 wire \yq[4] ;
 wire \yq[5] ;
 wire \yq[6] ;
 wire \yq[7] ;
 wire \yq[8] ;
 wire \yq[9] ;
 wire \yqo[0] ;
 wire \yqo[10] ;
 wire \yqo[11] ;
 wire \yqo[12] ;
 wire \yqo[1] ;
 wire \yqo[2] ;
 wire \yqo[3] ;
 wire \yqo[4] ;
 wire \yqo[5] ;
 wire \yqo[6] ;
 wire \yqo[7] ;
 wire \yqo[8] ;
 wire \yqo[9] ;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net1;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;

 sg13g2_inv_2 _1262_ (.Y(_0412_),
    .A(net172));
 sg13g2_inv_1 _1263_ (.Y(_0413_),
    .A(net377));
 sg13g2_inv_1 _1264_ (.Y(_0414_),
    .A(net437));
 sg13g2_inv_1 _1265_ (.Y(_0415_),
    .A(\Voice1.pulsewidth[8] ));
 sg13g2_inv_1 _1266_ (.Y(_0416_),
    .A(net188));
 sg13g2_inv_1 _1267_ (.Y(_0417_),
    .A(\Voice1.pulsewidth[5] ));
 sg13g2_inv_1 _1268_ (.Y(_0418_),
    .A(net369));
 sg13g2_inv_1 _1269_ (.Y(_0419_),
    .A(net466));
 sg13g2_inv_1 _1270_ (.Y(_0420_),
    .A(net258));
 sg13g2_inv_1 _1271_ (.Y(_0421_),
    .A(net286));
 sg13g2_inv_1 _1272_ (.Y(_0422_),
    .A(net451));
 sg13g2_inv_1 _1273_ (.Y(_0423_),
    .A(net299));
 sg13g2_inv_1 _1274_ (.Y(_0424_),
    .A(\yqo[11] ));
 sg13g2_inv_1 _1275_ (.Y(_0425_),
    .A(\yqo[9] ));
 sg13g2_inv_1 _1276_ (.Y(_0426_),
    .A(\yqo[7] ));
 sg13g2_inv_1 _1277_ (.Y(_0427_),
    .A(\ctr_clkdiv25[0] ));
 sg13g2_inv_1 _1278_ (.Y(_0428_),
    .A(net310));
 sg13g2_inv_1 _1279_ (.Y(_0429_),
    .A(\Voice1.accumulator[13] ));
 sg13g2_inv_1 _1280_ (.Y(_0430_),
    .A(\Voice1.accumulator[15] ));
 sg13g2_inv_1 _1281_ (.Y(_0431_),
    .A(\Voice1.accumulator[14] ));
 sg13g2_inv_1 _1282_ (.Y(_0432_),
    .A(net427));
 sg13g2_inv_1 _1283_ (.Y(_0433_),
    .A(net251));
 sg13g2_inv_1 _1284_ (.Y(_0434_),
    .A(net439));
 sg13g2_inv_1 _1285_ (.Y(_0435_),
    .A(net316));
 sg13g2_inv_1 _1286_ (.Y(_0436_),
    .A(net264));
 sg13g2_inv_1 _1287_ (.Y(_0437_),
    .A(\Voice1.accumulator[21] ));
 sg13g2_inv_1 _1288_ (.Y(_0438_),
    .A(net201));
 sg13g2_inv_1 _1289_ (.Y(_0439_),
    .A(net195));
 sg13g2_inv_1 _1290_ (.Y(_0440_),
    .A(\ctr_clkdiv25[3] ));
 sg13g2_inv_1 _1291_ (.Y(_0441_),
    .A(\ctr_clkdiv25[4] ));
 sg13g2_inv_1 _1292_ (.Y(_0442_),
    .A(\VAL[5] ));
 sg13g2_inv_1 _1293_ (.Y(_0443_),
    .A(\LFSR[5] ));
 sg13g2_inv_2 _1294_ (.Y(_0444_),
    .A(net394));
 sg13g2_inv_2 _1295_ (.Y(_0445_),
    .A(net340));
 sg13g2_inv_1 _1296_ (.Y(_0446_),
    .A(\VAL[3] ));
 sg13g2_inv_1 _1297_ (.Y(_0447_),
    .A(net429));
 sg13g2_inv_1 _1298_ (.Y(_0448_),
    .A(\LFSR[1] ));
 sg13g2_inv_1 _1299_ (.Y(_0449_),
    .A(\LFSR[0] ));
 sg13g2_inv_1 _1300_ (.Y(_0450_),
    .A(net361));
 sg13g2_inv_1 _1301_ (.Y(_0451_),
    .A(\VAL[13] ));
 sg13g2_inv_1 _1302_ (.Y(_0452_),
    .A(\VAL[11] ));
 sg13g2_inv_1 _1303_ (.Y(_0453_),
    .A(\VAL[9] ));
 sg13g2_inv_1 _1304_ (.Y(_0454_),
    .A(net249));
 sg13g2_inv_1 _1305_ (.Y(_0455_),
    .A(_0008_));
 sg13g2_inv_1 _1306_ (.Y(_0456_),
    .A(_0010_));
 sg13g2_inv_1 _1307_ (.Y(_0457_),
    .A(net331));
 sg13g2_inv_1 _1308_ (.Y(_0458_),
    .A(net302));
 sg13g2_inv_1 _1309_ (.Y(_0459_),
    .A(net410));
 sg13g2_inv_1 _1310_ (.Y(_0460_),
    .A(\counter[3] ));
 sg13g2_inv_1 _1311_ (.Y(_0461_),
    .A(\counter[8] ));
 sg13g2_inv_1 _1312_ (.Y(_0462_),
    .A(net358));
 sg13g2_inv_1 _1313_ (.Y(_0463_),
    .A(net454));
 sg13g2_inv_1 _1314_ (.Y(_0464_),
    .A(net372));
 sg13g2_nand4_1 _1315_ (.B(net178),
    .C(net179),
    .A(net176),
    .Y(_0465_),
    .D(net175));
 sg13g2_nand3b_1 _1316_ (.B(net183),
    .C(net389),
    .Y(_0466_),
    .A_N(net356));
 sg13g2_nor4_1 _1317_ (.A(net181),
    .B(\hvsync_gen.vpos[9] ),
    .C(_0465_),
    .D(net390),
    .Y(_0001_));
 sg13g2_nor3_1 _1318_ (.A(net193),
    .B(net195),
    .C(net194),
    .Y(_0467_));
 sg13g2_nor2b_1 _1319_ (.A(_0467_),
    .B_N(\hvsync_gen.hpos[9] ),
    .Y(_0468_));
 sg13g2_a22oi_1 _1320_ (.Y(_0469_),
    .B1(_0468_),
    .B2(net192),
    .A2(\hvsync_gen.hpos[9] ),
    .A1(net191));
 sg13g2_nand4_1 _1321_ (.B(net193),
    .C(net195),
    .A(\hvsync_gen.hpos[7] ),
    .Y(_0470_),
    .D(net194));
 sg13g2_nor2b_1 _1322_ (.A(net191),
    .B_N(net189),
    .Y(_0471_));
 sg13g2_a21oi_1 _1323_ (.A1(_0470_),
    .A2(_0471_),
    .Y(_0472_),
    .B1(net279));
 sg13g2_nor2_1 _1324_ (.A(_0469_),
    .B(net280),
    .Y(_0000_));
 sg13g2_a22oi_1 _1325_ (.Y(_0473_),
    .B1(_0444_),
    .B2(\VAL[4] ),
    .A2(_0443_),
    .A1(\VAL[5] ));
 sg13g2_nand2b_1 _1326_ (.Y(_0474_),
    .B(\LFSR[1] ),
    .A_N(\VAL[1] ));
 sg13g2_a22oi_1 _1327_ (.Y(_0475_),
    .B1(\VAL[0] ),
    .B2(_0449_),
    .A2(\VAL[1] ),
    .A1(_0448_));
 sg13g2_o21ai_1 _1328_ (.B1(_0474_),
    .Y(_0476_),
    .A1(net169),
    .A2(\VAL[2] ));
 sg13g2_or2_1 _1329_ (.X(_0477_),
    .B(_0476_),
    .A(_0475_));
 sg13g2_a22oi_1 _1330_ (.Y(_0478_),
    .B1(net169),
    .B2(\VAL[2] ),
    .A2(\VAL[3] ),
    .A1(_0445_));
 sg13g2_a22oi_1 _1331_ (.Y(_0479_),
    .B1(_0477_),
    .B2(_0478_),
    .A2(_0446_),
    .A1(\LFSR[3] ));
 sg13g2_o21ai_1 _1332_ (.B1(_0479_),
    .Y(_0480_),
    .A1(_0444_),
    .A2(\VAL[4] ));
 sg13g2_a22oi_1 _1333_ (.Y(_0481_),
    .B1(_0473_),
    .B2(_0480_),
    .A2(\LFSR[5] ),
    .A1(_0442_));
 sg13g2_and2_1 _1334_ (.A(\VAL[6] ),
    .B(_0481_),
    .X(_0482_));
 sg13g2_nor2_1 _1335_ (.A(net192),
    .B(net190),
    .Y(_0483_));
 sg13g2_nor2b_1 _1336_ (.A(\hvsync_gen.vpos[9] ),
    .B_N(_0465_),
    .Y(_0484_));
 sg13g2_o21ai_1 _1337_ (.B1(_0484_),
    .Y(_0485_),
    .A1(_0006_),
    .A2(_0483_));
 sg13g2_inv_1 _1338_ (.Y(_0486_),
    .A(_0485_));
 sg13g2_o21ai_1 _1339_ (.B1(_0486_),
    .Y(_0487_),
    .A1(\VAL[6] ),
    .A2(_0481_));
 sg13g2_nor2_1 _1340_ (.A(_0482_),
    .B(_0487_),
    .Y(uo_out[4]));
 sg13g2_xnor2_1 _1341_ (.Y(_0488_),
    .A(\VAL[7] ),
    .B(_0482_));
 sg13g2_nor2_1 _1342_ (.A(_0485_),
    .B(_0488_),
    .Y(uo_out[0]));
 sg13g2_a22oi_1 _1343_ (.Y(_0489_),
    .B1(\VAL[12] ),
    .B2(_0444_),
    .A2(\VAL[13] ),
    .A1(_0443_));
 sg13g2_a22oi_1 _1344_ (.Y(_0490_),
    .B1(\VAL[8] ),
    .B2(_0449_),
    .A2(\VAL[9] ),
    .A1(_0448_));
 sg13g2_a21oi_1 _1345_ (.A1(\LFSR[1] ),
    .A2(_0453_),
    .Y(_0491_),
    .B1(_0490_));
 sg13g2_o21ai_1 _1346_ (.B1(_0491_),
    .Y(_0492_),
    .A1(net169),
    .A2(\VAL[10] ));
 sg13g2_a22oi_1 _1347_ (.Y(_0493_),
    .B1(\VAL[10] ),
    .B2(net169),
    .A2(\VAL[11] ),
    .A1(_0445_));
 sg13g2_a22oi_1 _1348_ (.Y(_0494_),
    .B1(_0492_),
    .B2(_0493_),
    .A2(_0452_),
    .A1(\LFSR[3] ));
 sg13g2_o21ai_1 _1349_ (.B1(_0494_),
    .Y(_0495_),
    .A1(_0444_),
    .A2(\VAL[12] ));
 sg13g2_a22oi_1 _1350_ (.Y(_0496_),
    .B1(_0489_),
    .B2(_0495_),
    .A2(_0451_),
    .A1(\LFSR[5] ));
 sg13g2_xnor2_1 _1351_ (.Y(_0497_),
    .A(_0454_),
    .B(_0496_));
 sg13g2_nor2_1 _1352_ (.A(_0485_),
    .B(_0497_),
    .Y(uo_out[5]));
 sg13g2_and2_1 _1353_ (.A(\VAL[14] ),
    .B(_0496_),
    .X(_0498_));
 sg13g2_o21ai_1 _1354_ (.B1(_0486_),
    .Y(_0499_),
    .A1(\VAL[15] ),
    .A2(_0498_));
 sg13g2_a21oi_1 _1355_ (.A1(\VAL[15] ),
    .A2(_0498_),
    .Y(uo_out[1]),
    .B1(_0499_));
 sg13g2_nand2b_1 _1356_ (.Y(_0500_),
    .B(\VAL[17] ),
    .A_N(\LFSR[1] ));
 sg13g2_nand2b_1 _1357_ (.Y(_0501_),
    .B(\VAL[16] ),
    .A_N(\LFSR[0] ));
 sg13g2_nand2b_1 _1358_ (.Y(_0502_),
    .B(\LFSR[1] ),
    .A_N(\VAL[17] ));
 sg13g2_o21ai_1 _1359_ (.B1(_0502_),
    .Y(_0503_),
    .A1(net169),
    .A2(\VAL[18] ));
 sg13g2_a21oi_1 _1360_ (.A1(_0500_),
    .A2(_0501_),
    .Y(_0504_),
    .B1(_0503_));
 sg13g2_a221oi_1 _1361_ (.B2(net169),
    .C1(_0504_),
    .B1(\VAL[18] ),
    .A1(_0445_),
    .Y(_0505_),
    .A2(\VAL[19] ));
 sg13g2_nor2_1 _1362_ (.A(_0443_),
    .B(\VAL[21] ),
    .Y(_0506_));
 sg13g2_nand2b_1 _1363_ (.Y(_0507_),
    .B(\LFSR[4] ),
    .A_N(\VAL[20] ));
 sg13g2_o21ai_1 _1364_ (.B1(_0507_),
    .Y(_0508_),
    .A1(_0445_),
    .A2(\VAL[19] ));
 sg13g2_or3_1 _1365_ (.A(_0505_),
    .B(_0506_),
    .C(_0508_),
    .X(_0509_));
 sg13g2_a22oi_1 _1366_ (.Y(_0510_),
    .B1(\VAL[20] ),
    .B2(_0444_),
    .A2(\VAL[21] ),
    .A1(_0443_));
 sg13g2_o21ai_1 _1367_ (.B1(_0509_),
    .Y(_0511_),
    .A1(_0506_),
    .A2(_0510_));
 sg13g2_and2_1 _1368_ (.A(\VAL[22] ),
    .B(_0511_),
    .X(_0512_));
 sg13g2_o21ai_1 _1369_ (.B1(_0486_),
    .Y(_0513_),
    .A1(\VAL[22] ),
    .A2(_0511_));
 sg13g2_nor2_1 _1370_ (.A(_0512_),
    .B(_0513_),
    .Y(uo_out[6]));
 sg13g2_o21ai_1 _1371_ (.B1(_0486_),
    .Y(_0514_),
    .A1(\VAL[23] ),
    .A2(_0512_));
 sg13g2_a21oi_1 _1372_ (.A1(\VAL[23] ),
    .A2(_0512_),
    .Y(uo_out[2]),
    .B1(_0514_));
 sg13g2_and2_1 _1373_ (.A(\hvsync_gen.hpos[0] ),
    .B(net268),
    .X(_0515_));
 sg13g2_nand3_1 _1374_ (.B(\hvsync_gen.hpos[3] ),
    .C(_0515_),
    .A(net313),
    .Y(_0516_));
 sg13g2_inv_1 _1375_ (.Y(_0517_),
    .A(_0516_));
 sg13g2_nor4_1 _1376_ (.A(net192),
    .B(net193),
    .C(_0439_),
    .D(net194),
    .Y(_0518_));
 sg13g2_nand4_1 _1377_ (.B(net189),
    .C(_0517_),
    .A(net190),
    .Y(_0519_),
    .D(_0518_));
 sg13g2_and2_2 _1378_ (.A(net207),
    .B(_0519_),
    .X(_0520_));
 sg13g2_nand2_1 _1379_ (.Y(_0521_),
    .A(net207),
    .B(_0519_));
 sg13g2_and2_1 _1380_ (.A(net235),
    .B(_0520_),
    .X(_0021_));
 sg13g2_nor2_1 _1381_ (.A(\hvsync_gen.hpos[0] ),
    .B(net268),
    .Y(_0522_));
 sg13g2_nor3_1 _1382_ (.A(net197),
    .B(_0515_),
    .C(net269),
    .Y(_0022_));
 sg13g2_o21ai_1 _1383_ (.B1(net203),
    .Y(_0523_),
    .A1(net313),
    .A2(_0515_));
 sg13g2_a21oi_1 _1384_ (.A1(net313),
    .A2(_0515_),
    .Y(_0023_),
    .B1(_0523_));
 sg13g2_nor2b_1 _1385_ (.A(net338),
    .B_N(_0515_),
    .Y(_0524_));
 sg13g2_xnor2_1 _1386_ (.Y(_0525_),
    .A(net405),
    .B(_0524_));
 sg13g2_nor2_1 _1387_ (.A(net159),
    .B(_0525_),
    .Y(_0024_));
 sg13g2_xor2_1 _1388_ (.B(_0516_),
    .A(net195),
    .X(_0526_));
 sg13g2_nor2_1 _1389_ (.A(net159),
    .B(net476),
    .Y(_0025_));
 sg13g2_nor2_1 _1390_ (.A(net294),
    .B(_0516_),
    .Y(_0527_));
 sg13g2_xnor2_1 _1391_ (.Y(_0528_),
    .A(net194),
    .B(net295));
 sg13g2_nor2_1 _1392_ (.A(net159),
    .B(net296),
    .Y(_0026_));
 sg13g2_nand3_1 _1393_ (.B(net194),
    .C(_0517_),
    .A(net195),
    .Y(_0529_));
 sg13g2_xor2_1 _1394_ (.B(_0529_),
    .A(net193),
    .X(_0530_));
 sg13g2_nor2_1 _1395_ (.A(net159),
    .B(_0530_),
    .Y(_0027_));
 sg13g2_nor2_1 _1396_ (.A(net408),
    .B(_0529_),
    .Y(_0531_));
 sg13g2_xnor2_1 _1397_ (.Y(_0532_),
    .A(\hvsync_gen.hpos[7] ),
    .B(_0531_));
 sg13g2_nor2_1 _1398_ (.A(net159),
    .B(net409),
    .Y(_0028_));
 sg13g2_nor2_1 _1399_ (.A(_0470_),
    .B(_0516_),
    .Y(_0533_));
 sg13g2_nor2_1 _1400_ (.A(net191),
    .B(_0533_),
    .Y(_0534_));
 sg13g2_nand3_1 _1401_ (.B(net193),
    .C(net190),
    .A(\hvsync_gen.hpos[7] ),
    .Y(_0535_));
 sg13g2_nor2_1 _1402_ (.A(_0529_),
    .B(_0535_),
    .Y(_0536_));
 sg13g2_nor3_1 _1403_ (.A(net159),
    .B(net461),
    .C(_0536_),
    .Y(_0029_));
 sg13g2_o21ai_1 _1404_ (.B1(_0520_),
    .Y(_0537_),
    .A1(net189),
    .A2(_0536_));
 sg13g2_a21oi_1 _1405_ (.A1(net189),
    .A2(_0536_),
    .Y(_0030_),
    .B1(_0537_));
 sg13g2_and2_1 _1406_ (.A(net206),
    .B(_0019_),
    .X(_0031_));
 sg13g2_o21ai_1 _1407_ (.B1(net205),
    .Y(_0538_),
    .A1(\counter[0] ),
    .A2(\counter[1] ));
 sg13g2_a21oi_1 _1408_ (.A1(\counter[0] ),
    .A2(\counter[1] ),
    .Y(_0032_),
    .B1(_0538_));
 sg13g2_a21oi_1 _1409_ (.A1(\counter[0] ),
    .A2(\counter[1] ),
    .Y(_0539_),
    .B1(\counter[2] ));
 sg13g2_nand3_1 _1410_ (.B(\counter[1] ),
    .C(\counter[2] ),
    .A(\counter[0] ),
    .Y(_0540_));
 sg13g2_nand2_1 _1411_ (.Y(_0541_),
    .A(net205),
    .B(_0540_));
 sg13g2_nor2_1 _1412_ (.A(_0539_),
    .B(_0541_),
    .Y(_0033_));
 sg13g2_and2_1 _1413_ (.A(_0460_),
    .B(_0540_),
    .X(_0542_));
 sg13g2_nor2_1 _1414_ (.A(_0460_),
    .B(_0540_),
    .Y(_0543_));
 sg13g2_nor3_1 _1415_ (.A(net200),
    .B(_0542_),
    .C(_0543_),
    .Y(_0034_));
 sg13g2_and2_2 _1416_ (.A(\counter[4] ),
    .B(_0543_),
    .X(_0544_));
 sg13g2_o21ai_1 _1417_ (.B1(net206),
    .Y(_0545_),
    .A1(\counter[4] ),
    .A2(_0543_));
 sg13g2_nor2_1 _1418_ (.A(_0544_),
    .B(_0545_),
    .Y(_0035_));
 sg13g2_xnor2_1 _1419_ (.Y(_0546_),
    .A(net163),
    .B(_0544_));
 sg13g2_nor2_1 _1420_ (.A(net200),
    .B(_0546_),
    .Y(_0036_));
 sg13g2_a21oi_1 _1421_ (.A1(net163),
    .A2(_0544_),
    .Y(_0547_),
    .B1(\counter[6] ));
 sg13g2_nand3_1 _1422_ (.B(\counter[6] ),
    .C(_0544_),
    .A(net163),
    .Y(_0548_));
 sg13g2_nand2_1 _1423_ (.Y(_0549_),
    .A(net202),
    .B(_0548_));
 sg13g2_nor2_1 _1424_ (.A(_0547_),
    .B(_0549_),
    .Y(_0037_));
 sg13g2_nand2b_1 _1425_ (.Y(_0550_),
    .B(_0548_),
    .A_N(\counter[7] ));
 sg13g2_nand4_1 _1426_ (.B(\counter[6] ),
    .C(\counter[7] ),
    .A(net163),
    .Y(_0551_),
    .D(_0544_));
 sg13g2_and3_1 _1427_ (.X(_0038_),
    .A(net202),
    .B(_0550_),
    .C(_0551_));
 sg13g2_o21ai_1 _1428_ (.B1(net202),
    .Y(_0552_),
    .A1(_0461_),
    .A2(_0551_));
 sg13g2_a21oi_1 _1429_ (.A1(_0461_),
    .A2(_0551_),
    .Y(_0039_),
    .B1(_0552_));
 sg13g2_nand2b_1 _1430_ (.Y(_0553_),
    .B(\yq[5] ),
    .A_N(\xq[4] ));
 sg13g2_xor2_1 _1431_ (.B(\xq[4] ),
    .A(\yq[5] ),
    .X(_0554_));
 sg13g2_nand2b_1 _1432_ (.Y(_0555_),
    .B(\xq[10] ),
    .A_N(\yq[11] ));
 sg13g2_nand2b_1 _1433_ (.Y(_0556_),
    .B(\yq[8] ),
    .A_N(\xq[7] ));
 sg13g2_nor2b_1 _1434_ (.A(\yq[6] ),
    .B_N(\xq[5] ),
    .Y(_0557_));
 sg13g2_xnor2_1 _1435_ (.Y(_0558_),
    .A(\yq[6] ),
    .B(\xq[5] ));
 sg13g2_a21oi_2 _1436_ (.B1(_0557_),
    .Y(_0559_),
    .A2(_0558_),
    .A1(_0553_));
 sg13g2_nor2b_1 _1437_ (.A(\yq[7] ),
    .B_N(\xq[6] ),
    .Y(_0560_));
 sg13g2_xnor2_1 _1438_ (.Y(_0561_),
    .A(\yq[7] ),
    .B(\xq[6] ));
 sg13g2_nor2b_1 _1439_ (.A(_0559_),
    .B_N(_0561_),
    .Y(_0562_));
 sg13g2_nor2b_1 _1440_ (.A(\yq[8] ),
    .B_N(\xq[7] ),
    .Y(_0563_));
 sg13g2_a21oi_1 _1441_ (.A1(_0556_),
    .A2(_0560_),
    .Y(_0564_),
    .B1(_0563_));
 sg13g2_xnor2_1 _1442_ (.Y(_0565_),
    .A(\yq[8] ),
    .B(\xq[7] ));
 sg13g2_nand2_1 _1443_ (.Y(_0566_),
    .A(_0561_),
    .B(_0565_));
 sg13g2_o21ai_1 _1444_ (.B1(_0564_),
    .Y(_0567_),
    .A1(_0559_),
    .A2(_0566_));
 sg13g2_nor2b_1 _1445_ (.A(\yq[10] ),
    .B_N(\xq[9] ),
    .Y(_0568_));
 sg13g2_nand2b_1 _1446_ (.Y(_0569_),
    .B(\yq[10] ),
    .A_N(\xq[9] ));
 sg13g2_nand2b_1 _1447_ (.Y(_0570_),
    .B(_0569_),
    .A_N(_0568_));
 sg13g2_nor2b_1 _1448_ (.A(\yq[9] ),
    .B_N(\xq[8] ),
    .Y(_0571_));
 sg13g2_nand2b_1 _1449_ (.Y(_0572_),
    .B(\yq[9] ),
    .A_N(\xq[8] ));
 sg13g2_nand2b_1 _1450_ (.Y(_0573_),
    .B(_0572_),
    .A_N(_0571_));
 sg13g2_nor2_1 _1451_ (.A(_0570_),
    .B(_0573_),
    .Y(_0574_));
 sg13g2_a221oi_1 _1452_ (.B2(_0567_),
    .C1(_0568_),
    .B1(_0574_),
    .A1(_0569_),
    .Y(_0575_),
    .A2(_0571_));
 sg13g2_nor2b_1 _1453_ (.A(\xq[10] ),
    .B_N(\yq[11] ),
    .Y(_0576_));
 sg13g2_xnor2_1 _1454_ (.Y(_0577_),
    .A(\yq[11] ),
    .B(\xq[10] ));
 sg13g2_o21ai_1 _1455_ (.B1(_0555_),
    .Y(_0578_),
    .A1(_0575_),
    .A2(_0576_));
 sg13g2_xnor2_1 _1456_ (.Y(_0579_),
    .A(\yq[12] ),
    .B(\xq[11] ));
 sg13g2_xnor2_1 _1457_ (.Y(_0580_),
    .A(_0578_),
    .B(_0579_));
 sg13g2_xnor2_1 _1458_ (.Y(_0581_),
    .A(_0554_),
    .B(_0580_));
 sg13g2_nor2_1 _1459_ (.A(net183),
    .B(_0581_),
    .Y(_0582_));
 sg13g2_xor2_1 _1460_ (.B(_0581_),
    .A(net183),
    .X(_0583_));
 sg13g2_nor2b_1 _1461_ (.A(_0583_),
    .B_N(net338),
    .Y(_0584_));
 sg13g2_nor2b_1 _1462_ (.A(net338),
    .B_N(_0583_),
    .Y(_0585_));
 sg13g2_a21oi_1 _1463_ (.A1(net192),
    .A2(net193),
    .Y(_0586_),
    .B1(net190));
 sg13g2_and2_1 _1464_ (.A(net204),
    .B(_0535_),
    .X(_0587_));
 sg13g2_nor2_1 _1465_ (.A(net189),
    .B(_0586_),
    .Y(_0588_));
 sg13g2_nand2_2 _1466_ (.Y(_0589_),
    .A(_0587_),
    .B(_0588_));
 sg13g2_nor3_1 _1467_ (.A(_0584_),
    .B(_0585_),
    .C(_0589_),
    .Y(_0040_));
 sg13g2_xnor2_1 _1468_ (.Y(_0590_),
    .A(_0553_),
    .B(_0558_));
 sg13g2_xnor2_1 _1469_ (.Y(_0591_),
    .A(_0580_),
    .B(_0590_));
 sg13g2_xnor2_1 _1470_ (.Y(_0592_),
    .A(net181),
    .B(_0591_));
 sg13g2_xnor2_1 _1471_ (.Y(_0593_),
    .A(net405),
    .B(_0592_));
 sg13g2_a21oi_1 _1472_ (.A1(net183),
    .A2(_0581_),
    .Y(_0594_),
    .B1(net313));
 sg13g2_nor2_1 _1473_ (.A(_0582_),
    .B(_0594_),
    .Y(_0595_));
 sg13g2_inv_1 _1474_ (.Y(_0596_),
    .A(_0595_));
 sg13g2_nand2b_1 _1475_ (.Y(_0597_),
    .B(_0595_),
    .A_N(_0593_));
 sg13g2_nand2b_1 _1476_ (.Y(_0598_),
    .B(_0597_),
    .A_N(_0589_));
 sg13g2_a21oi_1 _1477_ (.A1(_0593_),
    .A2(_0596_),
    .Y(_0041_),
    .B1(_0598_));
 sg13g2_nor2_1 _1478_ (.A(_0014_),
    .B(_0591_),
    .Y(_0599_));
 sg13g2_a21oi_1 _1479_ (.A1(\hvsync_gen.hpos[3] ),
    .A2(_0592_),
    .Y(_0600_),
    .B1(_0599_));
 sg13g2_xnor2_1 _1480_ (.Y(_0601_),
    .A(_0559_),
    .B(_0561_));
 sg13g2_xnor2_1 _1481_ (.Y(_0602_),
    .A(_0580_),
    .B(_0601_));
 sg13g2_nor2_1 _1482_ (.A(net179),
    .B(_0602_),
    .Y(_0603_));
 sg13g2_xnor2_1 _1483_ (.Y(_0604_),
    .A(net179),
    .B(_0602_));
 sg13g2_nor2b_1 _1484_ (.A(_0600_),
    .B_N(_0604_),
    .Y(_0605_));
 sg13g2_xnor2_1 _1485_ (.Y(_0606_),
    .A(_0600_),
    .B(_0604_));
 sg13g2_xnor2_1 _1486_ (.Y(_0607_),
    .A(net475),
    .B(_0606_));
 sg13g2_and2_1 _1487_ (.A(_0597_),
    .B(_0607_),
    .X(_0608_));
 sg13g2_nor2_1 _1488_ (.A(_0597_),
    .B(_0607_),
    .Y(_0609_));
 sg13g2_nor3_1 _1489_ (.A(_0589_),
    .B(_0608_),
    .C(_0609_),
    .Y(_0042_));
 sg13g2_nor2_1 _1490_ (.A(_0560_),
    .B(_0562_),
    .Y(_0610_));
 sg13g2_xnor2_1 _1491_ (.Y(_0611_),
    .A(_0565_),
    .B(_0610_));
 sg13g2_xnor2_1 _1492_ (.Y(_0612_),
    .A(_0580_),
    .B(_0611_));
 sg13g2_xor2_1 _1493_ (.B(_0612_),
    .A(_0015_),
    .X(_0613_));
 sg13g2_nor2b_1 _1494_ (.A(_0603_),
    .B_N(_0613_),
    .Y(_0614_));
 sg13g2_xnor2_1 _1495_ (.Y(_0615_),
    .A(_0603_),
    .B(_0613_));
 sg13g2_xnor2_1 _1496_ (.Y(_0616_),
    .A(\hvsync_gen.hpos[5] ),
    .B(_0615_));
 sg13g2_a21oi_1 _1497_ (.A1(net195),
    .A2(_0606_),
    .Y(_0617_),
    .B1(_0605_));
 sg13g2_nor2_1 _1498_ (.A(_0616_),
    .B(_0617_),
    .Y(_0618_));
 sg13g2_nand2_1 _1499_ (.Y(_0619_),
    .A(_0616_),
    .B(_0617_));
 sg13g2_nand2b_1 _1500_ (.Y(_0620_),
    .B(_0619_),
    .A_N(_0618_));
 sg13g2_nor2b_1 _1501_ (.A(_0609_),
    .B_N(_0620_),
    .Y(_0621_));
 sg13g2_nor3_1 _1502_ (.A(_0597_),
    .B(_0607_),
    .C(_0620_),
    .Y(_0622_));
 sg13g2_nor3_1 _1503_ (.A(_0589_),
    .B(_0621_),
    .C(_0622_),
    .Y(_0043_));
 sg13g2_a21oi_2 _1504_ (.B1(_0618_),
    .Y(_0623_),
    .A2(_0619_),
    .A1(_0609_));
 sg13g2_nor2_1 _1505_ (.A(net178),
    .B(_0612_),
    .Y(_0624_));
 sg13g2_xnor2_1 _1506_ (.Y(_0625_),
    .A(_0567_),
    .B(_0573_));
 sg13g2_xnor2_1 _1507_ (.Y(_0626_),
    .A(_0580_),
    .B(_0625_));
 sg13g2_nand2_1 _1508_ (.Y(_0627_),
    .A(net176),
    .B(_0626_));
 sg13g2_xor2_1 _1509_ (.B(_0626_),
    .A(net176),
    .X(_0628_));
 sg13g2_xnor2_1 _1510_ (.Y(_0629_),
    .A(_0003_),
    .B(_0628_));
 sg13g2_nand2b_1 _1511_ (.Y(_0630_),
    .B(_0629_),
    .A_N(_0624_));
 sg13g2_xnor2_1 _1512_ (.Y(_0631_),
    .A(_0624_),
    .B(_0629_));
 sg13g2_a21o_1 _1513_ (.A2(_0615_),
    .A1(net194),
    .B1(_0614_),
    .X(_0632_));
 sg13g2_and2_1 _1514_ (.A(_0631_),
    .B(_0632_),
    .X(_0633_));
 sg13g2_nand2_1 _1515_ (.Y(_0634_),
    .A(_0631_),
    .B(_0632_));
 sg13g2_xor2_1 _1516_ (.B(_0632_),
    .A(_0631_),
    .X(_0635_));
 sg13g2_nand2b_1 _1517_ (.Y(_0636_),
    .B(_0635_),
    .A_N(_0623_));
 sg13g2_xor2_1 _1518_ (.B(_0635_),
    .A(_0623_),
    .X(_0637_));
 sg13g2_nor2_1 _1519_ (.A(_0589_),
    .B(_0637_),
    .Y(_0044_));
 sg13g2_a21o_1 _1520_ (.A2(_0572_),
    .A1(_0567_),
    .B1(_0571_),
    .X(_0638_));
 sg13g2_xnor2_1 _1521_ (.Y(_0639_),
    .A(_0570_),
    .B(_0638_));
 sg13g2_xnor2_1 _1522_ (.Y(_0640_),
    .A(_0580_),
    .B(_0639_));
 sg13g2_nor2_1 _1523_ (.A(net175),
    .B(_0640_),
    .Y(_0641_));
 sg13g2_xnor2_1 _1524_ (.Y(_0642_),
    .A(net175),
    .B(_0640_));
 sg13g2_o21ai_1 _1525_ (.B1(\hvsync_gen.hpos[6] ),
    .Y(_0643_),
    .A1(net176),
    .A2(_0626_));
 sg13g2_nand2_1 _1526_ (.Y(_0644_),
    .A(_0627_),
    .B(_0643_));
 sg13g2_and2_1 _1527_ (.A(_0642_),
    .B(_0644_),
    .X(_0645_));
 sg13g2_xor2_1 _1528_ (.B(_0644_),
    .A(_0642_),
    .X(_0646_));
 sg13g2_xnor2_1 _1529_ (.Y(_0647_),
    .A(net192),
    .B(_0646_));
 sg13g2_nor2_1 _1530_ (.A(_0630_),
    .B(_0647_),
    .Y(_0648_));
 sg13g2_nand2_1 _1531_ (.Y(_0649_),
    .A(_0630_),
    .B(_0647_));
 sg13g2_nand2b_1 _1532_ (.Y(_0650_),
    .B(_0649_),
    .A_N(_0648_));
 sg13g2_and3_1 _1533_ (.X(_0651_),
    .A(_0634_),
    .B(_0636_),
    .C(_0650_));
 sg13g2_a21oi_1 _1534_ (.A1(_0634_),
    .A2(_0636_),
    .Y(_0652_),
    .B1(_0650_));
 sg13g2_nor3_1 _1535_ (.A(_0589_),
    .B(_0651_),
    .C(_0652_),
    .Y(_0045_));
 sg13g2_nand3b_1 _1536_ (.B(_0649_),
    .C(_0635_),
    .Y(_0653_),
    .A_N(_0648_));
 sg13g2_a21oi_1 _1537_ (.A1(_0633_),
    .A2(_0649_),
    .Y(_0654_),
    .B1(_0648_));
 sg13g2_o21ai_1 _1538_ (.B1(_0654_),
    .Y(_0655_),
    .A1(_0623_),
    .A2(_0653_));
 sg13g2_xnor2_1 _1539_ (.Y(_0656_),
    .A(_0575_),
    .B(_0577_));
 sg13g2_xnor2_1 _1540_ (.Y(_0657_),
    .A(_0580_),
    .B(_0656_));
 sg13g2_nor2_1 _1541_ (.A(\hvsync_gen.vpos[9] ),
    .B(_0657_),
    .Y(_0658_));
 sg13g2_xnor2_1 _1542_ (.Y(_0659_),
    .A(\hvsync_gen.vpos[9] ),
    .B(_0657_));
 sg13g2_nor2b_1 _1543_ (.A(_0641_),
    .B_N(_0659_),
    .Y(_0660_));
 sg13g2_xnor2_1 _1544_ (.Y(_0661_),
    .A(_0641_),
    .B(_0659_));
 sg13g2_xnor2_1 _1545_ (.Y(_0662_),
    .A(net190),
    .B(_0661_));
 sg13g2_a21o_1 _1546_ (.A2(_0646_),
    .A1(net192),
    .B1(_0645_),
    .X(_0663_));
 sg13g2_nand2b_1 _1547_ (.Y(_0664_),
    .B(_0663_),
    .A_N(_0662_));
 sg13g2_xor2_1 _1548_ (.B(_0663_),
    .A(_0662_),
    .X(_0665_));
 sg13g2_nand2b_1 _1549_ (.Y(_0666_),
    .B(_0665_),
    .A_N(_0655_));
 sg13g2_nand2b_1 _1550_ (.Y(_0667_),
    .B(_0655_),
    .A_N(_0665_));
 sg13g2_and4_1 _1551_ (.A(_0587_),
    .B(_0588_),
    .C(_0666_),
    .D(_0667_),
    .X(_0046_));
 sg13g2_a21oi_1 _1552_ (.A1(net191),
    .A2(_0661_),
    .Y(_0668_),
    .B1(_0660_));
 sg13g2_xnor2_1 _1553_ (.Y(_0669_),
    .A(net189),
    .B(_0658_));
 sg13g2_xnor2_1 _1554_ (.Y(_0670_),
    .A(_0668_),
    .B(_0669_));
 sg13g2_and3_1 _1555_ (.X(_0671_),
    .A(_0664_),
    .B(_0667_),
    .C(_0670_));
 sg13g2_a21oi_1 _1556_ (.A1(_0664_),
    .A2(_0667_),
    .Y(_0672_),
    .B1(_0670_));
 sg13g2_nor3_1 _1557_ (.A(_0589_),
    .B(_0671_),
    .C(_0672_),
    .Y(_0047_));
 sg13g2_nand2_1 _1558_ (.Y(_0673_),
    .A(net182),
    .B(net386));
 sg13g2_o21ai_1 _1559_ (.B1(net208),
    .Y(_0674_),
    .A1(net182),
    .A2(net386));
 sg13g2_nor2b_1 _1560_ (.A(net387),
    .B_N(_0673_),
    .Y(_0048_));
 sg13g2_xnor2_1 _1561_ (.Y(_0675_),
    .A(net180),
    .B(net456));
 sg13g2_and2_1 _1562_ (.A(_0673_),
    .B(_0675_),
    .X(_0676_));
 sg13g2_nor2_1 _1563_ (.A(_0673_),
    .B(_0675_),
    .Y(_0677_));
 sg13g2_nor3_1 _1564_ (.A(net200),
    .B(net457),
    .C(_0677_),
    .Y(_0049_));
 sg13g2_xnor2_1 _1565_ (.Y(_0678_),
    .A(net178),
    .B(net480));
 sg13g2_a21oi_1 _1566_ (.A1(net180),
    .A2(net456),
    .Y(_0679_),
    .B1(_0677_));
 sg13g2_and2_1 _1567_ (.A(_0678_),
    .B(_0679_),
    .X(_0680_));
 sg13g2_nor2_1 _1568_ (.A(_0678_),
    .B(_0679_),
    .Y(_0681_));
 sg13g2_nor3_1 _1569_ (.A(net200),
    .B(_0680_),
    .C(_0681_),
    .Y(_0050_));
 sg13g2_xnor2_1 _1570_ (.Y(_0682_),
    .A(net177),
    .B(net440));
 sg13g2_a21oi_1 _1571_ (.A1(\hvsync_gen.vpos[6] ),
    .A2(\VAL[2] ),
    .Y(_0683_),
    .B1(_0681_));
 sg13g2_or2_1 _1572_ (.X(_0684_),
    .B(_0683_),
    .A(_0682_));
 sg13g2_inv_1 _1573_ (.Y(_0685_),
    .A(_0684_));
 sg13g2_nand2_1 _1574_ (.Y(_0686_),
    .A(net208),
    .B(_0684_));
 sg13g2_a21oi_1 _1575_ (.A1(net441),
    .A2(_0683_),
    .Y(_0051_),
    .B1(_0686_));
 sg13g2_xnor2_1 _1576_ (.Y(_0687_),
    .A(net473),
    .B(net474));
 sg13g2_a21oi_1 _1577_ (.A1(net177),
    .A2(net440),
    .Y(_0688_),
    .B1(_0685_));
 sg13g2_and2_1 _1578_ (.A(_0687_),
    .B(_0688_),
    .X(_0689_));
 sg13g2_nor2_1 _1579_ (.A(_0687_),
    .B(_0688_),
    .Y(_0690_));
 sg13g2_nor3_1 _1580_ (.A(net199),
    .B(_0689_),
    .C(_0690_),
    .Y(_0052_));
 sg13g2_a21oi_1 _1581_ (.A1(net483),
    .A2(\VAL[4] ),
    .Y(_0691_),
    .B1(_0690_));
 sg13g2_nor2_1 _1582_ (.A(net276),
    .B(_0691_),
    .Y(_0692_));
 sg13g2_a21oi_1 _1583_ (.A1(net276),
    .A2(_0691_),
    .Y(_0693_),
    .B1(net199));
 sg13g2_nor2b_1 _1584_ (.A(_0692_),
    .B_N(net277),
    .Y(_0053_));
 sg13g2_nand2_1 _1585_ (.Y(_0694_),
    .A(net421),
    .B(_0692_));
 sg13g2_o21ai_1 _1586_ (.B1(net207),
    .Y(_0695_),
    .A1(net421),
    .A2(_0692_));
 sg13g2_nor2b_1 _1587_ (.A(_0695_),
    .B_N(_0694_),
    .Y(_0054_));
 sg13g2_o21ai_1 _1588_ (.B1(net207),
    .Y(_0696_),
    .A1(_0450_),
    .A2(_0694_));
 sg13g2_a21oi_1 _1589_ (.A1(_0450_),
    .A2(_0694_),
    .Y(_0055_),
    .B1(_0696_));
 sg13g2_nand2_1 _1590_ (.Y(_0697_),
    .A(net181),
    .B(net422));
 sg13g2_o21ai_1 _1591_ (.B1(net207),
    .Y(_0698_),
    .A1(net181),
    .A2(net422));
 sg13g2_nor2b_1 _1592_ (.A(net423),
    .B_N(_0697_),
    .Y(_0056_));
 sg13g2_xnor2_1 _1593_ (.Y(_0699_),
    .A(net180),
    .B(net471));
 sg13g2_and2_1 _1594_ (.A(_0697_),
    .B(_0699_),
    .X(_0700_));
 sg13g2_nor2_1 _1595_ (.A(_0697_),
    .B(_0699_),
    .Y(_0701_));
 sg13g2_nor3_1 _1596_ (.A(net199),
    .B(_0700_),
    .C(_0701_),
    .Y(_0057_));
 sg13g2_xnor2_1 _1597_ (.Y(_0702_),
    .A(net472),
    .B(net479));
 sg13g2_a21oi_1 _1598_ (.A1(net180),
    .A2(net471),
    .Y(_0703_),
    .B1(_0701_));
 sg13g2_and2_1 _1599_ (.A(_0702_),
    .B(_0703_),
    .X(_0704_));
 sg13g2_nor2_1 _1600_ (.A(_0702_),
    .B(_0703_),
    .Y(_0705_));
 sg13g2_nor3_1 _1601_ (.A(net199),
    .B(_0704_),
    .C(_0705_),
    .Y(_0058_));
 sg13g2_xnor2_1 _1602_ (.Y(_0706_),
    .A(net177),
    .B(net447));
 sg13g2_a21oi_1 _1603_ (.A1(\hvsync_gen.vpos[6] ),
    .A2(\VAL[10] ),
    .Y(_0707_),
    .B1(_0705_));
 sg13g2_or2_1 _1604_ (.X(_0708_),
    .B(_0707_),
    .A(_0706_));
 sg13g2_inv_1 _1605_ (.Y(_0709_),
    .A(_0708_));
 sg13g2_nand2_1 _1606_ (.Y(_0710_),
    .A(net207),
    .B(_0708_));
 sg13g2_a21oi_1 _1607_ (.A1(net448),
    .A2(_0707_),
    .Y(_0059_),
    .B1(_0710_));
 sg13g2_xnor2_1 _1608_ (.Y(_0711_),
    .A(net175),
    .B(net477));
 sg13g2_a21oi_1 _1609_ (.A1(net177),
    .A2(net447),
    .Y(_0712_),
    .B1(_0709_));
 sg13g2_and2_1 _1610_ (.A(_0711_),
    .B(_0712_),
    .X(_0713_));
 sg13g2_nor2_1 _1611_ (.A(_0711_),
    .B(_0712_),
    .Y(_0714_));
 sg13g2_nor3_1 _1612_ (.A(net199),
    .B(_0713_),
    .C(_0714_),
    .Y(_0060_));
 sg13g2_a21oi_1 _1613_ (.A1(net175),
    .A2(net487),
    .Y(_0715_),
    .B1(_0714_));
 sg13g2_nor2_2 _1614_ (.A(net307),
    .B(_0715_),
    .Y(_0716_));
 sg13g2_a21oi_1 _1615_ (.A1(net307),
    .A2(_0715_),
    .Y(_0717_),
    .B1(net199));
 sg13g2_nor2b_1 _1616_ (.A(_0716_),
    .B_N(net308),
    .Y(_0061_));
 sg13g2_o21ai_1 _1617_ (.B1(net207),
    .Y(_0718_),
    .A1(_0454_),
    .A2(_0716_));
 sg13g2_a21oi_1 _1618_ (.A1(_0454_),
    .A2(_0716_),
    .Y(_0062_),
    .B1(_0718_));
 sg13g2_a21oi_1 _1619_ (.A1(\VAL[14] ),
    .A2(_0716_),
    .Y(_0719_),
    .B1(net323));
 sg13g2_and3_1 _1620_ (.X(_0720_),
    .A(\VAL[14] ),
    .B(net323),
    .C(_0716_));
 sg13g2_nor3_1 _1621_ (.A(net199),
    .B(net324),
    .C(_0720_),
    .Y(_0063_));
 sg13g2_nor2_2 _1622_ (.A(net200),
    .B(net174),
    .Y(_0721_));
 sg13g2_nand2b_2 _1623_ (.Y(_0722_),
    .B(net206),
    .A_N(net173));
 sg13g2_nand2_1 _1624_ (.Y(_0723_),
    .A(_0423_),
    .B(net300));
 sg13g2_nand2_1 _1625_ (.Y(_0724_),
    .A(\hvsync_gen.vpos[2] ),
    .B(\counter[0] ));
 sg13g2_nand2_1 _1626_ (.Y(_0725_),
    .A(\hvsync_gen.vpos[3] ),
    .B(\counter[1] ));
 sg13g2_xnor2_1 _1627_ (.Y(_0726_),
    .A(\hvsync_gen.vpos[3] ),
    .B(\counter[1] ));
 sg13g2_xnor2_1 _1628_ (.Y(_0727_),
    .A(_0724_),
    .B(_0726_));
 sg13g2_or2_1 _1629_ (.X(_0728_),
    .B(net163),
    .A(net176));
 sg13g2_nand2_1 _1630_ (.Y(_0729_),
    .A(\hvsync_gen.vpos[5] ),
    .B(\counter[3] ));
 sg13g2_and2_1 _1631_ (.A(net182),
    .B(\counter[2] ),
    .X(_0730_));
 sg13g2_xor2_1 _1632_ (.B(\counter[2] ),
    .A(net182),
    .X(_0731_));
 sg13g2_o21ai_1 _1633_ (.B1(_0725_),
    .Y(_0732_),
    .A1(_0724_),
    .A2(_0726_));
 sg13g2_a21oi_1 _1634_ (.A1(_0731_),
    .A2(_0732_),
    .Y(_0733_),
    .B1(_0730_));
 sg13g2_nor2_1 _1635_ (.A(net180),
    .B(\counter[3] ),
    .Y(_0734_));
 sg13g2_xor2_1 _1636_ (.B(\counter[3] ),
    .A(net180),
    .X(_0735_));
 sg13g2_o21ai_1 _1637_ (.B1(_0729_),
    .Y(_0736_),
    .A1(_0733_),
    .A2(_0734_));
 sg13g2_and2_1 _1638_ (.A(net178),
    .B(\counter[4] ),
    .X(_0737_));
 sg13g2_xor2_1 _1639_ (.B(\counter[4] ),
    .A(net178),
    .X(_0738_));
 sg13g2_inv_1 _1640_ (.Y(_0739_),
    .A(_0738_));
 sg13g2_and2_1 _1641_ (.A(net177),
    .B(\counter[5] ),
    .X(_0740_));
 sg13g2_xnor2_1 _1642_ (.Y(_0741_),
    .A(net176),
    .B(\counter[5] ));
 sg13g2_nor2_1 _1643_ (.A(_0739_),
    .B(_0741_),
    .Y(_0742_));
 sg13g2_a221oi_1 _1644_ (.B2(_0736_),
    .C1(_0740_),
    .B1(_0742_),
    .A1(_0728_),
    .Y(_0743_),
    .A2(_0737_));
 sg13g2_xor2_1 _1645_ (.B(\counter[6] ),
    .A(net175),
    .X(_0744_));
 sg13g2_xnor2_1 _1646_ (.Y(_0745_),
    .A(_0743_),
    .B(_0744_));
 sg13g2_xnor2_1 _1647_ (.Y(_0746_),
    .A(_0727_),
    .B(_0745_));
 sg13g2_nand2_1 _1648_ (.Y(_0747_),
    .A(net306),
    .B(_0746_));
 sg13g2_o21ai_1 _1649_ (.B1(net187),
    .Y(_0748_),
    .A1(net306),
    .A2(_0746_));
 sg13g2_nand2b_1 _1650_ (.Y(_0749_),
    .B(_0747_),
    .A_N(_0748_));
 sg13g2_a21oi_1 _1651_ (.A1(_0723_),
    .A2(_0749_),
    .Y(_0064_),
    .B1(net167));
 sg13g2_nand2_1 _1652_ (.Y(_0750_),
    .A(net171),
    .B(net303));
 sg13g2_xor2_1 _1653_ (.B(_0732_),
    .A(_0731_),
    .X(_0751_));
 sg13g2_xnor2_1 _1654_ (.Y(_0752_),
    .A(_0745_),
    .B(_0751_));
 sg13g2_nor2b_1 _1655_ (.A(\yqo[1] ),
    .B_N(_0752_),
    .Y(_0753_));
 sg13g2_xor2_1 _1656_ (.B(_0752_),
    .A(\yqo[1] ),
    .X(_0754_));
 sg13g2_nor2b_1 _1657_ (.A(_0747_),
    .B_N(_0754_),
    .Y(_0755_));
 sg13g2_nand2b_1 _1658_ (.Y(_0756_),
    .B(_0747_),
    .A_N(_0754_));
 sg13g2_nand3b_1 _1659_ (.B(_0756_),
    .C(net187),
    .Y(_0757_),
    .A_N(_0755_));
 sg13g2_a21oi_1 _1660_ (.A1(_0750_),
    .A2(_0757_),
    .Y(_0065_),
    .B1(_0722_));
 sg13g2_nand2_1 _1661_ (.Y(_0758_),
    .A(net171),
    .B(net309));
 sg13g2_xnor2_1 _1662_ (.Y(_0759_),
    .A(_0733_),
    .B(_0735_));
 sg13g2_xnor2_1 _1663_ (.Y(_0760_),
    .A(_0745_),
    .B(_0759_));
 sg13g2_nand2b_1 _1664_ (.Y(_0761_),
    .B(\yqo[2] ),
    .A_N(_0760_));
 sg13g2_xnor2_1 _1665_ (.Y(_0762_),
    .A(\yqo[2] ),
    .B(_0760_));
 sg13g2_nor2b_1 _1666_ (.A(_0753_),
    .B_N(_0762_),
    .Y(_0763_));
 sg13g2_nand2b_1 _1667_ (.Y(_0764_),
    .B(_0753_),
    .A_N(_0762_));
 sg13g2_nor2b_1 _1668_ (.A(_0763_),
    .B_N(_0764_),
    .Y(_0765_));
 sg13g2_o21ai_1 _1669_ (.B1(net187),
    .Y(_0766_),
    .A1(_0755_),
    .A2(_0765_));
 sg13g2_a21o_1 _1670_ (.A2(_0765_),
    .A1(_0755_),
    .B1(_0766_),
    .X(_0767_));
 sg13g2_a21oi_1 _1671_ (.A1(_0758_),
    .A2(_0767_),
    .Y(_0066_),
    .B1(net168));
 sg13g2_nand2_1 _1672_ (.Y(_0768_),
    .A(net171),
    .B(net335));
 sg13g2_a21oi_1 _1673_ (.A1(_0755_),
    .A2(_0764_),
    .Y(_0769_),
    .B1(_0763_));
 sg13g2_xnor2_1 _1674_ (.Y(_0770_),
    .A(_0736_),
    .B(_0738_));
 sg13g2_xnor2_1 _1675_ (.Y(_0771_),
    .A(_0745_),
    .B(_0770_));
 sg13g2_nor2_2 _1676_ (.A(\yqo[3] ),
    .B(_0771_),
    .Y(_0772_));
 sg13g2_xnor2_1 _1677_ (.Y(_0773_),
    .A(\yqo[3] ),
    .B(_0771_));
 sg13g2_nand2b_1 _1678_ (.Y(_0774_),
    .B(_0773_),
    .A_N(_0761_));
 sg13g2_xor2_1 _1679_ (.B(_0773_),
    .A(_0761_),
    .X(_0775_));
 sg13g2_xnor2_1 _1680_ (.Y(_0776_),
    .A(_0769_),
    .B(_0775_));
 sg13g2_o21ai_1 _1681_ (.B1(_0768_),
    .Y(_0777_),
    .A1(net171),
    .A2(_0776_));
 sg13g2_and2_1 _1682_ (.A(_0721_),
    .B(_0777_),
    .X(_0067_));
 sg13g2_nand2_1 _1683_ (.Y(_0778_),
    .A(net170),
    .B(net297));
 sg13g2_o21ai_1 _1684_ (.B1(_0774_),
    .Y(_0779_),
    .A1(_0769_),
    .A2(_0775_));
 sg13g2_a21oi_1 _1685_ (.A1(_0736_),
    .A2(_0738_),
    .Y(_0780_),
    .B1(_0737_));
 sg13g2_xnor2_1 _1686_ (.Y(_0781_),
    .A(_0741_),
    .B(_0780_));
 sg13g2_xnor2_1 _1687_ (.Y(_0782_),
    .A(_0745_),
    .B(_0781_));
 sg13g2_nand2_1 _1688_ (.Y(_0783_),
    .A(\yqo[4] ),
    .B(_0782_));
 sg13g2_xnor2_1 _1689_ (.Y(_0784_),
    .A(\yqo[4] ),
    .B(_0782_));
 sg13g2_nor2_1 _1690_ (.A(_0772_),
    .B(_0784_),
    .Y(_0785_));
 sg13g2_or2_1 _1691_ (.X(_0786_),
    .B(_0784_),
    .A(_0772_));
 sg13g2_xnor2_1 _1692_ (.Y(_0787_),
    .A(_0772_),
    .B(_0784_));
 sg13g2_nand2b_1 _1693_ (.Y(_0788_),
    .B(_0779_),
    .A_N(_0787_));
 sg13g2_nand2b_1 _1694_ (.Y(_0789_),
    .B(_0787_),
    .A_N(_0779_));
 sg13g2_nand3_1 _1695_ (.B(_0788_),
    .C(_0789_),
    .A(net185),
    .Y(_0790_));
 sg13g2_a21oi_1 _1696_ (.A1(_0778_),
    .A2(_0790_),
    .Y(_0068_),
    .B1(net167));
 sg13g2_nand2_1 _1697_ (.Y(_0791_),
    .A(net170),
    .B(net398));
 sg13g2_xor2_1 _1698_ (.B(_0783_),
    .A(_0002_),
    .X(_0792_));
 sg13g2_a21oi_1 _1699_ (.A1(_0786_),
    .A2(_0788_),
    .Y(_0793_),
    .B1(_0792_));
 sg13g2_nand3_1 _1700_ (.B(_0788_),
    .C(_0792_),
    .A(_0786_),
    .Y(_0794_));
 sg13g2_nand3b_1 _1701_ (.B(_0794_),
    .C(net186),
    .Y(_0795_),
    .A_N(_0793_));
 sg13g2_a21oi_1 _1702_ (.A1(_0791_),
    .A2(_0795_),
    .Y(_0069_),
    .B1(net167));
 sg13g2_nand2_1 _1703_ (.Y(_0796_),
    .A(net170),
    .B(net415));
 sg13g2_nand2b_1 _1704_ (.Y(_0797_),
    .B(\yqo[5] ),
    .A_N(\yqo[6] ));
 sg13g2_xnor2_1 _1705_ (.Y(_0798_),
    .A(\yqo[6] ),
    .B(\yqo[5] ));
 sg13g2_nor2_1 _1706_ (.A(\yqo[5] ),
    .B(_0783_),
    .Y(_0799_));
 sg13g2_o21ai_1 _1707_ (.B1(_0798_),
    .Y(_0800_),
    .A1(_0793_),
    .A2(_0799_));
 sg13g2_or3_1 _1708_ (.A(_0793_),
    .B(_0798_),
    .C(_0799_),
    .X(_0801_));
 sg13g2_nand3_1 _1709_ (.B(_0800_),
    .C(_0801_),
    .A(net185),
    .Y(_0802_));
 sg13g2_a21oi_1 _1710_ (.A1(_0796_),
    .A2(_0802_),
    .Y(_0070_),
    .B1(net165));
 sg13g2_nand2_1 _1711_ (.Y(_0803_),
    .A(net170),
    .B(net396));
 sg13g2_xor2_1 _1712_ (.B(\yqo[6] ),
    .A(\yqo[7] ),
    .X(_0804_));
 sg13g2_inv_1 _1713_ (.Y(_0805_),
    .A(_0804_));
 sg13g2_a21o_1 _1714_ (.A2(_0800_),
    .A1(_0797_),
    .B1(_0804_),
    .X(_0806_));
 sg13g2_nand3_1 _1715_ (.B(_0800_),
    .C(_0804_),
    .A(_0797_),
    .Y(_0807_));
 sg13g2_nand3_1 _1716_ (.B(_0806_),
    .C(_0807_),
    .A(net185),
    .Y(_0808_));
 sg13g2_a21oi_1 _1717_ (.A1(_0803_),
    .A2(_0808_),
    .Y(_0071_),
    .B1(net165));
 sg13g2_nand2_1 _1718_ (.Y(_0809_),
    .A(net171),
    .B(net436));
 sg13g2_nand2_1 _1719_ (.Y(_0810_),
    .A(_0798_),
    .B(_0805_));
 sg13g2_nor3_1 _1720_ (.A(_0787_),
    .B(_0792_),
    .C(_0810_),
    .Y(_0811_));
 sg13g2_a21oi_1 _1721_ (.A1(_0002_),
    .A2(_0785_),
    .Y(_0812_),
    .B1(_0799_));
 sg13g2_o21ai_1 _1722_ (.B1(_0426_),
    .Y(_0813_),
    .A1(\yqo[6] ),
    .A2(\yqo[5] ));
 sg13g2_o21ai_1 _1723_ (.B1(_0813_),
    .Y(_0814_),
    .A1(_0810_),
    .A2(_0812_));
 sg13g2_a21oi_1 _1724_ (.A1(_0779_),
    .A2(_0811_),
    .Y(_0815_),
    .B1(_0814_));
 sg13g2_xnor2_1 _1725_ (.Y(_0816_),
    .A(\yqo[8] ),
    .B(\yqo[7] ));
 sg13g2_nand2b_1 _1726_ (.Y(_0817_),
    .B(_0816_),
    .A_N(_0815_));
 sg13g2_nand2b_1 _1727_ (.Y(_0818_),
    .B(_0815_),
    .A_N(_0816_));
 sg13g2_nand3_1 _1728_ (.B(_0817_),
    .C(_0818_),
    .A(net184),
    .Y(_0819_));
 sg13g2_a21oi_1 _1729_ (.A1(_0809_),
    .A2(_0819_),
    .Y(_0072_),
    .B1(net165));
 sg13g2_nand2_1 _1730_ (.Y(_0820_),
    .A(net171),
    .B(net414));
 sg13g2_xor2_1 _1731_ (.B(\yqo[8] ),
    .A(\yqo[9] ),
    .X(_0821_));
 sg13g2_inv_1 _1732_ (.Y(_0822_),
    .A(_0821_));
 sg13g2_o21ai_1 _1733_ (.B1(_0817_),
    .Y(_0823_),
    .A1(\yqo[8] ),
    .A2(_0426_));
 sg13g2_xnor2_1 _1734_ (.Y(_0824_),
    .A(_0821_),
    .B(_0823_));
 sg13g2_nand2_1 _1735_ (.Y(_0825_),
    .A(net184),
    .B(_0824_));
 sg13g2_a21oi_1 _1736_ (.A1(_0820_),
    .A2(_0825_),
    .Y(_0073_),
    .B1(net166));
 sg13g2_nand2_1 _1737_ (.Y(_0826_),
    .A(net170),
    .B(net380));
 sg13g2_nand2_1 _1738_ (.Y(_0827_),
    .A(_0816_),
    .B(_0822_));
 sg13g2_o21ai_1 _1739_ (.B1(_0425_),
    .Y(_0828_),
    .A1(\yqo[8] ),
    .A2(\yqo[7] ));
 sg13g2_o21ai_1 _1740_ (.B1(_0828_),
    .Y(_0829_),
    .A1(_0815_),
    .A2(_0827_));
 sg13g2_nor2_1 _1741_ (.A(\yqo[10] ),
    .B(_0425_),
    .Y(_0830_));
 sg13g2_xnor2_1 _1742_ (.Y(_0831_),
    .A(\yqo[10] ),
    .B(\yqo[9] ));
 sg13g2_o21ai_1 _1743_ (.B1(net184),
    .Y(_0832_),
    .A1(_0829_),
    .A2(_0831_));
 sg13g2_a21o_1 _1744_ (.A2(_0831_),
    .A1(_0829_),
    .B1(_0832_),
    .X(_0833_));
 sg13g2_a21oi_1 _1745_ (.A1(_0826_),
    .A2(_0833_),
    .Y(_0074_),
    .B1(net166));
 sg13g2_nand2_1 _1746_ (.Y(_0834_),
    .A(net170),
    .B(net403));
 sg13g2_xor2_1 _1747_ (.B(\yqo[10] ),
    .A(\yqo[11] ),
    .X(_0835_));
 sg13g2_a21oi_1 _1748_ (.A1(_0829_),
    .A2(_0831_),
    .Y(_0836_),
    .B1(_0830_));
 sg13g2_a21oi_1 _1749_ (.A1(_0835_),
    .A2(_0836_),
    .Y(_0837_),
    .B1(net171));
 sg13g2_o21ai_1 _1750_ (.B1(_0837_),
    .Y(_0838_),
    .A1(_0835_),
    .A2(_0836_));
 sg13g2_a21oi_1 _1751_ (.A1(_0834_),
    .A2(_0838_),
    .Y(_0075_),
    .B1(net165));
 sg13g2_nand2_1 _1752_ (.Y(_0839_),
    .A(net339),
    .B(net170));
 sg13g2_nand3b_1 _1753_ (.B(_0829_),
    .C(_0831_),
    .Y(_0840_),
    .A_N(_0835_));
 sg13g2_o21ai_1 _1754_ (.B1(_0424_),
    .Y(_0841_),
    .A1(\yqo[10] ),
    .A2(\yqo[9] ));
 sg13g2_xor2_1 _1755_ (.B(\yqo[11] ),
    .A(\yqo[12] ),
    .X(_0842_));
 sg13g2_nand3_1 _1756_ (.B(_0841_),
    .C(_0842_),
    .A(_0840_),
    .Y(_0843_));
 sg13g2_a21o_1 _1757_ (.A2(_0841_),
    .A1(_0840_),
    .B1(_0842_),
    .X(_0844_));
 sg13g2_nand3_1 _1758_ (.B(_0843_),
    .C(_0844_),
    .A(net184),
    .Y(_0845_));
 sg13g2_a21oi_1 _1759_ (.A1(_0839_),
    .A2(_0845_),
    .Y(_0076_),
    .B1(net165));
 sg13g2_nand2_1 _1760_ (.Y(_0846_),
    .A(net187),
    .B(\yqo[0] ));
 sg13g2_a21oi_1 _1761_ (.A1(_0723_),
    .A2(_0846_),
    .Y(_0077_),
    .B1(net167));
 sg13g2_nand2_1 _1762_ (.Y(_0847_),
    .A(net187),
    .B(net345));
 sg13g2_a21oi_1 _1763_ (.A1(_0750_),
    .A2(_0847_),
    .Y(_0078_),
    .B1(net167));
 sg13g2_nand2_1 _1764_ (.Y(_0848_),
    .A(net187),
    .B(net311));
 sg13g2_a21oi_1 _1765_ (.A1(_0758_),
    .A2(_0848_),
    .Y(_0079_),
    .B1(net168));
 sg13g2_nand2_1 _1766_ (.Y(_0849_),
    .A(net187),
    .B(\yqo[3] ));
 sg13g2_a21oi_1 _1767_ (.A1(_0768_),
    .A2(_0849_),
    .Y(_0080_),
    .B1(_0722_));
 sg13g2_nand2_1 _1768_ (.Y(_0850_),
    .A(net185),
    .B(\yqo[4] ));
 sg13g2_a21oi_1 _1769_ (.A1(_0778_),
    .A2(_0850_),
    .Y(_0081_),
    .B1(net168));
 sg13g2_nand2_1 _1770_ (.Y(_0851_),
    .A(net186),
    .B(\yqo[5] ));
 sg13g2_a21oi_1 _1771_ (.A1(_0791_),
    .A2(_0851_),
    .Y(_0082_),
    .B1(net167));
 sg13g2_nand2_1 _1772_ (.Y(_0852_),
    .A(net185),
    .B(\yqo[6] ));
 sg13g2_a21oi_1 _1773_ (.A1(_0796_),
    .A2(_0852_),
    .Y(_0083_),
    .B1(net165));
 sg13g2_nand2_1 _1774_ (.Y(_0853_),
    .A(net184),
    .B(net397));
 sg13g2_a21oi_1 _1775_ (.A1(_0803_),
    .A2(_0853_),
    .Y(_0084_),
    .B1(net166));
 sg13g2_nand2_1 _1776_ (.Y(_0854_),
    .A(net185),
    .B(net432));
 sg13g2_a21oi_1 _1777_ (.A1(_0809_),
    .A2(_0854_),
    .Y(_0085_),
    .B1(net166));
 sg13g2_nand2_1 _1778_ (.Y(_0855_),
    .A(net184),
    .B(net424));
 sg13g2_a21oi_1 _1779_ (.A1(_0820_),
    .A2(_0855_),
    .Y(_0086_),
    .B1(net166));
 sg13g2_nand2_1 _1780_ (.Y(_0856_),
    .A(net184),
    .B(net401));
 sg13g2_a21oi_1 _1781_ (.A1(_0826_),
    .A2(_0856_),
    .Y(_0087_),
    .B1(net166));
 sg13g2_nand2_1 _1782_ (.Y(_0857_),
    .A(net184),
    .B(\yqo[11] ));
 sg13g2_a21oi_1 _1783_ (.A1(_0834_),
    .A2(_0857_),
    .Y(_0088_),
    .B1(net165));
 sg13g2_nand2_1 _1784_ (.Y(_0858_),
    .A(net332),
    .B(net185));
 sg13g2_a21oi_1 _1785_ (.A1(_0839_),
    .A2(_0858_),
    .Y(_0089_),
    .B1(net165));
 sg13g2_a21oi_1 _1786_ (.A1(_0447_),
    .A2(net419),
    .Y(_0859_),
    .B1(net168));
 sg13g2_o21ai_1 _1787_ (.B1(_0859_),
    .Y(_0090_),
    .A1(net169),
    .A2(net419));
 sg13g2_and2_1 _1788_ (.A(net266),
    .B(_0721_),
    .X(_0091_));
 sg13g2_and2_1 _1789_ (.A(net419),
    .B(_0721_),
    .X(_0092_));
 sg13g2_nor2_1 _1790_ (.A(net169),
    .B(net168),
    .Y(_0093_));
 sg13g2_nor2_1 _1791_ (.A(_0445_),
    .B(net168),
    .Y(_0094_));
 sg13g2_nor2_1 _1792_ (.A(_0444_),
    .B(net168),
    .Y(_0095_));
 sg13g2_and2_1 _1793_ (.A(net190),
    .B(net163),
    .X(_0860_));
 sg13g2_nand2_1 _1794_ (.Y(_0861_),
    .A(net190),
    .B(net163));
 sg13g2_nor2_1 _1795_ (.A(net190),
    .B(net163),
    .Y(_0862_));
 sg13g2_nor2_1 _1796_ (.A(net192),
    .B(\counter[4] ),
    .Y(_0863_));
 sg13g2_nor2_1 _1797_ (.A(net193),
    .B(\counter[3] ),
    .Y(_0864_));
 sg13g2_nor2_1 _1798_ (.A(net195),
    .B(\counter[1] ),
    .Y(_0865_));
 sg13g2_nor2_1 _1799_ (.A(net194),
    .B(\counter[2] ),
    .Y(_0866_));
 sg13g2_nor3_1 _1800_ (.A(_0864_),
    .B(_0865_),
    .C(_0866_),
    .Y(_0867_));
 sg13g2_a22oi_1 _1801_ (.Y(_0868_),
    .B1(\counter[1] ),
    .B2(net195),
    .A2(\counter[0] ),
    .A1(\hvsync_gen.hpos[3] ));
 sg13g2_a22oi_1 _1802_ (.Y(_0869_),
    .B1(\counter[3] ),
    .B2(net193),
    .A2(\counter[2] ),
    .A1(net194));
 sg13g2_nor2b_1 _1803_ (.A(_0868_),
    .B_N(_0869_),
    .Y(_0870_));
 sg13g2_nor2_1 _1804_ (.A(_0864_),
    .B(_0869_),
    .Y(_0871_));
 sg13g2_a221oi_1 _1805_ (.B2(_0870_),
    .C1(_0871_),
    .B1(_0867_),
    .A1(net192),
    .Y(_0872_),
    .A2(\counter[4] ));
 sg13g2_or2_1 _1806_ (.X(_0873_),
    .B(_0872_),
    .A(_0863_));
 sg13g2_or4_1 _1807_ (.A(_0860_),
    .B(_0862_),
    .C(_0863_),
    .D(_0872_),
    .X(_0874_));
 sg13g2_o21ai_1 _1808_ (.B1(_0873_),
    .Y(_0875_),
    .A1(_0860_),
    .A2(_0862_));
 sg13g2_and2_1 _1809_ (.A(_0874_),
    .B(_0875_),
    .X(_0876_));
 sg13g2_and2_1 _1810_ (.A(net189),
    .B(\counter[6] ),
    .X(_0877_));
 sg13g2_xnor2_1 _1811_ (.Y(_0878_),
    .A(net189),
    .B(\counter[6] ));
 sg13g2_a21oi_1 _1812_ (.A1(_0861_),
    .A2(_0874_),
    .Y(_0879_),
    .B1(_0878_));
 sg13g2_o21ai_1 _1813_ (.B1(\counter[7] ),
    .Y(_0880_),
    .A1(_0877_),
    .A2(_0879_));
 sg13g2_xnor2_1 _1814_ (.Y(_0881_),
    .A(_0461_),
    .B(_0880_));
 sg13g2_xnor2_1 _1815_ (.Y(_0882_),
    .A(_0876_),
    .B(_0881_));
 sg13g2_or2_1 _1816_ (.X(_0883_),
    .B(_0882_),
    .A(net438));
 sg13g2_nand2_1 _1817_ (.Y(_0884_),
    .A(net438),
    .B(_0882_));
 sg13g2_nor2_2 _1818_ (.A(net186),
    .B(net200),
    .Y(_0885_));
 sg13g2_nand2_2 _1819_ (.Y(_0886_),
    .A(net170),
    .B(net206));
 sg13g2_and3_1 _1820_ (.X(_0096_),
    .A(_0883_),
    .B(_0884_),
    .C(_0885_));
 sg13g2_nand3_1 _1821_ (.B(_0874_),
    .C(_0878_),
    .A(_0861_),
    .Y(_0887_));
 sg13g2_nor2b_1 _1822_ (.A(_0879_),
    .B_N(_0887_),
    .Y(_0888_));
 sg13g2_xnor2_1 _1823_ (.Y(_0889_),
    .A(_0881_),
    .B(_0888_));
 sg13g2_nor2_1 _1824_ (.A(net455),
    .B(_0889_),
    .Y(_0890_));
 sg13g2_xnor2_1 _1825_ (.Y(_0891_),
    .A(net455),
    .B(_0889_));
 sg13g2_nand2b_1 _1826_ (.Y(_0892_),
    .B(_0884_),
    .A_N(_0891_));
 sg13g2_nand2b_1 _1827_ (.Y(_0893_),
    .B(_0891_),
    .A_N(_0884_));
 sg13g2_and3_1 _1828_ (.X(_0097_),
    .A(_0885_),
    .B(_0892_),
    .C(_0893_));
 sg13g2_nor3_1 _1829_ (.A(\counter[7] ),
    .B(_0877_),
    .C(_0879_),
    .Y(_0894_));
 sg13g2_xnor2_1 _1830_ (.Y(_0895_),
    .A(\counter[8] ),
    .B(_0894_));
 sg13g2_nor2_1 _1831_ (.A(\xqo[2] ),
    .B(_0895_),
    .Y(_0896_));
 sg13g2_xor2_1 _1832_ (.B(_0895_),
    .A(\xqo[2] ),
    .X(_0897_));
 sg13g2_or2_1 _1833_ (.X(_0898_),
    .B(_0897_),
    .A(_0890_));
 sg13g2_xnor2_1 _1834_ (.Y(_0899_),
    .A(_0890_),
    .B(_0897_));
 sg13g2_o21ai_1 _1835_ (.B1(_0885_),
    .Y(_0900_),
    .A1(_0893_),
    .A2(_0899_));
 sg13g2_a21oi_1 _1836_ (.A1(_0893_),
    .A2(_0899_),
    .Y(_0098_),
    .B1(_0900_));
 sg13g2_o21ai_1 _1837_ (.B1(_0898_),
    .Y(_0901_),
    .A1(_0893_),
    .A2(_0899_));
 sg13g2_o21ai_1 _1838_ (.B1(\xqo[3] ),
    .Y(_0902_),
    .A1(\xqo[2] ),
    .A2(_0895_));
 sg13g2_inv_1 _1839_ (.Y(_0903_),
    .A(_0902_));
 sg13g2_xnor2_1 _1840_ (.Y(_0904_),
    .A(net481),
    .B(_0896_));
 sg13g2_or2_1 _1841_ (.X(_0905_),
    .B(_0904_),
    .A(_0901_));
 sg13g2_a21oi_1 _1842_ (.A1(_0901_),
    .A2(_0904_),
    .Y(_0906_),
    .B1(_0886_));
 sg13g2_and2_1 _1843_ (.A(_0905_),
    .B(_0906_),
    .X(_0099_));
 sg13g2_a21o_1 _1844_ (.A2(_0904_),
    .A1(_0901_),
    .B1(_0903_),
    .X(_0907_));
 sg13g2_or2_1 _1845_ (.X(_0908_),
    .B(_0907_),
    .A(net289));
 sg13g2_nand2_1 _1846_ (.Y(_0909_),
    .A(net289),
    .B(_0907_));
 sg13g2_a21oi_1 _1847_ (.A1(_0908_),
    .A2(net290),
    .Y(_0100_),
    .B1(_0886_));
 sg13g2_o21ai_1 _1848_ (.B1(net366),
    .Y(_0910_),
    .A1(net289),
    .A2(_0907_));
 sg13g2_and2_1 _1849_ (.A(_0885_),
    .B(_0910_),
    .X(_0911_));
 sg13g2_o21ai_1 _1850_ (.B1(_0911_),
    .Y(_0912_),
    .A1(net366),
    .A2(_0908_));
 sg13g2_inv_1 _1851_ (.Y(_0101_),
    .A(_0912_));
 sg13g2_or2_1 _1852_ (.X(_0913_),
    .B(_0910_),
    .A(_0462_));
 sg13g2_nand2_1 _1853_ (.Y(_0914_),
    .A(_0885_),
    .B(_0913_));
 sg13g2_a21oi_1 _1854_ (.A1(_0462_),
    .A2(_0910_),
    .Y(_0102_),
    .B1(_0914_));
 sg13g2_and2_1 _1855_ (.A(_0463_),
    .B(_0913_),
    .X(_0915_));
 sg13g2_nor2_1 _1856_ (.A(_0463_),
    .B(_0913_),
    .Y(_0916_));
 sg13g2_nor3_1 _1857_ (.A(_0886_),
    .B(_0915_),
    .C(_0916_),
    .Y(_0103_));
 sg13g2_nor4_2 _1858_ (.A(_0462_),
    .B(_0463_),
    .C(_0464_),
    .Y(_0917_),
    .D(_0910_));
 sg13g2_o21ai_1 _1859_ (.B1(_0885_),
    .Y(_0918_),
    .A1(net372),
    .A2(_0916_));
 sg13g2_nor2_1 _1860_ (.A(_0917_),
    .B(net373),
    .Y(_0104_));
 sg13g2_xnor2_1 _1861_ (.Y(_0919_),
    .A(net375),
    .B(_0917_));
 sg13g2_nor2_1 _1862_ (.A(_0886_),
    .B(net376),
    .Y(_0105_));
 sg13g2_a21oi_1 _1863_ (.A1(\xqo[9] ),
    .A2(_0917_),
    .Y(_0920_),
    .B1(net273));
 sg13g2_and3_1 _1864_ (.X(_0921_),
    .A(\xqo[9] ),
    .B(net273),
    .C(_0917_));
 sg13g2_nor3_1 _1865_ (.A(_0886_),
    .B(net274),
    .C(_0921_),
    .Y(_0106_));
 sg13g2_o21ai_1 _1866_ (.B1(_0885_),
    .Y(_0922_),
    .A1(net245),
    .A2(_0921_));
 sg13g2_a21oi_1 _1867_ (.A1(net245),
    .A2(_0921_),
    .Y(_0107_),
    .B1(_0922_));
 sg13g2_nor4_1 _1868_ (.A(\ctr_clkdiv25[5] ),
    .B(_0441_),
    .C(\ctr_clkdiv25[7] ),
    .D(net484),
    .Y(_0923_));
 sg13g2_nor4_1 _1869_ (.A(_0427_),
    .B(\ctr_clkdiv25[1] ),
    .C(\ctr_clkdiv25[2] ),
    .D(_0440_),
    .Y(_0924_));
 sg13g2_and2_1 _1870_ (.A(net485),
    .B(_0924_),
    .X(_0925_));
 sg13g2_nor2_1 _1871_ (.A(net196),
    .B(_0925_),
    .Y(_0926_));
 sg13g2_nand2b_2 _1872_ (.Y(_0927_),
    .B(net201),
    .A_N(_0925_));
 sg13g2_and2_1 _1873_ (.A(net201),
    .B(net486),
    .X(_0187_));
 sg13g2_a22oi_1 _1874_ (.Y(_0928_),
    .B1(_0187_),
    .B2(net237),
    .A2(_0926_),
    .A1(\ctr_audio[0] ));
 sg13g2_inv_1 _1875_ (.Y(_0108_),
    .A(net238));
 sg13g2_a21oi_1 _1876_ (.A1(\ctr_audio[0] ),
    .A2(_0925_),
    .Y(_0929_),
    .B1(net253));
 sg13g2_nand4_1 _1877_ (.B(\ctr_audio[0] ),
    .C(_0923_),
    .A(net253),
    .Y(_0930_),
    .D(_0924_));
 sg13g2_nand2_1 _1878_ (.Y(_0931_),
    .A(net201),
    .B(_0930_));
 sg13g2_nor2_1 _1879_ (.A(net254),
    .B(_0931_),
    .Y(_0109_));
 sg13g2_and2_1 _1880_ (.A(_0422_),
    .B(_0930_),
    .X(_0932_));
 sg13g2_nor2_1 _1881_ (.A(_0422_),
    .B(_0930_),
    .Y(_0933_));
 sg13g2_nor3_1 _1882_ (.A(net196),
    .B(net452),
    .C(_0933_),
    .Y(_0110_));
 sg13g2_o21ai_1 _1883_ (.B1(net201),
    .Y(_0934_),
    .A1(net286),
    .A2(_0933_));
 sg13g2_a21oi_1 _1884_ (.A1(net286),
    .A2(_0933_),
    .Y(_0111_),
    .B1(_0934_));
 sg13g2_a21oi_1 _1885_ (.A1(\ctr_audio[3] ),
    .A2(_0933_),
    .Y(_0935_),
    .B1(net258));
 sg13g2_nor4_2 _1886_ (.A(_0420_),
    .B(_0421_),
    .C(_0422_),
    .Y(_0936_),
    .D(_0930_));
 sg13g2_nor3_1 _1887_ (.A(net196),
    .B(net259),
    .C(_0936_),
    .Y(_0112_));
 sg13g2_and2_1 _1888_ (.A(net367),
    .B(_0936_),
    .X(_0937_));
 sg13g2_o21ai_1 _1889_ (.B1(net201),
    .Y(_0938_),
    .A1(net367),
    .A2(_0936_));
 sg13g2_nor2_1 _1890_ (.A(_0937_),
    .B(net368),
    .Y(_0113_));
 sg13g2_xnor2_1 _1891_ (.Y(_0939_),
    .A(net412),
    .B(_0937_));
 sg13g2_nor2_1 _1892_ (.A(net196),
    .B(_0939_),
    .Y(_0114_));
 sg13g2_a21oi_1 _1893_ (.A1(\ctr_audio[6] ),
    .A2(_0937_),
    .Y(_0940_),
    .B1(net291));
 sg13g2_nand3_1 _1894_ (.B(\ctr_audio[6] ),
    .C(_0937_),
    .A(net291),
    .Y(_0941_));
 sg13g2_nand2_1 _1895_ (.Y(_0942_),
    .A(net201),
    .B(_0941_));
 sg13g2_nor2_1 _1896_ (.A(net292),
    .B(_0942_),
    .Y(_0115_));
 sg13g2_nor2b_1 _1897_ (.A(net320),
    .B_N(_0941_),
    .Y(_0188_));
 sg13g2_and4_1 _1898_ (.A(net320),
    .B(net291),
    .C(\ctr_audio[6] ),
    .D(_0937_),
    .X(_0189_));
 sg13g2_nor3_1 _1899_ (.A(net196),
    .B(net321),
    .C(_0189_),
    .Y(_0116_));
 sg13g2_and2_1 _1900_ (.A(net384),
    .B(_0189_),
    .X(_0190_));
 sg13g2_o21ai_1 _1901_ (.B1(net203),
    .Y(_0191_),
    .A1(net384),
    .A2(_0189_));
 sg13g2_nor2_1 _1902_ (.A(_0190_),
    .B(net385),
    .Y(_0117_));
 sg13g2_xnor2_1 _1903_ (.Y(_0192_),
    .A(net402),
    .B(_0190_));
 sg13g2_nor2_1 _1904_ (.A(net196),
    .B(_0192_),
    .Y(_0118_));
 sg13g2_a21oi_1 _1905_ (.A1(\Voice1.pulsewidth[0] ),
    .A2(_0190_),
    .Y(_0193_),
    .B1(net341));
 sg13g2_and3_1 _1906_ (.X(_0194_),
    .A(net341),
    .B(\Voice1.pulsewidth[0] ),
    .C(_0190_));
 sg13g2_nor3_1 _1907_ (.A(net196),
    .B(net342),
    .C(_0194_),
    .Y(_0119_));
 sg13g2_or2_1 _1908_ (.X(_0195_),
    .B(_0194_),
    .A(net469));
 sg13g2_nand2_2 _1909_ (.Y(_0196_),
    .A(net469),
    .B(_0194_));
 sg13g2_and3_1 _1910_ (.X(_0120_),
    .A(net201),
    .B(_0195_),
    .C(_0196_));
 sg13g2_nor2_1 _1911_ (.A(_0419_),
    .B(_0196_),
    .Y(_0197_));
 sg13g2_a21oi_1 _1912_ (.A1(_0419_),
    .A2(_0196_),
    .Y(_0198_),
    .B1(net197));
 sg13g2_nor2b_1 _1913_ (.A(net467),
    .B_N(_0198_),
    .Y(_0121_));
 sg13g2_nor2_1 _1914_ (.A(net369),
    .B(_0197_),
    .Y(_0199_));
 sg13g2_nor3_2 _1915_ (.A(_0418_),
    .B(_0419_),
    .C(_0196_),
    .Y(_0200_));
 sg13g2_nor3_1 _1916_ (.A(net197),
    .B(net370),
    .C(_0200_),
    .Y(_0122_));
 sg13g2_and2_1 _1917_ (.A(net430),
    .B(_0200_),
    .X(_0201_));
 sg13g2_o21ai_1 _1918_ (.B1(net204),
    .Y(_0202_),
    .A1(net430),
    .A2(_0200_));
 sg13g2_nor2_1 _1919_ (.A(_0201_),
    .B(net431),
    .Y(_0123_));
 sg13g2_xnor2_1 _1920_ (.Y(_0203_),
    .A(net425),
    .B(_0201_));
 sg13g2_nor2_1 _1921_ (.A(net196),
    .B(net426),
    .Y(_0124_));
 sg13g2_a21oi_1 _1922_ (.A1(net425),
    .A2(_0201_),
    .Y(_0204_),
    .B1(net188));
 sg13g2_and3_1 _1923_ (.X(_0205_),
    .A(net188),
    .B(net425),
    .C(_0201_));
 sg13g2_nor3_1 _1924_ (.A(net198),
    .B(_0204_),
    .C(_0205_),
    .Y(_0125_));
 sg13g2_xnor2_1 _1925_ (.Y(_0206_),
    .A(net406),
    .B(_0205_));
 sg13g2_nor2_1 _1926_ (.A(net198),
    .B(net407),
    .Y(_0126_));
 sg13g2_a21oi_1 _1927_ (.A1(net406),
    .A2(_0205_),
    .Y(_0207_),
    .B1(net413));
 sg13g2_nand3_1 _1928_ (.B(net406),
    .C(_0205_),
    .A(net413),
    .Y(_0208_));
 sg13g2_nand2_1 _1929_ (.Y(_0209_),
    .A(net204),
    .B(_0208_));
 sg13g2_nor2_1 _1930_ (.A(_0207_),
    .B(_0209_),
    .Y(_0127_));
 sg13g2_and2_1 _1931_ (.A(_0414_),
    .B(_0208_),
    .X(_0210_));
 sg13g2_nor2_2 _1932_ (.A(_0414_),
    .B(_0208_),
    .Y(_0211_));
 sg13g2_nor3_1 _1933_ (.A(net198),
    .B(_0210_),
    .C(_0211_),
    .Y(_0128_));
 sg13g2_xnor2_1 _1934_ (.Y(_0212_),
    .A(net450),
    .B(_0211_));
 sg13g2_nor2_1 _1935_ (.A(net198),
    .B(_0212_),
    .Y(_0129_));
 sg13g2_a21o_1 _1936_ (.A2(_0211_),
    .A1(net450),
    .B1(net462),
    .X(_0213_));
 sg13g2_nand2_2 _1937_ (.Y(_0214_),
    .A(\ctr_audio[22] ),
    .B(\ctr_audio[21] ));
 sg13g2_nand3_1 _1938_ (.B(\ctr_audio[21] ),
    .C(_0211_),
    .A(net462),
    .Y(_0215_));
 sg13g2_and3_1 _1939_ (.X(_0130_),
    .A(net204),
    .B(_0213_),
    .C(_0215_));
 sg13g2_o21ai_1 _1940_ (.B1(net204),
    .Y(_0216_),
    .A1(_0413_),
    .A2(_0215_));
 sg13g2_a21oi_1 _1941_ (.A1(_0413_),
    .A2(_0215_),
    .Y(_0131_),
    .B1(_0216_));
 sg13g2_and2_1 _1942_ (.A(net203),
    .B(net242),
    .X(_0132_));
 sg13g2_and2_1 _1943_ (.A(net202),
    .B(net243),
    .X(_0133_));
 sg13g2_and2_1 _1944_ (.A(net202),
    .B(net244),
    .X(_0134_));
 sg13g2_and2_1 _1945_ (.A(net202),
    .B(net241),
    .X(_0135_));
 sg13g2_and2_1 _1946_ (.A(net202),
    .B(net344),
    .X(_0136_));
 sg13g2_and2_1 _1947_ (.A(net205),
    .B(net305),
    .X(_0137_));
 sg13g2_and2_1 _1948_ (.A(net205),
    .B(net288),
    .X(_0138_));
 sg13g2_and2_1 _1949_ (.A(net205),
    .B(net315),
    .X(_0139_));
 sg13g2_and2_1 _1950_ (.A(net202),
    .B(net282),
    .X(_0140_));
 sg13g2_and2_1 _1951_ (.A(net205),
    .B(net256),
    .X(_0141_));
 sg13g2_and2_1 _1952_ (.A(net205),
    .B(net337),
    .X(_0142_));
 sg13g2_and2_1 _1953_ (.A(net205),
    .B(net257),
    .X(_0143_));
 sg13g2_and2_1 _1954_ (.A(net236),
    .B(_0926_),
    .X(_0144_));
 sg13g2_xnor2_1 _1955_ (.Y(_0217_),
    .A(\ctr_clkdiv25[0] ),
    .B(net392));
 sg13g2_nor2_1 _1956_ (.A(_0927_),
    .B(net393),
    .Y(_0145_));
 sg13g2_and3_1 _1957_ (.X(_0218_),
    .A(\ctr_clkdiv25[0] ),
    .B(\ctr_clkdiv25[1] ),
    .C(net261));
 sg13g2_a21oi_1 _1958_ (.A1(\ctr_clkdiv25[0] ),
    .A2(\ctr_clkdiv25[1] ),
    .Y(_0219_),
    .B1(net261));
 sg13g2_nor3_1 _1959_ (.A(_0927_),
    .B(_0218_),
    .C(net262),
    .Y(_0146_));
 sg13g2_and2_1 _1960_ (.A(net329),
    .B(_0218_),
    .X(_0220_));
 sg13g2_nor2_1 _1961_ (.A(net329),
    .B(_0218_),
    .Y(_0221_));
 sg13g2_nor3_1 _1962_ (.A(_0927_),
    .B(_0220_),
    .C(net330),
    .Y(_0147_));
 sg13g2_and2_1 _1963_ (.A(net326),
    .B(_0220_),
    .X(_0222_));
 sg13g2_nor2_1 _1964_ (.A(net326),
    .B(_0220_),
    .Y(_0223_));
 sg13g2_nor3_1 _1965_ (.A(_0927_),
    .B(_0222_),
    .C(net327),
    .Y(_0148_));
 sg13g2_nor2_1 _1966_ (.A(net360),
    .B(_0222_),
    .Y(_0224_));
 sg13g2_and2_1 _1967_ (.A(net360),
    .B(_0222_),
    .X(_0225_));
 sg13g2_nor3_1 _1968_ (.A(_0927_),
    .B(_0224_),
    .C(_0225_),
    .Y(_0149_));
 sg13g2_nand2_1 _1969_ (.Y(_0226_),
    .A(net400),
    .B(_0225_));
 sg13g2_o21ai_1 _1970_ (.B1(_0926_),
    .Y(_0227_),
    .A1(net400),
    .A2(_0225_));
 sg13g2_nor2b_1 _1971_ (.A(_0227_),
    .B_N(_0226_),
    .Y(_0150_));
 sg13g2_xor2_1 _1972_ (.B(_0226_),
    .A(net381),
    .X(_0228_));
 sg13g2_nor2_1 _1973_ (.A(_0927_),
    .B(net382),
    .Y(_0151_));
 sg13g2_nand2_1 _1974_ (.Y(_0229_),
    .A(net188),
    .B(_0432_));
 sg13g2_nor2_1 _1975_ (.A(\Voice1.pulsewidth[6] ),
    .B(_0433_),
    .Y(_0230_));
 sg13g2_nor2_1 _1976_ (.A(\Voice1.pulsewidth[1] ),
    .B(_0429_),
    .Y(_0231_));
 sg13g2_nand2_1 _1977_ (.Y(_0232_),
    .A(\Voice1.pulsewidth[0] ),
    .B(_0428_));
 sg13g2_a22oi_1 _1978_ (.Y(_0233_),
    .B1(_0431_),
    .B2(\Voice1.pulsewidth[2] ),
    .A2(_0429_),
    .A1(\Voice1.pulsewidth[1] ));
 sg13g2_o21ai_1 _1979_ (.B1(_0233_),
    .Y(_0234_),
    .A1(_0231_),
    .A2(_0232_));
 sg13g2_o21ai_1 _1980_ (.B1(_0234_),
    .Y(_0235_),
    .A1(\Voice1.pulsewidth[2] ),
    .A2(_0431_));
 sg13g2_a21oi_1 _1981_ (.A1(_0419_),
    .A2(\Voice1.accumulator[15] ),
    .Y(_0236_),
    .B1(_0235_));
 sg13g2_a221oi_1 _1982_ (.B2(\Voice1.pulsewidth[4] ),
    .C1(_0236_),
    .B1(_0434_),
    .A1(\Voice1.pulsewidth[3] ),
    .Y(_0237_),
    .A2(_0430_));
 sg13g2_a221oi_1 _1983_ (.B2(_0417_),
    .C1(_0237_),
    .B1(\Voice1.accumulator[17] ),
    .A1(_0418_),
    .Y(_0238_),
    .A2(\Voice1.accumulator[16] ));
 sg13g2_a221oi_1 _1984_ (.B2(\Voice1.pulsewidth[5] ),
    .C1(_0238_),
    .B1(_0435_),
    .A1(\Voice1.pulsewidth[6] ),
    .Y(_0239_),
    .A2(_0433_));
 sg13g2_o21ai_1 _1985_ (.B1(_0229_),
    .Y(_0240_),
    .A1(_0230_),
    .A2(_0239_));
 sg13g2_a22oi_1 _1986_ (.Y(_0241_),
    .B1(\Voice1.accumulator[20] ),
    .B2(_0415_),
    .A2(\Voice1.accumulator[19] ),
    .A1(_0416_));
 sg13g2_o21ai_1 _1987_ (.B1(\Voice1.accumulator[21] ),
    .Y(_0242_),
    .A1(_0415_),
    .A2(\Voice1.accumulator[20] ));
 sg13g2_a221oi_1 _1988_ (.B2(_0241_),
    .C1(_0242_),
    .B1(_0240_),
    .A1(\Voice1.pulsewidth[10] ),
    .Y(_0243_),
    .A2(_0436_));
 sg13g2_nor2_1 _1989_ (.A(\Voice1.pulsewidth[10] ),
    .B(_0436_),
    .Y(_0244_));
 sg13g2_nor4_1 _1990_ (.A(_0412_),
    .B(net247),
    .C(_0243_),
    .D(_0244_),
    .Y(_0245_));
 sg13g2_o21ai_1 _1991_ (.B1(net204),
    .Y(_0246_),
    .A1(net363),
    .A2(net172));
 sg13g2_nor2_1 _1992_ (.A(_0245_),
    .B(net364),
    .Y(_0152_));
 sg13g2_nor2_1 _1993_ (.A(_0412_),
    .B(net198),
    .Y(_0247_));
 sg13g2_nand2_2 _1994_ (.Y(_0248_),
    .A(net172),
    .B(net204));
 sg13g2_nand2b_1 _1995_ (.Y(_0249_),
    .B(\ctr_audio[21] ),
    .A_N(\ctr_audio[22] ));
 sg13g2_a21o_1 _1996_ (.A2(_0249_),
    .A1(\Voice1.pulsewidth[7] ),
    .B1(\ctr_audio[19] ),
    .X(_0250_));
 sg13g2_nand3_1 _1997_ (.B(net188),
    .C(_0249_),
    .A(\ctr_audio[19] ),
    .Y(_0251_));
 sg13g2_nand2_2 _1998_ (.Y(_0252_),
    .A(_0250_),
    .B(_0251_));
 sg13g2_and2_1 _1999_ (.A(\ctr_audio[19] ),
    .B(net188),
    .X(_0253_));
 sg13g2_or3_2 _2000_ (.A(_0009_),
    .B(_0214_),
    .C(_0253_),
    .X(_0254_));
 sg13g2_and4_2 _2001_ (.A(\ctr_audio[22] ),
    .B(\ctr_audio[21] ),
    .C(\ctr_audio[19] ),
    .D(net188),
    .X(_0255_));
 sg13g2_nand2_1 _2002_ (.Y(_0256_),
    .A(_0009_),
    .B(_0255_));
 sg13g2_nand2_1 _2003_ (.Y(_0257_),
    .A(_0254_),
    .B(_0256_));
 sg13g2_nor2_1 _2004_ (.A(_0252_),
    .B(_0257_),
    .Y(_0258_));
 sg13g2_nand4_1 _2005_ (.B(_0251_),
    .C(_0254_),
    .A(_0250_),
    .Y(_0259_),
    .D(_0256_));
 sg13g2_nor2_2 _2006_ (.A(_0008_),
    .B(_0258_),
    .Y(_0260_));
 sg13g2_nand3_1 _2007_ (.B(_0456_),
    .C(_0259_),
    .A(_0455_),
    .Y(_0261_));
 sg13g2_o21ai_1 _2008_ (.B1(net160),
    .Y(_0262_),
    .A1(_0456_),
    .A2(_0260_));
 sg13g2_nor2b_1 _2009_ (.A(_0262_),
    .B_N(_0261_),
    .Y(_0263_));
 sg13g2_a21o_1 _2010_ (.A2(net164),
    .A1(net271),
    .B1(_0263_),
    .X(_0153_));
 sg13g2_o21ai_1 _2011_ (.B1(net188),
    .Y(_0264_),
    .A1(\ctr_audio[21] ),
    .A2(\ctr_audio[19] ));
 sg13g2_a21oi_1 _2012_ (.A1(_0214_),
    .A2(_0264_),
    .Y(_0265_),
    .B1(_0255_));
 sg13g2_a21o_1 _2013_ (.A2(_0264_),
    .A1(_0214_),
    .B1(_0255_),
    .X(_0266_));
 sg13g2_nand3_1 _2014_ (.B(_0251_),
    .C(_0266_),
    .A(_0250_),
    .Y(_0267_));
 sg13g2_nand2b_1 _2015_ (.Y(_0268_),
    .B(_0255_),
    .A_N(_0009_));
 sg13g2_and2_1 _2016_ (.A(_0455_),
    .B(_0268_),
    .X(_0269_));
 sg13g2_nand3_1 _2017_ (.B(_0267_),
    .C(_0269_),
    .A(net348),
    .Y(_0270_));
 sg13g2_a21oi_1 _2018_ (.A1(_0267_),
    .A2(_0269_),
    .Y(_0271_),
    .B1(\Voice1.accumulator[1] ));
 sg13g2_a21o_1 _2019_ (.A2(_0269_),
    .A1(_0267_),
    .B1(\Voice1.accumulator[1] ),
    .X(_0272_));
 sg13g2_nand2_1 _2020_ (.Y(_0273_),
    .A(_0270_),
    .B(_0272_));
 sg13g2_nor2_1 _2021_ (.A(net348),
    .B(net160),
    .Y(_0274_));
 sg13g2_xnor2_1 _2022_ (.Y(_0275_),
    .A(_0261_),
    .B(_0273_));
 sg13g2_a21oi_1 _2023_ (.A1(net160),
    .A2(_0275_),
    .Y(_0154_),
    .B1(_0274_));
 sg13g2_nor2_1 _2024_ (.A(net319),
    .B(net160),
    .Y(_0276_));
 sg13g2_a21oi_2 _2025_ (.B1(_0412_),
    .Y(_0277_),
    .A2(_0264_),
    .A1(_0214_));
 sg13g2_nand2_1 _2026_ (.Y(_0278_),
    .A(net319),
    .B(_0277_));
 sg13g2_inv_1 _2027_ (.Y(_0279_),
    .A(_0278_));
 sg13g2_or2_1 _2028_ (.X(_0280_),
    .B(_0277_),
    .A(\Voice1.accumulator[2] ));
 sg13g2_nand2_1 _2029_ (.Y(_0281_),
    .A(_0278_),
    .B(_0280_));
 sg13g2_o21ai_1 _2030_ (.B1(_0270_),
    .Y(_0282_),
    .A1(_0261_),
    .A2(_0271_));
 sg13g2_xor2_1 _2031_ (.B(_0282_),
    .A(_0281_),
    .X(_0283_));
 sg13g2_a21oi_1 _2032_ (.A1(net160),
    .A2(_0283_),
    .Y(_0155_),
    .B1(_0276_));
 sg13g2_nor2_1 _2033_ (.A(net350),
    .B(net160),
    .Y(_0284_));
 sg13g2_nand2b_1 _2034_ (.Y(_0285_),
    .B(_0257_),
    .A_N(_0250_));
 sg13g2_nand3_1 _2035_ (.B(_0260_),
    .C(_0285_),
    .A(net350),
    .Y(_0286_));
 sg13g2_a21oi_1 _2036_ (.A1(_0260_),
    .A2(_0285_),
    .Y(_0287_),
    .B1(\Voice1.accumulator[3] ));
 sg13g2_a21o_1 _2037_ (.A2(_0285_),
    .A1(_0260_),
    .B1(\Voice1.accumulator[3] ),
    .X(_0288_));
 sg13g2_nand2_1 _2038_ (.Y(_0289_),
    .A(_0286_),
    .B(_0288_));
 sg13g2_a21oi_1 _2039_ (.A1(_0280_),
    .A2(_0282_),
    .Y(_0290_),
    .B1(_0279_));
 sg13g2_xnor2_1 _2040_ (.Y(_0291_),
    .A(_0289_),
    .B(_0290_));
 sg13g2_a21oi_1 _2041_ (.A1(net160),
    .A2(_0291_),
    .Y(_0156_),
    .B1(_0284_));
 sg13g2_o21ai_1 _2042_ (.B1(_0286_),
    .Y(_0292_),
    .A1(_0287_),
    .A2(_0290_));
 sg13g2_nor2b_1 _2043_ (.A(_0254_),
    .B_N(_0277_),
    .Y(_0293_));
 sg13g2_nand2_1 _2044_ (.Y(_0294_),
    .A(\Voice1.accumulator[4] ),
    .B(_0293_));
 sg13g2_inv_1 _2045_ (.Y(_0295_),
    .A(_0294_));
 sg13g2_or2_1 _2046_ (.X(_0296_),
    .B(_0293_),
    .A(\Voice1.accumulator[4] ));
 sg13g2_and2_1 _2047_ (.A(_0294_),
    .B(_0296_),
    .X(_0297_));
 sg13g2_xor2_1 _2048_ (.B(_0297_),
    .A(_0292_),
    .X(_0298_));
 sg13g2_mux2_1 _2049_ (.A0(net312),
    .A1(_0298_),
    .S(net160),
    .X(_0157_));
 sg13g2_a21oi_1 _2050_ (.A1(_0292_),
    .A2(_0296_),
    .Y(_0299_),
    .B1(_0295_));
 sg13g2_nor2_1 _2051_ (.A(_0252_),
    .B(_0266_),
    .Y(_0300_));
 sg13g2_nand3_1 _2052_ (.B(_0256_),
    .C(_0265_),
    .A(_0254_),
    .Y(_0301_));
 sg13g2_nor3_2 _2053_ (.A(_0008_),
    .B(_0252_),
    .C(_0301_),
    .Y(_0302_));
 sg13g2_nand2_1 _2054_ (.Y(_0303_),
    .A(net482),
    .B(_0302_));
 sg13g2_xnor2_1 _2055_ (.Y(_0304_),
    .A(net334),
    .B(_0302_));
 sg13g2_xnor2_1 _2056_ (.Y(_0305_),
    .A(_0299_),
    .B(_0304_));
 sg13g2_nand2_1 _2057_ (.Y(_0306_),
    .A(net334),
    .B(net164));
 sg13g2_o21ai_1 _2058_ (.B1(_0306_),
    .Y(_0158_),
    .A1(net164),
    .A2(_0305_));
 sg13g2_a21o_1 _2059_ (.A2(_0301_),
    .A1(_0268_),
    .B1(_0412_),
    .X(_0307_));
 sg13g2_nor2_1 _2060_ (.A(_0457_),
    .B(_0307_),
    .Y(_0308_));
 sg13g2_nand2_1 _2061_ (.Y(_0309_),
    .A(_0457_),
    .B(_0307_));
 sg13g2_nand2b_1 _2062_ (.Y(_0310_),
    .B(_0309_),
    .A_N(_0308_));
 sg13g2_o21ai_1 _2063_ (.B1(_0303_),
    .Y(_0311_),
    .A1(_0299_),
    .A2(_0304_));
 sg13g2_xnor2_1 _2064_ (.Y(_0312_),
    .A(_0310_),
    .B(_0311_));
 sg13g2_nor2_1 _2065_ (.A(net164),
    .B(_0312_),
    .Y(_0313_));
 sg13g2_a21oi_1 _2066_ (.A1(_0457_),
    .A2(net164),
    .Y(_0159_),
    .B1(_0313_));
 sg13g2_o21ai_1 _2067_ (.B1(_0301_),
    .Y(_0314_),
    .A1(_0252_),
    .A2(_0266_));
 sg13g2_nor3_2 _2068_ (.A(_0009_),
    .B(_0008_),
    .C(_0214_),
    .Y(_0315_));
 sg13g2_a22oi_1 _2069_ (.Y(_0316_),
    .B1(_0315_),
    .B2(_0253_),
    .A2(_0314_),
    .A1(_0260_));
 sg13g2_nand2b_1 _2070_ (.Y(_0317_),
    .B(\Voice1.accumulator[7] ),
    .A_N(_0316_));
 sg13g2_nor2b_1 _2071_ (.A(\Voice1.accumulator[7] ),
    .B_N(_0316_),
    .Y(_0318_));
 sg13g2_xnor2_1 _2072_ (.Y(_0319_),
    .A(net383),
    .B(_0316_));
 sg13g2_a21oi_1 _2073_ (.A1(_0309_),
    .A2(_0311_),
    .Y(_0320_),
    .B1(_0308_));
 sg13g2_nand2b_1 _2074_ (.Y(_0321_),
    .B(_0319_),
    .A_N(_0320_));
 sg13g2_nor2b_1 _2075_ (.A(_0319_),
    .B_N(_0320_),
    .Y(_0322_));
 sg13g2_nor2_1 _2076_ (.A(net164),
    .B(_0322_),
    .Y(_0323_));
 sg13g2_a22oi_1 _2077_ (.Y(_0324_),
    .B1(_0321_),
    .B2(_0323_),
    .A2(net164),
    .A1(net383));
 sg13g2_inv_1 _2078_ (.Y(_0160_),
    .A(_0324_));
 sg13g2_nand3_1 _2079_ (.B(\Voice1.accumulator[8] ),
    .C(_0300_),
    .A(net172),
    .Y(_0325_));
 sg13g2_a21o_1 _2080_ (.A2(_0300_),
    .A1(net172),
    .B1(\Voice1.accumulator[8] ),
    .X(_0326_));
 sg13g2_nand2_1 _2081_ (.Y(_0327_),
    .A(_0325_),
    .B(_0326_));
 sg13g2_o21ai_1 _2082_ (.B1(_0317_),
    .Y(_0328_),
    .A1(_0318_),
    .A2(_0320_));
 sg13g2_nand2b_1 _2083_ (.Y(_0329_),
    .B(_0328_),
    .A_N(_0327_));
 sg13g2_nand2b_1 _2084_ (.Y(_0330_),
    .B(_0327_),
    .A_N(_0328_));
 sg13g2_a21oi_1 _2085_ (.A1(_0329_),
    .A2(_0330_),
    .Y(_0331_),
    .B1(_0248_));
 sg13g2_a21oi_1 _2086_ (.A1(_0458_),
    .A2(net164),
    .Y(_0161_),
    .B1(_0331_));
 sg13g2_nor2_1 _2087_ (.A(net379),
    .B(net161),
    .Y(_0332_));
 sg13g2_and3_1 _2088_ (.X(_0333_),
    .A(\Voice1.en ),
    .B(\Voice1.accumulator[9] ),
    .C(_0255_));
 sg13g2_nand3_1 _2089_ (.B(\Voice1.accumulator[9] ),
    .C(_0255_),
    .A(net172),
    .Y(_0334_));
 sg13g2_a21oi_1 _2090_ (.A1(net172),
    .A2(_0255_),
    .Y(_0335_),
    .B1(\Voice1.accumulator[9] ));
 sg13g2_nor2_1 _2091_ (.A(_0333_),
    .B(_0335_),
    .Y(_0336_));
 sg13g2_nand2_1 _2092_ (.Y(_0337_),
    .A(_0325_),
    .B(_0329_));
 sg13g2_xnor2_1 _2093_ (.Y(_0338_),
    .A(_0336_),
    .B(_0337_));
 sg13g2_a21oi_1 _2094_ (.A1(net161),
    .A2(_0338_),
    .Y(_0162_),
    .B1(_0332_));
 sg13g2_o21ai_1 _2095_ (.B1(_0301_),
    .Y(_0339_),
    .A1(_0258_),
    .A2(_0265_));
 sg13g2_nand3_1 _2096_ (.B(_0268_),
    .C(_0339_),
    .A(net172),
    .Y(_0340_));
 sg13g2_nor2_1 _2097_ (.A(_0459_),
    .B(_0340_),
    .Y(_0341_));
 sg13g2_xnor2_1 _2098_ (.Y(_0342_),
    .A(_0459_),
    .B(_0340_));
 sg13g2_nand3b_1 _2099_ (.B(_0328_),
    .C(_0336_),
    .Y(_0343_),
    .A_N(_0327_));
 sg13g2_a21o_1 _2100_ (.A2(_0334_),
    .A1(_0325_),
    .B1(_0335_),
    .X(_0344_));
 sg13g2_nand2_1 _2101_ (.Y(_0345_),
    .A(_0343_),
    .B(_0344_));
 sg13g2_a21oi_1 _2102_ (.A1(_0343_),
    .A2(_0344_),
    .Y(_0346_),
    .B1(_0342_));
 sg13g2_xnor2_1 _2103_ (.Y(_0347_),
    .A(_0342_),
    .B(_0345_));
 sg13g2_nor2_1 _2104_ (.A(_0248_),
    .B(_0347_),
    .Y(_0348_));
 sg13g2_a21oi_1 _2105_ (.A1(_0459_),
    .A2(_0248_),
    .Y(_0163_),
    .B1(_0348_));
 sg13g2_nor2_1 _2106_ (.A(net346),
    .B(net161),
    .Y(_0349_));
 sg13g2_or2_1 _2107_ (.X(_0350_),
    .B(_0315_),
    .A(\Voice1.accumulator[11] ));
 sg13g2_nand2_1 _2108_ (.Y(_0351_),
    .A(\Voice1.accumulator[11] ),
    .B(_0315_));
 sg13g2_nand2_1 _2109_ (.Y(_0352_),
    .A(_0350_),
    .B(_0351_));
 sg13g2_nor2_1 _2110_ (.A(_0341_),
    .B(_0346_),
    .Y(_0353_));
 sg13g2_xnor2_1 _2111_ (.Y(_0354_),
    .A(_0352_),
    .B(_0353_));
 sg13g2_a21oi_1 _2112_ (.A1(net161),
    .A2(_0354_),
    .Y(_0164_),
    .B1(_0349_));
 sg13g2_nand2_1 _2113_ (.Y(_0355_),
    .A(_0344_),
    .B(_0351_));
 sg13g2_a21oi_1 _2114_ (.A1(_0341_),
    .A2(_0350_),
    .Y(_0356_),
    .B1(_0355_));
 sg13g2_nand3_1 _2115_ (.B(_0340_),
    .C(_0351_),
    .A(_0459_),
    .Y(_0357_));
 sg13g2_nand2_1 _2116_ (.Y(_0358_),
    .A(_0350_),
    .B(_0357_));
 sg13g2_a21oi_2 _2117_ (.B1(_0358_),
    .Y(_0359_),
    .A2(_0356_),
    .A1(_0343_));
 sg13g2_nand2_1 _2118_ (.Y(_0360_),
    .A(net162),
    .B(_0359_));
 sg13g2_xnor2_1 _2119_ (.Y(_0165_),
    .A(net310),
    .B(_0360_));
 sg13g2_nand2_1 _2120_ (.Y(_0361_),
    .A(_0011_),
    .B(net162));
 sg13g2_a21oi_1 _2121_ (.A1(net310),
    .A2(_0359_),
    .Y(_0362_),
    .B1(_0361_));
 sg13g2_nor2_1 _2122_ (.A(net354),
    .B(net162),
    .Y(_0363_));
 sg13g2_nor3_2 _2123_ (.A(_0428_),
    .B(net417),
    .C(_0360_),
    .Y(_0364_));
 sg13g2_nor3_1 _2124_ (.A(_0362_),
    .B(_0363_),
    .C(_0364_),
    .Y(_0166_));
 sg13g2_xnor2_1 _2125_ (.Y(_0167_),
    .A(_0431_),
    .B(_0364_));
 sg13g2_nor4_1 _2126_ (.A(_0428_),
    .B(_0430_),
    .C(_0431_),
    .D(net417),
    .Y(_0365_));
 sg13g2_and3_2 _2127_ (.X(_0366_),
    .A(net162),
    .B(_0359_),
    .C(_0365_));
 sg13g2_a21oi_1 _2128_ (.A1(\Voice1.accumulator[14] ),
    .A2(_0364_),
    .Y(_0367_),
    .B1(net283));
 sg13g2_nor2_1 _2129_ (.A(_0366_),
    .B(net284),
    .Y(_0168_));
 sg13g2_xnor2_1 _2130_ (.Y(_0169_),
    .A(_0434_),
    .B(_0366_));
 sg13g2_a21oi_1 _2131_ (.A1(\Voice1.accumulator[16] ),
    .A2(_0366_),
    .Y(_0368_),
    .B1(net316));
 sg13g2_nand3_1 _2132_ (.B(net316),
    .C(_0366_),
    .A(\Voice1.accumulator[16] ),
    .Y(_0369_));
 sg13g2_nor2b_1 _2133_ (.A(net317),
    .B_N(_0369_),
    .Y(_0170_));
 sg13g2_or2_1 _2134_ (.X(_0370_),
    .B(_0369_),
    .A(_0433_));
 sg13g2_xnor2_1 _2135_ (.Y(_0171_),
    .A(net251),
    .B(_0369_));
 sg13g2_nor4_2 _2136_ (.A(_0432_),
    .B(_0433_),
    .C(_0434_),
    .Y(_0371_),
    .D(_0435_));
 sg13g2_a22oi_1 _2137_ (.Y(_0172_),
    .B1(_0371_),
    .B2(_0366_),
    .A2(_0370_),
    .A1(_0432_));
 sg13g2_nand3_1 _2138_ (.B(_0366_),
    .C(_0371_),
    .A(net459),
    .Y(_0372_));
 sg13g2_a21o_1 _2139_ (.A2(_0371_),
    .A1(_0366_),
    .B1(net459),
    .X(_0373_));
 sg13g2_and2_1 _2140_ (.A(_0372_),
    .B(_0373_),
    .X(_0173_));
 sg13g2_nand4_1 _2141_ (.B(\Voice1.accumulator[21] ),
    .C(_0366_),
    .A(\Voice1.accumulator[20] ),
    .Y(_0374_),
    .D(_0371_));
 sg13g2_xnor2_1 _2142_ (.Y(_0174_),
    .A(net352),
    .B(_0372_));
 sg13g2_nor3_1 _2143_ (.A(_0436_),
    .B(_0437_),
    .C(_0372_),
    .Y(_0375_));
 sg13g2_xnor2_1 _2144_ (.Y(_0175_),
    .A(net264),
    .B(_0374_));
 sg13g2_xor2_1 _2145_ (.B(_0375_),
    .A(net247),
    .X(_0176_));
 sg13g2_nor3_1 _2146_ (.A(net179),
    .B(net181),
    .C(net175),
    .Y(_0376_));
 sg13g2_nor2_1 _2147_ (.A(net176),
    .B(net178),
    .Y(_0377_));
 sg13g2_nand3_1 _2148_ (.B(\hvsync_gen.vpos[2] ),
    .C(_0377_),
    .A(net183),
    .Y(_0378_));
 sg13g2_nor2_1 _2149_ (.A(net389),
    .B(net395),
    .Y(_0379_));
 sg13g2_nand3_1 _2150_ (.B(_0376_),
    .C(_0379_),
    .A(\hvsync_gen.vpos[9] ),
    .Y(_0380_));
 sg13g2_o21ai_1 _2151_ (.B1(net207),
    .Y(_0381_),
    .A1(_0378_),
    .A2(_0380_));
 sg13g2_or2_2 _2152_ (.X(_0382_),
    .B(_0381_),
    .A(_0519_));
 sg13g2_inv_1 _2153_ (.Y(_0383_),
    .A(_0382_));
 sg13g2_a22oi_1 _2154_ (.Y(_0384_),
    .B1(_0383_),
    .B2(net239),
    .A2(_0520_),
    .A1(\hvsync_gen.vpos[0] ));
 sg13g2_inv_1 _2155_ (.Y(_0177_),
    .A(net240));
 sg13g2_and2_1 _2156_ (.A(net389),
    .B(net395),
    .X(_0385_));
 sg13g2_nor3_1 _2157_ (.A(_0379_),
    .B(_0382_),
    .C(_0385_),
    .Y(_0386_));
 sg13g2_a21o_1 _2158_ (.A2(_0520_),
    .A1(net389),
    .B1(_0386_),
    .X(_0178_));
 sg13g2_a21oi_1 _2159_ (.A1(_0521_),
    .A2(_0385_),
    .Y(_0387_),
    .B1(net356));
 sg13g2_and2_1 _2160_ (.A(net159),
    .B(_0381_),
    .X(_0388_));
 sg13g2_nand2_1 _2161_ (.Y(_0389_),
    .A(net356),
    .B(_0385_));
 sg13g2_inv_1 _2162_ (.Y(_0390_),
    .A(_0389_));
 sg13g2_o21ai_1 _2163_ (.B1(net159),
    .Y(_0391_),
    .A1(_0381_),
    .A2(_0390_));
 sg13g2_nor2b_1 _2164_ (.A(net357),
    .B_N(_0391_),
    .Y(_0179_));
 sg13g2_nor3_1 _2165_ (.A(net183),
    .B(_0382_),
    .C(_0389_),
    .Y(_0392_));
 sg13g2_a21o_1 _2166_ (.A2(_0391_),
    .A1(net183),
    .B1(_0392_),
    .X(_0180_));
 sg13g2_nand2_1 _2167_ (.Y(_0393_),
    .A(net183),
    .B(_0390_));
 sg13g2_nor2_1 _2168_ (.A(_0520_),
    .B(_0393_),
    .Y(_0394_));
 sg13g2_nand2_1 _2169_ (.Y(_0395_),
    .A(net181),
    .B(_0394_));
 sg13g2_inv_1 _2170_ (.Y(_0396_),
    .A(_0395_));
 sg13g2_nand2b_1 _2171_ (.Y(_0397_),
    .B(_0395_),
    .A_N(_0388_));
 sg13g2_nor2_1 _2172_ (.A(net181),
    .B(_0394_),
    .Y(_0398_));
 sg13g2_nor2_1 _2173_ (.A(_0397_),
    .B(_0398_),
    .Y(_0181_));
 sg13g2_nand2_1 _2174_ (.Y(_0399_),
    .A(net179),
    .B(_0520_));
 sg13g2_nor2_1 _2175_ (.A(net434),
    .B(_0393_),
    .Y(_0400_));
 sg13g2_xnor2_1 _2176_ (.Y(_0401_),
    .A(net179),
    .B(_0400_));
 sg13g2_o21ai_1 _2177_ (.B1(_0399_),
    .Y(_0182_),
    .A1(_0382_),
    .A2(_0401_));
 sg13g2_nand2_1 _2178_ (.Y(_0402_),
    .A(net179),
    .B(net181));
 sg13g2_a21oi_1 _2179_ (.A1(net179),
    .A2(_0396_),
    .Y(_0403_),
    .B1(net178));
 sg13g2_and3_1 _2180_ (.X(_0404_),
    .A(net178),
    .B(net180),
    .C(_0396_));
 sg13g2_nor3_1 _2181_ (.A(_0388_),
    .B(_0403_),
    .C(_0404_),
    .Y(_0183_));
 sg13g2_nand2_1 _2182_ (.Y(_0405_),
    .A(net177),
    .B(_0520_));
 sg13g2_nor3_1 _2183_ (.A(net443),
    .B(_0393_),
    .C(_0402_),
    .Y(_0406_));
 sg13g2_xnor2_1 _2184_ (.Y(_0407_),
    .A(net177),
    .B(_0406_));
 sg13g2_o21ai_1 _2185_ (.B1(_0405_),
    .Y(_0184_),
    .A1(_0382_),
    .A2(net444));
 sg13g2_nand2b_1 _2186_ (.Y(_0408_),
    .B(_0465_),
    .A_N(_0381_));
 sg13g2_nand2_1 _2187_ (.Y(_0409_),
    .A(_0397_),
    .B(_0408_));
 sg13g2_a21oi_1 _2188_ (.A1(net176),
    .A2(_0404_),
    .Y(_0410_),
    .B1(net175));
 sg13g2_a21oi_1 _2189_ (.A1(_0397_),
    .A2(_0408_),
    .Y(_0185_),
    .B1(_0410_));
 sg13g2_nor4_1 _2190_ (.A(net199),
    .B(net446),
    .C(_0465_),
    .D(_0395_),
    .Y(_0411_));
 sg13g2_a21o_1 _2191_ (.A2(_0409_),
    .A1(net446),
    .B1(_0411_),
    .X(_0186_));
 sg13g2_dfrbp_1 _2192_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net221),
    .D(_0021_),
    .Q_N(_0020_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 _2193_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net216),
    .D(net270),
    .Q_N(_1090_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 _2194_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net215),
    .D(net314),
    .Q_N(_0005_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 _2195_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net214),
    .D(_0024_),
    .Q_N(_1089_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 _2196_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net213),
    .D(_0025_),
    .Q_N(_0004_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 _2197_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net212),
    .D(_0026_),
    .Q_N(_1088_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 _2198_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net211),
    .D(_0027_),
    .Q_N(_0003_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 _2199_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net210),
    .D(_0028_),
    .Q_N(_1087_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 _2200_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net209),
    .D(_0029_),
    .Q_N(_1086_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 _2201_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net158),
    .D(net465),
    .Q_N(_0006_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _2202_ (.CLK(net173),
    .RESET_B(net157),
    .D(_0031_),
    .Q_N(_0019_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _2203_ (.CLK(net174),
    .RESET_B(net156),
    .D(_0032_),
    .Q_N(_1085_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _2204_ (.CLK(net174),
    .RESET_B(net155),
    .D(_0033_),
    .Q_N(_1084_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _2205_ (.CLK(net173),
    .RESET_B(net154),
    .D(_0034_),
    .Q_N(_1083_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _2206_ (.CLK(net173),
    .RESET_B(net153),
    .D(_0035_),
    .Q_N(_1082_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _2207_ (.CLK(net173),
    .RESET_B(net152),
    .D(_0036_),
    .Q_N(_1081_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _2208_ (.CLK(net173),
    .RESET_B(net151),
    .D(_0037_),
    .Q_N(_1080_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _2209_ (.CLK(net173),
    .RESET_B(net150),
    .D(_0038_),
    .Q_N(_1079_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 _2210_ (.CLK(net173),
    .RESET_B(net149),
    .D(_0039_),
    .Q_N(_1078_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 _2211_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net148),
    .D(_0040_),
    .Q_N(_1077_),
    .Q(\VAL[0] ));
 sg13g2_dfrbp_1 _2212_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net147),
    .D(_0041_),
    .Q_N(_1076_),
    .Q(\VAL[1] ));
 sg13g2_dfrbp_1 _2213_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net146),
    .D(_0042_),
    .Q_N(_1075_),
    .Q(\VAL[2] ));
 sg13g2_dfrbp_1 _2214_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net145),
    .D(_0043_),
    .Q_N(_1074_),
    .Q(\VAL[3] ));
 sg13g2_dfrbp_1 _2215_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net144),
    .D(_0044_),
    .Q_N(_1073_),
    .Q(\VAL[4] ));
 sg13g2_dfrbp_1 _2216_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net143),
    .D(_0045_),
    .Q_N(_0012_),
    .Q(\VAL[5] ));
 sg13g2_dfrbp_1 _2217_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net142),
    .D(_0046_),
    .Q_N(_1072_),
    .Q(\VAL[6] ));
 sg13g2_dfrbp_1 _2218_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net141),
    .D(_0047_),
    .Q_N(_1071_),
    .Q(\VAL[7] ));
 sg13g2_dfrbp_1 _2219_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net140),
    .D(net388),
    .Q_N(_1070_),
    .Q(\VAL[8] ));
 sg13g2_dfrbp_1 _2220_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net139),
    .D(_0049_),
    .Q_N(_1069_),
    .Q(\VAL[9] ));
 sg13g2_dfrbp_1 _2221_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net138),
    .D(_0050_),
    .Q_N(_1068_),
    .Q(\VAL[10] ));
 sg13g2_dfrbp_1 _2222_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net137),
    .D(net442),
    .Q_N(_1067_),
    .Q(\VAL[11] ));
 sg13g2_dfrbp_1 _2223_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net136),
    .D(_0052_),
    .Q_N(_1066_),
    .Q(\VAL[12] ));
 sg13g2_dfrbp_1 _2224_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net135),
    .D(net278),
    .Q_N(_0013_),
    .Q(\VAL[13] ));
 sg13g2_dfrbp_1 _2225_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net134),
    .D(_0054_),
    .Q_N(_0007_),
    .Q(\VAL[14] ));
 sg13g2_dfrbp_1 _2226_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net133),
    .D(net362),
    .Q_N(_1065_),
    .Q(\VAL[15] ));
 sg13g2_dfrbp_1 _2227_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net132),
    .D(_0056_),
    .Q_N(_1064_),
    .Q(\VAL[16] ));
 sg13g2_dfrbp_1 _2228_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net131),
    .D(_0057_),
    .Q_N(_1063_),
    .Q(\VAL[17] ));
 sg13g2_dfrbp_1 _2229_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net130),
    .D(_0058_),
    .Q_N(_1062_),
    .Q(\VAL[18] ));
 sg13g2_dfrbp_1 _2230_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net129),
    .D(net449),
    .Q_N(_1061_),
    .Q(\VAL[19] ));
 sg13g2_dfrbp_1 _2231_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net128),
    .D(_0060_),
    .Q_N(_1060_),
    .Q(\VAL[20] ));
 sg13g2_dfrbp_1 _2232_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net127),
    .D(_0061_),
    .Q_N(_1059_),
    .Q(\VAL[21] ));
 sg13g2_dfrbp_1 _2233_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net126),
    .D(net250),
    .Q_N(_1058_),
    .Q(\VAL[22] ));
 sg13g2_dfrbp_1 _2234_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net125),
    .D(net325),
    .Q_N(_1057_),
    .Q(\VAL[23] ));
 sg13g2_dfrbp_1 _2235_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net124),
    .D(_0064_),
    .Q_N(_1056_),
    .Q(\yq[0] ));
 sg13g2_dfrbp_1 _2236_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net122),
    .D(net304),
    .Q_N(_1055_),
    .Q(\yq[1] ));
 sg13g2_dfrbp_1 _2237_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net120),
    .D(_0066_),
    .Q_N(_1054_),
    .Q(\yq[2] ));
 sg13g2_dfrbp_1 _2238_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net118),
    .D(_0067_),
    .Q_N(_1053_),
    .Q(\yq[3] ));
 sg13g2_dfrbp_1 _2239_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net116),
    .D(_0068_),
    .Q_N(_1052_),
    .Q(\yq[4] ));
 sg13g2_dfrbp_1 _2240_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net114),
    .D(_0069_),
    .Q_N(_1051_),
    .Q(\yq[5] ));
 sg13g2_dfrbp_1 _2241_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net112),
    .D(_0070_),
    .Q_N(_1050_),
    .Q(\yq[6] ));
 sg13g2_dfrbp_1 _2242_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net110),
    .D(_0071_),
    .Q_N(_1049_),
    .Q(\yq[7] ));
 sg13g2_dfrbp_1 _2243_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net108),
    .D(_0072_),
    .Q_N(_1048_),
    .Q(\yq[8] ));
 sg13g2_dfrbp_1 _2244_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net106),
    .D(_0073_),
    .Q_N(_1047_),
    .Q(\yq[9] ));
 sg13g2_dfrbp_1 _2245_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net104),
    .D(_0074_),
    .Q_N(_1046_),
    .Q(\yq[10] ));
 sg13g2_dfrbp_1 _2246_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net102),
    .D(_0075_),
    .Q_N(_1045_),
    .Q(\yq[11] ));
 sg13g2_dfrbp_1 _2247_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net100),
    .D(_0076_),
    .Q_N(_1044_),
    .Q(\yq[12] ));
 sg13g2_dfrbp_1 _2248_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net98),
    .D(net301),
    .Q_N(_1043_),
    .Q(\yqo[0] ));
 sg13g2_dfrbp_1 _2249_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net96),
    .D(_0078_),
    .Q_N(_1042_),
    .Q(\yqo[1] ));
 sg13g2_dfrbp_1 _2250_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net94),
    .D(_0079_),
    .Q_N(_1041_),
    .Q(\yqo[2] ));
 sg13g2_dfrbp_1 _2251_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net92),
    .D(net336),
    .Q_N(_1040_),
    .Q(\yqo[3] ));
 sg13g2_dfrbp_1 _2252_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net90),
    .D(net298),
    .Q_N(_1039_),
    .Q(\yqo[4] ));
 sg13g2_dfrbp_1 _2253_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net88),
    .D(net399),
    .Q_N(_0002_),
    .Q(\yqo[5] ));
 sg13g2_dfrbp_1 _2254_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net86),
    .D(net416),
    .Q_N(_1038_),
    .Q(\yqo[6] ));
 sg13g2_dfrbp_1 _2255_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net84),
    .D(_0084_),
    .Q_N(_1037_),
    .Q(\yqo[7] ));
 sg13g2_dfrbp_1 _2256_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net82),
    .D(net433),
    .Q_N(_1036_),
    .Q(\yqo[8] ));
 sg13g2_dfrbp_1 _2257_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net80),
    .D(_0086_),
    .Q_N(_1035_),
    .Q(\yqo[9] ));
 sg13g2_dfrbp_1 _2258_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net78),
    .D(_0087_),
    .Q_N(_1034_),
    .Q(\yqo[10] ));
 sg13g2_dfrbp_1 _2259_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net76),
    .D(net404),
    .Q_N(_1033_),
    .Q(\yqo[11] ));
 sg13g2_dfrbp_1 _2260_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net74),
    .D(net333),
    .Q_N(_1032_),
    .Q(\yqo[12] ));
 sg13g2_dfrbp_1 _2261_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net72),
    .D(_0090_),
    .Q_N(_1031_),
    .Q(\LFSR[0] ));
 sg13g2_dfrbp_1 _2262_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net71),
    .D(net267),
    .Q_N(_1030_),
    .Q(\LFSR[1] ));
 sg13g2_dfrbp_1 _2263_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net70),
    .D(net420),
    .Q_N(_1029_),
    .Q(\LFSR[2] ));
 sg13g2_dfrbp_1 _2264_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net69),
    .D(_0093_),
    .Q_N(_1028_),
    .Q(\LFSR[3] ));
 sg13g2_dfrbp_1 _2265_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net68),
    .D(_0094_),
    .Q_N(_1027_),
    .Q(\LFSR[4] ));
 sg13g2_dfrbp_1 _2266_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net67),
    .D(_0095_),
    .Q_N(_1026_),
    .Q(\LFSR[5] ));
 sg13g2_dfrbp_1 _2267_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net66),
    .D(_0096_),
    .Q_N(_1025_),
    .Q(\xq[0] ));
 sg13g2_dfrbp_1 _2268_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net65),
    .D(_0097_),
    .Q_N(_1024_),
    .Q(\xq[1] ));
 sg13g2_dfrbp_1 _2269_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net64),
    .D(_0098_),
    .Q_N(_1023_),
    .Q(\xq[2] ));
 sg13g2_dfrbp_1 _2270_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net63),
    .D(_0099_),
    .Q_N(_1022_),
    .Q(\xq[3] ));
 sg13g2_dfrbp_1 _2271_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net62),
    .D(_0100_),
    .Q_N(_1021_),
    .Q(\xq[4] ));
 sg13g2_dfrbp_1 _2272_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net61),
    .D(_0101_),
    .Q_N(_1020_),
    .Q(\xq[5] ));
 sg13g2_dfrbp_1 _2273_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net60),
    .D(net359),
    .Q_N(_1019_),
    .Q(\xq[6] ));
 sg13g2_dfrbp_1 _2274_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net59),
    .D(_0103_),
    .Q_N(_1018_),
    .Q(\xq[7] ));
 sg13g2_dfrbp_1 _2275_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net58),
    .D(net374),
    .Q_N(_1017_),
    .Q(\xq[8] ));
 sg13g2_dfrbp_1 _2276_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net57),
    .D(_0105_),
    .Q_N(_1016_),
    .Q(\xq[9] ));
 sg13g2_dfrbp_1 _2277_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net56),
    .D(net275),
    .Q_N(_1015_),
    .Q(\xq[10] ));
 sg13g2_dfrbp_1 _2278_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net55),
    .D(net246),
    .Q_N(_1014_),
    .Q(\xq[11] ));
 sg13g2_dfrbp_1 _2279_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net54),
    .D(_0108_),
    .Q_N(_0018_),
    .Q(\ctr_audio[0] ));
 sg13g2_dfrbp_1 _2280_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net52),
    .D(net255),
    .Q_N(_1013_),
    .Q(\ctr_audio[1] ));
 sg13g2_dfrbp_1 _2281_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net50),
    .D(_0110_),
    .Q_N(_1012_),
    .Q(\ctr_audio[2] ));
 sg13g2_dfrbp_1 _2282_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net48),
    .D(net287),
    .Q_N(_1011_),
    .Q(\ctr_audio[3] ));
 sg13g2_dfrbp_1 _2283_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net46),
    .D(net260),
    .Q_N(_1010_),
    .Q(\ctr_audio[4] ));
 sg13g2_dfrbp_1 _2284_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net44),
    .D(_0113_),
    .Q_N(_1009_),
    .Q(\ctr_audio[5] ));
 sg13g2_dfrbp_1 _2285_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net42),
    .D(_0114_),
    .Q_N(_1008_),
    .Q(\ctr_audio[6] ));
 sg13g2_dfrbp_1 _2286_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net40),
    .D(net293),
    .Q_N(_1007_),
    .Q(\ctr_audio[7] ));
 sg13g2_dfrbp_1 _2287_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net38),
    .D(net322),
    .Q_N(_1006_),
    .Q(\ctr_audio[8] ));
 sg13g2_dfrbp_1 _2288_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net36),
    .D(_0117_),
    .Q_N(_1005_),
    .Q(\ctr_audio[9] ));
 sg13g2_dfrbp_1 _2289_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net34),
    .D(_0118_),
    .Q_N(_1004_),
    .Q(\Voice1.pulsewidth[0] ));
 sg13g2_dfrbp_1 _2290_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net32),
    .D(net343),
    .Q_N(_1003_),
    .Q(\Voice1.pulsewidth[1] ));
 sg13g2_dfrbp_1 _2291_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net30),
    .D(_0120_),
    .Q_N(_1002_),
    .Q(\Voice1.pulsewidth[2] ));
 sg13g2_dfrbp_1 _2292_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net28),
    .D(net468),
    .Q_N(_1001_),
    .Q(\Voice1.pulsewidth[3] ));
 sg13g2_dfrbp_1 _2293_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net26),
    .D(net371),
    .Q_N(_1000_),
    .Q(\Voice1.pulsewidth[4] ));
 sg13g2_dfrbp_1 _2294_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net24),
    .D(_0123_),
    .Q_N(_0999_),
    .Q(\Voice1.pulsewidth[5] ));
 sg13g2_dfrbp_1 _2295_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net22),
    .D(_0124_),
    .Q_N(_0998_),
    .Q(\Voice1.pulsewidth[6] ));
 sg13g2_dfrbp_1 _2296_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net20),
    .D(_0125_),
    .Q_N(_0997_),
    .Q(\Voice1.pulsewidth[7] ));
 sg13g2_dfrbp_1 _2297_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net18),
    .D(_0126_),
    .Q_N(_0996_),
    .Q(\Voice1.pulsewidth[8] ));
 sg13g2_dfrbp_1 _2298_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net16),
    .D(_0127_),
    .Q_N(_0995_),
    .Q(\ctr_audio[19] ));
 sg13g2_dfrbp_1 _2299_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net233),
    .D(_0128_),
    .Q_N(_0994_),
    .Q(\ctr_audio[20] ));
 sg13g2_dfrbp_1 _2300_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net230),
    .D(_0129_),
    .Q_N(_0993_),
    .Q(\ctr_audio[21] ));
 sg13g2_dfrbp_1 _2301_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net228),
    .D(net463),
    .Q_N(_0992_),
    .Q(\ctr_audio[22] ));
 sg13g2_dfrbp_1 _2302_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net226),
    .D(net378),
    .Q_N(_0009_),
    .Q(\Voice1.pulsewidth[10] ));
 sg13g2_dfrbp_1 _2303_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net224),
    .D(_0132_),
    .Q_N(_0991_),
    .Q(\xqo[0] ));
 sg13g2_dfrbp_1 _2304_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net223),
    .D(_0133_),
    .Q_N(_0990_),
    .Q(\xqo[1] ));
 sg13g2_dfrbp_1 _2305_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net222),
    .D(_0134_),
    .Q_N(_0989_),
    .Q(\xqo[2] ));
 sg13g2_dfrbp_1 _2306_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net220),
    .D(_0135_),
    .Q_N(_0988_),
    .Q(\xqo[3] ));
 sg13g2_dfrbp_1 _2307_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net219),
    .D(_0136_),
    .Q_N(_0987_),
    .Q(\xqo[4] ));
 sg13g2_dfrbp_1 _2308_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net218),
    .D(_0137_),
    .Q_N(_0986_),
    .Q(\xqo[5] ));
 sg13g2_dfrbp_1 _2309_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net217),
    .D(_0138_),
    .Q_N(_0985_),
    .Q(\xqo[6] ));
 sg13g2_dfrbp_1 _2310_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net123),
    .D(_0139_),
    .Q_N(_0984_),
    .Q(\xqo[7] ));
 sg13g2_dfrbp_1 _2311_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net121),
    .D(_0140_),
    .Q_N(_0983_),
    .Q(\xqo[8] ));
 sg13g2_dfrbp_1 _2312_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net119),
    .D(_0141_),
    .Q_N(_0982_),
    .Q(\xqo[9] ));
 sg13g2_dfrbp_1 _2313_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net117),
    .D(_0142_),
    .Q_N(_0981_),
    .Q(\xqo[10] ));
 sg13g2_dfrbp_1 _2314_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net115),
    .D(_0143_),
    .Q_N(_0980_),
    .Q(\xqo[11] ));
 sg13g2_dfrbp_1 _2315_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net113),
    .D(_0144_),
    .Q_N(_0017_),
    .Q(\ctr_clkdiv25[0] ));
 sg13g2_dfrbp_1 _2316_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net111),
    .D(_0145_),
    .Q_N(_0979_),
    .Q(\ctr_clkdiv25[1] ));
 sg13g2_dfrbp_1 _2317_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net109),
    .D(net263),
    .Q_N(_0978_),
    .Q(\ctr_clkdiv25[2] ));
 sg13g2_dfrbp_1 _2318_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net107),
    .D(_0147_),
    .Q_N(_0977_),
    .Q(\ctr_clkdiv25[3] ));
 sg13g2_dfrbp_1 _2319_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net105),
    .D(net328),
    .Q_N(_0976_),
    .Q(\ctr_clkdiv25[4] ));
 sg13g2_dfrbp_1 _2320_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net103),
    .D(_0149_),
    .Q_N(_0975_),
    .Q(\ctr_clkdiv25[5] ));
 sg13g2_dfrbp_1 _2321_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net101),
    .D(_0150_),
    .Q_N(_0974_),
    .Q(\ctr_clkdiv25[6] ));
 sg13g2_dfrbp_1 _2322_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net99),
    .D(_0151_),
    .Q_N(_0973_),
    .Q(\ctr_clkdiv25[7] ));
 sg13g2_dfrbp_1 _2323_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net97),
    .D(net365),
    .Q_N(_0972_),
    .Q(\Voice1.pulse ));
 sg13g2_dfrbp_1 _2324_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net93),
    .D(net272),
    .Q_N(_0010_),
    .Q(\Voice1.accumulator[0] ));
 sg13g2_dfrbp_1 _2325_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net91),
    .D(net349),
    .Q_N(_0971_),
    .Q(\Voice1.accumulator[1] ));
 sg13g2_dfrbp_1 _2326_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net89),
    .D(_0155_),
    .Q_N(_0970_),
    .Q(\Voice1.accumulator[2] ));
 sg13g2_dfrbp_1 _2327_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net87),
    .D(net351),
    .Q_N(_0969_),
    .Q(\Voice1.accumulator[3] ));
 sg13g2_dfrbp_1 _2328_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net85),
    .D(_0157_),
    .Q_N(_0968_),
    .Q(\Voice1.accumulator[4] ));
 sg13g2_dfrbp_1 _2329_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net83),
    .D(_0158_),
    .Q_N(_0967_),
    .Q(\Voice1.accumulator[5] ));
 sg13g2_dfrbp_1 _2330_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net81),
    .D(_0159_),
    .Q_N(_0966_),
    .Q(\Voice1.accumulator[6] ));
 sg13g2_dfrbp_1 _2331_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net79),
    .D(_0160_),
    .Q_N(_0965_),
    .Q(\Voice1.accumulator[7] ));
 sg13g2_dfrbp_1 _2332_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net77),
    .D(_0161_),
    .Q_N(_0964_),
    .Q(\Voice1.accumulator[8] ));
 sg13g2_dfrbp_1 _2333_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net75),
    .D(_0162_),
    .Q_N(_0963_),
    .Q(\Voice1.accumulator[9] ));
 sg13g2_dfrbp_1 _2334_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net73),
    .D(net411),
    .Q_N(_0962_),
    .Q(\Voice1.accumulator[10] ));
 sg13g2_dfrbp_1 _2335_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net53),
    .D(net347),
    .Q_N(_0961_),
    .Q(\Voice1.accumulator[11] ));
 sg13g2_dfrbp_1 _2336_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net51),
    .D(_0165_),
    .Q_N(_0960_),
    .Q(\Voice1.accumulator[12] ));
 sg13g2_dfrbp_1 _2337_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net49),
    .D(net355),
    .Q_N(_0011_),
    .Q(\Voice1.accumulator[13] ));
 sg13g2_dfrbp_1 _2338_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net47),
    .D(net418),
    .Q_N(_0959_),
    .Q(\Voice1.accumulator[14] ));
 sg13g2_dfrbp_1 _2339_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net45),
    .D(net285),
    .Q_N(_0958_),
    .Q(\Voice1.accumulator[15] ));
 sg13g2_dfrbp_1 _2340_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net43),
    .D(_0169_),
    .Q_N(_0957_),
    .Q(\Voice1.accumulator[16] ));
 sg13g2_dfrbp_1 _2341_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net41),
    .D(net318),
    .Q_N(_0956_),
    .Q(\Voice1.accumulator[17] ));
 sg13g2_dfrbp_1 _2342_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net39),
    .D(net252),
    .Q_N(_0955_),
    .Q(\Voice1.accumulator[18] ));
 sg13g2_dfrbp_1 _2343_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net37),
    .D(net428),
    .Q_N(_0954_),
    .Q(\Voice1.accumulator[19] ));
 sg13g2_dfrbp_1 _2344_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net35),
    .D(_0173_),
    .Q_N(_0953_),
    .Q(\Voice1.accumulator[20] ));
 sg13g2_dfrbp_1 _2345_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net33),
    .D(net353),
    .Q_N(_0952_),
    .Q(\Voice1.accumulator[21] ));
 sg13g2_dfrbp_1 _2346_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net31),
    .D(net265),
    .Q_N(_0951_),
    .Q(\Voice1.accumulator[22] ));
 sg13g2_dfrbp_1 _2347_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net232),
    .D(net248),
    .Q_N(_1091_),
    .Q(\Voice1.accumulator[23] ));
 sg13g2_dfrbp_1 _2348_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net29),
    .D(net281),
    .Q_N(_0950_),
    .Q(hsync));
 sg13g2_dfrbp_1 _2349_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net27),
    .D(_0177_),
    .Q_N(_0016_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _2350_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net23),
    .D(_0178_),
    .Q_N(_0949_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _2351_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net19),
    .D(_0179_),
    .Q_N(_0948_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _2352_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net15),
    .D(_0180_),
    .Q_N(_0947_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _2353_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net229),
    .D(_0181_),
    .Q_N(_0014_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _2354_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net225),
    .D(_0182_),
    .Q_N(_0946_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _2355_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net25),
    .D(_0183_),
    .Q_N(_0015_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _2356_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net17),
    .D(net445),
    .Q_N(_0945_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _2357_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net227),
    .D(_0185_),
    .Q_N(_0944_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _2358_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net231),
    .D(_0186_),
    .Q_N(_1092_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _2359_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net21),
    .D(net391),
    .Q_N(_0943_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 _2360_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net95),
    .D(_0187_),
    .Q_N(_0008_),
    .Q(\Voice1.en ));
 sg13g2_tiehi _2298__16 (.L_HI(net16));
 sg13g2_tiehi _2356__17 (.L_HI(net17));
 sg13g2_tiehi _2297__18 (.L_HI(net18));
 sg13g2_tiehi _2351__19 (.L_HI(net19));
 sg13g2_tiehi _2296__20 (.L_HI(net20));
 sg13g2_tiehi _2359__21 (.L_HI(net21));
 sg13g2_tiehi _2295__22 (.L_HI(net22));
 sg13g2_tiehi _2350__23 (.L_HI(net23));
 sg13g2_tiehi _2294__24 (.L_HI(net24));
 sg13g2_tiehi _2355__25 (.L_HI(net25));
 sg13g2_tiehi _2293__26 (.L_HI(net26));
 sg13g2_tiehi _2349__27 (.L_HI(net27));
 sg13g2_tiehi _2292__28 (.L_HI(net28));
 sg13g2_tiehi _2348__29 (.L_HI(net29));
 sg13g2_tiehi _2291__30 (.L_HI(net30));
 sg13g2_tiehi _2346__31 (.L_HI(net31));
 sg13g2_tiehi _2290__32 (.L_HI(net32));
 sg13g2_tiehi _2345__33 (.L_HI(net33));
 sg13g2_tiehi _2289__34 (.L_HI(net34));
 sg13g2_tiehi _2344__35 (.L_HI(net35));
 sg13g2_tiehi _2288__36 (.L_HI(net36));
 sg13g2_tiehi _2343__37 (.L_HI(net37));
 sg13g2_tiehi _2287__38 (.L_HI(net38));
 sg13g2_tiehi _2342__39 (.L_HI(net39));
 sg13g2_tiehi _2286__40 (.L_HI(net40));
 sg13g2_tiehi _2341__41 (.L_HI(net41));
 sg13g2_tiehi _2285__42 (.L_HI(net42));
 sg13g2_tiehi _2340__43 (.L_HI(net43));
 sg13g2_tiehi _2284__44 (.L_HI(net44));
 sg13g2_tiehi _2339__45 (.L_HI(net45));
 sg13g2_tiehi _2283__46 (.L_HI(net46));
 sg13g2_tiehi _2338__47 (.L_HI(net47));
 sg13g2_tiehi _2282__48 (.L_HI(net48));
 sg13g2_tiehi _2337__49 (.L_HI(net49));
 sg13g2_tiehi _2281__50 (.L_HI(net50));
 sg13g2_tiehi _2336__51 (.L_HI(net51));
 sg13g2_tiehi _2280__52 (.L_HI(net52));
 sg13g2_tiehi _2335__53 (.L_HI(net53));
 sg13g2_tiehi _2279__54 (.L_HI(net54));
 sg13g2_tiehi _2278__55 (.L_HI(net55));
 sg13g2_tiehi _2277__56 (.L_HI(net56));
 sg13g2_tiehi _2276__57 (.L_HI(net57));
 sg13g2_tiehi _2275__58 (.L_HI(net58));
 sg13g2_tiehi _2274__59 (.L_HI(net59));
 sg13g2_tiehi _2273__60 (.L_HI(net60));
 sg13g2_tiehi _2272__61 (.L_HI(net61));
 sg13g2_tiehi _2271__62 (.L_HI(net62));
 sg13g2_tiehi _2270__63 (.L_HI(net63));
 sg13g2_tiehi _2269__64 (.L_HI(net64));
 sg13g2_tiehi _2268__65 (.L_HI(net65));
 sg13g2_tiehi _2267__66 (.L_HI(net66));
 sg13g2_tiehi _2266__67 (.L_HI(net67));
 sg13g2_tiehi _2265__68 (.L_HI(net68));
 sg13g2_tiehi _2264__69 (.L_HI(net69));
 sg13g2_tiehi _2263__70 (.L_HI(net70));
 sg13g2_tiehi _2262__71 (.L_HI(net71));
 sg13g2_tiehi _2261__72 (.L_HI(net72));
 sg13g2_tiehi _2334__73 (.L_HI(net73));
 sg13g2_tiehi _2260__74 (.L_HI(net74));
 sg13g2_tiehi _2333__75 (.L_HI(net75));
 sg13g2_tiehi _2259__76 (.L_HI(net76));
 sg13g2_tiehi _2332__77 (.L_HI(net77));
 sg13g2_tiehi _2258__78 (.L_HI(net78));
 sg13g2_tiehi _2331__79 (.L_HI(net79));
 sg13g2_tiehi _2257__80 (.L_HI(net80));
 sg13g2_tiehi _2330__81 (.L_HI(net81));
 sg13g2_tiehi _2256__82 (.L_HI(net82));
 sg13g2_tiehi _2329__83 (.L_HI(net83));
 sg13g2_tiehi _2255__84 (.L_HI(net84));
 sg13g2_tiehi _2328__85 (.L_HI(net85));
 sg13g2_tiehi _2254__86 (.L_HI(net86));
 sg13g2_tiehi _2327__87 (.L_HI(net87));
 sg13g2_tiehi _2253__88 (.L_HI(net88));
 sg13g2_tiehi _2326__89 (.L_HI(net89));
 sg13g2_tiehi _2252__90 (.L_HI(net90));
 sg13g2_tiehi _2325__91 (.L_HI(net91));
 sg13g2_tiehi _2251__92 (.L_HI(net92));
 sg13g2_tiehi _2324__93 (.L_HI(net93));
 sg13g2_tiehi _2250__94 (.L_HI(net94));
 sg13g2_tiehi _2360__95 (.L_HI(net95));
 sg13g2_tiehi _2249__96 (.L_HI(net96));
 sg13g2_tiehi _2323__97 (.L_HI(net97));
 sg13g2_tiehi _2248__98 (.L_HI(net98));
 sg13g2_tiehi _2322__99 (.L_HI(net99));
 sg13g2_tiehi _2247__100 (.L_HI(net100));
 sg13g2_tiehi _2321__101 (.L_HI(net101));
 sg13g2_tiehi _2246__102 (.L_HI(net102));
 sg13g2_tiehi _2320__103 (.L_HI(net103));
 sg13g2_tiehi _2245__104 (.L_HI(net104));
 sg13g2_tiehi _2319__105 (.L_HI(net105));
 sg13g2_tiehi _2244__106 (.L_HI(net106));
 sg13g2_tiehi _2318__107 (.L_HI(net107));
 sg13g2_tiehi _2243__108 (.L_HI(net108));
 sg13g2_tiehi _2317__109 (.L_HI(net109));
 sg13g2_tiehi _2242__110 (.L_HI(net110));
 sg13g2_tiehi _2316__111 (.L_HI(net111));
 sg13g2_tiehi _2241__112 (.L_HI(net112));
 sg13g2_tiehi _2315__113 (.L_HI(net113));
 sg13g2_tiehi _2240__114 (.L_HI(net114));
 sg13g2_tiehi _2314__115 (.L_HI(net115));
 sg13g2_tiehi _2239__116 (.L_HI(net116));
 sg13g2_tiehi _2313__117 (.L_HI(net117));
 sg13g2_tiehi _2238__118 (.L_HI(net118));
 sg13g2_tiehi _2312__119 (.L_HI(net119));
 sg13g2_tiehi _2237__120 (.L_HI(net120));
 sg13g2_tiehi _2311__121 (.L_HI(net121));
 sg13g2_tiehi _2236__122 (.L_HI(net122));
 sg13g2_tiehi _2310__123 (.L_HI(net123));
 sg13g2_tiehi _2235__124 (.L_HI(net124));
 sg13g2_tiehi _2234__125 (.L_HI(net125));
 sg13g2_tiehi _2233__126 (.L_HI(net126));
 sg13g2_tiehi _2232__127 (.L_HI(net127));
 sg13g2_tiehi _2231__128 (.L_HI(net128));
 sg13g2_tiehi _2230__129 (.L_HI(net129));
 sg13g2_tiehi _2229__130 (.L_HI(net130));
 sg13g2_tiehi _2228__131 (.L_HI(net131));
 sg13g2_tiehi _2227__132 (.L_HI(net132));
 sg13g2_tiehi _2226__133 (.L_HI(net133));
 sg13g2_tiehi _2225__134 (.L_HI(net134));
 sg13g2_tiehi _2224__135 (.L_HI(net135));
 sg13g2_tiehi _2223__136 (.L_HI(net136));
 sg13g2_tiehi _2222__137 (.L_HI(net137));
 sg13g2_tiehi _2221__138 (.L_HI(net138));
 sg13g2_tiehi _2220__139 (.L_HI(net139));
 sg13g2_tiehi _2219__140 (.L_HI(net140));
 sg13g2_tiehi _2218__141 (.L_HI(net141));
 sg13g2_tiehi _2217__142 (.L_HI(net142));
 sg13g2_tiehi _2216__143 (.L_HI(net143));
 sg13g2_tiehi _2215__144 (.L_HI(net144));
 sg13g2_tiehi _2214__145 (.L_HI(net145));
 sg13g2_tiehi _2213__146 (.L_HI(net146));
 sg13g2_tiehi _2212__147 (.L_HI(net147));
 sg13g2_tiehi _2211__148 (.L_HI(net148));
 sg13g2_tiehi _2210__149 (.L_HI(net149));
 sg13g2_tiehi _2209__150 (.L_HI(net150));
 sg13g2_tiehi _2208__151 (.L_HI(net151));
 sg13g2_tiehi _2207__152 (.L_HI(net152));
 sg13g2_tiehi _2206__153 (.L_HI(net153));
 sg13g2_tiehi _2205__154 (.L_HI(net154));
 sg13g2_tiehi _2204__155 (.L_HI(net155));
 sg13g2_tiehi _2203__156 (.L_HI(net156));
 sg13g2_tiehi _2202__157 (.L_HI(net157));
 sg13g2_tiehi _2201__158 (.L_HI(net158));
 sg13g2_tiehi _2200__159 (.L_HI(net209));
 sg13g2_tiehi _2199__160 (.L_HI(net210));
 sg13g2_tiehi _2198__161 (.L_HI(net211));
 sg13g2_tiehi _2197__162 (.L_HI(net212));
 sg13g2_tiehi _2196__163 (.L_HI(net213));
 sg13g2_tiehi _2195__164 (.L_HI(net214));
 sg13g2_tiehi _2194__165 (.L_HI(net215));
 sg13g2_tiehi _2193__166 (.L_HI(net216));
 sg13g2_tiehi _2309__167 (.L_HI(net217));
 sg13g2_tiehi _2308__168 (.L_HI(net218));
 sg13g2_tiehi _2307__169 (.L_HI(net219));
 sg13g2_tiehi _2306__170 (.L_HI(net220));
 sg13g2_tiehi _2192__171 (.L_HI(net221));
 sg13g2_tiehi _2305__172 (.L_HI(net222));
 sg13g2_tiehi _2304__173 (.L_HI(net223));
 sg13g2_tiehi _2303__174 (.L_HI(net224));
 sg13g2_tiehi _2354__175 (.L_HI(net225));
 sg13g2_tiehi _2302__176 (.L_HI(net226));
 sg13g2_tiehi _2357__177 (.L_HI(net227));
 sg13g2_tiehi _2301__178 (.L_HI(net228));
 sg13g2_tiehi _2353__179 (.L_HI(net229));
 sg13g2_tiehi _2300__180 (.L_HI(net230));
 sg13g2_tiehi _2358__181 (.L_HI(net231));
 sg13g2_tiehi _2347__182 (.L_HI(net232));
 sg13g2_tiehi _2299__183 (.L_HI(net233));
 sg13g2_tiehi tt_um_top_184 (.L_HI(net234));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_top_2 (.L_LO(net2));
 sg13g2_tielo tt_um_top_3 (.L_LO(net3));
 sg13g2_tielo tt_um_top_4 (.L_LO(net4));
 sg13g2_tielo tt_um_top_5 (.L_LO(net5));
 sg13g2_tielo tt_um_top_6 (.L_LO(net6));
 sg13g2_tielo tt_um_top_7 (.L_LO(net7));
 sg13g2_tielo tt_um_top_8 (.L_LO(net8));
 sg13g2_tielo tt_um_top_9 (.L_LO(net9));
 sg13g2_tielo tt_um_top_10 (.L_LO(net10));
 sg13g2_tielo tt_um_top_11 (.L_LO(net11));
 sg13g2_tielo tt_um_top_12 (.L_LO(net12));
 sg13g2_tielo tt_um_top_13 (.L_LO(net13));
 sg13g2_tielo tt_um_top_14 (.L_LO(net14));
 sg13g2_tiehi _2352__15 (.L_HI(net15));
 sg13g2_buf_1 _2545_ (.A(\Voice1.pulse ),
    .X(uio_out[7]));
 sg13g2_buf_2 _2546_ (.A(net174),
    .X(uo_out[3]));
 sg13g2_buf_2 _2547_ (.A(net187),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout159 (.X(net159),
    .A(_0521_));
 sg13g2_buf_2 fanout160 (.A(net162),
    .X(net160));
 sg13g2_buf_1 fanout161 (.A(net162),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_0247_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(\counter[5] ),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_0248_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(net167),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(net167),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(net168),
    .X(net167));
 sg13g2_buf_4 fanout168 (.X(net168),
    .A(_0722_));
 sg13g2_buf_2 fanout169 (.A(_0447_),
    .X(net169));
 sg13g2_buf_4 fanout170 (.X(net170),
    .A(net171));
 sg13g2_buf_4 fanout171 (.X(net171),
    .A(_0423_));
 sg13g2_buf_2 fanout172 (.A(\Voice1.en ),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(net174),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(net453),
    .X(net174));
 sg13g2_buf_4 fanout175 (.X(net175),
    .A(net473));
 sg13g2_buf_2 fanout176 (.A(net177),
    .X(net176));
 sg13g2_buf_4 fanout177 (.X(net177),
    .A(\hvsync_gen.vpos[7] ));
 sg13g2_buf_4 fanout178 (.X(net178),
    .A(net472));
 sg13g2_buf_2 fanout179 (.A(net180),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(\hvsync_gen.vpos[5] ),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(net470),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(\hvsync_gen.vpos[4] ),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(net458),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(net185),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(net186),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(net299),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(net299),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(net435),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(net464),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(\hvsync_gen.hpos[8] ),
    .X(net190));
 sg13g2_buf_1 fanout191 (.A(net460),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(\hvsync_gen.hpos[7] ),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(net478),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(\hvsync_gen.hpos[5] ),
    .X(net194));
 sg13g2_buf_4 fanout195 (.X(net195),
    .A(net475));
 sg13g2_buf_2 fanout196 (.A(net197),
    .X(net196));
 sg13g2_buf_1 fanout197 (.A(net198),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_0438_),
    .X(net198));
 sg13g2_buf_4 fanout199 (.X(net199),
    .A(net200));
 sg13g2_buf_4 fanout200 (.X(net200),
    .A(_0438_));
 sg13g2_buf_2 fanout201 (.A(net203),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(net203),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(net204),
    .X(net203));
 sg13g2_buf_4 fanout204 (.X(net204),
    .A(rst_n));
 sg13g2_buf_2 fanout205 (.A(net206),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(net208),
    .X(net206));
 sg13g2_buf_4 fanout207 (.X(net207),
    .A(net208));
 sg13g2_buf_2 fanout208 (.A(rst_n),
    .X(net208));
 sg13g2_tielo tt_um_top_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0020_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0017_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0018_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0928_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0016_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0384_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold7 (.A(\xq[3] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold8 (.A(\xq[0] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold9 (.A(\xq[1] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold10 (.A(\xq[2] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold11 (.A(\xqo[11] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0107_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold13 (.A(\Voice1.accumulator[23] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0176_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0007_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0062_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold17 (.A(\Voice1.accumulator[18] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0171_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold19 (.A(\ctr_audio[1] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0929_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0109_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold22 (.A(\xq[9] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold23 (.A(\xq[11] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold24 (.A(\ctr_audio[4] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0935_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0112_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold27 (.A(\ctr_clkdiv25[2] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0219_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0146_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold30 (.A(\Voice1.accumulator[22] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0175_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold32 (.A(\LFSR[0] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0091_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold34 (.A(\hvsync_gen.hpos[1] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0522_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0022_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold37 (.A(\Voice1.accumulator[0] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0153_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold39 (.A(\xqo[10] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0920_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0106_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0012_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0693_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0053_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0006_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0472_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0000_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold48 (.A(\xq[8] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold49 (.A(\Voice1.accumulator[15] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0367_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0168_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold52 (.A(\ctr_audio[3] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0111_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold54 (.A(\xq[6] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold55 (.A(\xqo[4] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0909_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold57 (.A(\ctr_audio[7] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0940_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0115_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0004_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0527_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0528_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold63 (.A(\yq[4] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0081_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold65 (.A(hsync),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold66 (.A(\yq[0] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0077_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold68 (.A(\Voice1.accumulator[8] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold69 (.A(\yq[1] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0065_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold71 (.A(\xq[5] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold72 (.A(\yqo[0] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0013_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0717_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold75 (.A(\yq[2] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold76 (.A(\Voice1.accumulator[12] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold77 (.A(\yqo[2] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold78 (.A(\Voice1.accumulator[4] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold79 (.A(\hvsync_gen.hpos[2] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0023_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold81 (.A(\xq[7] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold82 (.A(\Voice1.accumulator[17] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0368_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0170_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold85 (.A(\Voice1.accumulator[2] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold86 (.A(\ctr_audio[8] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0188_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0116_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold89 (.A(\VAL[15] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0719_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0063_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold92 (.A(\ctr_clkdiv25[4] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0223_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0148_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold95 (.A(\ctr_clkdiv25[3] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0221_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold97 (.A(\Voice1.accumulator[6] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold98 (.A(\yqo[12] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0089_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold100 (.A(\Voice1.accumulator[5] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold101 (.A(\yq[3] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0080_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold103 (.A(\xq[10] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0005_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold105 (.A(\yq[12] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold106 (.A(\LFSR[3] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold107 (.A(\Voice1.pulsewidth[1] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0193_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0119_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold110 (.A(\xq[4] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold111 (.A(\yqo[1] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold112 (.A(\Voice1.accumulator[11] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0164_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold114 (.A(\Voice1.accumulator[1] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0154_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold116 (.A(\Voice1.accumulator[3] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0156_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold118 (.A(\Voice1.accumulator[21] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0174_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold120 (.A(\Voice1.accumulator[13] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0166_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold122 (.A(\hvsync_gen.vpos[2] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0387_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold124 (.A(\xqo[6] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0102_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold126 (.A(\ctr_clkdiv25[5] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold127 (.A(\VAL[7] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0055_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold129 (.A(\Voice1.pulse ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0246_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0152_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold132 (.A(\xqo[5] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold133 (.A(\ctr_audio[5] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0938_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold135 (.A(\Voice1.pulsewidth[4] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0199_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0122_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold138 (.A(\xqo[8] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0918_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0104_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold141 (.A(\xqo[9] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0919_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold143 (.A(\Voice1.pulsewidth[10] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0131_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold145 (.A(\Voice1.accumulator[9] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold146 (.A(\yq[10] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold147 (.A(\ctr_clkdiv25[7] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0228_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold149 (.A(\Voice1.accumulator[7] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold150 (.A(\ctr_audio[9] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0191_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold152 (.A(\VAL[0] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0674_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0048_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold155 (.A(\hvsync_gen.vpos[1] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0466_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0001_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold158 (.A(\ctr_clkdiv25[1] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0217_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold160 (.A(\LFSR[4] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold161 (.A(\hvsync_gen.vpos[0] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold162 (.A(\yq[7] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold163 (.A(\yqo[7] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold164 (.A(\yq[5] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0082_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold166 (.A(\ctr_clkdiv25[6] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold167 (.A(\yqo[10] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold168 (.A(\Voice1.pulsewidth[0] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold169 (.A(\yq[11] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0088_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold171 (.A(\hvsync_gen.hpos[3] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold172 (.A(\Voice1.pulsewidth[8] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0206_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0003_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0532_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold176 (.A(\Voice1.accumulator[10] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0163_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold178 (.A(\ctr_audio[6] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold179 (.A(\ctr_audio[19] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold180 (.A(\yq[9] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold181 (.A(\yq[6] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0083_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0011_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0167_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold185 (.A(\LFSR[1] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0092_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold187 (.A(\VAL[6] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold188 (.A(\VAL[8] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0698_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold190 (.A(\yqo[9] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold191 (.A(\Voice1.pulsewidth[6] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0203_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold193 (.A(\Voice1.accumulator[19] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0172_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold195 (.A(\LFSR[2] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold196 (.A(\Voice1.pulsewidth[5] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0202_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold198 (.A(\yqo[8] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0085_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0014_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold201 (.A(\Voice1.pulsewidth[7] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold202 (.A(\yq[8] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold203 (.A(\ctr_audio[20] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold204 (.A(\xqo[0] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold205 (.A(\Voice1.accumulator[16] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold206 (.A(\VAL[3] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0682_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0051_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0015_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0407_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0184_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold212 (.A(\hvsync_gen.vpos[9] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold213 (.A(\VAL[11] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0706_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0059_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold216 (.A(\ctr_audio[21] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold217 (.A(\ctr_audio[2] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0932_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold219 (.A(\hvsync_gen.vsync ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold220 (.A(\xqo[7] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold221 (.A(\xqo[1] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold222 (.A(\VAL[1] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0676_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold224 (.A(\hvsync_gen.vpos[3] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold225 (.A(\Voice1.accumulator[20] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold226 (.A(\hvsync_gen.hpos[8] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0534_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold228 (.A(\ctr_audio[22] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0130_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold230 (.A(\hvsync_gen.hpos[9] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0030_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold232 (.A(\Voice1.pulsewidth[3] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0197_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0121_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold235 (.A(\Voice1.pulsewidth[2] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold236 (.A(\hvsync_gen.vpos[4] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold237 (.A(\VAL[9] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold238 (.A(\hvsync_gen.vpos[6] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold239 (.A(\hvsync_gen.vpos[8] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold240 (.A(\VAL[4] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold241 (.A(\hvsync_gen.hpos[4] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0526_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold243 (.A(\VAL[12] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold244 (.A(\hvsync_gen.hpos[6] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold245 (.A(\VAL[10] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold246 (.A(\VAL[2] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold247 (.A(\xqo[3] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold248 (.A(\Voice1.accumulator[5] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold249 (.A(\hvsync_gen.vpos[8] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold250 (.A(\ctr_clkdiv25[6] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0923_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0925_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold253 (.A(\VAL[12] ),
    .X(net487));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_fill_2 FILLER_0_280 ();
 sg13g2_fill_1 FILLER_0_282 ();
 sg13g2_fill_2 FILLER_0_292 ();
 sg13g2_fill_2 FILLER_0_303 ();
 sg13g2_fill_2 FILLER_0_309 ();
 sg13g2_decap_8 FILLER_0_319 ();
 sg13g2_decap_8 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_fill_2 FILLER_1_175 ();
 sg13g2_fill_1 FILLER_1_181 ();
 sg13g2_decap_8 FILLER_1_187 ();
 sg13g2_decap_8 FILLER_1_194 ();
 sg13g2_decap_8 FILLER_1_201 ();
 sg13g2_fill_2 FILLER_1_208 ();
 sg13g2_decap_8 FILLER_1_214 ();
 sg13g2_fill_2 FILLER_1_221 ();
 sg13g2_decap_8 FILLER_1_232 ();
 sg13g2_decap_8 FILLER_1_239 ();
 sg13g2_decap_8 FILLER_1_246 ();
 sg13g2_fill_1 FILLER_1_253 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_fill_2 FILLER_1_329 ();
 sg13g2_fill_1 FILLER_1_331 ();
 sg13g2_decap_8 FILLER_1_347 ();
 sg13g2_decap_8 FILLER_1_354 ();
 sg13g2_decap_8 FILLER_1_361 ();
 sg13g2_decap_8 FILLER_1_368 ();
 sg13g2_decap_8 FILLER_1_375 ();
 sg13g2_decap_8 FILLER_1_382 ();
 sg13g2_decap_8 FILLER_1_389 ();
 sg13g2_decap_8 FILLER_1_396 ();
 sg13g2_decap_4 FILLER_1_403 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_4 FILLER_2_154 ();
 sg13g2_fill_2 FILLER_2_192 ();
 sg13g2_fill_2 FILLER_2_295 ();
 sg13g2_fill_1 FILLER_2_297 ();
 sg13g2_fill_2 FILLER_2_316 ();
 sg13g2_fill_1 FILLER_2_335 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_4 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_4 FILLER_3_133 ();
 sg13g2_fill_2 FILLER_3_137 ();
 sg13g2_fill_1 FILLER_3_165 ();
 sg13g2_fill_2 FILLER_3_175 ();
 sg13g2_fill_1 FILLER_3_186 ();
 sg13g2_decap_4 FILLER_3_212 ();
 sg13g2_fill_2 FILLER_3_253 ();
 sg13g2_fill_2 FILLER_3_287 ();
 sg13g2_fill_1 FILLER_3_289 ();
 sg13g2_fill_1 FILLER_3_331 ();
 sg13g2_fill_2 FILLER_3_393 ();
 sg13g2_fill_1 FILLER_3_395 ();
 sg13g2_decap_8 FILLER_3_400 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_4 FILLER_4_133 ();
 sg13g2_fill_1 FILLER_4_137 ();
 sg13g2_fill_1 FILLER_4_146 ();
 sg13g2_fill_2 FILLER_4_164 ();
 sg13g2_fill_1 FILLER_4_246 ();
 sg13g2_fill_1 FILLER_4_268 ();
 sg13g2_decap_4 FILLER_4_299 ();
 sg13g2_fill_1 FILLER_4_303 ();
 sg13g2_fill_2 FILLER_4_317 ();
 sg13g2_decap_4 FILLER_4_323 ();
 sg13g2_fill_1 FILLER_4_327 ();
 sg13g2_decap_4 FILLER_4_337 ();
 sg13g2_fill_1 FILLER_4_341 ();
 sg13g2_fill_2 FILLER_4_370 ();
 sg13g2_fill_2 FILLER_4_376 ();
 sg13g2_fill_1 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_fill_2 FILLER_5_35 ();
 sg13g2_fill_1 FILLER_5_37 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_4 FILLER_5_126 ();
 sg13g2_fill_1 FILLER_5_130 ();
 sg13g2_fill_2 FILLER_5_157 ();
 sg13g2_fill_2 FILLER_5_174 ();
 sg13g2_decap_4 FILLER_5_216 ();
 sg13g2_fill_1 FILLER_5_220 ();
 sg13g2_decap_8 FILLER_5_246 ();
 sg13g2_fill_1 FILLER_5_296 ();
 sg13g2_fill_1 FILLER_5_358 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_fill_2 FILLER_6_21 ();
 sg13g2_fill_1 FILLER_6_23 ();
 sg13g2_fill_1 FILLER_6_32 ();
 sg13g2_fill_2 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_69 ();
 sg13g2_decap_8 FILLER_6_76 ();
 sg13g2_decap_8 FILLER_6_83 ();
 sg13g2_decap_8 FILLER_6_90 ();
 sg13g2_decap_8 FILLER_6_97 ();
 sg13g2_decap_8 FILLER_6_104 ();
 sg13g2_decap_8 FILLER_6_111 ();
 sg13g2_decap_8 FILLER_6_118 ();
 sg13g2_fill_1 FILLER_6_125 ();
 sg13g2_fill_1 FILLER_6_166 ();
 sg13g2_fill_1 FILLER_6_224 ();
 sg13g2_fill_1 FILLER_6_267 ();
 sg13g2_fill_2 FILLER_6_299 ();
 sg13g2_fill_1 FILLER_6_306 ();
 sg13g2_fill_1 FILLER_6_320 ();
 sg13g2_fill_1 FILLER_6_330 ();
 sg13g2_decap_4 FILLER_6_335 ();
 sg13g2_fill_2 FILLER_6_339 ();
 sg13g2_fill_2 FILLER_6_344 ();
 sg13g2_fill_1 FILLER_6_354 ();
 sg13g2_fill_2 FILLER_6_380 ();
 sg13g2_fill_1 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_fill_2 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_87 ();
 sg13g2_decap_8 FILLER_7_94 ();
 sg13g2_decap_8 FILLER_7_101 ();
 sg13g2_decap_8 FILLER_7_108 ();
 sg13g2_decap_8 FILLER_7_115 ();
 sg13g2_decap_8 FILLER_7_122 ();
 sg13g2_fill_2 FILLER_7_129 ();
 sg13g2_fill_2 FILLER_7_157 ();
 sg13g2_decap_4 FILLER_7_218 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_fill_1 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_4 FILLER_7_280 ();
 sg13g2_fill_2 FILLER_7_284 ();
 sg13g2_fill_1 FILLER_7_291 ();
 sg13g2_fill_2 FILLER_7_321 ();
 sg13g2_fill_2 FILLER_7_334 ();
 sg13g2_decap_8 FILLER_7_341 ();
 sg13g2_decap_4 FILLER_7_348 ();
 sg13g2_fill_2 FILLER_7_352 ();
 sg13g2_decap_8 FILLER_7_358 ();
 sg13g2_fill_2 FILLER_7_379 ();
 sg13g2_fill_1 FILLER_7_381 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_94 ();
 sg13g2_decap_8 FILLER_8_101 ();
 sg13g2_decap_8 FILLER_8_108 ();
 sg13g2_decap_8 FILLER_8_115 ();
 sg13g2_decap_8 FILLER_8_122 ();
 sg13g2_decap_8 FILLER_8_129 ();
 sg13g2_decap_8 FILLER_8_136 ();
 sg13g2_fill_1 FILLER_8_143 ();
 sg13g2_fill_1 FILLER_8_257 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_4 FILLER_8_273 ();
 sg13g2_fill_1 FILLER_8_307 ();
 sg13g2_fill_2 FILLER_8_337 ();
 sg13g2_decap_4 FILLER_8_344 ();
 sg13g2_fill_1 FILLER_8_348 ();
 sg13g2_fill_1 FILLER_8_374 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_fill_2 FILLER_9_35 ();
 sg13g2_fill_1 FILLER_9_106 ();
 sg13g2_decap_8 FILLER_9_111 ();
 sg13g2_decap_8 FILLER_9_118 ();
 sg13g2_decap_8 FILLER_9_125 ();
 sg13g2_decap_4 FILLER_9_132 ();
 sg13g2_decap_8 FILLER_9_223 ();
 sg13g2_decap_8 FILLER_9_230 ();
 sg13g2_fill_2 FILLER_9_237 ();
 sg13g2_fill_1 FILLER_9_239 ();
 sg13g2_fill_2 FILLER_9_261 ();
 sg13g2_fill_1 FILLER_9_263 ();
 sg13g2_fill_1 FILLER_9_309 ();
 sg13g2_decap_8 FILLER_9_317 ();
 sg13g2_decap_8 FILLER_9_324 ();
 sg13g2_fill_1 FILLER_9_331 ();
 sg13g2_fill_2 FILLER_9_349 ();
 sg13g2_fill_1 FILLER_9_373 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_24 ();
 sg13g2_fill_1 FILLER_10_60 ();
 sg13g2_fill_2 FILLER_10_122 ();
 sg13g2_fill_1 FILLER_10_124 ();
 sg13g2_fill_2 FILLER_10_134 ();
 sg13g2_decap_4 FILLER_10_141 ();
 sg13g2_fill_2 FILLER_10_145 ();
 sg13g2_decap_4 FILLER_10_151 ();
 sg13g2_fill_2 FILLER_10_155 ();
 sg13g2_fill_2 FILLER_10_206 ();
 sg13g2_fill_2 FILLER_10_247 ();
 sg13g2_fill_1 FILLER_10_265 ();
 sg13g2_fill_2 FILLER_10_276 ();
 sg13g2_fill_1 FILLER_10_278 ();
 sg13g2_fill_2 FILLER_10_288 ();
 sg13g2_fill_2 FILLER_10_303 ();
 sg13g2_fill_1 FILLER_10_305 ();
 sg13g2_fill_2 FILLER_10_337 ();
 sg13g2_fill_1 FILLER_10_365 ();
 sg13g2_fill_2 FILLER_10_370 ();
 sg13g2_fill_1 FILLER_10_372 ();
 sg13g2_fill_1 FILLER_10_382 ();
 sg13g2_fill_2 FILLER_11_26 ();
 sg13g2_fill_1 FILLER_11_89 ();
 sg13g2_fill_2 FILLER_11_109 ();
 sg13g2_decap_4 FILLER_11_163 ();
 sg13g2_fill_2 FILLER_11_167 ();
 sg13g2_decap_4 FILLER_11_195 ();
 sg13g2_fill_1 FILLER_11_199 ();
 sg13g2_decap_4 FILLER_11_209 ();
 sg13g2_fill_2 FILLER_11_213 ();
 sg13g2_decap_4 FILLER_11_228 ();
 sg13g2_fill_2 FILLER_11_232 ();
 sg13g2_fill_2 FILLER_11_274 ();
 sg13g2_fill_1 FILLER_11_276 ();
 sg13g2_fill_2 FILLER_11_303 ();
 sg13g2_fill_1 FILLER_11_305 ();
 sg13g2_decap_8 FILLER_11_328 ();
 sg13g2_fill_2 FILLER_11_335 ();
 sg13g2_fill_2 FILLER_11_342 ();
 sg13g2_fill_1 FILLER_11_344 ();
 sg13g2_fill_2 FILLER_11_358 ();
 sg13g2_fill_1 FILLER_11_360 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_40 ();
 sg13g2_fill_1 FILLER_12_50 ();
 sg13g2_decap_8 FILLER_12_139 ();
 sg13g2_decap_4 FILLER_12_146 ();
 sg13g2_fill_1 FILLER_12_150 ();
 sg13g2_fill_2 FILLER_12_160 ();
 sg13g2_fill_1 FILLER_12_191 ();
 sg13g2_decap_8 FILLER_12_218 ();
 sg13g2_decap_8 FILLER_12_225 ();
 sg13g2_decap_8 FILLER_12_232 ();
 sg13g2_decap_4 FILLER_12_239 ();
 sg13g2_fill_2 FILLER_12_243 ();
 sg13g2_fill_2 FILLER_12_254 ();
 sg13g2_fill_1 FILLER_12_256 ();
 sg13g2_fill_2 FILLER_12_267 ();
 sg13g2_decap_8 FILLER_12_274 ();
 sg13g2_fill_2 FILLER_12_281 ();
 sg13g2_fill_1 FILLER_12_283 ();
 sg13g2_fill_2 FILLER_12_310 ();
 sg13g2_decap_4 FILLER_13_132 ();
 sg13g2_fill_1 FILLER_13_136 ();
 sg13g2_decap_4 FILLER_13_163 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_fill_1 FILLER_13_182 ();
 sg13g2_fill_1 FILLER_13_208 ();
 sg13g2_fill_2 FILLER_13_261 ();
 sg13g2_fill_1 FILLER_13_263 ();
 sg13g2_fill_2 FILLER_13_270 ();
 sg13g2_fill_1 FILLER_13_272 ();
 sg13g2_fill_1 FILLER_13_281 ();
 sg13g2_decap_4 FILLER_13_291 ();
 sg13g2_decap_8 FILLER_13_299 ();
 sg13g2_decap_4 FILLER_13_306 ();
 sg13g2_fill_2 FILLER_13_354 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_4 ();
 sg13g2_fill_2 FILLER_14_36 ();
 sg13g2_fill_2 FILLER_14_64 ();
 sg13g2_fill_2 FILLER_14_155 ();
 sg13g2_fill_1 FILLER_14_157 ();
 sg13g2_decap_4 FILLER_14_186 ();
 sg13g2_fill_2 FILLER_14_190 ();
 sg13g2_fill_2 FILLER_14_197 ();
 sg13g2_fill_1 FILLER_14_199 ();
 sg13g2_decap_8 FILLER_14_212 ();
 sg13g2_fill_1 FILLER_14_219 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_4 FILLER_14_231 ();
 sg13g2_fill_1 FILLER_14_235 ();
 sg13g2_fill_1 FILLER_14_270 ();
 sg13g2_fill_1 FILLER_14_302 ();
 sg13g2_decap_8 FILLER_14_307 ();
 sg13g2_fill_1 FILLER_14_314 ();
 sg13g2_fill_2 FILLER_14_333 ();
 sg13g2_fill_1 FILLER_14_335 ();
 sg13g2_fill_1 FILLER_14_350 ();
 sg13g2_fill_1 FILLER_14_375 ();
 sg13g2_fill_2 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_7 ();
 sg13g2_fill_1 FILLER_15_9 ();
 sg13g2_fill_1 FILLER_15_66 ();
 sg13g2_fill_2 FILLER_15_89 ();
 sg13g2_fill_1 FILLER_15_91 ();
 sg13g2_fill_2 FILLER_15_118 ();
 sg13g2_fill_1 FILLER_15_120 ();
 sg13g2_fill_1 FILLER_15_134 ();
 sg13g2_fill_2 FILLER_15_145 ();
 sg13g2_fill_1 FILLER_15_147 ();
 sg13g2_fill_2 FILLER_15_156 ();
 sg13g2_fill_1 FILLER_15_158 ();
 sg13g2_fill_2 FILLER_15_194 ();
 sg13g2_fill_1 FILLER_15_242 ();
 sg13g2_fill_1 FILLER_15_256 ();
 sg13g2_decap_4 FILLER_15_261 ();
 sg13g2_fill_2 FILLER_15_269 ();
 sg13g2_fill_1 FILLER_15_271 ();
 sg13g2_fill_2 FILLER_15_277 ();
 sg13g2_fill_2 FILLER_15_284 ();
 sg13g2_fill_1 FILLER_15_286 ();
 sg13g2_fill_2 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_fill_1 FILLER_15_332 ();
 sg13g2_fill_2 FILLER_15_349 ();
 sg13g2_fill_1 FILLER_15_351 ();
 sg13g2_fill_1 FILLER_15_365 ();
 sg13g2_fill_2 FILLER_15_389 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_43 ();
 sg13g2_fill_2 FILLER_16_84 ();
 sg13g2_fill_2 FILLER_16_109 ();
 sg13g2_fill_2 FILLER_16_163 ();
 sg13g2_fill_2 FILLER_16_181 ();
 sg13g2_fill_1 FILLER_16_191 ();
 sg13g2_decap_4 FILLER_16_214 ();
 sg13g2_fill_2 FILLER_16_218 ();
 sg13g2_decap_8 FILLER_16_229 ();
 sg13g2_fill_2 FILLER_16_236 ();
 sg13g2_fill_1 FILLER_16_238 ();
 sg13g2_fill_1 FILLER_16_248 ();
 sg13g2_fill_2 FILLER_16_259 ();
 sg13g2_fill_1 FILLER_16_261 ();
 sg13g2_decap_8 FILLER_16_288 ();
 sg13g2_decap_4 FILLER_16_295 ();
 sg13g2_fill_2 FILLER_16_299 ();
 sg13g2_decap_4 FILLER_16_309 ();
 sg13g2_fill_2 FILLER_16_313 ();
 sg13g2_fill_2 FILLER_16_335 ();
 sg13g2_fill_1 FILLER_16_337 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_fill_1 FILLER_16_361 ();
 sg13g2_decap_4 FILLER_16_367 ();
 sg13g2_fill_2 FILLER_16_391 ();
 sg13g2_fill_1 FILLER_16_393 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_21 ();
 sg13g2_fill_2 FILLER_17_65 ();
 sg13g2_fill_1 FILLER_17_67 ();
 sg13g2_decap_8 FILLER_17_149 ();
 sg13g2_fill_2 FILLER_17_156 ();
 sg13g2_fill_1 FILLER_17_158 ();
 sg13g2_fill_2 FILLER_17_179 ();
 sg13g2_fill_1 FILLER_17_181 ();
 sg13g2_decap_4 FILLER_17_190 ();
 sg13g2_fill_2 FILLER_17_212 ();
 sg13g2_fill_2 FILLER_17_232 ();
 sg13g2_fill_1 FILLER_17_234 ();
 sg13g2_fill_2 FILLER_17_271 ();
 sg13g2_fill_1 FILLER_17_277 ();
 sg13g2_decap_4 FILLER_17_282 ();
 sg13g2_fill_1 FILLER_17_289 ();
 sg13g2_fill_1 FILLER_17_298 ();
 sg13g2_fill_2 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_337 ();
 sg13g2_decap_8 FILLER_17_349 ();
 sg13g2_fill_2 FILLER_17_380 ();
 sg13g2_fill_1 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_79 ();
 sg13g2_fill_1 FILLER_18_174 ();
 sg13g2_decap_4 FILLER_18_184 ();
 sg13g2_decap_4 FILLER_18_192 ();
 sg13g2_fill_2 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_202 ();
 sg13g2_decap_8 FILLER_18_209 ();
 sg13g2_fill_1 FILLER_18_216 ();
 sg13g2_fill_1 FILLER_18_227 ();
 sg13g2_decap_4 FILLER_18_254 ();
 sg13g2_decap_4 FILLER_18_263 ();
 sg13g2_fill_1 FILLER_18_267 ();
 sg13g2_decap_8 FILLER_18_306 ();
 sg13g2_decap_4 FILLER_18_313 ();
 sg13g2_fill_2 FILLER_18_317 ();
 sg13g2_fill_2 FILLER_18_327 ();
 sg13g2_decap_8 FILLER_18_342 ();
 sg13g2_fill_1 FILLER_18_349 ();
 sg13g2_decap_8 FILLER_18_366 ();
 sg13g2_decap_4 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_7 ();
 sg13g2_fill_1 FILLER_19_38 ();
 sg13g2_fill_2 FILLER_19_72 ();
 sg13g2_fill_1 FILLER_19_100 ();
 sg13g2_fill_2 FILLER_19_130 ();
 sg13g2_fill_1 FILLER_19_132 ();
 sg13g2_decap_4 FILLER_19_146 ();
 sg13g2_decap_8 FILLER_19_167 ();
 sg13g2_decap_8 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_fill_1 FILLER_19_190 ();
 sg13g2_decap_4 FILLER_19_234 ();
 sg13g2_fill_1 FILLER_19_248 ();
 sg13g2_decap_4 FILLER_19_255 ();
 sg13g2_fill_2 FILLER_19_289 ();
 sg13g2_decap_8 FILLER_19_317 ();
 sg13g2_fill_2 FILLER_19_324 ();
 sg13g2_fill_1 FILLER_19_326 ();
 sg13g2_fill_1 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_370 ();
 sg13g2_fill_1 FILLER_19_377 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_4 ();
 sg13g2_fill_2 FILLER_20_34 ();
 sg13g2_fill_1 FILLER_20_56 ();
 sg13g2_fill_1 FILLER_20_79 ();
 sg13g2_fill_1 FILLER_20_115 ();
 sg13g2_fill_1 FILLER_20_147 ();
 sg13g2_fill_2 FILLER_20_216 ();
 sg13g2_fill_1 FILLER_20_218 ();
 sg13g2_fill_1 FILLER_20_244 ();
 sg13g2_decap_8 FILLER_20_249 ();
 sg13g2_decap_4 FILLER_20_256 ();
 sg13g2_fill_2 FILLER_20_260 ();
 sg13g2_fill_2 FILLER_20_265 ();
 sg13g2_fill_1 FILLER_20_313 ();
 sg13g2_decap_8 FILLER_20_345 ();
 sg13g2_fill_2 FILLER_20_352 ();
 sg13g2_fill_1 FILLER_20_354 ();
 sg13g2_decap_8 FILLER_20_368 ();
 sg13g2_fill_2 FILLER_20_375 ();
 sg13g2_fill_1 FILLER_20_377 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_fill_2 FILLER_21_109 ();
 sg13g2_decap_4 FILLER_21_123 ();
 sg13g2_fill_2 FILLER_21_131 ();
 sg13g2_fill_1 FILLER_21_133 ();
 sg13g2_fill_1 FILLER_21_182 ();
 sg13g2_fill_2 FILLER_21_198 ();
 sg13g2_fill_1 FILLER_21_200 ();
 sg13g2_fill_2 FILLER_21_236 ();
 sg13g2_fill_1 FILLER_21_238 ();
 sg13g2_fill_2 FILLER_21_332 ();
 sg13g2_fill_2 FILLER_21_374 ();
 sg13g2_fill_1 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_21_383 ();
 sg13g2_fill_1 FILLER_21_390 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_4 ();
 sg13g2_fill_1 FILLER_22_22 ();
 sg13g2_fill_1 FILLER_22_73 ();
 sg13g2_fill_2 FILLER_22_102 ();
 sg13g2_fill_1 FILLER_22_104 ();
 sg13g2_fill_2 FILLER_22_135 ();
 sg13g2_fill_2 FILLER_22_151 ();
 sg13g2_fill_2 FILLER_22_171 ();
 sg13g2_fill_1 FILLER_22_260 ();
 sg13g2_decap_4 FILLER_22_265 ();
 sg13g2_fill_2 FILLER_22_269 ();
 sg13g2_fill_2 FILLER_22_302 ();
 sg13g2_fill_1 FILLER_22_304 ();
 sg13g2_fill_2 FILLER_22_317 ();
 sg13g2_fill_1 FILLER_22_323 ();
 sg13g2_fill_2 FILLER_22_337 ();
 sg13g2_fill_2 FILLER_22_369 ();
 sg13g2_fill_1 FILLER_22_371 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_fill_2 FILLER_23_26 ();
 sg13g2_fill_2 FILLER_23_63 ();
 sg13g2_fill_1 FILLER_23_109 ();
 sg13g2_fill_1 FILLER_23_147 ();
 sg13g2_fill_2 FILLER_23_169 ();
 sg13g2_fill_1 FILLER_23_171 ();
 sg13g2_fill_2 FILLER_23_195 ();
 sg13g2_fill_1 FILLER_23_197 ();
 sg13g2_fill_2 FILLER_23_206 ();
 sg13g2_fill_2 FILLER_23_232 ();
 sg13g2_fill_1 FILLER_23_234 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_fill_2 FILLER_23_252 ();
 sg13g2_fill_1 FILLER_23_254 ();
 sg13g2_fill_2 FILLER_23_276 ();
 sg13g2_fill_2 FILLER_23_283 ();
 sg13g2_fill_1 FILLER_23_285 ();
 sg13g2_fill_2 FILLER_23_301 ();
 sg13g2_fill_2 FILLER_23_312 ();
 sg13g2_fill_2 FILLER_23_322 ();
 sg13g2_fill_1 FILLER_23_324 ();
 sg13g2_fill_2 FILLER_23_372 ();
 sg13g2_fill_2 FILLER_23_388 ();
 sg13g2_fill_1 FILLER_23_390 ();
 sg13g2_fill_2 FILLER_23_395 ();
 sg13g2_fill_1 FILLER_23_397 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_19 ();
 sg13g2_fill_2 FILLER_24_92 ();
 sg13g2_fill_1 FILLER_24_199 ();
 sg13g2_fill_1 FILLER_24_226 ();
 sg13g2_decap_4 FILLER_24_261 ();
 sg13g2_decap_4 FILLER_24_273 ();
 sg13g2_fill_1 FILLER_24_277 ();
 sg13g2_fill_1 FILLER_24_288 ();
 sg13g2_fill_2 FILLER_24_321 ();
 sg13g2_fill_2 FILLER_24_344 ();
 sg13g2_fill_1 FILLER_24_346 ();
 sg13g2_fill_1 FILLER_24_378 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_69 ();
 sg13g2_fill_2 FILLER_25_138 ();
 sg13g2_fill_1 FILLER_25_144 ();
 sg13g2_decap_8 FILLER_25_149 ();
 sg13g2_fill_2 FILLER_25_156 ();
 sg13g2_fill_1 FILLER_25_180 ();
 sg13g2_fill_2 FILLER_25_203 ();
 sg13g2_decap_4 FILLER_25_221 ();
 sg13g2_decap_4 FILLER_25_242 ();
 sg13g2_fill_1 FILLER_25_246 ();
 sg13g2_fill_2 FILLER_25_264 ();
 sg13g2_decap_8 FILLER_25_276 ();
 sg13g2_fill_2 FILLER_25_283 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_fill_2 FILLER_25_308 ();
 sg13g2_fill_1 FILLER_25_310 ();
 sg13g2_fill_2 FILLER_25_316 ();
 sg13g2_fill_1 FILLER_25_339 ();
 sg13g2_fill_2 FILLER_25_370 ();
 sg13g2_fill_1 FILLER_25_372 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_60 ();
 sg13g2_fill_1 FILLER_26_73 ();
 sg13g2_fill_2 FILLER_26_95 ();
 sg13g2_fill_1 FILLER_26_116 ();
 sg13g2_decap_4 FILLER_26_155 ();
 sg13g2_fill_2 FILLER_26_215 ();
 sg13g2_fill_1 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_233 ();
 sg13g2_fill_1 FILLER_26_240 ();
 sg13g2_fill_1 FILLER_26_254 ();
 sg13g2_decap_4 FILLER_26_302 ();
 sg13g2_fill_2 FILLER_26_306 ();
 sg13g2_fill_2 FILLER_26_365 ();
 sg13g2_fill_1 FILLER_26_367 ();
 sg13g2_fill_1 FILLER_26_382 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_73 ();
 sg13g2_fill_2 FILLER_27_139 ();
 sg13g2_decap_4 FILLER_27_222 ();
 sg13g2_fill_1 FILLER_27_226 ();
 sg13g2_fill_1 FILLER_27_240 ();
 sg13g2_decap_8 FILLER_27_249 ();
 sg13g2_fill_2 FILLER_27_256 ();
 sg13g2_fill_2 FILLER_27_270 ();
 sg13g2_decap_8 FILLER_27_276 ();
 sg13g2_decap_4 FILLER_27_283 ();
 sg13g2_decap_4 FILLER_27_291 ();
 sg13g2_fill_1 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_304 ();
 sg13g2_fill_2 FILLER_27_311 ();
 sg13g2_fill_2 FILLER_27_342 ();
 sg13g2_fill_2 FILLER_27_357 ();
 sg13g2_fill_1 FILLER_27_359 ();
 sg13g2_fill_1 FILLER_28_32 ();
 sg13g2_fill_2 FILLER_28_75 ();
 sg13g2_fill_1 FILLER_28_90 ();
 sg13g2_fill_1 FILLER_28_130 ();
 sg13g2_decap_4 FILLER_28_164 ();
 sg13g2_fill_1 FILLER_28_181 ();
 sg13g2_fill_2 FILLER_28_186 ();
 sg13g2_fill_1 FILLER_28_188 ();
 sg13g2_fill_1 FILLER_28_208 ();
 sg13g2_fill_2 FILLER_28_222 ();
 sg13g2_decap_4 FILLER_28_249 ();
 sg13g2_fill_1 FILLER_28_253 ();
 sg13g2_fill_1 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_327 ();
 sg13g2_fill_2 FILLER_28_363 ();
 sg13g2_fill_2 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_68 ();
 sg13g2_fill_1 FILLER_29_85 ();
 sg13g2_fill_2 FILLER_29_89 ();
 sg13g2_fill_2 FILLER_29_136 ();
 sg13g2_fill_1 FILLER_29_151 ();
 sg13g2_fill_1 FILLER_29_187 ();
 sg13g2_decap_4 FILLER_29_204 ();
 sg13g2_fill_2 FILLER_29_215 ();
 sg13g2_fill_1 FILLER_29_232 ();
 sg13g2_decap_8 FILLER_29_248 ();
 sg13g2_fill_1 FILLER_29_255 ();
 sg13g2_fill_1 FILLER_29_264 ();
 sg13g2_decap_8 FILLER_29_275 ();
 sg13g2_fill_2 FILLER_29_286 ();
 sg13g2_fill_1 FILLER_29_288 ();
 sg13g2_fill_1 FILLER_29_306 ();
 sg13g2_fill_2 FILLER_29_343 ();
 sg13g2_fill_2 FILLER_29_350 ();
 sg13g2_fill_2 FILLER_29_370 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_25 ();
 sg13g2_fill_1 FILLER_30_48 ();
 sg13g2_fill_1 FILLER_30_103 ();
 sg13g2_fill_1 FILLER_30_113 ();
 sg13g2_fill_2 FILLER_30_181 ();
 sg13g2_fill_1 FILLER_30_209 ();
 sg13g2_decap_8 FILLER_30_220 ();
 sg13g2_fill_2 FILLER_30_227 ();
 sg13g2_fill_2 FILLER_30_259 ();
 sg13g2_decap_4 FILLER_30_266 ();
 sg13g2_fill_1 FILLER_30_270 ();
 sg13g2_fill_2 FILLER_30_297 ();
 sg13g2_fill_1 FILLER_30_308 ();
 sg13g2_fill_1 FILLER_30_335 ();
 sg13g2_fill_2 FILLER_30_366 ();
 sg13g2_fill_1 FILLER_31_94 ();
 sg13g2_fill_2 FILLER_31_121 ();
 sg13g2_fill_1 FILLER_31_123 ();
 sg13g2_fill_1 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_175 ();
 sg13g2_fill_2 FILLER_31_193 ();
 sg13g2_fill_1 FILLER_31_195 ();
 sg13g2_decap_8 FILLER_31_222 ();
 sg13g2_decap_8 FILLER_31_229 ();
 sg13g2_fill_1 FILLER_31_236 ();
 sg13g2_fill_2 FILLER_31_307 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_53 ();
 sg13g2_fill_1 FILLER_32_69 ();
 sg13g2_decap_4 FILLER_32_101 ();
 sg13g2_fill_1 FILLER_32_105 ();
 sg13g2_fill_1 FILLER_32_110 ();
 sg13g2_fill_1 FILLER_32_137 ();
 sg13g2_fill_2 FILLER_32_143 ();
 sg13g2_decap_8 FILLER_32_150 ();
 sg13g2_decap_4 FILLER_32_161 ();
 sg13g2_fill_1 FILLER_32_165 ();
 sg13g2_fill_2 FILLER_32_194 ();
 sg13g2_fill_2 FILLER_32_205 ();
 sg13g2_decap_4 FILLER_32_211 ();
 sg13g2_fill_1 FILLER_32_215 ();
 sg13g2_decap_4 FILLER_32_242 ();
 sg13g2_fill_1 FILLER_32_246 ();
 sg13g2_fill_1 FILLER_32_277 ();
 sg13g2_fill_2 FILLER_32_301 ();
 sg13g2_fill_2 FILLER_32_329 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_fill_2 FILLER_32_352 ();
 sg13g2_fill_1 FILLER_33_42 ();
 sg13g2_fill_1 FILLER_33_74 ();
 sg13g2_fill_2 FILLER_33_104 ();
 sg13g2_fill_2 FILLER_33_115 ();
 sg13g2_decap_8 FILLER_33_141 ();
 sg13g2_fill_2 FILLER_33_148 ();
 sg13g2_fill_1 FILLER_33_150 ();
 sg13g2_fill_2 FILLER_33_168 ();
 sg13g2_fill_1 FILLER_33_170 ();
 sg13g2_fill_2 FILLER_33_175 ();
 sg13g2_fill_1 FILLER_33_177 ();
 sg13g2_decap_8 FILLER_33_199 ();
 sg13g2_decap_4 FILLER_33_206 ();
 sg13g2_fill_2 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_216 ();
 sg13g2_decap_4 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_268 ();
 sg13g2_fill_1 FILLER_33_286 ();
 sg13g2_fill_2 FILLER_33_312 ();
 sg13g2_fill_1 FILLER_33_337 ();
 sg13g2_fill_1 FILLER_33_394 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_fill_2 FILLER_34_20 ();
 sg13g2_fill_1 FILLER_34_60 ();
 sg13g2_fill_2 FILLER_34_116 ();
 sg13g2_fill_1 FILLER_34_128 ();
 sg13g2_fill_2 FILLER_34_134 ();
 sg13g2_fill_1 FILLER_34_136 ();
 sg13g2_fill_2 FILLER_34_166 ();
 sg13g2_fill_2 FILLER_34_199 ();
 sg13g2_fill_1 FILLER_34_245 ();
 sg13g2_fill_1 FILLER_34_256 ();
 sg13g2_fill_1 FILLER_34_325 ();
 sg13g2_fill_1 FILLER_34_362 ();
 sg13g2_fill_2 FILLER_34_368 ();
 sg13g2_fill_2 FILLER_34_375 ();
 sg13g2_fill_1 FILLER_34_377 ();
 sg13g2_fill_2 FILLER_35_50 ();
 sg13g2_fill_1 FILLER_35_52 ();
 sg13g2_fill_1 FILLER_35_123 ();
 sg13g2_fill_2 FILLER_35_135 ();
 sg13g2_fill_2 FILLER_35_140 ();
 sg13g2_fill_1 FILLER_35_157 ();
 sg13g2_fill_2 FILLER_35_170 ();
 sg13g2_fill_2 FILLER_35_201 ();
 sg13g2_decap_8 FILLER_35_207 ();
 sg13g2_decap_4 FILLER_35_214 ();
 sg13g2_fill_1 FILLER_35_218 ();
 sg13g2_fill_2 FILLER_35_272 ();
 sg13g2_fill_2 FILLER_35_278 ();
 sg13g2_fill_1 FILLER_35_311 ();
 sg13g2_fill_2 FILLER_35_356 ();
 sg13g2_fill_1 FILLER_35_358 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_24 ();
 sg13g2_fill_2 FILLER_36_43 ();
 sg13g2_fill_1 FILLER_36_45 ();
 sg13g2_fill_2 FILLER_36_123 ();
 sg13g2_fill_2 FILLER_36_148 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_fill_1 FILLER_36_180 ();
 sg13g2_fill_2 FILLER_36_185 ();
 sg13g2_fill_1 FILLER_36_221 ();
 sg13g2_fill_1 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_338 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_98 ();
 sg13g2_fill_2 FILLER_37_160 ();
 sg13g2_decap_8 FILLER_37_193 ();
 sg13g2_decap_8 FILLER_37_200 ();
 sg13g2_decap_8 FILLER_37_207 ();
 sg13g2_decap_8 FILLER_37_214 ();
 sg13g2_fill_2 FILLER_37_234 ();
 sg13g2_fill_2 FILLER_37_255 ();
 sg13g2_fill_1 FILLER_37_285 ();
 sg13g2_fill_1 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_45 ();
 sg13g2_fill_2 FILLER_38_80 ();
 sg13g2_fill_1 FILLER_38_82 ();
 sg13g2_fill_2 FILLER_38_97 ();
 sg13g2_fill_1 FILLER_38_99 ();
 sg13g2_fill_1 FILLER_38_135 ();
 sg13g2_fill_2 FILLER_38_175 ();
 sg13g2_fill_1 FILLER_38_181 ();
 sg13g2_decap_8 FILLER_38_198 ();
 sg13g2_decap_8 FILLER_38_205 ();
 sg13g2_decap_8 FILLER_38_212 ();
 sg13g2_fill_2 FILLER_38_219 ();
 sg13g2_fill_1 FILLER_38_221 ();
 sg13g2_decap_4 FILLER_38_257 ();
 sg13g2_fill_1 FILLER_38_297 ();
 sg13g2_fill_2 FILLER_38_324 ();
 sg13g2_fill_1 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_361 ();
 sg13g2_fill_2 FILLER_38_371 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net234;
 assign uio_out[0] = net8;
 assign uio_out[1] = net9;
 assign uio_out[2] = net10;
 assign uio_out[3] = net11;
 assign uio_out[4] = net12;
 assign uio_out[5] = net13;
 assign uio_out[6] = net14;
endmodule

module tt_um_idann (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire f0p_o;
 wire \final_o[0] ;
 wire \final_o[10] ;
 wire \final_o[1] ;
 wire \final_o[2] ;
 wire \final_o[3] ;
 wire \final_o[4] ;
 wire \final_o[5] ;
 wire \final_o[6] ;
 wire \final_o[7] ;
 wire \final_o[8] ;
 wire \final_o[9] ;
 wire \hn0.hidden_neuron_o[0] ;
 wire \hn0.hidden_neuron_o[1] ;
 wire \hn0.hidden_neuron_o[2] ;
 wire \hn0.hidden_neuron_o[3] ;
 wire \hn1.hidden_neuron_o[0] ;
 wire \hn1.hidden_neuron_o[1] ;
 wire \hn1.hidden_neuron_o[2] ;
 wire \hn1.hidden_neuron_o[3] ;
 wire \hn2.hidden_neuron_o[0] ;
 wire \hn2.hidden_neuron_o[1] ;
 wire \hn2.hidden_neuron_o[2] ;
 wire \hn2.hidden_neuron_o[3] ;
 wire \hn3.hidden_neuron_o[0] ;
 wire \hn3.hidden_neuron_o[1] ;
 wire \hn3.hidden_neuron_o[2] ;
 wire \hn3.hidden_neuron_o[3] ;
 wire \hn4.hidden_neuron_o[0] ;
 wire \hn4.hidden_neuron_o[1] ;
 wire \hn4.hidden_neuron_o[2] ;
 wire \hn4.hidden_neuron_o[3] ;
 wire \hn4.hidden_neuron_o[4] ;
 wire \hn5.hidden_neuron_o[0] ;
 wire \hn5.hidden_neuron_o[1] ;
 wire \hn5.hidden_neuron_o[2] ;
 wire \hn5.hidden_neuron_o[3] ;
 wire \hn5.hidden_neuron_o[4] ;
 wire \hn6.hidden_neuron_o[0] ;
 wire \hn6.hidden_neuron_o[1] ;
 wire \hn6.hidden_neuron_o[2] ;
 wire \hn6.hidden_neuron_o[3] ;
 wire \hn6.hidden_neuron_o[4] ;
 wire \hn7.hidden_neuron_o[0] ;
 wire \hn7.hidden_neuron_o[1] ;
 wire \hn7.hidden_neuron_o[2] ;
 wire \hn7.hidden_neuron_o[3] ;
 wire \hn7.hidden_neuron_o[4] ;
 wire \sm0.state_d[1] ;
 wire clknet_0_clk;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;

 sg13g2_inv_1 _0492_ (.Y(_0055_),
    .A(\hn4.hidden_neuron_o[4] ));
 sg13g2_inv_1 _0493_ (.Y(_0056_),
    .A(net87));
 sg13g2_inv_1 _0494_ (.Y(_0057_),
    .A(net65));
 sg13g2_inv_1 _0495_ (.Y(_0058_),
    .A(net131));
 sg13g2_inv_1 _0496_ (.Y(_0059_),
    .A(\hn6.hidden_neuron_o[2] ));
 sg13g2_inv_1 _0497_ (.Y(_0060_),
    .A(\hn6.hidden_neuron_o[0] ));
 sg13g2_inv_1 _0498_ (.Y(_0061_),
    .A(uio_out[5]));
 sg13g2_inv_1 _0499_ (.Y(_0062_),
    .A(net110));
 sg13g2_inv_1 _0500_ (.Y(_0063_),
    .A(net99));
 sg13g2_inv_1 _0501_ (.Y(_0064_),
    .A(_0001_));
 sg13g2_inv_1 _0502_ (.Y(_0065_),
    .A(_0002_));
 sg13g2_inv_1 _0503_ (.Y(_0066_),
    .A(_0004_));
 sg13g2_inv_1 _0504_ (.Y(_0067_),
    .A(net105));
 sg13g2_nor2_1 _0505_ (.A(uio_out[6]),
    .B(_0061_),
    .Y(\sm0.state_d[1] ));
 sg13g2_and2_1 _0506_ (.A(net128),
    .B(net124),
    .X(_0000_));
 sg13g2_o21ai_1 _0507_ (.B1(net91),
    .Y(_0068_),
    .A1(net1),
    .A2(net3));
 sg13g2_a21o_2 _0508_ (.A2(net3),
    .A1(net1),
    .B1(_0068_),
    .X(_0069_));
 sg13g2_nand2_1 _0509_ (.Y(_0070_),
    .A(net82),
    .B(net123));
 sg13g2_a21oi_1 _0510_ (.A1(_0069_),
    .A2(_0070_),
    .Y(_0006_),
    .B1(net93));
 sg13g2_nor2_2 _0511_ (.A(net99),
    .B(net100),
    .Y(_0071_));
 sg13g2_nor2_1 _0512_ (.A(net86),
    .B(_0071_),
    .Y(_0072_));
 sg13g2_nor2_1 _0513_ (.A(net100),
    .B(net97),
    .Y(_0073_));
 sg13g2_or2_1 _0514_ (.X(_0074_),
    .B(net97),
    .A(net100));
 sg13g2_nand2_1 _0515_ (.Y(_0075_),
    .A(net100),
    .B(net97));
 sg13g2_nand3_1 _0516_ (.B(_0074_),
    .C(_0075_),
    .A(net99),
    .Y(_0076_));
 sg13g2_nand2_1 _0517_ (.Y(_0077_),
    .A(_0072_),
    .B(_0076_));
 sg13g2_nand2_1 _0518_ (.Y(_0078_),
    .A(net84),
    .B(net127));
 sg13g2_a21oi_1 _0519_ (.A1(_0077_),
    .A2(_0078_),
    .Y(_0007_),
    .B1(net95));
 sg13g2_nand2_1 _0520_ (.Y(_0079_),
    .A(net83),
    .B(net111));
 sg13g2_nor3_1 _0521_ (.A(net99),
    .B(net100),
    .C(net97),
    .Y(_0080_));
 sg13g2_nand3b_1 _0522_ (.B(net90),
    .C(_0075_),
    .Y(_0081_),
    .A_N(_0080_));
 sg13g2_a21oi_1 _0523_ (.A1(_0079_),
    .A2(_0081_),
    .Y(_0008_),
    .B1(net94));
 sg13g2_and2_2 _0524_ (.A(net97),
    .B(net98),
    .X(_0082_));
 sg13g2_nand2_1 _0525_ (.Y(_0083_),
    .A(net97),
    .B(net98));
 sg13g2_nor2_2 _0526_ (.A(_0071_),
    .B(_0083_),
    .Y(_0084_));
 sg13g2_nor2_2 _0527_ (.A(net97),
    .B(net98),
    .Y(_0085_));
 sg13g2_nand2_2 _0528_ (.Y(_0086_),
    .A(net99),
    .B(net100));
 sg13g2_or2_1 _0529_ (.X(_0087_),
    .B(net98),
    .A(net1));
 sg13g2_o21ai_1 _0530_ (.B1(_0086_),
    .Y(_0088_),
    .A1(net100),
    .A2(_0087_));
 sg13g2_nor3_1 _0531_ (.A(_0084_),
    .B(_0085_),
    .C(_0088_),
    .Y(_0089_));
 sg13g2_nor2_2 _0532_ (.A(_0082_),
    .B(_0085_),
    .Y(_0090_));
 sg13g2_o21ai_1 _0533_ (.B1(net89),
    .Y(_0091_),
    .A1(_0086_),
    .A2(_0090_));
 sg13g2_o21ai_1 _0534_ (.B1(net104),
    .Y(_0092_),
    .A1(_0089_),
    .A2(_0091_));
 sg13g2_a21oi_1 _0535_ (.A1(net83),
    .A2(_0062_),
    .Y(_0009_),
    .B1(_0092_));
 sg13g2_nand2_1 _0536_ (.Y(_0093_),
    .A(net81),
    .B(net79));
 sg13g2_nor2_1 _0537_ (.A(_0085_),
    .B(_0086_),
    .Y(_0094_));
 sg13g2_nand2_1 _0538_ (.Y(_0095_),
    .A(net90),
    .B(_0094_));
 sg13g2_o21ai_1 _0539_ (.B1(net90),
    .Y(_0096_),
    .A1(_0084_),
    .A2(_0094_));
 sg13g2_a21oi_1 _0540_ (.A1(_0093_),
    .A2(_0096_),
    .Y(_0010_),
    .B1(net93));
 sg13g2_nor4_1 _0541_ (.A(_0061_),
    .B(net61),
    .C(net59),
    .D(net60),
    .Y(_0097_));
 sg13g2_nor2_1 _0542_ (.A(_0074_),
    .B(_0087_),
    .Y(_0098_));
 sg13g2_nor4_1 _0543_ (.A(\final_o[6] ),
    .B(\final_o[9] ),
    .C(\final_o[8] ),
    .D(net56),
    .Y(_0099_));
 sg13g2_nor4_1 _0544_ (.A(\final_o[2] ),
    .B(\final_o[5] ),
    .C(net58),
    .D(net63),
    .Y(_0100_));
 sg13g2_nand4_1 _0545_ (.B(_0098_),
    .C(_0099_),
    .A(_0097_),
    .Y(_0101_),
    .D(_0100_));
 sg13g2_nand2b_1 _0546_ (.Y(_0102_),
    .B(_0101_),
    .A_N(net128));
 sg13g2_o21ai_1 _0547_ (.B1(net102),
    .Y(_0103_),
    .A1(net124),
    .A2(net4));
 sg13g2_nor2_1 _0548_ (.A(_0102_),
    .B(_0103_),
    .Y(_0011_));
 sg13g2_nand2_1 _0549_ (.Y(_0104_),
    .A(net102),
    .B(_0102_));
 sg13g2_nor2_1 _0550_ (.A(_0000_),
    .B(_0104_),
    .Y(_0012_));
 sg13g2_nand2_1 _0551_ (.Y(_0105_),
    .A(net82),
    .B(net120));
 sg13g2_a21oi_1 _0552_ (.A1(net101),
    .A2(net2),
    .Y(_0106_),
    .B1(net84));
 sg13g2_o21ai_1 _0553_ (.B1(_0106_),
    .Y(_0107_),
    .A1(net101),
    .A2(net98));
 sg13g2_a21oi_1 _0554_ (.A1(_0105_),
    .A2(_0107_),
    .Y(_0013_),
    .B1(net93));
 sg13g2_a21oi_1 _0555_ (.A1(net100),
    .A2(_0090_),
    .Y(_0108_),
    .B1(_0073_));
 sg13g2_nand2_1 _0556_ (.Y(_0109_),
    .A(net91),
    .B(_0108_));
 sg13g2_nand2_1 _0557_ (.Y(_0110_),
    .A(net82),
    .B(net114));
 sg13g2_a21oi_1 _0558_ (.A1(_0109_),
    .A2(_0110_),
    .Y(_0014_),
    .B1(net96));
 sg13g2_nor2_1 _0559_ (.A(net98),
    .B(_0074_),
    .Y(_0111_));
 sg13g2_o21ai_1 _0560_ (.B1(net90),
    .Y(_0112_),
    .A1(_0082_),
    .A2(_0111_));
 sg13g2_inv_1 _0561_ (.Y(_0113_),
    .A(_0112_));
 sg13g2_o21ai_1 _0562_ (.B1(net103),
    .Y(_0114_),
    .A1(net88),
    .A2(net130));
 sg13g2_nor2_1 _0563_ (.A(_0113_),
    .B(_0114_),
    .Y(_0015_));
 sg13g2_nor2_2 _0564_ (.A(_0071_),
    .B(_0094_),
    .Y(_0115_));
 sg13g2_nor2_1 _0565_ (.A(net97),
    .B(_0087_),
    .Y(_0116_));
 sg13g2_nand2b_1 _0566_ (.Y(_0117_),
    .B(_0115_),
    .A_N(_0116_));
 sg13g2_a22oi_1 _0567_ (.Y(_0118_),
    .B1(_0117_),
    .B2(_0083_),
    .A2(_0086_),
    .A1(_0084_));
 sg13g2_o21ai_1 _0568_ (.B1(net104),
    .Y(_0119_),
    .A1(net83),
    .A2(_0118_));
 sg13g2_a21oi_1 _0569_ (.A1(net81),
    .A2(_0058_),
    .Y(_0016_),
    .B1(_0119_));
 sg13g2_nand2_1 _0570_ (.Y(_0120_),
    .A(net81),
    .B(net119));
 sg13g2_a21oi_1 _0571_ (.A1(_0096_),
    .A2(_0120_),
    .Y(_0017_),
    .B1(net93));
 sg13g2_nand2_1 _0572_ (.Y(_0121_),
    .A(net82),
    .B(net76));
 sg13g2_a21oi_1 _0573_ (.A1(_0069_),
    .A2(_0121_),
    .Y(_0018_),
    .B1(net96));
 sg13g2_nand2_1 _0574_ (.Y(_0122_),
    .A(net99),
    .B(net98));
 sg13g2_nand2_1 _0575_ (.Y(_0123_),
    .A(net90),
    .B(_0122_));
 sg13g2_a21oi_1 _0576_ (.A1(_0063_),
    .A2(_0090_),
    .Y(_0124_),
    .B1(_0123_));
 sg13g2_o21ai_1 _0577_ (.B1(net103),
    .Y(_0125_),
    .A1(net87),
    .A2(net112));
 sg13g2_nor2_1 _0578_ (.A(_0124_),
    .B(_0125_),
    .Y(_0019_));
 sg13g2_nor2_1 _0579_ (.A(_0116_),
    .B(_0123_),
    .Y(_0126_));
 sg13g2_a21oi_1 _0580_ (.A1(net81),
    .A2(net106),
    .Y(_0127_),
    .B1(_0126_));
 sg13g2_nor2_1 _0581_ (.A(net93),
    .B(_0127_),
    .Y(_0020_));
 sg13g2_o21ai_1 _0582_ (.B1(net105),
    .Y(_0128_),
    .A1(net89),
    .A2(net117));
 sg13g2_nor2_1 _0583_ (.A(_0082_),
    .B(_0115_),
    .Y(_0129_));
 sg13g2_a221oi_1 _0584_ (.B2(net89),
    .C1(_0128_),
    .B1(_0129_),
    .A1(_0113_),
    .Y(_0021_),
    .A2(_0115_));
 sg13g2_nand2_1 _0585_ (.Y(_0130_),
    .A(net81),
    .B(net75));
 sg13g2_a21oi_1 _0586_ (.A1(_0096_),
    .A2(_0130_),
    .Y(_0022_),
    .B1(net93));
 sg13g2_nor2_1 _0587_ (.A(net92),
    .B(net59),
    .Y(_0131_));
 sg13g2_and2_1 _0588_ (.A(\hn4.hidden_neuron_o[0] ),
    .B(\hn0.hidden_neuron_o[0] ),
    .X(_0132_));
 sg13g2_xor2_1 _0589_ (.B(\hn0.hidden_neuron_o[0] ),
    .A(\hn4.hidden_neuron_o[0] ),
    .X(_0133_));
 sg13g2_xnor2_1 _0590_ (.Y(_0134_),
    .A(\hn2.hidden_neuron_o[0] ),
    .B(_0133_));
 sg13g2_nor2_1 _0591_ (.A(_0060_),
    .B(_0134_),
    .Y(_0135_));
 sg13g2_xnor2_1 _0592_ (.Y(_0136_),
    .A(_0060_),
    .B(_0134_));
 sg13g2_a21oi_1 _0593_ (.A1(net88),
    .A2(_0136_),
    .Y(_0023_),
    .B1(_0131_));
 sg13g2_xor2_1 _0594_ (.B(\hn6.hidden_neuron_o[0] ),
    .A(\hn6.hidden_neuron_o[1] ),
    .X(_0137_));
 sg13g2_nand2_1 _0595_ (.Y(_0138_),
    .A(\hn5.hidden_neuron_o[0] ),
    .B(_0137_));
 sg13g2_xnor2_1 _0596_ (.Y(_0139_),
    .A(\hn5.hidden_neuron_o[0] ),
    .B(_0137_));
 sg13g2_a21oi_1 _0597_ (.A1(\hn2.hidden_neuron_o[0] ),
    .A2(_0133_),
    .Y(_0140_),
    .B1(_0132_));
 sg13g2_xor2_1 _0598_ (.B(\hn2.hidden_neuron_o[0] ),
    .A(\hn2.hidden_neuron_o[1] ),
    .X(_0141_));
 sg13g2_nand2_1 _0599_ (.Y(_0142_),
    .A(\hn1.hidden_neuron_o[0] ),
    .B(\hn0.hidden_neuron_o[1] ));
 sg13g2_xor2_1 _0600_ (.B(\hn0.hidden_neuron_o[1] ),
    .A(\hn1.hidden_neuron_o[0] ),
    .X(_0143_));
 sg13g2_xnor2_1 _0601_ (.Y(_0144_),
    .A(_0001_),
    .B(_0143_));
 sg13g2_and2_1 _0602_ (.A(_0141_),
    .B(_0144_),
    .X(_0145_));
 sg13g2_xor2_1 _0603_ (.B(_0144_),
    .A(_0141_),
    .X(_0146_));
 sg13g2_inv_1 _0604_ (.Y(_0147_),
    .A(_0146_));
 sg13g2_xnor2_1 _0605_ (.Y(_0148_),
    .A(_0140_),
    .B(_0146_));
 sg13g2_nand2b_1 _0606_ (.Y(_0149_),
    .B(_0148_),
    .A_N(_0139_));
 sg13g2_xnor2_1 _0607_ (.Y(_0150_),
    .A(_0139_),
    .B(_0148_));
 sg13g2_nand2_1 _0608_ (.Y(_0151_),
    .A(_0135_),
    .B(_0150_));
 sg13g2_xnor2_1 _0609_ (.Y(_0152_),
    .A(_0135_),
    .B(_0150_));
 sg13g2_nor2_1 _0610_ (.A(net88),
    .B(net61),
    .Y(_0153_));
 sg13g2_a21oi_1 _0611_ (.A1(net88),
    .A2(_0152_),
    .Y(_0024_),
    .B1(_0153_));
 sg13g2_o21ai_1 _0612_ (.B1(_0149_),
    .Y(_0154_),
    .A1(_0140_),
    .A2(_0147_));
 sg13g2_xor2_1 _0613_ (.B(\hn5.hidden_neuron_o[0] ),
    .A(\hn5.hidden_neuron_o[1] ),
    .X(_0155_));
 sg13g2_nand2_1 _0614_ (.Y(_0156_),
    .A(\hn6.hidden_neuron_o[2] ),
    .B(\hn6.hidden_neuron_o[1] ));
 sg13g2_nor2_1 _0615_ (.A(\hn6.hidden_neuron_o[2] ),
    .B(\hn6.hidden_neuron_o[1] ),
    .Y(_0157_));
 sg13g2_nor2_1 _0616_ (.A(\hn6.hidden_neuron_o[0] ),
    .B(_0157_),
    .Y(_0158_));
 sg13g2_a22oi_1 _0617_ (.Y(_0159_),
    .B1(_0156_),
    .B2(_0158_),
    .A2(\hn6.hidden_neuron_o[0] ),
    .A1(_0059_));
 sg13g2_nor2b_1 _0618_ (.A(\hn2.hidden_neuron_o[0] ),
    .B_N(\hn2.hidden_neuron_o[1] ),
    .Y(_0160_));
 sg13g2_xnor2_1 _0619_ (.Y(_0161_),
    .A(\hn2.hidden_neuron_o[2] ),
    .B(_0160_));
 sg13g2_xor2_1 _0620_ (.B(_0161_),
    .A(_0159_),
    .X(_0162_));
 sg13g2_nand2_1 _0621_ (.Y(_0163_),
    .A(_0155_),
    .B(_0162_));
 sg13g2_xnor2_1 _0622_ (.Y(_0164_),
    .A(_0155_),
    .B(_0162_));
 sg13g2_a21oi_1 _0623_ (.A1(_0064_),
    .A2(_0143_),
    .Y(_0165_),
    .B1(_0145_));
 sg13g2_nand2_1 _0624_ (.Y(_0166_),
    .A(\hn4.hidden_neuron_o[2] ),
    .B(\hn4.hidden_neuron_o[0] ));
 sg13g2_xor2_1 _0625_ (.B(\hn4.hidden_neuron_o[0] ),
    .A(\hn4.hidden_neuron_o[2] ),
    .X(_0167_));
 sg13g2_nand2_1 _0626_ (.Y(_0168_),
    .A(\hn1.hidden_neuron_o[1] ),
    .B(\hn0.hidden_neuron_o[2] ));
 sg13g2_xnor2_1 _0627_ (.Y(_0169_),
    .A(\hn1.hidden_neuron_o[1] ),
    .B(\hn0.hidden_neuron_o[2] ));
 sg13g2_xor2_1 _0628_ (.B(_0169_),
    .A(_0142_),
    .X(_0170_));
 sg13g2_xnor2_1 _0629_ (.Y(_0171_),
    .A(_0002_),
    .B(_0170_));
 sg13g2_and2_1 _0630_ (.A(_0167_),
    .B(_0171_),
    .X(_0172_));
 sg13g2_xnor2_1 _0631_ (.Y(_0173_),
    .A(_0167_),
    .B(_0171_));
 sg13g2_nor2_1 _0632_ (.A(_0165_),
    .B(_0173_),
    .Y(_0174_));
 sg13g2_xnor2_1 _0633_ (.Y(_0175_),
    .A(_0165_),
    .B(_0173_));
 sg13g2_nor2_1 _0634_ (.A(_0164_),
    .B(_0175_),
    .Y(_0176_));
 sg13g2_xor2_1 _0635_ (.B(_0175_),
    .A(_0164_),
    .X(_0177_));
 sg13g2_nand2_1 _0636_ (.Y(_0178_),
    .A(_0154_),
    .B(_0177_));
 sg13g2_xnor2_1 _0637_ (.Y(_0179_),
    .A(_0154_),
    .B(_0177_));
 sg13g2_xor2_1 _0638_ (.B(_0179_),
    .A(_0138_),
    .X(_0180_));
 sg13g2_nand2b_1 _0639_ (.Y(_0181_),
    .B(_0180_),
    .A_N(_0151_));
 sg13g2_xnor2_1 _0640_ (.Y(_0182_),
    .A(_0151_),
    .B(_0180_));
 sg13g2_mux2_1 _0641_ (.A0(net69),
    .A1(_0182_),
    .S(net88),
    .X(_0025_));
 sg13g2_nand2_1 _0642_ (.Y(_0183_),
    .A(net82),
    .B(net60));
 sg13g2_o21ai_1 _0643_ (.B1(_0178_),
    .Y(_0184_),
    .A1(_0138_),
    .A2(_0179_));
 sg13g2_o21ai_1 _0644_ (.B1(_0163_),
    .Y(_0185_),
    .A1(_0159_),
    .A2(_0161_));
 sg13g2_nor2_1 _0645_ (.A(_0174_),
    .B(_0176_),
    .Y(_0186_));
 sg13g2_a21oi_2 _0646_ (.B1(_0172_),
    .Y(_0187_),
    .A2(_0170_),
    .A1(_0065_));
 sg13g2_nand2_1 _0647_ (.Y(_0188_),
    .A(\hn4.hidden_neuron_o[3] ),
    .B(\hn4.hidden_neuron_o[1] ));
 sg13g2_xnor2_1 _0648_ (.Y(_0189_),
    .A(\hn4.hidden_neuron_o[3] ),
    .B(\hn4.hidden_neuron_o[1] ));
 sg13g2_xnor2_1 _0649_ (.Y(_0190_),
    .A(_0166_),
    .B(_0189_));
 sg13g2_o21ai_1 _0650_ (.B1(_0168_),
    .Y(_0191_),
    .A1(_0142_),
    .A2(_0169_));
 sg13g2_and2_1 _0651_ (.A(\hn1.hidden_neuron_o[2] ),
    .B(\hn0.hidden_neuron_o[3] ),
    .X(_0192_));
 sg13g2_or2_1 _0652_ (.X(_0193_),
    .B(\hn0.hidden_neuron_o[3] ),
    .A(\hn1.hidden_neuron_o[2] ));
 sg13g2_nand2b_1 _0653_ (.Y(_0194_),
    .B(_0193_),
    .A_N(_0192_));
 sg13g2_xnor2_1 _0654_ (.Y(_0195_),
    .A(_0191_),
    .B(_0194_));
 sg13g2_nand2_1 _0655_ (.Y(_0196_),
    .A(\hn3.hidden_neuron_o[1] ),
    .B(_0195_));
 sg13g2_xnor2_1 _0656_ (.Y(_0197_),
    .A(\hn3.hidden_neuron_o[1] ),
    .B(_0195_));
 sg13g2_xnor2_1 _0657_ (.Y(_0198_),
    .A(_0190_),
    .B(_0197_));
 sg13g2_nor2_1 _0658_ (.A(_0187_),
    .B(_0198_),
    .Y(_0199_));
 sg13g2_xor2_1 _0659_ (.B(_0198_),
    .A(_0187_),
    .X(_0200_));
 sg13g2_nand2b_1 _0660_ (.Y(_0201_),
    .B(\hn5.hidden_neuron_o[1] ),
    .A_N(\hn5.hidden_neuron_o[0] ));
 sg13g2_xor2_1 _0661_ (.B(_0201_),
    .A(\hn5.hidden_neuron_o[2] ),
    .X(_0202_));
 sg13g2_a21oi_1 _0662_ (.A1(\hn2.hidden_neuron_o[1] ),
    .A2(\hn2.hidden_neuron_o[0] ),
    .Y(_0203_),
    .B1(\hn2.hidden_neuron_o[2] ));
 sg13g2_a21oi_1 _0663_ (.A1(\hn2.hidden_neuron_o[2] ),
    .A2(\hn2.hidden_neuron_o[1] ),
    .Y(_0204_),
    .B1(_0203_));
 sg13g2_xnor2_1 _0664_ (.Y(_0205_),
    .A(\hn2.hidden_neuron_o[3] ),
    .B(_0204_));
 sg13g2_xnor2_1 _0665_ (.Y(_0206_),
    .A(\hn6.hidden_neuron_o[3] ),
    .B(_0158_));
 sg13g2_xor2_1 _0666_ (.B(_0206_),
    .A(_0205_),
    .X(_0207_));
 sg13g2_nand2b_1 _0667_ (.Y(_0208_),
    .B(_0207_),
    .A_N(_0202_));
 sg13g2_xnor2_1 _0668_ (.Y(_0209_),
    .A(_0202_),
    .B(_0207_));
 sg13g2_xnor2_1 _0669_ (.Y(_0210_),
    .A(_0200_),
    .B(_0209_));
 sg13g2_nor2_1 _0670_ (.A(_0186_),
    .B(_0210_),
    .Y(_0211_));
 sg13g2_xor2_1 _0671_ (.B(_0210_),
    .A(_0186_),
    .X(_0212_));
 sg13g2_xnor2_1 _0672_ (.Y(_0213_),
    .A(_0185_),
    .B(_0212_));
 sg13g2_nand2b_1 _0673_ (.Y(_0214_),
    .B(_0184_),
    .A_N(_0213_));
 sg13g2_xnor2_1 _0674_ (.Y(_0215_),
    .A(_0184_),
    .B(_0213_));
 sg13g2_nand2_1 _0675_ (.Y(_0216_),
    .A(\hn7.hidden_neuron_o[0] ),
    .B(_0215_));
 sg13g2_xnor2_1 _0676_ (.Y(_0217_),
    .A(\hn7.hidden_neuron_o[0] ),
    .B(_0215_));
 sg13g2_nor2_2 _0677_ (.A(_0181_),
    .B(_0217_),
    .Y(_0218_));
 sg13g2_a21o_1 _0678_ (.A2(_0217_),
    .A1(_0181_),
    .B1(net82),
    .X(_0219_));
 sg13g2_o21ai_1 _0679_ (.B1(_0183_),
    .Y(_0026_),
    .A1(_0218_),
    .A2(_0219_));
 sg13g2_a21oi_1 _0680_ (.A1(_0185_),
    .A2(_0212_),
    .Y(_0220_),
    .B1(_0211_));
 sg13g2_o21ai_1 _0681_ (.B1(_0208_),
    .Y(_0221_),
    .A1(_0205_),
    .A2(_0206_));
 sg13g2_a21oi_1 _0682_ (.A1(_0200_),
    .A2(_0209_),
    .Y(_0222_),
    .B1(_0199_));
 sg13g2_nand2b_2 _0683_ (.Y(_0223_),
    .B(\hn2.hidden_neuron_o[3] ),
    .A_N(_0203_));
 sg13g2_a21o_1 _0684_ (.A2(\hn2.hidden_neuron_o[1] ),
    .A1(\hn2.hidden_neuron_o[2] ),
    .B1(\hn2.hidden_neuron_o[3] ),
    .X(_0224_));
 sg13g2_and2_1 _0685_ (.A(_0223_),
    .B(_0224_),
    .X(_0225_));
 sg13g2_nor2_1 _0686_ (.A(\hn6.hidden_neuron_o[4] ),
    .B(\hn6.hidden_neuron_o[3] ),
    .Y(_0226_));
 sg13g2_nand2_1 _0687_ (.Y(_0227_),
    .A(\hn6.hidden_neuron_o[4] ),
    .B(\hn6.hidden_neuron_o[3] ));
 sg13g2_nand2_1 _0688_ (.Y(_0228_),
    .A(\hn6.hidden_neuron_o[4] ),
    .B(_0058_));
 sg13g2_xor2_1 _0689_ (.B(\hn6.hidden_neuron_o[3] ),
    .A(\hn6.hidden_neuron_o[4] ),
    .X(_0229_));
 sg13g2_xnor2_1 _0690_ (.Y(_0230_),
    .A(\hn6.hidden_neuron_o[2] ),
    .B(_0229_));
 sg13g2_o21ai_1 _0691_ (.B1(_0156_),
    .Y(_0231_),
    .A1(_0058_),
    .A2(_0157_));
 sg13g2_nor2b_1 _0692_ (.A(_0230_),
    .B_N(_0231_),
    .Y(_0232_));
 sg13g2_xnor2_1 _0693_ (.Y(_0233_),
    .A(_0230_),
    .B(_0231_));
 sg13g2_nand2b_1 _0694_ (.Y(_0234_),
    .B(\hn6.hidden_neuron_o[0] ),
    .A_N(\hn6.hidden_neuron_o[3] ));
 sg13g2_nand3_1 _0695_ (.B(\hn6.hidden_neuron_o[2] ),
    .C(\hn6.hidden_neuron_o[1] ),
    .A(\hn6.hidden_neuron_o[3] ),
    .Y(_0235_));
 sg13g2_o21ai_1 _0696_ (.B1(_0235_),
    .Y(_0236_),
    .A1(_0157_),
    .A2(_0234_));
 sg13g2_xor2_1 _0697_ (.B(_0236_),
    .A(_0233_),
    .X(_0237_));
 sg13g2_nand2_1 _0698_ (.Y(_0238_),
    .A(_0225_),
    .B(_0237_));
 sg13g2_xnor2_1 _0699_ (.Y(_0239_),
    .A(_0225_),
    .B(_0237_));
 sg13g2_a21oi_1 _0700_ (.A1(\hn5.hidden_neuron_o[1] ),
    .A2(\hn5.hidden_neuron_o[0] ),
    .Y(_0240_),
    .B1(\hn5.hidden_neuron_o[2] ));
 sg13g2_a21oi_1 _0701_ (.A1(\hn5.hidden_neuron_o[2] ),
    .A2(\hn5.hidden_neuron_o[1] ),
    .Y(_0241_),
    .B1(_0240_));
 sg13g2_xnor2_1 _0702_ (.Y(_0242_),
    .A(\hn5.hidden_neuron_o[3] ),
    .B(_0241_));
 sg13g2_xor2_1 _0703_ (.B(_0242_),
    .A(_0239_),
    .X(_0243_));
 sg13g2_inv_1 _0704_ (.Y(_0244_),
    .A(_0243_));
 sg13g2_o21ai_1 _0705_ (.B1(_0196_),
    .Y(_0245_),
    .A1(_0190_),
    .A2(_0197_));
 sg13g2_and2_1 _0706_ (.A(\hn4.hidden_neuron_o[4] ),
    .B(\hn4.hidden_neuron_o[2] ),
    .X(_0246_));
 sg13g2_or2_1 _0707_ (.X(_0247_),
    .B(\hn4.hidden_neuron_o[2] ),
    .A(\hn4.hidden_neuron_o[4] ));
 sg13g2_nand2b_1 _0708_ (.Y(_0248_),
    .B(_0247_),
    .A_N(_0246_));
 sg13g2_o21ai_1 _0709_ (.B1(_0188_),
    .Y(_0249_),
    .A1(_0166_),
    .A2(_0189_));
 sg13g2_nand2b_1 _0710_ (.Y(_0250_),
    .B(_0249_),
    .A_N(_0248_));
 sg13g2_xnor2_1 _0711_ (.Y(_0251_),
    .A(_0248_),
    .B(_0249_));
 sg13g2_a21o_2 _0712_ (.A2(_0193_),
    .A1(_0191_),
    .B1(_0192_),
    .X(_0252_));
 sg13g2_nand2_1 _0713_ (.Y(_0253_),
    .A(\hn1.hidden_neuron_o[3] ),
    .B(_0252_));
 sg13g2_xor2_1 _0714_ (.B(_0252_),
    .A(\hn1.hidden_neuron_o[3] ),
    .X(_0254_));
 sg13g2_nor2b_1 _0715_ (.A(_0003_),
    .B_N(_0254_),
    .Y(_0255_));
 sg13g2_xnor2_1 _0716_ (.Y(_0256_),
    .A(_0003_),
    .B(_0254_));
 sg13g2_xor2_1 _0717_ (.B(_0256_),
    .A(_0251_),
    .X(_0257_));
 sg13g2_nand2_1 _0718_ (.Y(_0258_),
    .A(_0245_),
    .B(_0257_));
 sg13g2_xnor2_1 _0719_ (.Y(_0259_),
    .A(_0245_),
    .B(_0257_));
 sg13g2_xnor2_1 _0720_ (.Y(_0260_),
    .A(_0244_),
    .B(_0259_));
 sg13g2_nor2_1 _0721_ (.A(_0222_),
    .B(_0260_),
    .Y(_0261_));
 sg13g2_xor2_1 _0722_ (.B(_0260_),
    .A(_0222_),
    .X(_0262_));
 sg13g2_xnor2_1 _0723_ (.Y(_0263_),
    .A(_0221_),
    .B(_0262_));
 sg13g2_xor2_1 _0724_ (.B(_0263_),
    .A(_0220_),
    .X(_0264_));
 sg13g2_nand2_1 _0725_ (.Y(_0265_),
    .A(\hn7.hidden_neuron_o[1] ),
    .B(_0264_));
 sg13g2_xnor2_1 _0726_ (.Y(_0266_),
    .A(\hn7.hidden_neuron_o[1] ),
    .B(_0264_));
 sg13g2_a21oi_1 _0727_ (.A1(_0214_),
    .A2(_0216_),
    .Y(_0267_),
    .B1(_0266_));
 sg13g2_nand3_1 _0728_ (.B(_0216_),
    .C(_0266_),
    .A(_0214_),
    .Y(_0268_));
 sg13g2_nand2b_1 _0729_ (.Y(_0269_),
    .B(_0268_),
    .A_N(_0267_));
 sg13g2_xor2_1 _0730_ (.B(_0269_),
    .A(_0218_),
    .X(_0270_));
 sg13g2_nor2_1 _0731_ (.A(net88),
    .B(net58),
    .Y(_0271_));
 sg13g2_a21oi_1 _0732_ (.A1(net88),
    .A2(_0270_),
    .Y(_0027_),
    .B1(_0271_));
 sg13g2_a21oi_1 _0733_ (.A1(_0218_),
    .A2(_0268_),
    .Y(_0272_),
    .B1(_0267_));
 sg13g2_o21ai_1 _0734_ (.B1(_0265_),
    .Y(_0273_),
    .A1(_0220_),
    .A2(_0263_));
 sg13g2_a21oi_2 _0735_ (.B1(_0261_),
    .Y(_0274_),
    .A2(_0262_),
    .A1(_0221_));
 sg13g2_o21ai_1 _0736_ (.B1(_0238_),
    .Y(_0275_),
    .A1(_0239_),
    .A2(_0242_));
 sg13g2_o21ai_1 _0737_ (.B1(_0258_),
    .Y(_0276_),
    .A1(_0244_),
    .A2(_0259_));
 sg13g2_a21oi_1 _0738_ (.A1(_0251_),
    .A2(_0256_),
    .Y(_0277_),
    .B1(_0255_));
 sg13g2_nand3_1 _0739_ (.B(_0066_),
    .C(_0252_),
    .A(\hn1.hidden_neuron_o[3] ),
    .Y(_0278_));
 sg13g2_a21oi_1 _0740_ (.A1(\hn1.hidden_neuron_o[3] ),
    .A2(_0252_),
    .Y(_0279_),
    .B1(_0066_));
 sg13g2_xnor2_1 _0741_ (.Y(_0280_),
    .A(_0004_),
    .B(_0253_));
 sg13g2_a21oi_1 _0742_ (.A1(_0247_),
    .A2(_0249_),
    .Y(_0281_),
    .B1(_0246_));
 sg13g2_xnor2_1 _0743_ (.Y(_0282_),
    .A(_0005_),
    .B(_0281_));
 sg13g2_xnor2_1 _0744_ (.Y(_0283_),
    .A(_0280_),
    .B(_0282_));
 sg13g2_nor2_1 _0745_ (.A(_0277_),
    .B(_0283_),
    .Y(_0284_));
 sg13g2_xor2_1 _0746_ (.B(_0283_),
    .A(_0277_),
    .X(_0285_));
 sg13g2_a21oi_1 _0747_ (.A1(\hn5.hidden_neuron_o[2] ),
    .A2(\hn5.hidden_neuron_o[1] ),
    .Y(_0286_),
    .B1(\hn5.hidden_neuron_o[3] ));
 sg13g2_nor2_1 _0748_ (.A(_0240_),
    .B(_0286_),
    .Y(_0287_));
 sg13g2_xor2_1 _0749_ (.B(\hn5.hidden_neuron_o[3] ),
    .A(\hn5.hidden_neuron_o[4] ),
    .X(_0288_));
 sg13g2_xnor2_1 _0750_ (.Y(_0289_),
    .A(_0287_),
    .B(_0288_));
 sg13g2_a21oi_1 _0751_ (.A1(_0233_),
    .A2(_0236_),
    .Y(_0290_),
    .B1(_0232_));
 sg13g2_a21oi_1 _0752_ (.A1(\hn6.hidden_neuron_o[2] ),
    .A2(_0227_),
    .Y(_0291_),
    .B1(_0226_));
 sg13g2_xor2_1 _0753_ (.B(_0291_),
    .A(_0290_),
    .X(_0292_));
 sg13g2_xor2_1 _0754_ (.B(_0292_),
    .A(_0223_),
    .X(_0293_));
 sg13g2_nand2b_1 _0755_ (.Y(_0294_),
    .B(_0293_),
    .A_N(_0289_));
 sg13g2_xnor2_1 _0756_ (.Y(_0295_),
    .A(_0289_),
    .B(_0293_));
 sg13g2_xnor2_1 _0757_ (.Y(_0296_),
    .A(_0285_),
    .B(_0295_));
 sg13g2_nor2b_1 _0758_ (.A(_0296_),
    .B_N(_0276_),
    .Y(_0297_));
 sg13g2_xnor2_1 _0759_ (.Y(_0298_),
    .A(_0276_),
    .B(_0296_));
 sg13g2_xnor2_1 _0760_ (.Y(_0299_),
    .A(_0275_),
    .B(_0298_));
 sg13g2_nor2_1 _0761_ (.A(_0274_),
    .B(_0299_),
    .Y(_0300_));
 sg13g2_xor2_1 _0762_ (.B(_0299_),
    .A(_0274_),
    .X(_0301_));
 sg13g2_xnor2_1 _0763_ (.Y(_0302_),
    .A(\hn7.hidden_neuron_o[2] ),
    .B(_0301_));
 sg13g2_inv_1 _0764_ (.Y(_0303_),
    .A(_0302_));
 sg13g2_nor2_2 _0765_ (.A(_0273_),
    .B(_0303_),
    .Y(_0304_));
 sg13g2_xor2_1 _0766_ (.B(_0302_),
    .A(_0273_),
    .X(_0305_));
 sg13g2_xor2_1 _0767_ (.B(_0305_),
    .A(_0272_),
    .X(_0306_));
 sg13g2_a221oi_1 _0768_ (.B2(_0303_),
    .C1(_0267_),
    .B1(_0273_),
    .A1(_0218_),
    .Y(_0307_),
    .A2(_0268_));
 sg13g2_mux2_1 _0769_ (.A0(net66),
    .A1(_0306_),
    .S(net87),
    .X(_0028_));
 sg13g2_a21oi_2 _0770_ (.B1(_0297_),
    .Y(_0308_),
    .A2(_0298_),
    .A1(_0275_));
 sg13g2_o21ai_1 _0771_ (.B1(_0294_),
    .Y(_0309_),
    .A1(_0223_),
    .A2(_0292_));
 sg13g2_a21oi_1 _0772_ (.A1(_0285_),
    .A2(_0295_),
    .Y(_0310_),
    .B1(_0284_));
 sg13g2_nor2b_2 _0773_ (.A(_0286_),
    .B_N(\hn5.hidden_neuron_o[4] ),
    .Y(_0311_));
 sg13g2_a21oi_1 _0774_ (.A1(\hn5.hidden_neuron_o[3] ),
    .A2(_0287_),
    .Y(_0312_),
    .B1(\hn5.hidden_neuron_o[4] ));
 sg13g2_nor2_1 _0775_ (.A(_0311_),
    .B(_0312_),
    .Y(_0313_));
 sg13g2_nand3b_1 _0776_ (.B(_0231_),
    .C(_0291_),
    .Y(_0314_),
    .A_N(_0230_));
 sg13g2_a22oi_1 _0777_ (.Y(_0315_),
    .B1(_0236_),
    .B2(\hn6.hidden_neuron_o[4] ),
    .A2(_0229_),
    .A1(\hn6.hidden_neuron_o[2] ));
 sg13g2_nand2_1 _0778_ (.Y(_0316_),
    .A(_0314_),
    .B(_0315_));
 sg13g2_xor2_1 _0779_ (.B(_0316_),
    .A(_0228_),
    .X(_0317_));
 sg13g2_or3_1 _0780_ (.A(_0311_),
    .B(_0312_),
    .C(_0317_),
    .X(_0318_));
 sg13g2_xor2_1 _0781_ (.B(_0317_),
    .A(_0313_),
    .X(_0319_));
 sg13g2_nor2_1 _0782_ (.A(_0005_),
    .B(_0250_),
    .Y(_0320_));
 sg13g2_nor4_1 _0783_ (.A(_0055_),
    .B(\hn4.hidden_neuron_o[2] ),
    .C(_0005_),
    .D(_0188_),
    .Y(_0321_));
 sg13g2_a21oi_2 _0784_ (.B1(_0321_),
    .Y(_0322_),
    .A2(_0246_),
    .A1(\hn4.hidden_neuron_o[3] ));
 sg13g2_o21ai_1 _0785_ (.B1(_0322_),
    .Y(_0323_),
    .A1(\hn4.hidden_neuron_o[4] ),
    .A2(_0320_));
 sg13g2_o21ai_1 _0786_ (.B1(_0278_),
    .Y(_0324_),
    .A1(_0279_),
    .A2(_0282_));
 sg13g2_nor2b_1 _0787_ (.A(_0323_),
    .B_N(_0324_),
    .Y(_0325_));
 sg13g2_xor2_1 _0788_ (.B(_0324_),
    .A(_0323_),
    .X(_0326_));
 sg13g2_nor2_1 _0789_ (.A(_0319_),
    .B(_0326_),
    .Y(_0327_));
 sg13g2_xnor2_1 _0790_ (.Y(_0328_),
    .A(_0319_),
    .B(_0326_));
 sg13g2_nor2_1 _0791_ (.A(_0310_),
    .B(_0328_),
    .Y(_0329_));
 sg13g2_xor2_1 _0792_ (.B(_0328_),
    .A(_0310_),
    .X(_0330_));
 sg13g2_xnor2_1 _0793_ (.Y(_0331_),
    .A(_0309_),
    .B(_0330_));
 sg13g2_nor2_1 _0794_ (.A(_0308_),
    .B(_0331_),
    .Y(_0332_));
 sg13g2_xor2_1 _0795_ (.B(_0331_),
    .A(_0308_),
    .X(_0333_));
 sg13g2_xnor2_1 _0796_ (.Y(_0334_),
    .A(\hn7.hidden_neuron_o[3] ),
    .B(_0333_));
 sg13g2_a21oi_1 _0797_ (.A1(\hn7.hidden_neuron_o[2] ),
    .A2(_0301_),
    .Y(_0335_),
    .B1(_0300_));
 sg13g2_nor2_1 _0798_ (.A(_0334_),
    .B(_0335_),
    .Y(_0336_));
 sg13g2_xnor2_1 _0799_ (.Y(_0337_),
    .A(_0334_),
    .B(_0335_));
 sg13g2_nor3_1 _0800_ (.A(_0304_),
    .B(_0307_),
    .C(_0337_),
    .Y(_0338_));
 sg13g2_o21ai_1 _0801_ (.B1(_0337_),
    .Y(_0339_),
    .A1(_0304_),
    .A2(_0307_));
 sg13g2_nand2_1 _0802_ (.Y(_0340_),
    .A(net82),
    .B(net62));
 sg13g2_nand2_1 _0803_ (.Y(_0341_),
    .A(net87),
    .B(_0339_));
 sg13g2_o21ai_1 _0804_ (.B1(_0340_),
    .Y(_0029_),
    .A1(_0338_),
    .A2(_0341_));
 sg13g2_a21oi_2 _0805_ (.B1(_0332_),
    .Y(_0342_),
    .A2(_0333_),
    .A1(\hn7.hidden_neuron_o[3] ));
 sg13g2_a21oi_2 _0806_ (.B1(_0329_),
    .Y(_0343_),
    .A2(_0330_),
    .A1(_0309_));
 sg13g2_nor2_1 _0807_ (.A(_0325_),
    .B(_0327_),
    .Y(_0344_));
 sg13g2_o21ai_1 _0808_ (.B1(\hn6.hidden_neuron_o[4] ),
    .Y(_0345_),
    .A1(\hn6.hidden_neuron_o[3] ),
    .A2(_0316_));
 sg13g2_nand2b_1 _0809_ (.Y(_0346_),
    .B(_0311_),
    .A_N(_0345_));
 sg13g2_xor2_1 _0810_ (.B(_0345_),
    .A(_0311_),
    .X(_0347_));
 sg13g2_xor2_1 _0811_ (.B(_0347_),
    .A(_0322_),
    .X(_0348_));
 sg13g2_o21ai_1 _0812_ (.B1(_0348_),
    .Y(_0349_),
    .A1(_0325_),
    .A2(_0327_));
 sg13g2_xnor2_1 _0813_ (.Y(_0350_),
    .A(_0344_),
    .B(_0348_));
 sg13g2_nand2b_1 _0814_ (.Y(_0351_),
    .B(_0350_),
    .A_N(_0318_));
 sg13g2_xnor2_1 _0815_ (.Y(_0352_),
    .A(_0318_),
    .B(_0350_));
 sg13g2_nand2b_1 _0816_ (.Y(_0353_),
    .B(_0352_),
    .A_N(_0343_));
 sg13g2_xnor2_1 _0817_ (.Y(_0354_),
    .A(_0343_),
    .B(_0352_));
 sg13g2_nand2_1 _0818_ (.Y(_0355_),
    .A(\hn7.hidden_neuron_o[4] ),
    .B(_0354_));
 sg13g2_xnor2_1 _0819_ (.Y(_0356_),
    .A(\hn7.hidden_neuron_o[4] ),
    .B(_0354_));
 sg13g2_nand2_1 _0820_ (.Y(_0357_),
    .A(_0342_),
    .B(_0356_));
 sg13g2_xor2_1 _0821_ (.B(_0356_),
    .A(_0342_),
    .X(_0358_));
 sg13g2_inv_1 _0822_ (.Y(_0359_),
    .A(_0358_));
 sg13g2_nor2_1 _0823_ (.A(_0336_),
    .B(_0338_),
    .Y(_0360_));
 sg13g2_xnor2_1 _0824_ (.Y(_0361_),
    .A(_0359_),
    .B(_0360_));
 sg13g2_nor2_1 _0825_ (.A(net87),
    .B(net63),
    .Y(_0362_));
 sg13g2_a21oi_1 _0826_ (.A1(net87),
    .A2(_0361_),
    .Y(_0030_),
    .B1(_0362_));
 sg13g2_nand2_1 _0827_ (.Y(_0363_),
    .A(net81),
    .B(net67));
 sg13g2_o21ai_1 _0828_ (.B1(_0346_),
    .Y(_0364_),
    .A1(_0322_),
    .A2(_0347_));
 sg13g2_nand2_1 _0829_ (.Y(_0365_),
    .A(_0349_),
    .B(_0351_));
 sg13g2_xnor2_1 _0830_ (.Y(_0366_),
    .A(_0364_),
    .B(_0365_));
 sg13g2_and3_1 _0831_ (.X(_0367_),
    .A(_0353_),
    .B(_0355_),
    .C(_0366_));
 sg13g2_a21oi_1 _0832_ (.A1(_0353_),
    .A2(_0355_),
    .Y(_0368_),
    .B1(_0366_));
 sg13g2_nor2_1 _0833_ (.A(_0367_),
    .B(_0368_),
    .Y(_0369_));
 sg13g2_nor4_2 _0834_ (.A(_0304_),
    .B(_0307_),
    .C(_0337_),
    .Y(_0370_),
    .D(_0359_));
 sg13g2_nand2_1 _0835_ (.Y(_0371_),
    .A(_0336_),
    .B(_0357_));
 sg13g2_o21ai_1 _0836_ (.B1(_0371_),
    .Y(_0372_),
    .A1(_0342_),
    .A2(_0356_));
 sg13g2_nor3_1 _0837_ (.A(_0369_),
    .B(_0370_),
    .C(_0372_),
    .Y(_0373_));
 sg13g2_o21ai_1 _0838_ (.B1(_0369_),
    .Y(_0374_),
    .A1(_0370_),
    .A2(_0372_));
 sg13g2_nand2_1 _0839_ (.Y(_0375_),
    .A(net87),
    .B(_0374_));
 sg13g2_o21ai_1 _0840_ (.B1(_0363_),
    .Y(_0031_),
    .A1(_0373_),
    .A2(_0375_));
 sg13g2_a21oi_1 _0841_ (.A1(_0364_),
    .A2(_0365_),
    .Y(_0376_),
    .B1(_0368_));
 sg13g2_a21oi_1 _0842_ (.A1(_0374_),
    .A2(_0376_),
    .Y(_0377_),
    .B1(net81));
 sg13g2_a21o_1 _0843_ (.A2(net78),
    .A1(net81),
    .B1(_0377_),
    .X(_0032_));
 sg13g2_nor2b_1 _0844_ (.A(net87),
    .B_N(net56),
    .Y(_0033_));
 sg13g2_nand2_1 _0845_ (.Y(_0378_),
    .A(net85),
    .B(net73));
 sg13g2_a21oi_1 _0846_ (.A1(_0107_),
    .A2(_0378_),
    .Y(_0034_),
    .B1(net95));
 sg13g2_nand2_1 _0847_ (.Y(_0379_),
    .A(net84),
    .B(net68));
 sg13g2_nand2_1 _0848_ (.Y(_0380_),
    .A(_0087_),
    .B(_0122_));
 sg13g2_o21ai_1 _0849_ (.B1(_0086_),
    .Y(_0381_),
    .A1(net101),
    .A2(_0380_));
 sg13g2_nand2_1 _0850_ (.Y(_0382_),
    .A(net91),
    .B(_0381_));
 sg13g2_a21oi_1 _0851_ (.A1(_0379_),
    .A2(_0382_),
    .Y(_0035_),
    .B1(net95));
 sg13g2_nor3_1 _0852_ (.A(_0080_),
    .B(_0084_),
    .C(_0085_),
    .Y(_0383_));
 sg13g2_o21ai_1 _0853_ (.B1(net104),
    .Y(_0384_),
    .A1(net84),
    .A2(_0383_));
 sg13g2_a21oi_1 _0854_ (.A1(net84),
    .A2(_0057_),
    .Y(_0036_),
    .B1(_0384_));
 sg13g2_a22oi_1 _0855_ (.Y(_0385_),
    .B1(_0072_),
    .B2(_0082_),
    .A2(net72),
    .A1(net86));
 sg13g2_nor2_1 _0856_ (.A(net94),
    .B(_0385_),
    .Y(_0037_));
 sg13g2_nand2_1 _0857_ (.Y(_0386_),
    .A(net84),
    .B(net77));
 sg13g2_a21oi_1 _0858_ (.A1(_0069_),
    .A2(_0386_),
    .Y(_0038_),
    .B1(net95));
 sg13g2_nand2_1 _0859_ (.Y(_0387_),
    .A(net85),
    .B(net74));
 sg13g2_a21oi_1 _0860_ (.A1(_0077_),
    .A2(_0387_),
    .Y(_0039_),
    .B1(net95));
 sg13g2_o21ai_1 _0861_ (.B1(net89),
    .Y(_0388_),
    .A1(_0073_),
    .A2(_0122_));
 sg13g2_a21oi_1 _0862_ (.A1(net99),
    .A2(_0074_),
    .Y(_0389_),
    .B1(net98));
 sg13g2_nor2_1 _0863_ (.A(net83),
    .B(_0111_),
    .Y(_0390_));
 sg13g2_nor2_1 _0864_ (.A(_0388_),
    .B(_0389_),
    .Y(_0391_));
 sg13g2_a21oi_1 _0865_ (.A1(net83),
    .A2(net71),
    .Y(_0392_),
    .B1(_0391_));
 sg13g2_nor2_1 _0866_ (.A(net94),
    .B(_0392_),
    .Y(_0040_));
 sg13g2_o21ai_1 _0867_ (.B1(net104),
    .Y(_0393_),
    .A1(net89),
    .A2(net122));
 sg13g2_nor2b_1 _0868_ (.A(_0393_),
    .B_N(_0388_),
    .Y(_0041_));
 sg13g2_nand2_1 _0869_ (.Y(_0394_),
    .A(net85),
    .B(net118));
 sg13g2_a21oi_1 _0870_ (.A1(_0107_),
    .A2(_0394_),
    .Y(_0042_),
    .B1(net93));
 sg13g2_nand2_1 _0871_ (.Y(_0395_),
    .A(net85),
    .B(net113));
 sg13g2_a21oi_1 _0872_ (.A1(_0109_),
    .A2(_0395_),
    .Y(_0043_),
    .B1(net93));
 sg13g2_o21ai_1 _0873_ (.B1(net104),
    .Y(_0396_),
    .A1(net92),
    .A2(net121));
 sg13g2_a21oi_1 _0874_ (.A1(net90),
    .A2(_0117_),
    .Y(_0044_),
    .B1(_0396_));
 sg13g2_nand2_1 _0875_ (.Y(_0397_),
    .A(net83),
    .B(net108));
 sg13g2_a21oi_1 _0876_ (.A1(_0095_),
    .A2(_0397_),
    .Y(_0045_),
    .B1(net94));
 sg13g2_o21ai_1 _0877_ (.B1(net104),
    .Y(_0398_),
    .A1(net91),
    .A2(net64));
 sg13g2_a21oi_1 _0878_ (.A1(net91),
    .A2(_0380_),
    .Y(_0046_),
    .B1(_0398_));
 sg13g2_a21oi_1 _0879_ (.A1(net99),
    .A2(_0090_),
    .Y(_0399_),
    .B1(_0068_));
 sg13g2_a21oi_1 _0880_ (.A1(net84),
    .A2(net80),
    .Y(_0400_),
    .B1(_0399_));
 sg13g2_nor2_1 _0881_ (.A(net95),
    .B(_0400_),
    .Y(_0047_));
 sg13g2_a22oi_1 _0882_ (.Y(_0401_),
    .B1(_0115_),
    .B2(_0390_),
    .A2(net70),
    .A1(net86));
 sg13g2_nor2_1 _0883_ (.A(net94),
    .B(_0401_),
    .Y(_0048_));
 sg13g2_nand2_1 _0884_ (.Y(_0402_),
    .A(net83),
    .B(net57));
 sg13g2_a21oi_1 _0885_ (.A1(_0095_),
    .A2(_0402_),
    .Y(_0049_),
    .B1(net94));
 sg13g2_nand2_1 _0886_ (.Y(_0403_),
    .A(net84),
    .B(net115));
 sg13g2_a21oi_1 _0887_ (.A1(_0107_),
    .A2(_0403_),
    .Y(_0050_),
    .B1(net94));
 sg13g2_nand2_1 _0888_ (.Y(_0404_),
    .A(net85),
    .B(net109));
 sg13g2_a21oi_1 _0889_ (.A1(_0382_),
    .A2(_0404_),
    .Y(_0051_),
    .B1(net95));
 sg13g2_o21ai_1 _0890_ (.B1(net104),
    .Y(_0405_),
    .A1(net89),
    .A2(net126));
 sg13g2_a21oi_1 _0891_ (.A1(net89),
    .A2(_0088_),
    .Y(_0052_),
    .B1(_0405_));
 sg13g2_a21oi_1 _0892_ (.A1(_0086_),
    .A2(_0383_),
    .Y(_0406_),
    .B1(_0091_));
 sg13g2_o21ai_1 _0893_ (.B1(net104),
    .Y(_0407_),
    .A1(net89),
    .A2(net116));
 sg13g2_nor2_1 _0894_ (.A(_0406_),
    .B(_0407_),
    .Y(_0053_));
 sg13g2_nand2_1 _0895_ (.Y(_0408_),
    .A(net107),
    .B(net83));
 sg13g2_a21oi_1 _0896_ (.A1(_0096_),
    .A2(_0408_),
    .Y(_0054_),
    .B1(net94));
 sg13g2_dfrbp_1 _0897_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net36),
    .D(_0006_),
    .Q_N(_0452_),
    .Q(\hn5.hidden_neuron_o[0] ));
 sg13g2_dfrbp_1 _0898_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net48),
    .D(_0007_),
    .Q_N(_0451_),
    .Q(\hn5.hidden_neuron_o[1] ));
 sg13g2_dfrbp_1 _0899_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net46),
    .D(_0008_),
    .Q_N(_0450_),
    .Q(\hn5.hidden_neuron_o[2] ));
 sg13g2_dfrbp_1 _0900_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net44),
    .D(_0009_),
    .Q_N(_0449_),
    .Q(\hn5.hidden_neuron_o[3] ));
 sg13g2_dfrbp_1 _0901_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net41),
    .D(_0010_),
    .Q_N(_0448_),
    .Q(\hn5.hidden_neuron_o[4] ));
 sg13g2_dfrbp_1 _0902_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net39),
    .D(net125),
    .Q_N(_0447_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _0903_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net37),
    .D(net129),
    .Q_N(_0446_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _0904_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net35),
    .D(_0013_),
    .Q_N(_0445_),
    .Q(\hn6.hidden_neuron_o[0] ));
 sg13g2_dfrbp_1 _0905_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net33),
    .D(_0014_),
    .Q_N(_0444_),
    .Q(\hn6.hidden_neuron_o[1] ));
 sg13g2_dfrbp_1 _0906_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net31),
    .D(_0015_),
    .Q_N(_0443_),
    .Q(\hn6.hidden_neuron_o[2] ));
 sg13g2_dfrbp_1 _0907_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net29),
    .D(_0016_),
    .Q_N(_0442_),
    .Q(\hn6.hidden_neuron_o[3] ));
 sg13g2_dfrbp_1 _0908_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net27),
    .D(_0017_),
    .Q_N(_0441_),
    .Q(\hn6.hidden_neuron_o[4] ));
 sg13g2_dfrbp_1 _0909_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net25),
    .D(_0018_),
    .Q_N(_0440_),
    .Q(\hn7.hidden_neuron_o[0] ));
 sg13g2_dfrbp_1 _0910_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net23),
    .D(_0019_),
    .Q_N(_0439_),
    .Q(\hn7.hidden_neuron_o[1] ));
 sg13g2_dfrbp_1 _0911_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net21),
    .D(_0020_),
    .Q_N(_0438_),
    .Q(\hn7.hidden_neuron_o[2] ));
 sg13g2_dfrbp_1 _0912_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net19),
    .D(_0021_),
    .Q_N(_0437_),
    .Q(\hn7.hidden_neuron_o[3] ));
 sg13g2_dfrbp_1 _0913_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net17),
    .D(_0022_),
    .Q_N(_0436_),
    .Q(\hn7.hidden_neuron_o[4] ));
 sg13g2_dfrbp_1 _0914_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net103),
    .D(_0023_),
    .Q_N(_0435_),
    .Q(\final_o[0] ));
 sg13g2_dfrbp_1 _0915_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net103),
    .D(_0024_),
    .Q_N(_0434_),
    .Q(\final_o[1] ));
 sg13g2_dfrbp_1 _0916_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net103),
    .D(_0025_),
    .Q_N(_0433_),
    .Q(\final_o[2] ));
 sg13g2_dfrbp_1 _0917_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net102),
    .D(_0026_),
    .Q_N(_0432_),
    .Q(\final_o[3] ));
 sg13g2_dfrbp_1 _0918_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net102),
    .D(_0027_),
    .Q_N(_0431_),
    .Q(\final_o[4] ));
 sg13g2_dfrbp_1 _0919_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net102),
    .D(_0028_),
    .Q_N(_0430_),
    .Q(\final_o[5] ));
 sg13g2_dfrbp_1 _0920_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net102),
    .D(_0029_),
    .Q_N(_0429_),
    .Q(\final_o[6] ));
 sg13g2_dfrbp_1 _0921_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net103),
    .D(_0030_),
    .Q_N(_0428_),
    .Q(\final_o[7] ));
 sg13g2_dfrbp_1 _0922_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net102),
    .D(_0031_),
    .Q_N(_0427_),
    .Q(\final_o[8] ));
 sg13g2_dfrbp_1 _0923_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net102),
    .D(_0032_),
    .Q_N(_0426_),
    .Q(\final_o[9] ));
 sg13g2_dfrbp_1 _0924_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net103),
    .D(_0033_),
    .Q_N(_0425_),
    .Q(\final_o[10] ));
 sg13g2_dllrq_1 _0925_ (.D(\sm0.state_d[1] ),
    .GATE_N(_0000_),
    .RESET_B(net42),
    .Q(f0p_o));
 sg13g2_dfrbp_1 _0926_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net54),
    .D(_0034_),
    .Q_N(_0424_),
    .Q(\hn0.hidden_neuron_o[0] ));
 sg13g2_dfrbp_1 _0927_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net52),
    .D(_0035_),
    .Q_N(_0423_),
    .Q(\hn0.hidden_neuron_o[1] ));
 sg13g2_dfrbp_1 _0928_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net50),
    .D(_0036_),
    .Q_N(_0422_),
    .Q(\hn0.hidden_neuron_o[2] ));
 sg13g2_dfrbp_1 _0929_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net47),
    .D(_0037_),
    .Q_N(_0421_),
    .Q(\hn0.hidden_neuron_o[3] ));
 sg13g2_dfrbp_1 _0930_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net43),
    .D(_0038_),
    .Q_N(_0420_),
    .Q(\hn1.hidden_neuron_o[0] ));
 sg13g2_dfrbp_1 _0931_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net38),
    .D(_0039_),
    .Q_N(_0419_),
    .Q(\hn1.hidden_neuron_o[1] ));
 sg13g2_dfrbp_1 _0932_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net34),
    .D(_0040_),
    .Q_N(_0418_),
    .Q(\hn1.hidden_neuron_o[2] ));
 sg13g2_dfrbp_1 _0933_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net30),
    .D(_0041_),
    .Q_N(_0417_),
    .Q(\hn1.hidden_neuron_o[3] ));
 sg13g2_dfrbp_1 _0934_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net26),
    .D(_0042_),
    .Q_N(_0416_),
    .Q(\hn2.hidden_neuron_o[0] ));
 sg13g2_dfrbp_1 _0935_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net22),
    .D(_0043_),
    .Q_N(_0415_),
    .Q(\hn2.hidden_neuron_o[1] ));
 sg13g2_dfrbp_1 _0936_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net18),
    .D(_0044_),
    .Q_N(_0414_),
    .Q(\hn2.hidden_neuron_o[2] ));
 sg13g2_dfrbp_1 _0937_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net53),
    .D(_0045_),
    .Q_N(_0413_),
    .Q(\hn2.hidden_neuron_o[3] ));
 sg13g2_dfrbp_1 _0938_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net49),
    .D(_0046_),
    .Q_N(_0002_),
    .Q(\hn3.hidden_neuron_o[0] ));
 sg13g2_dfrbp_1 _0939_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net40),
    .D(_0047_),
    .Q_N(_0412_),
    .Q(\hn3.hidden_neuron_o[1] ));
 sg13g2_dfrbp_1 _0940_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net32),
    .D(_0048_),
    .Q_N(_0003_),
    .Q(\hn3.hidden_neuron_o[2] ));
 sg13g2_dfrbp_1 _0941_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net24),
    .D(_0049_),
    .Q_N(_0004_),
    .Q(\hn3.hidden_neuron_o[3] ));
 sg13g2_dfrbp_1 _0942_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net16),
    .D(_0050_),
    .Q_N(_0411_),
    .Q(\hn4.hidden_neuron_o[0] ));
 sg13g2_dfrbp_1 _0943_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net45),
    .D(_0051_),
    .Q_N(_0001_),
    .Q(\hn4.hidden_neuron_o[1] ));
 sg13g2_dfrbp_1 _0944_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net28),
    .D(_0052_),
    .Q_N(_0410_),
    .Q(\hn4.hidden_neuron_o[2] ));
 sg13g2_dfrbp_1 _0945_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net51),
    .D(_0053_),
    .Q_N(_0005_),
    .Q(\hn4.hidden_neuron_o[3] ));
 sg13g2_dfrbp_1 _0946_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net20),
    .D(_0054_),
    .Q_N(_0409_),
    .Q(\hn4.hidden_neuron_o[4] ));
 sg13g2_tiehi _0913__17 (.L_HI(net17));
 sg13g2_tiehi _0936__18 (.L_HI(net18));
 sg13g2_tiehi _0912__19 (.L_HI(net19));
 sg13g2_tiehi _0946__20 (.L_HI(net20));
 sg13g2_tiehi _0911__21 (.L_HI(net21));
 sg13g2_tiehi _0935__22 (.L_HI(net22));
 sg13g2_tiehi _0910__23 (.L_HI(net23));
 sg13g2_tiehi _0941__24 (.L_HI(net24));
 sg13g2_tiehi _0909__25 (.L_HI(net25));
 sg13g2_tiehi _0934__26 (.L_HI(net26));
 sg13g2_tiehi _0908__27 (.L_HI(net27));
 sg13g2_tiehi _0944__28 (.L_HI(net28));
 sg13g2_tiehi _0907__29 (.L_HI(net29));
 sg13g2_tiehi _0933__30 (.L_HI(net30));
 sg13g2_tiehi _0906__31 (.L_HI(net31));
 sg13g2_tiehi _0940__32 (.L_HI(net32));
 sg13g2_tiehi _0905__33 (.L_HI(net33));
 sg13g2_tiehi _0932__34 (.L_HI(net34));
 sg13g2_tiehi _0904__35 (.L_HI(net35));
 sg13g2_tiehi _0897__36 (.L_HI(net36));
 sg13g2_tiehi _0903__37 (.L_HI(net37));
 sg13g2_tiehi _0931__38 (.L_HI(net38));
 sg13g2_tiehi _0902__39 (.L_HI(net39));
 sg13g2_tiehi _0939__40 (.L_HI(net40));
 sg13g2_tiehi _0901__41 (.L_HI(net41));
 sg13g2_tiehi _0925__42 (.L_HI(net42));
 sg13g2_tiehi _0930__43 (.L_HI(net43));
 sg13g2_tiehi _0900__44 (.L_HI(net44));
 sg13g2_tiehi _0943__45 (.L_HI(net45));
 sg13g2_tiehi _0899__46 (.L_HI(net46));
 sg13g2_tiehi _0929__47 (.L_HI(net47));
 sg13g2_tiehi _0898__48 (.L_HI(net48));
 sg13g2_tiehi _0938__49 (.L_HI(net49));
 sg13g2_tiehi _0928__50 (.L_HI(net50));
 sg13g2_tiehi _0945__51 (.L_HI(net51));
 sg13g2_tiehi _0927__52 (.L_HI(net52));
 sg13g2_tiehi _0937__53 (.L_HI(net53));
 sg13g2_tiehi _0926__54 (.L_HI(net54));
 sg13g2_tiehi tt_um_idann_55 (.L_HI(net55));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_idann_6 (.L_LO(net6));
 sg13g2_tielo tt_um_idann_7 (.L_LO(net7));
 sg13g2_tielo tt_um_idann_8 (.L_LO(net8));
 sg13g2_tielo tt_um_idann_9 (.L_LO(net9));
 sg13g2_tielo tt_um_idann_10 (.L_LO(net10));
 sg13g2_tielo tt_um_idann_11 (.L_LO(net11));
 sg13g2_tielo tt_um_idann_12 (.L_LO(net12));
 sg13g2_tielo tt_um_idann_13 (.L_LO(net13));
 sg13g2_tielo tt_um_idann_14 (.L_LO(net14));
 sg13g2_tielo tt_um_idann_15 (.L_LO(net15));
 sg13g2_tiehi _0942__16 (.L_HI(net16));
 sg13g2_buf_1 _0998_ (.A(\final_o[8] ),
    .X(uio_out[0]));
 sg13g2_buf_1 _0999_ (.A(\final_o[9] ),
    .X(uio_out[1]));
 sg13g2_buf_1 _1000_ (.A(\final_o[0] ),
    .X(uo_out[0]));
 sg13g2_buf_1 _1001_ (.A(\final_o[1] ),
    .X(uo_out[1]));
 sg13g2_buf_1 _1002_ (.A(\final_o[2] ),
    .X(uo_out[2]));
 sg13g2_buf_1 _1003_ (.A(\final_o[3] ),
    .X(uo_out[3]));
 sg13g2_buf_1 _1004_ (.A(\final_o[4] ),
    .X(uo_out[4]));
 sg13g2_buf_1 _1005_ (.A(\final_o[5] ),
    .X(uo_out[5]));
 sg13g2_buf_1 _1006_ (.A(\final_o[6] ),
    .X(uo_out[6]));
 sg13g2_buf_1 _1007_ (.A(\final_o[7] ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout81 (.A(_0056_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0056_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(net86),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(net85),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(net86),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0056_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(net88),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(net92),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(net90),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(net91),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(net92),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(f0p_o),
    .X(net92));
 sg13g2_buf_4 fanout93 (.X(net93),
    .A(net96));
 sg13g2_buf_4 fanout94 (.X(net94),
    .A(net96));
 sg13g2_buf_2 fanout95 (.A(net96),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_0067_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(net3),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(net2),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(net1),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(net101),
    .X(net100));
 sg13g2_buf_1 fanout101 (.A(ui_in[0]),
    .X(net101));
 sg13g2_buf_4 fanout102 (.X(net102),
    .A(net103));
 sg13g2_buf_4 fanout103 (.X(net103),
    .A(net105));
 sg13g2_buf_2 fanout104 (.A(net105),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(rst_n),
    .X(net105));
 sg13g2_buf_1 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[7]),
    .X(net4));
 sg13g2_tielo tt_um_idann_5 (.L_LO(net5));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_3_4__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\final_o[10] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold2 (.A(\hn3.hidden_neuron_o[3] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold3 (.A(\final_o[4] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold4 (.A(\final_o[0] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold5 (.A(\final_o[3] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold6 (.A(\final_o[1] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold7 (.A(\final_o[6] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold8 (.A(\final_o[7] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold9 (.A(\hn3.hidden_neuron_o[0] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold10 (.A(\hn0.hidden_neuron_o[2] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold11 (.A(\final_o[5] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold12 (.A(\final_o[8] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold13 (.A(\hn0.hidden_neuron_o[1] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold14 (.A(\final_o[2] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold15 (.A(\hn3.hidden_neuron_o[2] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold16 (.A(\hn1.hidden_neuron_o[2] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold17 (.A(\hn0.hidden_neuron_o[3] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold18 (.A(\hn0.hidden_neuron_o[0] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold19 (.A(\hn1.hidden_neuron_o[1] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold20 (.A(\hn7.hidden_neuron_o[4] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold21 (.A(\hn7.hidden_neuron_o[0] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold22 (.A(\hn1.hidden_neuron_o[0] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold23 (.A(\final_o[9] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold24 (.A(\hn5.hidden_neuron_o[4] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold25 (.A(\hn3.hidden_neuron_o[1] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold26 (.A(\hn7.hidden_neuron_o[2] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold27 (.A(\hn4.hidden_neuron_o[4] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold28 (.A(\hn2.hidden_neuron_o[3] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold29 (.A(\hn4.hidden_neuron_o[1] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold30 (.A(\hn5.hidden_neuron_o[3] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold31 (.A(\hn5.hidden_neuron_o[2] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold32 (.A(\hn7.hidden_neuron_o[1] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold33 (.A(\hn2.hidden_neuron_o[1] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold34 (.A(\hn6.hidden_neuron_o[1] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold35 (.A(\hn4.hidden_neuron_o[0] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold36 (.A(\hn4.hidden_neuron_o[3] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold37 (.A(\hn7.hidden_neuron_o[3] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold38 (.A(\hn2.hidden_neuron_o[0] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold39 (.A(\hn6.hidden_neuron_o[4] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold40 (.A(\hn6.hidden_neuron_o[0] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold41 (.A(\hn2.hidden_neuron_o[2] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold42 (.A(\hn1.hidden_neuron_o[3] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold43 (.A(\hn5.hidden_neuron_o[0] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold44 (.A(uio_out[5]),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0011_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold46 (.A(\hn4.hidden_neuron_o[2] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold47 (.A(\hn5.hidden_neuron_o[1] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold48 (.A(uio_out[6]),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0012_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold50 (.A(\hn6.hidden_neuron_o[2] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold51 (.A(\hn6.hidden_neuron_o[3] ),
    .X(net131));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_4 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_254 ();
 sg13g2_decap_8 FILLER_18_261 ();
 sg13g2_decap_8 FILLER_18_268 ();
 sg13g2_decap_8 FILLER_18_275 ();
 sg13g2_decap_8 FILLER_18_282 ();
 sg13g2_decap_8 FILLER_18_289 ();
 sg13g2_decap_8 FILLER_18_296 ();
 sg13g2_decap_8 FILLER_18_303 ();
 sg13g2_decap_8 FILLER_18_310 ();
 sg13g2_decap_8 FILLER_18_317 ();
 sg13g2_decap_8 FILLER_18_324 ();
 sg13g2_decap_8 FILLER_18_331 ();
 sg13g2_decap_8 FILLER_18_338 ();
 sg13g2_decap_8 FILLER_18_345 ();
 sg13g2_decap_8 FILLER_18_352 ();
 sg13g2_decap_8 FILLER_18_359 ();
 sg13g2_decap_8 FILLER_18_366 ();
 sg13g2_decap_8 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_fill_2 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_186 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_decap_8 FILLER_19_200 ();
 sg13g2_decap_8 FILLER_19_207 ();
 sg13g2_decap_8 FILLER_19_214 ();
 sg13g2_decap_4 FILLER_19_221 ();
 sg13g2_fill_2 FILLER_19_225 ();
 sg13g2_decap_8 FILLER_19_232 ();
 sg13g2_decap_4 FILLER_19_239 ();
 sg13g2_fill_1 FILLER_19_243 ();
 sg13g2_fill_2 FILLER_19_265 ();
 sg13g2_decap_4 FILLER_19_271 ();
 sg13g2_fill_1 FILLER_19_275 ();
 sg13g2_decap_8 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_291 ();
 sg13g2_decap_8 FILLER_19_298 ();
 sg13g2_decap_8 FILLER_19_305 ();
 sg13g2_decap_8 FILLER_19_312 ();
 sg13g2_decap_8 FILLER_19_319 ();
 sg13g2_decap_8 FILLER_19_326 ();
 sg13g2_decap_8 FILLER_19_333 ();
 sg13g2_decap_8 FILLER_19_340 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_decap_8 FILLER_19_361 ();
 sg13g2_decap_8 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_fill_2 FILLER_20_168 ();
 sg13g2_fill_1 FILLER_20_170 ();
 sg13g2_fill_2 FILLER_20_195 ();
 sg13g2_fill_1 FILLER_20_210 ();
 sg13g2_decap_4 FILLER_20_215 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_decap_4 FILLER_20_241 ();
 sg13g2_fill_2 FILLER_20_245 ();
 sg13g2_fill_2 FILLER_20_263 ();
 sg13g2_decap_8 FILLER_20_289 ();
 sg13g2_fill_2 FILLER_20_296 ();
 sg13g2_fill_1 FILLER_20_298 ();
 sg13g2_decap_4 FILLER_20_316 ();
 sg13g2_fill_2 FILLER_20_320 ();
 sg13g2_decap_8 FILLER_20_327 ();
 sg13g2_decap_4 FILLER_20_334 ();
 sg13g2_fill_2 FILLER_20_338 ();
 sg13g2_fill_1 FILLER_20_344 ();
 sg13g2_decap_8 FILLER_20_358 ();
 sg13g2_decap_4 FILLER_20_365 ();
 sg13g2_decap_8 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_fill_1 FILLER_21_147 ();
 sg13g2_decap_4 FILLER_21_191 ();
 sg13g2_decap_8 FILLER_21_226 ();
 sg13g2_decap_4 FILLER_21_233 ();
 sg13g2_fill_2 FILLER_21_237 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_4 FILLER_21_266 ();
 sg13g2_fill_1 FILLER_21_270 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_4 FILLER_21_292 ();
 sg13g2_fill_2 FILLER_21_322 ();
 sg13g2_fill_2 FILLER_21_359 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_fill_1 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_146 ();
 sg13g2_decap_4 FILLER_22_153 ();
 sg13g2_fill_2 FILLER_22_157 ();
 sg13g2_decap_4 FILLER_22_177 ();
 sg13g2_fill_2 FILLER_22_211 ();
 sg13g2_fill_1 FILLER_22_213 ();
 sg13g2_fill_2 FILLER_22_240 ();
 sg13g2_fill_2 FILLER_22_265 ();
 sg13g2_fill_1 FILLER_22_267 ();
 sg13g2_fill_1 FILLER_22_284 ();
 sg13g2_fill_2 FILLER_22_305 ();
 sg13g2_fill_2 FILLER_22_311 ();
 sg13g2_decap_8 FILLER_22_317 ();
 sg13g2_fill_2 FILLER_22_324 ();
 sg13g2_fill_1 FILLER_22_326 ();
 sg13g2_fill_2 FILLER_22_332 ();
 sg13g2_fill_1 FILLER_22_334 ();
 sg13g2_decap_8 FILLER_22_339 ();
 sg13g2_decap_4 FILLER_22_346 ();
 sg13g2_fill_1 FILLER_22_360 ();
 sg13g2_decap_4 FILLER_22_366 ();
 sg13g2_fill_2 FILLER_22_370 ();
 sg13g2_decap_4 FILLER_22_376 ();
 sg13g2_fill_1 FILLER_22_380 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_4 FILLER_23_119 ();
 sg13g2_fill_2 FILLER_23_165 ();
 sg13g2_decap_4 FILLER_23_186 ();
 sg13g2_fill_2 FILLER_23_190 ();
 sg13g2_fill_1 FILLER_23_196 ();
 sg13g2_fill_2 FILLER_23_201 ();
 sg13g2_fill_2 FILLER_23_234 ();
 sg13g2_fill_2 FILLER_23_248 ();
 sg13g2_fill_1 FILLER_23_255 ();
 sg13g2_decap_8 FILLER_23_264 ();
 sg13g2_fill_1 FILLER_23_271 ();
 sg13g2_decap_8 FILLER_23_277 ();
 sg13g2_decap_4 FILLER_23_284 ();
 sg13g2_fill_2 FILLER_23_288 ();
 sg13g2_decap_4 FILLER_23_295 ();
 sg13g2_fill_2 FILLER_23_345 ();
 sg13g2_fill_1 FILLER_23_347 ();
 sg13g2_fill_2 FILLER_23_361 ();
 sg13g2_fill_2 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_4 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_183 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_decap_4 FILLER_24_244 ();
 sg13g2_decap_4 FILLER_24_258 ();
 sg13g2_fill_1 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_267 ();
 sg13g2_fill_2 FILLER_24_276 ();
 sg13g2_decap_4 FILLER_24_291 ();
 sg13g2_fill_1 FILLER_24_314 ();
 sg13g2_decap_4 FILLER_24_338 ();
 sg13g2_fill_1 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_decap_4 FILLER_24_373 ();
 sg13g2_fill_1 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_fill_2 FILLER_25_112 ();
 sg13g2_fill_2 FILLER_25_150 ();
 sg13g2_fill_1 FILLER_25_152 ();
 sg13g2_fill_2 FILLER_25_158 ();
 sg13g2_fill_2 FILLER_25_164 ();
 sg13g2_fill_1 FILLER_25_166 ();
 sg13g2_fill_1 FILLER_25_172 ();
 sg13g2_decap_8 FILLER_25_184 ();
 sg13g2_fill_1 FILLER_25_191 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_fill_2 FILLER_25_210 ();
 sg13g2_fill_1 FILLER_25_226 ();
 sg13g2_fill_2 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_237 ();
 sg13g2_decap_8 FILLER_25_246 ();
 sg13g2_fill_2 FILLER_25_253 ();
 sg13g2_decap_4 FILLER_25_276 ();
 sg13g2_fill_1 FILLER_25_280 ();
 sg13g2_fill_1 FILLER_25_284 ();
 sg13g2_decap_8 FILLER_25_293 ();
 sg13g2_decap_4 FILLER_25_300 ();
 sg13g2_decap_8 FILLER_25_335 ();
 sg13g2_fill_1 FILLER_25_342 ();
 sg13g2_fill_2 FILLER_25_347 ();
 sg13g2_fill_1 FILLER_25_349 ();
 sg13g2_decap_8 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_377 ();
 sg13g2_fill_1 FILLER_25_384 ();
 sg13g2_fill_2 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_fill_1 FILLER_26_112 ();
 sg13g2_fill_1 FILLER_26_144 ();
 sg13g2_fill_1 FILLER_26_154 ();
 sg13g2_fill_1 FILLER_26_159 ();
 sg13g2_fill_1 FILLER_26_188 ();
 sg13g2_decap_8 FILLER_26_234 ();
 sg13g2_decap_4 FILLER_26_241 ();
 sg13g2_fill_1 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_fill_1 FILLER_26_279 ();
 sg13g2_decap_8 FILLER_26_306 ();
 sg13g2_fill_1 FILLER_26_313 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_fill_2 FILLER_27_131 ();
 sg13g2_fill_1 FILLER_27_133 ();
 sg13g2_fill_2 FILLER_27_165 ();
 sg13g2_fill_2 FILLER_27_176 ();
 sg13g2_fill_1 FILLER_27_178 ();
 sg13g2_decap_8 FILLER_27_184 ();
 sg13g2_fill_1 FILLER_27_191 ();
 sg13g2_fill_1 FILLER_27_200 ();
 sg13g2_decap_4 FILLER_27_210 ();
 sg13g2_fill_2 FILLER_27_235 ();
 sg13g2_fill_1 FILLER_27_237 ();
 sg13g2_fill_1 FILLER_27_259 ();
 sg13g2_fill_2 FILLER_27_276 ();
 sg13g2_fill_1 FILLER_27_290 ();
 sg13g2_decap_8 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_307 ();
 sg13g2_decap_4 FILLER_27_314 ();
 sg13g2_fill_2 FILLER_27_331 ();
 sg13g2_fill_1 FILLER_27_333 ();
 sg13g2_fill_1 FILLER_27_379 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_4 FILLER_28_105 ();
 sg13g2_fill_2 FILLER_28_208 ();
 sg13g2_fill_2 FILLER_28_215 ();
 sg13g2_fill_1 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_235 ();
 sg13g2_decap_4 FILLER_28_242 ();
 sg13g2_fill_1 FILLER_28_246 ();
 sg13g2_decap_8 FILLER_28_256 ();
 sg13g2_decap_4 FILLER_28_272 ();
 sg13g2_fill_2 FILLER_28_295 ();
 sg13g2_fill_1 FILLER_28_297 ();
 sg13g2_fill_2 FILLER_28_329 ();
 sg13g2_fill_1 FILLER_28_331 ();
 sg13g2_fill_2 FILLER_28_346 ();
 sg13g2_fill_1 FILLER_28_353 ();
 sg13g2_fill_2 FILLER_28_362 ();
 sg13g2_fill_1 FILLER_28_364 ();
 sg13g2_fill_2 FILLER_28_370 ();
 sg13g2_fill_2 FILLER_28_382 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_fill_2 FILLER_29_105 ();
 sg13g2_fill_1 FILLER_29_107 ();
 sg13g2_fill_1 FILLER_29_134 ();
 sg13g2_decap_8 FILLER_29_158 ();
 sg13g2_fill_1 FILLER_29_174 ();
 sg13g2_decap_8 FILLER_29_193 ();
 sg13g2_decap_8 FILLER_29_200 ();
 sg13g2_fill_1 FILLER_29_233 ();
 sg13g2_fill_2 FILLER_29_276 ();
 sg13g2_fill_2 FILLER_29_283 ();
 sg13g2_decap_4 FILLER_29_303 ();
 sg13g2_fill_2 FILLER_29_317 ();
 sg13g2_fill_2 FILLER_29_325 ();
 sg13g2_decap_4 FILLER_29_343 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_fill_2 FILLER_29_352 ();
 sg13g2_fill_1 FILLER_29_354 ();
 sg13g2_fill_1 FILLER_29_359 ();
 sg13g2_fill_2 FILLER_29_368 ();
 sg13g2_fill_1 FILLER_29_370 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_fill_1 FILLER_30_98 ();
 sg13g2_fill_2 FILLER_30_117 ();
 sg13g2_decap_4 FILLER_30_122 ();
 sg13g2_fill_1 FILLER_30_126 ();
 sg13g2_decap_4 FILLER_30_136 ();
 sg13g2_fill_2 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_184 ();
 sg13g2_fill_2 FILLER_30_191 ();
 sg13g2_fill_2 FILLER_30_198 ();
 sg13g2_fill_2 FILLER_30_217 ();
 sg13g2_fill_1 FILLER_30_219 ();
 sg13g2_fill_2 FILLER_30_233 ();
 sg13g2_fill_2 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_255 ();
 sg13g2_fill_2 FILLER_30_262 ();
 sg13g2_fill_1 FILLER_30_264 ();
 sg13g2_decap_8 FILLER_30_269 ();
 sg13g2_decap_8 FILLER_30_276 ();
 sg13g2_fill_2 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_290 ();
 sg13g2_fill_1 FILLER_30_310 ();
 sg13g2_fill_2 FILLER_30_323 ();
 sg13g2_fill_2 FILLER_30_331 ();
 sg13g2_decap_4 FILLER_30_338 ();
 sg13g2_fill_1 FILLER_30_342 ();
 sg13g2_fill_2 FILLER_30_348 ();
 sg13g2_fill_1 FILLER_30_350 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_fill_2 FILLER_31_84 ();
 sg13g2_fill_1 FILLER_31_86 ();
 sg13g2_fill_1 FILLER_31_113 ();
 sg13g2_fill_1 FILLER_31_140 ();
 sg13g2_fill_1 FILLER_31_161 ();
 sg13g2_fill_2 FILLER_31_175 ();
 sg13g2_fill_2 FILLER_31_187 ();
 sg13g2_decap_4 FILLER_31_227 ();
 sg13g2_fill_1 FILLER_31_231 ();
 sg13g2_fill_2 FILLER_31_252 ();
 sg13g2_fill_2 FILLER_31_280 ();
 sg13g2_fill_2 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_306 ();
 sg13g2_fill_2 FILLER_31_313 ();
 sg13g2_decap_4 FILLER_31_334 ();
 sg13g2_decap_4 FILLER_31_373 ();
 sg13g2_fill_2 FILLER_31_377 ();
 sg13g2_fill_2 FILLER_31_392 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_fill_2 FILLER_32_102 ();
 sg13g2_fill_2 FILLER_32_159 ();
 sg13g2_fill_1 FILLER_32_161 ();
 sg13g2_fill_1 FILLER_32_167 ();
 sg13g2_fill_2 FILLER_32_179 ();
 sg13g2_decap_8 FILLER_32_202 ();
 sg13g2_decap_4 FILLER_32_209 ();
 sg13g2_fill_1 FILLER_32_213 ();
 sg13g2_fill_2 FILLER_32_227 ();
 sg13g2_fill_1 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_243 ();
 sg13g2_decap_4 FILLER_32_256 ();
 sg13g2_fill_2 FILLER_32_260 ();
 sg13g2_decap_4 FILLER_32_275 ();
 sg13g2_fill_2 FILLER_32_293 ();
 sg13g2_fill_2 FILLER_32_312 ();
 sg13g2_decap_8 FILLER_32_340 ();
 sg13g2_fill_2 FILLER_32_347 ();
 sg13g2_decap_4 FILLER_32_353 ();
 sg13g2_decap_4 FILLER_32_366 ();
 sg13g2_fill_1 FILLER_32_370 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_91 ();
 sg13g2_fill_2 FILLER_33_105 ();
 sg13g2_fill_1 FILLER_33_116 ();
 sg13g2_fill_2 FILLER_33_133 ();
 sg13g2_fill_2 FILLER_33_140 ();
 sg13g2_fill_1 FILLER_33_157 ();
 sg13g2_fill_1 FILLER_33_167 ();
 sg13g2_fill_1 FILLER_33_179 ();
 sg13g2_fill_1 FILLER_33_188 ();
 sg13g2_fill_2 FILLER_33_220 ();
 sg13g2_fill_1 FILLER_33_222 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_247 ();
 sg13g2_fill_1 FILLER_33_254 ();
 sg13g2_decap_8 FILLER_33_263 ();
 sg13g2_decap_8 FILLER_33_270 ();
 sg13g2_fill_1 FILLER_33_277 ();
 sg13g2_fill_2 FILLER_33_302 ();
 sg13g2_decap_4 FILLER_33_309 ();
 sg13g2_fill_2 FILLER_33_318 ();
 sg13g2_fill_1 FILLER_33_320 ();
 sg13g2_decap_8 FILLER_33_334 ();
 sg13g2_fill_1 FILLER_33_341 ();
 sg13g2_fill_1 FILLER_33_389 ();
 sg13g2_fill_1 FILLER_33_399 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_84 ();
 sg13g2_fill_2 FILLER_34_156 ();
 sg13g2_fill_1 FILLER_34_176 ();
 sg13g2_decap_8 FILLER_34_186 ();
 sg13g2_fill_1 FILLER_34_193 ();
 sg13g2_fill_1 FILLER_34_203 ();
 sg13g2_fill_2 FILLER_34_222 ();
 sg13g2_fill_1 FILLER_34_224 ();
 sg13g2_fill_1 FILLER_34_229 ();
 sg13g2_fill_2 FILLER_34_235 ();
 sg13g2_fill_1 FILLER_34_249 ();
 sg13g2_fill_2 FILLER_34_281 ();
 sg13g2_fill_1 FILLER_34_283 ();
 sg13g2_fill_2 FILLER_34_292 ();
 sg13g2_fill_1 FILLER_34_294 ();
 sg13g2_fill_2 FILLER_34_303 ();
 sg13g2_decap_4 FILLER_34_309 ();
 sg13g2_decap_4 FILLER_34_318 ();
 sg13g2_fill_2 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_333 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_4 FILLER_35_105 ();
 sg13g2_fill_2 FILLER_35_109 ();
 sg13g2_fill_2 FILLER_35_120 ();
 sg13g2_fill_1 FILLER_35_122 ();
 sg13g2_fill_2 FILLER_35_154 ();
 sg13g2_fill_1 FILLER_35_156 ();
 sg13g2_fill_1 FILLER_35_225 ();
 sg13g2_fill_2 FILLER_35_234 ();
 sg13g2_fill_1 FILLER_35_236 ();
 sg13g2_decap_8 FILLER_35_253 ();
 sg13g2_fill_2 FILLER_35_264 ();
 sg13g2_fill_2 FILLER_35_283 ();
 sg13g2_decap_4 FILLER_35_297 ();
 sg13g2_fill_1 FILLER_35_301 ();
 sg13g2_fill_2 FILLER_35_355 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_4 FILLER_36_147 ();
 sg13g2_fill_1 FILLER_36_193 ();
 sg13g2_fill_2 FILLER_36_199 ();
 sg13g2_decap_4 FILLER_36_208 ();
 sg13g2_fill_1 FILLER_36_212 ();
 sg13g2_decap_8 FILLER_36_255 ();
 sg13g2_fill_2 FILLER_36_262 ();
 sg13g2_fill_1 FILLER_36_268 ();
 sg13g2_decap_4 FILLER_36_274 ();
 sg13g2_fill_2 FILLER_36_278 ();
 sg13g2_fill_2 FILLER_36_288 ();
 sg13g2_fill_1 FILLER_36_307 ();
 sg13g2_fill_1 FILLER_36_322 ();
 sg13g2_fill_2 FILLER_36_327 ();
 sg13g2_fill_1 FILLER_36_329 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_fill_1 FILLER_36_348 ();
 sg13g2_fill_1 FILLER_36_372 ();
 sg13g2_fill_1 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_4 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_162 ();
 sg13g2_decap_8 FILLER_37_169 ();
 sg13g2_decap_8 FILLER_37_176 ();
 sg13g2_fill_2 FILLER_37_183 ();
 sg13g2_fill_1 FILLER_37_185 ();
 sg13g2_fill_1 FILLER_37_224 ();
 sg13g2_fill_2 FILLER_37_229 ();
 sg13g2_fill_1 FILLER_37_245 ();
 sg13g2_decap_4 FILLER_37_249 ();
 sg13g2_fill_1 FILLER_37_258 ();
 sg13g2_fill_2 FILLER_37_271 ();
 sg13g2_fill_1 FILLER_37_286 ();
 sg13g2_fill_1 FILLER_37_399 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_8 FILLER_38_124 ();
 sg13g2_decap_8 FILLER_38_131 ();
 sg13g2_decap_4 FILLER_38_138 ();
 sg13g2_fill_2 FILLER_38_142 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_8 FILLER_38_164 ();
 sg13g2_decap_8 FILLER_38_171 ();
 sg13g2_decap_8 FILLER_38_178 ();
 sg13g2_decap_8 FILLER_38_185 ();
 sg13g2_fill_2 FILLER_38_192 ();
 sg13g2_fill_2 FILLER_38_198 ();
 sg13g2_fill_1 FILLER_38_213 ();
 sg13g2_decap_8 FILLER_38_240 ();
 sg13g2_decap_4 FILLER_38_286 ();
 sg13g2_decap_4 FILLER_38_320 ();
 sg13g2_decap_8 FILLER_38_328 ();
 sg13g2_fill_2 FILLER_38_335 ();
 sg13g2_fill_1 FILLER_38_358 ();
 sg13g2_fill_2 FILLER_38_368 ();
 sg13g2_fill_2 FILLER_38_374 ();
 sg13g2_fill_2 FILLER_38_397 ();
 sg13g2_fill_1 FILLER_38_399 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net55;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[7] = net15;
endmodule

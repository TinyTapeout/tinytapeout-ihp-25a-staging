module tt_um_tommythorn_cgates (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire Qc;
 wire Ql;
 wire R16c;
 wire R16ct;
 wire R16l;
 wire R16lt;
 wire R4c;
 wire R4ct;
 wire R4l;
 wire R4lt;
 wire RBigc;
 wire RBigct;
 wire RBigl;
 wire RBiglt;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire \r16ci.genblk1[0].genblk1.combcgate_inst.A ;
 wire \r16ci.genblk1[10].genblk1.combcgate_inst.A ;
 wire \r16ci.genblk1[10].genblk1.combcgate_inst.Q ;
 wire \r16ci.genblk1[11].genblk1.combcgate_inst.Q ;
 wire \r16ci.genblk1[12].genblk1.combcgate_inst.Q ;
 wire \r16ci.genblk1[13].genblk1.combcgate_inst.Q ;
 wire \r16ci.genblk1[14].genblk1.combcgate_inst.Q ;
 wire \r16ci.genblk1[1].genblk1.combcgate_inst.Q ;
 wire \r16ci.genblk1[2].genblk1.combcgate_inst.Q ;
 wire \r16ci.genblk1[3].genblk1.combcgate_inst.Q ;
 wire \r16ci.genblk1[4].genblk1.combcgate_inst.Q ;
 wire \r16ci.genblk1[5].genblk1.combcgate_inst.Q ;
 wire \r16ci.genblk1[6].genblk1.combcgate_inst.Q ;
 wire \r16ci.genblk1[7].genblk1.combcgate_inst.Q ;
 wire \r16ci.genblk1[8].genblk1.combcgate_inst.Q ;
 wire \r16li.genblk1[0].latchcgate_inst.A ;
 wire \r16li.genblk1[10].latchcgate_inst.A ;
 wire \r16li.genblk1[10].latchcgate_inst.Q ;
 wire \r16li.genblk1[11].latchcgate_inst.Q ;
 wire \r16li.genblk1[12].latchcgate_inst.Q ;
 wire \r16li.genblk1[13].latchcgate_inst.Q ;
 wire \r16li.genblk1[14].latchcgate_inst.Q ;
 wire \r16li.genblk1[1].latchcgate_inst.Q ;
 wire \r16li.genblk1[2].latchcgate_inst.Q ;
 wire \r16li.genblk1[3].latchcgate_inst.Q ;
 wire \r16li.genblk1[4].latchcgate_inst.Q ;
 wire \r16li.genblk1[5].latchcgate_inst.Q ;
 wire \r16li.genblk1[6].latchcgate_inst.Q ;
 wire \r16li.genblk1[7].latchcgate_inst.Q ;
 wire \r16li.genblk1[8].latchcgate_inst.Q ;
 wire \r4ci.genblk1[0].genblk1.combcgate_inst.A ;
 wire \r4ci.genblk1[1].genblk1.combcgate_inst.Q ;
 wire \r4ci.genblk1[2].genblk1.combcgate_inst.Q ;
 wire \r4li.genblk1[0].latchcgate_inst.A ;
 wire \r4li.genblk1[1].latchcgate_inst.Q ;
 wire \r4li.genblk1[2].latchcgate_inst.Q ;
 wire \rtbdci.genblk1[0].genblk1.combcgate_inst.A ;
 wire \rtbdci.genblk1[10].genblk1.combcgate_inst.A ;
 wire \rtbdci.genblk1[10].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[11].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[12].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[13].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[14].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[15].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[16].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[17].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[18].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[19].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[1].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[20].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[21].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[22].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[23].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[24].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[25].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[26].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[27].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[28].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[29].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[2].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[30].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[31].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[32].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[33].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[34].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[35].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[36].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[37].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[38].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[39].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[3].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[40].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[41].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[42].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[43].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[44].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[45].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[46].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[47].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[48].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[49].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[4].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[50].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[51].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[52].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[53].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[54].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[55].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[56].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[57].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[58].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[59].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[5].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[60].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[61].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[62].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[6].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[7].genblk1.combcgate_inst.Q ;
 wire \rtbdci.genblk1[8].genblk1.combcgate_inst.Q ;
 wire \rtbdli.genblk1[0].latchcgate_inst.A ;
 wire \rtbdli.genblk1[10].latchcgate_inst.A ;
 wire \rtbdli.genblk1[10].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[11].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[12].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[13].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[14].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[15].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[16].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[17].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[18].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[19].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[1].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[20].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[21].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[22].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[23].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[24].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[25].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[26].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[27].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[28].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[29].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[2].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[30].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[31].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[32].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[33].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[34].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[35].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[36].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[37].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[38].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[39].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[3].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[40].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[41].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[42].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[43].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[44].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[45].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[46].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[47].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[48].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[49].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[4].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[50].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[51].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[52].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[53].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[54].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[55].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[56].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[57].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[58].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[59].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[5].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[60].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[61].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[62].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[6].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[7].latchcgate_inst.Q ;
 wire \rtbdli.genblk1[8].latchcgate_inst.Q ;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net1;
 wire net2;
 wire net3;

 sg13g2_inv_1 _0518_ (.Y(_0174_),
    .A(net172));
 sg13g2_inv_1 _0519_ (.Y(_0175_),
    .A(\rtbdli.genblk1[0].latchcgate_inst.A ));
 sg13g2_inv_1 _0520_ (.Y(_0176_),
    .A(\r4li.genblk1[0].latchcgate_inst.A ));
 sg13g2_inv_1 _0521_ (.Y(_0177_),
    .A(\r16li.genblk1[0].latchcgate_inst.A ));
 sg13g2_inv_1 _0522_ (.Y(_0178_),
    .A(\r16ci.genblk1[1].genblk1.combcgate_inst.Q ));
 sg13g2_inv_1 _0523_ (.Y(_0179_),
    .A(\rtbdci.genblk1[1].genblk1.combcgate_inst.Q ));
 sg13g2_inv_1 _0524_ (.Y(_0180_),
    .A(\r4ci.genblk1[0].genblk1.combcgate_inst.A ));
 sg13g2_inv_1 _0525_ (.Y(_0181_),
    .A(\r4ci.genblk1[2].genblk1.combcgate_inst.Q ));
 sg13g2_inv_1 _0526_ (.Y(_0182_),
    .A(Qc));
 sg13g2_nand2_1 _0527_ (.Y(_0183_),
    .A(\r16ci.genblk1[5].genblk1.combcgate_inst.Q ),
    .B(\r16ci.genblk1[6].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0528_ (.B1(net164),
    .Y(_0184_),
    .A1(\r16ci.genblk1[5].genblk1.combcgate_inst.Q ),
    .A2(\r16ci.genblk1[6].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0529_ (.B1(_0184_),
    .Y(\r16ci.genblk1[6].genblk1.combcgate_inst.Q ),
    .A2(_0183_),
    .A1(\r16ci.genblk1[7].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0530_ (.Y(_0185_),
    .A(\r16ci.genblk1[3].genblk1.combcgate_inst.Q ),
    .B(\r16ci.genblk1[4].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0531_ (.B1(net163),
    .Y(_0186_),
    .A1(\r16ci.genblk1[3].genblk1.combcgate_inst.Q ),
    .A2(\r16ci.genblk1[4].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0532_ (.B1(_0186_),
    .Y(\r16ci.genblk1[4].genblk1.combcgate_inst.Q ),
    .A2(_0185_),
    .A1(\r16ci.genblk1[5].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0533_ (.Y(_0187_),
    .A(\r16ci.genblk1[4].genblk1.combcgate_inst.Q ),
    .B(\r16ci.genblk1[5].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0534_ (.B1(net163),
    .Y(_0188_),
    .A1(\r16ci.genblk1[4].genblk1.combcgate_inst.Q ),
    .A2(\r16ci.genblk1[5].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0535_ (.B1(_0188_),
    .Y(\r16ci.genblk1[5].genblk1.combcgate_inst.Q ),
    .A2(_0187_),
    .A1(\r16ci.genblk1[6].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0536_ (.Y(_0189_),
    .A(\r16ci.genblk1[2].genblk1.combcgate_inst.Q ),
    .B(\r16ci.genblk1[3].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0537_ (.B1(net163),
    .Y(_0190_),
    .A1(\r16ci.genblk1[2].genblk1.combcgate_inst.Q ),
    .A2(\r16ci.genblk1[3].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0538_ (.B1(_0190_),
    .Y(\r16ci.genblk1[3].genblk1.combcgate_inst.Q ),
    .A2(_0189_),
    .A1(\r16ci.genblk1[4].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0539_ (.Y(_0191_),
    .A(\r16ci.genblk1[1].genblk1.combcgate_inst.Q ),
    .B(\r16ci.genblk1[2].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0540_ (.B1(net163),
    .Y(_0192_),
    .A1(\r16ci.genblk1[1].genblk1.combcgate_inst.Q ),
    .A2(\r16ci.genblk1[2].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0541_ (.B1(_0192_),
    .Y(\r16ci.genblk1[2].genblk1.combcgate_inst.Q ),
    .A2(_0191_),
    .A1(\r16ci.genblk1[3].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0542_ (.Y(_0193_),
    .A(R16c),
    .B(\r16ci.genblk1[1].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0543_ (.B1(net165),
    .Y(_0194_),
    .A1(R16c),
    .A2(\r16ci.genblk1[1].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0544_ (.B1(_0194_),
    .Y(\r16ci.genblk1[1].genblk1.combcgate_inst.Q ),
    .A2(_0193_),
    .A1(\r16ci.genblk1[2].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0545_ (.B1(R16c),
    .Y(_0195_),
    .A1(\r16ci.genblk1[0].genblk1.combcgate_inst.A ),
    .A2(_0178_));
 sg13g2_nand2_1 _0546_ (.Y(_0196_),
    .A(\r16ci.genblk1[0].genblk1.combcgate_inst.A ),
    .B(_0178_));
 sg13g2_nand3_1 _0547_ (.B(_0195_),
    .C(_0196_),
    .A(net165),
    .Y(R16c));
 sg13g2_nand2_1 _0548_ (.Y(_0197_),
    .A(\rtbdci.genblk1[0].genblk1.combcgate_inst.A ),
    .B(\rtbdci.genblk1[62].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0549_ (.B1(net162),
    .Y(_0198_),
    .A1(\rtbdci.genblk1[0].genblk1.combcgate_inst.A ),
    .A2(\rtbdci.genblk1[62].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0550_ (.B1(_0198_),
    .Y(\rtbdci.genblk1[0].genblk1.combcgate_inst.A ),
    .A2(_0197_),
    .A1(RBigc));
 sg13g2_nand2_1 _0551_ (.Y(_0199_),
    .A(RBigc),
    .B(\rtbdci.genblk1[1].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0552_ (.B1(net163),
    .Y(_0200_),
    .A1(RBigc),
    .A2(\rtbdci.genblk1[1].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0553_ (.B1(_0200_),
    .Y(\rtbdci.genblk1[1].genblk1.combcgate_inst.Q ),
    .A2(_0199_),
    .A1(\rtbdci.genblk1[2].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0554_ (.B1(RBigc),
    .Y(_0201_),
    .A1(\rtbdci.genblk1[0].genblk1.combcgate_inst.A ),
    .A2(_0179_));
 sg13g2_nand2_1 _0555_ (.Y(_0202_),
    .A(\rtbdci.genblk1[0].genblk1.combcgate_inst.A ),
    .B(_0179_));
 sg13g2_nand3_1 _0556_ (.B(_0201_),
    .C(_0202_),
    .A(net162),
    .Y(RBigc));
 sg13g2_nand2_1 _0557_ (.Y(_0203_),
    .A(\rtbdci.genblk1[61].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[62].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0558_ (.B1(net162),
    .Y(_0204_),
    .A1(\rtbdci.genblk1[61].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[62].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0559_ (.B1(_0204_),
    .Y(\rtbdci.genblk1[62].genblk1.combcgate_inst.Q ),
    .A2(_0203_),
    .A1(\rtbdci.genblk1[0].genblk1.combcgate_inst.A ));
 sg13g2_nand2_1 _0560_ (.Y(_0205_),
    .A(\rtbdci.genblk1[60].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[61].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0561_ (.B1(net162),
    .Y(_0206_),
    .A1(\rtbdci.genblk1[60].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[61].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0562_ (.B1(_0206_),
    .Y(\rtbdci.genblk1[61].genblk1.combcgate_inst.Q ),
    .A2(_0205_),
    .A1(\rtbdci.genblk1[62].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0563_ (.Y(_0207_),
    .A(\rtbdci.genblk1[59].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[60].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0564_ (.B1(net159),
    .Y(_0208_),
    .A1(\rtbdci.genblk1[59].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[60].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0565_ (.B1(_0208_),
    .Y(\rtbdci.genblk1[60].genblk1.combcgate_inst.Q ),
    .A2(_0207_),
    .A1(\rtbdci.genblk1[61].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0566_ (.Y(_0209_),
    .A(\rtbdci.genblk1[58].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[59].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0567_ (.B1(net160),
    .Y(_0210_),
    .A1(\rtbdci.genblk1[58].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[59].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0568_ (.B1(_0210_),
    .Y(\rtbdci.genblk1[59].genblk1.combcgate_inst.Q ),
    .A2(_0209_),
    .A1(\rtbdci.genblk1[60].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0569_ (.Y(_0211_),
    .A(\rtbdci.genblk1[57].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[58].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0570_ (.B1(net159),
    .Y(_0212_),
    .A1(\rtbdci.genblk1[57].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[58].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0571_ (.B1(_0212_),
    .Y(\rtbdci.genblk1[58].genblk1.combcgate_inst.Q ),
    .A2(_0211_),
    .A1(\rtbdci.genblk1[59].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0572_ (.Y(_0213_),
    .A(\rtbdci.genblk1[56].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[57].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0573_ (.B1(net161),
    .Y(_0214_),
    .A1(\rtbdci.genblk1[56].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[57].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0574_ (.B1(_0214_),
    .Y(\rtbdci.genblk1[57].genblk1.combcgate_inst.Q ),
    .A2(_0213_),
    .A1(\rtbdci.genblk1[58].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0575_ (.Y(_0215_),
    .A(\rtbdci.genblk1[55].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[56].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0576_ (.B1(net161),
    .Y(_0216_),
    .A1(\rtbdci.genblk1[55].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[56].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0577_ (.B1(_0216_),
    .Y(\rtbdci.genblk1[56].genblk1.combcgate_inst.Q ),
    .A2(_0215_),
    .A1(\rtbdci.genblk1[57].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0578_ (.Y(_0217_),
    .A(\rtbdci.genblk1[54].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[55].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0579_ (.B1(net161),
    .Y(_0218_),
    .A1(\rtbdci.genblk1[54].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[55].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0580_ (.B1(_0218_),
    .Y(\rtbdci.genblk1[55].genblk1.combcgate_inst.Q ),
    .A2(_0217_),
    .A1(\rtbdci.genblk1[56].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0581_ (.Y(_0219_),
    .A(\rtbdci.genblk1[53].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[54].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0582_ (.B1(net160),
    .Y(_0220_),
    .A1(\rtbdci.genblk1[53].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[54].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0583_ (.B1(_0220_),
    .Y(\rtbdci.genblk1[54].genblk1.combcgate_inst.Q ),
    .A2(_0219_),
    .A1(\rtbdci.genblk1[55].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0584_ (.Y(_0221_),
    .A(\rtbdci.genblk1[52].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[53].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0585_ (.B1(net161),
    .Y(_0222_),
    .A1(\rtbdci.genblk1[52].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[53].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0586_ (.B1(_0222_),
    .Y(\rtbdci.genblk1[53].genblk1.combcgate_inst.Q ),
    .A2(_0221_),
    .A1(\rtbdci.genblk1[54].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0587_ (.Y(_0223_),
    .A(\rtbdci.genblk1[51].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[52].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0588_ (.B1(net155),
    .Y(_0224_),
    .A1(\rtbdci.genblk1[51].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[52].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0589_ (.B1(_0224_),
    .Y(\rtbdci.genblk1[52].genblk1.combcgate_inst.Q ),
    .A2(_0223_),
    .A1(\rtbdci.genblk1[53].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0590_ (.Y(_0225_),
    .A(\rtbdci.genblk1[50].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[51].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0591_ (.B1(net154),
    .Y(_0226_),
    .A1(\rtbdci.genblk1[50].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[51].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0592_ (.B1(_0226_),
    .Y(\rtbdci.genblk1[51].genblk1.combcgate_inst.Q ),
    .A2(_0225_),
    .A1(\rtbdci.genblk1[52].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0593_ (.Y(_0227_),
    .A(\rtbdci.genblk1[49].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[50].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0594_ (.B1(net154),
    .Y(_0228_),
    .A1(\rtbdci.genblk1[49].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[50].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0595_ (.B1(_0228_),
    .Y(\rtbdci.genblk1[50].genblk1.combcgate_inst.Q ),
    .A2(_0227_),
    .A1(\rtbdci.genblk1[51].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0596_ (.Y(_0229_),
    .A(\rtbdci.genblk1[48].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[49].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0597_ (.B1(net154),
    .Y(_0230_),
    .A1(\rtbdci.genblk1[48].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[49].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0598_ (.B1(_0230_),
    .Y(\rtbdci.genblk1[49].genblk1.combcgate_inst.Q ),
    .A2(_0229_),
    .A1(\rtbdci.genblk1[50].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0599_ (.Y(_0231_),
    .A(\rtbdci.genblk1[47].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[48].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0600_ (.B1(net154),
    .Y(_0232_),
    .A1(\rtbdci.genblk1[47].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[48].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0601_ (.B1(_0232_),
    .Y(\rtbdci.genblk1[48].genblk1.combcgate_inst.Q ),
    .A2(_0231_),
    .A1(\rtbdci.genblk1[49].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0602_ (.Y(_0233_),
    .A(\rtbdci.genblk1[46].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[47].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0603_ (.B1(net154),
    .Y(_0234_),
    .A1(\rtbdci.genblk1[46].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[47].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0604_ (.B1(_0234_),
    .Y(\rtbdci.genblk1[47].genblk1.combcgate_inst.Q ),
    .A2(_0233_),
    .A1(\rtbdci.genblk1[48].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0605_ (.Y(_0235_),
    .A(\rtbdci.genblk1[45].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[46].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0606_ (.B1(net154),
    .Y(_0236_),
    .A1(\rtbdci.genblk1[45].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[46].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0607_ (.B1(_0236_),
    .Y(\rtbdci.genblk1[46].genblk1.combcgate_inst.Q ),
    .A2(_0235_),
    .A1(\rtbdci.genblk1[47].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0608_ (.Y(_0237_),
    .A(\rtbdci.genblk1[44].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[45].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0609_ (.B1(net154),
    .Y(_0238_),
    .A1(\rtbdci.genblk1[44].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[45].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0610_ (.B1(_0238_),
    .Y(\rtbdci.genblk1[45].genblk1.combcgate_inst.Q ),
    .A2(_0237_),
    .A1(\rtbdci.genblk1[46].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0611_ (.Y(_0239_),
    .A(\rtbdci.genblk1[43].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[44].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0612_ (.B1(net154),
    .Y(_0240_),
    .A1(\rtbdci.genblk1[43].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[44].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0613_ (.B1(_0240_),
    .Y(\rtbdci.genblk1[44].genblk1.combcgate_inst.Q ),
    .A2(_0239_),
    .A1(\rtbdci.genblk1[45].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0614_ (.Y(_0241_),
    .A(\rtbdci.genblk1[42].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[43].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0615_ (.B1(net151),
    .Y(_0242_),
    .A1(\rtbdci.genblk1[42].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[43].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0616_ (.B1(_0242_),
    .Y(\rtbdci.genblk1[43].genblk1.combcgate_inst.Q ),
    .A2(_0241_),
    .A1(\rtbdci.genblk1[44].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0617_ (.Y(_0243_),
    .A(\rtbdci.genblk1[41].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[42].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0618_ (.B1(net151),
    .Y(_0244_),
    .A1(\rtbdci.genblk1[41].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[42].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0619_ (.B1(_0244_),
    .Y(\rtbdci.genblk1[42].genblk1.combcgate_inst.Q ),
    .A2(_0243_),
    .A1(\rtbdci.genblk1[43].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0620_ (.Y(_0245_),
    .A(\rtbdci.genblk1[40].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[41].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0621_ (.B1(net151),
    .Y(_0246_),
    .A1(\rtbdci.genblk1[40].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[41].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0622_ (.B1(_0246_),
    .Y(\rtbdci.genblk1[41].genblk1.combcgate_inst.Q ),
    .A2(_0245_),
    .A1(\rtbdci.genblk1[42].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0623_ (.Y(_0247_),
    .A(\rtbdci.genblk1[39].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[40].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0624_ (.B1(net151),
    .Y(_0248_),
    .A1(\rtbdci.genblk1[39].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[40].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0625_ (.B1(_0248_),
    .Y(\rtbdci.genblk1[40].genblk1.combcgate_inst.Q ),
    .A2(_0247_),
    .A1(\rtbdci.genblk1[41].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0626_ (.Y(_0249_),
    .A(\rtbdci.genblk1[38].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[39].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0627_ (.B1(net152),
    .Y(_0250_),
    .A1(\rtbdci.genblk1[38].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[39].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0628_ (.B1(_0250_),
    .Y(\rtbdci.genblk1[39].genblk1.combcgate_inst.Q ),
    .A2(_0249_),
    .A1(\rtbdci.genblk1[40].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0629_ (.Y(_0251_),
    .A(\rtbdci.genblk1[37].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[38].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0630_ (.B1(net151),
    .Y(_0252_),
    .A1(\rtbdci.genblk1[37].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[38].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0631_ (.B1(_0252_),
    .Y(\rtbdci.genblk1[38].genblk1.combcgate_inst.Q ),
    .A2(_0251_),
    .A1(\rtbdci.genblk1[39].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0632_ (.Y(_0253_),
    .A(\rtbdci.genblk1[36].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[37].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0633_ (.B1(net151),
    .Y(_0254_),
    .A1(\rtbdci.genblk1[36].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[37].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0634_ (.B1(_0254_),
    .Y(\rtbdci.genblk1[37].genblk1.combcgate_inst.Q ),
    .A2(_0253_),
    .A1(\rtbdci.genblk1[38].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0635_ (.Y(_0255_),
    .A(\rtbdci.genblk1[35].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[36].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0636_ (.B1(net151),
    .Y(_0256_),
    .A1(\rtbdci.genblk1[35].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[36].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0637_ (.B1(_0256_),
    .Y(\rtbdci.genblk1[36].genblk1.combcgate_inst.Q ),
    .A2(_0255_),
    .A1(\rtbdci.genblk1[37].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0638_ (.Y(_0257_),
    .A(\rtbdci.genblk1[34].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[35].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0639_ (.B1(net151),
    .Y(_0258_),
    .A1(\rtbdci.genblk1[34].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[35].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0640_ (.B1(_0258_),
    .Y(\rtbdci.genblk1[35].genblk1.combcgate_inst.Q ),
    .A2(_0257_),
    .A1(\rtbdci.genblk1[36].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0641_ (.Y(_0259_),
    .A(\rtbdci.genblk1[33].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[34].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0642_ (.B1(net150),
    .Y(_0260_),
    .A1(\rtbdci.genblk1[33].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[34].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0643_ (.B1(_0260_),
    .Y(\rtbdci.genblk1[34].genblk1.combcgate_inst.Q ),
    .A2(_0259_),
    .A1(\rtbdci.genblk1[35].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0644_ (.Y(_0261_),
    .A(\rtbdci.genblk1[32].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[33].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0645_ (.B1(net150),
    .Y(_0262_),
    .A1(\rtbdci.genblk1[32].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[33].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0646_ (.B1(_0262_),
    .Y(\rtbdci.genblk1[33].genblk1.combcgate_inst.Q ),
    .A2(_0261_),
    .A1(\rtbdci.genblk1[34].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0647_ (.Y(_0263_),
    .A(\rtbdci.genblk1[31].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[32].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0648_ (.B1(net150),
    .Y(_0264_),
    .A1(\rtbdci.genblk1[31].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[32].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0649_ (.B1(_0264_),
    .Y(\rtbdci.genblk1[32].genblk1.combcgate_inst.Q ),
    .A2(_0263_),
    .A1(\rtbdci.genblk1[33].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0650_ (.Y(_0265_),
    .A(\rtbdci.genblk1[30].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[31].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0651_ (.B1(net150),
    .Y(_0266_),
    .A1(\rtbdci.genblk1[30].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[31].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0652_ (.B1(_0266_),
    .Y(\rtbdci.genblk1[31].genblk1.combcgate_inst.Q ),
    .A2(_0265_),
    .A1(\rtbdci.genblk1[32].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0653_ (.Y(_0267_),
    .A(\rtbdci.genblk1[29].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[30].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0654_ (.B1(net150),
    .Y(_0268_),
    .A1(\rtbdci.genblk1[29].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[30].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0655_ (.B1(_0268_),
    .Y(\rtbdci.genblk1[30].genblk1.combcgate_inst.Q ),
    .A2(_0267_),
    .A1(\rtbdci.genblk1[31].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0656_ (.Y(_0269_),
    .A(\rtbdci.genblk1[28].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[29].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0657_ (.B1(net150),
    .Y(_0270_),
    .A1(\rtbdci.genblk1[28].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[29].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0658_ (.B1(_0270_),
    .Y(\rtbdci.genblk1[29].genblk1.combcgate_inst.Q ),
    .A2(_0269_),
    .A1(\rtbdci.genblk1[30].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0659_ (.Y(_0271_),
    .A(\rtbdci.genblk1[27].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[28].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0660_ (.B1(net152),
    .Y(_0272_),
    .A1(\rtbdci.genblk1[27].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[28].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0661_ (.B1(_0272_),
    .Y(\rtbdci.genblk1[28].genblk1.combcgate_inst.Q ),
    .A2(_0271_),
    .A1(\rtbdci.genblk1[29].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0662_ (.Y(_0273_),
    .A(\rtbdci.genblk1[26].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[27].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0663_ (.B1(net152),
    .Y(_0274_),
    .A1(\rtbdci.genblk1[26].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[27].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0664_ (.B1(_0274_),
    .Y(\rtbdci.genblk1[27].genblk1.combcgate_inst.Q ),
    .A2(_0273_),
    .A1(\rtbdci.genblk1[28].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0665_ (.Y(_0275_),
    .A(\rtbdci.genblk1[25].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[26].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0666_ (.B1(net150),
    .Y(_0276_),
    .A1(\rtbdci.genblk1[25].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[26].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0667_ (.B1(_0276_),
    .Y(\rtbdci.genblk1[26].genblk1.combcgate_inst.Q ),
    .A2(_0275_),
    .A1(\rtbdci.genblk1[27].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0668_ (.Y(_0277_),
    .A(\rtbdci.genblk1[24].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[25].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0669_ (.B1(net152),
    .Y(_0278_),
    .A1(\rtbdci.genblk1[24].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[25].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0670_ (.B1(_0278_),
    .Y(\rtbdci.genblk1[25].genblk1.combcgate_inst.Q ),
    .A2(_0277_),
    .A1(\rtbdci.genblk1[26].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0671_ (.Y(_0279_),
    .A(\rtbdci.genblk1[23].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[24].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0672_ (.B1(net150),
    .Y(_0280_),
    .A1(\rtbdci.genblk1[23].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[24].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0673_ (.B1(_0280_),
    .Y(\rtbdci.genblk1[24].genblk1.combcgate_inst.Q ),
    .A2(_0279_),
    .A1(\rtbdci.genblk1[25].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0674_ (.Y(_0281_),
    .A(\rtbdci.genblk1[22].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[23].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0675_ (.B1(net153),
    .Y(_0282_),
    .A1(\rtbdci.genblk1[22].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[23].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0676_ (.B1(_0282_),
    .Y(\rtbdci.genblk1[23].genblk1.combcgate_inst.Q ),
    .A2(_0281_),
    .A1(\rtbdci.genblk1[24].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0677_ (.Y(_0283_),
    .A(\rtbdci.genblk1[21].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[22].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0678_ (.B1(net153),
    .Y(_0284_),
    .A1(\rtbdci.genblk1[21].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[22].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0679_ (.B1(_0284_),
    .Y(\rtbdci.genblk1[22].genblk1.combcgate_inst.Q ),
    .A2(_0283_),
    .A1(\rtbdci.genblk1[23].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0680_ (.Y(_0285_),
    .A(\rtbdci.genblk1[20].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[21].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0681_ (.B1(net153),
    .Y(_0286_),
    .A1(\rtbdci.genblk1[20].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[21].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0682_ (.B1(_0286_),
    .Y(\rtbdci.genblk1[21].genblk1.combcgate_inst.Q ),
    .A2(_0285_),
    .A1(\rtbdci.genblk1[22].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0683_ (.Y(_0287_),
    .A(\rtbdci.genblk1[19].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[20].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0684_ (.B1(net153),
    .Y(_0288_),
    .A1(\rtbdci.genblk1[19].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[20].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0685_ (.B1(_0288_),
    .Y(\rtbdci.genblk1[20].genblk1.combcgate_inst.Q ),
    .A2(_0287_),
    .A1(\rtbdci.genblk1[21].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0686_ (.Y(_0289_),
    .A(\rtbdci.genblk1[18].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[19].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0687_ (.B1(net155),
    .Y(_0290_),
    .A1(\rtbdci.genblk1[18].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[19].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0688_ (.B1(_0290_),
    .Y(\rtbdci.genblk1[19].genblk1.combcgate_inst.Q ),
    .A2(_0289_),
    .A1(\rtbdci.genblk1[20].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0689_ (.Y(_0291_),
    .A(\rtbdci.genblk1[17].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[18].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0690_ (.B1(net153),
    .Y(_0292_),
    .A1(\rtbdci.genblk1[17].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[18].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0691_ (.B1(_0292_),
    .Y(\rtbdci.genblk1[18].genblk1.combcgate_inst.Q ),
    .A2(_0291_),
    .A1(\rtbdci.genblk1[19].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0692_ (.Y(_0293_),
    .A(\rtbdci.genblk1[16].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[17].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0693_ (.B1(net153),
    .Y(_0294_),
    .A1(\rtbdci.genblk1[16].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[17].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0694_ (.B1(_0294_),
    .Y(\rtbdci.genblk1[17].genblk1.combcgate_inst.Q ),
    .A2(_0293_),
    .A1(\rtbdci.genblk1[18].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0695_ (.Y(_0295_),
    .A(\rtbdci.genblk1[15].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[16].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0696_ (.B1(net153),
    .Y(_0296_),
    .A1(\rtbdci.genblk1[15].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[16].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0697_ (.B1(_0296_),
    .Y(\rtbdci.genblk1[16].genblk1.combcgate_inst.Q ),
    .A2(_0295_),
    .A1(\rtbdci.genblk1[17].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0698_ (.Y(_0297_),
    .A(\rtbdci.genblk1[14].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[15].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0699_ (.B1(net153),
    .Y(_0298_),
    .A1(\rtbdci.genblk1[14].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[15].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0700_ (.B1(_0298_),
    .Y(\rtbdci.genblk1[15].genblk1.combcgate_inst.Q ),
    .A2(_0297_),
    .A1(\rtbdci.genblk1[16].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0701_ (.Y(_0299_),
    .A(\rtbdci.genblk1[13].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[14].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0702_ (.B1(net159),
    .Y(_0300_),
    .A1(\rtbdci.genblk1[13].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[14].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0703_ (.B1(_0300_),
    .Y(\rtbdci.genblk1[14].genblk1.combcgate_inst.Q ),
    .A2(_0299_),
    .A1(\rtbdci.genblk1[15].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0704_ (.Y(_0301_),
    .A(\rtbdci.genblk1[12].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[13].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0705_ (.B1(net159),
    .Y(_0302_),
    .A1(\rtbdci.genblk1[12].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[13].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0706_ (.B1(_0302_),
    .Y(\rtbdci.genblk1[13].genblk1.combcgate_inst.Q ),
    .A2(_0301_),
    .A1(\rtbdci.genblk1[14].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0707_ (.Y(_0303_),
    .A(\rtbdci.genblk1[11].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[12].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0708_ (.B1(net159),
    .Y(_0304_),
    .A1(\rtbdci.genblk1[11].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[12].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0709_ (.B1(_0304_),
    .Y(\rtbdci.genblk1[12].genblk1.combcgate_inst.Q ),
    .A2(_0303_),
    .A1(\rtbdci.genblk1[13].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0710_ (.Y(_0305_),
    .A(\rtbdci.genblk1[10].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[11].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0711_ (.B1(net159),
    .Y(_0306_),
    .A1(\rtbdci.genblk1[10].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[11].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0712_ (.B1(_0306_),
    .Y(\rtbdci.genblk1[11].genblk1.combcgate_inst.Q ),
    .A2(_0305_),
    .A1(\rtbdci.genblk1[12].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0713_ (.Y(_0307_),
    .A(\rtbdci.genblk1[10].genblk1.combcgate_inst.A ),
    .B(\rtbdci.genblk1[10].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0714_ (.B1(net159),
    .Y(_0308_),
    .A1(\rtbdci.genblk1[10].genblk1.combcgate_inst.A ),
    .A2(\rtbdci.genblk1[10].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0715_ (.B1(_0308_),
    .Y(\rtbdci.genblk1[10].genblk1.combcgate_inst.Q ),
    .A2(_0307_),
    .A1(\rtbdci.genblk1[11].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0716_ (.Y(_0309_),
    .A(\rtbdci.genblk1[10].genblk1.combcgate_inst.A ),
    .B(\rtbdci.genblk1[8].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0717_ (.B1(net160),
    .Y(_0310_),
    .A1(\rtbdci.genblk1[10].genblk1.combcgate_inst.A ),
    .A2(\rtbdci.genblk1[8].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0718_ (.B1(_0310_),
    .Y(\rtbdci.genblk1[10].genblk1.combcgate_inst.A ),
    .A2(_0309_),
    .A1(\rtbdci.genblk1[10].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0719_ (.Y(_0311_),
    .A(\rtbdci.genblk1[7].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[8].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0720_ (.B1(net160),
    .Y(_0312_),
    .A1(\rtbdci.genblk1[7].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[8].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0721_ (.B1(_0312_),
    .Y(\rtbdci.genblk1[8].genblk1.combcgate_inst.Q ),
    .A2(_0311_),
    .A1(\rtbdci.genblk1[10].genblk1.combcgate_inst.A ));
 sg13g2_nand2_1 _0722_ (.Y(_0313_),
    .A(\rtbdci.genblk1[6].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[7].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0723_ (.B1(net159),
    .Y(_0314_),
    .A1(\rtbdci.genblk1[6].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[7].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0724_ (.B1(_0314_),
    .Y(\rtbdci.genblk1[7].genblk1.combcgate_inst.Q ),
    .A2(_0313_),
    .A1(\rtbdci.genblk1[8].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0725_ (.Y(_0315_),
    .A(\rtbdci.genblk1[5].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[6].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0726_ (.B1(net162),
    .Y(_0316_),
    .A1(\rtbdci.genblk1[5].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[6].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0727_ (.B1(_0316_),
    .Y(\rtbdci.genblk1[6].genblk1.combcgate_inst.Q ),
    .A2(_0315_),
    .A1(\rtbdci.genblk1[7].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0728_ (.Y(_0317_),
    .A(\rtbdci.genblk1[4].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[5].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0729_ (.B1(net162),
    .Y(_0318_),
    .A1(\rtbdci.genblk1[4].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[5].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0730_ (.B1(_0318_),
    .Y(\rtbdci.genblk1[5].genblk1.combcgate_inst.Q ),
    .A2(_0317_),
    .A1(\rtbdci.genblk1[6].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0731_ (.Y(_0319_),
    .A(\rtbdci.genblk1[3].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[4].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0732_ (.B1(net162),
    .Y(_0320_),
    .A1(\rtbdci.genblk1[3].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[4].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0733_ (.B1(_0320_),
    .Y(\rtbdci.genblk1[4].genblk1.combcgate_inst.Q ),
    .A2(_0319_),
    .A1(\rtbdci.genblk1[5].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0734_ (.Y(_0321_),
    .A(\rtbdci.genblk1[2].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[3].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0735_ (.B1(net162),
    .Y(_0322_),
    .A1(\rtbdci.genblk1[2].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[3].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0736_ (.B1(_0322_),
    .Y(\rtbdci.genblk1[3].genblk1.combcgate_inst.Q ),
    .A2(_0321_),
    .A1(\rtbdci.genblk1[4].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0737_ (.Y(_0323_),
    .A(\rtbdci.genblk1[1].genblk1.combcgate_inst.Q ),
    .B(\rtbdci.genblk1[2].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0738_ (.B1(net163),
    .Y(_0324_),
    .A1(\rtbdci.genblk1[1].genblk1.combcgate_inst.Q ),
    .A2(\rtbdci.genblk1[2].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0739_ (.B1(_0324_),
    .Y(\rtbdci.genblk1[2].genblk1.combcgate_inst.Q ),
    .A2(_0323_),
    .A1(\rtbdci.genblk1[3].genblk1.combcgate_inst.Q ));
 sg13g2_nor2b_1 _0740_ (.A(R4c),
    .B_N(\r4ci.genblk1[2].genblk1.combcgate_inst.Q ),
    .Y(_0325_));
 sg13g2_nor2_1 _0741_ (.A(\r4ci.genblk1[0].genblk1.combcgate_inst.A ),
    .B(_0325_),
    .Y(_0326_));
 sg13g2_nor2b_1 _0742_ (.A(\r4ci.genblk1[2].genblk1.combcgate_inst.Q ),
    .B_N(R4c),
    .Y(_0327_));
 sg13g2_nor3_1 _0743_ (.A(net140),
    .B(_0326_),
    .C(_0327_),
    .Y(\r4ci.genblk1[0].genblk1.combcgate_inst.A ));
 sg13g2_nor2_1 _0744_ (.A(\r4ci.genblk1[1].genblk1.combcgate_inst.Q ),
    .B(_0327_),
    .Y(_0328_));
 sg13g2_nor3_1 _0745_ (.A(net140),
    .B(_0325_),
    .C(_0328_),
    .Y(\r4ci.genblk1[1].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0746_ (.B1(net165),
    .Y(_0329_),
    .A1(_0180_),
    .A2(\r4ci.genblk1[1].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0747_ (.Y(_0330_),
    .A(_0180_),
    .B(\r4ci.genblk1[1].genblk1.combcgate_inst.Q ));
 sg13g2_a21o_1 _0748_ (.A2(_0330_),
    .A1(R4c),
    .B1(_0329_),
    .X(R4c));
 sg13g2_a21oi_1 _0749_ (.A1(_0181_),
    .A2(_0330_),
    .Y(\r4ci.genblk1[2].genblk1.combcgate_inst.Q ),
    .B1(_0329_));
 sg13g2_nand2_1 _0750_ (.Y(_0331_),
    .A(\r16ci.genblk1[0].genblk1.combcgate_inst.A ),
    .B(\r16ci.genblk1[14].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0751_ (.B1(net165),
    .Y(_0332_),
    .A1(\r16ci.genblk1[0].genblk1.combcgate_inst.A ),
    .A2(\r16ci.genblk1[14].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0752_ (.B1(_0332_),
    .Y(\r16ci.genblk1[0].genblk1.combcgate_inst.A ),
    .A2(_0331_),
    .A1(R16c));
 sg13g2_nand2_1 _0753_ (.Y(_0333_),
    .A(\r16ci.genblk1[13].genblk1.combcgate_inst.Q ),
    .B(\r16ci.genblk1[14].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0754_ (.B1(net165),
    .Y(_0334_),
    .A1(\r16ci.genblk1[13].genblk1.combcgate_inst.Q ),
    .A2(\r16ci.genblk1[14].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0755_ (.B1(_0334_),
    .Y(\r16ci.genblk1[14].genblk1.combcgate_inst.Q ),
    .A2(_0333_),
    .A1(\r16ci.genblk1[0].genblk1.combcgate_inst.A ));
 sg13g2_nand2_1 _0756_ (.Y(_0335_),
    .A(\r16ci.genblk1[12].genblk1.combcgate_inst.Q ),
    .B(\r16ci.genblk1[13].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0757_ (.B1(net165),
    .Y(_0336_),
    .A1(\r16ci.genblk1[12].genblk1.combcgate_inst.Q ),
    .A2(\r16ci.genblk1[13].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0758_ (.B1(_0336_),
    .Y(\r16ci.genblk1[13].genblk1.combcgate_inst.Q ),
    .A2(_0335_),
    .A1(\r16ci.genblk1[14].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0759_ (.Y(_0337_),
    .A(\r16ci.genblk1[11].genblk1.combcgate_inst.Q ),
    .B(\r16ci.genblk1[12].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0760_ (.B1(net166),
    .Y(_0338_),
    .A1(\r16ci.genblk1[11].genblk1.combcgate_inst.Q ),
    .A2(\r16ci.genblk1[12].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0761_ (.B1(_0338_),
    .Y(\r16ci.genblk1[12].genblk1.combcgate_inst.Q ),
    .A2(_0337_),
    .A1(\r16ci.genblk1[13].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0762_ (.Y(_0339_),
    .A(\r16ci.genblk1[10].genblk1.combcgate_inst.Q ),
    .B(\r16ci.genblk1[11].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0763_ (.B1(net160),
    .Y(_0340_),
    .A1(\r16ci.genblk1[10].genblk1.combcgate_inst.Q ),
    .A2(\r16ci.genblk1[11].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0764_ (.B1(_0340_),
    .Y(\r16ci.genblk1[11].genblk1.combcgate_inst.Q ),
    .A2(_0339_),
    .A1(\r16ci.genblk1[12].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0765_ (.Y(_0341_),
    .A(\r16ci.genblk1[10].genblk1.combcgate_inst.A ),
    .B(\r16ci.genblk1[10].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0766_ (.B1(net160),
    .Y(_0342_),
    .A1(\r16ci.genblk1[10].genblk1.combcgate_inst.A ),
    .A2(\r16ci.genblk1[10].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0767_ (.B1(_0342_),
    .Y(\r16ci.genblk1[10].genblk1.combcgate_inst.Q ),
    .A2(_0341_),
    .A1(\r16ci.genblk1[11].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0768_ (.Y(_0343_),
    .A(\r16ci.genblk1[10].genblk1.combcgate_inst.A ),
    .B(\r16ci.genblk1[8].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0769_ (.B1(net160),
    .Y(_0344_),
    .A1(\r16ci.genblk1[10].genblk1.combcgate_inst.A ),
    .A2(\r16ci.genblk1[8].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0770_ (.B1(_0344_),
    .Y(\r16ci.genblk1[10].genblk1.combcgate_inst.A ),
    .A2(_0343_),
    .A1(\r16ci.genblk1[10].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0771_ (.Y(_0345_),
    .A(\r16ci.genblk1[7].genblk1.combcgate_inst.Q ),
    .B(\r16ci.genblk1[8].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0772_ (.B1(net164),
    .Y(_0346_),
    .A1(\r16ci.genblk1[7].genblk1.combcgate_inst.Q ),
    .A2(\r16ci.genblk1[8].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0773_ (.B1(_0346_),
    .Y(\r16ci.genblk1[8].genblk1.combcgate_inst.Q ),
    .A2(_0345_),
    .A1(\r16ci.genblk1[10].genblk1.combcgate_inst.A ));
 sg13g2_nand2_1 _0774_ (.Y(_0347_),
    .A(\r16ci.genblk1[6].genblk1.combcgate_inst.Q ),
    .B(\r16ci.genblk1[7].genblk1.combcgate_inst.Q ));
 sg13g2_o21ai_1 _0775_ (.B1(net164),
    .Y(_0348_),
    .A1(\r16ci.genblk1[6].genblk1.combcgate_inst.Q ),
    .A2(\r16ci.genblk1[7].genblk1.combcgate_inst.Q ));
 sg13g2_a21oi_2 _0776_ (.B1(_0348_),
    .Y(\r16ci.genblk1[7].genblk1.combcgate_inst.Q ),
    .A2(_0347_),
    .A1(\r16ci.genblk1[8].genblk1.combcgate_inst.Q ));
 sg13g2_nand2_1 _0777_ (.Y(_0046_),
    .A(net166),
    .B(_0175_));
 sg13g2_nand2_1 _0778_ (.Y(_0040_),
    .A(net174),
    .B(_0176_));
 sg13g2_nand2_1 _0779_ (.Y(_0008_),
    .A(net175),
    .B(_0177_));
 sg13g2_and2_1 _0780_ (.A(net166),
    .B(\rtbdli.genblk1[62].latchcgate_inst.Q ),
    .X(_0164_));
 sg13g2_xor2_1 _0781_ (.B(RBigl),
    .A(\rtbdli.genblk1[62].latchcgate_inst.Q ),
    .X(_0349_));
 sg13g2_nor2_1 _0782_ (.A(net140),
    .B(_0349_),
    .Y(_0165_));
 sg13g2_nand2_1 _0783_ (.Y(_0350_),
    .A(net166),
    .B(\rtbdli.genblk1[61].latchcgate_inst.Q ));
 sg13g2_inv_1 _0784_ (.Y(_0162_),
    .A(_0350_));
 sg13g2_a22oi_1 _0785_ (.Y(_0163_),
    .B1(_0046_),
    .B2(_0350_),
    .A2(\rtbdli.genblk1[61].latchcgate_inst.Q ),
    .A1(_0175_));
 sg13g2_and2_1 _0786_ (.A(net166),
    .B(\rtbdli.genblk1[60].latchcgate_inst.Q ),
    .X(_0160_));
 sg13g2_xor2_1 _0787_ (.B(\rtbdli.genblk1[60].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[62].latchcgate_inst.Q ),
    .X(_0351_));
 sg13g2_nor2_1 _0788_ (.A(net140),
    .B(_0351_),
    .Y(_0161_));
 sg13g2_and2_1 _0789_ (.A(net166),
    .B(\rtbdli.genblk1[59].latchcgate_inst.Q ),
    .X(_0158_));
 sg13g2_xor2_1 _0790_ (.B(\rtbdli.genblk1[59].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[61].latchcgate_inst.Q ),
    .X(_0352_));
 sg13g2_nor2_1 _0791_ (.A(net140),
    .B(_0352_),
    .Y(_0159_));
 sg13g2_and2_1 _0792_ (.A(net157),
    .B(\rtbdli.genblk1[58].latchcgate_inst.Q ),
    .X(_0154_));
 sg13g2_xor2_1 _0793_ (.B(\rtbdli.genblk1[58].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[60].latchcgate_inst.Q ),
    .X(_0353_));
 sg13g2_nor2_1 _0794_ (.A(net140),
    .B(_0353_),
    .Y(_0155_));
 sg13g2_and2_1 _0795_ (.A(net157),
    .B(\rtbdli.genblk1[57].latchcgate_inst.Q ),
    .X(_0152_));
 sg13g2_xor2_1 _0796_ (.B(\rtbdli.genblk1[57].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[59].latchcgate_inst.Q ),
    .X(_0354_));
 sg13g2_nor2_1 _0797_ (.A(net137),
    .B(_0354_),
    .Y(_0153_));
 sg13g2_and2_1 _0798_ (.A(net157),
    .B(\rtbdli.genblk1[56].latchcgate_inst.Q ),
    .X(_0150_));
 sg13g2_xor2_1 _0799_ (.B(\rtbdli.genblk1[56].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[58].latchcgate_inst.Q ),
    .X(_0355_));
 sg13g2_nor2_1 _0800_ (.A(net137),
    .B(_0355_),
    .Y(_0151_));
 sg13g2_and2_1 _0801_ (.A(net158),
    .B(\rtbdli.genblk1[55].latchcgate_inst.Q ),
    .X(_0148_));
 sg13g2_xor2_1 _0802_ (.B(\rtbdli.genblk1[55].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[57].latchcgate_inst.Q ),
    .X(_0356_));
 sg13g2_nor2_1 _0803_ (.A(net137),
    .B(_0356_),
    .Y(_0149_));
 sg13g2_and2_1 _0804_ (.A(net158),
    .B(\rtbdli.genblk1[54].latchcgate_inst.Q ),
    .X(_0146_));
 sg13g2_xor2_1 _0805_ (.B(\rtbdli.genblk1[54].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[56].latchcgate_inst.Q ),
    .X(_0357_));
 sg13g2_nor2_1 _0806_ (.A(net137),
    .B(_0357_),
    .Y(_0147_));
 sg13g2_and2_1 _0807_ (.A(net157),
    .B(\rtbdli.genblk1[53].latchcgate_inst.Q ),
    .X(_0144_));
 sg13g2_xor2_1 _0808_ (.B(\rtbdli.genblk1[53].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[55].latchcgate_inst.Q ),
    .X(_0358_));
 sg13g2_nor2_1 _0809_ (.A(net137),
    .B(_0358_),
    .Y(_0145_));
 sg13g2_and2_1 _0810_ (.A(net157),
    .B(\rtbdli.genblk1[52].latchcgate_inst.Q ),
    .X(_0142_));
 sg13g2_xor2_1 _0811_ (.B(\rtbdli.genblk1[52].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[54].latchcgate_inst.Q ),
    .X(_0359_));
 sg13g2_nor2_1 _0812_ (.A(net137),
    .B(_0359_),
    .Y(_0143_));
 sg13g2_and2_1 _0813_ (.A(net156),
    .B(\rtbdli.genblk1[51].latchcgate_inst.Q ),
    .X(_0140_));
 sg13g2_xor2_1 _0814_ (.B(\rtbdli.genblk1[51].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[53].latchcgate_inst.Q ),
    .X(_0360_));
 sg13g2_nor2_1 _0815_ (.A(net136),
    .B(_0360_),
    .Y(_0141_));
 sg13g2_and2_1 _0816_ (.A(net156),
    .B(\rtbdli.genblk1[50].latchcgate_inst.Q ),
    .X(_0138_));
 sg13g2_xor2_1 _0817_ (.B(\rtbdli.genblk1[50].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[52].latchcgate_inst.Q ),
    .X(_0361_));
 sg13g2_nor2_1 _0818_ (.A(net136),
    .B(_0361_),
    .Y(_0139_));
 sg13g2_and2_1 _0819_ (.A(net156),
    .B(\rtbdli.genblk1[49].latchcgate_inst.Q ),
    .X(_0136_));
 sg13g2_xor2_1 _0820_ (.B(\rtbdli.genblk1[49].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[51].latchcgate_inst.Q ),
    .X(_0362_));
 sg13g2_nor2_1 _0821_ (.A(net136),
    .B(_0362_),
    .Y(_0137_));
 sg13g2_and2_1 _0822_ (.A(net156),
    .B(\rtbdli.genblk1[48].latchcgate_inst.Q ),
    .X(_0132_));
 sg13g2_xor2_1 _0823_ (.B(\rtbdli.genblk1[48].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[50].latchcgate_inst.Q ),
    .X(_0363_));
 sg13g2_nor2_1 _0824_ (.A(net136),
    .B(_0363_),
    .Y(_0133_));
 sg13g2_and2_1 _0825_ (.A(net156),
    .B(\rtbdli.genblk1[47].latchcgate_inst.Q ),
    .X(_0130_));
 sg13g2_xor2_1 _0826_ (.B(\rtbdli.genblk1[47].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[49].latchcgate_inst.Q ),
    .X(_0364_));
 sg13g2_nor2_1 _0827_ (.A(net136),
    .B(_0364_),
    .Y(_0131_));
 sg13g2_and2_1 _0828_ (.A(net156),
    .B(\rtbdli.genblk1[46].latchcgate_inst.Q ),
    .X(_0128_));
 sg13g2_xor2_1 _0829_ (.B(\rtbdli.genblk1[46].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[48].latchcgate_inst.Q ),
    .X(_0365_));
 sg13g2_nor2_1 _0830_ (.A(net136),
    .B(_0365_),
    .Y(_0129_));
 sg13g2_and2_1 _0831_ (.A(net156),
    .B(\rtbdli.genblk1[45].latchcgate_inst.Q ),
    .X(_0126_));
 sg13g2_xor2_1 _0832_ (.B(\rtbdli.genblk1[45].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[47].latchcgate_inst.Q ),
    .X(_0366_));
 sg13g2_nor2_1 _0833_ (.A(net136),
    .B(_0366_),
    .Y(_0127_));
 sg13g2_and2_1 _0834_ (.A(net156),
    .B(\rtbdli.genblk1[44].latchcgate_inst.Q ),
    .X(_0124_));
 sg13g2_xor2_1 _0835_ (.B(\rtbdli.genblk1[44].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[46].latchcgate_inst.Q ),
    .X(_0367_));
 sg13g2_nor2_1 _0836_ (.A(net137),
    .B(_0367_),
    .Y(_0125_));
 sg13g2_and2_1 _0837_ (.A(net157),
    .B(\rtbdli.genblk1[43].latchcgate_inst.Q ),
    .X(_0122_));
 sg13g2_xor2_1 _0838_ (.B(\rtbdli.genblk1[43].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[45].latchcgate_inst.Q ),
    .X(_0368_));
 sg13g2_nor2_1 _0839_ (.A(net136),
    .B(_0368_),
    .Y(_0123_));
 sg13g2_and2_1 _0840_ (.A(net168),
    .B(\rtbdli.genblk1[42].latchcgate_inst.Q ),
    .X(_0120_));
 sg13g2_xor2_1 _0841_ (.B(\rtbdli.genblk1[42].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[44].latchcgate_inst.Q ),
    .X(_0369_));
 sg13g2_nor2_1 _0842_ (.A(net138),
    .B(_0369_),
    .Y(_0121_));
 sg13g2_and2_1 _0843_ (.A(net168),
    .B(\rtbdli.genblk1[41].latchcgate_inst.Q ),
    .X(_0118_));
 sg13g2_xor2_1 _0844_ (.B(\rtbdli.genblk1[41].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[43].latchcgate_inst.Q ),
    .X(_0370_));
 sg13g2_nor2_1 _0845_ (.A(net138),
    .B(_0370_),
    .Y(_0119_));
 sg13g2_and2_1 _0846_ (.A(net168),
    .B(\rtbdli.genblk1[40].latchcgate_inst.Q ),
    .X(_0116_));
 sg13g2_xor2_1 _0847_ (.B(\rtbdli.genblk1[40].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[42].latchcgate_inst.Q ),
    .X(_0371_));
 sg13g2_nor2_1 _0848_ (.A(net138),
    .B(_0371_),
    .Y(_0117_));
 sg13g2_and2_1 _0849_ (.A(net168),
    .B(\rtbdli.genblk1[39].latchcgate_inst.Q ),
    .X(_0114_));
 sg13g2_xor2_1 _0850_ (.B(\rtbdli.genblk1[39].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[41].latchcgate_inst.Q ),
    .X(_0372_));
 sg13g2_nor2_1 _0851_ (.A(net138),
    .B(_0372_),
    .Y(_0115_));
 sg13g2_and2_1 _0852_ (.A(net168),
    .B(\rtbdli.genblk1[38].latchcgate_inst.Q ),
    .X(_0110_));
 sg13g2_xor2_1 _0853_ (.B(\rtbdli.genblk1[38].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[40].latchcgate_inst.Q ),
    .X(_0373_));
 sg13g2_nor2_1 _0854_ (.A(net138),
    .B(_0373_),
    .Y(_0111_));
 sg13g2_and2_1 _0855_ (.A(net168),
    .B(\rtbdli.genblk1[37].latchcgate_inst.Q ),
    .X(_0108_));
 sg13g2_xor2_1 _0856_ (.B(\rtbdli.genblk1[37].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[39].latchcgate_inst.Q ),
    .X(_0374_));
 sg13g2_nor2_1 _0857_ (.A(net138),
    .B(_0374_),
    .Y(_0109_));
 sg13g2_and2_1 _0858_ (.A(net169),
    .B(\rtbdli.genblk1[36].latchcgate_inst.Q ),
    .X(_0106_));
 sg13g2_xor2_1 _0859_ (.B(\rtbdli.genblk1[36].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[38].latchcgate_inst.Q ),
    .X(_0375_));
 sg13g2_nor2_1 _0860_ (.A(net139),
    .B(_0375_),
    .Y(_0107_));
 sg13g2_and2_1 _0861_ (.A(net169),
    .B(\rtbdli.genblk1[35].latchcgate_inst.Q ),
    .X(_0104_));
 sg13g2_xor2_1 _0862_ (.B(\rtbdli.genblk1[35].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[37].latchcgate_inst.Q ),
    .X(_0376_));
 sg13g2_nor2_1 _0863_ (.A(net145),
    .B(_0376_),
    .Y(_0105_));
 sg13g2_and2_1 _0864_ (.A(net169),
    .B(\rtbdli.genblk1[34].latchcgate_inst.Q ),
    .X(_0102_));
 sg13g2_xor2_1 _0865_ (.B(\rtbdli.genblk1[34].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[36].latchcgate_inst.Q ),
    .X(_0377_));
 sg13g2_nor2_1 _0866_ (.A(net145),
    .B(_0377_),
    .Y(_0103_));
 sg13g2_and2_1 _0867_ (.A(net171),
    .B(\rtbdli.genblk1[33].latchcgate_inst.Q ),
    .X(_0100_));
 sg13g2_xor2_1 _0868_ (.B(\rtbdli.genblk1[33].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[35].latchcgate_inst.Q ),
    .X(_0378_));
 sg13g2_nor2_1 _0869_ (.A(net142),
    .B(_0378_),
    .Y(_0101_));
 sg13g2_and2_1 _0870_ (.A(net170),
    .B(\rtbdli.genblk1[32].latchcgate_inst.Q ),
    .X(_0098_));
 sg13g2_xor2_1 _0871_ (.B(\rtbdli.genblk1[32].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[34].latchcgate_inst.Q ),
    .X(_0379_));
 sg13g2_nor2_1 _0872_ (.A(net142),
    .B(_0379_),
    .Y(_0099_));
 sg13g2_and2_1 _0873_ (.A(net170),
    .B(\rtbdli.genblk1[31].latchcgate_inst.Q ),
    .X(_0096_));
 sg13g2_xor2_1 _0874_ (.B(\rtbdli.genblk1[31].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[33].latchcgate_inst.Q ),
    .X(_0380_));
 sg13g2_nor2_1 _0875_ (.A(net142),
    .B(_0380_),
    .Y(_0097_));
 sg13g2_and2_1 _0876_ (.A(net170),
    .B(\rtbdli.genblk1[30].latchcgate_inst.Q ),
    .X(_0094_));
 sg13g2_xor2_1 _0877_ (.B(\rtbdli.genblk1[30].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[32].latchcgate_inst.Q ),
    .X(_0381_));
 sg13g2_nor2_1 _0878_ (.A(net142),
    .B(_0381_),
    .Y(_0095_));
 sg13g2_and2_1 _0879_ (.A(net170),
    .B(\rtbdli.genblk1[29].latchcgate_inst.Q ),
    .X(_0092_));
 sg13g2_xor2_1 _0880_ (.B(\rtbdli.genblk1[29].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[31].latchcgate_inst.Q ),
    .X(_0382_));
 sg13g2_nor2_1 _0881_ (.A(net142),
    .B(_0382_),
    .Y(_0093_));
 sg13g2_and2_1 _0882_ (.A(net170),
    .B(\rtbdli.genblk1[28].latchcgate_inst.Q ),
    .X(_0088_));
 sg13g2_xor2_1 _0883_ (.B(\rtbdli.genblk1[28].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[30].latchcgate_inst.Q ),
    .X(_0383_));
 sg13g2_nor2_1 _0884_ (.A(net143),
    .B(_0383_),
    .Y(_0089_));
 sg13g2_and2_1 _0885_ (.A(net172),
    .B(\rtbdli.genblk1[27].latchcgate_inst.Q ),
    .X(_0086_));
 sg13g2_xor2_1 _0886_ (.B(\rtbdli.genblk1[27].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[29].latchcgate_inst.Q ),
    .X(_0384_));
 sg13g2_nor2_1 _0887_ (.A(net143),
    .B(_0384_),
    .Y(_0087_));
 sg13g2_and2_1 _0888_ (.A(net170),
    .B(\rtbdli.genblk1[26].latchcgate_inst.Q ),
    .X(_0084_));
 sg13g2_xor2_1 _0889_ (.B(\rtbdli.genblk1[26].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[28].latchcgate_inst.Q ),
    .X(_0385_));
 sg13g2_nor2_1 _0890_ (.A(net143),
    .B(_0385_),
    .Y(_0085_));
 sg13g2_and2_1 _0891_ (.A(net172),
    .B(\rtbdli.genblk1[25].latchcgate_inst.Q ),
    .X(_0082_));
 sg13g2_xor2_1 _0892_ (.B(\rtbdli.genblk1[25].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[27].latchcgate_inst.Q ),
    .X(_0386_));
 sg13g2_nor2_1 _0893_ (.A(net143),
    .B(_0386_),
    .Y(_0083_));
 sg13g2_and2_1 _0894_ (.A(net170),
    .B(\rtbdli.genblk1[24].latchcgate_inst.Q ),
    .X(_0080_));
 sg13g2_xor2_1 _0895_ (.B(\rtbdli.genblk1[24].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[26].latchcgate_inst.Q ),
    .X(_0387_));
 sg13g2_nor2_1 _0896_ (.A(net143),
    .B(_0387_),
    .Y(_0081_));
 sg13g2_and2_1 _0897_ (.A(net170),
    .B(\rtbdli.genblk1[23].latchcgate_inst.Q ),
    .X(_0078_));
 sg13g2_xor2_1 _0898_ (.B(\rtbdli.genblk1[23].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[25].latchcgate_inst.Q ),
    .X(_0388_));
 sg13g2_nor2_1 _0899_ (.A(net143),
    .B(_0388_),
    .Y(_0079_));
 sg13g2_and2_1 _0900_ (.A(net171),
    .B(\rtbdli.genblk1[22].latchcgate_inst.Q ),
    .X(_0076_));
 sg13g2_xor2_1 _0901_ (.B(\rtbdli.genblk1[22].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[24].latchcgate_inst.Q ),
    .X(_0389_));
 sg13g2_nor2_1 _0902_ (.A(net143),
    .B(_0389_),
    .Y(_0077_));
 sg13g2_and2_1 _0903_ (.A(net172),
    .B(\rtbdli.genblk1[21].latchcgate_inst.Q ),
    .X(_0074_));
 sg13g2_xor2_1 _0904_ (.B(\rtbdli.genblk1[21].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[23].latchcgate_inst.Q ),
    .X(_0390_));
 sg13g2_nor2_1 _0905_ (.A(net144),
    .B(_0390_),
    .Y(_0075_));
 sg13g2_and2_1 _0906_ (.A(net171),
    .B(\rtbdli.genblk1[20].latchcgate_inst.Q ),
    .X(_0072_));
 sg13g2_xor2_1 _0907_ (.B(\rtbdli.genblk1[20].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[22].latchcgate_inst.Q ),
    .X(_0391_));
 sg13g2_nor2_1 _0908_ (.A(net144),
    .B(_0391_),
    .Y(_0073_));
 sg13g2_and2_1 _0909_ (.A(net171),
    .B(\rtbdli.genblk1[19].latchcgate_inst.Q ),
    .X(_0070_));
 sg13g2_xor2_1 _0910_ (.B(\rtbdli.genblk1[19].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[21].latchcgate_inst.Q ),
    .X(_0392_));
 sg13g2_nor2_1 _0911_ (.A(net144),
    .B(_0392_),
    .Y(_0071_));
 sg13g2_and2_1 _0912_ (.A(net171),
    .B(\rtbdli.genblk1[18].latchcgate_inst.Q ),
    .X(_0066_));
 sg13g2_xor2_1 _0913_ (.B(\rtbdli.genblk1[18].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[20].latchcgate_inst.Q ),
    .X(_0393_));
 sg13g2_nor2_1 _0914_ (.A(net144),
    .B(_0393_),
    .Y(_0067_));
 sg13g2_and2_1 _0915_ (.A(net176),
    .B(\rtbdli.genblk1[17].latchcgate_inst.Q ),
    .X(_0064_));
 sg13g2_xor2_1 _0916_ (.B(\rtbdli.genblk1[17].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[19].latchcgate_inst.Q ),
    .X(_0394_));
 sg13g2_nor2_1 _0917_ (.A(net146),
    .B(_0394_),
    .Y(_0065_));
 sg13g2_and2_1 _0918_ (.A(net176),
    .B(\rtbdli.genblk1[16].latchcgate_inst.Q ),
    .X(_0062_));
 sg13g2_xor2_1 _0919_ (.B(\rtbdli.genblk1[16].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[18].latchcgate_inst.Q ),
    .X(_0395_));
 sg13g2_nor2_1 _0920_ (.A(net146),
    .B(_0395_),
    .Y(_0063_));
 sg13g2_and2_1 _0921_ (.A(net171),
    .B(\rtbdli.genblk1[15].latchcgate_inst.Q ),
    .X(_0060_));
 sg13g2_xor2_1 _0922_ (.B(\rtbdli.genblk1[15].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[17].latchcgate_inst.Q ),
    .X(_0396_));
 sg13g2_nor2_1 _0923_ (.A(net143),
    .B(_0396_),
    .Y(_0061_));
 sg13g2_and2_1 _0924_ (.A(net171),
    .B(\rtbdli.genblk1[14].latchcgate_inst.Q ),
    .X(_0058_));
 sg13g2_xor2_1 _0925_ (.B(\rtbdli.genblk1[14].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[16].latchcgate_inst.Q ),
    .X(_0397_));
 sg13g2_nor2_1 _0926_ (.A(net146),
    .B(_0397_),
    .Y(_0059_));
 sg13g2_and2_1 _0927_ (.A(net171),
    .B(\rtbdli.genblk1[13].latchcgate_inst.Q ),
    .X(_0056_));
 sg13g2_xor2_1 _0928_ (.B(\rtbdli.genblk1[13].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[15].latchcgate_inst.Q ),
    .X(_0398_));
 sg13g2_nor2_1 _0929_ (.A(net142),
    .B(_0398_),
    .Y(_0057_));
 sg13g2_and2_1 _0930_ (.A(net168),
    .B(\rtbdli.genblk1[12].latchcgate_inst.Q ),
    .X(_0054_));
 sg13g2_xor2_1 _0931_ (.B(\rtbdli.genblk1[12].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[14].latchcgate_inst.Q ),
    .X(_0399_));
 sg13g2_nor2_1 _0932_ (.A(net142),
    .B(_0399_),
    .Y(_0055_));
 sg13g2_and2_1 _0933_ (.A(net173),
    .B(\rtbdli.genblk1[11].latchcgate_inst.Q ),
    .X(_0052_));
 sg13g2_xor2_1 _0934_ (.B(\rtbdli.genblk1[11].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[13].latchcgate_inst.Q ),
    .X(_0400_));
 sg13g2_nor2_1 _0935_ (.A(net148),
    .B(_0400_),
    .Y(_0053_));
 sg13g2_and2_1 _0936_ (.A(net168),
    .B(\rtbdli.genblk1[10].latchcgate_inst.Q ),
    .X(_0050_));
 sg13g2_xor2_1 _0937_ (.B(\rtbdli.genblk1[10].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[12].latchcgate_inst.Q ),
    .X(_0401_));
 sg13g2_nor2_1 _0938_ (.A(net142),
    .B(_0401_),
    .Y(_0051_));
 sg13g2_and2_1 _0939_ (.A(net169),
    .B(\rtbdli.genblk1[10].latchcgate_inst.A ),
    .X(_0048_));
 sg13g2_xor2_1 _0940_ (.B(\rtbdli.genblk1[10].latchcgate_inst.A ),
    .A(\rtbdli.genblk1[11].latchcgate_inst.Q ),
    .X(_0402_));
 sg13g2_nor2_1 _0941_ (.A(net139),
    .B(_0402_),
    .Y(_0049_));
 sg13g2_and2_1 _0942_ (.A(net169),
    .B(\rtbdli.genblk1[8].latchcgate_inst.Q ),
    .X(_0172_));
 sg13g2_xor2_1 _0943_ (.B(\rtbdli.genblk1[8].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[10].latchcgate_inst.Q ),
    .X(_0403_));
 sg13g2_nor2_1 _0944_ (.A(net138),
    .B(_0403_),
    .Y(_0173_));
 sg13g2_and2_1 _0945_ (.A(net157),
    .B(\rtbdli.genblk1[7].latchcgate_inst.Q ),
    .X(_0170_));
 sg13g2_xor2_1 _0946_ (.B(\rtbdli.genblk1[7].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[10].latchcgate_inst.A ),
    .X(_0404_));
 sg13g2_nor2_1 _0947_ (.A(net139),
    .B(_0404_),
    .Y(_0171_));
 sg13g2_and2_1 _0948_ (.A(net166),
    .B(\rtbdli.genblk1[6].latchcgate_inst.Q ),
    .X(_0168_));
 sg13g2_xor2_1 _0949_ (.B(\rtbdli.genblk1[6].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[8].latchcgate_inst.Q ),
    .X(_0405_));
 sg13g2_nor2_1 _0950_ (.A(net138),
    .B(_0405_),
    .Y(_0169_));
 sg13g2_and2_1 _0951_ (.A(net173),
    .B(\rtbdli.genblk1[5].latchcgate_inst.Q ),
    .X(_0166_));
 sg13g2_xor2_1 _0952_ (.B(\rtbdli.genblk1[5].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[7].latchcgate_inst.Q ),
    .X(_0406_));
 sg13g2_nor2_1 _0953_ (.A(net141),
    .B(_0406_),
    .Y(_0167_));
 sg13g2_and2_1 _0954_ (.A(net173),
    .B(\rtbdli.genblk1[4].latchcgate_inst.Q ),
    .X(_0156_));
 sg13g2_xor2_1 _0955_ (.B(\rtbdli.genblk1[4].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[6].latchcgate_inst.Q ),
    .X(_0407_));
 sg13g2_nor2_1 _0956_ (.A(net140),
    .B(_0407_),
    .Y(_0157_));
 sg13g2_and2_1 _0957_ (.A(net173),
    .B(\rtbdli.genblk1[3].latchcgate_inst.Q ),
    .X(_0134_));
 sg13g2_xor2_1 _0958_ (.B(\rtbdli.genblk1[3].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[5].latchcgate_inst.Q ),
    .X(_0408_));
 sg13g2_nor2_1 _0959_ (.A(net141),
    .B(_0408_),
    .Y(_0135_));
 sg13g2_and2_1 _0960_ (.A(net173),
    .B(\rtbdli.genblk1[2].latchcgate_inst.Q ),
    .X(_0112_));
 sg13g2_xor2_1 _0961_ (.B(\rtbdli.genblk1[2].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[4].latchcgate_inst.Q ),
    .X(_0409_));
 sg13g2_nor2_1 _0962_ (.A(net141),
    .B(_0409_),
    .Y(_0113_));
 sg13g2_nand2_1 _0963_ (.Y(_0410_),
    .A(net166),
    .B(\rtbdli.genblk1[1].latchcgate_inst.Q ));
 sg13g2_inv_1 _0964_ (.Y(_0090_),
    .A(_0410_));
 sg13g2_xor2_1 _0965_ (.B(\rtbdli.genblk1[1].latchcgate_inst.Q ),
    .A(\rtbdli.genblk1[3].latchcgate_inst.Q ),
    .X(_0411_));
 sg13g2_nor2_1 _0966_ (.A(net141),
    .B(_0411_),
    .Y(_0091_));
 sg13g2_and2_1 _0967_ (.A(net167),
    .B(RBigl),
    .X(_0068_));
 sg13g2_xor2_1 _0968_ (.B(\rtbdli.genblk1[2].latchcgate_inst.Q ),
    .A(RBigl),
    .X(_0412_));
 sg13g2_nor2_1 _0969_ (.A(net141),
    .B(_0412_),
    .Y(_0069_));
 sg13g2_a22oi_1 _0970_ (.Y(_0047_),
    .B1(_0046_),
    .B2(_0410_),
    .A2(\rtbdli.genblk1[1].latchcgate_inst.Q ),
    .A1(_0175_));
 sg13g2_a21oi_1 _0971_ (.A1(net2),
    .A2(net1),
    .Y(_0413_),
    .B1(net147));
 sg13g2_nor2_1 _0972_ (.A(net2),
    .B(net1),
    .Y(_0414_));
 sg13g2_nor2b_1 _0973_ (.A(_0414_),
    .B_N(_0413_),
    .Y(_0007_));
 sg13g2_and2_1 _0974_ (.A(net175),
    .B(net1),
    .X(_0006_));
 sg13g2_o21ai_1 _0975_ (.B1(_0413_),
    .Y(Qc),
    .A1(_0182_),
    .A2(_0414_));
 sg13g2_and2_1 _0976_ (.A(net174),
    .B(\r4li.genblk1[2].latchcgate_inst.Q ),
    .X(_0045_));
 sg13g2_xor2_1 _0977_ (.B(R4l),
    .A(\r4li.genblk1[2].latchcgate_inst.Q ),
    .X(_0415_));
 sg13g2_nor2_1 _0978_ (.A(net140),
    .B(_0415_),
    .Y(_0043_));
 sg13g2_nand2_1 _0979_ (.Y(_0416_),
    .A(net174),
    .B(\r4li.genblk1[1].latchcgate_inst.Q ));
 sg13g2_inv_1 _0980_ (.Y(_0044_),
    .A(_0416_));
 sg13g2_a22oi_1 _0981_ (.Y(_0041_),
    .B1(_0040_),
    .B2(_0416_),
    .A2(\r4li.genblk1[1].latchcgate_inst.Q ),
    .A1(_0176_));
 sg13g2_and2_1 _0982_ (.A(net173),
    .B(R4l),
    .X(_0042_));
 sg13g2_and2_1 _0983_ (.A(net174),
    .B(\r16li.genblk1[14].latchcgate_inst.Q ),
    .X(_0020_));
 sg13g2_xor2_1 _0984_ (.B(R16l),
    .A(\r16li.genblk1[14].latchcgate_inst.Q ),
    .X(_0417_));
 sg13g2_nor2_1 _0985_ (.A(net148),
    .B(_0417_),
    .Y(_0021_));
 sg13g2_nand2_1 _0986_ (.Y(_0418_),
    .A(net173),
    .B(\r16li.genblk1[13].latchcgate_inst.Q ));
 sg13g2_inv_1 _0987_ (.Y(_0018_),
    .A(_0418_));
 sg13g2_a22oi_1 _0988_ (.Y(_0019_),
    .B1(_0008_),
    .B2(_0418_),
    .A2(\r16li.genblk1[13].latchcgate_inst.Q ),
    .A1(_0177_));
 sg13g2_and2_1 _0989_ (.A(net173),
    .B(\r16li.genblk1[12].latchcgate_inst.Q ),
    .X(_0016_));
 sg13g2_xor2_1 _0990_ (.B(\r16li.genblk1[12].latchcgate_inst.Q ),
    .A(\r16li.genblk1[14].latchcgate_inst.Q ),
    .X(_0419_));
 sg13g2_nor2_1 _0991_ (.A(net148),
    .B(_0419_),
    .Y(_0017_));
 sg13g2_and2_1 _0992_ (.A(net176),
    .B(\r16li.genblk1[11].latchcgate_inst.Q ),
    .X(_0014_));
 sg13g2_xor2_1 _0993_ (.B(\r16li.genblk1[11].latchcgate_inst.Q ),
    .A(\r16li.genblk1[13].latchcgate_inst.Q ),
    .X(_0420_));
 sg13g2_nor2_1 _0994_ (.A(net148),
    .B(_0420_),
    .Y(_0015_));
 sg13g2_and2_1 _0995_ (.A(net176),
    .B(\r16li.genblk1[10].latchcgate_inst.Q ),
    .X(_0012_));
 sg13g2_xor2_1 _0996_ (.B(\r16li.genblk1[10].latchcgate_inst.Q ),
    .A(\r16li.genblk1[12].latchcgate_inst.Q ),
    .X(_0421_));
 sg13g2_nor2_1 _0997_ (.A(net148),
    .B(_0421_),
    .Y(_0013_));
 sg13g2_and2_1 _0998_ (.A(net176),
    .B(\r16li.genblk1[10].latchcgate_inst.A ),
    .X(_0010_));
 sg13g2_xor2_1 _0999_ (.B(\r16li.genblk1[10].latchcgate_inst.A ),
    .A(\r16li.genblk1[11].latchcgate_inst.Q ),
    .X(_0422_));
 sg13g2_nor2_1 _1000_ (.A(net146),
    .B(_0422_),
    .Y(_0011_));
 sg13g2_and2_1 _1001_ (.A(net176),
    .B(\r16li.genblk1[8].latchcgate_inst.Q ),
    .X(_0038_));
 sg13g2_xor2_1 _1002_ (.B(\r16li.genblk1[8].latchcgate_inst.Q ),
    .A(\r16li.genblk1[10].latchcgate_inst.Q ),
    .X(_0423_));
 sg13g2_nor2_1 _1003_ (.A(net146),
    .B(_0423_),
    .Y(_0039_));
 sg13g2_and2_1 _1004_ (.A(net176),
    .B(\r16li.genblk1[7].latchcgate_inst.Q ),
    .X(_0036_));
 sg13g2_xor2_1 _1005_ (.B(\r16li.genblk1[7].latchcgate_inst.Q ),
    .A(\r16li.genblk1[10].latchcgate_inst.A ),
    .X(_0424_));
 sg13g2_nor2_1 _1006_ (.A(net146),
    .B(_0424_),
    .Y(_0037_));
 sg13g2_and2_1 _1007_ (.A(net177),
    .B(\r16li.genblk1[6].latchcgate_inst.Q ),
    .X(_0034_));
 sg13g2_xor2_1 _1008_ (.B(\r16li.genblk1[6].latchcgate_inst.Q ),
    .A(\r16li.genblk1[8].latchcgate_inst.Q ),
    .X(_0425_));
 sg13g2_nor2_1 _1009_ (.A(net146),
    .B(_0425_),
    .Y(_0035_));
 sg13g2_and2_1 _1010_ (.A(net175),
    .B(\r16li.genblk1[5].latchcgate_inst.Q ),
    .X(_0032_));
 sg13g2_xor2_1 _1011_ (.B(\r16li.genblk1[5].latchcgate_inst.Q ),
    .A(\r16li.genblk1[7].latchcgate_inst.Q ),
    .X(_0426_));
 sg13g2_nor2_1 _1012_ (.A(net147),
    .B(_0426_),
    .Y(_0033_));
 sg13g2_and2_1 _1013_ (.A(net175),
    .B(\r16li.genblk1[4].latchcgate_inst.Q ),
    .X(_0030_));
 sg13g2_xor2_1 _1014_ (.B(\r16li.genblk1[4].latchcgate_inst.Q ),
    .A(\r16li.genblk1[6].latchcgate_inst.Q ),
    .X(_0427_));
 sg13g2_nor2_1 _1015_ (.A(net146),
    .B(_0427_),
    .Y(_0031_));
 sg13g2_and2_1 _1016_ (.A(net175),
    .B(\r16li.genblk1[3].latchcgate_inst.Q ),
    .X(_0028_));
 sg13g2_xor2_1 _1017_ (.B(\r16li.genblk1[3].latchcgate_inst.Q ),
    .A(\r16li.genblk1[5].latchcgate_inst.Q ),
    .X(_0428_));
 sg13g2_nor2_1 _1018_ (.A(net147),
    .B(_0428_),
    .Y(_0029_));
 sg13g2_and2_1 _1019_ (.A(net175),
    .B(\r16li.genblk1[2].latchcgate_inst.Q ),
    .X(_0026_));
 sg13g2_xor2_1 _1020_ (.B(\r16li.genblk1[2].latchcgate_inst.Q ),
    .A(\r16li.genblk1[4].latchcgate_inst.Q ),
    .X(_0429_));
 sg13g2_nor2_1 _1021_ (.A(net147),
    .B(_0429_),
    .Y(_0027_));
 sg13g2_nand2_1 _1022_ (.Y(_0430_),
    .A(net175),
    .B(\r16li.genblk1[1].latchcgate_inst.Q ));
 sg13g2_inv_1 _1023_ (.Y(_0024_),
    .A(_0430_));
 sg13g2_xor2_1 _1024_ (.B(\r16li.genblk1[1].latchcgate_inst.Q ),
    .A(\r16li.genblk1[3].latchcgate_inst.Q ),
    .X(_0431_));
 sg13g2_nor2_1 _1025_ (.A(net147),
    .B(_0431_),
    .Y(_0025_));
 sg13g2_and2_1 _1026_ (.A(net175),
    .B(R16l),
    .X(_0022_));
 sg13g2_xor2_1 _1027_ (.B(\r16li.genblk1[2].latchcgate_inst.Q ),
    .A(R16l),
    .X(_0432_));
 sg13g2_nor2_1 _1028_ (.A(net148),
    .B(_0432_),
    .Y(_0023_));
 sg13g2_a22oi_1 _1029_ (.Y(_0009_),
    .B1(_0008_),
    .B2(_0430_),
    .A2(\r16li.genblk1[1].latchcgate_inst.Q ),
    .A1(_0177_));
 sg13g2_dllrq_1 _1030_ (.D(_0164_),
    .GATE_N(_0165_),
    .RESET_B(net19),
    .Q(\rtbdli.genblk1[0].latchcgate_inst.A ));
 sg13g2_dllrq_1 _1031_ (.D(_0162_),
    .GATE_N(_0163_),
    .RESET_B(net20),
    .Q(\rtbdli.genblk1[62].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1032_ (.D(_0160_),
    .GATE_N(_0161_),
    .RESET_B(net21),
    .Q(\rtbdli.genblk1[61].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1033_ (.D(_0158_),
    .GATE_N(_0159_),
    .RESET_B(net22),
    .Q(\rtbdli.genblk1[60].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1034_ (.D(_0154_),
    .GATE_N(_0155_),
    .RESET_B(net23),
    .Q(\rtbdli.genblk1[59].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1035_ (.D(_0152_),
    .GATE_N(_0153_),
    .RESET_B(net24),
    .Q(\rtbdli.genblk1[58].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1036_ (.D(_0150_),
    .GATE_N(_0151_),
    .RESET_B(net25),
    .Q(\rtbdli.genblk1[57].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1037_ (.D(_0148_),
    .GATE_N(_0149_),
    .RESET_B(net26),
    .Q(\rtbdli.genblk1[56].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1038_ (.D(_0146_),
    .GATE_N(_0147_),
    .RESET_B(net27),
    .Q(\rtbdli.genblk1[55].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1039_ (.D(_0144_),
    .GATE_N(_0145_),
    .RESET_B(net28),
    .Q(\rtbdli.genblk1[54].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1040_ (.D(_0142_),
    .GATE_N(_0143_),
    .RESET_B(net29),
    .Q(\rtbdli.genblk1[53].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1041_ (.D(_0140_),
    .GATE_N(_0141_),
    .RESET_B(net30),
    .Q(\rtbdli.genblk1[52].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1042_ (.D(_0138_),
    .GATE_N(_0139_),
    .RESET_B(net31),
    .Q(\rtbdli.genblk1[51].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1043_ (.D(_0136_),
    .GATE_N(_0137_),
    .RESET_B(net32),
    .Q(\rtbdli.genblk1[50].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1044_ (.D(_0132_),
    .GATE_N(_0133_),
    .RESET_B(net33),
    .Q(\rtbdli.genblk1[49].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1045_ (.D(_0130_),
    .GATE_N(_0131_),
    .RESET_B(net34),
    .Q(\rtbdli.genblk1[48].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1046_ (.D(_0128_),
    .GATE_N(_0129_),
    .RESET_B(net35),
    .Q(\rtbdli.genblk1[47].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1047_ (.D(_0126_),
    .GATE_N(_0127_),
    .RESET_B(net36),
    .Q(\rtbdli.genblk1[46].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1048_ (.D(_0124_),
    .GATE_N(_0125_),
    .RESET_B(net37),
    .Q(\rtbdli.genblk1[45].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1049_ (.D(_0122_),
    .GATE_N(_0123_),
    .RESET_B(net38),
    .Q(\rtbdli.genblk1[44].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1050_ (.D(_0120_),
    .GATE_N(_0121_),
    .RESET_B(net39),
    .Q(\rtbdli.genblk1[43].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1051_ (.D(_0118_),
    .GATE_N(_0119_),
    .RESET_B(net40),
    .Q(\rtbdli.genblk1[42].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1052_ (.D(_0116_),
    .GATE_N(_0117_),
    .RESET_B(net41),
    .Q(\rtbdli.genblk1[41].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1053_ (.D(_0114_),
    .GATE_N(_0115_),
    .RESET_B(net42),
    .Q(\rtbdli.genblk1[40].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1054_ (.D(_0110_),
    .GATE_N(_0111_),
    .RESET_B(net43),
    .Q(\rtbdli.genblk1[39].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1055_ (.D(_0108_),
    .GATE_N(_0109_),
    .RESET_B(net44),
    .Q(\rtbdli.genblk1[38].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1056_ (.D(_0106_),
    .GATE_N(_0107_),
    .RESET_B(net45),
    .Q(\rtbdli.genblk1[37].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1057_ (.D(_0104_),
    .GATE_N(_0105_),
    .RESET_B(net46),
    .Q(\rtbdli.genblk1[36].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1058_ (.D(_0102_),
    .GATE_N(_0103_),
    .RESET_B(net47),
    .Q(\rtbdli.genblk1[35].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1059_ (.D(_0100_),
    .GATE_N(_0101_),
    .RESET_B(net48),
    .Q(\rtbdli.genblk1[34].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1060_ (.D(_0098_),
    .GATE_N(_0099_),
    .RESET_B(net49),
    .Q(\rtbdli.genblk1[33].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1061_ (.D(_0096_),
    .GATE_N(_0097_),
    .RESET_B(net50),
    .Q(\rtbdli.genblk1[32].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1062_ (.D(_0094_),
    .GATE_N(_0095_),
    .RESET_B(net51),
    .Q(\rtbdli.genblk1[31].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1063_ (.D(_0092_),
    .GATE_N(_0093_),
    .RESET_B(net52),
    .Q(\rtbdli.genblk1[30].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1064_ (.D(_0088_),
    .GATE_N(_0089_),
    .RESET_B(net53),
    .Q(\rtbdli.genblk1[29].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1065_ (.D(_0086_),
    .GATE_N(_0087_),
    .RESET_B(net54),
    .Q(\rtbdli.genblk1[28].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1066_ (.D(_0084_),
    .GATE_N(_0085_),
    .RESET_B(net55),
    .Q(\rtbdli.genblk1[27].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1067_ (.D(_0082_),
    .GATE_N(_0083_),
    .RESET_B(net56),
    .Q(\rtbdli.genblk1[26].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1068_ (.D(_0080_),
    .GATE_N(_0081_),
    .RESET_B(net57),
    .Q(\rtbdli.genblk1[25].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1069_ (.D(_0078_),
    .GATE_N(_0079_),
    .RESET_B(net58),
    .Q(\rtbdli.genblk1[24].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1070_ (.D(_0076_),
    .GATE_N(_0077_),
    .RESET_B(net59),
    .Q(\rtbdli.genblk1[23].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1071_ (.D(_0074_),
    .GATE_N(_0075_),
    .RESET_B(net60),
    .Q(\rtbdli.genblk1[22].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1072_ (.D(_0072_),
    .GATE_N(_0073_),
    .RESET_B(net61),
    .Q(\rtbdli.genblk1[21].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1073_ (.D(_0070_),
    .GATE_N(_0071_),
    .RESET_B(net62),
    .Q(\rtbdli.genblk1[20].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1074_ (.D(_0066_),
    .GATE_N(_0067_),
    .RESET_B(net63),
    .Q(\rtbdli.genblk1[19].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1075_ (.D(_0064_),
    .GATE_N(_0065_),
    .RESET_B(net64),
    .Q(\rtbdli.genblk1[18].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1076_ (.D(_0062_),
    .GATE_N(_0063_),
    .RESET_B(net65),
    .Q(\rtbdli.genblk1[17].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1077_ (.D(_0060_),
    .GATE_N(_0061_),
    .RESET_B(net66),
    .Q(\rtbdli.genblk1[16].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1078_ (.D(_0058_),
    .GATE_N(_0059_),
    .RESET_B(net67),
    .Q(\rtbdli.genblk1[15].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1079_ (.D(_0056_),
    .GATE_N(_0057_),
    .RESET_B(net68),
    .Q(\rtbdli.genblk1[14].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1080_ (.D(_0054_),
    .GATE_N(_0055_),
    .RESET_B(net69),
    .Q(\rtbdli.genblk1[13].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1081_ (.D(_0052_),
    .GATE_N(_0053_),
    .RESET_B(net70),
    .Q(\rtbdli.genblk1[12].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1082_ (.D(_0050_),
    .GATE_N(_0051_),
    .RESET_B(net71),
    .Q(\rtbdli.genblk1[11].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1083_ (.D(_0048_),
    .GATE_N(_0049_),
    .RESET_B(net72),
    .Q(\rtbdli.genblk1[10].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1084_ (.D(_0172_),
    .GATE_N(_0173_),
    .RESET_B(net73),
    .Q(\rtbdli.genblk1[10].latchcgate_inst.A ));
 sg13g2_dllrq_1 _1085_ (.D(_0170_),
    .GATE_N(_0171_),
    .RESET_B(net74),
    .Q(\rtbdli.genblk1[8].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1086_ (.D(_0168_),
    .GATE_N(_0169_),
    .RESET_B(net75),
    .Q(\rtbdli.genblk1[7].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1087_ (.D(_0166_),
    .GATE_N(_0167_),
    .RESET_B(net76),
    .Q(\rtbdli.genblk1[6].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1088_ (.D(_0156_),
    .GATE_N(_0157_),
    .RESET_B(net77),
    .Q(\rtbdli.genblk1[5].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1089_ (.D(_0134_),
    .GATE_N(_0135_),
    .RESET_B(net78),
    .Q(\rtbdli.genblk1[4].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1090_ (.D(_0112_),
    .GATE_N(_0113_),
    .RESET_B(net79),
    .Q(\rtbdli.genblk1[3].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1091_ (.D(_0090_),
    .GATE_N(_0091_),
    .RESET_B(net80),
    .Q(\rtbdli.genblk1[2].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1092_ (.D(_0068_),
    .GATE_N(_0069_),
    .RESET_B(net81),
    .Q(\rtbdli.genblk1[1].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1093_ (.D(_0046_),
    .GATE_N(_0047_),
    .RESET_B(net82),
    .Q(RBigl));
 sg13g2_dfrbp_1 _1094_ (.CLK(RBigc),
    .RESET_B(net163),
    .D(_0004_),
    .Q_N(_0004_),
    .Q(RBigct));
 sg13g2_dfrbp_1 _1095_ (.CLK(RBigl),
    .RESET_B(net167),
    .D(_0005_),
    .Q_N(_0005_),
    .Q(RBiglt));
 sg13g2_dfrbp_1 _1096_ (.CLK(R16c),
    .RESET_B(net165),
    .D(_0000_),
    .Q_N(_0000_),
    .Q(R16ct));
 sg13g2_dfrbp_1 _1097_ (.CLK(R16l),
    .RESET_B(net174),
    .D(_0001_),
    .Q_N(_0001_),
    .Q(R16lt));
 sg13g2_dfrbp_1 _1098_ (.CLK(R4c),
    .RESET_B(net165),
    .D(_0002_),
    .Q_N(_0002_),
    .Q(R4ct));
 sg13g2_dfrbp_1 _1099_ (.CLK(R4l),
    .RESET_B(net174),
    .D(_0003_),
    .Q_N(_0003_),
    .Q(R4lt));
 sg13g2_dllrq_1 _1100_ (.D(_0006_),
    .GATE_N(_0007_),
    .RESET_B(net83),
    .Q(Ql));
 sg13g2_dllrq_1 _1101_ (.D(_0045_),
    .GATE_N(_0043_),
    .RESET_B(net84),
    .Q(\r4li.genblk1[0].latchcgate_inst.A ));
 sg13g2_dllrq_1 _1102_ (.D(_0044_),
    .GATE_N(_0041_),
    .RESET_B(net85),
    .Q(\r4li.genblk1[2].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1103_ (.D(_0042_),
    .GATE_N(_0043_),
    .RESET_B(net86),
    .Q(\r4li.genblk1[1].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1104_ (.D(_0040_),
    .GATE_N(_0041_),
    .RESET_B(net87),
    .Q(R4l));
 sg13g2_dllrq_1 _1105_ (.D(_0020_),
    .GATE_N(_0021_),
    .RESET_B(net88),
    .Q(\r16li.genblk1[0].latchcgate_inst.A ));
 sg13g2_dllrq_1 _1106_ (.D(_0018_),
    .GATE_N(_0019_),
    .RESET_B(net89),
    .Q(\r16li.genblk1[14].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1107_ (.D(_0016_),
    .GATE_N(_0017_),
    .RESET_B(net90),
    .Q(\r16li.genblk1[13].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1108_ (.D(_0014_),
    .GATE_N(_0015_),
    .RESET_B(net91),
    .Q(\r16li.genblk1[12].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1109_ (.D(_0012_),
    .GATE_N(_0013_),
    .RESET_B(net92),
    .Q(\r16li.genblk1[11].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1110_ (.D(_0010_),
    .GATE_N(_0011_),
    .RESET_B(net93),
    .Q(\r16li.genblk1[10].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1111_ (.D(_0038_),
    .GATE_N(_0039_),
    .RESET_B(net94),
    .Q(\r16li.genblk1[10].latchcgate_inst.A ));
 sg13g2_dllrq_1 _1112_ (.D(_0036_),
    .GATE_N(_0037_),
    .RESET_B(net95),
    .Q(\r16li.genblk1[8].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1113_ (.D(_0034_),
    .GATE_N(_0035_),
    .RESET_B(net96),
    .Q(\r16li.genblk1[7].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1114_ (.D(_0032_),
    .GATE_N(_0033_),
    .RESET_B(net97),
    .Q(\r16li.genblk1[6].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1115_ (.D(_0030_),
    .GATE_N(_0031_),
    .RESET_B(net98),
    .Q(\r16li.genblk1[5].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1116_ (.D(_0028_),
    .GATE_N(_0029_),
    .RESET_B(net99),
    .Q(\r16li.genblk1[4].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1117_ (.D(_0026_),
    .GATE_N(_0027_),
    .RESET_B(net100),
    .Q(\r16li.genblk1[3].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1118_ (.D(_0024_),
    .GATE_N(_0025_),
    .RESET_B(net101),
    .Q(\r16li.genblk1[2].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1119_ (.D(_0022_),
    .GATE_N(_0023_),
    .RESET_B(net102),
    .Q(\r16li.genblk1[1].latchcgate_inst.Q ));
 sg13g2_dllrq_1 _1120_ (.D(_0008_),
    .GATE_N(_0009_),
    .RESET_B(net103),
    .Q(R16l));
 sg13g2_tiehi _1031__20 (.L_HI(net20));
 sg13g2_tiehi _1032__21 (.L_HI(net21));
 sg13g2_tiehi _1033__22 (.L_HI(net22));
 sg13g2_tiehi _1034__23 (.L_HI(net23));
 sg13g2_tiehi _1035__24 (.L_HI(net24));
 sg13g2_tiehi _1036__25 (.L_HI(net25));
 sg13g2_tiehi _1037__26 (.L_HI(net26));
 sg13g2_tiehi _1038__27 (.L_HI(net27));
 sg13g2_tiehi _1039__28 (.L_HI(net28));
 sg13g2_tiehi _1040__29 (.L_HI(net29));
 sg13g2_tiehi _1041__30 (.L_HI(net30));
 sg13g2_tiehi _1042__31 (.L_HI(net31));
 sg13g2_tiehi _1043__32 (.L_HI(net32));
 sg13g2_tiehi _1044__33 (.L_HI(net33));
 sg13g2_tiehi _1045__34 (.L_HI(net34));
 sg13g2_tiehi _1046__35 (.L_HI(net35));
 sg13g2_tiehi _1047__36 (.L_HI(net36));
 sg13g2_tiehi _1048__37 (.L_HI(net37));
 sg13g2_tiehi _1049__38 (.L_HI(net38));
 sg13g2_tiehi _1050__39 (.L_HI(net39));
 sg13g2_tiehi _1051__40 (.L_HI(net40));
 sg13g2_tiehi _1052__41 (.L_HI(net41));
 sg13g2_tiehi _1053__42 (.L_HI(net42));
 sg13g2_tiehi _1054__43 (.L_HI(net43));
 sg13g2_tiehi _1055__44 (.L_HI(net44));
 sg13g2_tiehi _1056__45 (.L_HI(net45));
 sg13g2_tiehi _1057__46 (.L_HI(net46));
 sg13g2_tiehi _1058__47 (.L_HI(net47));
 sg13g2_tiehi _1059__48 (.L_HI(net48));
 sg13g2_tiehi _1060__49 (.L_HI(net49));
 sg13g2_tiehi _1061__50 (.L_HI(net50));
 sg13g2_tiehi _1062__51 (.L_HI(net51));
 sg13g2_tiehi _1063__52 (.L_HI(net52));
 sg13g2_tiehi _1064__53 (.L_HI(net53));
 sg13g2_tiehi _1065__54 (.L_HI(net54));
 sg13g2_tiehi _1066__55 (.L_HI(net55));
 sg13g2_tiehi _1067__56 (.L_HI(net56));
 sg13g2_tiehi _1068__57 (.L_HI(net57));
 sg13g2_tiehi _1069__58 (.L_HI(net58));
 sg13g2_tiehi _1070__59 (.L_HI(net59));
 sg13g2_tiehi _1071__60 (.L_HI(net60));
 sg13g2_tiehi _1072__61 (.L_HI(net61));
 sg13g2_tiehi _1073__62 (.L_HI(net62));
 sg13g2_tiehi _1074__63 (.L_HI(net63));
 sg13g2_tiehi _1075__64 (.L_HI(net64));
 sg13g2_tiehi _1076__65 (.L_HI(net65));
 sg13g2_tiehi _1077__66 (.L_HI(net66));
 sg13g2_tiehi _1078__67 (.L_HI(net67));
 sg13g2_tiehi _1079__68 (.L_HI(net68));
 sg13g2_tiehi _1080__69 (.L_HI(net69));
 sg13g2_tiehi _1081__70 (.L_HI(net70));
 sg13g2_tiehi _1082__71 (.L_HI(net71));
 sg13g2_tiehi _1083__72 (.L_HI(net72));
 sg13g2_tiehi _1084__73 (.L_HI(net73));
 sg13g2_tiehi _1085__74 (.L_HI(net74));
 sg13g2_tiehi _1086__75 (.L_HI(net75));
 sg13g2_tiehi _1087__76 (.L_HI(net76));
 sg13g2_tiehi _1088__77 (.L_HI(net77));
 sg13g2_tiehi _1089__78 (.L_HI(net78));
 sg13g2_tiehi _1090__79 (.L_HI(net79));
 sg13g2_tiehi _1091__80 (.L_HI(net80));
 sg13g2_tiehi _1092__81 (.L_HI(net81));
 sg13g2_tiehi _1093__82 (.L_HI(net82));
 sg13g2_tiehi _1100__83 (.L_HI(net83));
 sg13g2_tiehi _1101__84 (.L_HI(net84));
 sg13g2_tiehi _1102__85 (.L_HI(net85));
 sg13g2_tiehi _1103__86 (.L_HI(net86));
 sg13g2_tiehi _1104__87 (.L_HI(net87));
 sg13g2_tiehi _1105__88 (.L_HI(net88));
 sg13g2_tiehi _1106__89 (.L_HI(net89));
 sg13g2_tiehi _1107__90 (.L_HI(net90));
 sg13g2_tiehi _1108__91 (.L_HI(net91));
 sg13g2_tiehi _1109__92 (.L_HI(net92));
 sg13g2_tiehi _1110__93 (.L_HI(net93));
 sg13g2_tiehi _1111__94 (.L_HI(net94));
 sg13g2_tiehi _1112__95 (.L_HI(net95));
 sg13g2_tiehi _1113__96 (.L_HI(net96));
 sg13g2_tiehi _1114__97 (.L_HI(net97));
 sg13g2_tiehi _1115__98 (.L_HI(net98));
 sg13g2_tiehi _1116__99 (.L_HI(net99));
 sg13g2_tiehi _1117__100 (.L_HI(net100));
 sg13g2_tiehi _1118__101 (.L_HI(net101));
 sg13g2_tiehi _1119__102 (.L_HI(net102));
 sg13g2_tiehi _1120__103 (.L_HI(net103));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_tielo tt_um_tommythorn_cgates_4 (.L_LO(net4));
 sg13g2_tielo tt_um_tommythorn_cgates_5 (.L_LO(net5));
 sg13g2_tielo tt_um_tommythorn_cgates_6 (.L_LO(net6));
 sg13g2_tielo tt_um_tommythorn_cgates_7 (.L_LO(net7));
 sg13g2_tielo tt_um_tommythorn_cgates_8 (.L_LO(net8));
 sg13g2_tielo tt_um_tommythorn_cgates_9 (.L_LO(net9));
 sg13g2_tielo tt_um_tommythorn_cgates_10 (.L_LO(net10));
 sg13g2_tielo tt_um_tommythorn_cgates_11 (.L_LO(net11));
 sg13g2_tielo tt_um_tommythorn_cgates_12 (.L_LO(net12));
 sg13g2_tielo tt_um_tommythorn_cgates_13 (.L_LO(net13));
 sg13g2_tielo tt_um_tommythorn_cgates_14 (.L_LO(net14));
 sg13g2_tielo tt_um_tommythorn_cgates_15 (.L_LO(net15));
 sg13g2_tielo tt_um_tommythorn_cgates_16 (.L_LO(net16));
 sg13g2_tielo tt_um_tommythorn_cgates_17 (.L_LO(net17));
 sg13g2_tielo tt_um_tommythorn_cgates_18 (.L_LO(net18));
 sg13g2_tiehi _1030__19 (.L_HI(net19));
 sg13g2_buf_1 _1222_ (.A(Ql),
    .X(uo_out[0]));
 sg13g2_buf_1 _1223_ (.A(Qc),
    .X(uo_out[1]));
 sg13g2_buf_1 _1224_ (.A(R4lt),
    .X(uo_out[2]));
 sg13g2_buf_1 _1225_ (.A(R4ct),
    .X(uo_out[3]));
 sg13g2_buf_1 _1226_ (.A(R16lt),
    .X(uo_out[4]));
 sg13g2_buf_1 _1227_ (.A(R16ct),
    .X(uo_out[5]));
 sg13g2_buf_1 _1228_ (.A(RBiglt),
    .X(uo_out[6]));
 sg13g2_buf_1 _1229_ (.A(RBigct),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout136 (.A(net137),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(net139),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(net139),
    .X(net138));
 sg13g2_buf_1 fanout139 (.A(net149),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(net149),
    .X(net140));
 sg13g2_buf_1 fanout141 (.A(net149),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(net145),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(net145),
    .X(net143));
 sg13g2_buf_1 fanout144 (.A(net145),
    .X(net144));
 sg13g2_buf_1 fanout145 (.A(net149),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(net148),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(net149),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_0174_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(net152),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(net152),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(net158),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(net155),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(net155),
    .X(net154));
 sg13g2_buf_1 fanout155 (.A(net158),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(net157),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(net158),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(rst_n),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(net160),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(net164),
    .X(net160));
 sg13g2_buf_1 fanout161 (.A(net164),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(net163),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(net164),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(net167),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(net167),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(net167),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(rst_n),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(net178),
    .X(net168));
 sg13g2_buf_1 fanout169 (.A(net178),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(net172),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(net172),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(net178),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(net177),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(net177),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(net176),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(net177),
    .X(net176));
 sg13g2_buf_1 fanout177 (.A(net178),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(rst_n),
    .X(net178));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_tielo tt_um_tommythorn_cgates_3 (.L_LO(net3));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_fill_1 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_117 ();
 sg13g2_decap_8 FILLER_16_124 ();
 sg13g2_decap_8 FILLER_16_131 ();
 sg13g2_decap_8 FILLER_16_138 ();
 sg13g2_decap_4 FILLER_16_145 ();
 sg13g2_fill_2 FILLER_16_149 ();
 sg13g2_decap_8 FILLER_16_167 ();
 sg13g2_fill_2 FILLER_16_174 ();
 sg13g2_decap_8 FILLER_16_181 ();
 sg13g2_fill_2 FILLER_16_188 ();
 sg13g2_decap_4 FILLER_16_194 ();
 sg13g2_fill_2 FILLER_16_198 ();
 sg13g2_fill_2 FILLER_16_216 ();
 sg13g2_decap_8 FILLER_16_227 ();
 sg13g2_decap_8 FILLER_16_234 ();
 sg13g2_decap_8 FILLER_16_241 ();
 sg13g2_decap_8 FILLER_16_248 ();
 sg13g2_decap_8 FILLER_16_255 ();
 sg13g2_decap_8 FILLER_16_262 ();
 sg13g2_decap_8 FILLER_16_269 ();
 sg13g2_decap_8 FILLER_16_276 ();
 sg13g2_decap_8 FILLER_16_283 ();
 sg13g2_decap_8 FILLER_16_290 ();
 sg13g2_decap_8 FILLER_16_297 ();
 sg13g2_decap_8 FILLER_16_304 ();
 sg13g2_decap_8 FILLER_16_311 ();
 sg13g2_decap_8 FILLER_16_318 ();
 sg13g2_decap_8 FILLER_16_325 ();
 sg13g2_decap_8 FILLER_16_332 ();
 sg13g2_decap_8 FILLER_16_339 ();
 sg13g2_decap_8 FILLER_16_346 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_367 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_fill_2 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_123 ();
 sg13g2_decap_8 FILLER_17_130 ();
 sg13g2_decap_8 FILLER_17_137 ();
 sg13g2_fill_2 FILLER_17_144 ();
 sg13g2_fill_1 FILLER_17_163 ();
 sg13g2_fill_1 FILLER_17_168 ();
 sg13g2_fill_2 FILLER_17_193 ();
 sg13g2_fill_1 FILLER_17_208 ();
 sg13g2_decap_8 FILLER_17_241 ();
 sg13g2_decap_8 FILLER_17_248 ();
 sg13g2_decap_8 FILLER_17_255 ();
 sg13g2_decap_8 FILLER_17_262 ();
 sg13g2_decap_8 FILLER_17_269 ();
 sg13g2_decap_8 FILLER_17_276 ();
 sg13g2_decap_8 FILLER_17_283 ();
 sg13g2_decap_8 FILLER_17_290 ();
 sg13g2_decap_8 FILLER_17_297 ();
 sg13g2_decap_8 FILLER_17_304 ();
 sg13g2_decap_8 FILLER_17_311 ();
 sg13g2_decap_8 FILLER_17_318 ();
 sg13g2_decap_8 FILLER_17_325 ();
 sg13g2_decap_8 FILLER_17_332 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_367 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_fill_2 FILLER_18_84 ();
 sg13g2_decap_4 FILLER_18_111 ();
 sg13g2_fill_2 FILLER_18_115 ();
 sg13g2_fill_2 FILLER_18_134 ();
 sg13g2_fill_1 FILLER_18_136 ();
 sg13g2_fill_2 FILLER_18_162 ();
 sg13g2_decap_8 FILLER_18_180 ();
 sg13g2_decap_8 FILLER_18_187 ();
 sg13g2_decap_4 FILLER_18_194 ();
 sg13g2_fill_1 FILLER_18_198 ();
 sg13g2_fill_1 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_212 ();
 sg13g2_decap_4 FILLER_18_219 ();
 sg13g2_decap_8 FILLER_18_235 ();
 sg13g2_fill_2 FILLER_18_242 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_4 FILLER_18_259 ();
 sg13g2_fill_2 FILLER_18_263 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_4 FILLER_18_294 ();
 sg13g2_fill_2 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_fill_2 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_344 ();
 sg13g2_decap_4 FILLER_18_351 ();
 sg13g2_fill_1 FILLER_18_355 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_4 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_102 ();
 sg13g2_decap_8 FILLER_19_109 ();
 sg13g2_fill_2 FILLER_19_116 ();
 sg13g2_decap_8 FILLER_19_135 ();
 sg13g2_decap_4 FILLER_19_142 ();
 sg13g2_fill_2 FILLER_19_146 ();
 sg13g2_fill_1 FILLER_19_165 ();
 sg13g2_decap_8 FILLER_19_187 ();
 sg13g2_fill_2 FILLER_19_225 ();
 sg13g2_fill_1 FILLER_19_227 ();
 sg13g2_decap_8 FILLER_19_286 ();
 sg13g2_decap_4 FILLER_19_293 ();
 sg13g2_fill_1 FILLER_19_334 ();
 sg13g2_fill_1 FILLER_19_356 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_4 FILLER_20_77 ();
 sg13g2_fill_2 FILLER_20_81 ();
 sg13g2_fill_1 FILLER_20_112 ();
 sg13g2_fill_1 FILLER_20_135 ();
 sg13g2_fill_1 FILLER_20_141 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_fill_1 FILLER_20_207 ();
 sg13g2_decap_8 FILLER_20_212 ();
 sg13g2_decap_4 FILLER_20_219 ();
 sg13g2_fill_1 FILLER_20_223 ();
 sg13g2_decap_4 FILLER_20_233 ();
 sg13g2_decap_8 FILLER_20_253 ();
 sg13g2_fill_2 FILLER_20_260 ();
 sg13g2_decap_4 FILLER_20_266 ();
 sg13g2_fill_2 FILLER_20_274 ();
 sg13g2_fill_2 FILLER_20_281 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_4 FILLER_20_294 ();
 sg13g2_decap_4 FILLER_20_314 ();
 sg13g2_fill_1 FILLER_20_318 ();
 sg13g2_decap_8 FILLER_20_323 ();
 sg13g2_fill_2 FILLER_20_330 ();
 sg13g2_decap_4 FILLER_20_336 ();
 sg13g2_fill_2 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_346 ();
 sg13g2_decap_8 FILLER_20_366 ();
 sg13g2_fill_1 FILLER_20_373 ();
 sg13g2_fill_2 FILLER_20_378 ();
 sg13g2_fill_1 FILLER_20_380 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_fill_1 FILLER_21_84 ();
 sg13g2_decap_4 FILLER_21_102 ();
 sg13g2_fill_2 FILLER_21_106 ();
 sg13g2_decap_8 FILLER_21_157 ();
 sg13g2_fill_1 FILLER_21_164 ();
 sg13g2_decap_8 FILLER_21_178 ();
 sg13g2_fill_1 FILLER_21_185 ();
 sg13g2_fill_2 FILLER_21_200 ();
 sg13g2_decap_4 FILLER_21_227 ();
 sg13g2_fill_1 FILLER_21_231 ();
 sg13g2_fill_2 FILLER_21_253 ();
 sg13g2_fill_1 FILLER_21_255 ();
 sg13g2_decap_4 FILLER_21_264 ();
 sg13g2_fill_2 FILLER_21_268 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_4 FILLER_21_301 ();
 sg13g2_decap_4 FILLER_21_318 ();
 sg13g2_fill_1 FILLER_21_335 ();
 sg13g2_decap_8 FILLER_21_341 ();
 sg13g2_fill_1 FILLER_21_348 ();
 sg13g2_fill_2 FILLER_21_362 ();
 sg13g2_decap_4 FILLER_21_380 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_4 FILLER_21_399 ();
 sg13g2_fill_1 FILLER_21_403 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_4 FILLER_22_77 ();
 sg13g2_fill_1 FILLER_22_81 ();
 sg13g2_decap_4 FILLER_22_99 ();
 sg13g2_decap_4 FILLER_22_107 ();
 sg13g2_fill_1 FILLER_22_111 ();
 sg13g2_fill_2 FILLER_22_117 ();
 sg13g2_fill_1 FILLER_22_119 ();
 sg13g2_decap_4 FILLER_22_129 ();
 sg13g2_fill_2 FILLER_22_133 ();
 sg13g2_decap_4 FILLER_22_157 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_178 ();
 sg13g2_fill_1 FILLER_22_187 ();
 sg13g2_fill_2 FILLER_22_220 ();
 sg13g2_decap_4 FILLER_22_234 ();
 sg13g2_fill_1 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_243 ();
 sg13g2_fill_1 FILLER_22_275 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_fill_1 FILLER_22_291 ();
 sg13g2_fill_2 FILLER_22_296 ();
 sg13g2_fill_2 FILLER_22_322 ();
 sg13g2_fill_1 FILLER_22_324 ();
 sg13g2_decap_4 FILLER_22_345 ();
 sg13g2_decap_8 FILLER_22_366 ();
 sg13g2_fill_1 FILLER_22_373 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_4 FILLER_23_77 ();
 sg13g2_fill_2 FILLER_23_81 ();
 sg13g2_fill_1 FILLER_23_100 ();
 sg13g2_decap_4 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_128 ();
 sg13g2_decap_4 FILLER_23_135 ();
 sg13g2_fill_2 FILLER_23_139 ();
 sg13g2_decap_8 FILLER_23_153 ();
 sg13g2_decap_8 FILLER_23_160 ();
 sg13g2_decap_8 FILLER_23_167 ();
 sg13g2_fill_2 FILLER_23_183 ();
 sg13g2_decap_4 FILLER_23_197 ();
 sg13g2_fill_1 FILLER_23_201 ();
 sg13g2_decap_4 FILLER_23_206 ();
 sg13g2_decap_8 FILLER_23_215 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_fill_1 FILLER_23_249 ();
 sg13g2_decap_4 FILLER_23_255 ();
 sg13g2_fill_1 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_264 ();
 sg13g2_fill_1 FILLER_23_271 ();
 sg13g2_fill_2 FILLER_23_296 ();
 sg13g2_fill_1 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_304 ();
 sg13g2_decap_4 FILLER_23_311 ();
 sg13g2_fill_1 FILLER_23_319 ();
 sg13g2_decap_4 FILLER_23_334 ();
 sg13g2_fill_2 FILLER_23_338 ();
 sg13g2_decap_4 FILLER_23_344 ();
 sg13g2_fill_2 FILLER_23_352 ();
 sg13g2_fill_1 FILLER_23_354 ();
 sg13g2_decap_4 FILLER_23_375 ();
 sg13g2_fill_1 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_105 ();
 sg13g2_decap_4 FILLER_24_127 ();
 sg13g2_fill_1 FILLER_24_131 ();
 sg13g2_decap_4 FILLER_24_161 ();
 sg13g2_fill_1 FILLER_24_165 ();
 sg13g2_decap_4 FILLER_24_190 ();
 sg13g2_decap_8 FILLER_24_199 ();
 sg13g2_decap_4 FILLER_24_206 ();
 sg13g2_decap_4 FILLER_24_223 ();
 sg13g2_fill_2 FILLER_24_227 ();
 sg13g2_decap_4 FILLER_24_234 ();
 sg13g2_fill_1 FILLER_24_238 ();
 sg13g2_fill_1 FILLER_24_243 ();
 sg13g2_decap_4 FILLER_24_272 ();
 sg13g2_fill_2 FILLER_24_276 ();
 sg13g2_fill_2 FILLER_24_287 ();
 sg13g2_fill_1 FILLER_24_289 ();
 sg13g2_fill_2 FILLER_24_352 ();
 sg13g2_decap_4 FILLER_24_378 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_4 FILLER_25_91 ();
 sg13g2_fill_2 FILLER_25_95 ();
 sg13g2_decap_4 FILLER_25_135 ();
 sg13g2_fill_1 FILLER_25_139 ();
 sg13g2_fill_2 FILLER_25_145 ();
 sg13g2_fill_1 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_165 ();
 sg13g2_decap_4 FILLER_25_172 ();
 sg13g2_fill_1 FILLER_25_176 ();
 sg13g2_decap_4 FILLER_25_181 ();
 sg13g2_fill_2 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_215 ();
 sg13g2_fill_2 FILLER_25_232 ();
 sg13g2_fill_2 FILLER_25_239 ();
 sg13g2_fill_1 FILLER_25_250 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_290 ();
 sg13g2_fill_1 FILLER_25_297 ();
 sg13g2_decap_8 FILLER_25_306 ();
 sg13g2_fill_2 FILLER_25_313 ();
 sg13g2_decap_8 FILLER_25_332 ();
 sg13g2_fill_2 FILLER_25_339 ();
 sg13g2_fill_1 FILLER_25_341 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_fill_1 FILLER_25_357 ();
 sg13g2_decap_4 FILLER_25_371 ();
 sg13g2_fill_2 FILLER_25_379 ();
 sg13g2_fill_1 FILLER_25_381 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_fill_2 FILLER_26_112 ();
 sg13g2_fill_1 FILLER_26_114 ();
 sg13g2_fill_2 FILLER_26_136 ();
 sg13g2_decap_8 FILLER_26_164 ();
 sg13g2_decap_4 FILLER_26_171 ();
 sg13g2_fill_2 FILLER_26_175 ();
 sg13g2_fill_2 FILLER_26_190 ();
 sg13g2_fill_1 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_201 ();
 sg13g2_decap_8 FILLER_26_208 ();
 sg13g2_fill_1 FILLER_26_228 ();
 sg13g2_fill_1 FILLER_26_233 ();
 sg13g2_fill_1 FILLER_26_276 ();
 sg13g2_fill_1 FILLER_26_290 ();
 sg13g2_fill_1 FILLER_26_315 ();
 sg13g2_fill_2 FILLER_26_332 ();
 sg13g2_fill_1 FILLER_26_334 ();
 sg13g2_fill_1 FILLER_26_356 ();
 sg13g2_decap_4 FILLER_26_381 ();
 sg13g2_fill_1 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_395 ();
 sg13g2_fill_2 FILLER_26_402 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_fill_2 FILLER_27_84 ();
 sg13g2_fill_1 FILLER_27_86 ();
 sg13g2_fill_2 FILLER_27_113 ();
 sg13g2_fill_1 FILLER_27_115 ();
 sg13g2_fill_2 FILLER_27_120 ();
 sg13g2_fill_1 FILLER_27_122 ();
 sg13g2_decap_8 FILLER_27_135 ();
 sg13g2_fill_1 FILLER_27_180 ();
 sg13g2_fill_2 FILLER_27_205 ();
 sg13g2_fill_1 FILLER_27_223 ();
 sg13g2_fill_1 FILLER_27_236 ();
 sg13g2_fill_2 FILLER_27_253 ();
 sg13g2_fill_1 FILLER_27_267 ();
 sg13g2_decap_8 FILLER_27_293 ();
 sg13g2_decap_4 FILLER_27_300 ();
 sg13g2_fill_1 FILLER_27_304 ();
 sg13g2_decap_8 FILLER_27_309 ();
 sg13g2_fill_2 FILLER_27_316 ();
 sg13g2_fill_1 FILLER_27_318 ();
 sg13g2_decap_8 FILLER_27_335 ();
 sg13g2_fill_2 FILLER_27_342 ();
 sg13g2_decap_4 FILLER_27_348 ();
 sg13g2_fill_1 FILLER_27_352 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_369 ();
 sg13g2_fill_2 FILLER_27_376 ();
 sg13g2_fill_1 FILLER_27_378 ();
 sg13g2_fill_2 FILLER_27_383 ();
 sg13g2_decap_8 FILLER_27_397 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_4 FILLER_28_74 ();
 sg13g2_fill_1 FILLER_28_78 ();
 sg13g2_fill_2 FILLER_28_88 ();
 sg13g2_fill_2 FILLER_28_103 ();
 sg13g2_fill_1 FILLER_28_140 ();
 sg13g2_fill_1 FILLER_28_146 ();
 sg13g2_decap_8 FILLER_28_164 ();
 sg13g2_fill_2 FILLER_28_171 ();
 sg13g2_decap_4 FILLER_28_186 ();
 sg13g2_decap_8 FILLER_28_198 ();
 sg13g2_fill_1 FILLER_28_205 ();
 sg13g2_fill_2 FILLER_28_211 ();
 sg13g2_fill_1 FILLER_28_213 ();
 sg13g2_fill_1 FILLER_28_219 ();
 sg13g2_fill_2 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_230 ();
 sg13g2_decap_8 FILLER_28_241 ();
 sg13g2_decap_4 FILLER_28_248 ();
 sg13g2_decap_8 FILLER_28_265 ();
 sg13g2_fill_2 FILLER_28_272 ();
 sg13g2_fill_1 FILLER_28_274 ();
 sg13g2_decap_8 FILLER_28_279 ();
 sg13g2_fill_1 FILLER_28_286 ();
 sg13g2_fill_1 FILLER_28_291 ();
 sg13g2_decap_8 FILLER_28_300 ();
 sg13g2_decap_8 FILLER_28_307 ();
 sg13g2_decap_8 FILLER_28_335 ();
 sg13g2_fill_2 FILLER_28_342 ();
 sg13g2_fill_1 FILLER_28_344 ();
 sg13g2_fill_2 FILLER_28_353 ();
 sg13g2_fill_1 FILLER_28_355 ();
 sg13g2_fill_2 FILLER_28_360 ();
 sg13g2_fill_1 FILLER_28_362 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_decap_4 FILLER_28_378 ();
 sg13g2_fill_2 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_fill_2 FILLER_29_63 ();
 sg13g2_fill_1 FILLER_29_65 ();
 sg13g2_fill_2 FILLER_29_79 ();
 sg13g2_decap_4 FILLER_29_102 ();
 sg13g2_fill_1 FILLER_29_106 ();
 sg13g2_decap_8 FILLER_29_111 ();
 sg13g2_decap_4 FILLER_29_123 ();
 sg13g2_fill_2 FILLER_29_132 ();
 sg13g2_decap_4 FILLER_29_143 ();
 sg13g2_fill_2 FILLER_29_164 ();
 sg13g2_fill_1 FILLER_29_166 ();
 sg13g2_fill_2 FILLER_29_191 ();
 sg13g2_decap_4 FILLER_29_201 ();
 sg13g2_fill_1 FILLER_29_205 ();
 sg13g2_decap_4 FILLER_29_216 ();
 sg13g2_fill_2 FILLER_29_252 ();
 sg13g2_fill_1 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_285 ();
 sg13g2_fill_1 FILLER_29_320 ();
 sg13g2_decap_8 FILLER_29_325 ();
 sg13g2_fill_2 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_384 ();
 sg13g2_decap_8 FILLER_29_391 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_4 FILLER_30_56 ();
 sg13g2_fill_2 FILLER_30_60 ();
 sg13g2_decap_4 FILLER_30_79 ();
 sg13g2_fill_1 FILLER_30_87 ();
 sg13g2_decap_8 FILLER_30_92 ();
 sg13g2_fill_1 FILLER_30_99 ();
 sg13g2_fill_2 FILLER_30_113 ();
 sg13g2_fill_1 FILLER_30_115 ();
 sg13g2_fill_1 FILLER_30_124 ();
 sg13g2_fill_2 FILLER_30_133 ();
 sg13g2_fill_1 FILLER_30_143 ();
 sg13g2_decap_8 FILLER_30_164 ();
 sg13g2_fill_2 FILLER_30_171 ();
 sg13g2_fill_1 FILLER_30_173 ();
 sg13g2_fill_2 FILLER_30_182 ();
 sg13g2_fill_1 FILLER_30_184 ();
 sg13g2_decap_8 FILLER_30_214 ();
 sg13g2_fill_2 FILLER_30_221 ();
 sg13g2_fill_1 FILLER_30_223 ();
 sg13g2_fill_2 FILLER_30_228 ();
 sg13g2_fill_1 FILLER_30_230 ();
 sg13g2_decap_4 FILLER_30_236 ();
 sg13g2_fill_1 FILLER_30_240 ();
 sg13g2_decap_4 FILLER_30_245 ();
 sg13g2_fill_2 FILLER_30_249 ();
 sg13g2_fill_2 FILLER_30_256 ();
 sg13g2_decap_8 FILLER_30_263 ();
 sg13g2_decap_8 FILLER_30_270 ();
 sg13g2_decap_4 FILLER_30_277 ();
 sg13g2_fill_1 FILLER_30_281 ();
 sg13g2_decap_4 FILLER_30_303 ();
 sg13g2_decap_4 FILLER_30_328 ();
 sg13g2_decap_4 FILLER_30_341 ();
 sg13g2_fill_1 FILLER_30_345 ();
 sg13g2_decap_4 FILLER_30_358 ();
 sg13g2_fill_2 FILLER_30_362 ();
 sg13g2_decap_8 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_30_375 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_63 ();
 sg13g2_decap_4 FILLER_31_81 ();
 sg13g2_fill_2 FILLER_31_85 ();
 sg13g2_decap_4 FILLER_31_92 ();
 sg13g2_fill_1 FILLER_31_96 ();
 sg13g2_decap_4 FILLER_31_114 ();
 sg13g2_fill_1 FILLER_31_118 ();
 sg13g2_decap_4 FILLER_31_123 ();
 sg13g2_decap_8 FILLER_31_131 ();
 sg13g2_decap_8 FILLER_31_138 ();
 sg13g2_fill_2 FILLER_31_145 ();
 sg13g2_fill_2 FILLER_31_152 ();
 sg13g2_fill_2 FILLER_31_159 ();
 sg13g2_fill_2 FILLER_31_215 ();
 sg13g2_fill_2 FILLER_31_249 ();
 sg13g2_fill_1 FILLER_31_251 ();
 sg13g2_decap_4 FILLER_31_280 ();
 sg13g2_decap_4 FILLER_31_296 ();
 sg13g2_fill_1 FILLER_31_300 ();
 sg13g2_fill_2 FILLER_31_305 ();
 sg13g2_fill_2 FILLER_31_319 ();
 sg13g2_fill_1 FILLER_31_321 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_4 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_4 FILLER_32_91 ();
 sg13g2_fill_1 FILLER_32_95 ();
 sg13g2_fill_2 FILLER_32_118 ();
 sg13g2_fill_2 FILLER_32_129 ();
 sg13g2_fill_1 FILLER_32_131 ();
 sg13g2_fill_2 FILLER_32_157 ();
 sg13g2_decap_8 FILLER_32_164 ();
 sg13g2_decap_4 FILLER_32_171 ();
 sg13g2_decap_4 FILLER_32_179 ();
 sg13g2_fill_1 FILLER_32_183 ();
 sg13g2_decap_4 FILLER_32_188 ();
 sg13g2_fill_2 FILLER_32_192 ();
 sg13g2_decap_4 FILLER_32_198 ();
 sg13g2_fill_1 FILLER_32_202 ();
 sg13g2_fill_2 FILLER_32_207 ();
 sg13g2_decap_4 FILLER_32_213 ();
 sg13g2_fill_1 FILLER_32_217 ();
 sg13g2_decap_4 FILLER_32_226 ();
 sg13g2_fill_2 FILLER_32_234 ();
 sg13g2_decap_8 FILLER_32_269 ();
 sg13g2_fill_1 FILLER_32_276 ();
 sg13g2_decap_8 FILLER_32_282 ();
 sg13g2_fill_2 FILLER_32_289 ();
 sg13g2_fill_1 FILLER_32_291 ();
 sg13g2_decap_4 FILLER_32_296 ();
 sg13g2_fill_2 FILLER_32_300 ();
 sg13g2_decap_8 FILLER_32_307 ();
 sg13g2_fill_2 FILLER_32_314 ();
 sg13g2_fill_1 FILLER_32_316 ();
 sg13g2_decap_8 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_328 ();
 sg13g2_fill_1 FILLER_32_330 ();
 sg13g2_decap_8 FILLER_32_339 ();
 sg13g2_fill_1 FILLER_32_346 ();
 sg13g2_decap_4 FILLER_32_351 ();
 sg13g2_fill_1 FILLER_32_355 ();
 sg13g2_decap_8 FILLER_32_360 ();
 sg13g2_fill_1 FILLER_32_367 ();
 sg13g2_decap_8 FILLER_32_372 ();
 sg13g2_decap_8 FILLER_32_379 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_decap_8 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_4 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_60 ();
 sg13g2_decap_4 FILLER_33_87 ();
 sg13g2_fill_1 FILLER_33_91 ();
 sg13g2_decap_4 FILLER_33_113 ();
 sg13g2_fill_2 FILLER_33_117 ();
 sg13g2_fill_2 FILLER_33_140 ();
 sg13g2_fill_1 FILLER_33_142 ();
 sg13g2_decap_8 FILLER_33_148 ();
 sg13g2_fill_1 FILLER_33_155 ();
 sg13g2_decap_8 FILLER_33_233 ();
 sg13g2_decap_8 FILLER_33_248 ();
 sg13g2_decap_8 FILLER_33_255 ();
 sg13g2_fill_2 FILLER_33_262 ();
 sg13g2_fill_1 FILLER_33_264 ();
 sg13g2_fill_2 FILLER_33_268 ();
 sg13g2_fill_1 FILLER_33_270 ();
 sg13g2_fill_1 FILLER_33_295 ();
 sg13g2_fill_1 FILLER_33_351 ();
 sg13g2_decap_8 FILLER_33_361 ();
 sg13g2_decap_8 FILLER_33_368 ();
 sg13g2_decap_8 FILLER_33_375 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_fill_2 FILLER_34_63 ();
 sg13g2_fill_1 FILLER_34_65 ();
 sg13g2_decap_8 FILLER_34_82 ();
 sg13g2_decap_4 FILLER_34_89 ();
 sg13g2_fill_1 FILLER_34_93 ();
 sg13g2_decap_8 FILLER_34_111 ();
 sg13g2_fill_2 FILLER_34_118 ();
 sg13g2_fill_1 FILLER_34_120 ();
 sg13g2_decap_8 FILLER_34_138 ();
 sg13g2_fill_1 FILLER_34_145 ();
 sg13g2_decap_8 FILLER_34_155 ();
 sg13g2_fill_2 FILLER_34_162 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_4 FILLER_34_196 ();
 sg13g2_fill_2 FILLER_34_200 ();
 sg13g2_decap_8 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_221 ();
 sg13g2_decap_4 FILLER_34_226 ();
 sg13g2_fill_1 FILLER_34_259 ();
 sg13g2_fill_2 FILLER_34_289 ();
 sg13g2_fill_2 FILLER_34_301 ();
 sg13g2_fill_1 FILLER_34_311 ();
 sg13g2_decap_4 FILLER_34_316 ();
 sg13g2_fill_1 FILLER_34_320 ();
 sg13g2_fill_1 FILLER_34_333 ();
 sg13g2_fill_1 FILLER_34_338 ();
 sg13g2_decap_4 FILLER_34_343 ();
 sg13g2_fill_1 FILLER_34_347 ();
 sg13g2_decap_8 FILLER_34_376 ();
 sg13g2_decap_8 FILLER_34_383 ();
 sg13g2_decap_8 FILLER_34_390 ();
 sg13g2_decap_8 FILLER_34_397 ();
 sg13g2_decap_4 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_4 FILLER_35_56 ();
 sg13g2_fill_1 FILLER_35_60 ();
 sg13g2_decap_4 FILLER_35_87 ();
 sg13g2_fill_2 FILLER_35_91 ();
 sg13g2_fill_2 FILLER_35_118 ();
 sg13g2_fill_1 FILLER_35_120 ();
 sg13g2_fill_1 FILLER_35_139 ();
 sg13g2_decap_8 FILLER_35_165 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_decap_8 FILLER_35_178 ();
 sg13g2_decap_8 FILLER_35_185 ();
 sg13g2_fill_1 FILLER_35_192 ();
 sg13g2_decap_8 FILLER_35_221 ();
 sg13g2_fill_2 FILLER_35_228 ();
 sg13g2_fill_1 FILLER_35_230 ();
 sg13g2_fill_2 FILLER_35_237 ();
 sg13g2_decap_8 FILLER_35_247 ();
 sg13g2_fill_2 FILLER_35_254 ();
 sg13g2_fill_1 FILLER_35_256 ();
 sg13g2_decap_8 FILLER_35_260 ();
 sg13g2_fill_1 FILLER_35_267 ();
 sg13g2_fill_1 FILLER_35_292 ();
 sg13g2_fill_1 FILLER_35_320 ();
 sg13g2_decap_4 FILLER_35_350 ();
 sg13g2_fill_2 FILLER_35_354 ();
 sg13g2_decap_4 FILLER_35_360 ();
 sg13g2_fill_1 FILLER_35_368 ();
 sg13g2_decap_8 FILLER_35_374 ();
 sg13g2_decap_8 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_35_395 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_fill_1 FILLER_36_63 ();
 sg13g2_decap_4 FILLER_36_81 ();
 sg13g2_fill_1 FILLER_36_85 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_115 ();
 sg13g2_decap_4 FILLER_36_122 ();
 sg13g2_fill_1 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_131 ();
 sg13g2_decap_8 FILLER_36_138 ();
 sg13g2_decap_4 FILLER_36_162 ();
 sg13g2_decap_8 FILLER_36_188 ();
 sg13g2_decap_4 FILLER_36_195 ();
 sg13g2_fill_1 FILLER_36_199 ();
 sg13g2_decap_8 FILLER_36_215 ();
 sg13g2_fill_1 FILLER_36_241 ();
 sg13g2_decap_4 FILLER_36_267 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_fill_2 FILLER_36_306 ();
 sg13g2_decap_8 FILLER_36_319 ();
 sg13g2_decap_8 FILLER_36_326 ();
 sg13g2_fill_1 FILLER_36_337 ();
 sg13g2_fill_2 FILLER_36_359 ();
 sg13g2_fill_1 FILLER_36_361 ();
 sg13g2_fill_1 FILLER_36_372 ();
 sg13g2_decap_8 FILLER_36_397 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_fill_2 FILLER_37_63 ();
 sg13g2_fill_2 FILLER_37_82 ();
 sg13g2_decap_4 FILLER_37_115 ();
 sg13g2_fill_1 FILLER_37_119 ();
 sg13g2_decap_4 FILLER_37_124 ();
 sg13g2_fill_1 FILLER_37_174 ();
 sg13g2_decap_8 FILLER_37_183 ();
 sg13g2_decap_4 FILLER_37_190 ();
 sg13g2_fill_2 FILLER_37_194 ();
 sg13g2_decap_8 FILLER_37_226 ();
 sg13g2_fill_2 FILLER_37_233 ();
 sg13g2_decap_8 FILLER_37_247 ();
 sg13g2_decap_8 FILLER_37_254 ();
 sg13g2_fill_2 FILLER_37_261 ();
 sg13g2_fill_1 FILLER_37_263 ();
 sg13g2_fill_2 FILLER_37_290 ();
 sg13g2_fill_1 FILLER_37_292 ();
 sg13g2_fill_2 FILLER_37_309 ();
 sg13g2_fill_1 FILLER_37_311 ();
 sg13g2_fill_2 FILLER_37_341 ();
 sg13g2_fill_1 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_348 ();
 sg13g2_fill_1 FILLER_37_355 ();
 sg13g2_decap_8 FILLER_37_360 ();
 sg13g2_fill_1 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_380 ();
 sg13g2_decap_8 FILLER_37_387 ();
 sg13g2_decap_8 FILLER_37_394 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_4 FILLER_38_49 ();
 sg13g2_fill_2 FILLER_38_85 ();
 sg13g2_fill_2 FILLER_38_103 ();
 sg13g2_fill_2 FILLER_38_135 ();
 sg13g2_fill_1 FILLER_38_137 ();
 sg13g2_decap_8 FILLER_38_204 ();
 sg13g2_decap_8 FILLER_38_211 ();
 sg13g2_decap_8 FILLER_38_218 ();
 sg13g2_decap_4 FILLER_38_225 ();
 sg13g2_decap_8 FILLER_38_275 ();
 sg13g2_decap_4 FILLER_38_282 ();
 sg13g2_fill_1 FILLER_38_286 ();
 sg13g2_fill_2 FILLER_38_291 ();
 sg13g2_fill_1 FILLER_38_293 ();
 sg13g2_fill_2 FILLER_38_303 ();
 sg13g2_fill_1 FILLER_38_305 ();
 sg13g2_decap_4 FILLER_38_310 ();
 sg13g2_fill_2 FILLER_38_314 ();
 sg13g2_decap_4 FILLER_38_320 ();
 sg13g2_fill_1 FILLER_38_324 ();
 sg13g2_decap_4 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_353 ();
 sg13g2_decap_4 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uio_out[7] = net18;
endmodule

module tt_um_dff_mem (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \RAM[0][0] ;
 wire \RAM[0][1] ;
 wire \RAM[0][2] ;
 wire \RAM[0][3] ;
 wire \RAM[0][4] ;
 wire \RAM[0][5] ;
 wire \RAM[0][6] ;
 wire \RAM[0][7] ;
 wire \RAM[10][0] ;
 wire \RAM[10][1] ;
 wire \RAM[10][2] ;
 wire \RAM[10][3] ;
 wire \RAM[10][4] ;
 wire \RAM[10][5] ;
 wire \RAM[10][6] ;
 wire \RAM[10][7] ;
 wire \RAM[11][0] ;
 wire \RAM[11][1] ;
 wire \RAM[11][2] ;
 wire \RAM[11][3] ;
 wire \RAM[11][4] ;
 wire \RAM[11][5] ;
 wire \RAM[11][6] ;
 wire \RAM[11][7] ;
 wire \RAM[12][0] ;
 wire \RAM[12][1] ;
 wire \RAM[12][2] ;
 wire \RAM[12][3] ;
 wire \RAM[12][4] ;
 wire \RAM[12][5] ;
 wire \RAM[12][6] ;
 wire \RAM[12][7] ;
 wire \RAM[13][0] ;
 wire \RAM[13][1] ;
 wire \RAM[13][2] ;
 wire \RAM[13][3] ;
 wire \RAM[13][4] ;
 wire \RAM[13][5] ;
 wire \RAM[13][6] ;
 wire \RAM[13][7] ;
 wire \RAM[14][0] ;
 wire \RAM[14][1] ;
 wire \RAM[14][2] ;
 wire \RAM[14][3] ;
 wire \RAM[14][4] ;
 wire \RAM[14][5] ;
 wire \RAM[14][6] ;
 wire \RAM[14][7] ;
 wire \RAM[15][0] ;
 wire \RAM[15][1] ;
 wire \RAM[15][2] ;
 wire \RAM[15][3] ;
 wire \RAM[15][4] ;
 wire \RAM[15][5] ;
 wire \RAM[15][6] ;
 wire \RAM[15][7] ;
 wire \RAM[1][0] ;
 wire \RAM[1][1] ;
 wire \RAM[1][2] ;
 wire \RAM[1][3] ;
 wire \RAM[1][4] ;
 wire \RAM[1][5] ;
 wire \RAM[1][6] ;
 wire \RAM[1][7] ;
 wire \RAM[2][0] ;
 wire \RAM[2][1] ;
 wire \RAM[2][2] ;
 wire \RAM[2][3] ;
 wire \RAM[2][4] ;
 wire \RAM[2][5] ;
 wire \RAM[2][6] ;
 wire \RAM[2][7] ;
 wire \RAM[3][0] ;
 wire \RAM[3][1] ;
 wire \RAM[3][2] ;
 wire \RAM[3][3] ;
 wire \RAM[3][4] ;
 wire \RAM[3][5] ;
 wire \RAM[3][6] ;
 wire \RAM[3][7] ;
 wire \RAM[4][0] ;
 wire \RAM[4][1] ;
 wire \RAM[4][2] ;
 wire \RAM[4][3] ;
 wire \RAM[4][4] ;
 wire \RAM[4][5] ;
 wire \RAM[4][6] ;
 wire \RAM[4][7] ;
 wire \RAM[5][0] ;
 wire \RAM[5][1] ;
 wire \RAM[5][2] ;
 wire \RAM[5][3] ;
 wire \RAM[5][4] ;
 wire \RAM[5][5] ;
 wire \RAM[5][6] ;
 wire \RAM[5][7] ;
 wire \RAM[6][0] ;
 wire \RAM[6][1] ;
 wire \RAM[6][2] ;
 wire \RAM[6][3] ;
 wire \RAM[6][4] ;
 wire \RAM[6][5] ;
 wire \RAM[6][6] ;
 wire \RAM[6][7] ;
 wire \RAM[7][0] ;
 wire \RAM[7][1] ;
 wire \RAM[7][2] ;
 wire \RAM[7][3] ;
 wire \RAM[7][4] ;
 wire \RAM[7][5] ;
 wire \RAM[7][6] ;
 wire \RAM[7][7] ;
 wire \RAM[8][0] ;
 wire \RAM[8][1] ;
 wire \RAM[8][2] ;
 wire \RAM[8][3] ;
 wire \RAM[8][4] ;
 wire \RAM[8][5] ;
 wire \RAM[8][6] ;
 wire \RAM[8][7] ;
 wire \RAM[9][0] ;
 wire \RAM[9][1] ;
 wire \RAM[9][2] ;
 wire \RAM[9][3] ;
 wire \RAM[9][4] ;
 wire \RAM[9][5] ;
 wire \RAM[9][6] ;
 wire \RAM[9][7] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire clknet_0_clk;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;

 sg13g2_inv_1 _0660_ (.Y(_0136_),
    .A(net13));
 sg13g2_inv_1 _0661_ (.Y(_0137_),
    .A(net12));
 sg13g2_inv_1 _0662_ (.Y(_0138_),
    .A(net11));
 sg13g2_inv_1 _0663_ (.Y(_0139_),
    .A(net10));
 sg13g2_inv_1 _0664_ (.Y(_0140_),
    .A(net9));
 sg13g2_inv_2 _0665_ (.Y(_0141_),
    .A(net8));
 sg13g2_inv_1 _0666_ (.Y(_0142_),
    .A(net7));
 sg13g2_inv_1 _0667_ (.Y(_0143_),
    .A(net6));
 sg13g2_nor2b_1 _0668_ (.A(net2),
    .B_N(net1),
    .Y(_0144_));
 sg13g2_nor2_1 _0669_ (.A(net1),
    .B(net2),
    .Y(_0145_));
 sg13g2_a22oi_1 _0670_ (.Y(_0146_),
    .B1(net350),
    .B2(\RAM[4][0] ),
    .A2(net356),
    .A1(\RAM[5][0] ));
 sg13g2_and2_1 _0671_ (.A(net1),
    .B(net2),
    .X(_0147_));
 sg13g2_nor2b_1 _0672_ (.A(net1),
    .B_N(net2),
    .Y(_0148_));
 sg13g2_a22oi_1 _0673_ (.Y(_0149_),
    .B1(net339),
    .B2(\RAM[6][0] ),
    .A2(net345),
    .A1(\RAM[7][0] ));
 sg13g2_nor2b_2 _0674_ (.A(net4),
    .B_N(net3),
    .Y(_0150_));
 sg13g2_nand2b_2 _0675_ (.Y(_0151_),
    .B(net377),
    .A_N(net376));
 sg13g2_a21oi_1 _0676_ (.A1(_0146_),
    .A2(_0149_),
    .Y(_0152_),
    .B1(_0151_));
 sg13g2_a22oi_1 _0677_ (.Y(_0153_),
    .B1(net353),
    .B2(\RAM[0][0] ),
    .A2(net359),
    .A1(\RAM[1][0] ));
 sg13g2_a22oi_1 _0678_ (.Y(_0154_),
    .B1(net341),
    .B2(\RAM[2][0] ),
    .A2(net347),
    .A1(\RAM[3][0] ));
 sg13g2_nor2_2 _0679_ (.A(net376),
    .B(net377),
    .Y(_0155_));
 sg13g2_or2_2 _0680_ (.X(_0156_),
    .B(net377),
    .A(net376));
 sg13g2_a21oi_1 _0681_ (.A1(_0153_),
    .A2(_0154_),
    .Y(_0157_),
    .B1(_0156_));
 sg13g2_a22oi_1 _0682_ (.Y(_0158_),
    .B1(net351),
    .B2(\RAM[12][0] ),
    .A2(net357),
    .A1(\RAM[13][0] ));
 sg13g2_a22oi_1 _0683_ (.Y(_0159_),
    .B1(net341),
    .B2(\RAM[14][0] ),
    .A2(net347),
    .A1(\RAM[15][0] ));
 sg13g2_nand2_2 _0684_ (.Y(_0160_),
    .A(net4),
    .B(net377));
 sg13g2_a21oi_1 _0685_ (.A1(_0158_),
    .A2(_0159_),
    .Y(_0161_),
    .B1(_0160_));
 sg13g2_a22oi_1 _0686_ (.Y(_0162_),
    .B1(net349),
    .B2(\RAM[8][0] ),
    .A2(net355),
    .A1(\RAM[9][0] ));
 sg13g2_a22oi_1 _0687_ (.Y(_0163_),
    .B1(net338),
    .B2(\RAM[10][0] ),
    .A2(net344),
    .A1(\RAM[11][0] ));
 sg13g2_nor2b_2 _0688_ (.A(net377),
    .B_N(net376),
    .Y(_0164_));
 sg13g2_nand2b_2 _0689_ (.Y(_0165_),
    .B(net376),
    .A_N(net377));
 sg13g2_a21oi_1 _0690_ (.A1(_0162_),
    .A2(_0163_),
    .Y(_0166_),
    .B1(_0165_));
 sg13g2_or4_1 _0691_ (.A(_0152_),
    .B(_0157_),
    .C(_0161_),
    .D(_0166_),
    .X(_0000_));
 sg13g2_a22oi_1 _0692_ (.Y(_0167_),
    .B1(net350),
    .B2(\RAM[4][1] ),
    .A2(net356),
    .A1(\RAM[5][1] ));
 sg13g2_a22oi_1 _0693_ (.Y(_0168_),
    .B1(net339),
    .B2(\RAM[6][1] ),
    .A2(net345),
    .A1(\RAM[7][1] ));
 sg13g2_a21oi_1 _0694_ (.A1(_0167_),
    .A2(_0168_),
    .Y(_0169_),
    .B1(_0151_));
 sg13g2_a22oi_1 _0695_ (.Y(_0170_),
    .B1(net353),
    .B2(\RAM[0][1] ),
    .A2(net359),
    .A1(\RAM[1][1] ));
 sg13g2_a22oi_1 _0696_ (.Y(_0171_),
    .B1(net341),
    .B2(\RAM[2][1] ),
    .A2(net347),
    .A1(\RAM[3][1] ));
 sg13g2_a21oi_2 _0697_ (.B1(_0156_),
    .Y(_0172_),
    .A2(_0171_),
    .A1(_0170_));
 sg13g2_a22oi_1 _0698_ (.Y(_0173_),
    .B1(net351),
    .B2(\RAM[12][1] ),
    .A2(net357),
    .A1(\RAM[13][1] ));
 sg13g2_a22oi_1 _0699_ (.Y(_0174_),
    .B1(net339),
    .B2(\RAM[14][1] ),
    .A2(net345),
    .A1(\RAM[15][1] ));
 sg13g2_a21oi_1 _0700_ (.A1(_0173_),
    .A2(_0174_),
    .Y(_0175_),
    .B1(_0160_));
 sg13g2_a22oi_1 _0701_ (.Y(_0176_),
    .B1(net349),
    .B2(\RAM[8][1] ),
    .A2(net355),
    .A1(\RAM[9][1] ));
 sg13g2_a22oi_1 _0702_ (.Y(_0177_),
    .B1(net338),
    .B2(\RAM[10][1] ),
    .A2(net344),
    .A1(\RAM[11][1] ));
 sg13g2_a21oi_2 _0703_ (.B1(_0165_),
    .Y(_0178_),
    .A2(_0177_),
    .A1(_0176_));
 sg13g2_or4_1 _0704_ (.A(_0169_),
    .B(_0172_),
    .C(_0175_),
    .D(_0178_),
    .X(_0001_));
 sg13g2_a22oi_1 _0705_ (.Y(_0179_),
    .B1(net350),
    .B2(\RAM[4][2] ),
    .A2(net356),
    .A1(\RAM[5][2] ));
 sg13g2_a22oi_1 _0706_ (.Y(_0180_),
    .B1(net339),
    .B2(\RAM[6][2] ),
    .A2(net345),
    .A1(\RAM[7][2] ));
 sg13g2_a21oi_1 _0707_ (.A1(_0179_),
    .A2(_0180_),
    .Y(_0181_),
    .B1(_0151_));
 sg13g2_a22oi_1 _0708_ (.Y(_0182_),
    .B1(net348),
    .B2(\RAM[0][2] ),
    .A2(net354),
    .A1(\RAM[1][2] ));
 sg13g2_a22oi_1 _0709_ (.Y(_0183_),
    .B1(net336),
    .B2(\RAM[2][2] ),
    .A2(net342),
    .A1(\RAM[3][2] ));
 sg13g2_a21oi_2 _0710_ (.B1(_0156_),
    .Y(_0184_),
    .A2(_0183_),
    .A1(_0182_));
 sg13g2_a22oi_1 _0711_ (.Y(_0185_),
    .B1(net351),
    .B2(\RAM[12][2] ),
    .A2(net357),
    .A1(\RAM[13][2] ));
 sg13g2_a22oi_1 _0712_ (.Y(_0186_),
    .B1(net339),
    .B2(\RAM[14][2] ),
    .A2(net345),
    .A1(\RAM[15][2] ));
 sg13g2_a21oi_1 _0713_ (.A1(_0185_),
    .A2(_0186_),
    .Y(_0187_),
    .B1(_0160_));
 sg13g2_a22oi_1 _0714_ (.Y(_0188_),
    .B1(net348),
    .B2(\RAM[8][2] ),
    .A2(net354),
    .A1(\RAM[9][2] ));
 sg13g2_a22oi_1 _0715_ (.Y(_0189_),
    .B1(net336),
    .B2(\RAM[10][2] ),
    .A2(net342),
    .A1(\RAM[11][2] ));
 sg13g2_a21oi_2 _0716_ (.B1(_0165_),
    .Y(_0190_),
    .A2(_0189_),
    .A1(_0188_));
 sg13g2_or4_1 _0717_ (.A(_0181_),
    .B(_0184_),
    .C(_0187_),
    .D(_0190_),
    .X(_0002_));
 sg13g2_a22oi_1 _0718_ (.Y(_0191_),
    .B1(net350),
    .B2(\RAM[4][3] ),
    .A2(net356),
    .A1(\RAM[5][3] ));
 sg13g2_a22oi_1 _0719_ (.Y(_0192_),
    .B1(net340),
    .B2(\RAM[6][3] ),
    .A2(net346),
    .A1(\RAM[7][3] ));
 sg13g2_a21oi_1 _0720_ (.A1(_0191_),
    .A2(_0192_),
    .Y(_0193_),
    .B1(_0151_));
 sg13g2_a22oi_1 _0721_ (.Y(_0194_),
    .B1(net348),
    .B2(\RAM[0][3] ),
    .A2(net354),
    .A1(\RAM[1][3] ));
 sg13g2_a22oi_1 _0722_ (.Y(_0195_),
    .B1(net336),
    .B2(\RAM[2][3] ),
    .A2(net342),
    .A1(\RAM[3][3] ));
 sg13g2_a21oi_2 _0723_ (.B1(_0156_),
    .Y(_0196_),
    .A2(_0195_),
    .A1(_0194_));
 sg13g2_a22oi_1 _0724_ (.Y(_0197_),
    .B1(net350),
    .B2(\RAM[12][3] ),
    .A2(net356),
    .A1(\RAM[13][3] ));
 sg13g2_a22oi_1 _0725_ (.Y(_0198_),
    .B1(net339),
    .B2(\RAM[14][3] ),
    .A2(net345),
    .A1(\RAM[15][3] ));
 sg13g2_a21oi_1 _0726_ (.A1(_0197_),
    .A2(_0198_),
    .Y(_0199_),
    .B1(_0160_));
 sg13g2_a22oi_1 _0727_ (.Y(_0200_),
    .B1(net349),
    .B2(\RAM[8][3] ),
    .A2(net355),
    .A1(\RAM[9][3] ));
 sg13g2_a22oi_1 _0728_ (.Y(_0201_),
    .B1(net337),
    .B2(\RAM[10][3] ),
    .A2(net343),
    .A1(\RAM[11][3] ));
 sg13g2_a21oi_1 _0729_ (.A1(_0200_),
    .A2(_0201_),
    .Y(_0202_),
    .B1(_0165_));
 sg13g2_or4_1 _0730_ (.A(_0193_),
    .B(_0196_),
    .C(_0199_),
    .D(_0202_),
    .X(_0003_));
 sg13g2_a22oi_1 _0731_ (.Y(_0203_),
    .B1(net350),
    .B2(\RAM[4][4] ),
    .A2(net356),
    .A1(\RAM[5][4] ));
 sg13g2_a22oi_1 _0732_ (.Y(_0204_),
    .B1(net339),
    .B2(\RAM[6][4] ),
    .A2(net345),
    .A1(\RAM[7][4] ));
 sg13g2_a21oi_1 _0733_ (.A1(_0203_),
    .A2(_0204_),
    .Y(_0205_),
    .B1(_0151_));
 sg13g2_a22oi_1 _0734_ (.Y(_0206_),
    .B1(net348),
    .B2(\RAM[0][4] ),
    .A2(net354),
    .A1(\RAM[1][4] ));
 sg13g2_a22oi_1 _0735_ (.Y(_0207_),
    .B1(net336),
    .B2(\RAM[2][4] ),
    .A2(net342),
    .A1(\RAM[3][4] ));
 sg13g2_a21oi_1 _0736_ (.A1(_0206_),
    .A2(_0207_),
    .Y(_0208_),
    .B1(_0156_));
 sg13g2_a22oi_1 _0737_ (.Y(_0209_),
    .B1(net350),
    .B2(\RAM[12][4] ),
    .A2(net356),
    .A1(\RAM[13][4] ));
 sg13g2_a22oi_1 _0738_ (.Y(_0210_),
    .B1(net340),
    .B2(\RAM[14][4] ),
    .A2(net346),
    .A1(\RAM[15][4] ));
 sg13g2_a21oi_1 _0739_ (.A1(_0209_),
    .A2(_0210_),
    .Y(_0211_),
    .B1(_0160_));
 sg13g2_a22oi_1 _0740_ (.Y(_0212_),
    .B1(net349),
    .B2(\RAM[8][4] ),
    .A2(net355),
    .A1(\RAM[9][4] ));
 sg13g2_a22oi_1 _0741_ (.Y(_0213_),
    .B1(net337),
    .B2(\RAM[10][4] ),
    .A2(net343),
    .A1(\RAM[11][4] ));
 sg13g2_a21oi_1 _0742_ (.A1(_0212_),
    .A2(_0213_),
    .Y(_0214_),
    .B1(_0165_));
 sg13g2_or4_1 _0743_ (.A(_0205_),
    .B(_0208_),
    .C(_0211_),
    .D(_0214_),
    .X(_0004_));
 sg13g2_a22oi_1 _0744_ (.Y(_0215_),
    .B1(net352),
    .B2(\RAM[4][5] ),
    .A2(net358),
    .A1(\RAM[5][5] ));
 sg13g2_a22oi_1 _0745_ (.Y(_0216_),
    .B1(net340),
    .B2(\RAM[6][5] ),
    .A2(net346),
    .A1(\RAM[7][5] ));
 sg13g2_a21oi_1 _0746_ (.A1(_0215_),
    .A2(_0216_),
    .Y(_0217_),
    .B1(_0151_));
 sg13g2_a22oi_1 _0747_ (.Y(_0218_),
    .B1(net349),
    .B2(\RAM[0][5] ),
    .A2(net359),
    .A1(\RAM[1][5] ));
 sg13g2_a22oi_1 _0748_ (.Y(_0219_),
    .B1(net336),
    .B2(\RAM[2][5] ),
    .A2(net342),
    .A1(\RAM[3][5] ));
 sg13g2_a21oi_1 _0749_ (.A1(_0218_),
    .A2(_0219_),
    .Y(_0220_),
    .B1(_0156_));
 sg13g2_a22oi_1 _0750_ (.Y(_0221_),
    .B1(net352),
    .B2(\RAM[12][5] ),
    .A2(net358),
    .A1(\RAM[13][5] ));
 sg13g2_a22oi_1 _0751_ (.Y(_0222_),
    .B1(net340),
    .B2(\RAM[14][5] ),
    .A2(net346),
    .A1(\RAM[15][5] ));
 sg13g2_a21oi_1 _0752_ (.A1(_0221_),
    .A2(_0222_),
    .Y(_0223_),
    .B1(_0160_));
 sg13g2_a22oi_1 _0753_ (.Y(_0224_),
    .B1(net349),
    .B2(\RAM[8][5] ),
    .A2(net355),
    .A1(\RAM[9][5] ));
 sg13g2_a22oi_1 _0754_ (.Y(_0225_),
    .B1(net337),
    .B2(\RAM[10][5] ),
    .A2(net343),
    .A1(\RAM[11][5] ));
 sg13g2_a21oi_1 _0755_ (.A1(_0224_),
    .A2(_0225_),
    .Y(_0226_),
    .B1(_0165_));
 sg13g2_or4_1 _0756_ (.A(_0217_),
    .B(_0220_),
    .C(_0223_),
    .D(_0226_),
    .X(_0005_));
 sg13g2_a22oi_1 _0757_ (.Y(_0227_),
    .B1(net352),
    .B2(\RAM[4][6] ),
    .A2(net358),
    .A1(\RAM[5][6] ));
 sg13g2_a22oi_1 _0758_ (.Y(_0228_),
    .B1(net338),
    .B2(\RAM[6][6] ),
    .A2(net344),
    .A1(\RAM[7][6] ));
 sg13g2_a21oi_1 _0759_ (.A1(_0227_),
    .A2(_0228_),
    .Y(_0229_),
    .B1(_0151_));
 sg13g2_a22oi_1 _0760_ (.Y(_0230_),
    .B1(net348),
    .B2(\RAM[0][6] ),
    .A2(net354),
    .A1(\RAM[1][6] ));
 sg13g2_a22oi_1 _0761_ (.Y(_0231_),
    .B1(net336),
    .B2(\RAM[2][6] ),
    .A2(net342),
    .A1(\RAM[3][6] ));
 sg13g2_a21oi_1 _0762_ (.A1(_0230_),
    .A2(_0231_),
    .Y(_0232_),
    .B1(_0156_));
 sg13g2_a22oi_1 _0763_ (.Y(_0233_),
    .B1(net352),
    .B2(\RAM[12][6] ),
    .A2(net358),
    .A1(\RAM[13][6] ));
 sg13g2_a22oi_1 _0764_ (.Y(_0234_),
    .B1(net340),
    .B2(\RAM[14][6] ),
    .A2(net346),
    .A1(\RAM[15][6] ));
 sg13g2_a21oi_1 _0765_ (.A1(_0233_),
    .A2(_0234_),
    .Y(_0235_),
    .B1(_0160_));
 sg13g2_a22oi_1 _0766_ (.Y(_0236_),
    .B1(net348),
    .B2(\RAM[8][6] ),
    .A2(net354),
    .A1(\RAM[9][6] ));
 sg13g2_a22oi_1 _0767_ (.Y(_0237_),
    .B1(net337),
    .B2(\RAM[10][6] ),
    .A2(net343),
    .A1(\RAM[11][6] ));
 sg13g2_a21oi_1 _0768_ (.A1(_0236_),
    .A2(_0237_),
    .Y(_0238_),
    .B1(_0165_));
 sg13g2_or4_1 _0769_ (.A(_0229_),
    .B(_0232_),
    .C(_0235_),
    .D(_0238_),
    .X(_0006_));
 sg13g2_a22oi_1 _0770_ (.Y(_0239_),
    .B1(net352),
    .B2(\RAM[4][7] ),
    .A2(net358),
    .A1(\RAM[5][7] ));
 sg13g2_a22oi_1 _0771_ (.Y(_0240_),
    .B1(net338),
    .B2(\RAM[6][7] ),
    .A2(net344),
    .A1(\RAM[7][7] ));
 sg13g2_a21oi_1 _0772_ (.A1(_0239_),
    .A2(_0240_),
    .Y(_0241_),
    .B1(_0151_));
 sg13g2_a22oi_1 _0773_ (.Y(_0242_),
    .B1(net348),
    .B2(\RAM[0][7] ),
    .A2(net354),
    .A1(\RAM[1][7] ));
 sg13g2_a22oi_1 _0774_ (.Y(_0243_),
    .B1(net336),
    .B2(\RAM[2][7] ),
    .A2(net342),
    .A1(\RAM[3][7] ));
 sg13g2_a21oi_1 _0775_ (.A1(_0242_),
    .A2(_0243_),
    .Y(_0244_),
    .B1(_0156_));
 sg13g2_a22oi_1 _0776_ (.Y(_0245_),
    .B1(net352),
    .B2(\RAM[12][7] ),
    .A2(net358),
    .A1(\RAM[13][7] ));
 sg13g2_a22oi_1 _0777_ (.Y(_0246_),
    .B1(net340),
    .B2(\RAM[14][7] ),
    .A2(net346),
    .A1(\RAM[15][7] ));
 sg13g2_a21oi_1 _0778_ (.A1(_0245_),
    .A2(_0246_),
    .Y(_0247_),
    .B1(_0160_));
 sg13g2_a22oi_1 _0779_ (.Y(_0248_),
    .B1(net348),
    .B2(\RAM[8][7] ),
    .A2(net354),
    .A1(\RAM[9][7] ));
 sg13g2_a22oi_1 _0780_ (.Y(_0249_),
    .B1(net336),
    .B2(\RAM[10][7] ),
    .A2(net342),
    .A1(\RAM[11][7] ));
 sg13g2_a21oi_1 _0781_ (.A1(_0248_),
    .A2(_0249_),
    .Y(_0250_),
    .B1(_0165_));
 sg13g2_or4_1 _0782_ (.A(_0241_),
    .B(_0244_),
    .C(_0247_),
    .D(_0250_),
    .X(_0007_));
 sg13g2_nor2b_1 _0783_ (.A(net5),
    .B_N(net397),
    .Y(_0251_));
 sg13g2_nand3_1 _0784_ (.B(_0164_),
    .C(net334),
    .A(net349),
    .Y(_0252_));
 sg13g2_nand3_1 _0785_ (.B(net253),
    .C(net333),
    .A(net386),
    .Y(_0253_));
 sg13g2_o21ai_1 _0786_ (.B1(_0253_),
    .Y(_0008_),
    .A1(net360),
    .A2(_0252_));
 sg13g2_nand3_1 _0787_ (.B(net266),
    .C(net333),
    .A(net386),
    .Y(_0254_));
 sg13g2_o21ai_1 _0788_ (.B1(_0254_),
    .Y(_0009_),
    .A1(net362),
    .A2(net333));
 sg13g2_nand3_1 _0789_ (.B(net160),
    .C(net332),
    .A(net384),
    .Y(_0255_));
 sg13g2_o21ai_1 _0790_ (.B1(_0255_),
    .Y(_0010_),
    .A1(net364),
    .A2(net332));
 sg13g2_nand3_1 _0791_ (.B(net274),
    .C(net332),
    .A(net384),
    .Y(_0256_));
 sg13g2_o21ai_1 _0792_ (.B1(_0256_),
    .Y(_0011_),
    .A1(net366),
    .A2(net332));
 sg13g2_nand3_1 _0793_ (.B(net232),
    .C(net333),
    .A(net384),
    .Y(_0257_));
 sg13g2_o21ai_1 _0794_ (.B1(_0257_),
    .Y(_0012_),
    .A1(net368),
    .A2(net333));
 sg13g2_nand3_1 _0795_ (.B(net240),
    .C(net333),
    .A(net386),
    .Y(_0258_));
 sg13g2_o21ai_1 _0796_ (.B1(_0258_),
    .Y(_0013_),
    .A1(net371),
    .A2(net333));
 sg13g2_nand3_1 _0797_ (.B(net257),
    .C(net332),
    .A(net384),
    .Y(_0259_));
 sg13g2_o21ai_1 _0798_ (.B1(_0259_),
    .Y(_0014_),
    .A1(net372),
    .A2(net332));
 sg13g2_nand3_1 _0799_ (.B(net271),
    .C(net332),
    .A(net385),
    .Y(_0260_));
 sg13g2_o21ai_1 _0800_ (.B1(_0260_),
    .Y(_0015_),
    .A1(net374),
    .A2(net332));
 sg13g2_nand4_1 _0801_ (.B(net377),
    .C(net346),
    .A(net4),
    .Y(_0261_),
    .D(net335));
 sg13g2_nand3_1 _0802_ (.B(net275),
    .C(net330),
    .A(net397),
    .Y(_0262_));
 sg13g2_o21ai_1 _0803_ (.B1(_0262_),
    .Y(_0016_),
    .A1(net361),
    .A2(net330));
 sg13g2_nand3_1 _0804_ (.B(net184),
    .C(net330),
    .A(net396),
    .Y(_0263_));
 sg13g2_o21ai_1 _0805_ (.B1(_0263_),
    .Y(_0017_),
    .A1(net363),
    .A2(net330));
 sg13g2_nand3_1 _0806_ (.B(net159),
    .C(net330),
    .A(net398),
    .Y(_0264_));
 sg13g2_o21ai_1 _0807_ (.B1(_0264_),
    .Y(_0018_),
    .A1(net365),
    .A2(_0261_));
 sg13g2_nand3_1 _0808_ (.B(net211),
    .C(net330),
    .A(net396),
    .Y(_0265_));
 sg13g2_o21ai_1 _0809_ (.B1(_0265_),
    .Y(_0019_),
    .A1(net367),
    .A2(net331));
 sg13g2_nand3_1 _0810_ (.B(net218),
    .C(net330),
    .A(net397),
    .Y(_0266_));
 sg13g2_o21ai_1 _0811_ (.B1(_0266_),
    .Y(_0020_),
    .A1(net369),
    .A2(net330));
 sg13g2_nand3_1 _0812_ (.B(net231),
    .C(net331),
    .A(net395),
    .Y(_0267_));
 sg13g2_o21ai_1 _0813_ (.B1(_0267_),
    .Y(_0021_),
    .A1(net371),
    .A2(net331));
 sg13g2_nand3_1 _0814_ (.B(net239),
    .C(net331),
    .A(net395),
    .Y(_0268_));
 sg13g2_o21ai_1 _0815_ (.B1(_0268_),
    .Y(_0022_),
    .A1(net373),
    .A2(net331));
 sg13g2_nand3_1 _0816_ (.B(net180),
    .C(net331),
    .A(net394),
    .Y(_0269_));
 sg13g2_o21ai_1 _0817_ (.B1(_0269_),
    .Y(_0023_),
    .A1(net375),
    .A2(net331));
 sg13g2_nand4_1 _0818_ (.B(net3),
    .C(net351),
    .A(net376),
    .Y(_0270_),
    .D(net335));
 sg13g2_nand3_1 _0819_ (.B(net270),
    .C(net329),
    .A(net396),
    .Y(_0271_));
 sg13g2_o21ai_1 _0820_ (.B1(_0271_),
    .Y(_0024_),
    .A1(net361),
    .A2(net329));
 sg13g2_nand3_1 _0821_ (.B(net198),
    .C(net329),
    .A(net398),
    .Y(_0272_));
 sg13g2_o21ai_1 _0822_ (.B1(_0272_),
    .Y(_0025_),
    .A1(net363),
    .A2(net329));
 sg13g2_nand3_1 _0823_ (.B(net176),
    .C(net329),
    .A(net396),
    .Y(_0273_));
 sg13g2_o21ai_1 _0824_ (.B1(_0273_),
    .Y(_0026_),
    .A1(net365),
    .A2(net329));
 sg13g2_nand3_1 _0825_ (.B(net246),
    .C(net328),
    .A(net396),
    .Y(_0274_));
 sg13g2_o21ai_1 _0826_ (.B1(_0274_),
    .Y(_0027_),
    .A1(net367),
    .A2(net328));
 sg13g2_nand3_1 _0827_ (.B(net281),
    .C(net329),
    .A(net397),
    .Y(_0275_));
 sg13g2_o21ai_1 _0828_ (.B1(_0275_),
    .Y(_0028_),
    .A1(net369),
    .A2(net329));
 sg13g2_nand3_1 _0829_ (.B(net258),
    .C(net328),
    .A(net394),
    .Y(_0276_));
 sg13g2_o21ai_1 _0830_ (.B1(_0276_),
    .Y(_0029_),
    .A1(net371),
    .A2(net328));
 sg13g2_nand3_1 _0831_ (.B(net269),
    .C(net328),
    .A(net394),
    .Y(_0277_));
 sg13g2_o21ai_1 _0832_ (.B1(_0277_),
    .Y(_0030_),
    .A1(net373),
    .A2(net328));
 sg13g2_nand3_1 _0833_ (.B(net261),
    .C(net328),
    .A(net394),
    .Y(_0278_));
 sg13g2_o21ai_1 _0834_ (.B1(_0278_),
    .Y(_0031_),
    .A1(net375),
    .A2(net328));
 sg13g2_nand4_1 _0835_ (.B(net3),
    .C(net357),
    .A(net376),
    .Y(_0279_),
    .D(net335));
 sg13g2_nand3_1 _0836_ (.B(net208),
    .C(net326),
    .A(net396),
    .Y(_0280_));
 sg13g2_o21ai_1 _0837_ (.B1(_0280_),
    .Y(_0032_),
    .A1(net361),
    .A2(net326));
 sg13g2_nand3_1 _0838_ (.B(net182),
    .C(_0279_),
    .A(net398),
    .Y(_0281_));
 sg13g2_o21ai_1 _0839_ (.B1(_0281_),
    .Y(_0033_),
    .A1(net363),
    .A2(net326));
 sg13g2_nand3_1 _0840_ (.B(net256),
    .C(net326),
    .A(net398),
    .Y(_0282_));
 sg13g2_o21ai_1 _0841_ (.B1(_0282_),
    .Y(_0034_),
    .A1(net365),
    .A2(net326));
 sg13g2_nand3_1 _0842_ (.B(net161),
    .C(net326),
    .A(net396),
    .Y(_0283_));
 sg13g2_o21ai_1 _0843_ (.B1(_0283_),
    .Y(_0035_),
    .A1(net367),
    .A2(net327));
 sg13g2_nand3_1 _0844_ (.B(net169),
    .C(net326),
    .A(net396),
    .Y(_0284_));
 sg13g2_o21ai_1 _0845_ (.B1(_0284_),
    .Y(_0036_),
    .A1(net369),
    .A2(net326));
 sg13g2_nand3_1 _0846_ (.B(net224),
    .C(net327),
    .A(net394),
    .Y(_0285_));
 sg13g2_o21ai_1 _0847_ (.B1(_0285_),
    .Y(_0037_),
    .A1(net371),
    .A2(net327));
 sg13g2_nand3_1 _0848_ (.B(net173),
    .C(net327),
    .A(net394),
    .Y(_0286_));
 sg13g2_o21ai_1 _0849_ (.B1(_0286_),
    .Y(_0038_),
    .A1(net373),
    .A2(net327));
 sg13g2_nand3_1 _0850_ (.B(net171),
    .C(net327),
    .A(net394),
    .Y(_0287_));
 sg13g2_o21ai_1 _0851_ (.B1(_0287_),
    .Y(_0039_),
    .A1(net375),
    .A2(net327));
 sg13g2_nand3_1 _0852_ (.B(_0155_),
    .C(net334),
    .A(net353),
    .Y(_0288_));
 sg13g2_nand3_1 _0853_ (.B(net191),
    .C(net325),
    .A(net381),
    .Y(_0289_));
 sg13g2_o21ai_1 _0854_ (.B1(_0289_),
    .Y(_0040_),
    .A1(net360),
    .A2(net325));
 sg13g2_nand3_1 _0855_ (.B(net172),
    .C(net325),
    .A(net381),
    .Y(_0290_));
 sg13g2_o21ai_1 _0856_ (.B1(_0290_),
    .Y(_0041_),
    .A1(net362),
    .A2(_0288_));
 sg13g2_nand3_1 _0857_ (.B(net263),
    .C(net324),
    .A(net378),
    .Y(_0291_));
 sg13g2_o21ai_1 _0858_ (.B1(_0291_),
    .Y(_0042_),
    .A1(net364),
    .A2(net324));
 sg13g2_nand3_1 _0859_ (.B(net236),
    .C(net324),
    .A(net378),
    .Y(_0292_));
 sg13g2_o21ai_1 _0860_ (.B1(_0292_),
    .Y(_0043_),
    .A1(net366),
    .A2(net324));
 sg13g2_nand3_1 _0861_ (.B(net226),
    .C(net325),
    .A(net379),
    .Y(_0293_));
 sg13g2_o21ai_1 _0862_ (.B1(_0293_),
    .Y(_0044_),
    .A1(net368),
    .A2(net325));
 sg13g2_nand3_1 _0863_ (.B(net207),
    .C(net325),
    .A(net381),
    .Y(_0294_));
 sg13g2_o21ai_1 _0864_ (.B1(_0294_),
    .Y(_0045_),
    .A1(net370),
    .A2(net325));
 sg13g2_nand3_1 _0865_ (.B(net277),
    .C(net324),
    .A(net378),
    .Y(_0295_));
 sg13g2_o21ai_1 _0866_ (.B1(_0295_),
    .Y(_0046_),
    .A1(net372),
    .A2(net324));
 sg13g2_nand3_1 _0867_ (.B(net189),
    .C(net324),
    .A(net380),
    .Y(_0296_));
 sg13g2_o21ai_1 _0868_ (.B1(_0296_),
    .Y(_0047_),
    .A1(net374),
    .A2(net324));
 sg13g2_nand3_1 _0869_ (.B(_0164_),
    .C(net334),
    .A(net338),
    .Y(_0297_));
 sg13g2_nand3_1 _0870_ (.B(net259),
    .C(net323),
    .A(net387),
    .Y(_0298_));
 sg13g2_o21ai_1 _0871_ (.B1(_0298_),
    .Y(_0048_),
    .A1(net360),
    .A2(net323));
 sg13g2_nand3_1 _0872_ (.B(net282),
    .C(net323),
    .A(net387),
    .Y(_0299_));
 sg13g2_o21ai_1 _0873_ (.B1(_0299_),
    .Y(_0049_),
    .A1(net362),
    .A2(net323));
 sg13g2_nand3_1 _0874_ (.B(net280),
    .C(net321),
    .A(net386),
    .Y(_0300_));
 sg13g2_o21ai_1 _0875_ (.B1(_0300_),
    .Y(_0050_),
    .A1(net364),
    .A2(net321));
 sg13g2_nand3_1 _0876_ (.B(net174),
    .C(net321),
    .A(net385),
    .Y(_0301_));
 sg13g2_o21ai_1 _0877_ (.B1(_0301_),
    .Y(_0051_),
    .A1(net366),
    .A2(net321));
 sg13g2_nand3_1 _0878_ (.B(net221),
    .C(net321),
    .A(net387),
    .Y(_0302_));
 sg13g2_o21ai_1 _0879_ (.B1(_0302_),
    .Y(_0052_),
    .A1(net368),
    .A2(net321));
 sg13g2_nand3_1 _0880_ (.B(net196),
    .C(net321),
    .A(net387),
    .Y(_0303_));
 sg13g2_o21ai_1 _0881_ (.B1(_0303_),
    .Y(_0053_),
    .A1(net371),
    .A2(net322));
 sg13g2_nand3_1 _0882_ (.B(net272),
    .C(net322),
    .A(net385),
    .Y(_0304_));
 sg13g2_o21ai_1 _0883_ (.B1(_0304_),
    .Y(_0054_),
    .A1(net372),
    .A2(net322));
 sg13g2_nand3_1 _0884_ (.B(net283),
    .C(net322),
    .A(net385),
    .Y(_0305_));
 sg13g2_o21ai_1 _0885_ (.B1(_0305_),
    .Y(_0055_),
    .A1(net374),
    .A2(net321));
 sg13g2_nand3_1 _0886_ (.B(_0164_),
    .C(net334),
    .A(net344),
    .Y(_0306_));
 sg13g2_nand3_1 _0887_ (.B(net279),
    .C(net320),
    .A(net387),
    .Y(_0307_));
 sg13g2_o21ai_1 _0888_ (.B1(_0307_),
    .Y(_0056_),
    .A1(net360),
    .A2(net320));
 sg13g2_nand3_1 _0889_ (.B(net165),
    .C(net320),
    .A(net386),
    .Y(_0308_));
 sg13g2_o21ai_1 _0890_ (.B1(_0308_),
    .Y(_0057_),
    .A1(net362),
    .A2(net320));
 sg13g2_nand3_1 _0891_ (.B(net183),
    .C(net319),
    .A(net384),
    .Y(_0309_));
 sg13g2_o21ai_1 _0892_ (.B1(_0309_),
    .Y(_0058_),
    .A1(net364),
    .A2(net319));
 sg13g2_nand3_1 _0893_ (.B(net215),
    .C(net319),
    .A(net384),
    .Y(_0310_));
 sg13g2_o21ai_1 _0894_ (.B1(_0310_),
    .Y(_0059_),
    .A1(net366),
    .A2(net319));
 sg13g2_nand3_1 _0895_ (.B(net252),
    .C(net320),
    .A(net387),
    .Y(_0311_));
 sg13g2_o21ai_1 _0896_ (.B1(_0311_),
    .Y(_0060_),
    .A1(net368),
    .A2(_0306_));
 sg13g2_nand3_1 _0897_ (.B(net216),
    .C(net319),
    .A(net387),
    .Y(_0312_));
 sg13g2_o21ai_1 _0898_ (.B1(_0312_),
    .Y(_0061_),
    .A1(net371),
    .A2(net320));
 sg13g2_nand3_1 _0899_ (.B(net225),
    .C(net320),
    .A(net385),
    .Y(_0313_));
 sg13g2_o21ai_1 _0900_ (.B1(_0313_),
    .Y(_0062_),
    .A1(net372),
    .A2(net319));
 sg13g2_nand3_1 _0901_ (.B(net285),
    .C(net319),
    .A(net385),
    .Y(_0314_));
 sg13g2_o21ai_1 _0902_ (.B1(_0314_),
    .Y(_0063_),
    .A1(net374),
    .A2(net319));
 sg13g2_nand3_1 _0903_ (.B(_0155_),
    .C(net334),
    .A(net355),
    .Y(_0315_));
 sg13g2_nand3_1 _0904_ (.B(net245),
    .C(net318),
    .A(net381),
    .Y(_0316_));
 sg13g2_o21ai_1 _0905_ (.B1(_0316_),
    .Y(_0064_),
    .A1(net360),
    .A2(_0315_));
 sg13g2_nand3_1 _0906_ (.B(net242),
    .C(net318),
    .A(net381),
    .Y(_0317_));
 sg13g2_o21ai_1 _0907_ (.B1(_0317_),
    .Y(_0065_),
    .A1(net362),
    .A2(net318));
 sg13g2_nand3_1 _0908_ (.B(net200),
    .C(net317),
    .A(net378),
    .Y(_0318_));
 sg13g2_o21ai_1 _0909_ (.B1(_0318_),
    .Y(_0066_),
    .A1(net364),
    .A2(net317));
 sg13g2_nand3_1 _0910_ (.B(net268),
    .C(net317),
    .A(net378),
    .Y(_0319_));
 sg13g2_o21ai_1 _0911_ (.B1(_0319_),
    .Y(_0067_),
    .A1(net366),
    .A2(net317));
 sg13g2_nand3_1 _0912_ (.B(net276),
    .C(net318),
    .A(net379),
    .Y(_0320_));
 sg13g2_o21ai_1 _0913_ (.B1(_0320_),
    .Y(_0068_),
    .A1(net368),
    .A2(net318));
 sg13g2_nand3_1 _0914_ (.B(net204),
    .C(net318),
    .A(net381),
    .Y(_0321_));
 sg13g2_o21ai_1 _0915_ (.B1(_0321_),
    .Y(_0069_),
    .A1(net370),
    .A2(net318));
 sg13g2_nand3_1 _0916_ (.B(net243),
    .C(net317),
    .A(net378),
    .Y(_0322_));
 sg13g2_o21ai_1 _0917_ (.B1(_0322_),
    .Y(_0070_),
    .A1(net372),
    .A2(net317));
 sg13g2_nand3_1 _0918_ (.B(net162),
    .C(net317),
    .A(net383),
    .Y(_0323_));
 sg13g2_o21ai_1 _0919_ (.B1(_0323_),
    .Y(_0071_),
    .A1(net374),
    .A2(net317));
 sg13g2_nand4_1 _0920_ (.B(net377),
    .C(net340),
    .A(net376),
    .Y(_0324_),
    .D(net335));
 sg13g2_nand3_1 _0921_ (.B(net284),
    .C(net316),
    .A(net397),
    .Y(_0325_));
 sg13g2_o21ai_1 _0922_ (.B1(_0325_),
    .Y(_0072_),
    .A1(net361),
    .A2(net316));
 sg13g2_nand3_1 _0923_ (.B(net260),
    .C(net316),
    .A(net397),
    .Y(_0326_));
 sg13g2_o21ai_1 _0924_ (.B1(_0326_),
    .Y(_0073_),
    .A1(net363),
    .A2(net316));
 sg13g2_nand3_1 _0925_ (.B(net192),
    .C(net316),
    .A(net398),
    .Y(_0327_));
 sg13g2_o21ai_1 _0926_ (.B1(_0327_),
    .Y(_0074_),
    .A1(net365),
    .A2(net316));
 sg13g2_nand3_1 _0927_ (.B(net195),
    .C(net315),
    .A(net397),
    .Y(_0328_));
 sg13g2_o21ai_1 _0928_ (.B1(_0328_),
    .Y(_0075_),
    .A1(net367),
    .A2(net315));
 sg13g2_nand3_1 _0929_ (.B(net219),
    .C(net316),
    .A(net397),
    .Y(_0329_));
 sg13g2_o21ai_1 _0930_ (.B1(_0329_),
    .Y(_0076_),
    .A1(net369),
    .A2(net316));
 sg13g2_nand3_1 _0931_ (.B(net250),
    .C(net315),
    .A(net395),
    .Y(_0330_));
 sg13g2_o21ai_1 _0932_ (.B1(_0330_),
    .Y(_0077_),
    .A1(net371),
    .A2(net315));
 sg13g2_nand3_1 _0933_ (.B(net212),
    .C(net315),
    .A(net394),
    .Y(_0331_));
 sg13g2_o21ai_1 _0934_ (.B1(_0331_),
    .Y(_0078_),
    .A1(net373),
    .A2(net315));
 sg13g2_nand3_1 _0935_ (.B(net199),
    .C(net315),
    .A(net395),
    .Y(_0332_));
 sg13g2_o21ai_1 _0936_ (.B1(_0332_),
    .Y(_0079_),
    .A1(net375),
    .A2(net315));
 sg13g2_nand3_1 _0937_ (.B(_0155_),
    .C(net334),
    .A(net338),
    .Y(_0333_));
 sg13g2_nand3_1 _0938_ (.B(net244),
    .C(_0333_),
    .A(net382),
    .Y(_0334_));
 sg13g2_o21ai_1 _0939_ (.B1(_0334_),
    .Y(_0080_),
    .A1(net360),
    .A2(net314));
 sg13g2_nand3_1 _0940_ (.B(net229),
    .C(net314),
    .A(net381),
    .Y(_0335_));
 sg13g2_o21ai_1 _0941_ (.B1(_0335_),
    .Y(_0081_),
    .A1(net362),
    .A2(net314));
 sg13g2_nand3_1 _0942_ (.B(net249),
    .C(net313),
    .A(net379),
    .Y(_0336_));
 sg13g2_o21ai_1 _0943_ (.B1(_0336_),
    .Y(_0082_),
    .A1(net364),
    .A2(net313));
 sg13g2_nand3_1 _0944_ (.B(net262),
    .C(net313),
    .A(net379),
    .Y(_0337_));
 sg13g2_o21ai_1 _0945_ (.B1(_0337_),
    .Y(_0083_),
    .A1(net366),
    .A2(net313));
 sg13g2_nand3_1 _0946_ (.B(net238),
    .C(net313),
    .A(net378),
    .Y(_0338_));
 sg13g2_o21ai_1 _0947_ (.B1(_0338_),
    .Y(_0084_),
    .A1(net368),
    .A2(net313));
 sg13g2_nand3_1 _0948_ (.B(net255),
    .C(net314),
    .A(net382),
    .Y(_0339_));
 sg13g2_o21ai_1 _0949_ (.B1(_0339_),
    .Y(_0085_),
    .A1(net370),
    .A2(net314));
 sg13g2_nand3_1 _0950_ (.B(net265),
    .C(net314),
    .A(net380),
    .Y(_0340_));
 sg13g2_o21ai_1 _0951_ (.B1(_0340_),
    .Y(_0086_),
    .A1(net372),
    .A2(net313));
 sg13g2_nand3_1 _0952_ (.B(net194),
    .C(net313),
    .A(net380),
    .Y(_0341_));
 sg13g2_o21ai_1 _0953_ (.B1(_0341_),
    .Y(_0087_),
    .A1(net374),
    .A2(net314));
 sg13g2_nand3_1 _0954_ (.B(_0150_),
    .C(net335),
    .A(net345),
    .Y(_0342_));
 sg13g2_nand3_1 _0955_ (.B(net220),
    .C(net312),
    .A(net392),
    .Y(_0343_));
 sg13g2_o21ai_1 _0956_ (.B1(_0343_),
    .Y(_0088_),
    .A1(net361),
    .A2(net312));
 sg13g2_nand3_1 _0957_ (.B(net167),
    .C(net312),
    .A(net393),
    .Y(_0344_));
 sg13g2_o21ai_1 _0958_ (.B1(_0344_),
    .Y(_0089_),
    .A1(net363),
    .A2(net312));
 sg13g2_nand3_1 _0959_ (.B(net202),
    .C(net312),
    .A(net393),
    .Y(_0345_));
 sg13g2_o21ai_1 _0960_ (.B1(_0345_),
    .Y(_0090_),
    .A1(net365),
    .A2(net312));
 sg13g2_nand3_1 _0961_ (.B(net214),
    .C(net311),
    .A(net390),
    .Y(_0346_));
 sg13g2_o21ai_1 _0962_ (.B1(_0346_),
    .Y(_0091_),
    .A1(net367),
    .A2(net311));
 sg13g2_nand3_1 _0963_ (.B(net201),
    .C(net312),
    .A(net391),
    .Y(_0347_));
 sg13g2_o21ai_1 _0964_ (.B1(_0347_),
    .Y(_0092_),
    .A1(net369),
    .A2(net312));
 sg13g2_nand3_1 _0965_ (.B(net228),
    .C(net311),
    .A(net390),
    .Y(_0348_));
 sg13g2_o21ai_1 _0966_ (.B1(_0348_),
    .Y(_0093_),
    .A1(net370),
    .A2(net311));
 sg13g2_nand3_1 _0967_ (.B(net177),
    .C(net311),
    .A(net389),
    .Y(_0349_));
 sg13g2_o21ai_1 _0968_ (.B1(_0349_),
    .Y(_0094_),
    .A1(net373),
    .A2(net311));
 sg13g2_nand3_1 _0969_ (.B(net166),
    .C(net311),
    .A(net390),
    .Y(_0350_));
 sg13g2_o21ai_1 _0970_ (.B1(_0350_),
    .Y(_0095_),
    .A1(net375),
    .A2(net311));
 sg13g2_nand3_1 _0971_ (.B(_0164_),
    .C(net334),
    .A(net355),
    .Y(_0351_));
 sg13g2_nand3_1 _0972_ (.B(net163),
    .C(net310),
    .A(net386),
    .Y(_0352_));
 sg13g2_o21ai_1 _0973_ (.B1(_0352_),
    .Y(_0096_),
    .A1(net360),
    .A2(_0351_));
 sg13g2_nand3_1 _0974_ (.B(net217),
    .C(net310),
    .A(net386),
    .Y(_0353_));
 sg13g2_o21ai_1 _0975_ (.B1(_0353_),
    .Y(_0097_),
    .A1(net362),
    .A2(net310));
 sg13g2_nand3_1 _0976_ (.B(net210),
    .C(net309),
    .A(net384),
    .Y(_0354_));
 sg13g2_o21ai_1 _0977_ (.B1(_0354_),
    .Y(_0098_),
    .A1(net364),
    .A2(net309));
 sg13g2_nand3_1 _0978_ (.B(net170),
    .C(net309),
    .A(net380),
    .Y(_0355_));
 sg13g2_o21ai_1 _0979_ (.B1(_0355_),
    .Y(_0099_),
    .A1(net366),
    .A2(net309));
 sg13g2_nand3_1 _0980_ (.B(net179),
    .C(net310),
    .A(net388),
    .Y(_0356_));
 sg13g2_o21ai_1 _0981_ (.B1(_0356_),
    .Y(_0100_),
    .A1(net368),
    .A2(net309));
 sg13g2_nand3_1 _0982_ (.B(net222),
    .C(net310),
    .A(net386),
    .Y(_0357_));
 sg13g2_o21ai_1 _0983_ (.B1(_0357_),
    .Y(_0101_),
    .A1(net371),
    .A2(net310));
 sg13g2_nand3_1 _0984_ (.B(net209),
    .C(net310),
    .A(net384),
    .Y(_0358_));
 sg13g2_o21ai_1 _0985_ (.B1(_0358_),
    .Y(_0102_),
    .A1(net372),
    .A2(net309));
 sg13g2_nand3_1 _0986_ (.B(net188),
    .C(net309),
    .A(net385),
    .Y(_0359_));
 sg13g2_o21ai_1 _0987_ (.B1(_0359_),
    .Y(_0103_),
    .A1(net374),
    .A2(net309));
 sg13g2_nand3_1 _0988_ (.B(_0150_),
    .C(net335),
    .A(net339),
    .Y(_0360_));
 sg13g2_nand3_1 _0989_ (.B(net175),
    .C(net308),
    .A(net392),
    .Y(_0361_));
 sg13g2_o21ai_1 _0990_ (.B1(_0361_),
    .Y(_0104_),
    .A1(net361),
    .A2(net308));
 sg13g2_nand3_1 _0991_ (.B(net264),
    .C(net308),
    .A(net393),
    .Y(_0362_));
 sg13g2_o21ai_1 _0992_ (.B1(_0362_),
    .Y(_0105_),
    .A1(net363),
    .A2(net308));
 sg13g2_nand3_1 _0993_ (.B(net267),
    .C(net308),
    .A(net392),
    .Y(_0363_));
 sg13g2_o21ai_1 _0994_ (.B1(_0363_),
    .Y(_0106_),
    .A1(net365),
    .A2(net308));
 sg13g2_nand3_1 _0995_ (.B(net247),
    .C(net307),
    .A(net390),
    .Y(_0364_));
 sg13g2_o21ai_1 _0996_ (.B1(_0364_),
    .Y(_0107_),
    .A1(net367),
    .A2(net307));
 sg13g2_nand3_1 _0997_ (.B(net254),
    .C(net308),
    .A(net392),
    .Y(_0365_));
 sg13g2_o21ai_1 _0998_ (.B1(_0365_),
    .Y(_0108_),
    .A1(net369),
    .A2(net308));
 sg13g2_nand3_1 _0999_ (.B(net203),
    .C(net307),
    .A(net390),
    .Y(_0366_));
 sg13g2_o21ai_1 _1000_ (.B1(_0366_),
    .Y(_0109_),
    .A1(net370),
    .A2(net307));
 sg13g2_nand3_1 _1001_ (.B(net241),
    .C(net307),
    .A(net389),
    .Y(_0367_));
 sg13g2_o21ai_1 _1002_ (.B1(_0367_),
    .Y(_0110_),
    .A1(net373),
    .A2(net307));
 sg13g2_nand3_1 _1003_ (.B(net248),
    .C(net307),
    .A(net390),
    .Y(_0368_));
 sg13g2_o21ai_1 _1004_ (.B1(_0368_),
    .Y(_0111_),
    .A1(net375),
    .A2(net307));
 sg13g2_nand3_1 _1005_ (.B(_0155_),
    .C(net334),
    .A(net344),
    .Y(_0369_));
 sg13g2_nand3_1 _1006_ (.B(net178),
    .C(_0369_),
    .A(net382),
    .Y(_0370_));
 sg13g2_o21ai_1 _1007_ (.B1(_0370_),
    .Y(_0112_),
    .A1(net360),
    .A2(net306));
 sg13g2_nand3_1 _1008_ (.B(net190),
    .C(net306),
    .A(net381),
    .Y(_0371_));
 sg13g2_o21ai_1 _1009_ (.B1(_0371_),
    .Y(_0113_),
    .A1(net362),
    .A2(net306));
 sg13g2_nand3_1 _1010_ (.B(net206),
    .C(net305),
    .A(net379),
    .Y(_0372_));
 sg13g2_o21ai_1 _1011_ (.B1(_0372_),
    .Y(_0114_),
    .A1(net364),
    .A2(net305));
 sg13g2_nand3_1 _1012_ (.B(net186),
    .C(net305),
    .A(net383),
    .Y(_0373_));
 sg13g2_o21ai_1 _1013_ (.B1(_0373_),
    .Y(_0115_),
    .A1(net366),
    .A2(net306));
 sg13g2_nand3_1 _1014_ (.B(net230),
    .C(net305),
    .A(net378),
    .Y(_0374_));
 sg13g2_o21ai_1 _1015_ (.B1(_0374_),
    .Y(_0116_),
    .A1(net368),
    .A2(net305));
 sg13g2_nand3_1 _1016_ (.B(net234),
    .C(net306),
    .A(net382),
    .Y(_0375_));
 sg13g2_o21ai_1 _1017_ (.B1(_0375_),
    .Y(_0117_),
    .A1(net370),
    .A2(net306));
 sg13g2_nand3_1 _1018_ (.B(net168),
    .C(net305),
    .A(net380),
    .Y(_0376_));
 sg13g2_o21ai_1 _1019_ (.B1(_0376_),
    .Y(_0118_),
    .A1(net372),
    .A2(net305));
 sg13g2_nand3_1 _1020_ (.B(net164),
    .C(net305),
    .A(net380),
    .Y(_0377_));
 sg13g2_o21ai_1 _1021_ (.B1(_0377_),
    .Y(_0119_),
    .A1(net374),
    .A2(net306));
 sg13g2_nand3_1 _1022_ (.B(_0150_),
    .C(net335),
    .A(net350),
    .Y(_0378_));
 sg13g2_nand3_1 _1023_ (.B(net278),
    .C(net304),
    .A(net392),
    .Y(_0379_));
 sg13g2_o21ai_1 _1024_ (.B1(_0379_),
    .Y(_0120_),
    .A1(net361),
    .A2(net304));
 sg13g2_nand3_1 _1025_ (.B(net251),
    .C(net304),
    .A(net391),
    .Y(_0380_));
 sg13g2_o21ai_1 _1026_ (.B1(_0380_),
    .Y(_0121_),
    .A1(net363),
    .A2(net304));
 sg13g2_nand3_1 _1027_ (.B(net181),
    .C(net304),
    .A(net391),
    .Y(_0381_));
 sg13g2_o21ai_1 _1028_ (.B1(_0381_),
    .Y(_0122_),
    .A1(net365),
    .A2(net303));
 sg13g2_nand3_1 _1029_ (.B(net213),
    .C(net304),
    .A(net391),
    .Y(_0382_));
 sg13g2_o21ai_1 _1030_ (.B1(_0382_),
    .Y(_0123_),
    .A1(net367),
    .A2(net303));
 sg13g2_nand3_1 _1031_ (.B(net237),
    .C(net304),
    .A(net392),
    .Y(_0383_));
 sg13g2_o21ai_1 _1032_ (.B1(_0383_),
    .Y(_0124_),
    .A1(net369),
    .A2(net304));
 sg13g2_nand3_1 _1033_ (.B(net273),
    .C(net303),
    .A(net389),
    .Y(_0384_));
 sg13g2_o21ai_1 _1034_ (.B1(_0384_),
    .Y(_0125_),
    .A1(net370),
    .A2(net303));
 sg13g2_nand3_1 _1035_ (.B(net233),
    .C(net303),
    .A(net389),
    .Y(_0385_));
 sg13g2_o21ai_1 _1036_ (.B1(_0385_),
    .Y(_0126_),
    .A1(net373),
    .A2(net303));
 sg13g2_nand3_1 _1037_ (.B(net187),
    .C(net303),
    .A(net389),
    .Y(_0386_));
 sg13g2_o21ai_1 _1038_ (.B1(_0386_),
    .Y(_0127_),
    .A1(net375),
    .A2(net303));
 sg13g2_nand3_1 _1039_ (.B(_0150_),
    .C(net335),
    .A(net356),
    .Y(_0387_));
 sg13g2_nand3_1 _1040_ (.B(net235),
    .C(net302),
    .A(net391),
    .Y(_0388_));
 sg13g2_o21ai_1 _1041_ (.B1(_0388_),
    .Y(_0128_),
    .A1(net361),
    .A2(net302));
 sg13g2_nand3_1 _1042_ (.B(net227),
    .C(net302),
    .A(net391),
    .Y(_0389_));
 sg13g2_o21ai_1 _1043_ (.B1(_0389_),
    .Y(_0129_),
    .A1(net363),
    .A2(net302));
 sg13g2_nand3_1 _1044_ (.B(net185),
    .C(net302),
    .A(net391),
    .Y(_0390_));
 sg13g2_o21ai_1 _1045_ (.B1(_0390_),
    .Y(_0130_),
    .A1(net365),
    .A2(net301));
 sg13g2_nand3_1 _1046_ (.B(net193),
    .C(net302),
    .A(net391),
    .Y(_0391_));
 sg13g2_o21ai_1 _1047_ (.B1(_0391_),
    .Y(_0131_),
    .A1(net367),
    .A2(net301));
 sg13g2_nand3_1 _1048_ (.B(net223),
    .C(net302),
    .A(net392),
    .Y(_0392_));
 sg13g2_o21ai_1 _1049_ (.B1(_0392_),
    .Y(_0132_),
    .A1(net369),
    .A2(_0387_));
 sg13g2_nand3_1 _1050_ (.B(net205),
    .C(net301),
    .A(net389),
    .Y(_0393_));
 sg13g2_o21ai_1 _1051_ (.B1(_0393_),
    .Y(_0133_),
    .A1(net370),
    .A2(net301));
 sg13g2_nand3_1 _1052_ (.B(net158),
    .C(net301),
    .A(net389),
    .Y(_0394_));
 sg13g2_o21ai_1 _1053_ (.B1(_0394_),
    .Y(_0134_),
    .A1(net373),
    .A2(net301));
 sg13g2_nand3_1 _1054_ (.B(net197),
    .C(net301),
    .A(net389),
    .Y(_0395_));
 sg13g2_o21ai_1 _1055_ (.B1(_0395_),
    .Y(_0135_),
    .A1(net375),
    .A2(net301));
 sg13g2_buf_1 _1056_ (.A(ui_in[6]),
    .X(_0403_));
 sg13g2_buf_1 _1057_ (.A(ui_in[6]),
    .X(_0402_));
 sg13g2_buf_1 _1058_ (.A(ui_in[6]),
    .X(_0401_));
 sg13g2_buf_1 _1059_ (.A(ui_in[6]),
    .X(_0400_));
 sg13g2_buf_1 _1060_ (.A(ui_in[6]),
    .X(_0399_));
 sg13g2_buf_1 _1061_ (.A(ui_in[6]),
    .X(_0398_));
 sg13g2_buf_1 _1062_ (.A(ui_in[6]),
    .X(_0397_));
 sg13g2_buf_1 _1063_ (.A(ui_in[6]),
    .X(_0396_));
 sg13g2_dfrbp_1 _1064_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net98),
    .D(_0008_),
    .Q_N(_0531_),
    .Q(\RAM[8][0] ));
 sg13g2_dfrbp_1 _1065_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net97),
    .D(_0009_),
    .Q_N(_0530_),
    .Q(\RAM[8][1] ));
 sg13g2_dfrbp_1 _1066_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net95),
    .D(_0010_),
    .Q_N(_0529_),
    .Q(\RAM[8][2] ));
 sg13g2_dfrbp_1 _1067_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net93),
    .D(_0011_),
    .Q_N(_0528_),
    .Q(\RAM[8][3] ));
 sg13g2_dfrbp_1 _1068_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net91),
    .D(_0012_),
    .Q_N(_0527_),
    .Q(\RAM[8][4] ));
 sg13g2_dfrbp_1 _1069_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net89),
    .D(_0013_),
    .Q_N(_0526_),
    .Q(\RAM[8][5] ));
 sg13g2_dfrbp_1 _1070_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net87),
    .D(_0014_),
    .Q_N(_0525_),
    .Q(\RAM[8][6] ));
 sg13g2_dfrbp_1 _1071_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net85),
    .D(_0015_),
    .Q_N(_0524_),
    .Q(\RAM[8][7] ));
 sg13g2_dfrbp_1 _1072_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net83),
    .D(_0016_),
    .Q_N(_0523_),
    .Q(\RAM[15][0] ));
 sg13g2_dfrbp_1 _1073_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net81),
    .D(_0017_),
    .Q_N(_0522_),
    .Q(\RAM[15][1] ));
 sg13g2_dfrbp_1 _1074_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net79),
    .D(_0018_),
    .Q_N(_0521_),
    .Q(\RAM[15][2] ));
 sg13g2_dfrbp_1 _1075_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net77),
    .D(_0019_),
    .Q_N(_0520_),
    .Q(\RAM[15][3] ));
 sg13g2_dfrbp_1 _1076_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net75),
    .D(_0020_),
    .Q_N(_0519_),
    .Q(\RAM[15][4] ));
 sg13g2_dfrbp_1 _1077_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net73),
    .D(_0021_),
    .Q_N(_0518_),
    .Q(\RAM[15][5] ));
 sg13g2_dfrbp_1 _1078_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net71),
    .D(_0022_),
    .Q_N(_0517_),
    .Q(\RAM[15][6] ));
 sg13g2_dfrbp_1 _1079_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net69),
    .D(_0023_),
    .Q_N(_0516_),
    .Q(\RAM[15][7] ));
 sg13g2_dfrbp_1 _1080_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net67),
    .D(_0024_),
    .Q_N(_0515_),
    .Q(\RAM[12][0] ));
 sg13g2_dfrbp_1 _1081_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net65),
    .D(_0025_),
    .Q_N(_0514_),
    .Q(\RAM[12][1] ));
 sg13g2_dfrbp_1 _1082_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net63),
    .D(_0026_),
    .Q_N(_0513_),
    .Q(\RAM[12][2] ));
 sg13g2_dfrbp_1 _1083_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net61),
    .D(_0027_),
    .Q_N(_0512_),
    .Q(\RAM[12][3] ));
 sg13g2_dfrbp_1 _1084_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net59),
    .D(_0028_),
    .Q_N(_0511_),
    .Q(\RAM[12][4] ));
 sg13g2_dfrbp_1 _1085_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net57),
    .D(_0029_),
    .Q_N(_0510_),
    .Q(\RAM[12][5] ));
 sg13g2_dfrbp_1 _1086_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net55),
    .D(_0030_),
    .Q_N(_0509_),
    .Q(\RAM[12][6] ));
 sg13g2_dfrbp_1 _1087_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net53),
    .D(_0031_),
    .Q_N(_0508_),
    .Q(\RAM[12][7] ));
 sg13g2_dfrbp_1 _1088_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net51),
    .D(_0032_),
    .Q_N(_0507_),
    .Q(\RAM[13][0] ));
 sg13g2_dfrbp_1 _1089_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net49),
    .D(_0033_),
    .Q_N(_0506_),
    .Q(\RAM[13][1] ));
 sg13g2_dfrbp_1 _1090_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net47),
    .D(_0034_),
    .Q_N(_0505_),
    .Q(\RAM[13][2] ));
 sg13g2_dfrbp_1 _1091_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net45),
    .D(_0035_),
    .Q_N(_0504_),
    .Q(\RAM[13][3] ));
 sg13g2_dfrbp_1 _1092_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net43),
    .D(_0036_),
    .Q_N(_0503_),
    .Q(\RAM[13][4] ));
 sg13g2_dfrbp_1 _1093_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net41),
    .D(_0037_),
    .Q_N(_0502_),
    .Q(\RAM[13][5] ));
 sg13g2_dfrbp_1 _1094_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net39),
    .D(_0038_),
    .Q_N(_0501_),
    .Q(\RAM[13][6] ));
 sg13g2_dfrbp_1 _1095_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net37),
    .D(_0039_),
    .Q_N(_0500_),
    .Q(\RAM[13][7] ));
 sg13g2_dfrbp_1 _1096_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net35),
    .D(_0040_),
    .Q_N(_0499_),
    .Q(\RAM[0][0] ));
 sg13g2_dfrbp_1 _1097_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net33),
    .D(_0041_),
    .Q_N(_0498_),
    .Q(\RAM[0][1] ));
 sg13g2_dfrbp_1 _1098_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net31),
    .D(_0042_),
    .Q_N(_0497_),
    .Q(\RAM[0][2] ));
 sg13g2_dfrbp_1 _1099_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net157),
    .D(_0043_),
    .Q_N(_0496_),
    .Q(\RAM[0][3] ));
 sg13g2_dfrbp_1 _1100_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net155),
    .D(_0044_),
    .Q_N(_0495_),
    .Q(\RAM[0][4] ));
 sg13g2_dfrbp_1 _1101_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net153),
    .D(_0045_),
    .Q_N(_0494_),
    .Q(\RAM[0][5] ));
 sg13g2_dfrbp_1 _1102_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net151),
    .D(_0046_),
    .Q_N(_0493_),
    .Q(\RAM[0][6] ));
 sg13g2_dfrbp_1 _1103_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net149),
    .D(_0047_),
    .Q_N(_0492_),
    .Q(\RAM[0][7] ));
 sg13g2_dfrbp_1 _1104_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net147),
    .D(_0048_),
    .Q_N(_0491_),
    .Q(\RAM[10][0] ));
 sg13g2_dfrbp_1 _1105_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net145),
    .D(_0049_),
    .Q_N(_0490_),
    .Q(\RAM[10][1] ));
 sg13g2_dfrbp_1 _1106_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net143),
    .D(_0050_),
    .Q_N(_0489_),
    .Q(\RAM[10][2] ));
 sg13g2_dfrbp_1 _1107_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net141),
    .D(_0051_),
    .Q_N(_0488_),
    .Q(\RAM[10][3] ));
 sg13g2_dfrbp_1 _1108_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net139),
    .D(_0052_),
    .Q_N(_0487_),
    .Q(\RAM[10][4] ));
 sg13g2_dfrbp_1 _1109_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net137),
    .D(_0053_),
    .Q_N(_0486_),
    .Q(\RAM[10][5] ));
 sg13g2_dfrbp_1 _1110_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net135),
    .D(_0054_),
    .Q_N(_0485_),
    .Q(\RAM[10][6] ));
 sg13g2_dfrbp_1 _1111_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net133),
    .D(_0055_),
    .Q_N(_0484_),
    .Q(\RAM[10][7] ));
 sg13g2_dfrbp_1 _1112_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net131),
    .D(_0056_),
    .Q_N(_0483_),
    .Q(\RAM[11][0] ));
 sg13g2_dfrbp_1 _1113_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net129),
    .D(_0057_),
    .Q_N(_0482_),
    .Q(\RAM[11][1] ));
 sg13g2_dfrbp_1 _1114_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net127),
    .D(_0058_),
    .Q_N(_0481_),
    .Q(\RAM[11][2] ));
 sg13g2_dfrbp_1 _1115_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net125),
    .D(_0059_),
    .Q_N(_0480_),
    .Q(\RAM[11][3] ));
 sg13g2_dfrbp_1 _1116_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net123),
    .D(_0060_),
    .Q_N(_0479_),
    .Q(\RAM[11][4] ));
 sg13g2_dfrbp_1 _1117_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net121),
    .D(_0061_),
    .Q_N(_0478_),
    .Q(\RAM[11][5] ));
 sg13g2_dfrbp_1 _1118_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net119),
    .D(_0062_),
    .Q_N(_0477_),
    .Q(\RAM[11][6] ));
 sg13g2_dfrbp_1 _1119_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net117),
    .D(_0063_),
    .Q_N(_0476_),
    .Q(\RAM[11][7] ));
 sg13g2_dfrbp_1 _1120_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net115),
    .D(_0064_),
    .Q_N(_0475_),
    .Q(\RAM[1][0] ));
 sg13g2_dfrbp_1 _1121_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net113),
    .D(_0065_),
    .Q_N(_0474_),
    .Q(\RAM[1][1] ));
 sg13g2_dfrbp_1 _1122_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net111),
    .D(_0066_),
    .Q_N(_0473_),
    .Q(\RAM[1][2] ));
 sg13g2_dfrbp_1 _1123_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net109),
    .D(_0067_),
    .Q_N(_0472_),
    .Q(\RAM[1][3] ));
 sg13g2_dfrbp_1 _1124_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net107),
    .D(_0068_),
    .Q_N(_0471_),
    .Q(\RAM[1][4] ));
 sg13g2_dfrbp_1 _1125_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net105),
    .D(_0069_),
    .Q_N(_0470_),
    .Q(\RAM[1][5] ));
 sg13g2_dfrbp_1 _1126_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net103),
    .D(_0070_),
    .Q_N(_0469_),
    .Q(\RAM[1][6] ));
 sg13g2_dfrbp_1 _1127_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net101),
    .D(_0071_),
    .Q_N(_0468_),
    .Q(\RAM[1][7] ));
 sg13g2_dfrbp_1 _1128_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net99),
    .D(_0072_),
    .Q_N(_0467_),
    .Q(\RAM[14][0] ));
 sg13g2_dfrbp_1 _1129_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net96),
    .D(_0073_),
    .Q_N(_0466_),
    .Q(\RAM[14][1] ));
 sg13g2_dfrbp_1 _1130_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net92),
    .D(_0074_),
    .Q_N(_0465_),
    .Q(\RAM[14][2] ));
 sg13g2_dfrbp_1 _1131_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net88),
    .D(_0075_),
    .Q_N(_0464_),
    .Q(\RAM[14][3] ));
 sg13g2_dfrbp_1 _1132_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net84),
    .D(_0076_),
    .Q_N(_0463_),
    .Q(\RAM[14][4] ));
 sg13g2_dfrbp_1 _1133_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net80),
    .D(_0077_),
    .Q_N(_0462_),
    .Q(\RAM[14][5] ));
 sg13g2_dfrbp_1 _1134_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net76),
    .D(_0078_),
    .Q_N(_0461_),
    .Q(\RAM[14][6] ));
 sg13g2_dfrbp_1 _1135_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net72),
    .D(_0079_),
    .Q_N(_0460_),
    .Q(\RAM[14][7] ));
 sg13g2_dfrbp_1 _1136_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net68),
    .D(_0080_),
    .Q_N(_0459_),
    .Q(\RAM[2][0] ));
 sg13g2_dfrbp_1 _1137_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net64),
    .D(_0081_),
    .Q_N(_0458_),
    .Q(\RAM[2][1] ));
 sg13g2_dfrbp_1 _1138_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net60),
    .D(_0082_),
    .Q_N(_0457_),
    .Q(\RAM[2][2] ));
 sg13g2_dfrbp_1 _1139_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net56),
    .D(_0083_),
    .Q_N(_0456_),
    .Q(\RAM[2][3] ));
 sg13g2_dfrbp_1 _1140_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net52),
    .D(_0084_),
    .Q_N(_0455_),
    .Q(\RAM[2][4] ));
 sg13g2_dfrbp_1 _1141_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net48),
    .D(_0085_),
    .Q_N(_0454_),
    .Q(\RAM[2][5] ));
 sg13g2_dfrbp_1 _1142_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net44),
    .D(_0086_),
    .Q_N(_0453_),
    .Q(\RAM[2][6] ));
 sg13g2_dfrbp_1 _1143_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net40),
    .D(_0087_),
    .Q_N(_0452_),
    .Q(\RAM[2][7] ));
 sg13g2_dfrbp_1 _1144_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net36),
    .D(_0088_),
    .Q_N(_0451_),
    .Q(\RAM[7][0] ));
 sg13g2_dfrbp_1 _1145_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net32),
    .D(_0089_),
    .Q_N(_0450_),
    .Q(\RAM[7][1] ));
 sg13g2_dfrbp_1 _1146_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net156),
    .D(_0090_),
    .Q_N(_0449_),
    .Q(\RAM[7][2] ));
 sg13g2_dfrbp_1 _1147_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net152),
    .D(_0091_),
    .Q_N(_0448_),
    .Q(\RAM[7][3] ));
 sg13g2_dfrbp_1 _1148_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net148),
    .D(_0092_),
    .Q_N(_0447_),
    .Q(\RAM[7][4] ));
 sg13g2_dfrbp_1 _1149_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net144),
    .D(_0093_),
    .Q_N(_0446_),
    .Q(\RAM[7][5] ));
 sg13g2_dfrbp_1 _1150_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net140),
    .D(_0094_),
    .Q_N(_0445_),
    .Q(\RAM[7][6] ));
 sg13g2_dfrbp_1 _1151_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net136),
    .D(_0095_),
    .Q_N(_0444_),
    .Q(\RAM[7][7] ));
 sg13g2_dfrbp_1 _1152_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net132),
    .D(_0096_),
    .Q_N(_0443_),
    .Q(\RAM[9][0] ));
 sg13g2_dfrbp_1 _1153_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net128),
    .D(_0097_),
    .Q_N(_0442_),
    .Q(\RAM[9][1] ));
 sg13g2_dfrbp_1 _1154_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net124),
    .D(_0098_),
    .Q_N(_0441_),
    .Q(\RAM[9][2] ));
 sg13g2_dfrbp_1 _1155_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net120),
    .D(_0099_),
    .Q_N(_0440_),
    .Q(\RAM[9][3] ));
 sg13g2_dfrbp_1 _1156_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net116),
    .D(_0100_),
    .Q_N(_0439_),
    .Q(\RAM[9][4] ));
 sg13g2_dfrbp_1 _1157_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net112),
    .D(_0101_),
    .Q_N(_0438_),
    .Q(\RAM[9][5] ));
 sg13g2_dfrbp_1 _1158_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net108),
    .D(_0102_),
    .Q_N(_0437_),
    .Q(\RAM[9][6] ));
 sg13g2_dfrbp_1 _1159_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net104),
    .D(_0103_),
    .Q_N(_0436_),
    .Q(\RAM[9][7] ));
 sg13g2_dfrbp_1 _1160_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net100),
    .D(_0104_),
    .Q_N(_0435_),
    .Q(\RAM[6][0] ));
 sg13g2_dfrbp_1 _1161_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net94),
    .D(_0105_),
    .Q_N(_0434_),
    .Q(\RAM[6][1] ));
 sg13g2_dfrbp_1 _1162_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net86),
    .D(_0106_),
    .Q_N(_0433_),
    .Q(\RAM[6][2] ));
 sg13g2_dfrbp_1 _1163_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net78),
    .D(_0107_),
    .Q_N(_0432_),
    .Q(\RAM[6][3] ));
 sg13g2_dfrbp_1 _1164_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net70),
    .D(_0108_),
    .Q_N(_0431_),
    .Q(\RAM[6][4] ));
 sg13g2_dfrbp_1 _1165_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net62),
    .D(_0109_),
    .Q_N(_0430_),
    .Q(\RAM[6][5] ));
 sg13g2_dfrbp_1 _1166_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net54),
    .D(_0110_),
    .Q_N(_0429_),
    .Q(\RAM[6][6] ));
 sg13g2_dfrbp_1 _1167_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net46),
    .D(_0111_),
    .Q_N(_0428_),
    .Q(\RAM[6][7] ));
 sg13g2_dfrbp_1 _1168_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net38),
    .D(_0112_),
    .Q_N(_0427_),
    .Q(\RAM[3][0] ));
 sg13g2_dfrbp_1 _1169_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net30),
    .D(_0113_),
    .Q_N(_0426_),
    .Q(\RAM[3][1] ));
 sg13g2_dfrbp_1 _1170_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net150),
    .D(_0114_),
    .Q_N(_0425_),
    .Q(\RAM[3][2] ));
 sg13g2_dfrbp_1 _1171_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net142),
    .D(_0115_),
    .Q_N(_0424_),
    .Q(\RAM[3][3] ));
 sg13g2_dfrbp_1 _1172_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net134),
    .D(_0116_),
    .Q_N(_0423_),
    .Q(\RAM[3][4] ));
 sg13g2_dfrbp_1 _1173_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net126),
    .D(_0117_),
    .Q_N(_0422_),
    .Q(\RAM[3][5] ));
 sg13g2_dfrbp_1 _1174_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net118),
    .D(_0118_),
    .Q_N(_0421_),
    .Q(\RAM[3][6] ));
 sg13g2_dfrbp_1 _1175_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net110),
    .D(_0119_),
    .Q_N(_0420_),
    .Q(\RAM[3][7] ));
 sg13g2_dfrbp_1 _1176_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net102),
    .D(_0120_),
    .Q_N(_0419_),
    .Q(\RAM[4][0] ));
 sg13g2_dfrbp_1 _1177_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net90),
    .D(_0121_),
    .Q_N(_0418_),
    .Q(\RAM[4][1] ));
 sg13g2_dfrbp_1 _1178_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net74),
    .D(_0122_),
    .Q_N(_0417_),
    .Q(\RAM[4][2] ));
 sg13g2_dfrbp_1 _1179_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net58),
    .D(_0123_),
    .Q_N(_0416_),
    .Q(\RAM[4][3] ));
 sg13g2_dfrbp_1 _1180_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net42),
    .D(_0124_),
    .Q_N(_0415_),
    .Q(\RAM[4][4] ));
 sg13g2_dfrbp_1 _1181_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net154),
    .D(_0125_),
    .Q_N(_0414_),
    .Q(\RAM[4][5] ));
 sg13g2_dfrbp_1 _1182_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net138),
    .D(_0126_),
    .Q_N(_0413_),
    .Q(\RAM[4][6] ));
 sg13g2_dfrbp_1 _1183_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net122),
    .D(_0127_),
    .Q_N(_0412_),
    .Q(\RAM[4][7] ));
 sg13g2_dfrbp_1 _1184_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net106),
    .D(_0128_),
    .Q_N(_0411_),
    .Q(\RAM[5][0] ));
 sg13g2_dfrbp_1 _1185_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net82),
    .D(_0129_),
    .Q_N(_0410_),
    .Q(\RAM[5][1] ));
 sg13g2_dfrbp_1 _1186_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net50),
    .D(_0130_),
    .Q_N(_0409_),
    .Q(\RAM[5][2] ));
 sg13g2_dfrbp_1 _1187_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net146),
    .D(_0131_),
    .Q_N(_0408_),
    .Q(\RAM[5][3] ));
 sg13g2_dfrbp_1 _1188_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net114),
    .D(_0132_),
    .Q_N(_0407_),
    .Q(\RAM[5][4] ));
 sg13g2_dfrbp_1 _1189_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net66),
    .D(_0133_),
    .Q_N(_0406_),
    .Q(\RAM[5][5] ));
 sg13g2_dfrbp_1 _1190_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net130),
    .D(_0134_),
    .Q_N(_0405_),
    .Q(\RAM[5][6] ));
 sg13g2_dfrbp_1 _1191_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net34),
    .D(_0135_),
    .Q_N(_0404_),
    .Q(\RAM[5][7] ));
 sg13g2_tiehi _1098__31 (.L_HI(net31));
 sg13g2_tiehi _1145__32 (.L_HI(net32));
 sg13g2_tiehi _1097__33 (.L_HI(net33));
 sg13g2_tiehi _1191__34 (.L_HI(net34));
 sg13g2_tiehi _1096__35 (.L_HI(net35));
 sg13g2_tiehi _1144__36 (.L_HI(net36));
 sg13g2_tiehi _1095__37 (.L_HI(net37));
 sg13g2_tiehi _1168__38 (.L_HI(net38));
 sg13g2_tiehi _1094__39 (.L_HI(net39));
 sg13g2_tiehi _1143__40 (.L_HI(net40));
 sg13g2_tiehi _1093__41 (.L_HI(net41));
 sg13g2_tiehi _1180__42 (.L_HI(net42));
 sg13g2_tiehi _1092__43 (.L_HI(net43));
 sg13g2_tiehi _1142__44 (.L_HI(net44));
 sg13g2_tiehi _1091__45 (.L_HI(net45));
 sg13g2_tiehi _1167__46 (.L_HI(net46));
 sg13g2_tiehi _1090__47 (.L_HI(net47));
 sg13g2_tiehi _1141__48 (.L_HI(net48));
 sg13g2_tiehi _1089__49 (.L_HI(net49));
 sg13g2_tiehi _1186__50 (.L_HI(net50));
 sg13g2_tiehi _1088__51 (.L_HI(net51));
 sg13g2_tiehi _1140__52 (.L_HI(net52));
 sg13g2_tiehi _1087__53 (.L_HI(net53));
 sg13g2_tiehi _1166__54 (.L_HI(net54));
 sg13g2_tiehi _1086__55 (.L_HI(net55));
 sg13g2_tiehi _1139__56 (.L_HI(net56));
 sg13g2_tiehi _1085__57 (.L_HI(net57));
 sg13g2_tiehi _1179__58 (.L_HI(net58));
 sg13g2_tiehi _1084__59 (.L_HI(net59));
 sg13g2_tiehi _1138__60 (.L_HI(net60));
 sg13g2_tiehi _1083__61 (.L_HI(net61));
 sg13g2_tiehi _1165__62 (.L_HI(net62));
 sg13g2_tiehi _1082__63 (.L_HI(net63));
 sg13g2_tiehi _1137__64 (.L_HI(net64));
 sg13g2_tiehi _1081__65 (.L_HI(net65));
 sg13g2_tiehi _1189__66 (.L_HI(net66));
 sg13g2_tiehi _1080__67 (.L_HI(net67));
 sg13g2_tiehi _1136__68 (.L_HI(net68));
 sg13g2_tiehi _1079__69 (.L_HI(net69));
 sg13g2_tiehi _1164__70 (.L_HI(net70));
 sg13g2_tiehi _1078__71 (.L_HI(net71));
 sg13g2_tiehi _1135__72 (.L_HI(net72));
 sg13g2_tiehi _1077__73 (.L_HI(net73));
 sg13g2_tiehi _1178__74 (.L_HI(net74));
 sg13g2_tiehi _1076__75 (.L_HI(net75));
 sg13g2_tiehi _1134__76 (.L_HI(net76));
 sg13g2_tiehi _1075__77 (.L_HI(net77));
 sg13g2_tiehi _1163__78 (.L_HI(net78));
 sg13g2_tiehi _1074__79 (.L_HI(net79));
 sg13g2_tiehi _1133__80 (.L_HI(net80));
 sg13g2_tiehi _1073__81 (.L_HI(net81));
 sg13g2_tiehi _1185__82 (.L_HI(net82));
 sg13g2_tiehi _1072__83 (.L_HI(net83));
 sg13g2_tiehi _1132__84 (.L_HI(net84));
 sg13g2_tiehi _1071__85 (.L_HI(net85));
 sg13g2_tiehi _1162__86 (.L_HI(net86));
 sg13g2_tiehi _1070__87 (.L_HI(net87));
 sg13g2_tiehi _1131__88 (.L_HI(net88));
 sg13g2_tiehi _1069__89 (.L_HI(net89));
 sg13g2_tiehi _1177__90 (.L_HI(net90));
 sg13g2_tiehi _1068__91 (.L_HI(net91));
 sg13g2_tiehi _1130__92 (.L_HI(net92));
 sg13g2_tiehi _1067__93 (.L_HI(net93));
 sg13g2_tiehi _1161__94 (.L_HI(net94));
 sg13g2_tiehi _1066__95 (.L_HI(net95));
 sg13g2_tiehi _1129__96 (.L_HI(net96));
 sg13g2_tiehi _1065__97 (.L_HI(net97));
 sg13g2_tiehi _1064__98 (.L_HI(net98));
 sg13g2_tiehi _1128__99 (.L_HI(net99));
 sg13g2_tiehi _1160__100 (.L_HI(net100));
 sg13g2_tiehi _1127__101 (.L_HI(net101));
 sg13g2_tiehi _1176__102 (.L_HI(net102));
 sg13g2_tiehi _1126__103 (.L_HI(net103));
 sg13g2_tiehi _1159__104 (.L_HI(net104));
 sg13g2_tiehi _1125__105 (.L_HI(net105));
 sg13g2_tiehi _1184__106 (.L_HI(net106));
 sg13g2_tiehi _1124__107 (.L_HI(net107));
 sg13g2_tiehi _1158__108 (.L_HI(net108));
 sg13g2_tiehi _1123__109 (.L_HI(net109));
 sg13g2_tiehi _1175__110 (.L_HI(net110));
 sg13g2_tiehi _1122__111 (.L_HI(net111));
 sg13g2_tiehi _1157__112 (.L_HI(net112));
 sg13g2_tiehi _1121__113 (.L_HI(net113));
 sg13g2_tiehi _1188__114 (.L_HI(net114));
 sg13g2_tiehi _1120__115 (.L_HI(net115));
 sg13g2_tiehi _1156__116 (.L_HI(net116));
 sg13g2_tiehi _1119__117 (.L_HI(net117));
 sg13g2_tiehi _1174__118 (.L_HI(net118));
 sg13g2_tiehi _1118__119 (.L_HI(net119));
 sg13g2_tiehi _1155__120 (.L_HI(net120));
 sg13g2_tiehi _1117__121 (.L_HI(net121));
 sg13g2_tiehi _1183__122 (.L_HI(net122));
 sg13g2_tiehi _1116__123 (.L_HI(net123));
 sg13g2_tiehi _1154__124 (.L_HI(net124));
 sg13g2_tiehi _1115__125 (.L_HI(net125));
 sg13g2_tiehi _1173__126 (.L_HI(net126));
 sg13g2_tiehi _1114__127 (.L_HI(net127));
 sg13g2_tiehi _1153__128 (.L_HI(net128));
 sg13g2_tiehi _1113__129 (.L_HI(net129));
 sg13g2_tiehi _1190__130 (.L_HI(net130));
 sg13g2_tiehi _1112__131 (.L_HI(net131));
 sg13g2_tiehi _1152__132 (.L_HI(net132));
 sg13g2_tiehi _1111__133 (.L_HI(net133));
 sg13g2_tiehi _1172__134 (.L_HI(net134));
 sg13g2_tiehi _1110__135 (.L_HI(net135));
 sg13g2_tiehi _1151__136 (.L_HI(net136));
 sg13g2_tiehi _1109__137 (.L_HI(net137));
 sg13g2_tiehi _1182__138 (.L_HI(net138));
 sg13g2_tiehi _1108__139 (.L_HI(net139));
 sg13g2_tiehi _1150__140 (.L_HI(net140));
 sg13g2_tiehi _1107__141 (.L_HI(net141));
 sg13g2_tiehi _1171__142 (.L_HI(net142));
 sg13g2_tiehi _1106__143 (.L_HI(net143));
 sg13g2_tiehi _1149__144 (.L_HI(net144));
 sg13g2_tiehi _1105__145 (.L_HI(net145));
 sg13g2_tiehi _1187__146 (.L_HI(net146));
 sg13g2_tiehi _1104__147 (.L_HI(net147));
 sg13g2_tiehi _1148__148 (.L_HI(net148));
 sg13g2_tiehi _1103__149 (.L_HI(net149));
 sg13g2_tiehi _1170__150 (.L_HI(net150));
 sg13g2_tiehi _1102__151 (.L_HI(net151));
 sg13g2_tiehi _1147__152 (.L_HI(net152));
 sg13g2_tiehi _1101__153 (.L_HI(net153));
 sg13g2_tiehi _1181__154 (.L_HI(net154));
 sg13g2_tiehi _1100__155 (.L_HI(net155));
 sg13g2_tiehi _1146__156 (.L_HI(net156));
 sg13g2_tiehi _1099__157 (.L_HI(net157));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_dff_mem_15 (.L_LO(net15));
 sg13g2_tielo tt_um_dff_mem_16 (.L_LO(net16));
 sg13g2_tielo tt_um_dff_mem_17 (.L_LO(net17));
 sg13g2_tielo tt_um_dff_mem_18 (.L_LO(net18));
 sg13g2_tielo tt_um_dff_mem_19 (.L_LO(net19));
 sg13g2_tielo tt_um_dff_mem_20 (.L_LO(net20));
 sg13g2_tielo tt_um_dff_mem_21 (.L_LO(net21));
 sg13g2_tielo tt_um_dff_mem_22 (.L_LO(net22));
 sg13g2_tielo tt_um_dff_mem_23 (.L_LO(net23));
 sg13g2_tielo tt_um_dff_mem_24 (.L_LO(net24));
 sg13g2_tielo tt_um_dff_mem_25 (.L_LO(net25));
 sg13g2_tielo tt_um_dff_mem_26 (.L_LO(net26));
 sg13g2_tielo tt_um_dff_mem_27 (.L_LO(net27));
 sg13g2_tielo tt_um_dff_mem_28 (.L_LO(net28));
 sg13g2_tielo tt_um_dff_mem_29 (.L_LO(net29));
 sg13g2_tiehi _1169__30 (.L_HI(net30));
 sg13g2_ebufn_2 _1336_ (.TE_B(_0396_),
    .A(_0000_),
    .Z(uo_out[0]));
 sg13g2_ebufn_4 _1337_ (.A(_0001_),
    .TE_B(_0397_),
    .Z(uo_out[1]));
 sg13g2_ebufn_4 _1338_ (.A(_0002_),
    .TE_B(_0398_),
    .Z(uo_out[2]));
 sg13g2_ebufn_2 _1339_ (.TE_B(_0399_),
    .A(_0003_),
    .Z(uo_out[3]));
 sg13g2_ebufn_2 _1340_ (.TE_B(_0400_),
    .A(_0004_),
    .Z(uo_out[4]));
 sg13g2_ebufn_2 _1341_ (.TE_B(_0401_),
    .A(_0005_),
    .Z(uo_out[5]));
 sg13g2_ebufn_2 _1342_ (.TE_B(_0402_),
    .A(_0006_),
    .Z(uo_out[6]));
 sg13g2_ebufn_2 _1343_ (.TE_B(_0403_),
    .A(_0007_),
    .Z(uo_out[7]));
 sg13g2_buf_2 fanout301 (.A(net302),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_0387_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_0378_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_0378_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(net306),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_0369_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_0360_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_0360_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(net310),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_0351_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_0342_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_0342_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(net314),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_0333_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_0324_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_0324_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(net318),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_0315_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(net320),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_0306_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(net323),
    .X(net321));
 sg13g2_buf_1 fanout322 (.A(net323),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_0297_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(net325),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_0288_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(net327),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_0279_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_0270_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_0270_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(net331),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_0261_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(net333),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_0252_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_0251_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_0251_),
    .X(net335));
 sg13g2_buf_4 fanout336 (.X(net336),
    .A(net338));
 sg13g2_buf_2 fanout337 (.A(net338),
    .X(net337));
 sg13g2_buf_4 fanout338 (.X(net338),
    .A(net341));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(net340));
 sg13g2_buf_4 fanout340 (.X(net340),
    .A(net341));
 sg13g2_buf_2 fanout341 (.A(_0148_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(net344),
    .X(net342));
 sg13g2_buf_1 fanout343 (.A(net344),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(net347),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(net346),
    .X(net345));
 sg13g2_buf_4 fanout346 (.X(net346),
    .A(net347));
 sg13g2_buf_2 fanout347 (.A(_0147_),
    .X(net347));
 sg13g2_buf_4 fanout348 (.X(net348),
    .A(net349));
 sg13g2_buf_4 fanout349 (.X(net349),
    .A(net353));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(net352));
 sg13g2_buf_2 fanout351 (.A(net352),
    .X(net351));
 sg13g2_buf_4 fanout352 (.X(net352),
    .A(net353));
 sg13g2_buf_2 fanout353 (.A(_0145_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(net355),
    .X(net354));
 sg13g2_buf_4 fanout355 (.X(net355),
    .A(net359));
 sg13g2_buf_2 fanout356 (.A(net358),
    .X(net356));
 sg13g2_buf_1 fanout357 (.A(net358),
    .X(net357));
 sg13g2_buf_4 fanout358 (.X(net358),
    .A(net359));
 sg13g2_buf_2 fanout359 (.A(_0144_),
    .X(net359));
 sg13g2_buf_4 fanout360 (.X(net360),
    .A(_0143_));
 sg13g2_buf_4 fanout361 (.X(net361),
    .A(_0143_));
 sg13g2_buf_4 fanout362 (.X(net362),
    .A(_0142_));
 sg13g2_buf_4 fanout363 (.X(net363),
    .A(_0142_));
 sg13g2_buf_4 fanout364 (.X(net364),
    .A(_0141_));
 sg13g2_buf_4 fanout365 (.X(net365),
    .A(_0141_));
 sg13g2_buf_4 fanout366 (.X(net366),
    .A(_0140_));
 sg13g2_buf_4 fanout367 (.X(net367),
    .A(_0140_));
 sg13g2_buf_4 fanout368 (.X(net368),
    .A(_0139_));
 sg13g2_buf_4 fanout369 (.X(net369),
    .A(_0139_));
 sg13g2_buf_4 fanout370 (.X(net370),
    .A(_0138_));
 sg13g2_buf_4 fanout371 (.X(net371),
    .A(_0138_));
 sg13g2_buf_4 fanout372 (.X(net372),
    .A(_0137_));
 sg13g2_buf_4 fanout373 (.X(net373),
    .A(_0137_));
 sg13g2_buf_4 fanout374 (.X(net374),
    .A(_0136_));
 sg13g2_buf_4 fanout375 (.X(net375),
    .A(_0136_));
 sg13g2_buf_4 fanout376 (.X(net376),
    .A(net4));
 sg13g2_buf_4 fanout377 (.X(net377),
    .A(net3));
 sg13g2_buf_2 fanout378 (.A(net380),
    .X(net378));
 sg13g2_buf_1 fanout379 (.A(net380),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(net383),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(net383),
    .X(net381));
 sg13g2_buf_1 fanout382 (.A(net383),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(rst_n),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(net385),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(net388),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(net388),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(net388),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(rst_n),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(net393),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(net393),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(net392),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(net393),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(net399),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(net399),
    .X(net394));
 sg13g2_buf_1 fanout395 (.A(net399),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(net398),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(net398),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(net399),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(rst_n),
    .X(net399));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[7]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[0]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[1]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[2]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[4]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[5]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[6]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[7]),
    .X(net13));
 sg13g2_tielo tt_um_dff_mem_14 (.L_LO(net14));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\RAM[5][6] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold2 (.A(\RAM[15][2] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold3 (.A(\RAM[8][2] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold4 (.A(\RAM[13][3] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold5 (.A(\RAM[1][7] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold6 (.A(\RAM[9][0] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold7 (.A(\RAM[3][7] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold8 (.A(\RAM[11][1] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold9 (.A(\RAM[7][7] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold10 (.A(\RAM[7][1] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold11 (.A(\RAM[3][6] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold12 (.A(\RAM[13][4] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold13 (.A(\RAM[9][3] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold14 (.A(\RAM[13][7] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold15 (.A(\RAM[0][1] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold16 (.A(\RAM[13][6] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold17 (.A(\RAM[10][3] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold18 (.A(\RAM[6][0] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold19 (.A(\RAM[12][2] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold20 (.A(\RAM[7][6] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold21 (.A(\RAM[3][0] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold22 (.A(\RAM[9][4] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold23 (.A(\RAM[15][7] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold24 (.A(\RAM[4][2] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold25 (.A(\RAM[13][1] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold26 (.A(\RAM[11][2] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold27 (.A(\RAM[15][1] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold28 (.A(\RAM[5][2] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold29 (.A(\RAM[3][3] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold30 (.A(\RAM[4][7] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold31 (.A(\RAM[9][7] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold32 (.A(\RAM[0][7] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold33 (.A(\RAM[3][1] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold34 (.A(\RAM[0][0] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold35 (.A(\RAM[14][2] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold36 (.A(\RAM[5][3] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold37 (.A(\RAM[2][7] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold38 (.A(\RAM[14][3] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold39 (.A(\RAM[10][5] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold40 (.A(\RAM[5][7] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold41 (.A(\RAM[12][1] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold42 (.A(\RAM[14][7] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold43 (.A(\RAM[1][2] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold44 (.A(\RAM[7][4] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold45 (.A(\RAM[7][2] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold46 (.A(\RAM[6][5] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold47 (.A(\RAM[1][5] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold48 (.A(\RAM[5][5] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold49 (.A(\RAM[3][2] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold50 (.A(\RAM[0][5] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold51 (.A(\RAM[13][0] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold52 (.A(\RAM[9][6] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold53 (.A(\RAM[9][2] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold54 (.A(\RAM[15][3] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold55 (.A(\RAM[14][6] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold56 (.A(\RAM[4][3] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold57 (.A(\RAM[7][3] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold58 (.A(\RAM[11][3] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold59 (.A(\RAM[11][5] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold60 (.A(\RAM[9][1] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold61 (.A(\RAM[15][4] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold62 (.A(\RAM[14][4] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold63 (.A(\RAM[7][0] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold64 (.A(\RAM[10][4] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold65 (.A(\RAM[9][5] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold66 (.A(\RAM[5][4] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold67 (.A(\RAM[13][5] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold68 (.A(\RAM[11][6] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold69 (.A(\RAM[0][4] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold70 (.A(\RAM[5][1] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold71 (.A(\RAM[7][5] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold72 (.A(\RAM[2][1] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold73 (.A(\RAM[3][4] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold74 (.A(\RAM[15][5] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold75 (.A(\RAM[8][4] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold76 (.A(\RAM[4][6] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold77 (.A(\RAM[3][5] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold78 (.A(\RAM[5][0] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold79 (.A(\RAM[0][3] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold80 (.A(\RAM[4][4] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold81 (.A(\RAM[2][4] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold82 (.A(\RAM[15][6] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold83 (.A(\RAM[8][5] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold84 (.A(\RAM[6][6] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold85 (.A(\RAM[1][1] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold86 (.A(\RAM[1][6] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold87 (.A(\RAM[2][0] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold88 (.A(\RAM[1][0] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold89 (.A(\RAM[12][3] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold90 (.A(\RAM[6][3] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold91 (.A(\RAM[6][7] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold92 (.A(\RAM[2][2] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold93 (.A(\RAM[14][5] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold94 (.A(\RAM[4][1] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold95 (.A(\RAM[11][4] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold96 (.A(\RAM[8][0] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold97 (.A(\RAM[6][4] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold98 (.A(\RAM[2][5] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold99 (.A(\RAM[13][2] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold100 (.A(\RAM[8][6] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold101 (.A(\RAM[12][5] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold102 (.A(\RAM[10][0] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold103 (.A(\RAM[14][1] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold104 (.A(\RAM[12][7] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold105 (.A(\RAM[2][3] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold106 (.A(\RAM[0][2] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold107 (.A(\RAM[6][1] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold108 (.A(\RAM[2][6] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold109 (.A(\RAM[8][1] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold110 (.A(\RAM[6][2] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold111 (.A(\RAM[1][3] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold112 (.A(\RAM[12][6] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold113 (.A(\RAM[12][0] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold114 (.A(\RAM[8][7] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold115 (.A(\RAM[10][6] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold116 (.A(\RAM[4][5] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold117 (.A(\RAM[8][3] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold118 (.A(\RAM[15][0] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold119 (.A(\RAM[1][4] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold120 (.A(\RAM[0][6] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold121 (.A(\RAM[4][0] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold122 (.A(\RAM[11][0] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold123 (.A(\RAM[10][2] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold124 (.A(\RAM[12][4] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold125 (.A(\RAM[10][1] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold126 (.A(\RAM[10][7] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold127 (.A(\RAM[14][0] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold128 (.A(\RAM[11][7] ),
    .X(net285));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_4 FILLER_14_175 ();
 sg13g2_fill_1 FILLER_14_179 ();
 sg13g2_fill_2 FILLER_14_185 ();
 sg13g2_fill_1 FILLER_14_187 ();
 sg13g2_decap_8 FILLER_14_192 ();
 sg13g2_decap_8 FILLER_14_199 ();
 sg13g2_decap_8 FILLER_14_206 ();
 sg13g2_decap_8 FILLER_14_213 ();
 sg13g2_decap_8 FILLER_14_220 ();
 sg13g2_decap_8 FILLER_14_227 ();
 sg13g2_decap_8 FILLER_14_234 ();
 sg13g2_decap_8 FILLER_14_241 ();
 sg13g2_decap_8 FILLER_14_248 ();
 sg13g2_decap_8 FILLER_14_255 ();
 sg13g2_decap_8 FILLER_14_262 ();
 sg13g2_decap_8 FILLER_14_269 ();
 sg13g2_decap_8 FILLER_14_276 ();
 sg13g2_decap_8 FILLER_14_283 ();
 sg13g2_decap_8 FILLER_14_290 ();
 sg13g2_decap_8 FILLER_14_297 ();
 sg13g2_decap_8 FILLER_14_304 ();
 sg13g2_decap_8 FILLER_14_311 ();
 sg13g2_decap_8 FILLER_14_318 ();
 sg13g2_decap_8 FILLER_14_325 ();
 sg13g2_decap_8 FILLER_14_332 ();
 sg13g2_decap_8 FILLER_14_339 ();
 sg13g2_decap_8 FILLER_14_346 ();
 sg13g2_decap_8 FILLER_14_353 ();
 sg13g2_decap_8 FILLER_14_360 ();
 sg13g2_decap_8 FILLER_14_367 ();
 sg13g2_decap_8 FILLER_14_374 ();
 sg13g2_decap_8 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_14_388 ();
 sg13g2_decap_8 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_fill_2 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_fill_2 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_fill_2 FILLER_15_84 ();
 sg13g2_decap_4 FILLER_15_100 ();
 sg13g2_fill_2 FILLER_15_104 ();
 sg13g2_decap_8 FILLER_15_111 ();
 sg13g2_decap_4 FILLER_15_118 ();
 sg13g2_decap_8 FILLER_15_130 ();
 sg13g2_fill_1 FILLER_15_137 ();
 sg13g2_decap_4 FILLER_15_148 ();
 sg13g2_decap_4 FILLER_15_157 ();
 sg13g2_fill_2 FILLER_15_161 ();
 sg13g2_decap_4 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_213 ();
 sg13g2_decap_8 FILLER_15_220 ();
 sg13g2_decap_8 FILLER_15_227 ();
 sg13g2_fill_2 FILLER_15_234 ();
 sg13g2_decap_8 FILLER_15_244 ();
 sg13g2_decap_8 FILLER_15_251 ();
 sg13g2_decap_4 FILLER_15_258 ();
 sg13g2_fill_1 FILLER_15_262 ();
 sg13g2_fill_2 FILLER_15_268 ();
 sg13g2_fill_1 FILLER_15_270 ();
 sg13g2_decap_8 FILLER_15_297 ();
 sg13g2_decap_4 FILLER_15_304 ();
 sg13g2_fill_2 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_314 ();
 sg13g2_decap_8 FILLER_15_321 ();
 sg13g2_decap_8 FILLER_15_328 ();
 sg13g2_decap_8 FILLER_15_335 ();
 sg13g2_decap_8 FILLER_15_342 ();
 sg13g2_decap_8 FILLER_15_349 ();
 sg13g2_decap_8 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_4 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_46 ();
 sg13g2_fill_2 FILLER_16_51 ();
 sg13g2_fill_2 FILLER_16_131 ();
 sg13g2_fill_1 FILLER_16_159 ();
 sg13g2_fill_2 FILLER_16_186 ();
 sg13g2_fill_1 FILLER_16_188 ();
 sg13g2_decap_8 FILLER_16_220 ();
 sg13g2_fill_2 FILLER_16_297 ();
 sg13g2_fill_1 FILLER_16_299 ();
 sg13g2_fill_2 FILLER_16_326 ();
 sg13g2_fill_1 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_338 ();
 sg13g2_decap_4 FILLER_16_345 ();
 sg13g2_fill_1 FILLER_16_349 ();
 sg13g2_decap_4 FILLER_16_355 ();
 sg13g2_decap_8 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_388 ();
 sg13g2_decap_8 FILLER_16_395 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_28 ();
 sg13g2_fill_2 FILLER_17_33 ();
 sg13g2_fill_1 FILLER_17_35 ();
 sg13g2_fill_2 FILLER_17_65 ();
 sg13g2_fill_1 FILLER_17_67 ();
 sg13g2_fill_1 FILLER_17_82 ();
 sg13g2_fill_2 FILLER_17_111 ();
 sg13g2_fill_1 FILLER_17_113 ();
 sg13g2_fill_2 FILLER_17_119 ();
 sg13g2_fill_1 FILLER_17_121 ();
 sg13g2_decap_4 FILLER_17_213 ();
 sg13g2_fill_1 FILLER_17_243 ();
 sg13g2_fill_2 FILLER_17_263 ();
 sg13g2_fill_2 FILLER_17_274 ();
 sg13g2_fill_2 FILLER_17_300 ();
 sg13g2_fill_2 FILLER_17_307 ();
 sg13g2_fill_2 FILLER_17_319 ();
 sg13g2_fill_1 FILLER_17_321 ();
 sg13g2_fill_1 FILLER_17_348 ();
 sg13g2_decap_8 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_11 ();
 sg13g2_fill_2 FILLER_18_17 ();
 sg13g2_fill_1 FILLER_18_45 ();
 sg13g2_fill_2 FILLER_18_55 ();
 sg13g2_fill_1 FILLER_18_57 ();
 sg13g2_fill_2 FILLER_18_104 ();
 sg13g2_fill_1 FILLER_18_137 ();
 sg13g2_fill_2 FILLER_18_219 ();
 sg13g2_fill_2 FILLER_18_231 ();
 sg13g2_fill_1 FILLER_18_233 ();
 sg13g2_fill_1 FILLER_18_264 ();
 sg13g2_fill_2 FILLER_18_280 ();
 sg13g2_fill_2 FILLER_18_313 ();
 sg13g2_fill_1 FILLER_18_315 ();
 sg13g2_fill_2 FILLER_18_336 ();
 sg13g2_fill_1 FILLER_18_338 ();
 sg13g2_fill_2 FILLER_18_363 ();
 sg13g2_fill_1 FILLER_18_365 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_fill_1 FILLER_19_44 ();
 sg13g2_fill_2 FILLER_19_56 ();
 sg13g2_decap_4 FILLER_19_85 ();
 sg13g2_decap_4 FILLER_19_98 ();
 sg13g2_decap_4 FILLER_19_122 ();
 sg13g2_fill_1 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_141 ();
 sg13g2_fill_1 FILLER_19_148 ();
 sg13g2_decap_4 FILLER_19_153 ();
 sg13g2_fill_1 FILLER_19_157 ();
 sg13g2_fill_2 FILLER_19_164 ();
 sg13g2_fill_1 FILLER_19_166 ();
 sg13g2_fill_2 FILLER_19_175 ();
 sg13g2_decap_4 FILLER_19_195 ();
 sg13g2_fill_1 FILLER_19_199 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_4 FILLER_19_217 ();
 sg13g2_fill_2 FILLER_19_242 ();
 sg13g2_fill_1 FILLER_19_244 ();
 sg13g2_fill_2 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_282 ();
 sg13g2_fill_1 FILLER_19_288 ();
 sg13g2_fill_1 FILLER_19_297 ();
 sg13g2_fill_1 FILLER_19_326 ();
 sg13g2_fill_2 FILLER_19_353 ();
 sg13g2_fill_1 FILLER_19_361 ();
 sg13g2_fill_2 FILLER_19_380 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_30 ();
 sg13g2_fill_1 FILLER_20_32 ();
 sg13g2_fill_2 FILLER_20_65 ();
 sg13g2_fill_2 FILLER_20_107 ();
 sg13g2_fill_1 FILLER_20_109 ();
 sg13g2_fill_1 FILLER_20_149 ();
 sg13g2_decap_4 FILLER_20_155 ();
 sg13g2_fill_1 FILLER_20_164 ();
 sg13g2_decap_4 FILLER_20_183 ();
 sg13g2_fill_1 FILLER_20_187 ();
 sg13g2_decap_4 FILLER_20_193 ();
 sg13g2_fill_2 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_223 ();
 sg13g2_fill_1 FILLER_20_229 ();
 sg13g2_fill_2 FILLER_20_240 ();
 sg13g2_fill_1 FILLER_20_242 ();
 sg13g2_fill_2 FILLER_20_304 ();
 sg13g2_fill_1 FILLER_20_306 ();
 sg13g2_fill_2 FILLER_20_350 ();
 sg13g2_fill_1 FILLER_20_361 ();
 sg13g2_fill_1 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_45 ();
 sg13g2_fill_1 FILLER_21_47 ();
 sg13g2_fill_1 FILLER_21_53 ();
 sg13g2_decap_4 FILLER_21_81 ();
 sg13g2_decap_4 FILLER_21_94 ();
 sg13g2_fill_1 FILLER_21_98 ();
 sg13g2_fill_1 FILLER_21_104 ();
 sg13g2_fill_2 FILLER_21_118 ();
 sg13g2_fill_1 FILLER_21_120 ();
 sg13g2_fill_2 FILLER_21_134 ();
 sg13g2_fill_2 FILLER_21_230 ();
 sg13g2_fill_1 FILLER_21_257 ();
 sg13g2_fill_2 FILLER_21_277 ();
 sg13g2_fill_1 FILLER_21_279 ();
 sg13g2_decap_8 FILLER_21_293 ();
 sg13g2_fill_2 FILLER_21_300 ();
 sg13g2_decap_4 FILLER_21_307 ();
 sg13g2_fill_2 FILLER_21_316 ();
 sg13g2_fill_1 FILLER_21_318 ();
 sg13g2_fill_1 FILLER_21_388 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_36 ();
 sg13g2_fill_1 FILLER_22_38 ();
 sg13g2_decap_8 FILLER_22_96 ();
 sg13g2_fill_2 FILLER_22_103 ();
 sg13g2_fill_1 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_132 ();
 sg13g2_fill_2 FILLER_22_167 ();
 sg13g2_decap_8 FILLER_22_198 ();
 sg13g2_fill_1 FILLER_22_251 ();
 sg13g2_fill_1 FILLER_22_329 ();
 sg13g2_fill_2 FILLER_22_334 ();
 sg13g2_fill_1 FILLER_22_336 ();
 sg13g2_fill_1 FILLER_22_368 ();
 sg13g2_fill_1 FILLER_22_374 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_4 ();
 sg13g2_fill_1 FILLER_23_44 ();
 sg13g2_fill_2 FILLER_23_133 ();
 sg13g2_fill_1 FILLER_23_135 ();
 sg13g2_fill_1 FILLER_23_149 ();
 sg13g2_fill_2 FILLER_23_217 ();
 sg13g2_fill_1 FILLER_23_219 ();
 sg13g2_decap_4 FILLER_23_225 ();
 sg13g2_fill_2 FILLER_23_229 ();
 sg13g2_fill_1 FILLER_23_235 ();
 sg13g2_fill_1 FILLER_23_241 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_fill_2 FILLER_23_280 ();
 sg13g2_fill_1 FILLER_23_310 ();
 sg13g2_fill_2 FILLER_23_337 ();
 sg13g2_fill_2 FILLER_23_367 ();
 sg13g2_fill_1 FILLER_23_369 ();
 sg13g2_fill_2 FILLER_23_380 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_18 ();
 sg13g2_decap_8 FILLER_24_24 ();
 sg13g2_fill_2 FILLER_24_55 ();
 sg13g2_fill_2 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_93 ();
 sg13g2_fill_1 FILLER_24_99 ();
 sg13g2_decap_4 FILLER_24_124 ();
 sg13g2_fill_1 FILLER_24_154 ();
 sg13g2_fill_1 FILLER_24_169 ();
 sg13g2_fill_1 FILLER_24_175 ();
 sg13g2_fill_1 FILLER_24_181 ();
 sg13g2_fill_2 FILLER_24_197 ();
 sg13g2_fill_1 FILLER_24_199 ();
 sg13g2_fill_1 FILLER_24_260 ();
 sg13g2_fill_2 FILLER_24_270 ();
 sg13g2_fill_1 FILLER_24_272 ();
 sg13g2_fill_1 FILLER_24_278 ();
 sg13g2_fill_1 FILLER_24_284 ();
 sg13g2_decap_8 FILLER_24_299 ();
 sg13g2_fill_2 FILLER_24_316 ();
 sg13g2_fill_2 FILLER_24_327 ();
 sg13g2_fill_2 FILLER_24_335 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_fill_1 FILLER_25_30 ();
 sg13g2_fill_2 FILLER_25_70 ();
 sg13g2_fill_2 FILLER_25_98 ();
 sg13g2_fill_1 FILLER_25_100 ();
 sg13g2_fill_2 FILLER_25_133 ();
 sg13g2_fill_1 FILLER_25_135 ();
 sg13g2_decap_8 FILLER_25_174 ();
 sg13g2_decap_4 FILLER_25_181 ();
 sg13g2_fill_2 FILLER_25_185 ();
 sg13g2_decap_4 FILLER_25_193 ();
 sg13g2_fill_1 FILLER_25_197 ();
 sg13g2_decap_4 FILLER_25_220 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_229 ();
 sg13g2_fill_1 FILLER_25_236 ();
 sg13g2_fill_2 FILLER_25_262 ();
 sg13g2_fill_1 FILLER_25_275 ();
 sg13g2_decap_4 FILLER_25_308 ();
 sg13g2_fill_2 FILLER_25_356 ();
 sg13g2_fill_2 FILLER_25_379 ();
 sg13g2_fill_1 FILLER_25_381 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_14 ();
 sg13g2_fill_2 FILLER_26_41 ();
 sg13g2_fill_1 FILLER_26_93 ();
 sg13g2_fill_2 FILLER_26_99 ();
 sg13g2_fill_1 FILLER_26_101 ();
 sg13g2_fill_2 FILLER_26_115 ();
 sg13g2_fill_1 FILLER_26_117 ();
 sg13g2_fill_2 FILLER_26_144 ();
 sg13g2_fill_1 FILLER_26_146 ();
 sg13g2_fill_1 FILLER_26_165 ();
 sg13g2_decap_8 FILLER_26_180 ();
 sg13g2_decap_8 FILLER_26_187 ();
 sg13g2_fill_2 FILLER_26_200 ();
 sg13g2_fill_2 FILLER_26_210 ();
 sg13g2_fill_1 FILLER_26_212 ();
 sg13g2_decap_8 FILLER_26_218 ();
 sg13g2_fill_1 FILLER_26_251 ();
 sg13g2_fill_1 FILLER_26_276 ();
 sg13g2_fill_1 FILLER_26_282 ();
 sg13g2_fill_1 FILLER_26_315 ();
 sg13g2_fill_2 FILLER_26_334 ();
 sg13g2_fill_2 FILLER_26_349 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_60 ();
 sg13g2_fill_2 FILLER_27_103 ();
 sg13g2_decap_4 FILLER_27_127 ();
 sg13g2_fill_1 FILLER_27_131 ();
 sg13g2_decap_4 FILLER_27_137 ();
 sg13g2_fill_2 FILLER_27_141 ();
 sg13g2_decap_8 FILLER_27_150 ();
 sg13g2_decap_8 FILLER_27_162 ();
 sg13g2_decap_8 FILLER_27_169 ();
 sg13g2_fill_2 FILLER_27_181 ();
 sg13g2_fill_2 FILLER_27_200 ();
 sg13g2_decap_8 FILLER_27_229 ();
 sg13g2_fill_2 FILLER_27_236 ();
 sg13g2_decap_8 FILLER_27_247 ();
 sg13g2_fill_1 FILLER_27_254 ();
 sg13g2_decap_4 FILLER_27_303 ();
 sg13g2_fill_1 FILLER_27_307 ();
 sg13g2_fill_2 FILLER_27_334 ();
 sg13g2_fill_2 FILLER_27_390 ();
 sg13g2_fill_1 FILLER_28_30 ();
 sg13g2_fill_1 FILLER_28_60 ();
 sg13g2_fill_1 FILLER_28_75 ();
 sg13g2_decap_8 FILLER_28_81 ();
 sg13g2_fill_2 FILLER_28_88 ();
 sg13g2_fill_2 FILLER_28_99 ();
 sg13g2_fill_1 FILLER_28_101 ();
 sg13g2_fill_1 FILLER_28_118 ();
 sg13g2_fill_1 FILLER_28_134 ();
 sg13g2_decap_4 FILLER_28_169 ();
 sg13g2_decap_8 FILLER_28_208 ();
 sg13g2_fill_1 FILLER_28_215 ();
 sg13g2_decap_8 FILLER_28_242 ();
 sg13g2_fill_2 FILLER_28_270 ();
 sg13g2_fill_1 FILLER_28_272 ();
 sg13g2_fill_1 FILLER_28_310 ();
 sg13g2_fill_2 FILLER_28_316 ();
 sg13g2_fill_1 FILLER_28_318 ();
 sg13g2_fill_2 FILLER_28_323 ();
 sg13g2_fill_1 FILLER_28_325 ();
 sg13g2_fill_2 FILLER_28_338 ();
 sg13g2_fill_1 FILLER_28_367 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_34 ();
 sg13g2_fill_2 FILLER_29_51 ();
 sg13g2_fill_2 FILLER_29_59 ();
 sg13g2_decap_4 FILLER_29_87 ();
 sg13g2_fill_1 FILLER_29_143 ();
 sg13g2_decap_8 FILLER_29_206 ();
 sg13g2_fill_2 FILLER_29_213 ();
 sg13g2_decap_4 FILLER_29_219 ();
 sg13g2_fill_1 FILLER_29_223 ();
 sg13g2_fill_1 FILLER_29_252 ();
 sg13g2_fill_2 FILLER_29_258 ();
 sg13g2_fill_1 FILLER_29_270 ();
 sg13g2_fill_1 FILLER_29_275 ();
 sg13g2_fill_2 FILLER_29_281 ();
 sg13g2_decap_4 FILLER_29_287 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_312 ();
 sg13g2_fill_1 FILLER_29_324 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_54 ();
 sg13g2_decap_8 FILLER_30_64 ();
 sg13g2_fill_2 FILLER_30_71 ();
 sg13g2_fill_2 FILLER_30_122 ();
 sg13g2_fill_1 FILLER_30_142 ();
 sg13g2_decap_4 FILLER_30_247 ();
 sg13g2_fill_2 FILLER_30_277 ();
 sg13g2_fill_1 FILLER_30_279 ();
 sg13g2_fill_2 FILLER_30_285 ();
 sg13g2_fill_1 FILLER_30_287 ();
 sg13g2_fill_1 FILLER_30_346 ();
 sg13g2_fill_1 FILLER_30_361 ();
 sg13g2_fill_2 FILLER_30_368 ();
 sg13g2_fill_1 FILLER_30_370 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_14 ();
 sg13g2_decap_4 FILLER_31_20 ();
 sg13g2_fill_1 FILLER_31_24 ();
 sg13g2_fill_2 FILLER_31_59 ();
 sg13g2_fill_2 FILLER_31_115 ();
 sg13g2_fill_2 FILLER_31_183 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_fill_2 FILLER_31_217 ();
 sg13g2_fill_2 FILLER_31_263 ();
 sg13g2_fill_1 FILLER_31_313 ();
 sg13g2_fill_2 FILLER_31_326 ();
 sg13g2_fill_2 FILLER_31_365 ();
 sg13g2_fill_1 FILLER_31_367 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_4 ();
 sg13g2_fill_2 FILLER_32_40 ();
 sg13g2_fill_2 FILLER_32_66 ();
 sg13g2_fill_2 FILLER_32_92 ();
 sg13g2_fill_1 FILLER_32_94 ();
 sg13g2_fill_2 FILLER_32_116 ();
 sg13g2_fill_2 FILLER_32_147 ();
 sg13g2_fill_2 FILLER_32_154 ();
 sg13g2_fill_2 FILLER_32_181 ();
 sg13g2_decap_4 FILLER_32_204 ();
 sg13g2_fill_2 FILLER_32_248 ();
 sg13g2_fill_1 FILLER_32_293 ();
 sg13g2_fill_2 FILLER_32_299 ();
 sg13g2_fill_1 FILLER_32_301 ();
 sg13g2_fill_1 FILLER_32_320 ();
 sg13g2_fill_2 FILLER_32_378 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_fill_2 FILLER_33_28 ();
 sg13g2_fill_2 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_157 ();
 sg13g2_decap_4 FILLER_33_203 ();
 sg13g2_fill_2 FILLER_33_207 ();
 sg13g2_fill_1 FILLER_33_239 ();
 sg13g2_fill_1 FILLER_33_260 ();
 sg13g2_fill_1 FILLER_33_266 ();
 sg13g2_fill_2 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_313 ();
 sg13g2_fill_1 FILLER_33_346 ();
 sg13g2_fill_1 FILLER_33_387 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_fill_2 FILLER_34_44 ();
 sg13g2_fill_1 FILLER_34_61 ();
 sg13g2_fill_1 FILLER_34_84 ();
 sg13g2_fill_2 FILLER_34_89 ();
 sg13g2_fill_2 FILLER_34_99 ();
 sg13g2_fill_2 FILLER_34_106 ();
 sg13g2_fill_1 FILLER_34_134 ();
 sg13g2_fill_2 FILLER_34_144 ();
 sg13g2_fill_1 FILLER_34_146 ();
 sg13g2_decap_4 FILLER_34_183 ();
 sg13g2_fill_1 FILLER_34_187 ();
 sg13g2_decap_4 FILLER_34_192 ();
 sg13g2_fill_2 FILLER_34_204 ();
 sg13g2_fill_2 FILLER_34_218 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_fill_2 FILLER_34_231 ();
 sg13g2_fill_1 FILLER_34_233 ();
 sg13g2_fill_2 FILLER_34_335 ();
 sg13g2_fill_2 FILLER_34_342 ();
 sg13g2_fill_2 FILLER_34_349 ();
 sg13g2_fill_1 FILLER_34_351 ();
 sg13g2_fill_2 FILLER_34_363 ();
 sg13g2_fill_1 FILLER_34_365 ();
 sg13g2_fill_1 FILLER_34_381 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_fill_2 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_51 ();
 sg13g2_decap_4 FILLER_35_78 ();
 sg13g2_fill_2 FILLER_35_123 ();
 sg13g2_fill_2 FILLER_35_154 ();
 sg13g2_fill_1 FILLER_35_156 ();
 sg13g2_fill_1 FILLER_35_255 ();
 sg13g2_fill_2 FILLER_35_290 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_fill_2 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_65 ();
 sg13g2_decap_4 FILLER_36_71 ();
 sg13g2_fill_1 FILLER_36_125 ();
 sg13g2_fill_2 FILLER_36_152 ();
 sg13g2_fill_1 FILLER_36_154 ();
 sg13g2_fill_2 FILLER_36_167 ();
 sg13g2_fill_2 FILLER_36_179 ();
 sg13g2_fill_1 FILLER_36_200 ();
 sg13g2_fill_2 FILLER_36_244 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_fill_2 FILLER_36_280 ();
 sg13g2_fill_2 FILLER_36_389 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_4 FILLER_37_63 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_fill_1 FILLER_37_95 ();
 sg13g2_fill_1 FILLER_37_124 ();
 sg13g2_fill_2 FILLER_37_148 ();
 sg13g2_fill_1 FILLER_37_202 ();
 sg13g2_decap_4 FILLER_37_214 ();
 sg13g2_fill_2 FILLER_37_218 ();
 sg13g2_fill_2 FILLER_37_349 ();
 sg13g2_fill_1 FILLER_37_351 ();
 sg13g2_fill_1 FILLER_37_371 ();
 sg13g2_fill_1 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_4 FILLER_38_49 ();
 sg13g2_fill_1 FILLER_38_120 ();
 sg13g2_fill_1 FILLER_38_172 ();
 sg13g2_fill_2 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_197 ();
 sg13g2_decap_8 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_211 ();
 sg13g2_fill_2 FILLER_38_245 ();
 sg13g2_fill_1 FILLER_38_247 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_fill_1 FILLER_38_285 ();
 sg13g2_fill_2 FILLER_38_336 ();
 sg13g2_fill_1 FILLER_38_338 ();
 sg13g2_fill_2 FILLER_38_360 ();
 sg13g2_fill_1 FILLER_38_362 ();
 sg13g2_fill_2 FILLER_38_389 ();
 sg13g2_fill_1 FILLER_38_391 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net14;
 assign uio_oe[1] = net15;
 assign uio_oe[2] = net16;
 assign uio_oe[3] = net17;
 assign uio_oe[4] = net18;
 assign uio_oe[5] = net19;
 assign uio_oe[6] = net20;
 assign uio_oe[7] = net21;
 assign uio_out[0] = net22;
 assign uio_out[1] = net23;
 assign uio_out[2] = net24;
 assign uio_out[3] = net25;
 assign uio_out[4] = net26;
 assign uio_out[5] = net27;
 assign uio_out[6] = net28;
 assign uio_out[7] = net29;
endmodule

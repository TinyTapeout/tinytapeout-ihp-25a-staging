module tt_um_bitty (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire clknet_leaf_0_clk;
 wire \addr[0] ;
 wire \addr[1] ;
 wire \addr[2] ;
 wire \addr[3] ;
 wire \addr[4] ;
 wire \addr[5] ;
 wire \addr[6] ;
 wire \addr[7] ;
 wire \bitty_inst.alu_inst.in_a[0] ;
 wire \bitty_inst.alu_inst.in_a[10] ;
 wire \bitty_inst.alu_inst.in_a[11] ;
 wire \bitty_inst.alu_inst.in_a[12] ;
 wire \bitty_inst.alu_inst.in_a[13] ;
 wire \bitty_inst.alu_inst.in_a[14] ;
 wire \bitty_inst.alu_inst.in_a[15] ;
 wire \bitty_inst.alu_inst.in_a[1] ;
 wire \bitty_inst.alu_inst.in_a[2] ;
 wire \bitty_inst.alu_inst.in_a[3] ;
 wire \bitty_inst.alu_inst.in_a[4] ;
 wire \bitty_inst.alu_inst.in_a[5] ;
 wire \bitty_inst.alu_inst.in_a[6] ;
 wire \bitty_inst.alu_inst.in_a[7] ;
 wire \bitty_inst.alu_inst.in_a[8] ;
 wire \bitty_inst.alu_inst.in_a[9] ;
 wire \bitty_inst.cpu_inst.cur_state[0] ;
 wire \bitty_inst.cpu_inst.cur_state[1] ;
 wire \bitty_inst.cpu_inst.cur_state[2] ;
 wire \bitty_inst.cpu_inst.d_inst[0] ;
 wire \bitty_inst.cpu_inst.d_inst[10] ;
 wire \bitty_inst.cpu_inst.d_inst[11] ;
 wire \bitty_inst.cpu_inst.d_inst[12] ;
 wire \bitty_inst.cpu_inst.d_inst[13] ;
 wire \bitty_inst.cpu_inst.d_inst[14] ;
 wire \bitty_inst.cpu_inst.d_inst[15] ;
 wire \bitty_inst.cpu_inst.d_inst[1] ;
 wire \bitty_inst.cpu_inst.d_inst[2] ;
 wire \bitty_inst.cpu_inst.d_inst[3] ;
 wire \bitty_inst.cpu_inst.d_inst[4] ;
 wire \bitty_inst.cpu_inst.d_inst[5] ;
 wire \bitty_inst.cpu_inst.d_inst[6] ;
 wire \bitty_inst.cpu_inst.d_inst[7] ;
 wire \bitty_inst.cpu_inst.d_inst[8] ;
 wire \bitty_inst.cpu_inst.d_inst[9] ;
 wire \bitty_inst.cpu_inst.run ;
 wire \bitty_inst.d_instr[0] ;
 wire \bitty_inst.d_instr[10] ;
 wire \bitty_inst.d_instr[11] ;
 wire \bitty_inst.d_instr[12] ;
 wire \bitty_inst.d_instr[13] ;
 wire \bitty_inst.d_instr[14] ;
 wire \bitty_inst.d_instr[15] ;
 wire \bitty_inst.d_instr[1] ;
 wire \bitty_inst.d_instr[2] ;
 wire \bitty_inst.d_instr[3] ;
 wire \bitty_inst.d_instr[4] ;
 wire \bitty_inst.d_instr[5] ;
 wire \bitty_inst.d_instr[6] ;
 wire \bitty_inst.d_instr[7] ;
 wire \bitty_inst.d_instr[8] ;
 wire \bitty_inst.d_instr[9] ;
 wire \bitty_inst.d_out[0] ;
 wire \bitty_inst.d_out[10] ;
 wire \bitty_inst.d_out[11] ;
 wire \bitty_inst.d_out[12] ;
 wire \bitty_inst.d_out[13] ;
 wire \bitty_inst.d_out[14] ;
 wire \bitty_inst.d_out[15] ;
 wire \bitty_inst.d_out[1] ;
 wire \bitty_inst.d_out[2] ;
 wire \bitty_inst.d_out[3] ;
 wire \bitty_inst.d_out[4] ;
 wire \bitty_inst.d_out[5] ;
 wire \bitty_inst.d_out[6] ;
 wire \bitty_inst.d_out[7] ;
 wire \bitty_inst.d_out[8] ;
 wire \bitty_inst.d_out[9] ;
 wire \bitty_inst.data_to_ld[0] ;
 wire \bitty_inst.data_to_ld[10] ;
 wire \bitty_inst.data_to_ld[11] ;
 wire \bitty_inst.data_to_ld[12] ;
 wire \bitty_inst.data_to_ld[13] ;
 wire \bitty_inst.data_to_ld[14] ;
 wire \bitty_inst.data_to_ld[15] ;
 wire \bitty_inst.data_to_ld[1] ;
 wire \bitty_inst.data_to_ld[2] ;
 wire \bitty_inst.data_to_ld[3] ;
 wire \bitty_inst.data_to_ld[4] ;
 wire \bitty_inst.data_to_ld[5] ;
 wire \bitty_inst.data_to_ld[6] ;
 wire \bitty_inst.data_to_ld[7] ;
 wire \bitty_inst.data_to_ld[8] ;
 wire \bitty_inst.data_to_ld[9] ;
 wire \bitty_inst.gen_dff[0].reg_out.mux_out[0] ;
 wire \bitty_inst.gen_dff[0].reg_out.mux_out[10] ;
 wire \bitty_inst.gen_dff[0].reg_out.mux_out[11] ;
 wire \bitty_inst.gen_dff[0].reg_out.mux_out[12] ;
 wire \bitty_inst.gen_dff[0].reg_out.mux_out[13] ;
 wire \bitty_inst.gen_dff[0].reg_out.mux_out[14] ;
 wire \bitty_inst.gen_dff[0].reg_out.mux_out[15] ;
 wire \bitty_inst.gen_dff[0].reg_out.mux_out[1] ;
 wire \bitty_inst.gen_dff[0].reg_out.mux_out[2] ;
 wire \bitty_inst.gen_dff[0].reg_out.mux_out[3] ;
 wire \bitty_inst.gen_dff[0].reg_out.mux_out[4] ;
 wire \bitty_inst.gen_dff[0].reg_out.mux_out[5] ;
 wire \bitty_inst.gen_dff[0].reg_out.mux_out[6] ;
 wire \bitty_inst.gen_dff[0].reg_out.mux_out[7] ;
 wire \bitty_inst.gen_dff[0].reg_out.mux_out[8] ;
 wire \bitty_inst.gen_dff[0].reg_out.mux_out[9] ;
 wire \bitty_inst.gen_dff[1].reg_out.mux_out[0] ;
 wire \bitty_inst.gen_dff[1].reg_out.mux_out[10] ;
 wire \bitty_inst.gen_dff[1].reg_out.mux_out[11] ;
 wire \bitty_inst.gen_dff[1].reg_out.mux_out[12] ;
 wire \bitty_inst.gen_dff[1].reg_out.mux_out[13] ;
 wire \bitty_inst.gen_dff[1].reg_out.mux_out[14] ;
 wire \bitty_inst.gen_dff[1].reg_out.mux_out[15] ;
 wire \bitty_inst.gen_dff[1].reg_out.mux_out[1] ;
 wire \bitty_inst.gen_dff[1].reg_out.mux_out[2] ;
 wire \bitty_inst.gen_dff[1].reg_out.mux_out[3] ;
 wire \bitty_inst.gen_dff[1].reg_out.mux_out[4] ;
 wire \bitty_inst.gen_dff[1].reg_out.mux_out[5] ;
 wire \bitty_inst.gen_dff[1].reg_out.mux_out[6] ;
 wire \bitty_inst.gen_dff[1].reg_out.mux_out[7] ;
 wire \bitty_inst.gen_dff[1].reg_out.mux_out[8] ;
 wire \bitty_inst.gen_dff[1].reg_out.mux_out[9] ;
 wire \bitty_inst.gen_dff[2].reg_out.mux_out[0] ;
 wire \bitty_inst.gen_dff[2].reg_out.mux_out[10] ;
 wire \bitty_inst.gen_dff[2].reg_out.mux_out[11] ;
 wire \bitty_inst.gen_dff[2].reg_out.mux_out[12] ;
 wire \bitty_inst.gen_dff[2].reg_out.mux_out[13] ;
 wire \bitty_inst.gen_dff[2].reg_out.mux_out[14] ;
 wire \bitty_inst.gen_dff[2].reg_out.mux_out[15] ;
 wire \bitty_inst.gen_dff[2].reg_out.mux_out[1] ;
 wire \bitty_inst.gen_dff[2].reg_out.mux_out[2] ;
 wire \bitty_inst.gen_dff[2].reg_out.mux_out[3] ;
 wire \bitty_inst.gen_dff[2].reg_out.mux_out[4] ;
 wire \bitty_inst.gen_dff[2].reg_out.mux_out[5] ;
 wire \bitty_inst.gen_dff[2].reg_out.mux_out[6] ;
 wire \bitty_inst.gen_dff[2].reg_out.mux_out[7] ;
 wire \bitty_inst.gen_dff[2].reg_out.mux_out[8] ;
 wire \bitty_inst.gen_dff[2].reg_out.mux_out[9] ;
 wire \bitty_inst.gen_dff[3].reg_out.mux_out[0] ;
 wire \bitty_inst.gen_dff[3].reg_out.mux_out[10] ;
 wire \bitty_inst.gen_dff[3].reg_out.mux_out[11] ;
 wire \bitty_inst.gen_dff[3].reg_out.mux_out[12] ;
 wire \bitty_inst.gen_dff[3].reg_out.mux_out[13] ;
 wire \bitty_inst.gen_dff[3].reg_out.mux_out[14] ;
 wire \bitty_inst.gen_dff[3].reg_out.mux_out[15] ;
 wire \bitty_inst.gen_dff[3].reg_out.mux_out[1] ;
 wire \bitty_inst.gen_dff[3].reg_out.mux_out[2] ;
 wire \bitty_inst.gen_dff[3].reg_out.mux_out[3] ;
 wire \bitty_inst.gen_dff[3].reg_out.mux_out[4] ;
 wire \bitty_inst.gen_dff[3].reg_out.mux_out[5] ;
 wire \bitty_inst.gen_dff[3].reg_out.mux_out[6] ;
 wire \bitty_inst.gen_dff[3].reg_out.mux_out[7] ;
 wire \bitty_inst.gen_dff[3].reg_out.mux_out[8] ;
 wire \bitty_inst.gen_dff[3].reg_out.mux_out[9] ;
 wire \bitty_inst.gen_dff[4].reg_out.mux_out[0] ;
 wire \bitty_inst.gen_dff[4].reg_out.mux_out[10] ;
 wire \bitty_inst.gen_dff[4].reg_out.mux_out[11] ;
 wire \bitty_inst.gen_dff[4].reg_out.mux_out[12] ;
 wire \bitty_inst.gen_dff[4].reg_out.mux_out[13] ;
 wire \bitty_inst.gen_dff[4].reg_out.mux_out[14] ;
 wire \bitty_inst.gen_dff[4].reg_out.mux_out[15] ;
 wire \bitty_inst.gen_dff[4].reg_out.mux_out[1] ;
 wire \bitty_inst.gen_dff[4].reg_out.mux_out[2] ;
 wire \bitty_inst.gen_dff[4].reg_out.mux_out[3] ;
 wire \bitty_inst.gen_dff[4].reg_out.mux_out[4] ;
 wire \bitty_inst.gen_dff[4].reg_out.mux_out[5] ;
 wire \bitty_inst.gen_dff[4].reg_out.mux_out[6] ;
 wire \bitty_inst.gen_dff[4].reg_out.mux_out[7] ;
 wire \bitty_inst.gen_dff[4].reg_out.mux_out[8] ;
 wire \bitty_inst.gen_dff[4].reg_out.mux_out[9] ;
 wire \bitty_inst.gen_dff[5].reg_out.mux_out[0] ;
 wire \bitty_inst.gen_dff[5].reg_out.mux_out[10] ;
 wire \bitty_inst.gen_dff[5].reg_out.mux_out[11] ;
 wire \bitty_inst.gen_dff[5].reg_out.mux_out[12] ;
 wire \bitty_inst.gen_dff[5].reg_out.mux_out[13] ;
 wire \bitty_inst.gen_dff[5].reg_out.mux_out[14] ;
 wire \bitty_inst.gen_dff[5].reg_out.mux_out[15] ;
 wire \bitty_inst.gen_dff[5].reg_out.mux_out[1] ;
 wire \bitty_inst.gen_dff[5].reg_out.mux_out[2] ;
 wire \bitty_inst.gen_dff[5].reg_out.mux_out[3] ;
 wire \bitty_inst.gen_dff[5].reg_out.mux_out[4] ;
 wire \bitty_inst.gen_dff[5].reg_out.mux_out[5] ;
 wire \bitty_inst.gen_dff[5].reg_out.mux_out[6] ;
 wire \bitty_inst.gen_dff[5].reg_out.mux_out[7] ;
 wire \bitty_inst.gen_dff[5].reg_out.mux_out[8] ;
 wire \bitty_inst.gen_dff[5].reg_out.mux_out[9] ;
 wire \bitty_inst.gen_dff[6].reg_out.mux_out[0] ;
 wire \bitty_inst.gen_dff[6].reg_out.mux_out[10] ;
 wire \bitty_inst.gen_dff[6].reg_out.mux_out[11] ;
 wire \bitty_inst.gen_dff[6].reg_out.mux_out[12] ;
 wire \bitty_inst.gen_dff[6].reg_out.mux_out[13] ;
 wire \bitty_inst.gen_dff[6].reg_out.mux_out[14] ;
 wire \bitty_inst.gen_dff[6].reg_out.mux_out[15] ;
 wire \bitty_inst.gen_dff[6].reg_out.mux_out[1] ;
 wire \bitty_inst.gen_dff[6].reg_out.mux_out[2] ;
 wire \bitty_inst.gen_dff[6].reg_out.mux_out[3] ;
 wire \bitty_inst.gen_dff[6].reg_out.mux_out[4] ;
 wire \bitty_inst.gen_dff[6].reg_out.mux_out[5] ;
 wire \bitty_inst.gen_dff[6].reg_out.mux_out[6] ;
 wire \bitty_inst.gen_dff[6].reg_out.mux_out[7] ;
 wire \bitty_inst.gen_dff[6].reg_out.mux_out[8] ;
 wire \bitty_inst.gen_dff[6].reg_out.mux_out[9] ;
 wire \bitty_inst.gen_dff[7].reg_out.mux_out[0] ;
 wire \bitty_inst.gen_dff[7].reg_out.mux_out[10] ;
 wire \bitty_inst.gen_dff[7].reg_out.mux_out[11] ;
 wire \bitty_inst.gen_dff[7].reg_out.mux_out[12] ;
 wire \bitty_inst.gen_dff[7].reg_out.mux_out[13] ;
 wire \bitty_inst.gen_dff[7].reg_out.mux_out[14] ;
 wire \bitty_inst.gen_dff[7].reg_out.mux_out[15] ;
 wire \bitty_inst.gen_dff[7].reg_out.mux_out[1] ;
 wire \bitty_inst.gen_dff[7].reg_out.mux_out[2] ;
 wire \bitty_inst.gen_dff[7].reg_out.mux_out[3] ;
 wire \bitty_inst.gen_dff[7].reg_out.mux_out[4] ;
 wire \bitty_inst.gen_dff[7].reg_out.mux_out[5] ;
 wire \bitty_inst.gen_dff[7].reg_out.mux_out[6] ;
 wire \bitty_inst.gen_dff[7].reg_out.mux_out[7] ;
 wire \bitty_inst.gen_dff[7].reg_out.mux_out[8] ;
 wire \bitty_inst.gen_dff[7].reg_out.mux_out[9] ;
 wire \bitty_inst.lsu_inst.next_state[0] ;
 wire \bitty_inst.lsu_inst.next_state[1] ;
 wire \bitty_inst.lsu_inst.next_state[2] ;
 wire \bitty_inst.lsu_inst.rx_data[0] ;
 wire \bitty_inst.lsu_inst.rx_data[1] ;
 wire \bitty_inst.lsu_inst.rx_data[2] ;
 wire \bitty_inst.lsu_inst.rx_data[3] ;
 wire \bitty_inst.lsu_inst.rx_data[4] ;
 wire \bitty_inst.lsu_inst.rx_data[5] ;
 wire \bitty_inst.lsu_inst.rx_data[6] ;
 wire \bitty_inst.lsu_inst.rx_data[7] ;
 wire \bitty_inst.lsu_inst.rx_do ;
 wire \bitty_inst.lsu_inst.state[0] ;
 wire \bitty_inst.lsu_inst.state[1] ;
 wire \bitty_inst.lsu_inst.state[2] ;
 wire \bitty_inst.lsu_inst.tx_done ;
 wire \cur_state[0] ;
 wire \cur_state[1] ;
 wire \cur_state[2] ;
 wire \cur_state[3] ;
 wire \cur_state[4] ;
 wire \cur_state[6] ;
 wire \cur_state[7] ;
 wire fetch_done;
 wire \fi_inst.state[0] ;
 wire \fi_inst.state[1] ;
 wire \fi_inst.state[2] ;
 wire \fi_inst.state[4] ;
 wire \fi_inst.state[5] ;
 wire tx_data_bit;
 wire \uart_inst.R0.PS[0] ;
 wire \uart_inst.R0.PS[1] ;
 wire \uart_inst.R0.PS[2] ;
 wire \uart_inst.R0.PS[3] ;
 wire \uart_inst.R0.PS[5] ;
 wire \uart_inst.R0.bit_counter[0] ;
 wire \uart_inst.R0.bit_counter[1] ;
 wire \uart_inst.R0.bit_counter[2] ;
 wire \uart_inst.R0.clk_counter[0] ;
 wire \uart_inst.R0.clk_counter[10] ;
 wire \uart_inst.R0.clk_counter[11] ;
 wire \uart_inst.R0.clk_counter[12] ;
 wire \uart_inst.R0.clk_counter[1] ;
 wire \uart_inst.R0.clk_counter[2] ;
 wire \uart_inst.R0.clk_counter[3] ;
 wire \uart_inst.R0.clk_counter[4] ;
 wire \uart_inst.R0.clk_counter[5] ;
 wire \uart_inst.R0.clk_counter[6] ;
 wire \uart_inst.R0.clk_counter[7] ;
 wire \uart_inst.R0.clk_counter[8] ;
 wire \uart_inst.R0.clk_counter[9] ;
 wire \uart_inst.T0.PS[0] ;
 wire \uart_inst.T0.PS[1] ;
 wire \uart_inst.T0.PS[2] ;
 wire \uart_inst.T0.PS[4] ;
 wire \uart_inst.T0.bit_counter[0] ;
 wire \uart_inst.T0.bit_counter[1] ;
 wire \uart_inst.T0.bit_counter[2] ;
 wire \uart_inst.T0.clk_counter[0] ;
 wire \uart_inst.T0.clk_counter[10] ;
 wire \uart_inst.T0.clk_counter[11] ;
 wire \uart_inst.T0.clk_counter[12] ;
 wire \uart_inst.T0.clk_counter[1] ;
 wire \uart_inst.T0.clk_counter[2] ;
 wire \uart_inst.T0.clk_counter[3] ;
 wire \uart_inst.T0.clk_counter[4] ;
 wire \uart_inst.T0.clk_counter[5] ;
 wire \uart_inst.T0.clk_counter[6] ;
 wire \uart_inst.T0.clk_counter[7] ;
 wire \uart_inst.T0.clk_counter[8] ;
 wire \uart_inst.T0.clk_counter[9] ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net1;
 wire net2;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;

 sg13g2_inv_1 _2188_ (.Y(_1341_),
    .A(net962));
 sg13g2_inv_1 _2189_ (.Y(_1342_),
    .A(net916));
 sg13g2_inv_2 _2190_ (.Y(_1343_),
    .A(net903));
 sg13g2_inv_1 _2191_ (.Y(_1344_),
    .A(net322));
 sg13g2_inv_1 _2192_ (.Y(_1345_),
    .A(\bitty_inst.d_instr[11] ));
 sg13g2_inv_1 _2193_ (.Y(_1346_),
    .A(net439));
 sg13g2_inv_1 _2194_ (.Y(_1347_),
    .A(\bitty_inst.d_instr[9] ));
 sg13g2_inv_1 _2195_ (.Y(_1348_),
    .A(net402));
 sg13g2_inv_1 _2196_ (.Y(_1349_),
    .A(\bitty_inst.d_instr[7] ));
 sg13g2_inv_1 _2197_ (.Y(_1350_),
    .A(net355));
 sg13g2_inv_1 _2198_ (.Y(_1351_),
    .A(\bitty_inst.d_instr[5] ));
 sg13g2_inv_1 _2199_ (.Y(_1352_),
    .A(net904));
 sg13g2_inv_1 _2200_ (.Y(_1353_),
    .A(\bitty_inst.d_instr[3] ));
 sg13g2_inv_1 _2201_ (.Y(_1354_),
    .A(net449));
 sg13g2_inv_1 _2202_ (.Y(_1355_),
    .A(net801));
 sg13g2_inv_1 _2203_ (.Y(_1356_),
    .A(net940));
 sg13g2_inv_1 _2204_ (.Y(_1357_),
    .A(\bitty_inst.alu_inst.in_a[15] ));
 sg13g2_inv_1 _2205_ (.Y(_1358_),
    .A(\bitty_inst.alu_inst.in_a[10] ));
 sg13g2_inv_1 _2206_ (.Y(_1359_),
    .A(\bitty_inst.alu_inst.in_a[9] ));
 sg13g2_inv_1 _2207_ (.Y(_1360_),
    .A(\bitty_inst.alu_inst.in_a[7] ));
 sg13g2_inv_1 _2208_ (.Y(_1361_),
    .A(\bitty_inst.alu_inst.in_a[6] ));
 sg13g2_inv_1 _2209_ (.Y(_1362_),
    .A(\bitty_inst.alu_inst.in_a[5] ));
 sg13g2_inv_1 _2210_ (.Y(_1363_),
    .A(\bitty_inst.alu_inst.in_a[4] ));
 sg13g2_inv_1 _2211_ (.Y(_1364_),
    .A(\bitty_inst.alu_inst.in_a[1] ));
 sg13g2_inv_1 _2212_ (.Y(_1365_),
    .A(\bitty_inst.alu_inst.in_a[0] ));
 sg13g2_inv_1 _2213_ (.Y(_1366_),
    .A(\bitty_inst.d_out[15] ));
 sg13g2_inv_1 _2214_ (.Y(_1367_),
    .A(net808));
 sg13g2_inv_2 _2215_ (.Y(_1368_),
    .A(net957));
 sg13g2_inv_1 _2216_ (.Y(_1369_),
    .A(\bitty_inst.d_out[13] ));
 sg13g2_inv_2 _2217_ (.Y(_1370_),
    .A(\bitty_inst.d_out[12] ));
 sg13g2_inv_1 _2218_ (.Y(_1371_),
    .A(\bitty_inst.d_out[11] ));
 sg13g2_inv_2 _2219_ (.Y(_1372_),
    .A(net947));
 sg13g2_inv_1 _2220_ (.Y(_1373_),
    .A(\bitty_inst.d_out[9] ));
 sg13g2_inv_2 _2221_ (.Y(_1374_),
    .A(net960));
 sg13g2_inv_1 _2222_ (.Y(_1375_),
    .A(\bitty_inst.d_out[7] ));
 sg13g2_inv_2 _2223_ (.Y(_1376_),
    .A(net963));
 sg13g2_inv_2 _2224_ (.Y(_1377_),
    .A(\bitty_inst.d_out[5] ));
 sg13g2_inv_2 _2225_ (.Y(_1378_),
    .A(net950));
 sg13g2_inv_4 _2226_ (.A(net939),
    .Y(_1379_));
 sg13g2_inv_2 _2227_ (.Y(_1380_),
    .A(net961));
 sg13g2_inv_2 _2228_ (.Y(_1381_),
    .A(\bitty_inst.d_out[1] ));
 sg13g2_inv_2 _2229_ (.Y(_1382_),
    .A(\bitty_inst.d_out[0] ));
 sg13g2_inv_1 _2230_ (.Y(_1383_),
    .A(net384));
 sg13g2_inv_1 _2231_ (.Y(_1384_),
    .A(net356));
 sg13g2_inv_1 _2232_ (.Y(_1385_),
    .A(net323));
 sg13g2_inv_1 _2233_ (.Y(_1386_),
    .A(net380));
 sg13g2_inv_1 _2234_ (.Y(_1387_),
    .A(net376));
 sg13g2_inv_1 _2235_ (.Y(_1388_),
    .A(net374));
 sg13g2_inv_1 _2236_ (.Y(_1389_),
    .A(net343));
 sg13g2_inv_1 _2237_ (.Y(_1390_),
    .A(net351));
 sg13g2_inv_1 _2238_ (.Y(_1391_),
    .A(net327));
 sg13g2_inv_1 _2239_ (.Y(_1392_),
    .A(net362));
 sg13g2_inv_1 _2240_ (.Y(_1393_),
    .A(net337));
 sg13g2_inv_1 _2241_ (.Y(_1394_),
    .A(net428));
 sg13g2_inv_1 _2242_ (.Y(_1395_),
    .A(net335));
 sg13g2_inv_1 _2243_ (.Y(_1396_),
    .A(net349));
 sg13g2_inv_1 _2244_ (.Y(_1397_),
    .A(net414));
 sg13g2_inv_1 _2245_ (.Y(_1398_),
    .A(net432));
 sg13g2_inv_1 _2246_ (.Y(_1399_),
    .A(net368));
 sg13g2_inv_1 _2247_ (.Y(_1400_),
    .A(net378));
 sg13g2_inv_1 _2248_ (.Y(_1401_),
    .A(net341));
 sg13g2_inv_1 _2249_ (.Y(_1402_),
    .A(net392));
 sg13g2_inv_1 _2250_ (.Y(_1403_),
    .A(net394));
 sg13g2_inv_1 _2251_ (.Y(_1404_),
    .A(net347));
 sg13g2_inv_1 _2252_ (.Y(_1405_),
    .A(net331));
 sg13g2_inv_1 _2253_ (.Y(_1406_),
    .A(net404));
 sg13g2_inv_1 _2254_ (.Y(_1407_),
    .A(net358));
 sg13g2_inv_1 _2255_ (.Y(_1408_),
    .A(net390));
 sg13g2_inv_1 _2256_ (.Y(_1409_),
    .A(net372));
 sg13g2_inv_1 _2257_ (.Y(_1410_),
    .A(net396));
 sg13g2_inv_1 _2258_ (.Y(_1411_),
    .A(net333));
 sg13g2_inv_1 _2259_ (.Y(_1412_),
    .A(net370));
 sg13g2_inv_1 _2260_ (.Y(_1413_),
    .A(net416));
 sg13g2_inv_1 _2261_ (.Y(_1414_),
    .A(net408));
 sg13g2_inv_1 _2262_ (.Y(_1415_),
    .A(net353));
 sg13g2_inv_1 _2263_ (.Y(_1416_),
    .A(net329));
 sg13g2_inv_1 _2264_ (.Y(_1417_),
    .A(net400));
 sg13g2_inv_1 _2265_ (.Y(_1418_),
    .A(net382));
 sg13g2_inv_1 _2266_ (.Y(_1419_),
    .A(net366));
 sg13g2_inv_1 _2267_ (.Y(_1420_),
    .A(net437));
 sg13g2_inv_1 _2268_ (.Y(_1421_),
    .A(net345));
 sg13g2_inv_1 _2269_ (.Y(_1422_),
    .A(net360));
 sg13g2_inv_1 _2270_ (.Y(_1423_),
    .A(net388));
 sg13g2_inv_1 _2271_ (.Y(_1424_),
    .A(net386));
 sg13g2_inv_1 _2272_ (.Y(_1425_),
    .A(net339));
 sg13g2_inv_1 _2273_ (.Y(_1426_),
    .A(net406));
 sg13g2_inv_1 _2274_ (.Y(_1427_),
    .A(net398));
 sg13g2_inv_1 _2275_ (.Y(_1428_),
    .A(net364));
 sg13g2_inv_1 _2276_ (.Y(_1429_),
    .A(net426));
 sg13g2_inv_1 _2277_ (.Y(_1430_),
    .A(net410));
 sg13g2_inv_2 _2278_ (.Y(_1431_),
    .A(net814));
 sg13g2_inv_1 _2279_ (.Y(_1432_),
    .A(net942));
 sg13g2_inv_1 _2280_ (.Y(_1433_),
    .A(net895));
 sg13g2_inv_1 _2281_ (.Y(_1434_),
    .A(\uart_inst.R0.bit_counter[2] ));
 sg13g2_inv_1 _2282_ (.Y(_1435_),
    .A(\uart_inst.R0.bit_counter[1] ));
 sg13g2_inv_1 _2283_ (.Y(_1436_),
    .A(net882));
 sg13g2_inv_1 _2284_ (.Y(_1437_),
    .A(\uart_inst.R0.clk_counter[0] ));
 sg13g2_inv_1 _2285_ (.Y(_1438_),
    .A(\uart_inst.T0.bit_counter[2] ));
 sg13g2_inv_1 _2286_ (.Y(_1439_),
    .A(net847));
 sg13g2_inv_1 _2287_ (.Y(_1440_),
    .A(net443));
 sg13g2_inv_2 _2288_ (.Y(_1441_),
    .A(\bitty_inst.lsu_inst.rx_do ));
 sg13g2_inv_1 _2289_ (.Y(_1442_),
    .A(\bitty_inst.cpu_inst.cur_state[1] ));
 sg13g2_inv_1 _2290_ (.Y(_1443_),
    .A(\bitty_inst.lsu_inst.tx_done ));
 sg13g2_inv_1 _2291_ (.Y(_1444_),
    .A(net824));
 sg13g2_inv_1 _2292_ (.Y(_1445_),
    .A(\uart_inst.T0.clk_counter[1] ));
 sg13g2_inv_1 _2293_ (.Y(_1446_),
    .A(net316));
 sg13g2_inv_1 _2294_ (.Y(_1447_),
    .A(\fi_inst.state[1] ));
 sg13g2_inv_1 _2295_ (.Y(_1448_),
    .A(net617));
 sg13g2_inv_1 _2296_ (.Y(_1449_),
    .A(net643));
 sg13g2_inv_1 _2297_ (.Y(_1450_),
    .A(net320));
 sg13g2_inv_2 _2298_ (.Y(_1451_),
    .A(net639));
 sg13g2_inv_1 _2299_ (.Y(_1452_),
    .A(_0033_));
 sg13g2_inv_1 _2300_ (.Y(_1453_),
    .A(_0036_));
 sg13g2_inv_1 _2301_ (.Y(_1454_),
    .A(net805));
 sg13g2_inv_2 _2302_ (.Y(_1455_),
    .A(_0042_));
 sg13g2_inv_2 _2303_ (.Y(_1456_),
    .A(_0044_));
 sg13g2_inv_2 _2304_ (.Y(_1457_),
    .A(_0046_));
 sg13g2_inv_2 _2305_ (.Y(_1458_),
    .A(_0048_));
 sg13g2_inv_1 _2306_ (.Y(_1459_),
    .A(\bitty_inst.data_to_ld[5] ));
 sg13g2_nand2b_2 _2307_ (.Y(_1460_),
    .B(net833),
    .A_N(net812));
 sg13g2_a22oi_1 _2308_ (.Y(_1461_),
    .B1(_1441_),
    .B2(net441),
    .A2(\fi_inst.state[2] ),
    .A1(_1440_));
 sg13g2_nor2_1 _2309_ (.A(_1460_),
    .B(net444),
    .Y(_0018_));
 sg13g2_nor2_1 _2310_ (.A(net819),
    .B(net483),
    .Y(_1462_));
 sg13g2_nand2_1 _2311_ (.Y(_1463_),
    .A(net434),
    .B(_1462_));
 sg13g2_nand2_1 _2312_ (.Y(_1464_),
    .A(\bitty_inst.d_instr[1] ),
    .B(\bitty_inst.d_instr[0] ));
 sg13g2_nand3_1 _2313_ (.B(\bitty_inst.cpu_inst.run ),
    .C(_1464_),
    .A(net828),
    .Y(_1465_));
 sg13g2_nand2_1 _2314_ (.Y(_0012_),
    .A(net435),
    .B(_1465_));
 sg13g2_a21oi_1 _2315_ (.A1(_1443_),
    .A2(\fi_inst.state[4] ),
    .Y(_1466_),
    .B1(net318));
 sg13g2_nor2_1 _2316_ (.A(_1460_),
    .B(net319),
    .Y(_0017_));
 sg13g2_xor2_1 _2317_ (.B(_0067_),
    .A(net1),
    .X(_1467_));
 sg13g2_and2_2 _2318_ (.A(net823),
    .B(net825),
    .X(_1468_));
 sg13g2_nand2_1 _2319_ (.Y(_1469_),
    .A(net824),
    .B(net1));
 sg13g2_nor2_1 _2320_ (.A(\uart_inst.T0.clk_counter[7] ),
    .B(net818),
    .Y(_1470_));
 sg13g2_a21oi_1 _2321_ (.A1(\uart_inst.T0.clk_counter[7] ),
    .A2(net818),
    .Y(_1471_),
    .B1(_1467_));
 sg13g2_nand2b_1 _2322_ (.Y(_1472_),
    .B(_1471_),
    .A_N(_1470_));
 sg13g2_nor2_2 _2323_ (.A(net824),
    .B(net825),
    .Y(_1473_));
 sg13g2_or2_2 _2324_ (.X(_1474_),
    .B(net825),
    .A(net824));
 sg13g2_nand2_2 _2325_ (.Y(_1475_),
    .A(_1469_),
    .B(_1474_));
 sg13g2_nor2_1 _2326_ (.A(_0068_),
    .B(net795),
    .Y(_1476_));
 sg13g2_a22oi_1 _2327_ (.Y(_1477_),
    .B1(_1475_),
    .B2(_0068_),
    .A2(net817),
    .A1(\uart_inst.T0.clk_counter[5] ));
 sg13g2_o21ai_1 _2328_ (.B1(_1477_),
    .Y(_1478_),
    .A1(\uart_inst.T0.clk_counter[5] ),
    .A2(_1473_));
 sg13g2_or3_1 _2329_ (.A(_1472_),
    .B(_1476_),
    .C(_1478_),
    .X(_1479_));
 sg13g2_nand2_2 _2330_ (.Y(_1480_),
    .A(_1444_),
    .B(net825));
 sg13g2_nor2_1 _2331_ (.A(\uart_inst.T0.clk_counter[9] ),
    .B(_1475_),
    .Y(_1481_));
 sg13g2_nand2b_1 _2332_ (.Y(_1482_),
    .B(_1473_),
    .A_N(\uart_inst.T0.clk_counter[12] ));
 sg13g2_o21ai_1 _2333_ (.B1(_1482_),
    .Y(_1483_),
    .A1(\uart_inst.T0.clk_counter[11] ),
    .A2(net794));
 sg13g2_a21oi_1 _2334_ (.A1(\uart_inst.T0.clk_counter[11] ),
    .A2(_1480_),
    .Y(_1484_),
    .B1(_1481_));
 sg13g2_xnor2_1 _2335_ (.Y(_1485_),
    .A(net936),
    .B(_1474_));
 sg13g2_nand3b_1 _2336_ (.B(_1484_),
    .C(_1485_),
    .Y(_1486_),
    .A_N(_1483_));
 sg13g2_xnor2_1 _2337_ (.Y(_1487_),
    .A(_0069_),
    .B(net817));
 sg13g2_and2_1 _2338_ (.A(\uart_inst.T0.clk_counter[3] ),
    .B(_1480_),
    .X(_1488_));
 sg13g2_nor2_1 _2339_ (.A(\uart_inst.T0.clk_counter[3] ),
    .B(net794),
    .Y(_1489_));
 sg13g2_nor3_1 _2340_ (.A(_1487_),
    .B(_1488_),
    .C(_1489_),
    .Y(_1490_));
 sg13g2_nand2_1 _2341_ (.Y(_1491_),
    .A(\uart_inst.T0.clk_counter[12] ),
    .B(_1474_));
 sg13g2_a22oi_1 _2342_ (.Y(_1492_),
    .B1(_1474_),
    .B2(\uart_inst.T0.clk_counter[12] ),
    .A2(_0066_),
    .A1(net824));
 sg13g2_o21ai_1 _2343_ (.B1(_1492_),
    .Y(_1493_),
    .A1(net824),
    .A2(_0066_));
 sg13g2_a21oi_1 _2344_ (.A1(\uart_inst.T0.clk_counter[9] ),
    .A2(_1475_),
    .Y(_1494_),
    .B1(_1493_));
 sg13g2_a21oi_1 _2345_ (.A1(_1445_),
    .A2(net818),
    .Y(_1495_),
    .B1(net316));
 sg13g2_nand2_1 _2346_ (.Y(_1496_),
    .A(\uart_inst.T0.clk_counter[1] ),
    .B(_1468_));
 sg13g2_nand4_1 _2347_ (.B(_1494_),
    .C(_1495_),
    .A(_1490_),
    .Y(_1497_),
    .D(_1496_));
 sg13g2_nor3_2 _2348_ (.A(_1479_),
    .B(_1486_),
    .C(_1497_),
    .Y(_1498_));
 sg13g2_nor2_1 _2349_ (.A(net821),
    .B(_1498_),
    .Y(_1499_));
 sg13g2_nand2_1 _2350_ (.Y(_1500_),
    .A(\uart_inst.T0.bit_counter[1] ),
    .B(net816));
 sg13g2_nor3_1 _2351_ (.A(_1438_),
    .B(net569),
    .C(_1500_),
    .Y(_1501_));
 sg13g2_o21ai_1 _2352_ (.B1(net848),
    .Y(_1502_),
    .A1(net569),
    .A2(net934));
 sg13g2_nor2_1 _2353_ (.A(_1501_),
    .B(_1502_),
    .Y(_1503_));
 sg13g2_a22oi_1 _2354_ (.Y(_1504_),
    .B1(_1503_),
    .B2(_1498_),
    .A2(_1499_),
    .A1(net920));
 sg13g2_inv_1 _2355_ (.Y(_0025_),
    .A(_1504_));
 sg13g2_nand2_2 _2356_ (.Y(_0031_),
    .A(\bitty_inst.lsu_inst.rx_do ),
    .B(\fi_inst.state[1] ));
 sg13g2_nand2_2 _2357_ (.Y(_0032_),
    .A(\bitty_inst.lsu_inst.rx_do ),
    .B(\fi_inst.state[5] ));
 sg13g2_a22oi_1 _2358_ (.Y(_1505_),
    .B1(net497),
    .B2(_1440_),
    .A2(_1443_),
    .A1(\fi_inst.state[2] ));
 sg13g2_nor2_1 _2359_ (.A(_1460_),
    .B(net498),
    .Y(_0016_));
 sg13g2_nor2_1 _2360_ (.A(\fi_inst.state[2] ),
    .B(\fi_inst.state[4] ),
    .Y(_1506_));
 sg13g2_nor3_1 _2361_ (.A(net811),
    .B(\fi_inst.state[2] ),
    .C(\fi_inst.state[4] ),
    .Y(_1507_));
 sg13g2_nor2b_1 _2362_ (.A(\bitty_inst.lsu_inst.state[1] ),
    .B_N(\bitty_inst.lsu_inst.state[0] ),
    .Y(_1508_));
 sg13g2_nand2_2 _2363_ (.Y(_1509_),
    .A(_0072_),
    .B(_1508_));
 sg13g2_nand3b_1 _2364_ (.B(\bitty_inst.lsu_inst.state[1] ),
    .C(_0072_),
    .Y(_1510_),
    .A_N(\bitty_inst.lsu_inst.state[0] ));
 sg13g2_nand2_1 _2365_ (.Y(_1511_),
    .A(_1509_),
    .B(_1510_));
 sg13g2_nor2_2 _2366_ (.A(net798),
    .B(_0035_),
    .Y(_1512_));
 sg13g2_nand2b_2 _2367_ (.Y(_1513_),
    .B(net808),
    .A_N(_0035_));
 sg13g2_nand2_1 _2368_ (.Y(_1514_),
    .A(net801),
    .B(\bitty_inst.cpu_inst.d_inst[0] ));
 sg13g2_nand3_1 _2369_ (.B(net801),
    .C(\bitty_inst.cpu_inst.d_inst[0] ),
    .A(\bitty_inst.cpu_inst.d_inst[2] ),
    .Y(_1515_));
 sg13g2_or2_1 _2370_ (.X(_1516_),
    .B(_1515_),
    .A(_1513_));
 sg13g2_nand3_1 _2371_ (.B(\bitty_inst.cpu_inst.d_inst[0] ),
    .C(_0035_),
    .A(net801),
    .Y(_1517_));
 sg13g2_or2_1 _2372_ (.X(_1518_),
    .B(_1517_),
    .A(net798));
 sg13g2_o21ai_1 _2373_ (.B1(_1516_),
    .Y(_1519_),
    .A1(\bitty_inst.cpu_inst.d_inst[2] ),
    .A2(_1518_));
 sg13g2_nand2_1 _2374_ (.Y(_1520_),
    .A(\bitty_inst.lsu_inst.state[2] ),
    .B(_1508_));
 sg13g2_nor2b_1 _2375_ (.A(\bitty_inst.lsu_inst.state[0] ),
    .B_N(\bitty_inst.lsu_inst.state[2] ),
    .Y(_1521_));
 sg13g2_and2_2 _2376_ (.A(\bitty_inst.lsu_inst.state[1] ),
    .B(_1521_),
    .X(_1522_));
 sg13g2_a21oi_1 _2377_ (.A1(\bitty_inst.lsu_inst.state[2] ),
    .A2(_1508_),
    .Y(_1523_),
    .B1(net788));
 sg13g2_o21ai_1 _2378_ (.B1(net811),
    .Y(_1524_),
    .A1(_1511_),
    .A2(_1523_));
 sg13g2_a21oi_1 _2379_ (.A1(_1511_),
    .A2(_1519_),
    .Y(_1525_),
    .B1(_1524_));
 sg13g2_nand2_1 _2380_ (.Y(_1526_),
    .A(net845),
    .B(net471));
 sg13g2_nor3_2 _2381_ (.A(_1507_),
    .B(_1525_),
    .C(_1526_),
    .Y(_1527_));
 sg13g2_a21o_1 _2382_ (.A2(_1499_),
    .A1(net569),
    .B1(_1527_),
    .X(_0026_));
 sg13g2_o21ai_1 _2383_ (.B1(net483),
    .Y(_1528_),
    .A1(\cur_state[7] ),
    .A2(net434));
 sg13g2_nand2b_1 _2384_ (.Y(_1529_),
    .B(net325),
    .A_N(fetch_done));
 sg13g2_nand3_1 _2385_ (.B(net484),
    .C(_1529_),
    .A(net830),
    .Y(_0011_));
 sg13g2_nand2_1 _2386_ (.Y(_1530_),
    .A(net421),
    .B(_1499_));
 sg13g2_nand4_1 _2387_ (.B(\uart_inst.T0.bit_counter[1] ),
    .C(net816),
    .A(\uart_inst.T0.bit_counter[2] ),
    .Y(_1531_),
    .D(\uart_inst.T0.PS[1] ));
 sg13g2_nand2_1 _2388_ (.Y(_1532_),
    .A(net847),
    .B(_1498_));
 sg13g2_o21ai_1 _2389_ (.B1(_1530_),
    .Y(_0027_),
    .A1(_1531_),
    .A2(_1532_));
 sg13g2_a22oi_1 _2390_ (.Y(_1533_),
    .B1(_1450_),
    .B2(net441),
    .A2(\fi_inst.state[1] ),
    .A1(_1441_));
 sg13g2_nor2_1 _2391_ (.A(_1460_),
    .B(net442),
    .Y(_0015_));
 sg13g2_or2_1 _2392_ (.X(_0014_),
    .B(_1460_),
    .A(net645));
 sg13g2_nand2_1 _2393_ (.Y(_1534_),
    .A(net609),
    .B(_1462_));
 sg13g2_nand4_1 _2394_ (.B(\bitty_inst.d_instr[0] ),
    .C(net828),
    .A(\bitty_inst.d_instr[1] ),
    .Y(_1535_),
    .D(net503));
 sg13g2_nand2_1 _2395_ (.Y(_0013_),
    .A(_1534_),
    .B(_1535_));
 sg13g2_o21ai_1 _2396_ (.B1(net471),
    .Y(_1536_),
    .A1(_1507_),
    .A2(_1525_));
 sg13g2_nand3_1 _2397_ (.B(_1443_),
    .C(_1536_),
    .A(net833),
    .Y(_0024_));
 sg13g2_nor2_1 _2398_ (.A(net820),
    .B(net827),
    .Y(_1537_));
 sg13g2_xor2_1 _2399_ (.B(_0059_),
    .A(net825),
    .X(_1538_));
 sg13g2_xnor2_1 _2400_ (.Y(_1539_),
    .A(\uart_inst.R0.clk_counter[7] ),
    .B(net818));
 sg13g2_nor2_1 _2401_ (.A(_1538_),
    .B(_1539_),
    .Y(_1540_));
 sg13g2_xnor2_1 _2402_ (.Y(_1541_),
    .A(_0060_),
    .B(net817));
 sg13g2_xor2_1 _2403_ (.B(net795),
    .A(_0061_),
    .X(_1542_));
 sg13g2_nand3_1 _2404_ (.B(_1541_),
    .C(_1542_),
    .A(_1540_),
    .Y(_1543_));
 sg13g2_xor2_1 _2405_ (.B(net795),
    .A(_0057_),
    .X(_1544_));
 sg13g2_nor2_1 _2406_ (.A(\uart_inst.R0.clk_counter[11] ),
    .B(net824),
    .Y(_1545_));
 sg13g2_nor2_1 _2407_ (.A(net825),
    .B(_0056_),
    .Y(_1546_));
 sg13g2_mux2_1 _2408_ (.A0(_0056_),
    .A1(_1546_),
    .S(_1545_),
    .X(_1547_));
 sg13g2_xnor2_1 _2409_ (.Y(_1548_),
    .A(_0055_),
    .B(net817));
 sg13g2_inv_1 _2410_ (.Y(_1549_),
    .A(_1548_));
 sg13g2_xnor2_1 _2411_ (.Y(_1550_),
    .A(net823),
    .B(_0058_));
 sg13g2_a21oi_1 _2412_ (.A1(\uart_inst.R0.clk_counter[11] ),
    .A2(net794),
    .Y(_1551_),
    .B1(_1550_));
 sg13g2_nand3_1 _2413_ (.B(_1549_),
    .C(_1551_),
    .A(_1547_),
    .Y(_1552_));
 sg13g2_or2_1 _2414_ (.X(_1553_),
    .B(_1552_),
    .A(_1544_));
 sg13g2_nand2_1 _2415_ (.Y(_1554_),
    .A(\uart_inst.R0.clk_counter[1] ),
    .B(_1468_));
 sg13g2_o21ai_1 _2416_ (.B1(_0063_),
    .Y(_1555_),
    .A1(\uart_inst.R0.clk_counter[3] ),
    .A2(net823));
 sg13g2_a21oi_1 _2417_ (.A1(\uart_inst.R0.clk_counter[3] ),
    .A2(net794),
    .Y(_1556_),
    .B1(_1555_));
 sg13g2_nor2_1 _2418_ (.A(\uart_inst.R0.clk_counter[3] ),
    .B(_0063_),
    .Y(_1557_));
 sg13g2_a21oi_1 _2419_ (.A1(net817),
    .A2(_1557_),
    .Y(_1558_),
    .B1(_1556_));
 sg13g2_nand2_1 _2420_ (.Y(_1559_),
    .A(\uart_inst.R0.clk_counter[1] ),
    .B(\uart_inst.R0.clk_counter[0] ));
 sg13g2_o21ai_1 _2421_ (.B1(\uart_inst.R0.clk_counter[0] ),
    .Y(_1560_),
    .A1(\uart_inst.R0.clk_counter[1] ),
    .A2(_1468_));
 sg13g2_a21o_1 _2422_ (.A2(_1468_),
    .A1(\uart_inst.R0.clk_counter[1] ),
    .B1(_1560_),
    .X(_1561_));
 sg13g2_nor4_2 _2423_ (.A(_1543_),
    .B(_1553_),
    .C(_1558_),
    .Y(_1562_),
    .D(_1561_));
 sg13g2_a21o_1 _2424_ (.A2(_1562_),
    .A1(net617),
    .B1(net910),
    .X(_1563_));
 sg13g2_nor2_1 _2425_ (.A(\uart_inst.R0.clk_counter[9] ),
    .B(_0061_),
    .Y(_1564_));
 sg13g2_a21oi_1 _2426_ (.A1(\uart_inst.R0.clk_counter[11] ),
    .A2(net817),
    .Y(_1565_),
    .B1(_1564_));
 sg13g2_nand3_1 _2427_ (.B(net823),
    .C(_0063_),
    .A(\uart_inst.R0.clk_counter[7] ),
    .Y(_1566_));
 sg13g2_or3_1 _2428_ (.A(\uart_inst.R0.clk_counter[7] ),
    .B(net823),
    .C(_0063_),
    .X(_1567_));
 sg13g2_or3_1 _2429_ (.A(\uart_inst.R0.clk_counter[8] ),
    .B(\uart_inst.R0.clk_counter[1] ),
    .C(_0062_),
    .X(_1568_));
 sg13g2_and3_1 _2430_ (.X(_1569_),
    .A(\uart_inst.R0.clk_counter[8] ),
    .B(\uart_inst.R0.clk_counter[1] ),
    .C(_0062_));
 sg13g2_xor2_1 _2431_ (.B(_0060_),
    .A(net825),
    .X(_1570_));
 sg13g2_nor2_1 _2432_ (.A(\uart_inst.R0.clk_counter[10] ),
    .B(net794),
    .Y(_1571_));
 sg13g2_a21oi_1 _2433_ (.A1(\uart_inst.R0.clk_counter[6] ),
    .A2(net818),
    .Y(_1572_),
    .B1(_1571_));
 sg13g2_nand2_1 _2434_ (.Y(_1573_),
    .A(\uart_inst.R0.clk_counter[9] ),
    .B(_0061_));
 sg13g2_o21ai_1 _2435_ (.B1(_1573_),
    .Y(_1574_),
    .A1(\uart_inst.R0.clk_counter[11] ),
    .A2(net817));
 sg13g2_a22oi_1 _2436_ (.Y(_1575_),
    .B1(net794),
    .B2(\uart_inst.R0.clk_counter[10] ),
    .A2(_1468_),
    .A1(_0064_));
 sg13g2_and2_1 _2437_ (.A(\uart_inst.R0.clk_counter[6] ),
    .B(net825),
    .X(_1576_));
 sg13g2_a21oi_1 _2438_ (.A1(net823),
    .A2(_1576_),
    .Y(_1577_),
    .B1(_0064_));
 sg13g2_o21ai_1 _2439_ (.B1(_1574_),
    .Y(_1578_),
    .A1(net795),
    .A2(_1569_));
 sg13g2_nor4_1 _2440_ (.A(\uart_inst.R0.clk_counter[12] ),
    .B(_1565_),
    .C(_1570_),
    .D(_1578_),
    .Y(_1579_));
 sg13g2_a221oi_1 _2441_ (.B2(net795),
    .C1(_1577_),
    .B1(_1568_),
    .A1(_1566_),
    .Y(_1580_),
    .A2(_1567_));
 sg13g2_and4_2 _2442_ (.A(_1572_),
    .B(_1575_),
    .C(_1579_),
    .D(_1580_),
    .X(_1581_));
 sg13g2_and2_1 _2443_ (.A(net643),
    .B(_1581_),
    .X(_1582_));
 sg13g2_nand2_2 _2444_ (.Y(_1583_),
    .A(net827),
    .B(_1582_));
 sg13g2_nor2_1 _2445_ (.A(net820),
    .B(_1583_),
    .Y(_1584_));
 sg13g2_a21o_1 _2446_ (.A2(_1563_),
    .A1(_1537_),
    .B1(net655),
    .X(_0021_));
 sg13g2_nor2_2 _2447_ (.A(_1449_),
    .B(_1581_),
    .Y(_1585_));
 sg13g2_a22oi_1 _2448_ (.Y(_1586_),
    .B1(_1585_),
    .B2(net845),
    .A2(_1537_),
    .A1(net596));
 sg13g2_inv_1 _2449_ (.Y(_0022_),
    .A(net597));
 sg13g2_nand2_2 _2450_ (.Y(_1587_),
    .A(\uart_inst.R0.bit_counter[1] ),
    .B(\uart_inst.R0.bit_counter[0] ));
 sg13g2_nor2_1 _2451_ (.A(net796),
    .B(_1587_),
    .Y(_1588_));
 sg13g2_nand2_1 _2452_ (.Y(_1589_),
    .A(net886),
    .B(_1588_));
 sg13g2_nand2_1 _2453_ (.Y(_1590_),
    .A(_1562_),
    .B(_1589_));
 sg13g2_o21ai_1 _2454_ (.B1(_1590_),
    .Y(_1591_),
    .A1(net617),
    .A2(_1562_));
 sg13g2_nor2_1 _2455_ (.A(net820),
    .B(_1591_),
    .Y(_0023_));
 sg13g2_nand2_1 _2456_ (.Y(_1592_),
    .A(net807),
    .B(net828));
 sg13g2_nand3_1 _2457_ (.B(\bitty_inst.lsu_inst.state[0] ),
    .C(\bitty_inst.lsu_inst.state[1] ),
    .A(\bitty_inst.lsu_inst.state[2] ),
    .Y(_1593_));
 sg13g2_nand2b_2 _2458_ (.Y(_1594_),
    .B(_1593_),
    .A_N(_1514_));
 sg13g2_nor2b_2 _2459_ (.A(\bitty_inst.cpu_inst.d_inst[0] ),
    .B_N(\bitty_inst.cpu_inst.d_inst[1] ),
    .Y(_1595_));
 sg13g2_nand2b_1 _2460_ (.Y(_1596_),
    .B(net801),
    .A_N(\bitty_inst.cpu_inst.d_inst[0] ));
 sg13g2_nor2_1 _2461_ (.A(_1451_),
    .B(_1595_),
    .Y(_1597_));
 sg13g2_nand3_1 _2462_ (.B(net503),
    .C(net783),
    .A(net828),
    .Y(_1598_));
 sg13g2_o21ai_1 _2463_ (.B1(_1598_),
    .Y(_0010_),
    .A1(_1592_),
    .A2(_1594_));
 sg13g2_o21ai_1 _2464_ (.B1(_1462_),
    .Y(_0008_),
    .A1(net503),
    .A2(_1451_));
 sg13g2_o21ai_1 _2465_ (.B1(net826),
    .Y(_1599_),
    .A1(net910),
    .A2(net596));
 sg13g2_nand3_1 _2466_ (.B(_1441_),
    .C(_1599_),
    .A(net845),
    .Y(_0019_));
 sg13g2_and2_2 _2467_ (.A(net846),
    .B(\uart_inst.R0.PS[1] ),
    .X(_1600_));
 sg13g2_nand2_2 _2468_ (.Y(_1601_),
    .A(net845),
    .B(net886));
 sg13g2_a21oi_1 _2469_ (.A1(_1562_),
    .A2(_1588_),
    .Y(_1602_),
    .B1(_1601_));
 sg13g2_a21o_1 _2470_ (.A2(_1582_),
    .A1(_1537_),
    .B1(_1602_),
    .X(_0020_));
 sg13g2_nand2b_1 _2471_ (.Y(_1603_),
    .B(_1594_),
    .A_N(_1592_));
 sg13g2_nand3_1 _2472_ (.B(net503),
    .C(_1595_),
    .A(net828),
    .Y(_1604_));
 sg13g2_o21ai_1 _2473_ (.B1(_1603_),
    .Y(_0009_),
    .A1(_1451_),
    .A2(_1604_));
 sg13g2_nor2b_2 _2474_ (.A(\bitty_inst.lsu_inst.state[1] ),
    .B_N(_1521_),
    .Y(_1605_));
 sg13g2_inv_1 _2475_ (.Y(_1606_),
    .A(_1605_));
 sg13g2_nand2_2 _2476_ (.Y(_0030_),
    .A(\bitty_inst.lsu_inst.rx_do ),
    .B(_1605_));
 sg13g2_nand3_1 _2477_ (.B(\bitty_inst.lsu_inst.state[1] ),
    .C(_0072_),
    .A(\bitty_inst.lsu_inst.state[0] ),
    .Y(_1607_));
 sg13g2_or2_1 _2478_ (.X(_0029_),
    .B(_1607_),
    .A(_1441_));
 sg13g2_a21oi_1 _2479_ (.A1(_1515_),
    .A2(_1517_),
    .Y(_1608_),
    .B1(net798));
 sg13g2_nand2_1 _2480_ (.Y(_1609_),
    .A(\bitty_inst.lsu_inst.tx_done ),
    .B(_1608_));
 sg13g2_nand2b_1 _2481_ (.Y(_1610_),
    .B(_1609_),
    .A_N(_1509_));
 sg13g2_a21o_1 _2482_ (.A2(\bitty_inst.lsu_inst.state[1] ),
    .A1(\bitty_inst.lsu_inst.state[0] ),
    .B1(\bitty_inst.lsu_inst.state[2] ),
    .X(_1611_));
 sg13g2_a21oi_1 _2483_ (.A1(_1593_),
    .A2(_1611_),
    .Y(_1612_),
    .B1(_1511_));
 sg13g2_nand2_1 _2484_ (.Y(_1613_),
    .A(\bitty_inst.lsu_inst.tx_done ),
    .B(net788));
 sg13g2_o21ai_1 _2485_ (.B1(_1613_),
    .Y(_1614_),
    .A1(\bitty_inst.lsu_inst.tx_done ),
    .A2(net789));
 sg13g2_nor2_1 _2486_ (.A(_1510_),
    .B(_1516_),
    .Y(_1615_));
 sg13g2_o21ai_1 _2487_ (.B1(_1607_),
    .Y(_1616_),
    .A1(_0073_),
    .A2(_1606_));
 sg13g2_nor4_1 _2488_ (.A(_1612_),
    .B(_1614_),
    .C(_1615_),
    .D(_1616_),
    .Y(_1617_));
 sg13g2_nand2_1 _2489_ (.Y(_0304_),
    .A(_1610_),
    .B(_1617_));
 sg13g2_nor2_1 _2490_ (.A(_1509_),
    .B(_1609_),
    .Y(_1618_));
 sg13g2_nor2_1 _2491_ (.A(_0075_),
    .B(net789),
    .Y(_1619_));
 sg13g2_or2_1 _2492_ (.X(_1620_),
    .B(_1519_),
    .A(_1510_));
 sg13g2_nor4_1 _2493_ (.A(net788),
    .B(_1616_),
    .C(_1618_),
    .D(_1619_),
    .Y(_1621_));
 sg13g2_a21oi_1 _2494_ (.A1(_1620_),
    .A2(_1621_),
    .Y(_0305_),
    .B1(_1612_));
 sg13g2_nand2b_1 _2495_ (.Y(_1622_),
    .B(_1519_),
    .A_N(_1510_));
 sg13g2_inv_1 _2496_ (.Y(_1623_),
    .A(_1622_));
 sg13g2_nand2_1 _2497_ (.Y(_1624_),
    .A(_1523_),
    .B(_0029_));
 sg13g2_a21oi_1 _2498_ (.A1(_1441_),
    .A2(_1605_),
    .Y(_1625_),
    .B1(_1624_));
 sg13g2_a21oi_1 _2499_ (.A1(net729),
    .A2(_1625_),
    .Y(_0306_),
    .B1(_1612_));
 sg13g2_and2_1 _2500_ (.A(net830),
    .B(net317),
    .X(_0001_));
 sg13g2_nor3_1 _2501_ (.A(_1447_),
    .B(net320),
    .C(_1460_),
    .Y(_0005_));
 sg13g2_and3_1 _2502_ (.X(_0000_),
    .A(net814),
    .B(net830),
    .C(_1464_));
 sg13g2_and3_1 _2503_ (.X(_0007_),
    .A(net847),
    .B(net421),
    .C(_1498_));
 sg13g2_and4_1 _2504_ (.A(net846),
    .B(net617),
    .C(net826),
    .D(_1562_),
    .X(_0006_));
 sg13g2_and3_1 _2505_ (.X(_0002_),
    .A(net830),
    .B(fetch_done),
    .C(net325));
 sg13g2_nor2_1 _2506_ (.A(\bitty_inst.lsu_inst.tx_done ),
    .B(_1510_),
    .Y(_0028_));
 sg13g2_nor3_1 _2507_ (.A(_1431_),
    .B(net819),
    .C(_1464_),
    .Y(_0004_));
 sg13g2_o21ai_1 _2508_ (.B1(net830),
    .Y(_1626_),
    .A1(\cur_state[6] ),
    .A2(net447));
 sg13g2_inv_1 _2509_ (.Y(_0003_),
    .A(net448));
 sg13g2_nand2b_1 _2510_ (.Y(_0201_),
    .B(net845),
    .A_N(\bitty_inst.lsu_inst.next_state[0] ));
 sg13g2_and2_1 _2511_ (.A(net845),
    .B(\bitty_inst.lsu_inst.next_state[1] ),
    .X(_0202_));
 sg13g2_and2_1 _2512_ (.A(net845),
    .B(\bitty_inst.lsu_inst.next_state[2] ),
    .X(_0203_));
 sg13g2_a22oi_1 _2513_ (.Y(_1627_),
    .B1(net795),
    .B2(\uart_inst.T0.clk_counter[9] ),
    .A2(\uart_inst.T0.clk_counter[8] ),
    .A1(_1444_));
 sg13g2_nand2b_1 _2514_ (.Y(_1628_),
    .B(_1496_),
    .A_N(_1495_));
 sg13g2_nand3b_1 _2515_ (.B(\uart_inst.T0.clk_counter[2] ),
    .C(_1474_),
    .Y(_1629_),
    .A_N(_1489_));
 sg13g2_a21oi_1 _2516_ (.A1(_1490_),
    .A2(_1628_),
    .Y(_1630_),
    .B1(_1488_));
 sg13g2_a21oi_1 _2517_ (.A1(_1629_),
    .A2(_1630_),
    .Y(_1631_),
    .B1(_1479_));
 sg13g2_a22oi_1 _2518_ (.Y(_1632_),
    .B1(net818),
    .B2(\uart_inst.T0.clk_counter[7] ),
    .A2(\uart_inst.T0.clk_counter[6] ),
    .A1(net1));
 sg13g2_or2_1 _2519_ (.X(_1633_),
    .B(_1632_),
    .A(_1470_));
 sg13g2_o21ai_1 _2520_ (.B1(\uart_inst.T0.clk_counter[5] ),
    .Y(_1634_),
    .A1(_1473_),
    .A2(_1476_));
 sg13g2_o21ai_1 _2521_ (.B1(_1633_),
    .Y(_1635_),
    .A1(_1472_),
    .A2(_1634_));
 sg13g2_o21ai_1 _2522_ (.B1(_1494_),
    .Y(_1636_),
    .A1(_1631_),
    .A2(_1635_));
 sg13g2_a21o_1 _2523_ (.A2(_1636_),
    .A1(_1627_),
    .B1(_1486_),
    .X(_1637_));
 sg13g2_a22oi_1 _2524_ (.Y(_1638_),
    .B1(_1480_),
    .B2(\uart_inst.T0.clk_counter[11] ),
    .A2(_1474_),
    .A1(\uart_inst.T0.clk_counter[10] ));
 sg13g2_o21ai_1 _2525_ (.B1(_1491_),
    .Y(_1639_),
    .A1(_1483_),
    .A2(_1638_));
 sg13g2_nor2b_1 _2526_ (.A(_1639_),
    .B_N(_1637_),
    .Y(_1640_));
 sg13g2_a21oi_1 _2527_ (.A1(\uart_inst.T0.PS[1] ),
    .A2(_1640_),
    .Y(_1641_),
    .B1(\uart_inst.T0.PS[2] ));
 sg13g2_nand2b_1 _2528_ (.Y(_1642_),
    .B(_1641_),
    .A_N(\uart_inst.T0.PS[4] ));
 sg13g2_nor2b_2 _2529_ (.A(_1642_),
    .B_N(_1531_),
    .Y(_1643_));
 sg13g2_a21oi_1 _2530_ (.A1(net920),
    .A2(_1643_),
    .Y(_1644_),
    .B1(net816));
 sg13g2_a21oi_1 _2531_ (.A1(net816),
    .A2(_1643_),
    .Y(_1645_),
    .B1(net820));
 sg13g2_nor2b_1 _2532_ (.A(net921),
    .B_N(_1645_),
    .Y(_0204_));
 sg13g2_a21oi_1 _2533_ (.A1(net816),
    .A2(_1643_),
    .Y(_1646_),
    .B1(net887));
 sg13g2_nand2_1 _2534_ (.Y(_1647_),
    .A(\uart_inst.T0.PS[1] ),
    .B(_1500_));
 sg13g2_a21oi_1 _2535_ (.A1(_1643_),
    .A2(_1647_),
    .Y(_1648_),
    .B1(net820));
 sg13g2_nor2b_1 _2536_ (.A(net888),
    .B_N(_1648_),
    .Y(_0205_));
 sg13g2_nand2b_1 _2537_ (.Y(_1649_),
    .B(\uart_inst.T0.bit_counter[2] ),
    .A_N(_1643_));
 sg13g2_xor2_1 _2538_ (.B(_1500_),
    .A(net648),
    .X(_1650_));
 sg13g2_nand3_1 _2539_ (.B(_1643_),
    .C(_1650_),
    .A(\uart_inst.T0.PS[1] ),
    .Y(_1651_));
 sg13g2_a21oi_1 _2540_ (.A1(_1649_),
    .A2(net649),
    .Y(_0206_),
    .B1(net820));
 sg13g2_nand3_1 _2541_ (.B(_1640_),
    .C(_1642_),
    .A(net848),
    .Y(_1652_));
 sg13g2_nor2_1 _2542_ (.A(_1446_),
    .B(net654),
    .Y(_0207_));
 sg13g2_xnor2_1 _2543_ (.Y(_1653_),
    .A(net873),
    .B(\uart_inst.T0.clk_counter[1] ));
 sg13g2_nor2_1 _2544_ (.A(net654),
    .B(net874),
    .Y(_0208_));
 sg13g2_and3_1 _2545_ (.X(_1654_),
    .A(\uart_inst.T0.clk_counter[0] ),
    .B(\uart_inst.T0.clk_counter[1] ),
    .C(net418));
 sg13g2_a21oi_1 _2546_ (.A1(\uart_inst.T0.clk_counter[0] ),
    .A2(\uart_inst.T0.clk_counter[1] ),
    .Y(_1655_),
    .B1(net418));
 sg13g2_nor3_1 _2547_ (.A(net654),
    .B(_1654_),
    .C(net419),
    .Y(_0209_));
 sg13g2_nand3b_1 _2548_ (.B(\uart_inst.T0.clk_counter[1] ),
    .C(net873),
    .Y(_1656_),
    .A_N(net533));
 sg13g2_xor2_1 _2549_ (.B(_1656_),
    .A(net912),
    .X(_1657_));
 sg13g2_nor2_1 _2550_ (.A(net653),
    .B(net913),
    .Y(_0210_));
 sg13g2_and3_1 _2551_ (.X(_1658_),
    .A(net964),
    .B(net412),
    .C(_1654_));
 sg13g2_a21oi_1 _2552_ (.A1(\uart_inst.T0.clk_counter[3] ),
    .A2(_1654_),
    .Y(_1659_),
    .B1(net412));
 sg13g2_nor3_1 _2553_ (.A(net654),
    .B(_1658_),
    .C(net413),
    .Y(_0211_));
 sg13g2_nand3b_1 _2554_ (.B(_1654_),
    .C(net912),
    .Y(_1660_),
    .A_N(_0068_));
 sg13g2_xor2_1 _2555_ (.B(_1660_),
    .A(net917),
    .X(_1661_));
 sg13g2_nor2_1 _2556_ (.A(net653),
    .B(net918),
    .Y(_0212_));
 sg13g2_and3_1 _2557_ (.X(_1662_),
    .A(net423),
    .B(\uart_inst.T0.clk_counter[5] ),
    .C(_1658_));
 sg13g2_a21oi_1 _2558_ (.A1(\uart_inst.T0.clk_counter[5] ),
    .A2(_1658_),
    .Y(_1663_),
    .B1(net423));
 sg13g2_nor3_1 _2559_ (.A(net654),
    .B(_1662_),
    .C(net424),
    .Y(_0213_));
 sg13g2_nand3b_1 _2560_ (.B(\uart_inst.T0.clk_counter[5] ),
    .C(_1658_),
    .Y(_1664_),
    .A_N(_0067_));
 sg13g2_xor2_1 _2561_ (.B(_1664_),
    .A(net880),
    .X(_1665_));
 sg13g2_nor2_1 _2562_ (.A(net653),
    .B(net881),
    .Y(_0214_));
 sg13g2_and2_1 _2563_ (.A(\uart_inst.T0.clk_counter[7] ),
    .B(_1662_),
    .X(_1666_));
 sg13g2_nor2_1 _2564_ (.A(net454),
    .B(_1666_),
    .Y(_1667_));
 sg13g2_and2_1 _2565_ (.A(net454),
    .B(_1666_),
    .X(_1668_));
 sg13g2_nor3_1 _2566_ (.A(net653),
    .B(net455),
    .C(_1668_),
    .Y(_0215_));
 sg13g2_nor2b_1 _2567_ (.A(net637),
    .B_N(_1666_),
    .Y(_1669_));
 sg13g2_xnor2_1 _2568_ (.Y(_1670_),
    .A(\uart_inst.T0.clk_counter[9] ),
    .B(_1669_));
 sg13g2_nor2_1 _2569_ (.A(net653),
    .B(net638),
    .Y(_0216_));
 sg13g2_nand2_1 _2570_ (.Y(_1671_),
    .A(\uart_inst.T0.clk_counter[9] ),
    .B(_1668_));
 sg13g2_xor2_1 _2571_ (.B(_1671_),
    .A(net877),
    .X(_1672_));
 sg13g2_nor2_1 _2572_ (.A(net653),
    .B(net878),
    .Y(_0217_));
 sg13g2_nor2_1 _2573_ (.A(net651),
    .B(_1671_),
    .Y(_1673_));
 sg13g2_xnor2_1 _2574_ (.Y(_1674_),
    .A(\uart_inst.T0.clk_counter[11] ),
    .B(net863));
 sg13g2_nor2_1 _2575_ (.A(net653),
    .B(net864),
    .Y(_0218_));
 sg13g2_nand4_1 _2576_ (.B(net877),
    .C(\uart_inst.T0.clk_counter[9] ),
    .A(\uart_inst.T0.clk_counter[11] ),
    .Y(_1675_),
    .D(_1668_));
 sg13g2_xor2_1 _2577_ (.B(_1675_),
    .A(net890),
    .X(_1676_));
 sg13g2_nor2_1 _2578_ (.A(net653),
    .B(net891),
    .Y(_0219_));
 sg13g2_a21o_1 _2579_ (.A2(net794),
    .A1(\uart_inst.R0.clk_counter[3] ),
    .B1(\uart_inst.R0.clk_counter[2] ),
    .X(_1677_));
 sg13g2_o21ai_1 _2580_ (.B1(_1677_),
    .Y(_1678_),
    .A1(\uart_inst.R0.clk_counter[3] ),
    .A2(net823));
 sg13g2_a21o_1 _2581_ (.A2(_1560_),
    .A1(_1554_),
    .B1(_1558_),
    .X(_1679_));
 sg13g2_a21oi_1 _2582_ (.A1(_1678_),
    .A2(_1679_),
    .Y(_1680_),
    .B1(_1543_));
 sg13g2_nor3_1 _2583_ (.A(_0060_),
    .B(_0061_),
    .C(net795),
    .Y(_1681_));
 sg13g2_a21o_1 _2584_ (.A2(net817),
    .A1(\uart_inst.R0.clk_counter[5] ),
    .B1(_1681_),
    .X(_1682_));
 sg13g2_o21ai_1 _2585_ (.B1(_1576_),
    .Y(_1683_),
    .A1(\uart_inst.R0.clk_counter[7] ),
    .A2(net818));
 sg13g2_a221oi_1 _2586_ (.B2(_1682_),
    .C1(_1680_),
    .B1(_1540_),
    .A1(\uart_inst.R0.clk_counter[7] ),
    .Y(_0307_),
    .A2(net818));
 sg13g2_a21oi_1 _2587_ (.A1(_1683_),
    .A2(_0307_),
    .Y(_0308_),
    .B1(_1553_));
 sg13g2_nor3_1 _2588_ (.A(net823),
    .B(_0058_),
    .C(_1544_),
    .Y(_0309_));
 sg13g2_and2_1 _2589_ (.A(\uart_inst.R0.clk_counter[9] ),
    .B(net795),
    .X(_0310_));
 sg13g2_o21ai_1 _2590_ (.B1(_1547_),
    .Y(_0311_),
    .A1(_0309_),
    .A2(_0310_));
 sg13g2_a21oi_1 _2591_ (.A1(\uart_inst.R0.clk_counter[11] ),
    .A2(net794),
    .Y(_0312_),
    .B1(\uart_inst.R0.clk_counter[10] ));
 sg13g2_o21ai_1 _2592_ (.B1(_0311_),
    .Y(_0313_),
    .A1(_1545_),
    .A2(_0312_));
 sg13g2_a221oi_1 _2593_ (.B2(_0313_),
    .C1(_0308_),
    .B1(_1549_),
    .A1(\uart_inst.R0.clk_counter[12] ),
    .Y(_0314_),
    .A2(_1474_));
 sg13g2_nand2_1 _2594_ (.Y(_0315_),
    .A(_1448_),
    .B(_1449_));
 sg13g2_a21oi_2 _2595_ (.B1(_0315_),
    .Y(_0316_),
    .A2(_0314_),
    .A1(net948));
 sg13g2_inv_1 _2596_ (.Y(_0317_),
    .A(_0316_));
 sg13g2_nor4_2 _2597_ (.A(\bitty_inst.lsu_inst.rx_do ),
    .B(net910),
    .C(net596),
    .Y(_0318_),
    .D(_0317_));
 sg13g2_nor3_1 _2598_ (.A(\uart_inst.R0.bit_counter[2] ),
    .B(\uart_inst.R0.bit_counter[1] ),
    .C(\uart_inst.R0.bit_counter[0] ),
    .Y(_0319_));
 sg13g2_nor2_1 _2599_ (.A(\bitty_inst.lsu_inst.rx_data[0] ),
    .B(_0319_),
    .Y(_0320_));
 sg13g2_nor2b_1 _2600_ (.A(net827),
    .B_N(_0319_),
    .Y(_0321_));
 sg13g2_nor3_1 _2601_ (.A(_1601_),
    .B(_0320_),
    .C(_0321_),
    .Y(_0322_));
 sg13g2_nor2_2 _2602_ (.A(net820),
    .B(net652),
    .Y(_0323_));
 sg13g2_a22oi_1 _2603_ (.Y(_0324_),
    .B1(_0323_),
    .B2(\bitty_inst.lsu_inst.rx_data[0] ),
    .A2(_0322_),
    .A1(_0318_));
 sg13g2_inv_1 _2604_ (.Y(_0220_),
    .A(net911));
 sg13g2_nor2_1 _2605_ (.A(net928),
    .B(_0318_),
    .Y(_0325_));
 sg13g2_nand2_2 _2606_ (.Y(_0326_),
    .A(_1435_),
    .B(\uart_inst.R0.bit_counter[0] ));
 sg13g2_o21ai_1 _2607_ (.B1(\bitty_inst.lsu_inst.rx_data[1] ),
    .Y(_0327_),
    .A1(\uart_inst.R0.bit_counter[2] ),
    .A2(_0326_));
 sg13g2_nand2_1 _2608_ (.Y(_0328_),
    .A(_1434_),
    .B(net826));
 sg13g2_o21ai_1 _2609_ (.B1(_0327_),
    .Y(_0329_),
    .A1(_0326_),
    .A2(_0328_));
 sg13g2_a21oi_1 _2610_ (.A1(_1600_),
    .A2(_0329_),
    .Y(_0330_),
    .B1(_0323_));
 sg13g2_nor2_1 _2611_ (.A(_0325_),
    .B(_0330_),
    .Y(_0221_));
 sg13g2_nor2_1 _2612_ (.A(net924),
    .B(net652),
    .Y(_0331_));
 sg13g2_nand2_2 _2613_ (.Y(_0332_),
    .A(\uart_inst.R0.bit_counter[1] ),
    .B(_1436_));
 sg13g2_o21ai_1 _2614_ (.B1(\bitty_inst.lsu_inst.rx_data[2] ),
    .Y(_0333_),
    .A1(\uart_inst.R0.bit_counter[2] ),
    .A2(_0332_));
 sg13g2_o21ai_1 _2615_ (.B1(_0333_),
    .Y(_0334_),
    .A1(_0328_),
    .A2(_0332_));
 sg13g2_a21oi_1 _2616_ (.A1(_1600_),
    .A2(_0334_),
    .Y(_0335_),
    .B1(_0323_));
 sg13g2_nor2_1 _2617_ (.A(_0331_),
    .B(_0335_),
    .Y(_0222_));
 sg13g2_nor2_1 _2618_ (.A(\uart_inst.R0.bit_counter[2] ),
    .B(_1587_),
    .Y(_0336_));
 sg13g2_nor2_1 _2619_ (.A(\bitty_inst.lsu_inst.rx_data[3] ),
    .B(_0336_),
    .Y(_0337_));
 sg13g2_nor3_1 _2620_ (.A(\uart_inst.R0.bit_counter[2] ),
    .B(net826),
    .C(_1587_),
    .Y(_0338_));
 sg13g2_nor3_1 _2621_ (.A(_1601_),
    .B(_0337_),
    .C(_0338_),
    .Y(_0339_));
 sg13g2_a22oi_1 _2622_ (.Y(_0340_),
    .B1(_0339_),
    .B2(net652),
    .A2(_0323_),
    .A1(net953));
 sg13g2_inv_1 _2623_ (.Y(_0223_),
    .A(_0340_));
 sg13g2_nand2_1 _2624_ (.Y(_0341_),
    .A(net945),
    .B(_0323_));
 sg13g2_nor3_1 _2625_ (.A(net796),
    .B(\uart_inst.R0.bit_counter[1] ),
    .C(\uart_inst.R0.bit_counter[0] ),
    .Y(_0342_));
 sg13g2_mux2_1 _2626_ (.A0(\bitty_inst.lsu_inst.rx_data[4] ),
    .A1(net826),
    .S(_0342_),
    .X(_0343_));
 sg13g2_nand3_1 _2627_ (.B(net652),
    .C(_0343_),
    .A(_1600_),
    .Y(_0344_));
 sg13g2_nand2_1 _2628_ (.Y(_0224_),
    .A(_0341_),
    .B(_0344_));
 sg13g2_nor2_1 _2629_ (.A(net796),
    .B(_0326_),
    .Y(_0345_));
 sg13g2_nor2_1 _2630_ (.A(\bitty_inst.lsu_inst.rx_data[5] ),
    .B(_0345_),
    .Y(_0346_));
 sg13g2_nor3_1 _2631_ (.A(net796),
    .B(net826),
    .C(_0326_),
    .Y(_0347_));
 sg13g2_nor3_1 _2632_ (.A(_1601_),
    .B(_0346_),
    .C(_0347_),
    .Y(_0348_));
 sg13g2_a22oi_1 _2633_ (.Y(_0349_),
    .B1(_0348_),
    .B2(net652),
    .A2(_0323_),
    .A1(net959));
 sg13g2_inv_1 _2634_ (.Y(_0225_),
    .A(_0349_));
 sg13g2_nor2_1 _2635_ (.A(net796),
    .B(_0332_),
    .Y(_0350_));
 sg13g2_nor2_1 _2636_ (.A(\bitty_inst.lsu_inst.rx_data[6] ),
    .B(_0350_),
    .Y(_0351_));
 sg13g2_nor3_1 _2637_ (.A(net796),
    .B(net826),
    .C(_0332_),
    .Y(_0352_));
 sg13g2_nor3_1 _2638_ (.A(_1601_),
    .B(_0351_),
    .C(_0352_),
    .Y(_0353_));
 sg13g2_a22oi_1 _2639_ (.Y(_0354_),
    .B1(_0353_),
    .B2(net652),
    .A2(_0323_),
    .A1(net944));
 sg13g2_inv_1 _2640_ (.Y(_0226_),
    .A(_0354_));
 sg13g2_nor3_1 _2641_ (.A(net796),
    .B(net826),
    .C(_1587_),
    .Y(_0355_));
 sg13g2_o21ai_1 _2642_ (.B1(net886),
    .Y(_0356_),
    .A1(\bitty_inst.lsu_inst.rx_data[7] ),
    .A2(_1588_));
 sg13g2_o21ai_1 _2643_ (.B1(net652),
    .Y(_0357_),
    .A1(_0355_),
    .A2(_0356_));
 sg13g2_o21ai_1 _2644_ (.B1(net846),
    .Y(_0358_),
    .A1(net958),
    .A2(net652));
 sg13g2_nor2b_1 _2645_ (.A(_0358_),
    .B_N(_0357_),
    .Y(_0227_));
 sg13g2_nand2_2 _2646_ (.Y(_0359_),
    .A(net847),
    .B(_1583_));
 sg13g2_nor2_1 _2647_ (.A(\uart_inst.R0.PS[1] ),
    .B(net617),
    .Y(_0360_));
 sg13g2_nor2b_1 _2648_ (.A(_0360_),
    .B_N(_0314_),
    .Y(_0361_));
 sg13g2_a22oi_1 _2649_ (.Y(_0362_),
    .B1(_0361_),
    .B2(net602),
    .A2(_1585_),
    .A1(_1437_));
 sg13g2_nand2_1 _2650_ (.Y(_0363_),
    .A(\uart_inst.R0.clk_counter[0] ),
    .B(net655));
 sg13g2_o21ai_1 _2651_ (.B1(_0363_),
    .Y(_0228_),
    .A1(_0359_),
    .A2(net603));
 sg13g2_nor2_2 _2652_ (.A(_1585_),
    .B(_0361_),
    .Y(_0364_));
 sg13g2_and2_1 _2653_ (.A(_1583_),
    .B(_0364_),
    .X(_0365_));
 sg13g2_nand2b_2 _2654_ (.Y(_0366_),
    .B(net847),
    .A_N(_0365_));
 sg13g2_a21oi_1 _2655_ (.A1(net827),
    .A2(_1582_),
    .Y(_0367_),
    .B1(_1559_));
 sg13g2_a21oi_1 _2656_ (.A1(\uart_inst.R0.clk_counter[0] ),
    .A2(_1583_),
    .Y(_0368_),
    .B1(net898));
 sg13g2_nor3_1 _2657_ (.A(_0366_),
    .B(_0367_),
    .C(net899),
    .Y(_0229_));
 sg13g2_nor2_2 _2658_ (.A(_0359_),
    .B(_0364_),
    .Y(_0369_));
 sg13g2_nor2_1 _2659_ (.A(_0063_),
    .B(_1559_),
    .Y(_0370_));
 sg13g2_xor2_1 _2660_ (.B(_1559_),
    .A(_0063_),
    .X(_0371_));
 sg13g2_a22oi_1 _2661_ (.Y(_0372_),
    .B1(_0369_),
    .B2(_0371_),
    .A2(_1584_),
    .A1(net445));
 sg13g2_inv_1 _2662_ (.Y(_0230_),
    .A(net446));
 sg13g2_xor2_1 _2663_ (.B(_0370_),
    .A(_0062_),
    .X(_0373_));
 sg13g2_nor2_1 _2664_ (.A(_0359_),
    .B(_0373_),
    .Y(_0374_));
 sg13g2_a21oi_1 _2665_ (.A1(net875),
    .A2(_1584_),
    .Y(_0375_),
    .B1(_0374_));
 sg13g2_nor2_1 _2666_ (.A(_0365_),
    .B(net876),
    .Y(_0231_));
 sg13g2_nand4_1 _2667_ (.B(\uart_inst.R0.clk_counter[2] ),
    .C(\uart_inst.R0.clk_counter[1] ),
    .A(\uart_inst.R0.clk_counter[3] ),
    .Y(_0376_),
    .D(\uart_inst.R0.clk_counter[0] ));
 sg13g2_nor2_1 _2668_ (.A(_0061_),
    .B(_0376_),
    .Y(_0377_));
 sg13g2_xor2_1 _2669_ (.B(_0376_),
    .A(_0061_),
    .X(_0378_));
 sg13g2_a22oi_1 _2670_ (.Y(_0379_),
    .B1(_0369_),
    .B2(_0378_),
    .A2(net655),
    .A1(net430));
 sg13g2_inv_1 _2671_ (.Y(_0232_),
    .A(net431));
 sg13g2_xor2_1 _2672_ (.B(_0377_),
    .A(_0060_),
    .X(_0380_));
 sg13g2_nor2_1 _2673_ (.A(_0359_),
    .B(_0380_),
    .Y(_0381_));
 sg13g2_a21oi_1 _2674_ (.A1(net461),
    .A2(net655),
    .Y(_0382_),
    .B1(_0381_));
 sg13g2_nor2_1 _2675_ (.A(_0365_),
    .B(net462),
    .Y(_0233_));
 sg13g2_nand2_1 _2676_ (.Y(_0383_),
    .A(net461),
    .B(net430));
 sg13g2_nor2_2 _2677_ (.A(_0376_),
    .B(_0383_),
    .Y(_0384_));
 sg13g2_xnor2_1 _2678_ (.Y(_0385_),
    .A(_0059_),
    .B(_0384_));
 sg13g2_a22oi_1 _2679_ (.Y(_0386_),
    .B1(_0369_),
    .B2(_0385_),
    .A2(net655),
    .A1(net635));
 sg13g2_inv_1 _2680_ (.Y(_0234_),
    .A(net636));
 sg13g2_and3_1 _2681_ (.X(_0387_),
    .A(\uart_inst.R0.clk_counter[7] ),
    .B(\uart_inst.R0.clk_counter[6] ),
    .C(_0384_));
 sg13g2_a21oi_1 _2682_ (.A1(net635),
    .A2(_0384_),
    .Y(_0388_),
    .B1(net868));
 sg13g2_nor3_1 _2683_ (.A(_0366_),
    .B(_0387_),
    .C(_0388_),
    .Y(_0235_));
 sg13g2_nor2b_1 _2684_ (.A(_0058_),
    .B_N(_0387_),
    .Y(_0389_));
 sg13g2_xnor2_1 _2685_ (.Y(_0390_),
    .A(_0058_),
    .B(_0387_));
 sg13g2_a22oi_1 _2686_ (.Y(_0391_),
    .B1(_0369_),
    .B2(_0390_),
    .A2(net655),
    .A1(net581));
 sg13g2_inv_1 _2687_ (.Y(_0236_),
    .A(net582));
 sg13g2_xnor2_1 _2688_ (.Y(_0392_),
    .A(_0057_),
    .B(_0389_));
 sg13g2_a22oi_1 _2689_ (.Y(_0393_),
    .B1(_0369_),
    .B2(_0392_),
    .A2(net655),
    .A1(net618));
 sg13g2_inv_1 _2690_ (.Y(_0237_),
    .A(net619));
 sg13g2_and3_1 _2691_ (.X(_0394_),
    .A(\uart_inst.R0.clk_counter[9] ),
    .B(\uart_inst.R0.clk_counter[8] ),
    .C(_0387_));
 sg13g2_xnor2_1 _2692_ (.Y(_0395_),
    .A(_0056_),
    .B(_0394_));
 sg13g2_a22oi_1 _2693_ (.Y(_0396_),
    .B1(_0369_),
    .B2(_0395_),
    .A2(net655),
    .A1(net906));
 sg13g2_inv_1 _2694_ (.Y(_0238_),
    .A(net907));
 sg13g2_nand3_1 _2695_ (.B(net965),
    .C(_0394_),
    .A(\uart_inst.R0.clk_counter[11] ),
    .Y(_0397_));
 sg13g2_a21oi_1 _2696_ (.A1(net906),
    .A2(_0394_),
    .Y(_0398_),
    .B1(net955));
 sg13g2_nor2_1 _2697_ (.A(_0366_),
    .B(_0398_),
    .Y(_0399_));
 sg13g2_and2_1 _2698_ (.A(_0397_),
    .B(_0399_),
    .X(_0239_));
 sg13g2_xnor2_1 _2699_ (.Y(_0400_),
    .A(net492),
    .B(_0397_));
 sg13g2_nor3_1 _2700_ (.A(_0359_),
    .B(_0364_),
    .C(_0400_),
    .Y(_0240_));
 sg13g2_nand2_1 _2701_ (.Y(_0401_),
    .A(_1589_),
    .B(_0316_));
 sg13g2_a22oi_1 _2702_ (.Y(_0402_),
    .B1(_0401_),
    .B2(net845),
    .A2(_1600_),
    .A1(_1436_));
 sg13g2_a21oi_1 _2703_ (.A1(_1436_),
    .A2(_0401_),
    .Y(_0241_),
    .B1(_0402_));
 sg13g2_nand4_1 _2704_ (.B(net882),
    .C(_1600_),
    .A(_1435_),
    .Y(_0403_),
    .D(_0316_));
 sg13g2_o21ai_1 _2705_ (.B1(net883),
    .Y(_0242_),
    .A1(_1435_),
    .A2(_0402_));
 sg13g2_nand2b_1 _2706_ (.Y(_0404_),
    .B(_0316_),
    .A_N(_1587_));
 sg13g2_a221oi_1 _2707_ (.B2(net796),
    .C1(net820),
    .B1(_0404_),
    .A1(_1449_),
    .Y(_0243_),
    .A2(_0360_));
 sg13g2_nor2_1 _2708_ (.A(\bitty_inst.d_instr[2] ),
    .B(_1382_),
    .Y(_0405_));
 sg13g2_a22oi_1 _2709_ (.Y(_0406_),
    .B1(_1382_),
    .B2(\bitty_inst.d_instr[2] ),
    .A2(_1381_),
    .A1(\bitty_inst.d_instr[3] ));
 sg13g2_nor3_1 _2710_ (.A(\bitty_inst.d_out[15] ),
    .B(\bitty_inst.d_out[14] ),
    .C(_0405_),
    .Y(_0407_));
 sg13g2_nor4_1 _2711_ (.A(\bitty_inst.d_out[9] ),
    .B(\bitty_inst.d_out[8] ),
    .C(\bitty_inst.d_out[7] ),
    .D(\bitty_inst.d_out[6] ),
    .Y(_0408_));
 sg13g2_nor4_2 _2712_ (.A(\bitty_inst.d_out[13] ),
    .B(\bitty_inst.d_out[12] ),
    .C(\bitty_inst.d_out[11] ),
    .Y(_0409_),
    .D(\bitty_inst.d_out[10] ));
 sg13g2_and4_1 _2713_ (.A(_0406_),
    .B(_0407_),
    .C(_0408_),
    .D(_0409_),
    .X(_0410_));
 sg13g2_nand2b_1 _2714_ (.Y(_0411_),
    .B(\bitty_inst.d_instr[1] ),
    .A_N(\bitty_inst.d_instr[0] ));
 sg13g2_a21oi_2 _2715_ (.B1(_0411_),
    .Y(_0412_),
    .A2(\bitty_inst.d_instr[2] ),
    .A1(\bitty_inst.d_instr[3] ));
 sg13g2_o21ai_1 _2716_ (.B1(\bitty_inst.d_out[1] ),
    .Y(_0413_),
    .A1(_1353_),
    .A2(\bitty_inst.d_out[0] ));
 sg13g2_nor4_1 _2717_ (.A(\bitty_inst.d_out[5] ),
    .B(\bitty_inst.d_out[4] ),
    .C(\bitty_inst.d_out[3] ),
    .D(\bitty_inst.d_out[2] ),
    .Y(_0414_));
 sg13g2_mux2_1 _2718_ (.A0(_0054_),
    .A1(_1433_),
    .S(_0412_),
    .X(_0415_));
 sg13g2_nand4_1 _2719_ (.B(_0412_),
    .C(_0413_),
    .A(_0410_),
    .Y(_0416_),
    .D(_0414_));
 sg13g2_inv_2 _2720_ (.Y(_0417_),
    .A(net696));
 sg13g2_nand2_1 _2721_ (.Y(_0418_),
    .A(\bitty_inst.d_instr[4] ),
    .B(_0417_));
 sg13g2_a21oi_1 _2722_ (.A1(_0415_),
    .A2(net696),
    .Y(_0419_),
    .B1(_1431_));
 sg13g2_a221oi_1 _2723_ (.B2(_0419_),
    .C1(net819),
    .B1(_0418_),
    .A1(_1431_),
    .Y(_0244_),
    .A2(_1433_));
 sg13g2_nor2_1 _2724_ (.A(net813),
    .B(net908),
    .Y(_0420_));
 sg13g2_xor2_1 _2725_ (.B(net895),
    .A(net908),
    .X(_0421_));
 sg13g2_o21ai_1 _2726_ (.B1(net813),
    .Y(_0422_),
    .A1(_1351_),
    .A2(net696));
 sg13g2_a21oi_1 _2727_ (.A1(net696),
    .A2(_0421_),
    .Y(_0423_),
    .B1(_0422_));
 sg13g2_nor3_1 _2728_ (.A(net819),
    .B(_0420_),
    .C(_0423_),
    .Y(_0245_));
 sg13g2_nand3_1 _2729_ (.B(\addr[1] ),
    .C(\addr[0] ),
    .A(\addr[2] ),
    .Y(_0424_));
 sg13g2_a21o_1 _2730_ (.A2(\addr[0] ),
    .A1(\addr[1] ),
    .B1(\addr[2] ),
    .X(_0425_));
 sg13g2_nand2_1 _2731_ (.Y(_0426_),
    .A(_0424_),
    .B(_0425_));
 sg13g2_o21ai_1 _2732_ (.B1(net813),
    .Y(_0427_),
    .A1(_0417_),
    .A2(_0426_));
 sg13g2_a21oi_1 _2733_ (.A1(\bitty_inst.d_instr[6] ),
    .A2(_0417_),
    .Y(_0428_),
    .B1(_0427_));
 sg13g2_o21ai_1 _2734_ (.B1(net833),
    .Y(_0429_),
    .A1(net813),
    .A2(net914));
 sg13g2_nor2_1 _2735_ (.A(_0428_),
    .B(_0429_),
    .Y(_0246_));
 sg13g2_a21oi_1 _2736_ (.A1(\bitty_inst.d_instr[7] ),
    .A2(_0417_),
    .Y(_0430_),
    .B1(_1431_));
 sg13g2_nor2_2 _2737_ (.A(_1432_),
    .B(_0424_),
    .Y(_0431_));
 sg13g2_and2_1 _2738_ (.A(_1432_),
    .B(_0424_),
    .X(_0432_));
 sg13g2_or3_1 _2739_ (.A(_0417_),
    .B(_0431_),
    .C(_0432_),
    .X(_0433_));
 sg13g2_a221oi_1 _2740_ (.B2(_0433_),
    .C1(net819),
    .B1(_0430_),
    .A1(_1431_),
    .Y(_0247_),
    .A2(_1432_));
 sg13g2_nor3_1 _2741_ (.A(_1432_),
    .B(_0053_),
    .C(_0424_),
    .Y(_0434_));
 sg13g2_xnor2_1 _2742_ (.Y(_0435_),
    .A(_0053_),
    .B(_0431_));
 sg13g2_nand2_1 _2743_ (.Y(_0436_),
    .A(\bitty_inst.d_instr[8] ),
    .B(_0417_));
 sg13g2_a21oi_1 _2744_ (.A1(net696),
    .A2(_0435_),
    .Y(_0437_),
    .B1(_1431_));
 sg13g2_o21ai_1 _2745_ (.B1(net831),
    .Y(_0438_),
    .A1(net813),
    .A2(net926));
 sg13g2_a21oi_1 _2746_ (.A1(_0436_),
    .A2(_0437_),
    .Y(_0248_),
    .B1(_0438_));
 sg13g2_xor2_1 _2747_ (.B(_0434_),
    .A(\addr[5] ),
    .X(_0439_));
 sg13g2_o21ai_1 _2748_ (.B1(net813),
    .Y(_0440_),
    .A1(_1347_),
    .A2(net696));
 sg13g2_a21oi_1 _2749_ (.A1(_0416_),
    .A2(_0439_),
    .Y(_0441_),
    .B1(_0440_));
 sg13g2_o21ai_1 _2750_ (.B1(net831),
    .Y(_0442_),
    .A1(net814),
    .A2(net930));
 sg13g2_nor2_1 _2751_ (.A(_0441_),
    .B(_0442_),
    .Y(_0249_));
 sg13g2_a21oi_1 _2752_ (.A1(\bitty_inst.d_instr[10] ),
    .A2(_0417_),
    .Y(_0443_),
    .B1(_1431_));
 sg13g2_nand3_1 _2753_ (.B(\addr[4] ),
    .C(_0431_),
    .A(\addr[5] ),
    .Y(_0444_));
 sg13g2_nand4_1 _2754_ (.B(\addr[5] ),
    .C(\addr[4] ),
    .A(\addr[6] ),
    .Y(_0445_),
    .D(_0431_));
 sg13g2_nand2b_1 _2755_ (.Y(_0446_),
    .B(_0444_),
    .A_N(\addr[6] ));
 sg13g2_nand3_1 _2756_ (.B(_0445_),
    .C(_0446_),
    .A(net696),
    .Y(_0447_));
 sg13g2_o21ai_1 _2757_ (.B1(net831),
    .Y(_0448_),
    .A1(net813),
    .A2(net937));
 sg13g2_a21oi_1 _2758_ (.A1(_0443_),
    .A2(_0447_),
    .Y(_0250_),
    .B1(_0448_));
 sg13g2_xnor2_1 _2759_ (.Y(_0449_),
    .A(\addr[7] ),
    .B(_0445_));
 sg13g2_o21ai_1 _2760_ (.B1(net814),
    .Y(_0450_),
    .A1(_1345_),
    .A2(net696));
 sg13g2_a21oi_1 _2761_ (.A1(_0416_),
    .A2(_0449_),
    .Y(_0451_),
    .B1(_0450_));
 sg13g2_o21ai_1 _2762_ (.B1(net831),
    .Y(_0452_),
    .A1(net932),
    .A2(net813));
 sg13g2_nor2_1 _2763_ (.A(_0451_),
    .B(_0452_),
    .Y(_0251_));
 sg13g2_a21oi_2 _2764_ (.B1(_1442_),
    .Y(_0453_),
    .A2(_1517_),
    .A1(net801));
 sg13g2_nand2_1 _2765_ (.Y(_0454_),
    .A(\bitty_inst.cpu_inst.d_inst[14] ),
    .B(_0453_));
 sg13g2_nand4_1 _2766_ (.B(\bitty_inst.cpu_inst.d_inst[14] ),
    .C(\bitty_inst.cpu_inst.d_inst[13] ),
    .A(\bitty_inst.cpu_inst.d_inst[15] ),
    .Y(_0455_),
    .D(_0453_));
 sg13g2_o21ai_1 _2767_ (.B1(net836),
    .Y(_0456_),
    .A1(\bitty_inst.d_out[0] ),
    .A2(net771));
 sg13g2_a21oi_1 _2768_ (.A1(_1430_),
    .A2(net770),
    .Y(_0252_),
    .B1(_0456_));
 sg13g2_o21ai_1 _2769_ (.B1(net835),
    .Y(_0457_),
    .A1(\bitty_inst.d_out[1] ),
    .A2(net770));
 sg13g2_a21oi_1 _2770_ (.A1(_1429_),
    .A2(net770),
    .Y(_0253_),
    .B1(_0457_));
 sg13g2_o21ai_1 _2771_ (.B1(net834),
    .Y(_0458_),
    .A1(\bitty_inst.d_out[2] ),
    .A2(net770));
 sg13g2_a21oi_1 _2772_ (.A1(_1428_),
    .A2(net770),
    .Y(_0254_),
    .B1(_0458_));
 sg13g2_o21ai_1 _2773_ (.B1(net836),
    .Y(_0459_),
    .A1(\bitty_inst.d_out[3] ),
    .A2(net771));
 sg13g2_a21oi_1 _2774_ (.A1(_1427_),
    .A2(net770),
    .Y(_0255_),
    .B1(_0459_));
 sg13g2_o21ai_1 _2775_ (.B1(net841),
    .Y(_0460_),
    .A1(\bitty_inst.d_out[4] ),
    .A2(net771));
 sg13g2_a21oi_1 _2776_ (.A1(_1426_),
    .A2(net771),
    .Y(_0256_),
    .B1(_0460_));
 sg13g2_o21ai_1 _2777_ (.B1(net840),
    .Y(_0461_),
    .A1(\bitty_inst.d_out[5] ),
    .A2(net774));
 sg13g2_a21oi_1 _2778_ (.A1(_1425_),
    .A2(net771),
    .Y(_0257_),
    .B1(_0461_));
 sg13g2_o21ai_1 _2779_ (.B1(net838),
    .Y(_0462_),
    .A1(\bitty_inst.d_out[6] ),
    .A2(net770));
 sg13g2_a21oi_1 _2780_ (.A1(_1424_),
    .A2(net770),
    .Y(_0258_),
    .B1(_0462_));
 sg13g2_o21ai_1 _2781_ (.B1(net841),
    .Y(_0463_),
    .A1(\bitty_inst.d_out[7] ),
    .A2(net771));
 sg13g2_a21oi_1 _2782_ (.A1(_1423_),
    .A2(net771),
    .Y(_0259_),
    .B1(_0463_));
 sg13g2_o21ai_1 _2783_ (.B1(net857),
    .Y(_0464_),
    .A1(\bitty_inst.d_out[8] ),
    .A2(net772));
 sg13g2_a21oi_1 _2784_ (.A1(_1422_),
    .A2(net772),
    .Y(_0260_),
    .B1(_0464_));
 sg13g2_o21ai_1 _2785_ (.B1(net850),
    .Y(_0465_),
    .A1(\bitty_inst.d_out[9] ),
    .A2(net773));
 sg13g2_a21oi_1 _2786_ (.A1(_1421_),
    .A2(net773),
    .Y(_0261_),
    .B1(_0465_));
 sg13g2_o21ai_1 _2787_ (.B1(net855),
    .Y(_0466_),
    .A1(\bitty_inst.d_out[10] ),
    .A2(net773));
 sg13g2_a21oi_1 _2788_ (.A1(_1420_),
    .A2(net774),
    .Y(_0262_),
    .B1(_0466_));
 sg13g2_o21ai_1 _2789_ (.B1(net857),
    .Y(_0467_),
    .A1(\bitty_inst.d_out[11] ),
    .A2(net772));
 sg13g2_a21oi_1 _2790_ (.A1(_1419_),
    .A2(net772),
    .Y(_0263_),
    .B1(_0467_));
 sg13g2_o21ai_1 _2791_ (.B1(net854),
    .Y(_0468_),
    .A1(\bitty_inst.d_out[12] ),
    .A2(net772));
 sg13g2_a21oi_1 _2792_ (.A1(_1418_),
    .A2(net772),
    .Y(_0264_),
    .B1(_0468_));
 sg13g2_o21ai_1 _2793_ (.B1(net860),
    .Y(_0469_),
    .A1(\bitty_inst.d_out[13] ),
    .A2(net772));
 sg13g2_a21oi_1 _2794_ (.A1(_1417_),
    .A2(net772),
    .Y(_0265_),
    .B1(_0469_));
 sg13g2_o21ai_1 _2795_ (.B1(net851),
    .Y(_0470_),
    .A1(\bitty_inst.d_out[14] ),
    .A2(net773));
 sg13g2_a21oi_1 _2796_ (.A1(_1416_),
    .A2(net773),
    .Y(_0266_),
    .B1(_0470_));
 sg13g2_o21ai_1 _2797_ (.B1(net849),
    .Y(_0471_),
    .A1(\bitty_inst.d_out[15] ),
    .A2(net773));
 sg13g2_a21oi_1 _2798_ (.A1(_1415_),
    .A2(net773),
    .Y(_0267_),
    .B1(_0471_));
 sg13g2_nand4_1 _2799_ (.B(\bitty_inst.cpu_inst.d_inst[14] ),
    .C(_1343_),
    .A(\bitty_inst.cpu_inst.d_inst[15] ),
    .Y(_0472_),
    .D(_0453_));
 sg13g2_o21ai_1 _2800_ (.B1(net836),
    .Y(_0473_),
    .A1(\bitty_inst.d_out[0] ),
    .A2(net766));
 sg13g2_a21oi_1 _2801_ (.A1(_1414_),
    .A2(net766),
    .Y(_0268_),
    .B1(_0473_));
 sg13g2_o21ai_1 _2802_ (.B1(net835),
    .Y(_0474_),
    .A1(\bitty_inst.d_out[1] ),
    .A2(net765));
 sg13g2_a21oi_1 _2803_ (.A1(_1413_),
    .A2(net765),
    .Y(_0269_),
    .B1(_0474_));
 sg13g2_o21ai_1 _2804_ (.B1(net834),
    .Y(_0475_),
    .A1(\bitty_inst.d_out[2] ),
    .A2(net765));
 sg13g2_a21oi_1 _2805_ (.A1(_1412_),
    .A2(net765),
    .Y(_0270_),
    .B1(_0475_));
 sg13g2_o21ai_1 _2806_ (.B1(net843),
    .Y(_0476_),
    .A1(\bitty_inst.d_out[3] ),
    .A2(net765));
 sg13g2_a21oi_1 _2807_ (.A1(_1411_),
    .A2(net765),
    .Y(_0271_),
    .B1(_0476_));
 sg13g2_o21ai_1 _2808_ (.B1(net841),
    .Y(_0477_),
    .A1(\bitty_inst.d_out[4] ),
    .A2(net767));
 sg13g2_a21oi_1 _2809_ (.A1(_1410_),
    .A2(net767),
    .Y(_0272_),
    .B1(_0477_));
 sg13g2_o21ai_1 _2810_ (.B1(net839),
    .Y(_0478_),
    .A1(\bitty_inst.d_out[5] ),
    .A2(net766));
 sg13g2_a21oi_1 _2811_ (.A1(_1409_),
    .A2(net766),
    .Y(_0273_),
    .B1(_0478_));
 sg13g2_o21ai_1 _2812_ (.B1(net838),
    .Y(_0479_),
    .A1(\bitty_inst.d_out[6] ),
    .A2(net765));
 sg13g2_a21oi_1 _2813_ (.A1(_1408_),
    .A2(net765),
    .Y(_0274_),
    .B1(_0479_));
 sg13g2_o21ai_1 _2814_ (.B1(net841),
    .Y(_0480_),
    .A1(\bitty_inst.d_out[7] ),
    .A2(net767));
 sg13g2_a21oi_1 _2815_ (.A1(_1407_),
    .A2(net766),
    .Y(_0275_),
    .B1(_0480_));
 sg13g2_o21ai_1 _2816_ (.B1(net857),
    .Y(_0481_),
    .A1(\bitty_inst.d_out[8] ),
    .A2(net768));
 sg13g2_a21oi_1 _2817_ (.A1(_1406_),
    .A2(net768),
    .Y(_0276_),
    .B1(_0481_));
 sg13g2_o21ai_1 _2818_ (.B1(net851),
    .Y(_0482_),
    .A1(\bitty_inst.d_out[9] ),
    .A2(net769));
 sg13g2_a21oi_1 _2819_ (.A1(_1405_),
    .A2(net769),
    .Y(_0277_),
    .B1(_0482_));
 sg13g2_o21ai_1 _2820_ (.B1(net855),
    .Y(_0483_),
    .A1(\bitty_inst.d_out[10] ),
    .A2(net768));
 sg13g2_a21oi_1 _2821_ (.A1(_1404_),
    .A2(net768),
    .Y(_0278_),
    .B1(_0483_));
 sg13g2_o21ai_1 _2822_ (.B1(net861),
    .Y(_0484_),
    .A1(\bitty_inst.d_out[11] ),
    .A2(_0472_));
 sg13g2_a21oi_1 _2823_ (.A1(_1403_),
    .A2(net769),
    .Y(_0279_),
    .B1(_0484_));
 sg13g2_o21ai_1 _2824_ (.B1(net855),
    .Y(_0485_),
    .A1(\bitty_inst.d_out[12] ),
    .A2(net768));
 sg13g2_a21oi_1 _2825_ (.A1(_1402_),
    .A2(net768),
    .Y(_0280_),
    .B1(_0485_));
 sg13g2_o21ai_1 _2826_ (.B1(net859),
    .Y(_0486_),
    .A1(\bitty_inst.d_out[13] ),
    .A2(net768));
 sg13g2_a21oi_1 _2827_ (.A1(_1401_),
    .A2(net768),
    .Y(_0281_),
    .B1(_0486_));
 sg13g2_o21ai_1 _2828_ (.B1(net851),
    .Y(_0487_),
    .A1(\bitty_inst.d_out[14] ),
    .A2(net769));
 sg13g2_a21oi_1 _2829_ (.A1(_1400_),
    .A2(net769),
    .Y(_0282_),
    .B1(_0487_));
 sg13g2_o21ai_1 _2830_ (.B1(net850),
    .Y(_0488_),
    .A1(\bitty_inst.d_out[15] ),
    .A2(net769));
 sg13g2_a21oi_1 _2831_ (.A1(_1399_),
    .A2(net769),
    .Y(_0283_),
    .B1(_0488_));
 sg13g2_nor2_1 _2832_ (.A(\bitty_inst.cpu_inst.d_inst[14] ),
    .B(_1343_),
    .Y(_0489_));
 sg13g2_nand3_1 _2833_ (.B(_0453_),
    .C(_0489_),
    .A(\bitty_inst.cpu_inst.d_inst[15] ),
    .Y(_0490_));
 sg13g2_o21ai_1 _2834_ (.B1(net836),
    .Y(_0491_),
    .A1(\bitty_inst.d_out[0] ),
    .A2(net760));
 sg13g2_a21oi_1 _2835_ (.A1(_1398_),
    .A2(net760),
    .Y(_0284_),
    .B1(_0491_));
 sg13g2_o21ai_1 _2836_ (.B1(net837),
    .Y(_0492_),
    .A1(\bitty_inst.d_out[1] ),
    .A2(net760));
 sg13g2_a21oi_1 _2837_ (.A1(_1397_),
    .A2(net760),
    .Y(_0285_),
    .B1(_0492_));
 sg13g2_o21ai_1 _2838_ (.B1(net836),
    .Y(_0493_),
    .A1(\bitty_inst.d_out[2] ),
    .A2(net760));
 sg13g2_a21oi_1 _2839_ (.A1(_1396_),
    .A2(net760),
    .Y(_0286_),
    .B1(_0493_));
 sg13g2_o21ai_1 _2840_ (.B1(net843),
    .Y(_0494_),
    .A1(\bitty_inst.d_out[3] ),
    .A2(net761));
 sg13g2_a21oi_1 _2841_ (.A1(_1395_),
    .A2(net761),
    .Y(_0287_),
    .B1(_0494_));
 sg13g2_o21ai_1 _2842_ (.B1(net840),
    .Y(_0495_),
    .A1(\bitty_inst.d_out[4] ),
    .A2(net761));
 sg13g2_a21oi_1 _2843_ (.A1(_1394_),
    .A2(net761),
    .Y(_0288_),
    .B1(_0495_));
 sg13g2_o21ai_1 _2844_ (.B1(net840),
    .Y(_0496_),
    .A1(\bitty_inst.d_out[5] ),
    .A2(net761));
 sg13g2_a21oi_1 _2845_ (.A1(_1393_),
    .A2(net761),
    .Y(_0289_),
    .B1(_0496_));
 sg13g2_o21ai_1 _2846_ (.B1(net838),
    .Y(_0497_),
    .A1(\bitty_inst.d_out[6] ),
    .A2(net760));
 sg13g2_a21oi_1 _2847_ (.A1(_1392_),
    .A2(net760),
    .Y(_0290_),
    .B1(_0497_));
 sg13g2_o21ai_1 _2848_ (.B1(net842),
    .Y(_0498_),
    .A1(\bitty_inst.d_out[7] ),
    .A2(net762));
 sg13g2_a21oi_1 _2849_ (.A1(_1391_),
    .A2(net762),
    .Y(_0291_),
    .B1(_0498_));
 sg13g2_o21ai_1 _2850_ (.B1(net857),
    .Y(_0499_),
    .A1(\bitty_inst.d_out[8] ),
    .A2(net763));
 sg13g2_a21oi_1 _2851_ (.A1(_1390_),
    .A2(net763),
    .Y(_0292_),
    .B1(_0499_));
 sg13g2_o21ai_1 _2852_ (.B1(net851),
    .Y(_0500_),
    .A1(\bitty_inst.d_out[9] ),
    .A2(net764));
 sg13g2_a21oi_1 _2853_ (.A1(_1389_),
    .A2(net764),
    .Y(_0293_),
    .B1(_0500_));
 sg13g2_o21ai_1 _2854_ (.B1(net855),
    .Y(_0501_),
    .A1(\bitty_inst.d_out[10] ),
    .A2(net763));
 sg13g2_a21oi_1 _2855_ (.A1(_1388_),
    .A2(net763),
    .Y(_0294_),
    .B1(_0501_));
 sg13g2_o21ai_1 _2856_ (.B1(net859),
    .Y(_0502_),
    .A1(\bitty_inst.d_out[11] ),
    .A2(net763));
 sg13g2_a21oi_1 _2857_ (.A1(_1387_),
    .A2(net764),
    .Y(_0295_),
    .B1(_0502_));
 sg13g2_o21ai_1 _2858_ (.B1(net855),
    .Y(_0503_),
    .A1(\bitty_inst.d_out[12] ),
    .A2(net763));
 sg13g2_a21oi_1 _2859_ (.A1(_1386_),
    .A2(net763),
    .Y(_0296_),
    .B1(_0503_));
 sg13g2_o21ai_1 _2860_ (.B1(net860),
    .Y(_0504_),
    .A1(\bitty_inst.d_out[13] ),
    .A2(_0490_));
 sg13g2_a21oi_1 _2861_ (.A1(_1385_),
    .A2(net763),
    .Y(_0297_),
    .B1(_0504_));
 sg13g2_o21ai_1 _2862_ (.B1(net851),
    .Y(_0505_),
    .A1(\bitty_inst.d_out[14] ),
    .A2(net764));
 sg13g2_a21oi_1 _2863_ (.A1(_1384_),
    .A2(net764),
    .Y(_0298_),
    .B1(_0505_));
 sg13g2_o21ai_1 _2864_ (.B1(net850),
    .Y(_0506_),
    .A1(\bitty_inst.d_out[15] ),
    .A2(net764));
 sg13g2_a21oi_1 _2865_ (.A1(_1383_),
    .A2(net764),
    .Y(_0299_),
    .B1(_0506_));
 sg13g2_and4_1 _2866_ (.A(\bitty_inst.cpu_inst.d_inst[15] ),
    .B(_1342_),
    .C(_1343_),
    .D(_0453_),
    .X(_0507_));
 sg13g2_o21ai_1 _2867_ (.B1(net841),
    .Y(_0508_),
    .A1(net465),
    .A2(net759));
 sg13g2_a21oi_1 _2868_ (.A1(_1382_),
    .A2(net756),
    .Y(_0300_),
    .B1(_0508_));
 sg13g2_o21ai_1 _2869_ (.B1(net835),
    .Y(_0509_),
    .A1(net646),
    .A2(net755));
 sg13g2_a21oi_1 _2870_ (.A1(_1381_),
    .A2(net755),
    .Y(_0301_),
    .B1(_0509_));
 sg13g2_o21ai_1 _2871_ (.B1(net834),
    .Y(_0510_),
    .A1(net521),
    .A2(net755));
 sg13g2_a21oi_1 _2872_ (.A1(_1380_),
    .A2(net755),
    .Y(_0302_),
    .B1(_0510_));
 sg13g2_o21ai_1 _2873_ (.B1(net835),
    .Y(_0511_),
    .A1(net499),
    .A2(net755));
 sg13g2_a21oi_1 _2874_ (.A1(_1379_),
    .A2(net755),
    .Y(_0303_),
    .B1(_0511_));
 sg13g2_o21ai_1 _2875_ (.B1(net840),
    .Y(_0512_),
    .A1(net623),
    .A2(net756));
 sg13g2_a21oi_1 _2876_ (.A1(_1378_),
    .A2(net756),
    .Y(_0076_),
    .B1(_0512_));
 sg13g2_o21ai_1 _2877_ (.B1(net839),
    .Y(_0513_),
    .A1(net589),
    .A2(net755));
 sg13g2_a21oi_1 _2878_ (.A1(_1377_),
    .A2(net755),
    .Y(_0077_),
    .B1(_0513_));
 sg13g2_o21ai_1 _2879_ (.B1(net838),
    .Y(_0514_),
    .A1(net553),
    .A2(net756));
 sg13g2_a21oi_1 _2880_ (.A1(_1376_),
    .A2(net756),
    .Y(_0078_),
    .B1(_0514_));
 sg13g2_o21ai_1 _2881_ (.B1(net842),
    .Y(_0515_),
    .A1(net585),
    .A2(net756));
 sg13g2_a21oi_1 _2882_ (.A1(_1375_),
    .A2(net756),
    .Y(_0079_),
    .B1(_0515_));
 sg13g2_o21ai_1 _2883_ (.B1(net858),
    .Y(_0516_),
    .A1(net583),
    .A2(net758));
 sg13g2_a21oi_1 _2884_ (.A1(_1374_),
    .A2(net759),
    .Y(_0080_),
    .B1(_0516_));
 sg13g2_o21ai_1 _2885_ (.B1(net850),
    .Y(_0517_),
    .A1(net559),
    .A2(net758));
 sg13g2_a21oi_1 _2886_ (.A1(_1373_),
    .A2(net758),
    .Y(_0081_),
    .B1(_0517_));
 sg13g2_o21ai_1 _2887_ (.B1(net854),
    .Y(_0518_),
    .A1(net459),
    .A2(net757));
 sg13g2_a21oi_1 _2888_ (.A1(_1372_),
    .A2(net757),
    .Y(_0082_),
    .B1(_0518_));
 sg13g2_o21ai_1 _2889_ (.B1(net859),
    .Y(_0519_),
    .A1(net538),
    .A2(net757));
 sg13g2_a21oi_1 _2890_ (.A1(_1371_),
    .A2(net757),
    .Y(_0083_),
    .B1(_0519_));
 sg13g2_o21ai_1 _2891_ (.B1(net860),
    .Y(_0520_),
    .A1(net452),
    .A2(net757));
 sg13g2_a21oi_1 _2892_ (.A1(_1370_),
    .A2(net757),
    .Y(_0084_),
    .B1(_0520_));
 sg13g2_o21ai_1 _2893_ (.B1(net860),
    .Y(_0521_),
    .A1(net540),
    .A2(net757));
 sg13g2_a21oi_1 _2894_ (.A1(_1369_),
    .A2(net757),
    .Y(_0085_),
    .B1(_0521_));
 sg13g2_o21ai_1 _2895_ (.B1(net851),
    .Y(_0522_),
    .A1(net463),
    .A2(net758));
 sg13g2_a21oi_1 _2896_ (.A1(_1368_),
    .A2(net758),
    .Y(_0086_),
    .B1(_0522_));
 sg13g2_o21ai_1 _2897_ (.B1(net849),
    .Y(_0523_),
    .A1(net490),
    .A2(net758));
 sg13g2_a21oi_1 _2898_ (.A1(_1366_),
    .A2(net758),
    .Y(_0087_),
    .B1(_0523_));
 sg13g2_nor3_2 _2899_ (.A(\bitty_inst.cpu_inst.d_inst[15] ),
    .B(_1343_),
    .C(_0454_),
    .Y(_0524_));
 sg13g2_o21ai_1 _2900_ (.B1(net839),
    .Y(_0525_),
    .A1(net600),
    .A2(net725));
 sg13g2_a21oi_1 _2901_ (.A1(_1382_),
    .A2(net725),
    .Y(_0088_),
    .B1(_0525_));
 sg13g2_o21ai_1 _2902_ (.B1(net835),
    .Y(_0526_),
    .A1(net606),
    .A2(net724));
 sg13g2_a21oi_1 _2903_ (.A1(_1381_),
    .A2(net724),
    .Y(_0089_),
    .B1(_0526_));
 sg13g2_o21ai_1 _2904_ (.B1(net834),
    .Y(_0527_),
    .A1(net536),
    .A2(net724));
 sg13g2_a21oi_1 _2905_ (.A1(_1380_),
    .A2(net724),
    .Y(_0090_),
    .B1(_0527_));
 sg13g2_o21ai_1 _2906_ (.B1(net835),
    .Y(_0528_),
    .A1(net574),
    .A2(net724));
 sg13g2_a21oi_1 _2907_ (.A1(_1379_),
    .A2(net724),
    .Y(_0091_),
    .B1(_0528_));
 sg13g2_o21ai_1 _2908_ (.B1(net840),
    .Y(_0529_),
    .A1(net565),
    .A2(net726));
 sg13g2_a21oi_1 _2909_ (.A1(_1378_),
    .A2(net726),
    .Y(_0092_),
    .B1(_0529_));
 sg13g2_o21ai_1 _2910_ (.B1(net839),
    .Y(_0530_),
    .A1(net628),
    .A2(net725));
 sg13g2_a21oi_1 _2911_ (.A1(_1377_),
    .A2(net724),
    .Y(_0093_),
    .B1(_0530_));
 sg13g2_o21ai_1 _2912_ (.B1(net838),
    .Y(_0531_),
    .A1(net501),
    .A2(net724));
 sg13g2_a21oi_1 _2913_ (.A1(_1376_),
    .A2(net725),
    .Y(_0094_),
    .B1(_0531_));
 sg13g2_o21ai_1 _2914_ (.B1(net842),
    .Y(_0532_),
    .A1(net610),
    .A2(net726));
 sg13g2_a21oi_1 _2915_ (.A1(_1375_),
    .A2(net726),
    .Y(_0095_),
    .B1(_0532_));
 sg13g2_o21ai_1 _2916_ (.B1(net857),
    .Y(_0533_),
    .A1(net511),
    .A2(net728));
 sg13g2_a21oi_1 _2917_ (.A1(_1374_),
    .A2(_0524_),
    .Y(_0096_),
    .B1(_0533_));
 sg13g2_o21ai_1 _2918_ (.B1(net849),
    .Y(_0534_),
    .A1(net627),
    .A2(net728));
 sg13g2_a21oi_1 _2919_ (.A1(_1373_),
    .A2(net728),
    .Y(_0097_),
    .B1(_0534_));
 sg13g2_o21ai_1 _2920_ (.B1(net854),
    .Y(_0535_),
    .A1(net555),
    .A2(net727));
 sg13g2_a21oi_1 _2921_ (.A1(_1372_),
    .A2(net727),
    .Y(_0098_),
    .B1(_0535_));
 sg13g2_o21ai_1 _2922_ (.B1(net859),
    .Y(_0536_),
    .A1(net570),
    .A2(net727));
 sg13g2_a21oi_1 _2923_ (.A1(_1371_),
    .A2(net727),
    .Y(_0099_),
    .B1(_0536_));
 sg13g2_o21ai_1 _2924_ (.B1(net858),
    .Y(_0537_),
    .A1(net473),
    .A2(net727));
 sg13g2_a21oi_1 _2925_ (.A1(_1370_),
    .A2(net727),
    .Y(_0100_),
    .B1(_0537_));
 sg13g2_o21ai_1 _2926_ (.B1(net859),
    .Y(_0538_),
    .A1(net870),
    .A2(net727));
 sg13g2_a21oi_1 _2927_ (.A1(_1369_),
    .A2(net727),
    .Y(_0101_),
    .B1(_0538_));
 sg13g2_o21ai_1 _2928_ (.B1(net852),
    .Y(_0539_),
    .A1(net527),
    .A2(net728));
 sg13g2_a21oi_1 _2929_ (.A1(_1368_),
    .A2(net728),
    .Y(_0102_),
    .B1(_0539_));
 sg13g2_o21ai_1 _2930_ (.B1(net849),
    .Y(_0540_),
    .A1(net517),
    .A2(net728));
 sg13g2_a21oi_1 _2931_ (.A1(_1366_),
    .A2(net728),
    .Y(_0103_),
    .B1(_0540_));
 sg13g2_nor3_1 _2932_ (.A(\bitty_inst.cpu_inst.d_inst[15] ),
    .B(\bitty_inst.cpu_inst.d_inst[13] ),
    .C(_0454_),
    .Y(_0541_));
 sg13g2_o21ai_1 _2933_ (.B1(net839),
    .Y(_0542_),
    .A1(net519),
    .A2(net719));
 sg13g2_a21oi_1 _2934_ (.A1(_1382_),
    .A2(net719),
    .Y(_0104_),
    .B1(_0542_));
 sg13g2_o21ai_1 _2935_ (.B1(net835),
    .Y(_0543_),
    .A1(net531),
    .A2(net719));
 sg13g2_a21oi_1 _2936_ (.A1(_1381_),
    .A2(net719),
    .Y(_0105_),
    .B1(_0543_));
 sg13g2_o21ai_1 _2937_ (.B1(net834),
    .Y(_0544_),
    .A1(net481),
    .A2(net719));
 sg13g2_a21oi_1 _2938_ (.A1(_1380_),
    .A2(net719),
    .Y(_0106_),
    .B1(_0544_));
 sg13g2_o21ai_1 _2939_ (.B1(net843),
    .Y(_0545_),
    .A1(net486),
    .A2(net720));
 sg13g2_a21oi_1 _2940_ (.A1(_1379_),
    .A2(net720),
    .Y(_0107_),
    .B1(_0545_));
 sg13g2_o21ai_1 _2941_ (.B1(net842),
    .Y(_0546_),
    .A1(net475),
    .A2(net720));
 sg13g2_a21oi_1 _2942_ (.A1(_1378_),
    .A2(net720),
    .Y(_0108_),
    .B1(_0546_));
 sg13g2_o21ai_1 _2943_ (.B1(net840),
    .Y(_0547_),
    .A1(net560),
    .A2(net720));
 sg13g2_a21oi_1 _2944_ (.A1(_1377_),
    .A2(net720),
    .Y(_0109_),
    .B1(_0547_));
 sg13g2_o21ai_1 _2945_ (.B1(net838),
    .Y(_0548_),
    .A1(net612),
    .A2(net719));
 sg13g2_a21oi_1 _2946_ (.A1(_1376_),
    .A2(net719),
    .Y(_0110_),
    .B1(_0548_));
 sg13g2_o21ai_1 _2947_ (.B1(net841),
    .Y(_0549_),
    .A1(net631),
    .A2(net720));
 sg13g2_a21oi_1 _2948_ (.A1(_1375_),
    .A2(net720),
    .Y(_0111_),
    .B1(_0549_));
 sg13g2_o21ai_1 _2949_ (.B1(net858),
    .Y(_0550_),
    .A1(net625),
    .A2(net721));
 sg13g2_a21oi_1 _2950_ (.A1(_1374_),
    .A2(net721),
    .Y(_0112_),
    .B1(_0550_));
 sg13g2_o21ai_1 _2951_ (.B1(net852),
    .Y(_0551_),
    .A1(net608),
    .A2(net722));
 sg13g2_a21oi_1 _2952_ (.A1(_1373_),
    .A2(net722),
    .Y(_0113_),
    .B1(_0551_));
 sg13g2_o21ai_1 _2953_ (.B1(net854),
    .Y(_0552_),
    .A1(net525),
    .A2(net721));
 sg13g2_a21oi_1 _2954_ (.A1(_1372_),
    .A2(net721),
    .Y(_0114_),
    .B1(_0552_));
 sg13g2_o21ai_1 _2955_ (.B1(net857),
    .Y(_0553_),
    .A1(net567),
    .A2(net721));
 sg13g2_a21oi_1 _2956_ (.A1(_1371_),
    .A2(net721),
    .Y(_0115_),
    .B1(_0553_));
 sg13g2_o21ai_1 _2957_ (.B1(net858),
    .Y(_0554_),
    .A1(net469),
    .A2(net722));
 sg13g2_a21oi_1 _2958_ (.A1(_1370_),
    .A2(net723),
    .Y(_0116_),
    .B1(_0554_));
 sg13g2_o21ai_1 _2959_ (.B1(net859),
    .Y(_0555_),
    .A1(net507),
    .A2(net721));
 sg13g2_a21oi_1 _2960_ (.A1(_1369_),
    .A2(net721),
    .Y(_0117_),
    .B1(_0555_));
 sg13g2_o21ai_1 _2961_ (.B1(net851),
    .Y(_0556_),
    .A1(net529),
    .A2(net722));
 sg13g2_a21oi_1 _2962_ (.A1(_1368_),
    .A2(net722),
    .Y(_0118_),
    .B1(_0556_));
 sg13g2_o21ai_1 _2963_ (.B1(net849),
    .Y(_0557_),
    .A1(net547),
    .A2(net722));
 sg13g2_a21oi_1 _2964_ (.A1(_1366_),
    .A2(net722),
    .Y(_0119_),
    .B1(_0557_));
 sg13g2_and3_2 _2965_ (.X(_0558_),
    .A(_1341_),
    .B(_0453_),
    .C(_0489_));
 sg13g2_o21ai_1 _2966_ (.B1(net839),
    .Y(_0559_),
    .A1(net544),
    .A2(net750));
 sg13g2_a21oi_1 _2967_ (.A1(_1382_),
    .A2(net750),
    .Y(_0120_),
    .B1(_0559_));
 sg13g2_o21ai_1 _2968_ (.B1(net836),
    .Y(_0560_),
    .A1(net633),
    .A2(net750));
 sg13g2_a21oi_1 _2969_ (.A1(_1381_),
    .A2(net750),
    .Y(_0121_),
    .B1(_0560_));
 sg13g2_o21ai_1 _2970_ (.B1(net834),
    .Y(_0561_),
    .A1(net513),
    .A2(net750));
 sg13g2_a21oi_1 _2971_ (.A1(_1380_),
    .A2(net750),
    .Y(_0122_),
    .B1(_0561_));
 sg13g2_o21ai_1 _2972_ (.B1(net843),
    .Y(_0562_),
    .A1(net495),
    .A2(net750));
 sg13g2_a21oi_1 _2973_ (.A1(_1379_),
    .A2(net750),
    .Y(_0123_),
    .B1(_0562_));
 sg13g2_o21ai_1 _2974_ (.B1(net842),
    .Y(_0563_),
    .A1(net577),
    .A2(net752));
 sg13g2_a21oi_1 _2975_ (.A1(_1378_),
    .A2(net752),
    .Y(_0124_),
    .B1(_0563_));
 sg13g2_o21ai_1 _2976_ (.B1(net840),
    .Y(_0564_),
    .A1(net488),
    .A2(net751));
 sg13g2_a21oi_1 _2977_ (.A1(_1377_),
    .A2(net751),
    .Y(_0125_),
    .B1(_0564_));
 sg13g2_o21ai_1 _2978_ (.B1(net838),
    .Y(_0565_),
    .A1(net509),
    .A2(net751));
 sg13g2_a21oi_1 _2979_ (.A1(_1376_),
    .A2(net751),
    .Y(_0126_),
    .B1(_0565_));
 sg13g2_o21ai_1 _2980_ (.B1(net842),
    .Y(_0566_),
    .A1(net467),
    .A2(net752));
 sg13g2_a21oi_1 _2981_ (.A1(_1375_),
    .A2(net752),
    .Y(_0127_),
    .B1(_0566_));
 sg13g2_o21ai_1 _2982_ (.B1(net858),
    .Y(_0567_),
    .A1(net587),
    .A2(net753));
 sg13g2_a21oi_1 _2983_ (.A1(_1374_),
    .A2(net753),
    .Y(_0128_),
    .B1(_0567_));
 sg13g2_o21ai_1 _2984_ (.B1(net852),
    .Y(_0568_),
    .A1(net576),
    .A2(net754));
 sg13g2_a21oi_1 _2985_ (.A1(_1373_),
    .A2(net754),
    .Y(_0129_),
    .B1(_0568_));
 sg13g2_o21ai_1 _2986_ (.B1(net854),
    .Y(_0569_),
    .A1(net549),
    .A2(net753));
 sg13g2_a21oi_1 _2987_ (.A1(_1372_),
    .A2(net753),
    .Y(_0130_),
    .B1(_0569_));
 sg13g2_o21ai_1 _2988_ (.B1(net857),
    .Y(_0570_),
    .A1(net598),
    .A2(net754));
 sg13g2_a21oi_1 _2989_ (.A1(_1371_),
    .A2(net754),
    .Y(_0131_),
    .B1(_0570_));
 sg13g2_o21ai_1 _2990_ (.B1(net858),
    .Y(_0571_),
    .A1(net614),
    .A2(net753));
 sg13g2_a21oi_1 _2991_ (.A1(_1370_),
    .A2(net753),
    .Y(_0132_),
    .B1(_0571_));
 sg13g2_o21ai_1 _2992_ (.B1(net859),
    .Y(_0572_),
    .A1(net557),
    .A2(net753));
 sg13g2_a21oi_1 _2993_ (.A1(_1369_),
    .A2(net753),
    .Y(_0133_),
    .B1(_0572_));
 sg13g2_o21ai_1 _2994_ (.B1(net851),
    .Y(_0573_),
    .A1(net551),
    .A2(net754));
 sg13g2_a21oi_1 _2995_ (.A1(_1368_),
    .A2(net754),
    .Y(_0134_),
    .B1(_0573_));
 sg13g2_o21ai_1 _2996_ (.B1(net849),
    .Y(_0574_),
    .A1(net456),
    .A2(net752));
 sg13g2_a21oi_1 _2997_ (.A1(_1366_),
    .A2(net752),
    .Y(_0135_),
    .B1(_0574_));
 sg13g2_and4_1 _2998_ (.A(_1341_),
    .B(_1342_),
    .C(_1343_),
    .D(_0453_),
    .X(_0575_));
 sg13g2_o21ai_1 _2999_ (.B1(net841),
    .Y(_0576_),
    .A1(net592),
    .A2(net746));
 sg13g2_a21oi_1 _3000_ (.A1(_1382_),
    .A2(net746),
    .Y(_0136_),
    .B1(_0576_));
 sg13g2_o21ai_1 _3001_ (.B1(net835),
    .Y(_0577_),
    .A1(net523),
    .A2(net745));
 sg13g2_a21oi_1 _3002_ (.A1(_1381_),
    .A2(net745),
    .Y(_0137_),
    .B1(_0577_));
 sg13g2_o21ai_1 _3003_ (.B1(net834),
    .Y(_0578_),
    .A1(net515),
    .A2(net745));
 sg13g2_a21oi_1 _3004_ (.A1(_1380_),
    .A2(net745),
    .Y(_0138_),
    .B1(_0578_));
 sg13g2_o21ai_1 _3005_ (.B1(net834),
    .Y(_0579_),
    .A1(net542),
    .A2(net745));
 sg13g2_a21oi_1 _3006_ (.A1(_1379_),
    .A2(net745),
    .Y(_0139_),
    .B1(_0579_));
 sg13g2_o21ai_1 _3007_ (.B1(net840),
    .Y(_0580_),
    .A1(net534),
    .A2(net746));
 sg13g2_a21oi_1 _3008_ (.A1(_1378_),
    .A2(net746),
    .Y(_0140_),
    .B1(_0580_));
 sg13g2_o21ai_1 _3009_ (.B1(net839),
    .Y(_0581_),
    .A1(net572),
    .A2(net746));
 sg13g2_a21oi_1 _3010_ (.A1(_1377_),
    .A2(net746),
    .Y(_0141_),
    .B1(_0581_));
 sg13g2_o21ai_1 _3011_ (.B1(net838),
    .Y(_0582_),
    .A1(net505),
    .A2(net745));
 sg13g2_a21oi_1 _3012_ (.A1(_1376_),
    .A2(net745),
    .Y(_0142_),
    .B1(_0582_));
 sg13g2_o21ai_1 _3013_ (.B1(net842),
    .Y(_0583_),
    .A1(net493),
    .A2(net746));
 sg13g2_a21oi_1 _3014_ (.A1(_1375_),
    .A2(net746),
    .Y(_0143_),
    .B1(_0583_));
 sg13g2_o21ai_1 _3015_ (.B1(net858),
    .Y(_0584_),
    .A1(net579),
    .A2(net748));
 sg13g2_a21oi_1 _3016_ (.A1(_1374_),
    .A2(net749),
    .Y(_0144_),
    .B1(_0584_));
 sg13g2_o21ai_1 _3017_ (.B1(net849),
    .Y(_0585_),
    .A1(net616),
    .A2(net748));
 sg13g2_a21oi_1 _3018_ (.A1(_1373_),
    .A2(net748),
    .Y(_0145_),
    .B1(_0585_));
 sg13g2_o21ai_1 _3019_ (.B1(net854),
    .Y(_0586_),
    .A1(net620),
    .A2(net747));
 sg13g2_a21oi_1 _3020_ (.A1(_1372_),
    .A2(net747),
    .Y(_0146_),
    .B1(_0586_));
 sg13g2_o21ai_1 _3021_ (.B1(net857),
    .Y(_0587_),
    .A1(net479),
    .A2(net747));
 sg13g2_a21oi_1 _3022_ (.A1(_1371_),
    .A2(net747),
    .Y(_0147_),
    .B1(_0587_));
 sg13g2_o21ai_1 _3023_ (.B1(net858),
    .Y(_0588_),
    .A1(net594),
    .A2(net747));
 sg13g2_a21oi_1 _3024_ (.A1(_1370_),
    .A2(net747),
    .Y(_0148_),
    .B1(_0588_));
 sg13g2_o21ai_1 _3025_ (.B1(net859),
    .Y(_0589_),
    .A1(net450),
    .A2(net747));
 sg13g2_a21oi_1 _3026_ (.A1(_1369_),
    .A2(net747),
    .Y(_0149_),
    .B1(_0589_));
 sg13g2_o21ai_1 _3027_ (.B1(net852),
    .Y(_0590_),
    .A1(net563),
    .A2(net748));
 sg13g2_a21oi_1 _3028_ (.A1(_1368_),
    .A2(net748),
    .Y(_0150_),
    .B1(_0590_));
 sg13g2_o21ai_1 _3029_ (.B1(net849),
    .Y(_0591_),
    .A1(net477),
    .A2(net748));
 sg13g2_a21oi_1 _3030_ (.A1(_1366_),
    .A2(net748),
    .Y(_0151_),
    .B1(_0591_));
 sg13g2_nor3_1 _3031_ (.A(_1341_),
    .B(_1451_),
    .C(_1595_),
    .Y(_0592_));
 sg13g2_nand3_1 _3032_ (.B(\bitty_inst.cpu_inst.cur_state[0] ),
    .C(net793),
    .A(\bitty_inst.cpu_inst.d_inst[15] ),
    .Y(_0593_));
 sg13g2_nor2b_2 _3033_ (.A(net801),
    .B_N(\bitty_inst.cpu_inst.d_inst[0] ),
    .Y(_0594_));
 sg13g2_nor4_2 _3034_ (.A(_0052_),
    .B(_0033_),
    .C(_1595_),
    .Y(_0595_),
    .D(_0594_));
 sg13g2_or4_2 _3035_ (.A(_0052_),
    .B(_0033_),
    .C(_1595_),
    .D(_0594_),
    .X(_0596_));
 sg13g2_nand3b_1 _3036_ (.B(\bitty_inst.cpu_inst.d_inst[0] ),
    .C(net807),
    .Y(_0597_),
    .A_N(net801));
 sg13g2_nor2_1 _3037_ (.A(net807),
    .B(\bitty_inst.cpu_inst.cur_state[0] ),
    .Y(_0598_));
 sg13g2_or2_1 _3038_ (.X(_0599_),
    .B(\bitty_inst.cpu_inst.cur_state[0] ),
    .A(net807));
 sg13g2_and3_1 _3039_ (.X(_0600_),
    .A(net793),
    .B(_0597_),
    .C(_0599_));
 sg13g2_nand3_1 _3040_ (.B(_0597_),
    .C(_0599_),
    .A(net793),
    .Y(_0601_));
 sg13g2_a21oi_2 _3041_ (.B1(_0601_),
    .Y(_0602_),
    .A2(_0596_),
    .A1(_0593_));
 sg13g2_o21ai_1 _3042_ (.B1(_0600_),
    .Y(_0603_),
    .A1(_0592_),
    .A2(_0595_));
 sg13g2_a21oi_1 _3043_ (.A1(_1346_),
    .A2(net793),
    .Y(_0604_),
    .B1(_0594_));
 sg13g2_a21oi_1 _3044_ (.A1(_1343_),
    .A2(net793),
    .Y(_0605_),
    .B1(_1451_));
 sg13g2_a21oi_2 _3045_ (.B1(_0605_),
    .Y(_0606_),
    .A2(_0604_),
    .A1(net807));
 sg13g2_a21o_1 _3046_ (.A2(_0604_),
    .A1(net807),
    .B1(_0605_),
    .X(_0607_));
 sg13g2_nand3_1 _3047_ (.B(\bitty_inst.cpu_inst.cur_state[0] ),
    .C(net793),
    .A(\bitty_inst.cpu_inst.d_inst[14] ),
    .Y(_0608_));
 sg13g2_or4_2 _3048_ (.A(_0034_),
    .B(_0052_),
    .C(_1595_),
    .D(_0594_),
    .X(_0609_));
 sg13g2_and2_1 _3049_ (.A(_0608_),
    .B(_0609_),
    .X(_0610_));
 sg13g2_nand2_1 _3050_ (.Y(_0611_),
    .A(_0608_),
    .B(_0609_));
 sg13g2_nor3_1 _3051_ (.A(net743),
    .B(net739),
    .C(net735),
    .Y(_0612_));
 sg13g2_nor3_2 _3052_ (.A(net743),
    .B(net742),
    .C(net737),
    .Y(_0613_));
 sg13g2_nor3_2 _3053_ (.A(_0592_),
    .B(_0595_),
    .C(_0601_),
    .Y(_0614_));
 sg13g2_nand3_1 _3054_ (.B(_0596_),
    .C(_0600_),
    .A(_0593_),
    .Y(_0615_));
 sg13g2_nor3_1 _3055_ (.A(net739),
    .B(net735),
    .C(_0615_),
    .Y(_0616_));
 sg13g2_nor3_2 _3056_ (.A(net742),
    .B(net737),
    .C(_0615_),
    .Y(_0617_));
 sg13g2_a22oi_1 _3057_ (.Y(_0618_),
    .B1(net714),
    .B2(\bitty_inst.gen_dff[0].reg_out.mux_out[15] ),
    .A2(net717),
    .A1(\bitty_inst.gen_dff[4].reg_out.mux_out[15] ));
 sg13g2_a22oi_1 _3058_ (.Y(_0619_),
    .B1(net712),
    .B2(\bitty_inst.gen_dff[3].reg_out.mux_out[15] ),
    .A2(net716),
    .A1(\bitty_inst.gen_dff[7].reg_out.mux_out[15] ));
 sg13g2_a21oi_2 _3059_ (.B1(_0598_),
    .Y(_0620_),
    .A2(_0609_),
    .A1(_0608_));
 sg13g2_a21o_2 _3060_ (.A2(_0609_),
    .A1(_0608_),
    .B1(_0598_),
    .X(_0621_));
 sg13g2_nor3_1 _3061_ (.A(net743),
    .B(net739),
    .C(_0621_),
    .Y(_0622_));
 sg13g2_nor3_2 _3062_ (.A(net743),
    .B(net742),
    .C(_0620_),
    .Y(_0623_));
 sg13g2_nor3_2 _3063_ (.A(net739),
    .B(_0615_),
    .C(_0621_),
    .Y(_0624_));
 sg13g2_nor3_2 _3064_ (.A(net742),
    .B(_0615_),
    .C(_0620_),
    .Y(_0625_));
 sg13g2_a22oi_1 _3065_ (.Y(_0626_),
    .B1(net704),
    .B2(\bitty_inst.gen_dff[1].reg_out.mux_out[15] ),
    .A2(net706),
    .A1(\bitty_inst.gen_dff[2].reg_out.mux_out[15] ));
 sg13g2_nand3_1 _3066_ (.B(_0619_),
    .C(_0626_),
    .A(_0618_),
    .Y(_0627_));
 sg13g2_a221oi_1 _3067_ (.B2(\bitty_inst.gen_dff[5].reg_out.mux_out[15] ),
    .C1(_0627_),
    .B1(net709),
    .A1(\bitty_inst.gen_dff[6].reg_out.mux_out[15] ),
    .Y(_0628_),
    .A2(net711));
 sg13g2_nand2_1 _3068_ (.Y(_0629_),
    .A(_0036_),
    .B(_0628_));
 sg13g2_o21ai_1 _3069_ (.B1(_0629_),
    .Y(_0630_),
    .A1(_1357_),
    .A2(_0628_));
 sg13g2_a22oi_1 _3070_ (.Y(_0631_),
    .B1(net713),
    .B2(\bitty_inst.gen_dff[3].reg_out.mux_out[14] ),
    .A2(net718),
    .A1(\bitty_inst.gen_dff[4].reg_out.mux_out[14] ));
 sg13g2_a22oi_1 _3071_ (.Y(_0632_),
    .B1(net715),
    .B2(\bitty_inst.gen_dff[0].reg_out.mux_out[14] ),
    .A2(_0613_),
    .A1(\bitty_inst.gen_dff[7].reg_out.mux_out[14] ));
 sg13g2_a22oi_1 _3072_ (.Y(_0633_),
    .B1(net705),
    .B2(\bitty_inst.gen_dff[1].reg_out.mux_out[14] ),
    .A2(net709),
    .A1(\bitty_inst.gen_dff[5].reg_out.mux_out[14] ));
 sg13g2_nand3_1 _3073_ (.B(_0632_),
    .C(_0633_),
    .A(_0631_),
    .Y(_0634_));
 sg13g2_a221oi_1 _3074_ (.B2(\bitty_inst.gen_dff[2].reg_out.mux_out[14] ),
    .C1(_0634_),
    .B1(net707),
    .A1(\bitty_inst.gen_dff[6].reg_out.mux_out[14] ),
    .Y(_0635_),
    .A2(net711));
 sg13g2_inv_1 _3075_ (.Y(_0636_),
    .A(_0635_));
 sg13g2_mux2_1 _3076_ (.A0(\bitty_inst.alu_inst.in_a[14] ),
    .A1(_0037_),
    .S(_0635_),
    .X(_0637_));
 sg13g2_nand2_1 _3077_ (.Y(_0638_),
    .A(_0630_),
    .B(_0637_));
 sg13g2_a22oi_1 _3078_ (.Y(_0639_),
    .B1(_0613_),
    .B2(\bitty_inst.gen_dff[7].reg_out.mux_out[13] ),
    .A2(net718),
    .A1(\bitty_inst.gen_dff[4].reg_out.mux_out[13] ));
 sg13g2_a22oi_1 _3079_ (.Y(_0640_),
    .B1(net713),
    .B2(\bitty_inst.gen_dff[3].reg_out.mux_out[13] ),
    .A2(net715),
    .A1(\bitty_inst.gen_dff[0].reg_out.mux_out[13] ));
 sg13g2_a22oi_1 _3080_ (.Y(_0641_),
    .B1(net707),
    .B2(\bitty_inst.gen_dff[2].reg_out.mux_out[13] ),
    .A2(net709),
    .A1(\bitty_inst.gen_dff[5].reg_out.mux_out[13] ));
 sg13g2_nand3_1 _3081_ (.B(_0640_),
    .C(_0641_),
    .A(_0639_),
    .Y(_0642_));
 sg13g2_a221oi_1 _3082_ (.B2(\bitty_inst.gen_dff[1].reg_out.mux_out[13] ),
    .C1(_0642_),
    .B1(net705),
    .A1(\bitty_inst.gen_dff[6].reg_out.mux_out[13] ),
    .Y(_0643_),
    .A2(net711));
 sg13g2_inv_1 _3083_ (.Y(_0644_),
    .A(_0643_));
 sg13g2_mux2_1 _3084_ (.A0(\bitty_inst.alu_inst.in_a[13] ),
    .A1(_0038_),
    .S(_0643_),
    .X(_0645_));
 sg13g2_a22oi_1 _3085_ (.Y(_0646_),
    .B1(net713),
    .B2(\bitty_inst.gen_dff[3].reg_out.mux_out[12] ),
    .A2(net716),
    .A1(\bitty_inst.gen_dff[7].reg_out.mux_out[12] ));
 sg13g2_a22oi_1 _3086_ (.Y(_0647_),
    .B1(net715),
    .B2(\bitty_inst.gen_dff[0].reg_out.mux_out[12] ),
    .A2(net718),
    .A1(\bitty_inst.gen_dff[4].reg_out.mux_out[12] ));
 sg13g2_a22oi_1 _3087_ (.Y(_0648_),
    .B1(net707),
    .B2(\bitty_inst.gen_dff[2].reg_out.mux_out[12] ),
    .A2(net711),
    .A1(\bitty_inst.gen_dff[6].reg_out.mux_out[12] ));
 sg13g2_nand3_1 _3088_ (.B(_0647_),
    .C(_0648_),
    .A(_0646_),
    .Y(_0649_));
 sg13g2_a221oi_1 _3089_ (.B2(\bitty_inst.gen_dff[1].reg_out.mux_out[12] ),
    .C1(_0649_),
    .B1(net705),
    .A1(\bitty_inst.gen_dff[5].reg_out.mux_out[12] ),
    .Y(_0650_),
    .A2(net708));
 sg13g2_inv_1 _3090_ (.Y(_0651_),
    .A(_0650_));
 sg13g2_nor2_1 _3091_ (.A(\bitty_inst.alu_inst.in_a[12] ),
    .B(_0650_),
    .Y(_0652_));
 sg13g2_a22oi_1 _3092_ (.Y(_0653_),
    .B1(_0645_),
    .B2(_0652_),
    .A2(_0644_),
    .A1(net803));
 sg13g2_nor2_1 _3093_ (.A(_0638_),
    .B(_0653_),
    .Y(_0654_));
 sg13g2_nand3_1 _3094_ (.B(_0630_),
    .C(_0636_),
    .A(net802),
    .Y(_0655_));
 sg13g2_o21ai_1 _3095_ (.B1(_0655_),
    .Y(_0656_),
    .A1(\bitty_inst.alu_inst.in_a[15] ),
    .A2(_0628_));
 sg13g2_nor2_1 _3096_ (.A(_0654_),
    .B(_0656_),
    .Y(_0657_));
 sg13g2_mux2_1 _3097_ (.A0(\bitty_inst.alu_inst.in_a[12] ),
    .A1(_0039_),
    .S(_0650_),
    .X(_0658_));
 sg13g2_nand4_1 _3098_ (.B(_0637_),
    .C(_0645_),
    .A(_0630_),
    .Y(_0659_),
    .D(_0658_));
 sg13g2_a22oi_1 _3099_ (.Y(_0660_),
    .B1(net713),
    .B2(\bitty_inst.gen_dff[3].reg_out.mux_out[11] ),
    .A2(net718),
    .A1(\bitty_inst.gen_dff[4].reg_out.mux_out[11] ));
 sg13g2_a22oi_1 _3100_ (.Y(_0661_),
    .B1(net715),
    .B2(\bitty_inst.gen_dff[0].reg_out.mux_out[11] ),
    .A2(net716),
    .A1(\bitty_inst.gen_dff[7].reg_out.mux_out[11] ));
 sg13g2_a22oi_1 _3101_ (.Y(_0662_),
    .B1(net705),
    .B2(\bitty_inst.gen_dff[1].reg_out.mux_out[11] ),
    .A2(net707),
    .A1(\bitty_inst.gen_dff[2].reg_out.mux_out[11] ));
 sg13g2_nand3_1 _3102_ (.B(_0661_),
    .C(_0662_),
    .A(_0660_),
    .Y(_0663_));
 sg13g2_a221oi_1 _3103_ (.B2(\bitty_inst.gen_dff[5].reg_out.mux_out[11] ),
    .C1(_0663_),
    .B1(net709),
    .A1(\bitty_inst.gen_dff[6].reg_out.mux_out[11] ),
    .Y(_0664_),
    .A2(net710));
 sg13g2_inv_1 _3104_ (.Y(_0665_),
    .A(_0664_));
 sg13g2_nor2b_1 _3105_ (.A(_0664_),
    .B_N(\bitty_inst.alu_inst.in_a[11] ),
    .Y(_0666_));
 sg13g2_a21o_1 _3106_ (.A2(_0664_),
    .A1(_0040_),
    .B1(_0666_),
    .X(_0667_));
 sg13g2_a22oi_1 _3107_ (.Y(_0668_),
    .B1(net713),
    .B2(\bitty_inst.gen_dff[3].reg_out.mux_out[10] ),
    .A2(net716),
    .A1(\bitty_inst.gen_dff[7].reg_out.mux_out[10] ));
 sg13g2_a22oi_1 _3108_ (.Y(_0669_),
    .B1(net714),
    .B2(\bitty_inst.gen_dff[0].reg_out.mux_out[10] ),
    .A2(net718),
    .A1(\bitty_inst.gen_dff[4].reg_out.mux_out[10] ));
 sg13g2_a22oi_1 _3109_ (.Y(_0670_),
    .B1(net708),
    .B2(\bitty_inst.gen_dff[5].reg_out.mux_out[10] ),
    .A2(net710),
    .A1(\bitty_inst.gen_dff[6].reg_out.mux_out[10] ));
 sg13g2_nand3_1 _3110_ (.B(_0669_),
    .C(_0670_),
    .A(_0668_),
    .Y(_0671_));
 sg13g2_a221oi_1 _3111_ (.B2(\bitty_inst.gen_dff[1].reg_out.mux_out[10] ),
    .C1(_0671_),
    .B1(net705),
    .A1(\bitty_inst.gen_dff[2].reg_out.mux_out[10] ),
    .Y(_0672_),
    .A2(net707));
 sg13g2_nand2_1 _3112_ (.Y(_0673_),
    .A(_0041_),
    .B(net663));
 sg13g2_o21ai_1 _3113_ (.B1(_0673_),
    .Y(_0674_),
    .A1(_1358_),
    .A2(net663));
 sg13g2_nand2_1 _3114_ (.Y(_0675_),
    .A(_0667_),
    .B(_0674_));
 sg13g2_a22oi_1 _3115_ (.Y(_0676_),
    .B1(net712),
    .B2(\bitty_inst.gen_dff[3].reg_out.mux_out[9] ),
    .A2(net717),
    .A1(\bitty_inst.gen_dff[4].reg_out.mux_out[9] ));
 sg13g2_a22oi_1 _3116_ (.Y(_0677_),
    .B1(net714),
    .B2(\bitty_inst.gen_dff[0].reg_out.mux_out[9] ),
    .A2(net716),
    .A1(\bitty_inst.gen_dff[7].reg_out.mux_out[9] ));
 sg13g2_and2_1 _3117_ (.A(_0676_),
    .B(_0677_),
    .X(_0678_));
 sg13g2_a22oi_1 _3118_ (.Y(_0679_),
    .B1(net705),
    .B2(\bitty_inst.gen_dff[1].reg_out.mux_out[9] ),
    .A2(net706),
    .A1(\bitty_inst.gen_dff[2].reg_out.mux_out[9] ));
 sg13g2_a22oi_1 _3119_ (.Y(_0680_),
    .B1(net708),
    .B2(\bitty_inst.gen_dff[5].reg_out.mux_out[9] ),
    .A2(net711),
    .A1(\bitty_inst.gen_dff[6].reg_out.mux_out[9] ));
 sg13g2_and3_2 _3120_ (.X(_0681_),
    .A(_0678_),
    .B(_0679_),
    .C(_0680_));
 sg13g2_nand2_1 _3121_ (.Y(_0682_),
    .A(_0042_),
    .B(net662));
 sg13g2_o21ai_1 _3122_ (.B1(_0682_),
    .Y(_0683_),
    .A1(_1359_),
    .A2(net662));
 sg13g2_a22oi_1 _3123_ (.Y(_0684_),
    .B1(net712),
    .B2(\bitty_inst.gen_dff[3].reg_out.mux_out[8] ),
    .A2(net716),
    .A1(\bitty_inst.gen_dff[7].reg_out.mux_out[8] ));
 sg13g2_a22oi_1 _3124_ (.Y(_0685_),
    .B1(net714),
    .B2(\bitty_inst.gen_dff[0].reg_out.mux_out[8] ),
    .A2(net717),
    .A1(\bitty_inst.gen_dff[4].reg_out.mux_out[8] ));
 sg13g2_a22oi_1 _3125_ (.Y(_0686_),
    .B1(net709),
    .B2(\bitty_inst.gen_dff[5].reg_out.mux_out[8] ),
    .A2(net710),
    .A1(\bitty_inst.gen_dff[6].reg_out.mux_out[8] ));
 sg13g2_nand3_1 _3126_ (.B(_0685_),
    .C(_0686_),
    .A(_0684_),
    .Y(_0687_));
 sg13g2_a221oi_1 _3127_ (.B2(\bitty_inst.gen_dff[1].reg_out.mux_out[8] ),
    .C1(_0687_),
    .B1(net705),
    .A1(\bitty_inst.gen_dff[2].reg_out.mux_out[8] ),
    .Y(_0688_),
    .A2(net707));
 sg13g2_inv_1 _3128_ (.Y(_0689_),
    .A(_0688_));
 sg13g2_nand3_1 _3129_ (.B(_0683_),
    .C(_0689_),
    .A(_0043_),
    .Y(_0690_));
 sg13g2_o21ai_1 _3130_ (.B1(_0690_),
    .Y(_0691_),
    .A1(_1455_),
    .A2(net662));
 sg13g2_nor2b_1 _3131_ (.A(_0675_),
    .B_N(_0691_),
    .Y(_0692_));
 sg13g2_nor2b_1 _3132_ (.A(net663),
    .B_N(net806),
    .Y(_0693_));
 sg13g2_a221oi_1 _3133_ (.B2(_0693_),
    .C1(_0692_),
    .B1(_0667_),
    .A1(_0040_),
    .Y(_0694_),
    .A2(_0665_));
 sg13g2_a22oi_1 _3134_ (.Y(_0695_),
    .B1(net704),
    .B2(\bitty_inst.gen_dff[1].reg_out.mux_out[7] ),
    .A2(net708),
    .A1(\bitty_inst.gen_dff[5].reg_out.mux_out[7] ));
 sg13g2_nand3_1 _3135_ (.B(_0596_),
    .C(_0599_),
    .A(_0593_),
    .Y(_0696_));
 sg13g2_nor4_2 _3136_ (.A(_0600_),
    .B(net739),
    .C(_0611_),
    .Y(_0697_),
    .D(_0696_));
 sg13g2_nand2_1 _3137_ (.Y(_0698_),
    .A(\bitty_inst.gen_dff[3].reg_out.mux_out[7] ),
    .B(net712));
 sg13g2_nor4_1 _3138_ (.A(_1423_),
    .B(net743),
    .C(net742),
    .D(net737),
    .Y(_0699_));
 sg13g2_nor4_1 _3139_ (.A(_1407_),
    .B(net743),
    .C(net739),
    .D(_0621_),
    .Y(_0700_));
 sg13g2_a221oi_1 _3140_ (.B2(\bitty_inst.gen_dff[0].reg_out.mux_out[7] ),
    .C1(_0699_),
    .B1(net714),
    .A1(\bitty_inst.gen_dff[4].reg_out.mux_out[7] ),
    .Y(_0701_),
    .A2(net717));
 sg13g2_a221oi_1 _3141_ (.B2(_1452_),
    .C1(_0700_),
    .B1(_0697_),
    .A1(\bitty_inst.gen_dff[2].reg_out.mux_out[7] ),
    .Y(_0702_),
    .A2(net706));
 sg13g2_and4_2 _3142_ (.A(_0695_),
    .B(_0698_),
    .C(_0701_),
    .D(_0702_),
    .X(_0703_));
 sg13g2_nand4_1 _3143_ (.B(_0698_),
    .C(_0701_),
    .A(_0695_),
    .Y(_0704_),
    .D(_0702_));
 sg13g2_nand2_1 _3144_ (.Y(_0705_),
    .A(\bitty_inst.alu_inst.in_a[7] ),
    .B(_0704_));
 sg13g2_o21ai_1 _3145_ (.B1(_0705_),
    .Y(_0706_),
    .A1(_1456_),
    .A2(_0704_));
 sg13g2_nand4_1 _3146_ (.B(_0602_),
    .C(net738),
    .A(\bitty_inst.gen_dff[7].reg_out.mux_out[6] ),
    .Y(_0707_),
    .D(net735));
 sg13g2_nand4_1 _3147_ (.B(net744),
    .C(net740),
    .A(\bitty_inst.gen_dff[4].reg_out.mux_out[6] ),
    .Y(_0708_),
    .D(net736));
 sg13g2_nand4_1 _3148_ (.B(net738),
    .C(net735),
    .A(\bitty_inst.gen_dff[3].reg_out.mux_out[6] ),
    .Y(_0709_),
    .D(_0614_));
 sg13g2_nand2b_1 _3149_ (.Y(_0710_),
    .B(_0697_),
    .A_N(_0034_));
 sg13g2_nand4_1 _3150_ (.B(net741),
    .C(net736),
    .A(\bitty_inst.gen_dff[0].reg_out.mux_out[6] ),
    .Y(_0711_),
    .D(_0614_));
 sg13g2_a22oi_1 _3151_ (.Y(_0712_),
    .B1(net706),
    .B2(\bitty_inst.gen_dff[2].reg_out.mux_out[6] ),
    .A2(net708),
    .A1(\bitty_inst.gen_dff[5].reg_out.mux_out[6] ));
 sg13g2_a22oi_1 _3152_ (.Y(_0713_),
    .B1(net704),
    .B2(\bitty_inst.gen_dff[1].reg_out.mux_out[6] ),
    .A2(net710),
    .A1(\bitty_inst.gen_dff[6].reg_out.mux_out[6] ));
 sg13g2_and4_1 _3153_ (.A(_0707_),
    .B(_0708_),
    .C(_0709_),
    .D(_0711_),
    .X(_0714_));
 sg13g2_and4_2 _3154_ (.A(_0710_),
    .B(_0712_),
    .C(_0713_),
    .D(_0714_),
    .X(_0715_));
 sg13g2_nand2_1 _3155_ (.Y(_0716_),
    .A(_0045_),
    .B(net694));
 sg13g2_o21ai_1 _3156_ (.B1(_0716_),
    .Y(_0717_),
    .A1(_1361_),
    .A2(net695));
 sg13g2_and2_1 _3157_ (.A(_0706_),
    .B(_0717_),
    .X(_0718_));
 sg13g2_nand2_1 _3158_ (.Y(_0719_),
    .A(\bitty_inst.cpu_inst.d_inst[10] ),
    .B(_0697_));
 sg13g2_a22oi_1 _3159_ (.Y(_0720_),
    .B1(net714),
    .B2(\bitty_inst.gen_dff[0].reg_out.mux_out[5] ),
    .A2(net717),
    .A1(\bitty_inst.gen_dff[4].reg_out.mux_out[5] ));
 sg13g2_a22oi_1 _3160_ (.Y(_0721_),
    .B1(net710),
    .B2(\bitty_inst.gen_dff[6].reg_out.mux_out[5] ),
    .A2(net712),
    .A1(\bitty_inst.gen_dff[3].reg_out.mux_out[5] ));
 sg13g2_a22oi_1 _3161_ (.Y(_0722_),
    .B1(net706),
    .B2(\bitty_inst.gen_dff[2].reg_out.mux_out[5] ),
    .A2(net716),
    .A1(\bitty_inst.gen_dff[7].reg_out.mux_out[5] ));
 sg13g2_a22oi_1 _3162_ (.Y(_0723_),
    .B1(net704),
    .B2(\bitty_inst.gen_dff[1].reg_out.mux_out[5] ),
    .A2(net708),
    .A1(\bitty_inst.gen_dff[5].reg_out.mux_out[5] ));
 sg13g2_and3_1 _3163_ (.X(_0724_),
    .A(_0720_),
    .B(_0722_),
    .C(_0723_));
 sg13g2_and3_2 _3164_ (.X(_0725_),
    .A(_0719_),
    .B(_0721_),
    .C(_0724_));
 sg13g2_nand2_1 _3165_ (.Y(_0726_),
    .A(_0046_),
    .B(net660));
 sg13g2_o21ai_1 _3166_ (.B1(_0726_),
    .Y(_0727_),
    .A1(_1362_),
    .A2(net660));
 sg13g2_nand2_1 _3167_ (.Y(_0728_),
    .A(\bitty_inst.gen_dff[6].reg_out.mux_out[4] ),
    .B(net710));
 sg13g2_a22oi_1 _3168_ (.Y(_0729_),
    .B1(net704),
    .B2(\bitty_inst.gen_dff[1].reg_out.mux_out[4] ),
    .A2(net706),
    .A1(\bitty_inst.gen_dff[2].reg_out.mux_out[4] ));
 sg13g2_and2_1 _3169_ (.A(\bitty_inst.cpu_inst.d_inst[9] ),
    .B(_0697_),
    .X(_0730_));
 sg13g2_a221oi_1 _3170_ (.B2(\bitty_inst.gen_dff[0].reg_out.mux_out[4] ),
    .C1(_0730_),
    .B1(net714),
    .A1(\bitty_inst.gen_dff[4].reg_out.mux_out[4] ),
    .Y(_0731_),
    .A2(net717));
 sg13g2_and2_1 _3171_ (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[4] ),
    .B(net712),
    .X(_0732_));
 sg13g2_a221oi_1 _3172_ (.B2(\bitty_inst.gen_dff[5].reg_out.mux_out[4] ),
    .C1(_0732_),
    .B1(net708),
    .A1(\bitty_inst.gen_dff[7].reg_out.mux_out[4] ),
    .Y(_0733_),
    .A2(net716));
 sg13g2_and4_1 _3173_ (.A(_0728_),
    .B(_0729_),
    .C(_0731_),
    .D(_0733_),
    .X(_0734_));
 sg13g2_nand2_1 _3174_ (.Y(_0735_),
    .A(_0047_),
    .B(net658));
 sg13g2_o21ai_1 _3175_ (.B1(_0735_),
    .Y(_0736_),
    .A1(_1363_),
    .A2(net658));
 sg13g2_nand2_1 _3176_ (.Y(_0737_),
    .A(_0727_),
    .B(_0736_));
 sg13g2_nand4_1 _3177_ (.B(net740),
    .C(net736),
    .A(\bitty_inst.gen_dff[0].reg_out.mux_out[3] ),
    .Y(_0738_),
    .D(net734));
 sg13g2_nand4_1 _3178_ (.B(net738),
    .C(net735),
    .A(\bitty_inst.gen_dff[3].reg_out.mux_out[3] ),
    .Y(_0739_),
    .D(net734));
 sg13g2_nand4_1 _3179_ (.B(net744),
    .C(net738),
    .A(\bitty_inst.gen_dff[7].reg_out.mux_out[3] ),
    .Y(_0740_),
    .D(net735));
 sg13g2_nand4_1 _3180_ (.B(net744),
    .C(net740),
    .A(\bitty_inst.gen_dff[4].reg_out.mux_out[3] ),
    .Y(_0741_),
    .D(net736));
 sg13g2_nand2_1 _3181_ (.Y(_0742_),
    .A(\bitty_inst.cpu_inst.d_inst[8] ),
    .B(_0697_));
 sg13g2_a22oi_1 _3182_ (.Y(_0743_),
    .B1(net706),
    .B2(\bitty_inst.gen_dff[2].reg_out.mux_out[3] ),
    .A2(net708),
    .A1(\bitty_inst.gen_dff[5].reg_out.mux_out[3] ));
 sg13g2_a22oi_1 _3183_ (.Y(_0744_),
    .B1(net704),
    .B2(\bitty_inst.gen_dff[1].reg_out.mux_out[3] ),
    .A2(net710),
    .A1(\bitty_inst.gen_dff[6].reg_out.mux_out[3] ));
 sg13g2_and4_2 _3184_ (.A(_0738_),
    .B(_0739_),
    .C(_0740_),
    .D(_0741_),
    .X(_0745_));
 sg13g2_and4_2 _3185_ (.A(_0742_),
    .B(_0743_),
    .C(_0744_),
    .D(_0745_),
    .X(_0746_));
 sg13g2_nand4_1 _3186_ (.B(_0743_),
    .C(_0744_),
    .A(_0742_),
    .Y(_0747_),
    .D(_0745_));
 sg13g2_nand2_1 _3187_ (.Y(_0748_),
    .A(\bitty_inst.alu_inst.in_a[3] ),
    .B(net692));
 sg13g2_o21ai_1 _3188_ (.B1(_0748_),
    .Y(_0749_),
    .A1(_1458_),
    .A2(net692));
 sg13g2_nand4_1 _3189_ (.B(net744),
    .C(net738),
    .A(\bitty_inst.gen_dff[5].reg_out.mux_out[2] ),
    .Y(_0750_),
    .D(_0621_));
 sg13g2_nand4_1 _3190_ (.B(net744),
    .C(net740),
    .A(\bitty_inst.gen_dff[6].reg_out.mux_out[2] ),
    .Y(_0751_),
    .D(_0620_));
 sg13g2_nand4_1 _3191_ (.B(net738),
    .C(net734),
    .A(\bitty_inst.gen_dff[1].reg_out.mux_out[2] ),
    .Y(_0752_),
    .D(_0621_));
 sg13g2_nand3_1 _3192_ (.B(_0751_),
    .C(_0752_),
    .A(_0750_),
    .Y(_0753_));
 sg13g2_and2_1 _3193_ (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[2] ),
    .B(net717),
    .X(_0754_));
 sg13g2_and4_1 _3194_ (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[2] ),
    .B(net738),
    .C(net735),
    .D(net734),
    .X(_0755_));
 sg13g2_a21o_1 _3195_ (.A2(_0697_),
    .A1(\bitty_inst.cpu_inst.d_inst[7] ),
    .B1(_0755_),
    .X(_0756_));
 sg13g2_nand4_1 _3196_ (.B(net740),
    .C(net734),
    .A(\bitty_inst.gen_dff[2].reg_out.mux_out[2] ),
    .Y(_0757_),
    .D(_0620_));
 sg13g2_nand4_1 _3197_ (.B(net740),
    .C(net736),
    .A(\bitty_inst.gen_dff[0].reg_out.mux_out[2] ),
    .Y(_0758_),
    .D(net734));
 sg13g2_nand4_1 _3198_ (.B(net744),
    .C(net738),
    .A(\bitty_inst.gen_dff[7].reg_out.mux_out[2] ),
    .Y(_0759_),
    .D(net735));
 sg13g2_nand3_1 _3199_ (.B(_0758_),
    .C(_0759_),
    .A(_0757_),
    .Y(_0760_));
 sg13g2_nor4_2 _3200_ (.A(_0753_),
    .B(_0754_),
    .C(_0756_),
    .Y(_0761_),
    .D(_0760_));
 sg13g2_or4_1 _3201_ (.A(_0753_),
    .B(_0754_),
    .C(_0756_),
    .D(_0760_),
    .X(_0762_));
 sg13g2_mux2_1 _3202_ (.A0(\bitty_inst.alu_inst.in_a[2] ),
    .A1(_0049_),
    .S(net689),
    .X(_0763_));
 sg13g2_nand2_1 _3203_ (.Y(_0764_),
    .A(_0749_),
    .B(_0763_));
 sg13g2_nor4_1 _3204_ (.A(_1397_),
    .B(net743),
    .C(_0606_),
    .D(_0620_),
    .Y(_0765_));
 sg13g2_nand4_1 _3205_ (.B(net741),
    .C(net734),
    .A(\bitty_inst.gen_dff[2].reg_out.mux_out[1] ),
    .Y(_0766_),
    .D(_0620_));
 sg13g2_and2_1 _3206_ (.A(\bitty_inst.cpu_inst.d_inst[6] ),
    .B(_0697_),
    .X(_0767_));
 sg13g2_nand4_1 _3207_ (.B(net741),
    .C(net736),
    .A(\bitty_inst.gen_dff[0].reg_out.mux_out[1] ),
    .Y(_0768_),
    .D(net734));
 sg13g2_nand4_1 _3208_ (.B(net744),
    .C(net740),
    .A(\bitty_inst.gen_dff[6].reg_out.mux_out[1] ),
    .Y(_0769_),
    .D(_0620_));
 sg13g2_nor4_1 _3209_ (.A(_1429_),
    .B(net743),
    .C(net741),
    .D(net736),
    .Y(_0770_));
 sg13g2_nand4_1 _3210_ (.B(net744),
    .C(net740),
    .A(\bitty_inst.gen_dff[4].reg_out.mux_out[1] ),
    .Y(_0771_),
    .D(net736));
 sg13g2_a21o_1 _3211_ (.A2(net712),
    .A1(\bitty_inst.gen_dff[3].reg_out.mux_out[1] ),
    .B1(_0770_),
    .X(_0772_));
 sg13g2_a21o_1 _3212_ (.A2(net704),
    .A1(\bitty_inst.gen_dff[1].reg_out.mux_out[1] ),
    .B1(_0765_),
    .X(_0773_));
 sg13g2_nand4_1 _3213_ (.B(_0768_),
    .C(_0769_),
    .A(_0766_),
    .Y(_0774_),
    .D(_0771_));
 sg13g2_nor4_2 _3214_ (.A(_0767_),
    .B(_0772_),
    .C(_0773_),
    .Y(_0775_),
    .D(_0774_));
 sg13g2_or4_1 _3215_ (.A(_0767_),
    .B(_0772_),
    .C(_0773_),
    .D(_0774_),
    .X(_0776_));
 sg13g2_nand2_1 _3216_ (.Y(_0777_),
    .A(_0050_),
    .B(net676));
 sg13g2_nand3_1 _3217_ (.B(_0749_),
    .C(net686),
    .A(_0049_),
    .Y(_0778_));
 sg13g2_nand3b_1 _3218_ (.B(_0047_),
    .C(_0727_),
    .Y(_0779_),
    .A_N(net658));
 sg13g2_o21ai_1 _3219_ (.B1(_0779_),
    .Y(_0780_),
    .A1(_1457_),
    .A2(net660));
 sg13g2_nor4_1 _3220_ (.A(_1398_),
    .B(_0603_),
    .C(_0606_),
    .D(_0620_),
    .Y(_0781_));
 sg13g2_a221oi_1 _3221_ (.B2(\bitty_inst.gen_dff[1].reg_out.mux_out[0] ),
    .C1(_0781_),
    .B1(net704),
    .A1(\bitty_inst.gen_dff[6].reg_out.mux_out[0] ),
    .Y(_0782_),
    .A2(net710));
 sg13g2_nand2_1 _3222_ (.Y(_0783_),
    .A(\bitty_inst.cpu_inst.d_inst[5] ),
    .B(_0697_));
 sg13g2_a22oi_1 _3223_ (.Y(_0784_),
    .B1(net714),
    .B2(\bitty_inst.gen_dff[0].reg_out.mux_out[0] ),
    .A2(net717),
    .A1(\bitty_inst.gen_dff[4].reg_out.mux_out[0] ));
 sg13g2_nor4_1 _3224_ (.A(_1430_),
    .B(_0603_),
    .C(net742),
    .D(net737),
    .Y(_0785_));
 sg13g2_a221oi_1 _3225_ (.B2(\bitty_inst.gen_dff[2].reg_out.mux_out[0] ),
    .C1(_0785_),
    .B1(net706),
    .A1(\bitty_inst.gen_dff[3].reg_out.mux_out[0] ),
    .Y(_0786_),
    .A2(net712));
 sg13g2_and4_2 _3226_ (.A(_0782_),
    .B(_0783_),
    .C(_0784_),
    .D(_0786_),
    .X(_0787_));
 sg13g2_nand4_1 _3227_ (.B(_0783_),
    .C(_0784_),
    .A(_0782_),
    .Y(_0788_),
    .D(_0786_));
 sg13g2_nand2_1 _3228_ (.Y(_0789_),
    .A(_0050_),
    .B(net677));
 sg13g2_o21ai_1 _3229_ (.B1(_0789_),
    .Y(_0790_),
    .A1(_1364_),
    .A2(net677));
 sg13g2_o21ai_1 _3230_ (.B1(_0790_),
    .Y(_0791_),
    .A1(_1365_),
    .A2(net665));
 sg13g2_nor3_1 _3231_ (.A(_0737_),
    .B(_0764_),
    .C(_0791_),
    .Y(_0792_));
 sg13g2_a21oi_1 _3232_ (.A1(_0777_),
    .A2(_0791_),
    .Y(_0793_),
    .B1(_0764_));
 sg13g2_a21oi_1 _3233_ (.A1(_0048_),
    .A2(net692),
    .Y(_0794_),
    .B1(_0793_));
 sg13g2_a21oi_1 _3234_ (.A1(_0778_),
    .A2(_0794_),
    .Y(_0795_),
    .B1(_0737_));
 sg13g2_o21ai_1 _3235_ (.B1(_0718_),
    .Y(_0796_),
    .A1(_0780_),
    .A2(_0795_));
 sg13g2_nor2b_1 _3236_ (.A(net695),
    .B_N(_0045_),
    .Y(_0797_));
 sg13g2_a22oi_1 _3237_ (.Y(_0798_),
    .B1(_0706_),
    .B2(_0797_),
    .A2(_0704_),
    .A1(_0044_));
 sg13g2_nand2_1 _3238_ (.Y(_0799_),
    .A(_0796_),
    .B(_0798_));
 sg13g2_mux2_1 _3239_ (.A0(\bitty_inst.alu_inst.in_a[8] ),
    .A1(_0043_),
    .S(_0688_),
    .X(_0800_));
 sg13g2_nand2_1 _3240_ (.Y(_0801_),
    .A(_0683_),
    .B(_0800_));
 sg13g2_nor3_2 _3241_ (.A(_0659_),
    .B(_0675_),
    .C(_0801_),
    .Y(_0802_));
 sg13g2_o21ai_1 _3242_ (.B1(_0657_),
    .Y(_0803_),
    .A1(_0659_),
    .A2(_0694_));
 sg13g2_a21oi_1 _3243_ (.A1(_0799_),
    .A2(_0802_),
    .Y(_0804_),
    .B1(_0803_));
 sg13g2_nand2b_1 _3244_ (.Y(_0805_),
    .B(\bitty_inst.cpu_inst.d_inst[3] ),
    .A_N(_0052_));
 sg13g2_nand2b_2 _3245_ (.Y(_0806_),
    .B(_1596_),
    .A_N(_0805_));
 sg13g2_nor2_2 _3246_ (.A(_1513_),
    .B(_0806_),
    .Y(_0807_));
 sg13g2_nand2_2 _3247_ (.Y(_0808_),
    .A(_0051_),
    .B(net664));
 sg13g2_nand4_1 _3248_ (.B(_0792_),
    .C(_0802_),
    .A(_0718_),
    .Y(_0809_),
    .D(_0808_));
 sg13g2_nand3_1 _3249_ (.B(_0807_),
    .C(_0809_),
    .A(\bitty_inst.cpu_inst.d_inst[4] ),
    .Y(_0810_));
 sg13g2_nand4_1 _3250_ (.B(_0804_),
    .C(_0807_),
    .A(\bitty_inst.cpu_inst.d_inst[4] ),
    .Y(_0811_),
    .D(_0809_));
 sg13g2_nand2_1 _3251_ (.Y(_0812_),
    .A(_0047_),
    .B(net668));
 sg13g2_o21ai_1 _3252_ (.B1(_0812_),
    .Y(_0813_),
    .A1(_1457_),
    .A2(net669));
 sg13g2_nand2_1 _3253_ (.Y(_0814_),
    .A(_0045_),
    .B(net670));
 sg13g2_o21ai_1 _3254_ (.B1(_0814_),
    .Y(_0815_),
    .A1(_1456_),
    .A2(net669));
 sg13g2_mux2_1 _3255_ (.A0(_0813_),
    .A1(_0815_),
    .S(net674),
    .X(_0816_));
 sg13g2_nand2_1 _3256_ (.Y(_0817_),
    .A(net683),
    .B(_0816_));
 sg13g2_nor2_1 _3257_ (.A(_1512_),
    .B(_0806_),
    .Y(_0818_));
 sg13g2_nand3_1 _3258_ (.B(net808),
    .C(net793),
    .A(\bitty_inst.cpu_inst.d_inst[4] ),
    .Y(_0819_));
 sg13g2_nor3_2 _3259_ (.A(_1512_),
    .B(_0806_),
    .C(_0819_),
    .Y(_0820_));
 sg13g2_nand3_1 _3260_ (.B(net808),
    .C(_0818_),
    .A(\bitty_inst.cpu_inst.d_inst[4] ),
    .Y(_0821_));
 sg13g2_nor2_2 _3261_ (.A(net690),
    .B(_0821_),
    .Y(_0822_));
 sg13g2_nand2_2 _3262_ (.Y(_0823_),
    .A(_0746_),
    .B(_0820_));
 sg13g2_nand2_1 _3263_ (.Y(_0824_),
    .A(_0051_),
    .B(net673));
 sg13g2_and2_1 _3264_ (.A(_0050_),
    .B(net664),
    .X(_0825_));
 sg13g2_nor2_1 _3265_ (.A(net675),
    .B(_0825_),
    .Y(_0826_));
 sg13g2_nand2_1 _3266_ (.Y(_0827_),
    .A(_0049_),
    .B(net673));
 sg13g2_o21ai_1 _3267_ (.B1(_0827_),
    .Y(_0828_),
    .A1(_1458_),
    .A2(net673));
 sg13g2_o21ai_1 _3268_ (.B1(net688),
    .Y(_0829_),
    .A1(net682),
    .A2(_0828_));
 sg13g2_a21oi_1 _3269_ (.A1(_0824_),
    .A2(_0826_),
    .Y(_0830_),
    .B1(_0829_));
 sg13g2_nor2_1 _3270_ (.A(_0823_),
    .B(_0830_),
    .Y(_0831_));
 sg13g2_nand3_1 _3271_ (.B(net678),
    .C(net668),
    .A(net689),
    .Y(_0832_));
 sg13g2_nor2_1 _3272_ (.A(_0051_),
    .B(net664),
    .Y(_0833_));
 sg13g2_nor2_1 _3273_ (.A(_0051_),
    .B(_0832_),
    .Y(_0834_));
 sg13g2_nand2b_1 _3274_ (.Y(_0835_),
    .B(_0805_),
    .A_N(_0819_));
 sg13g2_nor2_2 _3275_ (.A(_0035_),
    .B(_0835_),
    .Y(_0836_));
 sg13g2_inv_2 _3276_ (.Y(_0837_),
    .A(_0836_));
 sg13g2_nor2_2 _3277_ (.A(net690),
    .B(_0837_),
    .Y(_0838_));
 sg13g2_nand2_2 _3278_ (.Y(_0839_),
    .A(_0746_),
    .B(_0836_));
 sg13g2_nand2_1 _3279_ (.Y(_0840_),
    .A(_0834_),
    .B(_0838_));
 sg13g2_nor2_2 _3280_ (.A(_1512_),
    .B(_0835_),
    .Y(_0841_));
 sg13g2_o21ai_1 _3281_ (.B1(net702),
    .Y(_0842_),
    .A1(_0051_),
    .A2(net673));
 sg13g2_nor2b_1 _3282_ (.A(_0842_),
    .B_N(_0824_),
    .Y(_0843_));
 sg13g2_nand2_2 _3283_ (.Y(_0844_),
    .A(_0818_),
    .B(_0819_));
 sg13g2_inv_2 _3284_ (.Y(_0845_),
    .A(_0844_));
 sg13g2_nor3_1 _3285_ (.A(_0051_),
    .B(net673),
    .C(net701),
    .Y(_0846_));
 sg13g2_and2_2 _3286_ (.A(_0806_),
    .B(_0819_),
    .X(_0847_));
 sg13g2_nand2_2 _3287_ (.Y(_0848_),
    .A(_0806_),
    .B(_0819_));
 sg13g2_nand2_2 _3288_ (.Y(_0849_),
    .A(_1352_),
    .B(_0807_));
 sg13g2_a21oi_1 _3289_ (.A1(_1365_),
    .A2(net668),
    .Y(_0850_),
    .B1(net699));
 sg13g2_nor4_1 _3290_ (.A(_0843_),
    .B(_0846_),
    .C(net732),
    .D(_0850_),
    .Y(_0851_));
 sg13g2_nor2_2 _3291_ (.A(net693),
    .B(_0821_),
    .Y(_0852_));
 sg13g2_mux2_1 _3292_ (.A0(_0038_),
    .A1(net804),
    .S(net671),
    .X(_0853_));
 sg13g2_nand2_1 _3293_ (.Y(_0854_),
    .A(net802),
    .B(net672));
 sg13g2_o21ai_1 _3294_ (.B1(_0854_),
    .Y(_0855_),
    .A1(_1453_),
    .A2(net671));
 sg13g2_mux2_1 _3295_ (.A0(_0853_),
    .A1(_0855_),
    .S(net674),
    .X(_0856_));
 sg13g2_nand2_1 _3296_ (.Y(_0857_),
    .A(_0043_),
    .B(net671));
 sg13g2_o21ai_1 _3297_ (.B1(_0857_),
    .Y(_0858_),
    .A1(_1455_),
    .A2(net671));
 sg13g2_nand2_1 _3298_ (.Y(_0859_),
    .A(net806),
    .B(net671));
 sg13g2_o21ai_1 _3299_ (.B1(_0859_),
    .Y(_0860_),
    .A1(_1454_),
    .A2(net671));
 sg13g2_mux2_1 _3300_ (.A0(_0858_),
    .A1(_0860_),
    .S(net674),
    .X(_0861_));
 sg13g2_mux2_1 _3301_ (.A0(_0856_),
    .A1(_0861_),
    .S(net687),
    .X(_0862_));
 sg13g2_inv_1 _3302_ (.Y(_0863_),
    .A(_0862_));
 sg13g2_a22oi_1 _3303_ (.Y(_0864_),
    .B1(_0852_),
    .B2(_0863_),
    .A2(_0831_),
    .A1(_0817_));
 sg13g2_nand4_1 _3304_ (.B(_0840_),
    .C(_0851_),
    .A(_0811_),
    .Y(_0865_),
    .D(_0864_));
 sg13g2_nor2_2 _3305_ (.A(_0052_),
    .B(_1514_),
    .Y(_0866_));
 sg13g2_or2_2 _3306_ (.X(_0867_),
    .B(_1514_),
    .A(_0052_));
 sg13g2_a21oi_1 _3307_ (.A1(\bitty_inst.alu_inst.in_a[0] ),
    .A2(net667),
    .Y(_0868_),
    .B1(net730));
 sg13g2_a21oi_1 _3308_ (.A1(_0808_),
    .A2(_0868_),
    .Y(_0869_),
    .B1(net778));
 sg13g2_a221oi_1 _3309_ (.B2(_0865_),
    .C1(net800),
    .B1(_0869_),
    .A1(\bitty_inst.data_to_ld[0] ),
    .Y(_0870_),
    .A2(net778));
 sg13g2_o21ai_1 _3310_ (.B1(net836),
    .Y(_0871_),
    .A1(net807),
    .A2(net919));
 sg13g2_nor2_1 _3311_ (.A(_0870_),
    .B(_0871_),
    .Y(_0152_));
 sg13g2_mux2_1 _3312_ (.A0(net802),
    .A1(net803),
    .S(net670),
    .X(_0872_));
 sg13g2_nand2b_1 _3313_ (.Y(_0873_),
    .B(net679),
    .A_N(_0872_));
 sg13g2_nand2_1 _3314_ (.Y(_0874_),
    .A(_1453_),
    .B(net672));
 sg13g2_o21ai_1 _3315_ (.B1(_0873_),
    .Y(_0875_),
    .A1(net681),
    .A2(_0874_));
 sg13g2_nor2_1 _3316_ (.A(net687),
    .B(_0875_),
    .Y(_0876_));
 sg13g2_nor2_1 _3317_ (.A(net806),
    .B(net673),
    .Y(_0877_));
 sg13g2_a21oi_2 _3318_ (.B1(_0877_),
    .Y(_0878_),
    .A2(net669),
    .A1(_1455_));
 sg13g2_mux2_1 _3319_ (.A0(net804),
    .A1(net805),
    .S(net670),
    .X(_0879_));
 sg13g2_mux2_1 _3320_ (.A0(_0878_),
    .A1(_0879_),
    .S(net675),
    .X(_0880_));
 sg13g2_a21oi_1 _3321_ (.A1(net689),
    .A2(_0880_),
    .Y(_0881_),
    .B1(_0876_));
 sg13g2_nand2_1 _3322_ (.Y(_0882_),
    .A(_0045_),
    .B(net665));
 sg13g2_o21ai_1 _3323_ (.B1(_0882_),
    .Y(_0883_),
    .A1(_1457_),
    .A2(net665));
 sg13g2_nor2_1 _3324_ (.A(_0043_),
    .B(net669),
    .Y(_0884_));
 sg13g2_a21oi_2 _3325_ (.B1(_0884_),
    .Y(_0885_),
    .A2(net669),
    .A1(_1456_));
 sg13g2_mux2_1 _3326_ (.A0(_0883_),
    .A1(_0885_),
    .S(net676),
    .X(_0886_));
 sg13g2_nand2_1 _3327_ (.Y(_0887_),
    .A(net683),
    .B(_0886_));
 sg13g2_nand2_1 _3328_ (.Y(_0888_),
    .A(_0047_),
    .B(net665));
 sg13g2_o21ai_1 _3329_ (.B1(_0888_),
    .Y(_0889_),
    .A1(_1458_),
    .A2(net665));
 sg13g2_nor2_1 _3330_ (.A(net678),
    .B(_0889_),
    .Y(_0890_));
 sg13g2_nand2_1 _3331_ (.Y(_0891_),
    .A(_0049_),
    .B(net664));
 sg13g2_nand2_1 _3332_ (.Y(_0892_),
    .A(_0050_),
    .B(net667));
 sg13g2_nand3_1 _3333_ (.B(_0891_),
    .C(_0892_),
    .A(net682),
    .Y(_0893_));
 sg13g2_nor2_1 _3334_ (.A(net686),
    .B(_0890_),
    .Y(_0894_));
 sg13g2_a21oi_1 _3335_ (.A1(_0893_),
    .A2(_0894_),
    .Y(_0895_),
    .B1(_0823_));
 sg13g2_o21ai_1 _3336_ (.B1(net702),
    .Y(_0896_),
    .A1(_0050_),
    .A2(net678));
 sg13g2_a22oi_1 _3337_ (.Y(_0897_),
    .B1(net699),
    .B2(_0896_),
    .A2(net678),
    .A1(_0050_));
 sg13g2_nand2_1 _3338_ (.Y(_0898_),
    .A(_0808_),
    .B(_0892_));
 sg13g2_nor2_1 _3339_ (.A(net675),
    .B(_0898_),
    .Y(_0899_));
 sg13g2_nand2_1 _3340_ (.Y(_0900_),
    .A(net689),
    .B(_0899_));
 sg13g2_nor3_1 _3341_ (.A(_1364_),
    .B(net677),
    .C(net701),
    .Y(_0901_));
 sg13g2_nor3_1 _3342_ (.A(net732),
    .B(_0897_),
    .C(_0901_),
    .Y(_0902_));
 sg13g2_o21ai_1 _3343_ (.B1(_0902_),
    .Y(_0903_),
    .A1(_0839_),
    .A2(_0900_));
 sg13g2_a221oi_1 _3344_ (.B2(_0895_),
    .C1(_0903_),
    .B1(_0887_),
    .A1(_0852_),
    .Y(_0904_),
    .A2(_0881_));
 sg13g2_o21ai_1 _3345_ (.B1(_0904_),
    .Y(_0905_),
    .A1(_0804_),
    .A2(_0810_));
 sg13g2_nor2_1 _3346_ (.A(\bitty_inst.alu_inst.in_a[0] ),
    .B(net667),
    .Y(_0906_));
 sg13g2_nor3_2 _3347_ (.A(_1513_),
    .B(_1595_),
    .C(net730),
    .Y(_0907_));
 sg13g2_nand3_1 _3348_ (.B(net793),
    .C(net732),
    .A(_1512_),
    .Y(_0908_));
 sg13g2_nor3_1 _3349_ (.A(net676),
    .B(net667),
    .C(_0907_),
    .Y(_0909_));
 sg13g2_nand3_1 _3350_ (.B(net665),
    .C(net697),
    .A(net677),
    .Y(_0910_));
 sg13g2_a21oi_1 _3351_ (.A1(net665),
    .A2(net697),
    .Y(_0911_),
    .B1(net677));
 sg13g2_o21ai_1 _3352_ (.B1(net676),
    .Y(_0912_),
    .A1(net667),
    .A2(_0907_));
 sg13g2_nor3_1 _3353_ (.A(_1364_),
    .B(_0909_),
    .C(_0911_),
    .Y(_0913_));
 sg13g2_a21oi_1 _3354_ (.A1(_0910_),
    .A2(_0912_),
    .Y(_0914_),
    .B1(\bitty_inst.alu_inst.in_a[1] ));
 sg13g2_or2_1 _3355_ (.X(_0915_),
    .B(_0914_),
    .A(_0913_));
 sg13g2_nor3_1 _3356_ (.A(_0906_),
    .B(_0913_),
    .C(_0914_),
    .Y(_0916_));
 sg13g2_xnor2_1 _3357_ (.Y(_0917_),
    .A(_0906_),
    .B(_0915_));
 sg13g2_a21oi_1 _3358_ (.A1(net732),
    .A2(_0917_),
    .Y(_0918_),
    .B1(net777));
 sg13g2_a221oi_1 _3359_ (.B2(_0918_),
    .C1(net797),
    .B1(_0905_),
    .A1(\bitty_inst.data_to_ld[1] ),
    .Y(_0919_),
    .A2(net777));
 sg13g2_o21ai_1 _3360_ (.B1(net836),
    .Y(_0920_),
    .A1(net807),
    .A2(net952));
 sg13g2_nor2_1 _3361_ (.A(_0919_),
    .B(_0920_),
    .Y(_0153_));
 sg13g2_nor3_1 _3362_ (.A(_0050_),
    .B(_0909_),
    .C(_0911_),
    .Y(_0921_));
 sg13g2_nor2_1 _3363_ (.A(_0916_),
    .B(_0921_),
    .Y(_0922_));
 sg13g2_a21oi_1 _3364_ (.A1(net677),
    .A2(net667),
    .Y(_0923_),
    .B1(_0907_));
 sg13g2_xnor2_1 _3365_ (.Y(_0924_),
    .A(net686),
    .B(_0923_));
 sg13g2_xnor2_1 _3366_ (.Y(_0925_),
    .A(_0049_),
    .B(_0924_));
 sg13g2_o21ai_1 _3367_ (.B1(_0925_),
    .Y(_0926_),
    .A1(_0916_),
    .A2(_0921_));
 sg13g2_xnor2_1 _3368_ (.Y(_0927_),
    .A(_0922_),
    .B(_0925_));
 sg13g2_mux2_1 _3369_ (.A0(_0815_),
    .A1(_0858_),
    .S(net674),
    .X(_0928_));
 sg13g2_nor2_1 _3370_ (.A(net680),
    .B(_0813_),
    .Y(_0929_));
 sg13g2_nor2_1 _3371_ (.A(net683),
    .B(_0929_),
    .Y(_0930_));
 sg13g2_o21ai_1 _3372_ (.B1(_0930_),
    .Y(_0931_),
    .A1(net674),
    .A2(_0828_));
 sg13g2_a21oi_1 _3373_ (.A1(net684),
    .A2(_0928_),
    .Y(_0932_),
    .B1(_0823_));
 sg13g2_mux2_1 _3374_ (.A0(_0853_),
    .A1(_0860_),
    .S(net681),
    .X(_0933_));
 sg13g2_nor2_1 _3375_ (.A(net688),
    .B(net674),
    .Y(_0934_));
 sg13g2_nor2_1 _3376_ (.A(net675),
    .B(_0855_),
    .Y(_0935_));
 sg13g2_nor2_1 _3377_ (.A(net687),
    .B(_0935_),
    .Y(_0936_));
 sg13g2_a21oi_1 _3378_ (.A1(net687),
    .A2(_0933_),
    .Y(_0937_),
    .B1(_0936_));
 sg13g2_nor2b_1 _3379_ (.A(_0825_),
    .B_N(_0827_),
    .Y(_0938_));
 sg13g2_mux2_1 _3380_ (.A0(_0833_),
    .A1(_0938_),
    .S(net682),
    .X(_0939_));
 sg13g2_nand2_1 _3381_ (.Y(_0940_),
    .A(net688),
    .B(_0939_));
 sg13g2_o21ai_1 _3382_ (.B1(net703),
    .Y(_0941_),
    .A1(_0049_),
    .A2(net688));
 sg13g2_a22oi_1 _3383_ (.Y(_0942_),
    .B1(net700),
    .B2(_0941_),
    .A2(net688),
    .A1(_0049_));
 sg13g2_and3_1 _3384_ (.X(_0943_),
    .A(\bitty_inst.alu_inst.in_a[2] ),
    .B(net684),
    .C(_0845_));
 sg13g2_nor3_1 _3385_ (.A(net733),
    .B(_0942_),
    .C(_0943_),
    .Y(_0944_));
 sg13g2_o21ai_1 _3386_ (.B1(_0944_),
    .Y(_0945_),
    .A1(_0839_),
    .A2(_0940_));
 sg13g2_a221oi_1 _3387_ (.B2(_0852_),
    .C1(_0945_),
    .B1(_0937_),
    .A1(_0931_),
    .Y(_0946_),
    .A2(_0932_));
 sg13g2_nor2_1 _3388_ (.A(net778),
    .B(_0946_),
    .Y(_0947_));
 sg13g2_o21ai_1 _3389_ (.B1(_0947_),
    .Y(_0948_),
    .A1(net730),
    .A2(_0927_));
 sg13g2_a21oi_1 _3390_ (.A1(\bitty_inst.data_to_ld[2] ),
    .A2(net777),
    .Y(_0949_),
    .B1(net797));
 sg13g2_a221oi_1 _3391_ (.B2(_0949_),
    .C1(net822),
    .B1(_0948_),
    .A1(net797),
    .Y(_0154_),
    .A2(_1380_));
 sg13g2_nand2_1 _3392_ (.Y(_0950_),
    .A(\bitty_inst.alu_inst.in_a[2] ),
    .B(_0924_));
 sg13g2_nand2_1 _3393_ (.Y(_0951_),
    .A(_0832_),
    .B(net697));
 sg13g2_xnor2_1 _3394_ (.Y(_0952_),
    .A(net692),
    .B(_0951_));
 sg13g2_nor2_1 _3395_ (.A(_0048_),
    .B(_0952_),
    .Y(_0953_));
 sg13g2_inv_1 _3396_ (.Y(_0954_),
    .A(_0953_));
 sg13g2_xnor2_1 _3397_ (.Y(_0955_),
    .A(_0048_),
    .B(_0952_));
 sg13g2_a21o_1 _3398_ (.A2(_0950_),
    .A1(_0926_),
    .B1(_0955_),
    .X(_0956_));
 sg13g2_nand3_1 _3399_ (.B(_0950_),
    .C(_0955_),
    .A(_0926_),
    .Y(_0957_));
 sg13g2_a21o_1 _3400_ (.A2(_0957_),
    .A1(_0956_),
    .B1(net730),
    .X(_0958_));
 sg13g2_mux2_1 _3401_ (.A0(_0878_),
    .A1(_0885_),
    .S(net679),
    .X(_0959_));
 sg13g2_nor2_1 _3402_ (.A(net689),
    .B(_0959_),
    .Y(_0960_));
 sg13g2_a21o_1 _3403_ (.A2(_0883_),
    .A1(net676),
    .B1(net686),
    .X(_0961_));
 sg13g2_a21oi_1 _3404_ (.A1(net678),
    .A2(_0889_),
    .Y(_0962_),
    .B1(_0961_));
 sg13g2_o21ai_1 _3405_ (.B1(_0822_),
    .Y(_0963_),
    .A1(_0960_),
    .A2(_0962_));
 sg13g2_nor2_2 _3406_ (.A(net675),
    .B(_0874_),
    .Y(_0964_));
 sg13g2_mux2_1 _3407_ (.A0(_0872_),
    .A1(_0879_),
    .S(net679),
    .X(_0965_));
 sg13g2_nor2_1 _3408_ (.A(net687),
    .B(_0964_),
    .Y(_0966_));
 sg13g2_a21oi_2 _3409_ (.B1(_0966_),
    .Y(_0967_),
    .A2(_0965_),
    .A1(net687));
 sg13g2_o21ai_1 _3410_ (.B1(net702),
    .Y(_0968_),
    .A1(_0048_),
    .A2(net693));
 sg13g2_a22oi_1 _3411_ (.Y(_0969_),
    .B1(net699),
    .B2(_0968_),
    .A2(net693),
    .A1(_0048_));
 sg13g2_o21ai_1 _3412_ (.B1(net730),
    .Y(_0970_),
    .A1(_0748_),
    .A2(net701));
 sg13g2_nor2_1 _3413_ (.A(_0969_),
    .B(_0970_),
    .Y(_0971_));
 sg13g2_o21ai_1 _3414_ (.B1(_0891_),
    .Y(_0972_),
    .A1(_1458_),
    .A2(net664));
 sg13g2_mux2_1 _3415_ (.A0(_0898_),
    .A1(_0972_),
    .S(net679),
    .X(_0973_));
 sg13g2_nor2_1 _3416_ (.A(net683),
    .B(_0973_),
    .Y(_0974_));
 sg13g2_a22oi_1 _3417_ (.Y(_0975_),
    .B1(_0974_),
    .B2(_0838_),
    .A2(_0967_),
    .A1(_0852_));
 sg13g2_nand3_1 _3418_ (.B(_0971_),
    .C(_0975_),
    .A(_0963_),
    .Y(_0976_));
 sg13g2_nand3_1 _3419_ (.B(_0958_),
    .C(_0976_),
    .A(net776),
    .Y(_0977_));
 sg13g2_a21oi_1 _3420_ (.A1(\bitty_inst.data_to_ld[3] ),
    .A2(net777),
    .Y(_0978_),
    .B1(net797));
 sg13g2_a221oi_1 _3421_ (.B2(_0978_),
    .C1(net822),
    .B1(_0977_),
    .A1(net797),
    .Y(_0155_),
    .A2(_1379_));
 sg13g2_and2_1 _3422_ (.A(_0954_),
    .B(_0956_),
    .X(_0979_));
 sg13g2_nor2_1 _3423_ (.A(net691),
    .B(net685),
    .Y(_0980_));
 sg13g2_nor4_2 _3424_ (.A(net692),
    .B(net686),
    .C(net676),
    .Y(_0981_),
    .D(net665));
 sg13g2_nor2_1 _3425_ (.A(_0907_),
    .B(_0981_),
    .Y(_0982_));
 sg13g2_xor2_1 _3426_ (.B(_0982_),
    .A(net659),
    .X(_0983_));
 sg13g2_nand2_1 _3427_ (.Y(_0984_),
    .A(_0047_),
    .B(_0983_));
 sg13g2_or2_1 _3428_ (.X(_0985_),
    .B(_0983_),
    .A(_0047_));
 sg13g2_nand2_1 _3429_ (.Y(_0986_),
    .A(_0984_),
    .B(_0985_));
 sg13g2_nand2b_1 _3430_ (.Y(_0987_),
    .B(_0986_),
    .A_N(_0979_));
 sg13g2_xor2_1 _3431_ (.B(_0986_),
    .A(_0979_),
    .X(_0988_));
 sg13g2_o21ai_1 _3432_ (.B1(net691),
    .Y(_0989_),
    .A1(net685),
    .A2(_0856_));
 sg13g2_o21ai_1 _3433_ (.B1(_0812_),
    .Y(_0990_),
    .A1(_1458_),
    .A2(net669));
 sg13g2_nor2_1 _3434_ (.A(net682),
    .B(_0938_),
    .Y(_0991_));
 sg13g2_a21oi_1 _3435_ (.A1(net682),
    .A2(_0990_),
    .Y(_0992_),
    .B1(_0991_));
 sg13g2_a22oi_1 _3436_ (.Y(_0993_),
    .B1(_0992_),
    .B2(net687),
    .A2(_0934_),
    .A1(_0833_));
 sg13g2_nand2_1 _3437_ (.Y(_0994_),
    .A(_0816_),
    .B(net657));
 sg13g2_nand2_1 _3438_ (.Y(_0995_),
    .A(net684),
    .B(_0861_));
 sg13g2_nand3_1 _3439_ (.B(_0994_),
    .C(_0995_),
    .A(_0820_),
    .Y(_0996_));
 sg13g2_o21ai_1 _3440_ (.B1(_0996_),
    .Y(_0997_),
    .A1(_0839_),
    .A2(_0993_));
 sg13g2_nand2_2 _3441_ (.Y(_0998_),
    .A(_0989_),
    .B(_0997_));
 sg13g2_o21ai_1 _3442_ (.B1(net702),
    .Y(_0999_),
    .A1(_0047_),
    .A2(net658));
 sg13g2_a22oi_1 _3443_ (.Y(_1000_),
    .B1(net699),
    .B2(_0999_),
    .A2(net658),
    .A1(_0047_));
 sg13g2_nor3_1 _3444_ (.A(_1363_),
    .B(net658),
    .C(net701),
    .Y(_1001_));
 sg13g2_nor3_1 _3445_ (.A(net732),
    .B(_1000_),
    .C(_1001_),
    .Y(_1002_));
 sg13g2_a22oi_1 _3446_ (.Y(_1003_),
    .B1(_0998_),
    .B2(_1002_),
    .A2(_0988_),
    .A1(net732));
 sg13g2_nand2_1 _3447_ (.Y(_1004_),
    .A(net776),
    .B(_1003_));
 sg13g2_a21oi_1 _3448_ (.A1(\bitty_inst.data_to_ld[4] ),
    .A2(net777),
    .Y(_1005_),
    .B1(net797));
 sg13g2_a221oi_1 _3449_ (.B2(_1005_),
    .C1(net822),
    .B1(_1004_),
    .A1(net798),
    .Y(_0156_),
    .A2(_1378_));
 sg13g2_a21oi_1 _3450_ (.A1(net659),
    .A2(_0981_),
    .Y(_1006_),
    .B1(_0907_));
 sg13g2_xor2_1 _3451_ (.B(_1006_),
    .A(net661),
    .X(_1007_));
 sg13g2_nor2_1 _3452_ (.A(\bitty_inst.alu_inst.in_a[5] ),
    .B(_1007_),
    .Y(_1008_));
 sg13g2_xnor2_1 _3453_ (.Y(_1009_),
    .A(\bitty_inst.alu_inst.in_a[5] ),
    .B(_1007_));
 sg13g2_nand2_1 _3454_ (.Y(_1010_),
    .A(\bitty_inst.alu_inst.in_a[4] ),
    .B(_0983_));
 sg13g2_nand2_1 _3455_ (.Y(_1011_),
    .A(_0987_),
    .B(_1010_));
 sg13g2_xor2_1 _3456_ (.B(_1011_),
    .A(_1009_),
    .X(_1012_));
 sg13g2_nand2_1 _3457_ (.Y(_1013_),
    .A(net687),
    .B(_0875_));
 sg13g2_nand2_1 _3458_ (.Y(_1014_),
    .A(net690),
    .B(_1013_));
 sg13g2_a221oi_1 _3459_ (.B2(net656),
    .C1(_0821_),
    .B1(_0886_),
    .A1(net683),
    .Y(_1015_),
    .A2(_0880_));
 sg13g2_o21ai_1 _3460_ (.B1(_0888_),
    .Y(_1016_),
    .A1(_1457_),
    .A2(net664));
 sg13g2_mux2_1 _3461_ (.A0(_0972_),
    .A1(_1016_),
    .S(net679),
    .X(_1017_));
 sg13g2_nor2_1 _3462_ (.A(net683),
    .B(_1017_),
    .Y(_1018_));
 sg13g2_a21oi_1 _3463_ (.A1(net683),
    .A2(_0899_),
    .Y(_1019_),
    .B1(_1018_));
 sg13g2_o21ai_1 _3464_ (.B1(net702),
    .Y(_1020_),
    .A1(_0046_),
    .A2(net661));
 sg13g2_a22oi_1 _3465_ (.Y(_1021_),
    .B1(net699),
    .B2(_1020_),
    .A2(net661),
    .A1(_0046_));
 sg13g2_nor3_1 _3466_ (.A(_1362_),
    .B(net660),
    .C(net701),
    .Y(_1022_));
 sg13g2_nor3_1 _3467_ (.A(net778),
    .B(_1021_),
    .C(_1022_),
    .Y(_1023_));
 sg13g2_o21ai_1 _3468_ (.B1(_1023_),
    .Y(_1024_),
    .A1(_0839_),
    .A2(_1019_));
 sg13g2_a21oi_2 _3469_ (.B1(_1024_),
    .Y(_1025_),
    .A2(_1015_),
    .A1(_1014_));
 sg13g2_o21ai_1 _3470_ (.B1(_1025_),
    .Y(_1026_),
    .A1(net730),
    .A2(_1012_));
 sg13g2_a21oi_1 _3471_ (.A1(_1459_),
    .A2(net777),
    .Y(_1027_),
    .B1(net797));
 sg13g2_a22oi_1 _3472_ (.Y(_1028_),
    .B1(_1026_),
    .B2(_1027_),
    .A2(net935),
    .A1(net798));
 sg13g2_nor2_1 _3473_ (.A(net819),
    .B(_1028_),
    .Y(_0157_));
 sg13g2_a22oi_1 _3474_ (.Y(_1029_),
    .B1(_1007_),
    .B2(\bitty_inst.alu_inst.in_a[5] ),
    .A2(_0983_),
    .A1(\bitty_inst.alu_inst.in_a[4] ));
 sg13g2_a221oi_1 _3475_ (.B2(_0985_),
    .C1(_1009_),
    .B1(_0984_),
    .A1(_0954_),
    .Y(_1030_),
    .A2(_0956_));
 sg13g2_a21o_1 _3476_ (.A2(_1029_),
    .A1(_0987_),
    .B1(_1008_),
    .X(_1031_));
 sg13g2_and3_1 _3477_ (.X(_1032_),
    .A(net660),
    .B(net659),
    .C(_0981_));
 sg13g2_o21ai_1 _3478_ (.B1(net694),
    .Y(_1033_),
    .A1(_0907_),
    .A2(_1032_));
 sg13g2_or3_1 _3479_ (.A(net694),
    .B(_0907_),
    .C(_1032_),
    .X(_1034_));
 sg13g2_and2_1 _3480_ (.A(_1033_),
    .B(_1034_),
    .X(_1035_));
 sg13g2_xnor2_1 _3481_ (.Y(_1036_),
    .A(_0045_),
    .B(_1035_));
 sg13g2_xor2_1 _3482_ (.B(_1036_),
    .A(_1031_),
    .X(_1037_));
 sg13g2_nand2_1 _3483_ (.Y(_1038_),
    .A(net684),
    .B(_0933_));
 sg13g2_nand2_1 _3484_ (.Y(_1039_),
    .A(net688),
    .B(_0935_));
 sg13g2_a221oi_1 _3485_ (.B2(net691),
    .C1(_0821_),
    .B1(_1039_),
    .A1(_0928_),
    .Y(_1040_),
    .A2(net657));
 sg13g2_o21ai_1 _3486_ (.B1(_0814_),
    .Y(_1041_),
    .A1(_1457_),
    .A2(net669));
 sg13g2_mux2_1 _3487_ (.A0(_0990_),
    .A1(_1041_),
    .S(net680),
    .X(_1042_));
 sg13g2_nand2_1 _3488_ (.Y(_1043_),
    .A(net684),
    .B(_0939_));
 sg13g2_o21ai_1 _3489_ (.B1(_1043_),
    .Y(_1044_),
    .A1(net684),
    .A2(_1042_));
 sg13g2_o21ai_1 _3490_ (.B1(net702),
    .Y(_1045_),
    .A1(_0045_),
    .A2(net695));
 sg13g2_a22oi_1 _3491_ (.Y(_1046_),
    .B1(net699),
    .B2(_1045_),
    .A2(net694),
    .A1(_0045_));
 sg13g2_nor3_1 _3492_ (.A(_1361_),
    .B(net695),
    .C(net701),
    .Y(_1047_));
 sg13g2_or3_1 _3493_ (.A(net732),
    .B(_1046_),
    .C(_1047_),
    .X(_1048_));
 sg13g2_a221oi_1 _3494_ (.B2(_0838_),
    .C1(_1048_),
    .B1(_1044_),
    .A1(_1038_),
    .Y(_1049_),
    .A2(_1040_));
 sg13g2_nor2_1 _3495_ (.A(net777),
    .B(_1049_),
    .Y(_1050_));
 sg13g2_o21ai_1 _3496_ (.B1(_1050_),
    .Y(_1051_),
    .A1(net730),
    .A2(_1037_));
 sg13g2_a21oi_1 _3497_ (.A1(\bitty_inst.data_to_ld[6] ),
    .A2(net777),
    .Y(_1052_),
    .B1(net797));
 sg13g2_a221oi_1 _3498_ (.B2(_1052_),
    .C1(net819),
    .B1(_1051_),
    .A1(net798),
    .Y(_0158_),
    .A2(_1376_));
 sg13g2_a21oi_1 _3499_ (.A1(_1033_),
    .A2(_1034_),
    .Y(_1053_),
    .B1(_1361_));
 sg13g2_nand2b_1 _3500_ (.Y(_1054_),
    .B(\bitty_inst.alu_inst.in_a[6] ),
    .A_N(_1035_));
 sg13g2_o21ai_1 _3501_ (.B1(_1054_),
    .Y(_1055_),
    .A1(_1031_),
    .A2(_1036_));
 sg13g2_nand4_1 _3502_ (.B(net661),
    .C(net659),
    .A(net694),
    .Y(_1056_),
    .D(_0981_));
 sg13g2_a21oi_1 _3503_ (.A1(net697),
    .A2(_1056_),
    .Y(_1057_),
    .B1(_0703_));
 sg13g2_and3_1 _3504_ (.X(_1058_),
    .A(_0703_),
    .B(net697),
    .C(_1056_));
 sg13g2_nor3_1 _3505_ (.A(_1360_),
    .B(_1057_),
    .C(_1058_),
    .Y(_1059_));
 sg13g2_o21ai_1 _3506_ (.B1(_1360_),
    .Y(_1060_),
    .A1(_1057_),
    .A2(_1058_));
 sg13g2_nand2b_1 _3507_ (.Y(_1061_),
    .B(_1060_),
    .A_N(_1059_));
 sg13g2_xnor2_1 _3508_ (.Y(_1062_),
    .A(_1055_),
    .B(_1061_));
 sg13g2_o21ai_1 _3509_ (.B1(_0882_),
    .Y(_1063_),
    .A1(_1456_),
    .A2(net666));
 sg13g2_mux2_1 _3510_ (.A0(_1016_),
    .A1(_1063_),
    .S(net679),
    .X(_1064_));
 sg13g2_mux2_1 _3511_ (.A0(_0973_),
    .A1(_1064_),
    .S(net689),
    .X(_1065_));
 sg13g2_a21oi_1 _3512_ (.A1(net689),
    .A2(_0964_),
    .Y(_1066_),
    .B1(_0746_));
 sg13g2_a21oi_1 _3513_ (.A1(_0959_),
    .A2(net656),
    .Y(_1067_),
    .B1(_1066_));
 sg13g2_nand2_1 _3514_ (.Y(_1068_),
    .A(_0820_),
    .B(_1067_));
 sg13g2_a21oi_1 _3515_ (.A1(net683),
    .A2(_0965_),
    .Y(_1069_),
    .B1(_1068_));
 sg13g2_o21ai_1 _3516_ (.B1(net702),
    .Y(_1070_),
    .A1(_0044_),
    .A2(_0703_));
 sg13g2_a22oi_1 _3517_ (.Y(_1071_),
    .B1(net699),
    .B2(_1070_),
    .A2(_0703_),
    .A1(_0044_));
 sg13g2_o21ai_1 _3518_ (.B1(net776),
    .Y(_1072_),
    .A1(_0705_),
    .A2(net701));
 sg13g2_nor3_1 _3519_ (.A(_1069_),
    .B(_1071_),
    .C(_1072_),
    .Y(_1073_));
 sg13g2_o21ai_1 _3520_ (.B1(_1073_),
    .Y(_1074_),
    .A1(_0839_),
    .A2(_1065_));
 sg13g2_a21oi_1 _3521_ (.A1(net732),
    .A2(_1062_),
    .Y(_1075_),
    .B1(_1074_));
 sg13g2_o21ai_1 _3522_ (.B1(net808),
    .Y(_1076_),
    .A1(\bitty_inst.data_to_ld[7] ),
    .A2(net776));
 sg13g2_nor2_1 _3523_ (.A(_1075_),
    .B(_1076_),
    .Y(_1077_));
 sg13g2_a21oi_1 _3524_ (.A1(net798),
    .A2(net893),
    .Y(_1078_),
    .B1(_1077_));
 sg13g2_nor2_1 _3525_ (.A(net819),
    .B(_1078_),
    .Y(_0159_));
 sg13g2_a21oi_1 _3526_ (.A1(_1053_),
    .A2(_1060_),
    .Y(_1079_),
    .B1(_1059_));
 sg13g2_o21ai_1 _3527_ (.B1(_1079_),
    .Y(_1080_),
    .A1(_1036_),
    .A2(_1061_));
 sg13g2_o21ai_1 _3528_ (.B1(_1079_),
    .Y(_1081_),
    .A1(_1008_),
    .A2(_1029_));
 sg13g2_o21ai_1 _3529_ (.B1(_1080_),
    .Y(_1082_),
    .A1(_1030_),
    .A2(_1081_));
 sg13g2_and2_1 _3530_ (.A(_0703_),
    .B(net694),
    .X(_1083_));
 sg13g2_nand4_1 _3531_ (.B(net659),
    .C(_0981_),
    .A(net660),
    .Y(_1084_),
    .D(_1083_));
 sg13g2_nand2_1 _3532_ (.Y(_1085_),
    .A(net698),
    .B(_1084_));
 sg13g2_xnor2_1 _3533_ (.Y(_1086_),
    .A(_0688_),
    .B(_1085_));
 sg13g2_xor2_1 _3534_ (.B(_1086_),
    .A(_0043_),
    .X(_1087_));
 sg13g2_nor2_1 _3535_ (.A(_1082_),
    .B(_1087_),
    .Y(_1088_));
 sg13g2_and2_1 _3536_ (.A(_1082_),
    .B(_1087_),
    .X(_1089_));
 sg13g2_o21ai_1 _3537_ (.B1(net733),
    .Y(_1090_),
    .A1(_1088_),
    .A2(_1089_));
 sg13g2_nand2_1 _3538_ (.Y(_1091_),
    .A(net693),
    .B(_0992_));
 sg13g2_nor2_1 _3539_ (.A(_0834_),
    .B(net657),
    .Y(_1092_));
 sg13g2_o21ai_1 _3540_ (.B1(_0857_),
    .Y(_1093_),
    .A1(_1456_),
    .A2(net671));
 sg13g2_mux2_1 _3541_ (.A0(_1041_),
    .A1(_1093_),
    .S(net680),
    .X(_1094_));
 sg13g2_a221oi_1 _3542_ (.B2(net657),
    .C1(_0837_),
    .B1(_1094_),
    .A1(_1091_),
    .Y(_1095_),
    .A2(_1092_));
 sg13g2_o21ai_1 _3543_ (.B1(net703),
    .Y(_1096_),
    .A1(_0043_),
    .A2(_0688_));
 sg13g2_a22oi_1 _3544_ (.Y(_1097_),
    .B1(net700),
    .B2(_1096_),
    .A2(_0688_),
    .A1(_0043_));
 sg13g2_and3_1 _3545_ (.X(_1098_),
    .A(\bitty_inst.alu_inst.in_a[8] ),
    .B(_0689_),
    .C(_0845_));
 sg13g2_nor4_1 _3546_ (.A(net733),
    .B(_1095_),
    .C(_1097_),
    .D(_1098_),
    .Y(_1099_));
 sg13g2_o21ai_1 _3547_ (.B1(_1099_),
    .Y(_1100_),
    .A1(_0823_),
    .A2(_0862_));
 sg13g2_nand3_1 _3548_ (.B(_1090_),
    .C(_1100_),
    .A(net776),
    .Y(_1101_));
 sg13g2_a21oi_1 _3549_ (.A1(\bitty_inst.data_to_ld[8] ),
    .A2(net779),
    .Y(_1102_),
    .B1(net800));
 sg13g2_a221oi_1 _3550_ (.B2(_1102_),
    .C1(net821),
    .B1(_1101_),
    .A1(net799),
    .Y(_0160_),
    .A2(_1374_));
 sg13g2_a21oi_1 _3551_ (.A1(\bitty_inst.alu_inst.in_a[8] ),
    .A2(_1086_),
    .Y(_1103_),
    .B1(_1088_));
 sg13g2_o21ai_1 _3552_ (.B1(net698),
    .Y(_1104_),
    .A1(_0689_),
    .A2(_1084_));
 sg13g2_xnor2_1 _3553_ (.Y(_1105_),
    .A(net662),
    .B(_1104_));
 sg13g2_nor2_1 _3554_ (.A(\bitty_inst.alu_inst.in_a[9] ),
    .B(_1105_),
    .Y(_1106_));
 sg13g2_xnor2_1 _3555_ (.Y(_1107_),
    .A(\bitty_inst.alu_inst.in_a[9] ),
    .B(_1105_));
 sg13g2_a21oi_1 _3556_ (.A1(_1103_),
    .A2(_1107_),
    .Y(_1108_),
    .B1(net731));
 sg13g2_o21ai_1 _3557_ (.B1(_1108_),
    .Y(_1109_),
    .A1(_1103_),
    .A2(_1107_));
 sg13g2_nor2_2 _3558_ (.A(net690),
    .B(_0761_),
    .Y(_1110_));
 sg13g2_a21oi_1 _3559_ (.A1(_1455_),
    .A2(net669),
    .Y(_1111_),
    .B1(_0884_));
 sg13g2_mux2_1 _3560_ (.A0(_1063_),
    .A1(_1111_),
    .S(net679),
    .X(_1112_));
 sg13g2_a22oi_1 _3561_ (.Y(_1113_),
    .B1(_1112_),
    .B2(net656),
    .A2(_1110_),
    .A1(_1017_));
 sg13g2_a22oi_1 _3562_ (.Y(_1114_),
    .B1(_1113_),
    .B2(_0836_),
    .A2(_0881_),
    .A1(_0822_));
 sg13g2_a21oi_2 _3563_ (.B1(_1114_),
    .Y(_1115_),
    .A2(_0900_),
    .A1(net690));
 sg13g2_o21ai_1 _3564_ (.B1(net703),
    .Y(_1116_),
    .A1(_0042_),
    .A2(net662));
 sg13g2_a22oi_1 _3565_ (.Y(_1117_),
    .B1(net700),
    .B2(_1116_),
    .A2(net662),
    .A1(_0042_));
 sg13g2_nor3_1 _3566_ (.A(_1359_),
    .B(net662),
    .C(_0844_),
    .Y(_1118_));
 sg13g2_nor4_1 _3567_ (.A(net779),
    .B(_1115_),
    .C(_1117_),
    .D(_1118_),
    .Y(_1119_));
 sg13g2_o21ai_1 _3568_ (.B1(net809),
    .Y(_1120_),
    .A1(\bitty_inst.data_to_ld[9] ),
    .A2(_0867_));
 sg13g2_a21oi_2 _3569_ (.B1(_1120_),
    .Y(_1121_),
    .A2(_1119_),
    .A1(_1109_));
 sg13g2_a21oi_1 _3570_ (.A1(net799),
    .A2(net941),
    .Y(_1122_),
    .B1(_1121_));
 sg13g2_nor2_1 _3571_ (.A(net821),
    .B(_1122_),
    .Y(_0161_));
 sg13g2_a22oi_1 _3572_ (.Y(_1123_),
    .B1(_1105_),
    .B2(\bitty_inst.alu_inst.in_a[9] ),
    .A2(_1086_),
    .A1(\bitty_inst.alu_inst.in_a[8] ));
 sg13g2_or2_1 _3573_ (.X(_1124_),
    .B(_1123_),
    .A(_1106_));
 sg13g2_or2_1 _3574_ (.X(_1125_),
    .B(_1107_),
    .A(_1087_));
 sg13g2_o21ai_1 _3575_ (.B1(_1124_),
    .Y(_1126_),
    .A1(_1082_),
    .A2(_1125_));
 sg13g2_nand2b_1 _3576_ (.Y(_1127_),
    .B(net698),
    .A_N(_0681_));
 sg13g2_nand2_1 _3577_ (.Y(_1128_),
    .A(_1104_),
    .B(_1127_));
 sg13g2_xor2_1 _3578_ (.B(_1128_),
    .A(_0672_),
    .X(_1129_));
 sg13g2_xor2_1 _3579_ (.B(_1129_),
    .A(net806),
    .X(_1130_));
 sg13g2_inv_1 _3580_ (.Y(_1131_),
    .A(_1130_));
 sg13g2_xnor2_1 _3581_ (.Y(_1132_),
    .A(_1126_),
    .B(_1130_));
 sg13g2_o21ai_1 _3582_ (.B1(_0859_),
    .Y(_1133_),
    .A1(_1455_),
    .A2(net671));
 sg13g2_mux2_1 _3583_ (.A0(_1093_),
    .A1(_1133_),
    .S(net680),
    .X(_1134_));
 sg13g2_a221oi_1 _3584_ (.B2(net657),
    .C1(_0837_),
    .B1(_1134_),
    .A1(net684),
    .Y(_1135_),
    .A2(_1042_));
 sg13g2_a21oi_1 _3585_ (.A1(_0822_),
    .A2(_0937_),
    .Y(_1136_),
    .B1(_1135_));
 sg13g2_a21oi_1 _3586_ (.A1(net691),
    .A2(_0940_),
    .Y(_1137_),
    .B1(_1136_));
 sg13g2_o21ai_1 _3587_ (.B1(net703),
    .Y(_1138_),
    .A1(net806),
    .A2(net663));
 sg13g2_a22oi_1 _3588_ (.Y(_1139_),
    .B1(net700),
    .B2(_1138_),
    .A2(net663),
    .A1(net806));
 sg13g2_nor3_1 _3589_ (.A(_1358_),
    .B(net663),
    .C(_0844_),
    .Y(_1140_));
 sg13g2_nor3_1 _3590_ (.A(_1137_),
    .B(_1139_),
    .C(_1140_),
    .Y(_1141_));
 sg13g2_a21oi_1 _3591_ (.A1(net731),
    .A2(_1141_),
    .Y(_1142_),
    .B1(net779));
 sg13g2_o21ai_1 _3592_ (.B1(_1142_),
    .Y(_1143_),
    .A1(net731),
    .A2(_1132_));
 sg13g2_a21oi_2 _3593_ (.B1(net800),
    .Y(_1144_),
    .A2(net779),
    .A1(\bitty_inst.data_to_ld[10] ));
 sg13g2_a221oi_1 _3594_ (.B2(_1144_),
    .C1(net821),
    .B1(_1143_),
    .A1(net799),
    .Y(_0162_),
    .A2(_1372_));
 sg13g2_nand2_1 _3595_ (.Y(_1145_),
    .A(net799),
    .B(net954));
 sg13g2_nand2_1 _3596_ (.Y(_1146_),
    .A(\bitty_inst.alu_inst.in_a[10] ),
    .B(_1129_));
 sg13g2_a22oi_1 _3597_ (.Y(_1147_),
    .B1(_1131_),
    .B2(_1126_),
    .A2(_1129_),
    .A1(\bitty_inst.alu_inst.in_a[10] ));
 sg13g2_nand2b_1 _3598_ (.Y(_1148_),
    .B(net698),
    .A_N(net663));
 sg13g2_nand3_1 _3599_ (.B(_1127_),
    .C(_1148_),
    .A(_1104_),
    .Y(_1149_));
 sg13g2_xnor2_1 _3600_ (.Y(_1150_),
    .A(_0665_),
    .B(_1149_));
 sg13g2_xnor2_1 _3601_ (.Y(_1151_),
    .A(\bitty_inst.alu_inst.in_a[11] ),
    .B(_1150_));
 sg13g2_o21ai_1 _3602_ (.B1(net733),
    .Y(_1152_),
    .A1(_1147_),
    .A2(_1151_));
 sg13g2_a21oi_1 _3603_ (.A1(_1147_),
    .A2(_1151_),
    .Y(_1153_),
    .B1(_1152_));
 sg13g2_mux2_1 _3604_ (.A0(net805),
    .A1(net806),
    .S(net664),
    .X(_1154_));
 sg13g2_mux2_1 _3605_ (.A0(_1111_),
    .A1(_1154_),
    .S(net680),
    .X(_1155_));
 sg13g2_a22oi_1 _3606_ (.Y(_1156_),
    .B1(_1155_),
    .B2(net656),
    .A2(_1064_),
    .A1(net685));
 sg13g2_o21ai_1 _3607_ (.B1(_1156_),
    .Y(_1157_),
    .A1(net693),
    .A2(_0974_));
 sg13g2_o21ai_1 _3608_ (.B1(net703),
    .Y(_1158_),
    .A1(net805),
    .A2(_0664_));
 sg13g2_a22oi_1 _3609_ (.Y(_1159_),
    .B1(net700),
    .B2(_1158_),
    .A2(_0664_),
    .A1(net805));
 sg13g2_a221oi_1 _3610_ (.B2(_0822_),
    .C1(_1159_),
    .B1(_0967_),
    .A1(_0666_),
    .Y(_1160_),
    .A2(_0845_));
 sg13g2_o21ai_1 _3611_ (.B1(_1160_),
    .Y(_1161_),
    .A1(_0837_),
    .A2(_1157_));
 sg13g2_nor3_1 _3612_ (.A(net779),
    .B(_1153_),
    .C(_1161_),
    .Y(_1162_));
 sg13g2_o21ai_1 _3613_ (.B1(net809),
    .Y(_1163_),
    .A1(\bitty_inst.data_to_ld[11] ),
    .A2(net776));
 sg13g2_o21ai_1 _3614_ (.B1(_1145_),
    .Y(_1164_),
    .A1(_1162_),
    .A2(_1163_));
 sg13g2_and2_1 _3615_ (.A(net854),
    .B(_1164_),
    .X(_0163_));
 sg13g2_or4_1 _3616_ (.A(_1082_),
    .B(_1125_),
    .C(_1130_),
    .D(_1151_),
    .X(_1165_));
 sg13g2_nor3_1 _3617_ (.A(_1124_),
    .B(_1130_),
    .C(_1151_),
    .Y(_1166_));
 sg13g2_nand2b_1 _3618_ (.Y(_1167_),
    .B(_1150_),
    .A_N(net805));
 sg13g2_o21ai_1 _3619_ (.B1(_1167_),
    .Y(_1168_),
    .A1(_1146_),
    .A2(_1151_));
 sg13g2_nor2_1 _3620_ (.A(_1166_),
    .B(_1168_),
    .Y(_1169_));
 sg13g2_nand2_1 _3621_ (.Y(_1170_),
    .A(_0665_),
    .B(net697));
 sg13g2_nand4_1 _3622_ (.B(_1127_),
    .C(_1148_),
    .A(_1104_),
    .Y(_1171_),
    .D(_1170_));
 sg13g2_xnor2_1 _3623_ (.Y(_1172_),
    .A(_0651_),
    .B(_1171_));
 sg13g2_xor2_1 _3624_ (.B(_1172_),
    .A(net804),
    .X(_1173_));
 sg13g2_a21oi_1 _3625_ (.A1(_1165_),
    .A2(_1169_),
    .Y(_1174_),
    .B1(_1173_));
 sg13g2_and3_1 _3626_ (.X(_1175_),
    .A(_1165_),
    .B(_1169_),
    .C(_1173_));
 sg13g2_o21ai_1 _3627_ (.B1(net733),
    .Y(_1176_),
    .A1(_1174_),
    .A2(_1175_));
 sg13g2_nor2_1 _3628_ (.A(net680),
    .B(_1133_),
    .Y(_1177_));
 sg13g2_mux2_1 _3629_ (.A0(net804),
    .A1(net805),
    .S(net666),
    .X(_1178_));
 sg13g2_o21ai_1 _3630_ (.B1(net656),
    .Y(_1179_),
    .A1(net674),
    .A2(_1178_));
 sg13g2_a21oi_1 _3631_ (.A1(_1094_),
    .A2(_1110_),
    .Y(_1180_),
    .B1(_0837_));
 sg13g2_o21ai_1 _3632_ (.B1(_1180_),
    .Y(_1181_),
    .A1(_1177_),
    .A2(_1179_));
 sg13g2_a21oi_1 _3633_ (.A1(net690),
    .A2(_0993_),
    .Y(_1182_),
    .B1(_1181_));
 sg13g2_nor3_1 _3634_ (.A(net684),
    .B(_0823_),
    .C(_0856_),
    .Y(_1183_));
 sg13g2_o21ai_1 _3635_ (.B1(net703),
    .Y(_1184_),
    .A1(net804),
    .A2(_0650_));
 sg13g2_a22oi_1 _3636_ (.Y(_1185_),
    .B1(net700),
    .B2(_1184_),
    .A2(_0650_),
    .A1(net804));
 sg13g2_and3_1 _3637_ (.X(_1186_),
    .A(\bitty_inst.alu_inst.in_a[12] ),
    .B(_0651_),
    .C(_0845_));
 sg13g2_nor4_1 _3638_ (.A(_1182_),
    .B(_1183_),
    .C(_1185_),
    .D(_1186_),
    .Y(_1187_));
 sg13g2_a21oi_1 _3639_ (.A1(net731),
    .A2(_1187_),
    .Y(_1188_),
    .B1(net779));
 sg13g2_a221oi_1 _3640_ (.B2(_1188_),
    .C1(net799),
    .B1(_1176_),
    .A1(\bitty_inst.data_to_ld[12] ),
    .Y(_1189_),
    .A2(net779));
 sg13g2_o21ai_1 _3641_ (.B1(net854),
    .Y(_1190_),
    .A1(net809),
    .A2(net951));
 sg13g2_nor2_1 _3642_ (.A(_1189_),
    .B(_1190_),
    .Y(_0164_));
 sg13g2_nand2_1 _3643_ (.Y(_1191_),
    .A(net799),
    .B(net902));
 sg13g2_nand2_1 _3644_ (.Y(_1192_),
    .A(\bitty_inst.alu_inst.in_a[12] ),
    .B(_1172_));
 sg13g2_nor2b_1 _3645_ (.A(_1174_),
    .B_N(_1192_),
    .Y(_1193_));
 sg13g2_o21ai_1 _3646_ (.B1(net697),
    .Y(_1194_),
    .A1(_0651_),
    .A2(_1171_));
 sg13g2_xnor2_1 _3647_ (.Y(_1195_),
    .A(_0644_),
    .B(_1194_));
 sg13g2_xnor2_1 _3648_ (.Y(_1196_),
    .A(net803),
    .B(_1195_));
 sg13g2_a21oi_1 _3649_ (.A1(_1193_),
    .A2(_1196_),
    .Y(_1197_),
    .B1(net730));
 sg13g2_o21ai_1 _3650_ (.B1(_1197_),
    .Y(_1198_),
    .A1(_1193_),
    .A2(_1196_));
 sg13g2_mux2_1 _3651_ (.A0(net803),
    .A1(net804),
    .S(net664),
    .X(_1199_));
 sg13g2_nor2_1 _3652_ (.A(net680),
    .B(_1154_),
    .Y(_1200_));
 sg13g2_o21ai_1 _3653_ (.B1(net656),
    .Y(_1201_),
    .A1(net675),
    .A2(_1199_));
 sg13g2_o21ai_1 _3654_ (.B1(_0836_),
    .Y(_1202_),
    .A1(_1200_),
    .A2(_1201_));
 sg13g2_a221oi_1 _3655_ (.B2(_1112_),
    .C1(_1202_),
    .B1(_1110_),
    .A1(net690),
    .Y(_1203_),
    .A2(_1019_));
 sg13g2_o21ai_1 _3656_ (.B1(net703),
    .Y(_1204_),
    .A1(net803),
    .A2(_0643_));
 sg13g2_a22oi_1 _3657_ (.Y(_1205_),
    .B1(net700),
    .B2(_1204_),
    .A2(_0643_),
    .A1(net803));
 sg13g2_nand3_1 _3658_ (.B(_0644_),
    .C(_0845_),
    .A(\bitty_inst.alu_inst.in_a[13] ),
    .Y(_1206_));
 sg13g2_o21ai_1 _3659_ (.B1(_1206_),
    .Y(_1207_),
    .A1(_0823_),
    .A2(_1013_));
 sg13g2_nor4_1 _3660_ (.A(net779),
    .B(_1203_),
    .C(_1205_),
    .D(_1207_),
    .Y(_1208_));
 sg13g2_o21ai_1 _3661_ (.B1(net809),
    .Y(_1209_),
    .A1(\bitty_inst.data_to_ld[13] ),
    .A2(net776));
 sg13g2_a21o_1 _3662_ (.A2(_1208_),
    .A1(_1198_),
    .B1(_1209_),
    .X(_1210_));
 sg13g2_a21oi_1 _3663_ (.A1(_1191_),
    .A2(_1210_),
    .Y(_0165_),
    .B1(net821));
 sg13g2_or2_1 _3664_ (.X(_1211_),
    .B(_1196_),
    .A(_1173_));
 sg13g2_a21oi_2 _3665_ (.B1(_1211_),
    .Y(_1212_),
    .A2(_1169_),
    .A1(_1165_));
 sg13g2_nand2b_1 _3666_ (.Y(_1213_),
    .B(\bitty_inst.alu_inst.in_a[13] ),
    .A_N(_1195_));
 sg13g2_o21ai_1 _3667_ (.B1(_1213_),
    .Y(_1214_),
    .A1(_1192_),
    .A2(_1196_));
 sg13g2_nor2_1 _3668_ (.A(_1212_),
    .B(_1214_),
    .Y(_1215_));
 sg13g2_a21oi_2 _3669_ (.B1(_0907_),
    .Y(_1216_),
    .A2(_1194_),
    .A1(_0643_));
 sg13g2_xnor2_1 _3670_ (.Y(_1217_),
    .A(_0635_),
    .B(_1216_));
 sg13g2_xor2_1 _3671_ (.B(_1217_),
    .A(net802),
    .X(_1218_));
 sg13g2_o21ai_1 _3672_ (.B1(_1218_),
    .Y(_1219_),
    .A1(_1212_),
    .A2(_1214_));
 sg13g2_xnor2_1 _3673_ (.Y(_1220_),
    .A(_1215_),
    .B(_1218_));
 sg13g2_a21oi_1 _3674_ (.A1(_1110_),
    .A2(_1134_),
    .Y(_1221_),
    .B1(_0837_));
 sg13g2_a21oi_1 _3675_ (.A1(net803),
    .A2(net666),
    .Y(_1222_),
    .B1(net674));
 sg13g2_o21ai_1 _3676_ (.B1(net656),
    .Y(_1223_),
    .A1(net680),
    .A2(_1178_));
 sg13g2_a21oi_1 _3677_ (.A1(_0854_),
    .A2(_1222_),
    .Y(_1224_),
    .B1(_1223_));
 sg13g2_nor2b_1 _3678_ (.A(_1224_),
    .B_N(_1221_),
    .Y(_1225_));
 sg13g2_o21ai_1 _3679_ (.B1(_1225_),
    .Y(_1226_),
    .A1(net693),
    .A2(_1044_));
 sg13g2_nor2_1 _3680_ (.A(_0823_),
    .B(_1039_),
    .Y(_1227_));
 sg13g2_o21ai_1 _3681_ (.B1(net703),
    .Y(_1228_),
    .A1(net802),
    .A2(_0635_));
 sg13g2_a22oi_1 _3682_ (.Y(_1229_),
    .B1(net700),
    .B2(_1228_),
    .A2(_0635_),
    .A1(net802));
 sg13g2_and3_1 _3683_ (.X(_1230_),
    .A(\bitty_inst.alu_inst.in_a[14] ),
    .B(_0636_),
    .C(_0845_));
 sg13g2_nor4_1 _3684_ (.A(net733),
    .B(_1227_),
    .C(_1229_),
    .D(_1230_),
    .Y(_1231_));
 sg13g2_a21oi_1 _3685_ (.A1(_1226_),
    .A2(_1231_),
    .Y(_1232_),
    .B1(net780));
 sg13g2_o21ai_1 _3686_ (.B1(_1232_),
    .Y(_1233_),
    .A1(net731),
    .A2(_1220_));
 sg13g2_a21oi_1 _3687_ (.A1(\bitty_inst.data_to_ld[14] ),
    .A2(net780),
    .Y(_1234_),
    .B1(net799));
 sg13g2_a221oi_1 _3688_ (.B2(_1234_),
    .C1(net821),
    .B1(_1233_),
    .A1(net799),
    .Y(_0166_),
    .A2(_1368_));
 sg13g2_nand2_1 _3689_ (.Y(_1235_),
    .A(net897),
    .B(net800));
 sg13g2_nand2b_1 _3690_ (.Y(_1236_),
    .B(\bitty_inst.alu_inst.in_a[14] ),
    .A_N(_1217_));
 sg13g2_o21ai_1 _3691_ (.B1(net697),
    .Y(_1237_),
    .A1(_0636_),
    .A2(_1216_));
 sg13g2_xnor2_1 _3692_ (.Y(_1238_),
    .A(\bitty_inst.alu_inst.in_a[15] ),
    .B(_0628_));
 sg13g2_xnor2_1 _3693_ (.Y(_1239_),
    .A(_1237_),
    .B(_1238_));
 sg13g2_nand3_1 _3694_ (.B(_1236_),
    .C(_1239_),
    .A(_1219_),
    .Y(_1240_));
 sg13g2_a21o_1 _3695_ (.A2(_1236_),
    .A1(_1219_),
    .B1(_1239_),
    .X(_1241_));
 sg13g2_nand3_1 _3696_ (.B(_1240_),
    .C(_1241_),
    .A(net733),
    .Y(_1242_));
 sg13g2_a21oi_1 _3697_ (.A1(_1110_),
    .A2(_1155_),
    .Y(_1243_),
    .B1(_0837_));
 sg13g2_nor3_1 _3698_ (.A(net802),
    .B(net675),
    .C(net670),
    .Y(_1244_));
 sg13g2_o21ai_1 _3699_ (.B1(net656),
    .Y(_1245_),
    .A1(net679),
    .A2(_1199_));
 sg13g2_nor3_1 _3700_ (.A(_0964_),
    .B(_1244_),
    .C(_1245_),
    .Y(_1246_));
 sg13g2_a21oi_1 _3701_ (.A1(net690),
    .A2(_1065_),
    .Y(_1247_),
    .B1(_1246_));
 sg13g2_o21ai_1 _3702_ (.B1(net702),
    .Y(_1248_),
    .A1(_0036_),
    .A2(_0628_));
 sg13g2_a22oi_1 _3703_ (.Y(_1249_),
    .B1(net699),
    .B2(_1248_),
    .A2(_0628_),
    .A1(_0036_));
 sg13g2_nor3_1 _3704_ (.A(_0036_),
    .B(_0823_),
    .C(_0832_),
    .Y(_1250_));
 sg13g2_nor3_1 _3705_ (.A(_1357_),
    .B(_0628_),
    .C(net701),
    .Y(_1251_));
 sg13g2_or4_1 _3706_ (.A(net780),
    .B(_1249_),
    .C(_1250_),
    .D(_1251_),
    .X(_1252_));
 sg13g2_a21oi_1 _3707_ (.A1(_1243_),
    .A2(_1247_),
    .Y(_1253_),
    .B1(_1252_));
 sg13g2_o21ai_1 _3708_ (.B1(net809),
    .Y(_1254_),
    .A1(\bitty_inst.data_to_ld[15] ),
    .A2(net776));
 sg13g2_a21o_1 _3709_ (.A2(_1253_),
    .A1(_1242_),
    .B1(_1254_),
    .X(_1255_));
 sg13g2_a21oi_1 _3710_ (.A1(_1235_),
    .A2(_1255_),
    .Y(_0167_),
    .B1(net821));
 sg13g2_o21ai_1 _3711_ (.B1(net846),
    .Y(_1256_),
    .A1(net909),
    .A2(net786));
 sg13g2_a21oi_1 _3712_ (.A1(net786),
    .A2(net667),
    .Y(_0168_),
    .B1(_1256_));
 sg13g2_o21ai_1 _3713_ (.B1(net832),
    .Y(_1257_),
    .A1(net866),
    .A2(net782));
 sg13g2_a21oi_1 _3714_ (.A1(net782),
    .A2(net677),
    .Y(_0169_),
    .B1(_1257_));
 sg13g2_o21ai_1 _3715_ (.B1(net846),
    .Y(_1258_),
    .A1(net923),
    .A2(net786));
 sg13g2_a21oi_1 _3716_ (.A1(net786),
    .A2(net688),
    .Y(_0170_),
    .B1(_1258_));
 sg13g2_o21ai_1 _3717_ (.B1(net846),
    .Y(_1259_),
    .A1(net591),
    .A2(net782));
 sg13g2_a21oi_1 _3718_ (.A1(net782),
    .A2(net693),
    .Y(_0171_),
    .B1(_1259_));
 sg13g2_o21ai_1 _3719_ (.B1(net843),
    .Y(_1260_),
    .A1(net900),
    .A2(net783));
 sg13g2_a21oi_1 _3720_ (.A1(net783),
    .A2(net658),
    .Y(_0172_),
    .B1(_1260_));
 sg13g2_o21ai_1 _3721_ (.B1(net843),
    .Y(_1261_),
    .A1(net915),
    .A2(net782));
 sg13g2_a21oi_1 _3722_ (.A1(net782),
    .A2(net660),
    .Y(_0173_),
    .B1(_1261_));
 sg13g2_o21ai_1 _3723_ (.B1(net853),
    .Y(_1262_),
    .A1(net885),
    .A2(net786));
 sg13g2_a21oi_1 _3724_ (.A1(net786),
    .A2(net694),
    .Y(_0174_),
    .B1(_1262_));
 sg13g2_o21ai_1 _3725_ (.B1(net853),
    .Y(_1263_),
    .A1(net901),
    .A2(net782));
 sg13g2_a21oi_1 _3726_ (.A1(net782),
    .A2(_0703_),
    .Y(_0175_),
    .B1(_1263_));
 sg13g2_o21ai_1 _3727_ (.B1(net848),
    .Y(_1264_),
    .A1(net872),
    .A2(net784));
 sg13g2_a21oi_1 _3728_ (.A1(net784),
    .A2(_0688_),
    .Y(_0176_),
    .B1(_1264_));
 sg13g2_o21ai_1 _3729_ (.B1(net847),
    .Y(_1265_),
    .A1(net905),
    .A2(net784));
 sg13g2_a21oi_1 _3730_ (.A1(net784),
    .A2(net662),
    .Y(_0177_),
    .B1(_1265_));
 sg13g2_o21ai_1 _3731_ (.B1(net847),
    .Y(_1266_),
    .A1(net865),
    .A2(net784));
 sg13g2_a21oi_1 _3732_ (.A1(net784),
    .A2(net663),
    .Y(_0178_),
    .B1(_1266_));
 sg13g2_o21ai_1 _3733_ (.B1(net847),
    .Y(_1267_),
    .A1(net642),
    .A2(net784));
 sg13g2_a21oi_1 _3734_ (.A1(net784),
    .A2(_0664_),
    .Y(_0179_),
    .B1(_1267_));
 sg13g2_o21ai_1 _3735_ (.B1(net856),
    .Y(_1268_),
    .A1(net879),
    .A2(net785));
 sg13g2_a21oi_1 _3736_ (.A1(net785),
    .A2(_0650_),
    .Y(_0180_),
    .B1(_1268_));
 sg13g2_o21ai_1 _3737_ (.B1(net856),
    .Y(_1269_),
    .A1(net867),
    .A2(net785));
 sg13g2_a21oi_1 _3738_ (.A1(net785),
    .A2(_0643_),
    .Y(_0181_),
    .B1(_1269_));
 sg13g2_o21ai_1 _3739_ (.B1(net853),
    .Y(_1270_),
    .A1(net605),
    .A2(net785));
 sg13g2_a21oi_1 _3740_ (.A1(net785),
    .A2(_0635_),
    .Y(_0182_),
    .B1(_1270_));
 sg13g2_o21ai_1 _3741_ (.B1(net853),
    .Y(_1271_),
    .A1(net892),
    .A2(net786));
 sg13g2_a21oi_1 _3742_ (.A1(net786),
    .A2(_0628_),
    .Y(_0183_),
    .B1(_1271_));
 sg13g2_nor2_2 _3743_ (.A(\bitty_inst.cpu_inst.cur_state[1] ),
    .B(\bitty_inst.cpu_inst.cur_state[0] ),
    .Y(_1272_));
 sg13g2_nand2_1 _3744_ (.Y(_1273_),
    .A(_1442_),
    .B(_1451_));
 sg13g2_o21ai_1 _3745_ (.B1(net828),
    .Y(_1274_),
    .A1(\bitty_inst.d_instr[0] ),
    .A2(net791));
 sg13g2_a21oi_1 _3746_ (.A1(_1356_),
    .A2(net790),
    .Y(_0184_),
    .B1(_1274_));
 sg13g2_o21ai_1 _3747_ (.B1(net829),
    .Y(_1275_),
    .A1(\bitty_inst.d_instr[1] ),
    .A2(net790));
 sg13g2_a21oi_1 _3748_ (.A1(_1355_),
    .A2(net790),
    .Y(_0185_),
    .B1(_1275_));
 sg13g2_o21ai_1 _3749_ (.B1(net831),
    .Y(_1276_),
    .A1(\bitty_inst.d_instr[2] ),
    .A2(net792));
 sg13g2_a21oi_1 _3750_ (.A1(_1354_),
    .A2(net792),
    .Y(_0186_),
    .B1(_1276_));
 sg13g2_o21ai_1 _3751_ (.B1(net831),
    .Y(_1277_),
    .A1(net562),
    .A2(net775));
 sg13g2_a21oi_1 _3752_ (.A1(_1353_),
    .A2(net775),
    .Y(_0187_),
    .B1(_1277_));
 sg13g2_o21ai_1 _3753_ (.B1(net831),
    .Y(_1278_),
    .A1(\bitty_inst.d_instr[4] ),
    .A2(net792));
 sg13g2_a21oi_1 _3754_ (.A1(_1352_),
    .A2(net792),
    .Y(_0188_),
    .B1(_1278_));
 sg13g2_o21ai_1 _3755_ (.B1(net829),
    .Y(_1279_),
    .A1(net622),
    .A2(_1273_));
 sg13g2_a21oi_1 _3756_ (.A1(_1351_),
    .A2(net775),
    .Y(_0189_),
    .B1(_1279_));
 sg13g2_o21ai_1 _3757_ (.B1(net828),
    .Y(_1280_),
    .A1(\bitty_inst.d_instr[6] ),
    .A2(net790));
 sg13g2_a21oi_1 _3758_ (.A1(_1350_),
    .A2(net790),
    .Y(_0190_),
    .B1(_1280_));
 sg13g2_o21ai_1 _3759_ (.B1(net829),
    .Y(_1281_),
    .A1(net630),
    .A2(net775));
 sg13g2_a21oi_1 _3760_ (.A1(_1349_),
    .A2(net775),
    .Y(_0191_),
    .B1(_1281_));
 sg13g2_o21ai_1 _3761_ (.B1(net831),
    .Y(_1282_),
    .A1(\bitty_inst.d_instr[8] ),
    .A2(net792));
 sg13g2_a21oi_1 _3762_ (.A1(_1348_),
    .A2(_1272_),
    .Y(_0192_),
    .B1(_1282_));
 sg13g2_o21ai_1 _3763_ (.B1(net832),
    .Y(_1283_),
    .A1(net641),
    .A2(_1273_));
 sg13g2_a21oi_1 _3764_ (.A1(_1347_),
    .A2(net775),
    .Y(_0193_),
    .B1(_1283_));
 sg13g2_o21ai_1 _3765_ (.B1(net832),
    .Y(_1284_),
    .A1(\bitty_inst.d_instr[10] ),
    .A2(_1272_));
 sg13g2_a21oi_1 _3766_ (.A1(_1346_),
    .A2(_1272_),
    .Y(_0194_),
    .B1(_1284_));
 sg13g2_o21ai_1 _3767_ (.B1(net829),
    .Y(_1285_),
    .A1(net458),
    .A2(net775));
 sg13g2_a21oi_1 _3768_ (.A1(_1345_),
    .A2(net775),
    .Y(_0195_),
    .B1(_1285_));
 sg13g2_o21ai_1 _3769_ (.B1(net828),
    .Y(_1286_),
    .A1(\bitty_inst.d_instr[12] ),
    .A2(net792));
 sg13g2_a21oi_1 _3770_ (.A1(_1344_),
    .A2(net792),
    .Y(_0196_),
    .B1(_1286_));
 sg13g2_o21ai_1 _3771_ (.B1(net829),
    .Y(_1287_),
    .A1(\bitty_inst.d_instr[13] ),
    .A2(net790));
 sg13g2_a21oi_1 _3772_ (.A1(_1343_),
    .A2(net791),
    .Y(_0197_),
    .B1(_1287_));
 sg13g2_o21ai_1 _3773_ (.B1(net829),
    .Y(_1288_),
    .A1(\bitty_inst.d_instr[14] ),
    .A2(net790));
 sg13g2_a21oi_1 _3774_ (.A1(_1342_),
    .A2(net791),
    .Y(_0198_),
    .B1(_1288_));
 sg13g2_o21ai_1 _3775_ (.B1(net829),
    .Y(_1289_),
    .A1(\bitty_inst.d_instr[15] ),
    .A2(net790));
 sg13g2_a21oi_1 _3776_ (.A1(_1341_),
    .A2(net791),
    .Y(_0199_),
    .B1(_1289_));
 sg13g2_nor2_1 _3777_ (.A(net804),
    .B(_1520_),
    .Y(_1290_));
 sg13g2_a21oi_1 _3778_ (.A1(\bitty_inst.alu_inst.in_a[4] ),
    .A2(_1522_),
    .Y(_1291_),
    .B1(_1290_));
 sg13g2_o21ai_1 _3779_ (.B1(_1291_),
    .Y(_1292_),
    .A1(net729),
    .A2(net658));
 sg13g2_nand2_1 _3780_ (.Y(_1293_),
    .A(net811),
    .B(_1292_));
 sg13g2_nor2b_2 _3781_ (.A(net810),
    .B_N(\fi_inst.state[2] ),
    .Y(_1294_));
 sg13g2_a21oi_1 _3782_ (.A1(\addr[4] ),
    .A2(_1294_),
    .Y(_1295_),
    .B1(net815));
 sg13g2_nor2_1 _3783_ (.A(net803),
    .B(_1520_),
    .Y(_1296_));
 sg13g2_a21oi_1 _3784_ (.A1(\bitty_inst.alu_inst.in_a[5] ),
    .A2(_1522_),
    .Y(_1297_),
    .B1(_1296_));
 sg13g2_o21ai_1 _3785_ (.B1(_1297_),
    .Y(_1298_),
    .A1(net729),
    .A2(net660));
 sg13g2_a22oi_1 _3786_ (.Y(_1299_),
    .B1(_1298_),
    .B2(net810),
    .A2(_1294_),
    .A1(\addr[5] ));
 sg13g2_a221oi_1 _3787_ (.B2(net815),
    .C1(\uart_inst.T0.bit_counter[1] ),
    .B1(_1299_),
    .A1(_1293_),
    .Y(_1300_),
    .A2(_1295_));
 sg13g2_nor2_1 _3788_ (.A(net802),
    .B(net789),
    .Y(_1301_));
 sg13g2_a21oi_1 _3789_ (.A1(\bitty_inst.alu_inst.in_a[6] ),
    .A2(_1522_),
    .Y(_1302_),
    .B1(_1301_));
 sg13g2_o21ai_1 _3790_ (.B1(_1302_),
    .Y(_1303_),
    .A1(net729),
    .A2(net694));
 sg13g2_a221oi_1 _3791_ (.B2(net810),
    .C1(net815),
    .B1(_1303_),
    .A1(\addr[6] ),
    .Y(_1304_),
    .A2(_1294_));
 sg13g2_a22oi_1 _3792_ (.Y(_1305_),
    .B1(_1623_),
    .B2(_0704_),
    .A2(net788),
    .A1(\bitty_inst.alu_inst.in_a[7] ));
 sg13g2_o21ai_1 _3793_ (.B1(_1305_),
    .Y(_1306_),
    .A1(_0036_),
    .A2(net789));
 sg13g2_a22oi_1 _3794_ (.Y(_1307_),
    .B1(_1306_),
    .B2(net810),
    .A2(_1294_),
    .A1(\addr[7] ));
 sg13g2_nand2_1 _3795_ (.Y(_1308_),
    .A(net815),
    .B(_1307_));
 sg13g2_nand2_1 _3796_ (.Y(_1309_),
    .A(\uart_inst.T0.bit_counter[1] ),
    .B(_1308_));
 sg13g2_o21ai_1 _3797_ (.B1(\uart_inst.T0.bit_counter[2] ),
    .Y(_1310_),
    .A1(_1304_),
    .A2(_1309_));
 sg13g2_nor2_1 _3798_ (.A(net805),
    .B(net789),
    .Y(_1311_));
 sg13g2_a21oi_1 _3799_ (.A1(\bitty_inst.alu_inst.in_a[3] ),
    .A2(net788),
    .Y(_1312_),
    .B1(_1311_));
 sg13g2_o21ai_1 _3800_ (.B1(_1312_),
    .Y(_1313_),
    .A1(net729),
    .A2(net693));
 sg13g2_a22oi_1 _3801_ (.Y(_1314_),
    .B1(_1313_),
    .B2(net810),
    .A2(_1294_),
    .A1(\addr[3] ));
 sg13g2_nor2_1 _3802_ (.A(net806),
    .B(net789),
    .Y(_1315_));
 sg13g2_a21oi_1 _3803_ (.A1(\bitty_inst.alu_inst.in_a[2] ),
    .A2(net788),
    .Y(_1316_),
    .B1(_1315_));
 sg13g2_o21ai_1 _3804_ (.B1(_1316_),
    .Y(_1317_),
    .A1(net729),
    .A2(net689));
 sg13g2_a221oi_1 _3805_ (.B2(net810),
    .C1(net815),
    .B1(_1317_),
    .A1(\addr[2] ),
    .Y(_1318_),
    .A2(_1294_));
 sg13g2_nand2b_1 _3806_ (.Y(_1319_),
    .B(\uart_inst.T0.bit_counter[1] ),
    .A_N(_1318_));
 sg13g2_a21oi_1 _3807_ (.A1(net815),
    .A2(_1314_),
    .Y(_1320_),
    .B1(_1319_));
 sg13g2_nand2_1 _3808_ (.Y(_1321_),
    .A(\bitty_inst.alu_inst.in_a[1] ),
    .B(net788));
 sg13g2_o21ai_1 _3809_ (.B1(net810),
    .Y(_1322_),
    .A1(_0042_),
    .A2(net789));
 sg13g2_o21ai_1 _3810_ (.B1(_1321_),
    .Y(_1323_),
    .A1(_1509_),
    .A2(_1516_));
 sg13g2_nor2_1 _3811_ (.A(_1322_),
    .B(_1323_),
    .Y(_1324_));
 sg13g2_o21ai_1 _3812_ (.B1(_1324_),
    .Y(_1325_),
    .A1(net729),
    .A2(net677));
 sg13g2_a21oi_1 _3813_ (.A1(\addr[1] ),
    .A2(\fi_inst.state[2] ),
    .Y(_1326_),
    .B1(net812));
 sg13g2_o21ai_1 _3814_ (.B1(_1326_),
    .Y(_1327_),
    .A1(_0074_),
    .A2(_1506_));
 sg13g2_nand3_1 _3815_ (.B(_1325_),
    .C(_1327_),
    .A(net815),
    .Y(_1328_));
 sg13g2_nor3_1 _3816_ (.A(\bitty_inst.cpu_inst.d_inst[2] ),
    .B(_1509_),
    .C(_1518_),
    .Y(_1329_));
 sg13g2_and2_1 _3817_ (.A(\bitty_inst.alu_inst.in_a[0] ),
    .B(net788),
    .X(_1330_));
 sg13g2_o21ai_1 _3818_ (.B1(net810),
    .Y(_1331_),
    .A1(_0043_),
    .A2(net789));
 sg13g2_nor3_1 _3819_ (.A(_1329_),
    .B(_1330_),
    .C(_1331_),
    .Y(_1332_));
 sg13g2_o21ai_1 _3820_ (.B1(_1332_),
    .Y(_1333_),
    .A1(net729),
    .A2(net667));
 sg13g2_a21oi_1 _3821_ (.A1(\addr[0] ),
    .A2(\fi_inst.state[2] ),
    .Y(_1334_),
    .B1(net812));
 sg13g2_o21ai_1 _3822_ (.B1(_1334_),
    .Y(_1335_),
    .A1(_0074_),
    .A2(_1506_));
 sg13g2_nand3b_1 _3823_ (.B(_1333_),
    .C(_1335_),
    .Y(_1336_),
    .A_N(net815));
 sg13g2_a21oi_1 _3824_ (.A1(_1328_),
    .A2(_1336_),
    .Y(_1337_),
    .B1(\uart_inst.T0.bit_counter[1] ));
 sg13g2_nor3_1 _3825_ (.A(\uart_inst.T0.bit_counter[2] ),
    .B(_1320_),
    .C(_1337_),
    .Y(_1338_));
 sg13g2_nor2b_1 _3826_ (.A(_1338_),
    .B_N(\uart_inst.T0.PS[1] ),
    .Y(_1339_));
 sg13g2_o21ai_1 _3827_ (.B1(_1339_),
    .Y(_1340_),
    .A1(_1300_),
    .A2(_1310_));
 sg13g2_nand2b_1 _3828_ (.Y(_0200_),
    .B(_1340_),
    .A_N(_1502_));
 sg13g2_dfrbp_1 _3829_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net27),
    .D(_0019_),
    .Q_N(_1873_),
    .Q(\uart_inst.R0.PS[0] ));
 sg13g2_dfrbp_1 _3830_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net28),
    .D(_0020_),
    .Q_N(_1874_),
    .Q(\uart_inst.R0.PS[1] ));
 sg13g2_dfrbp_1 _3831_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net29),
    .D(_0021_),
    .Q_N(_1875_),
    .Q(\uart_inst.R0.PS[2] ));
 sg13g2_dfrbp_1 _3832_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net30),
    .D(_0022_),
    .Q_N(_1876_),
    .Q(\uart_inst.R0.PS[3] ));
 sg13g2_dfrbp_1 _3833_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net74),
    .D(_0006_),
    .Q_N(_0073_),
    .Q(\bitty_inst.lsu_inst.rx_do ));
 sg13g2_dfrbp_1 _3834_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net26),
    .D(_0023_),
    .Q_N(_1872_),
    .Q(\uart_inst.R0.PS[5] ));
 sg13g2_dllrq_1 _3835_ (.D(\bitty_inst.lsu_inst.rx_data[0] ),
    .GATE_N(_0031_),
    .RESET_B(net31),
    .Q(\bitty_inst.d_instr[0] ));
 sg13g2_dllrq_1 _3836_ (.D(\bitty_inst.lsu_inst.rx_data[1] ),
    .GATE_N(_0031_),
    .RESET_B(net32),
    .Q(\bitty_inst.d_instr[1] ));
 sg13g2_dllrq_1 _3837_ (.D(\bitty_inst.lsu_inst.rx_data[2] ),
    .GATE_N(_0031_),
    .RESET_B(net33),
    .Q(\bitty_inst.d_instr[2] ));
 sg13g2_dllrq_1 _3838_ (.D(\bitty_inst.lsu_inst.rx_data[3] ),
    .GATE_N(_0031_),
    .RESET_B(net34),
    .Q(\bitty_inst.d_instr[3] ));
 sg13g2_dllrq_1 _3839_ (.D(\bitty_inst.lsu_inst.rx_data[4] ),
    .GATE_N(_0031_),
    .RESET_B(net35),
    .Q(\bitty_inst.d_instr[4] ));
 sg13g2_dllrq_1 _3840_ (.D(\bitty_inst.lsu_inst.rx_data[5] ),
    .GATE_N(_0031_),
    .RESET_B(net36),
    .Q(\bitty_inst.d_instr[5] ));
 sg13g2_dllrq_1 _3841_ (.D(\bitty_inst.lsu_inst.rx_data[6] ),
    .GATE_N(_0031_),
    .RESET_B(net37),
    .Q(\bitty_inst.d_instr[6] ));
 sg13g2_dllrq_1 _3842_ (.D(\bitty_inst.lsu_inst.rx_data[7] ),
    .GATE_N(_0031_),
    .RESET_B(net38),
    .Q(\bitty_inst.d_instr[7] ));
 sg13g2_dllrq_1 _3843_ (.D(\bitty_inst.lsu_inst.rx_data[0] ),
    .GATE_N(_0032_),
    .RESET_B(net39),
    .Q(\bitty_inst.d_instr[8] ));
 sg13g2_dllrq_1 _3844_ (.D(\bitty_inst.lsu_inst.rx_data[1] ),
    .GATE_N(_0032_),
    .RESET_B(net40),
    .Q(\bitty_inst.d_instr[9] ));
 sg13g2_dllrq_1 _3845_ (.D(\bitty_inst.lsu_inst.rx_data[2] ),
    .GATE_N(_0032_),
    .RESET_B(net41),
    .Q(\bitty_inst.d_instr[10] ));
 sg13g2_dllrq_1 _3846_ (.D(\bitty_inst.lsu_inst.rx_data[3] ),
    .GATE_N(_0032_),
    .RESET_B(net42),
    .Q(\bitty_inst.d_instr[11] ));
 sg13g2_dllrq_1 _3847_ (.D(\bitty_inst.lsu_inst.rx_data[4] ),
    .GATE_N(_0032_),
    .RESET_B(net43),
    .Q(\bitty_inst.d_instr[12] ));
 sg13g2_dllrq_1 _3848_ (.D(\bitty_inst.lsu_inst.rx_data[5] ),
    .GATE_N(_0032_),
    .RESET_B(net44),
    .Q(\bitty_inst.d_instr[13] ));
 sg13g2_dllrq_1 _3849_ (.D(\bitty_inst.lsu_inst.rx_data[6] ),
    .GATE_N(_0032_),
    .RESET_B(net45),
    .Q(\bitty_inst.d_instr[14] ));
 sg13g2_dllrq_1 _3850_ (.D(\bitty_inst.lsu_inst.rx_data[7] ),
    .GATE_N(_0032_),
    .RESET_B(net46),
    .Q(\bitty_inst.d_instr[15] ));
 sg13g2_dfrbp_1 _3851_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net270),
    .D(_0201_),
    .Q_N(_1871_),
    .Q(\bitty_inst.lsu_inst.state[0] ));
 sg13g2_dfrbp_1 _3852_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net269),
    .D(_0202_),
    .Q_N(_1870_),
    .Q(\bitty_inst.lsu_inst.state[1] ));
 sg13g2_dfrbp_1 _3853_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net268),
    .D(_0203_),
    .Q_N(_0072_),
    .Q(\bitty_inst.lsu_inst.state[2] ));
 sg13g2_dfrbp_1 _3854_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net267),
    .D(net922),
    .Q_N(_1869_),
    .Q(\uart_inst.T0.bit_counter[0] ));
 sg13g2_dfrbp_1 _3855_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net265),
    .D(net889),
    .Q_N(_1868_),
    .Q(\uart_inst.T0.bit_counter[1] ));
 sg13g2_dfrbp_1 _3856_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net263),
    .D(net650),
    .Q_N(_0071_),
    .Q(\uart_inst.T0.bit_counter[2] ));
 sg13g2_dfrbp_1 _3857_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net261),
    .D(_0207_),
    .Q_N(_0070_),
    .Q(\uart_inst.T0.clk_counter[0] ));
 sg13g2_dfrbp_1 _3858_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net260),
    .D(_0208_),
    .Q_N(_1867_),
    .Q(\uart_inst.T0.clk_counter[1] ));
 sg13g2_dfrbp_1 _3859_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net259),
    .D(net420),
    .Q_N(_0069_),
    .Q(\uart_inst.T0.clk_counter[2] ));
 sg13g2_dfrbp_1 _3860_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net258),
    .D(_0210_),
    .Q_N(_1866_),
    .Q(\uart_inst.T0.clk_counter[3] ));
 sg13g2_dfrbp_1 _3861_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net257),
    .D(_0211_),
    .Q_N(_0068_),
    .Q(\uart_inst.T0.clk_counter[4] ));
 sg13g2_dfrbp_1 _3862_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net256),
    .D(_0212_),
    .Q_N(_1865_),
    .Q(\uart_inst.T0.clk_counter[5] ));
 sg13g2_dfrbp_1 _3863_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net255),
    .D(net425),
    .Q_N(_0067_),
    .Q(\uart_inst.T0.clk_counter[6] ));
 sg13g2_dfrbp_1 _3864_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net254),
    .D(_0214_),
    .Q_N(_1864_),
    .Q(\uart_inst.T0.clk_counter[7] ));
 sg13g2_dfrbp_1 _3865_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net253),
    .D(_0215_),
    .Q_N(_0066_),
    .Q(\uart_inst.T0.clk_counter[8] ));
 sg13g2_dfrbp_1 _3866_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net252),
    .D(_0216_),
    .Q_N(_1863_),
    .Q(\uart_inst.T0.clk_counter[9] ));
 sg13g2_dfrbp_1 _3867_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net251),
    .D(_0217_),
    .Q_N(_0065_),
    .Q(\uart_inst.T0.clk_counter[10] ));
 sg13g2_dfrbp_1 _3868_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net250),
    .D(_0218_),
    .Q_N(_1862_),
    .Q(\uart_inst.T0.clk_counter[11] ));
 sg13g2_dfrbp_1 _3869_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net249),
    .D(_0219_),
    .Q_N(_1861_),
    .Q(\uart_inst.T0.clk_counter[12] ));
 sg13g2_dfrbp_1 _3870_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net248),
    .D(_0220_),
    .Q_N(_1860_),
    .Q(\bitty_inst.lsu_inst.rx_data[0] ));
 sg13g2_dfrbp_1 _3871_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net246),
    .D(net929),
    .Q_N(_1859_),
    .Q(\bitty_inst.lsu_inst.rx_data[1] ));
 sg13g2_dfrbp_1 _3872_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net244),
    .D(net925),
    .Q_N(_1858_),
    .Q(\bitty_inst.lsu_inst.rx_data[2] ));
 sg13g2_dfrbp_1 _3873_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net242),
    .D(_0223_),
    .Q_N(_1857_),
    .Q(\bitty_inst.lsu_inst.rx_data[3] ));
 sg13g2_dfrbp_1 _3874_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net240),
    .D(net946),
    .Q_N(_1856_),
    .Q(\bitty_inst.lsu_inst.rx_data[4] ));
 sg13g2_dfrbp_1 _3875_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net238),
    .D(_0225_),
    .Q_N(_1855_),
    .Q(\bitty_inst.lsu_inst.rx_data[5] ));
 sg13g2_dfrbp_1 _3876_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net236),
    .D(_0226_),
    .Q_N(_1854_),
    .Q(\bitty_inst.lsu_inst.rx_data[6] ));
 sg13g2_dfrbp_1 _3877_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net75),
    .D(_0227_),
    .Q_N(_1877_),
    .Q(\bitty_inst.lsu_inst.rx_data[7] ));
 sg13g2_dfrbp_1 _3878_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net76),
    .D(_0014_),
    .Q_N(_1878_),
    .Q(\fi_inst.state[0] ));
 sg13g2_dfrbp_1 _3879_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net77),
    .D(_0015_),
    .Q_N(_1879_),
    .Q(\fi_inst.state[1] ));
 sg13g2_dfrbp_1 _3880_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net78),
    .D(_0016_),
    .Q_N(_1880_),
    .Q(\fi_inst.state[2] ));
 sg13g2_dfrbp_1 _3881_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net79),
    .D(net321),
    .Q_N(_1881_),
    .Q(fetch_done));
 sg13g2_dfrbp_1 _3882_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net104),
    .D(_0017_),
    .Q_N(_0074_),
    .Q(\fi_inst.state[4] ));
 sg13g2_dfrbp_1 _3883_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net234),
    .D(_0018_),
    .Q_N(_1853_),
    .Q(\fi_inst.state[5] ));
 sg13g2_dfrbp_1 _3884_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net232),
    .D(net604),
    .Q_N(_0064_),
    .Q(\uart_inst.R0.clk_counter[0] ));
 sg13g2_dfrbp_1 _3885_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net230),
    .D(_0229_),
    .Q_N(_1852_),
    .Q(\uart_inst.R0.clk_counter[1] ));
 sg13g2_dfrbp_1 _3886_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net228),
    .D(_0230_),
    .Q_N(_0063_),
    .Q(\uart_inst.R0.clk_counter[2] ));
 sg13g2_dfrbp_1 _3887_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net226),
    .D(_0231_),
    .Q_N(_0062_),
    .Q(\uart_inst.R0.clk_counter[3] ));
 sg13g2_dfrbp_1 _3888_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net224),
    .D(_0232_),
    .Q_N(_0061_),
    .Q(\uart_inst.R0.clk_counter[4] ));
 sg13g2_dfrbp_1 _3889_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net222),
    .D(_0233_),
    .Q_N(_0060_),
    .Q(\uart_inst.R0.clk_counter[5] ));
 sg13g2_dfrbp_1 _3890_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net220),
    .D(_0234_),
    .Q_N(_0059_),
    .Q(\uart_inst.R0.clk_counter[6] ));
 sg13g2_dfrbp_1 _3891_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net218),
    .D(net869),
    .Q_N(_1851_),
    .Q(\uart_inst.R0.clk_counter[7] ));
 sg13g2_dfrbp_1 _3892_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net216),
    .D(_0236_),
    .Q_N(_0058_),
    .Q(\uart_inst.R0.clk_counter[8] ));
 sg13g2_dfrbp_1 _3893_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net214),
    .D(_0237_),
    .Q_N(_0057_),
    .Q(\uart_inst.R0.clk_counter[9] ));
 sg13g2_dfrbp_1 _3894_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net212),
    .D(_0238_),
    .Q_N(_0056_),
    .Q(\uart_inst.R0.clk_counter[10] ));
 sg13g2_dfrbp_1 _3895_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net210),
    .D(net956),
    .Q_N(_1850_),
    .Q(\uart_inst.R0.clk_counter[11] ));
 sg13g2_dfrbp_1 _3896_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net208),
    .D(_0240_),
    .Q_N(_0055_),
    .Q(\uart_inst.R0.clk_counter[12] ));
 sg13g2_dfrbp_1 _3897_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net206),
    .D(net949),
    .Q_N(_1849_),
    .Q(\uart_inst.R0.bit_counter[0] ));
 sg13g2_dfrbp_1 _3898_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net204),
    .D(net884),
    .Q_N(_1848_),
    .Q(\uart_inst.R0.bit_counter[1] ));
 sg13g2_dfrbp_1 _3899_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net202),
    .D(net644),
    .Q_N(_1847_),
    .Q(\uart_inst.R0.bit_counter[2] ));
 sg13g2_dfrbp_1 _3900_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net200),
    .D(net896),
    .Q_N(_0054_),
    .Q(\addr[0] ));
 sg13g2_dfrbp_1 _3901_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net198),
    .D(_0245_),
    .Q_N(_1846_),
    .Q(\addr[1] ));
 sg13g2_dfrbp_1 _3902_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net196),
    .D(_0246_),
    .Q_N(_1845_),
    .Q(\addr[2] ));
 sg13g2_dfrbp_1 _3903_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net194),
    .D(_0247_),
    .Q_N(_1844_),
    .Q(\addr[3] ));
 sg13g2_dfrbp_1 _3904_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net192),
    .D(net927),
    .Q_N(_0053_),
    .Q(\addr[4] ));
 sg13g2_dfrbp_1 _3905_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net190),
    .D(net931),
    .Q_N(_1843_),
    .Q(\addr[5] ));
 sg13g2_dfrbp_1 _3906_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net188),
    .D(net938),
    .Q_N(_1842_),
    .Q(\addr[6] ));
 sg13g2_dfrbp_1 _3907_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net105),
    .D(net933),
    .Q_N(_1882_),
    .Q(\addr[7] ));
 sg13g2_dfrbp_1 _3908_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net106),
    .D(net472),
    .Q_N(_1883_),
    .Q(\uart_inst.T0.PS[0] ));
 sg13g2_dfrbp_1 _3909_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net107),
    .D(_0025_),
    .Q_N(_1884_),
    .Q(\uart_inst.T0.PS[1] ));
 sg13g2_dfrbp_1 _3910_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net108),
    .D(_0026_),
    .Q_N(_1885_),
    .Q(\uart_inst.T0.PS[2] ));
 sg13g2_dfrbp_1 _3911_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net109),
    .D(_0007_),
    .Q_N(_0075_),
    .Q(\bitty_inst.lsu_inst.tx_done ));
 sg13g2_dfrbp_1 _3912_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net110),
    .D(net422),
    .Q_N(_1886_),
    .Q(\uart_inst.T0.PS[4] ));
 sg13g2_dfrbp_1 _3913_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net111),
    .D(net485),
    .Q_N(_1887_),
    .Q(\cur_state[0] ));
 sg13g2_dfrbp_1 _3914_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net112),
    .D(_0000_),
    .Q_N(_1888_),
    .Q(\cur_state[1] ));
 sg13g2_dfrbp_1 _3915_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net113),
    .D(_0001_),
    .Q_N(_1889_),
    .Q(\cur_state[2] ));
 sg13g2_dfrbp_1 _3916_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net114),
    .D(net436),
    .Q_N(_1890_),
    .Q(\cur_state[3] ));
 sg13g2_dfrbp_1 _3917_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net115),
    .D(net326),
    .Q_N(_1891_),
    .Q(\cur_state[4] ));
 sg13g2_dfrbp_1 _3918_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net116),
    .D(_0003_),
    .Q_N(_1892_),
    .Q(\bitty_inst.cpu_inst.run ));
 sg13g2_dfrbp_1 _3919_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net117),
    .D(_0004_),
    .Q_N(_1893_),
    .Q(\cur_state[6] ));
 sg13g2_dfrbp_1 _3920_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net118),
    .D(_0013_),
    .Q_N(_1894_),
    .Q(\cur_state[7] ));
 sg13g2_dfrbp_1 _3921_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net119),
    .D(net504),
    .Q_N(_1895_),
    .Q(\bitty_inst.cpu_inst.cur_state[0] ));
 sg13g2_dfrbp_1 _3922_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net63),
    .D(net640),
    .Q_N(_1896_),
    .Q(\bitty_inst.cpu_inst.cur_state[1] ));
 sg13g2_dfrbp_1 _3923_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net186),
    .D(_0010_),
    .Q_N(_0052_),
    .Q(\bitty_inst.cpu_inst.cur_state[2] ));
 sg13g2_dfrbp_1 _3924_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net184),
    .D(net411),
    .Q_N(_1841_),
    .Q(\bitty_inst.gen_dff[7].reg_out.mux_out[0] ));
 sg13g2_dfrbp_1 _3925_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net182),
    .D(net427),
    .Q_N(_1840_),
    .Q(\bitty_inst.gen_dff[7].reg_out.mux_out[1] ));
 sg13g2_dfrbp_1 _3926_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net180),
    .D(net365),
    .Q_N(_1839_),
    .Q(\bitty_inst.gen_dff[7].reg_out.mux_out[2] ));
 sg13g2_dfrbp_1 _3927_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net178),
    .D(net399),
    .Q_N(_1838_),
    .Q(\bitty_inst.gen_dff[7].reg_out.mux_out[3] ));
 sg13g2_dfrbp_1 _3928_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net176),
    .D(net407),
    .Q_N(_1837_),
    .Q(\bitty_inst.gen_dff[7].reg_out.mux_out[4] ));
 sg13g2_dfrbp_1 _3929_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net174),
    .D(net340),
    .Q_N(_1836_),
    .Q(\bitty_inst.gen_dff[7].reg_out.mux_out[5] ));
 sg13g2_dfrbp_1 _3930_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net172),
    .D(net387),
    .Q_N(_1835_),
    .Q(\bitty_inst.gen_dff[7].reg_out.mux_out[6] ));
 sg13g2_dfrbp_1 _3931_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net170),
    .D(net389),
    .Q_N(_1834_),
    .Q(\bitty_inst.gen_dff[7].reg_out.mux_out[7] ));
 sg13g2_dfrbp_1 _3932_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net168),
    .D(net361),
    .Q_N(_1833_),
    .Q(\bitty_inst.gen_dff[7].reg_out.mux_out[8] ));
 sg13g2_dfrbp_1 _3933_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net166),
    .D(net346),
    .Q_N(_1832_),
    .Q(\bitty_inst.gen_dff[7].reg_out.mux_out[9] ));
 sg13g2_dfrbp_1 _3934_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net164),
    .D(net438),
    .Q_N(_1831_),
    .Q(\bitty_inst.gen_dff[7].reg_out.mux_out[10] ));
 sg13g2_dfrbp_1 _3935_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net162),
    .D(net367),
    .Q_N(_1830_),
    .Q(\bitty_inst.gen_dff[7].reg_out.mux_out[11] ));
 sg13g2_dfrbp_1 _3936_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net160),
    .D(net383),
    .Q_N(_1829_),
    .Q(\bitty_inst.gen_dff[7].reg_out.mux_out[12] ));
 sg13g2_dfrbp_1 _3937_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net158),
    .D(net401),
    .Q_N(_1828_),
    .Q(\bitty_inst.gen_dff[7].reg_out.mux_out[13] ));
 sg13g2_dfrbp_1 _3938_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net156),
    .D(net330),
    .Q_N(_1827_),
    .Q(\bitty_inst.gen_dff[7].reg_out.mux_out[14] ));
 sg13g2_dfrbp_1 _3939_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net154),
    .D(net354),
    .Q_N(_1826_),
    .Q(\bitty_inst.gen_dff[7].reg_out.mux_out[15] ));
 sg13g2_dfrbp_1 _3940_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net152),
    .D(net409),
    .Q_N(_1825_),
    .Q(\bitty_inst.gen_dff[6].reg_out.mux_out[0] ));
 sg13g2_dfrbp_1 _3941_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net150),
    .D(net417),
    .Q_N(_1824_),
    .Q(\bitty_inst.gen_dff[6].reg_out.mux_out[1] ));
 sg13g2_dfrbp_1 _3942_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net148),
    .D(net371),
    .Q_N(_1823_),
    .Q(\bitty_inst.gen_dff[6].reg_out.mux_out[2] ));
 sg13g2_dfrbp_1 _3943_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net146),
    .D(net334),
    .Q_N(_1822_),
    .Q(\bitty_inst.gen_dff[6].reg_out.mux_out[3] ));
 sg13g2_dfrbp_1 _3944_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net144),
    .D(net397),
    .Q_N(_1821_),
    .Q(\bitty_inst.gen_dff[6].reg_out.mux_out[4] ));
 sg13g2_dfrbp_1 _3945_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net142),
    .D(net373),
    .Q_N(_1820_),
    .Q(\bitty_inst.gen_dff[6].reg_out.mux_out[5] ));
 sg13g2_dfrbp_1 _3946_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net140),
    .D(net391),
    .Q_N(_1819_),
    .Q(\bitty_inst.gen_dff[6].reg_out.mux_out[6] ));
 sg13g2_dfrbp_1 _3947_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net138),
    .D(net359),
    .Q_N(_1818_),
    .Q(\bitty_inst.gen_dff[6].reg_out.mux_out[7] ));
 sg13g2_dfrbp_1 _3948_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net136),
    .D(net405),
    .Q_N(_1817_),
    .Q(\bitty_inst.gen_dff[6].reg_out.mux_out[8] ));
 sg13g2_dfrbp_1 _3949_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net134),
    .D(net332),
    .Q_N(_1816_),
    .Q(\bitty_inst.gen_dff[6].reg_out.mux_out[9] ));
 sg13g2_dfrbp_1 _3950_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net132),
    .D(net348),
    .Q_N(_1815_),
    .Q(\bitty_inst.gen_dff[6].reg_out.mux_out[10] ));
 sg13g2_dfrbp_1 _3951_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net130),
    .D(net395),
    .Q_N(_1814_),
    .Q(\bitty_inst.gen_dff[6].reg_out.mux_out[11] ));
 sg13g2_dfrbp_1 _3952_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net128),
    .D(net393),
    .Q_N(_1813_),
    .Q(\bitty_inst.gen_dff[6].reg_out.mux_out[12] ));
 sg13g2_dfrbp_1 _3953_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net126),
    .D(net342),
    .Q_N(_1812_),
    .Q(\bitty_inst.gen_dff[6].reg_out.mux_out[13] ));
 sg13g2_dfrbp_1 _3954_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net124),
    .D(net379),
    .Q_N(_1811_),
    .Q(\bitty_inst.gen_dff[6].reg_out.mux_out[14] ));
 sg13g2_dfrbp_1 _3955_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net122),
    .D(net369),
    .Q_N(_1810_),
    .Q(\bitty_inst.gen_dff[6].reg_out.mux_out[15] ));
 sg13g2_dfrbp_1 _3956_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net120),
    .D(net433),
    .Q_N(_1809_),
    .Q(\bitty_inst.gen_dff[5].reg_out.mux_out[0] ));
 sg13g2_dfrbp_1 _3957_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net102),
    .D(net415),
    .Q_N(_1808_),
    .Q(\bitty_inst.gen_dff[5].reg_out.mux_out[1] ));
 sg13g2_dfrbp_1 _3958_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net100),
    .D(net350),
    .Q_N(_1807_),
    .Q(\bitty_inst.gen_dff[5].reg_out.mux_out[2] ));
 sg13g2_dfrbp_1 _3959_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net98),
    .D(net336),
    .Q_N(_1806_),
    .Q(\bitty_inst.gen_dff[5].reg_out.mux_out[3] ));
 sg13g2_dfrbp_1 _3960_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net96),
    .D(net429),
    .Q_N(_1805_),
    .Q(\bitty_inst.gen_dff[5].reg_out.mux_out[4] ));
 sg13g2_dfrbp_1 _3961_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net94),
    .D(net338),
    .Q_N(_1804_),
    .Q(\bitty_inst.gen_dff[5].reg_out.mux_out[5] ));
 sg13g2_dfrbp_1 _3962_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net92),
    .D(net363),
    .Q_N(_1803_),
    .Q(\bitty_inst.gen_dff[5].reg_out.mux_out[6] ));
 sg13g2_dfrbp_1 _3963_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net90),
    .D(net328),
    .Q_N(_1802_),
    .Q(\bitty_inst.gen_dff[5].reg_out.mux_out[7] ));
 sg13g2_dfrbp_1 _3964_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net88),
    .D(net352),
    .Q_N(_1801_),
    .Q(\bitty_inst.gen_dff[5].reg_out.mux_out[8] ));
 sg13g2_dfrbp_1 _3965_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net86),
    .D(net344),
    .Q_N(_1800_),
    .Q(\bitty_inst.gen_dff[5].reg_out.mux_out[9] ));
 sg13g2_dfrbp_1 _3966_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net84),
    .D(net375),
    .Q_N(_1799_),
    .Q(\bitty_inst.gen_dff[5].reg_out.mux_out[10] ));
 sg13g2_dfrbp_1 _3967_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net82),
    .D(net377),
    .Q_N(_1798_),
    .Q(\bitty_inst.gen_dff[5].reg_out.mux_out[11] ));
 sg13g2_dfrbp_1 _3968_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net80),
    .D(net381),
    .Q_N(_1797_),
    .Q(\bitty_inst.gen_dff[5].reg_out.mux_out[12] ));
 sg13g2_dfrbp_1 _3969_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net72),
    .D(net324),
    .Q_N(_1796_),
    .Q(\bitty_inst.gen_dff[5].reg_out.mux_out[13] ));
 sg13g2_dfrbp_1 _3970_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net70),
    .D(net357),
    .Q_N(_1795_),
    .Q(\bitty_inst.gen_dff[5].reg_out.mux_out[14] ));
 sg13g2_dfrbp_1 _3971_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net68),
    .D(net385),
    .Q_N(_1794_),
    .Q(\bitty_inst.gen_dff[5].reg_out.mux_out[15] ));
 sg13g2_dfrbp_1 _3972_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net66),
    .D(net466),
    .Q_N(_1793_),
    .Q(\bitty_inst.gen_dff[4].reg_out.mux_out[0] ));
 sg13g2_dfrbp_1 _3973_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net64),
    .D(net647),
    .Q_N(_1792_),
    .Q(\bitty_inst.gen_dff[4].reg_out.mux_out[1] ));
 sg13g2_dfrbp_1 _3974_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net62),
    .D(net522),
    .Q_N(_1791_),
    .Q(\bitty_inst.gen_dff[4].reg_out.mux_out[2] ));
 sg13g2_dfrbp_1 _3975_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net60),
    .D(net500),
    .Q_N(_1790_),
    .Q(\bitty_inst.gen_dff[4].reg_out.mux_out[3] ));
 sg13g2_dfrbp_1 _3976_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net58),
    .D(net624),
    .Q_N(_1789_),
    .Q(\bitty_inst.gen_dff[4].reg_out.mux_out[4] ));
 sg13g2_dfrbp_1 _3977_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net56),
    .D(net590),
    .Q_N(_1788_),
    .Q(\bitty_inst.gen_dff[4].reg_out.mux_out[5] ));
 sg13g2_dfrbp_1 _3978_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net54),
    .D(net554),
    .Q_N(_1787_),
    .Q(\bitty_inst.gen_dff[4].reg_out.mux_out[6] ));
 sg13g2_dfrbp_1 _3979_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net52),
    .D(net586),
    .Q_N(_1786_),
    .Q(\bitty_inst.gen_dff[4].reg_out.mux_out[7] ));
 sg13g2_dfrbp_1 _3980_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net50),
    .D(net584),
    .Q_N(_1785_),
    .Q(\bitty_inst.gen_dff[4].reg_out.mux_out[8] ));
 sg13g2_dfrbp_1 _3981_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net48),
    .D(_0081_),
    .Q_N(_1784_),
    .Q(\bitty_inst.gen_dff[4].reg_out.mux_out[9] ));
 sg13g2_dfrbp_1 _3982_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net25),
    .D(net460),
    .Q_N(_1783_),
    .Q(\bitty_inst.gen_dff[4].reg_out.mux_out[10] ));
 sg13g2_dfrbp_1 _3983_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net295),
    .D(net539),
    .Q_N(_1782_),
    .Q(\bitty_inst.gen_dff[4].reg_out.mux_out[11] ));
 sg13g2_dfrbp_1 _3984_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net293),
    .D(net453),
    .Q_N(_1781_),
    .Q(\bitty_inst.gen_dff[4].reg_out.mux_out[12] ));
 sg13g2_dfrbp_1 _3985_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net291),
    .D(net541),
    .Q_N(_1780_),
    .Q(\bitty_inst.gen_dff[4].reg_out.mux_out[13] ));
 sg13g2_dfrbp_1 _3986_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net289),
    .D(net464),
    .Q_N(_1779_),
    .Q(\bitty_inst.gen_dff[4].reg_out.mux_out[14] ));
 sg13g2_dfrbp_1 _3987_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net287),
    .D(net491),
    .Q_N(_1778_),
    .Q(\bitty_inst.gen_dff[4].reg_out.mux_out[15] ));
 sg13g2_dfrbp_1 _3988_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net285),
    .D(net601),
    .Q_N(_1777_),
    .Q(\bitty_inst.gen_dff[3].reg_out.mux_out[0] ));
 sg13g2_dfrbp_1 _3989_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net283),
    .D(net607),
    .Q_N(_1776_),
    .Q(\bitty_inst.gen_dff[3].reg_out.mux_out[1] ));
 sg13g2_dfrbp_1 _3990_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net281),
    .D(net537),
    .Q_N(_1775_),
    .Q(\bitty_inst.gen_dff[3].reg_out.mux_out[2] ));
 sg13g2_dfrbp_1 _3991_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net279),
    .D(net575),
    .Q_N(_1774_),
    .Q(\bitty_inst.gen_dff[3].reg_out.mux_out[3] ));
 sg13g2_dfrbp_1 _3992_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net277),
    .D(net566),
    .Q_N(_1773_),
    .Q(\bitty_inst.gen_dff[3].reg_out.mux_out[4] ));
 sg13g2_dfrbp_1 _3993_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net275),
    .D(net629),
    .Q_N(_1772_),
    .Q(\bitty_inst.gen_dff[3].reg_out.mux_out[5] ));
 sg13g2_dfrbp_1 _3994_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net273),
    .D(net502),
    .Q_N(_1771_),
    .Q(\bitty_inst.gen_dff[3].reg_out.mux_out[6] ));
 sg13g2_dfrbp_1 _3995_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net271),
    .D(net611),
    .Q_N(_1770_),
    .Q(\bitty_inst.gen_dff[3].reg_out.mux_out[7] ));
 sg13g2_dfrbp_1 _3996_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net264),
    .D(net512),
    .Q_N(_1769_),
    .Q(\bitty_inst.gen_dff[3].reg_out.mux_out[8] ));
 sg13g2_dfrbp_1 _3997_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net247),
    .D(_0097_),
    .Q_N(_1768_),
    .Q(\bitty_inst.gen_dff[3].reg_out.mux_out[9] ));
 sg13g2_dfrbp_1 _3998_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net243),
    .D(net556),
    .Q_N(_1767_),
    .Q(\bitty_inst.gen_dff[3].reg_out.mux_out[10] ));
 sg13g2_dfrbp_1 _3999_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net239),
    .D(net571),
    .Q_N(_1766_),
    .Q(\bitty_inst.gen_dff[3].reg_out.mux_out[11] ));
 sg13g2_dfrbp_1 _4000_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net235),
    .D(net474),
    .Q_N(_1765_),
    .Q(\bitty_inst.gen_dff[3].reg_out.mux_out[12] ));
 sg13g2_dfrbp_1 _4001_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net231),
    .D(net871),
    .Q_N(_1764_),
    .Q(\bitty_inst.gen_dff[3].reg_out.mux_out[13] ));
 sg13g2_dfrbp_1 _4002_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net227),
    .D(net528),
    .Q_N(_1763_),
    .Q(\bitty_inst.gen_dff[3].reg_out.mux_out[14] ));
 sg13g2_dfrbp_1 _4003_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net223),
    .D(net518),
    .Q_N(_1762_),
    .Q(\bitty_inst.gen_dff[3].reg_out.mux_out[15] ));
 sg13g2_dfrbp_1 _4004_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net219),
    .D(net520),
    .Q_N(_1761_),
    .Q(\bitty_inst.gen_dff[2].reg_out.mux_out[0] ));
 sg13g2_dfrbp_1 _4005_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net215),
    .D(net532),
    .Q_N(_1760_),
    .Q(\bitty_inst.gen_dff[2].reg_out.mux_out[1] ));
 sg13g2_dfrbp_1 _4006_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net211),
    .D(net482),
    .Q_N(_1759_),
    .Q(\bitty_inst.gen_dff[2].reg_out.mux_out[2] ));
 sg13g2_dfrbp_1 _4007_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net207),
    .D(net487),
    .Q_N(_1758_),
    .Q(\bitty_inst.gen_dff[2].reg_out.mux_out[3] ));
 sg13g2_dfrbp_1 _4008_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net203),
    .D(net476),
    .Q_N(_1757_),
    .Q(\bitty_inst.gen_dff[2].reg_out.mux_out[4] ));
 sg13g2_dfrbp_1 _4009_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net199),
    .D(net561),
    .Q_N(_1756_),
    .Q(\bitty_inst.gen_dff[2].reg_out.mux_out[5] ));
 sg13g2_dfrbp_1 _4010_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net195),
    .D(net613),
    .Q_N(_1755_),
    .Q(\bitty_inst.gen_dff[2].reg_out.mux_out[6] ));
 sg13g2_dfrbp_1 _4011_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net191),
    .D(net632),
    .Q_N(_1754_),
    .Q(\bitty_inst.gen_dff[2].reg_out.mux_out[7] ));
 sg13g2_dfrbp_1 _4012_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net187),
    .D(net626),
    .Q_N(_1753_),
    .Q(\bitty_inst.gen_dff[2].reg_out.mux_out[8] ));
 sg13g2_dfrbp_1 _4013_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net183),
    .D(_0113_),
    .Q_N(_1752_),
    .Q(\bitty_inst.gen_dff[2].reg_out.mux_out[9] ));
 sg13g2_dfrbp_1 _4014_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net179),
    .D(net526),
    .Q_N(_1751_),
    .Q(\bitty_inst.gen_dff[2].reg_out.mux_out[10] ));
 sg13g2_dfrbp_1 _4015_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net175),
    .D(net568),
    .Q_N(_1750_),
    .Q(\bitty_inst.gen_dff[2].reg_out.mux_out[11] ));
 sg13g2_dfrbp_1 _4016_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net171),
    .D(net470),
    .Q_N(_1749_),
    .Q(\bitty_inst.gen_dff[2].reg_out.mux_out[12] ));
 sg13g2_dfrbp_1 _4017_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net167),
    .D(net508),
    .Q_N(_1748_),
    .Q(\bitty_inst.gen_dff[2].reg_out.mux_out[13] ));
 sg13g2_dfrbp_1 _4018_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net163),
    .D(net530),
    .Q_N(_1747_),
    .Q(\bitty_inst.gen_dff[2].reg_out.mux_out[14] ));
 sg13g2_dfrbp_1 _4019_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net159),
    .D(net548),
    .Q_N(_1746_),
    .Q(\bitty_inst.gen_dff[2].reg_out.mux_out[15] ));
 sg13g2_dfrbp_1 _4020_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net155),
    .D(net545),
    .Q_N(_1745_),
    .Q(\bitty_inst.gen_dff[1].reg_out.mux_out[0] ));
 sg13g2_dfrbp_1 _4021_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net151),
    .D(net634),
    .Q_N(_1744_),
    .Q(\bitty_inst.gen_dff[1].reg_out.mux_out[1] ));
 sg13g2_dfrbp_1 _4022_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net147),
    .D(net514),
    .Q_N(_1743_),
    .Q(\bitty_inst.gen_dff[1].reg_out.mux_out[2] ));
 sg13g2_dfrbp_1 _4023_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net143),
    .D(net496),
    .Q_N(_1742_),
    .Q(\bitty_inst.gen_dff[1].reg_out.mux_out[3] ));
 sg13g2_dfrbp_1 _4024_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net139),
    .D(net578),
    .Q_N(_1741_),
    .Q(\bitty_inst.gen_dff[1].reg_out.mux_out[4] ));
 sg13g2_dfrbp_1 _4025_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net135),
    .D(net489),
    .Q_N(_1740_),
    .Q(\bitty_inst.gen_dff[1].reg_out.mux_out[5] ));
 sg13g2_dfrbp_1 _4026_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net131),
    .D(net510),
    .Q_N(_1739_),
    .Q(\bitty_inst.gen_dff[1].reg_out.mux_out[6] ));
 sg13g2_dfrbp_1 _4027_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net127),
    .D(net468),
    .Q_N(_1738_),
    .Q(\bitty_inst.gen_dff[1].reg_out.mux_out[7] ));
 sg13g2_dfrbp_1 _4028_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net123),
    .D(net588),
    .Q_N(_1737_),
    .Q(\bitty_inst.gen_dff[1].reg_out.mux_out[8] ));
 sg13g2_dfrbp_1 _4029_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net103),
    .D(_0129_),
    .Q_N(_1736_),
    .Q(\bitty_inst.gen_dff[1].reg_out.mux_out[9] ));
 sg13g2_dfrbp_1 _4030_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net99),
    .D(net550),
    .Q_N(_1735_),
    .Q(\bitty_inst.gen_dff[1].reg_out.mux_out[10] ));
 sg13g2_dfrbp_1 _4031_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net95),
    .D(net599),
    .Q_N(_1734_),
    .Q(\bitty_inst.gen_dff[1].reg_out.mux_out[11] ));
 sg13g2_dfrbp_1 _4032_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net91),
    .D(net615),
    .Q_N(_1733_),
    .Q(\bitty_inst.gen_dff[1].reg_out.mux_out[12] ));
 sg13g2_dfrbp_1 _4033_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net87),
    .D(net558),
    .Q_N(_1732_),
    .Q(\bitty_inst.gen_dff[1].reg_out.mux_out[13] ));
 sg13g2_dfrbp_1 _4034_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net83),
    .D(net552),
    .Q_N(_1731_),
    .Q(\bitty_inst.gen_dff[1].reg_out.mux_out[14] ));
 sg13g2_dfrbp_1 _4035_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net73),
    .D(net457),
    .Q_N(_1730_),
    .Q(\bitty_inst.gen_dff[1].reg_out.mux_out[15] ));
 sg13g2_dfrbp_1 _4036_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net69),
    .D(net593),
    .Q_N(_1729_),
    .Q(\bitty_inst.gen_dff[0].reg_out.mux_out[0] ));
 sg13g2_dfrbp_1 _4037_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net65),
    .D(net524),
    .Q_N(_1728_),
    .Q(\bitty_inst.gen_dff[0].reg_out.mux_out[1] ));
 sg13g2_dfrbp_1 _4038_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net61),
    .D(net516),
    .Q_N(_1727_),
    .Q(\bitty_inst.gen_dff[0].reg_out.mux_out[2] ));
 sg13g2_dfrbp_1 _4039_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net57),
    .D(net543),
    .Q_N(_1726_),
    .Q(\bitty_inst.gen_dff[0].reg_out.mux_out[3] ));
 sg13g2_dfrbp_1 _4040_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net53),
    .D(net535),
    .Q_N(_1725_),
    .Q(\bitty_inst.gen_dff[0].reg_out.mux_out[4] ));
 sg13g2_dfrbp_1 _4041_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net49),
    .D(net573),
    .Q_N(_1724_),
    .Q(\bitty_inst.gen_dff[0].reg_out.mux_out[5] ));
 sg13g2_dfrbp_1 _4042_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net315),
    .D(net506),
    .Q_N(_1723_),
    .Q(\bitty_inst.gen_dff[0].reg_out.mux_out[6] ));
 sg13g2_dfrbp_1 _4043_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net292),
    .D(net494),
    .Q_N(_1722_),
    .Q(\bitty_inst.gen_dff[0].reg_out.mux_out[7] ));
 sg13g2_dfrbp_1 _4044_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net288),
    .D(net580),
    .Q_N(_1721_),
    .Q(\bitty_inst.gen_dff[0].reg_out.mux_out[8] ));
 sg13g2_dfrbp_1 _4045_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net284),
    .D(_0145_),
    .Q_N(_1720_),
    .Q(\bitty_inst.gen_dff[0].reg_out.mux_out[9] ));
 sg13g2_dfrbp_1 _4046_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net280),
    .D(net621),
    .Q_N(_1719_),
    .Q(\bitty_inst.gen_dff[0].reg_out.mux_out[10] ));
 sg13g2_dfrbp_1 _4047_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net276),
    .D(net480),
    .Q_N(_1718_),
    .Q(\bitty_inst.gen_dff[0].reg_out.mux_out[11] ));
 sg13g2_dfrbp_1 _4048_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net272),
    .D(net595),
    .Q_N(_1717_),
    .Q(\bitty_inst.gen_dff[0].reg_out.mux_out[12] ));
 sg13g2_dfrbp_1 _4049_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net262),
    .D(net451),
    .Q_N(_1716_),
    .Q(\bitty_inst.gen_dff[0].reg_out.mux_out[13] ));
 sg13g2_dfrbp_1 _4050_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net241),
    .D(net564),
    .Q_N(_1715_),
    .Q(\bitty_inst.gen_dff[0].reg_out.mux_out[14] ));
 sg13g2_dfrbp_1 _4051_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net233),
    .D(net478),
    .Q_N(_1714_),
    .Q(\bitty_inst.gen_dff[0].reg_out.mux_out[15] ));
 sg13g2_dfrbp_1 _4052_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net225),
    .D(_0152_),
    .Q_N(_1713_),
    .Q(\bitty_inst.d_out[0] ));
 sg13g2_dfrbp_1 _4053_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net217),
    .D(_0153_),
    .Q_N(_1712_),
    .Q(\bitty_inst.d_out[1] ));
 sg13g2_dfrbp_1 _4054_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net209),
    .D(_0154_),
    .Q_N(_1711_),
    .Q(\bitty_inst.d_out[2] ));
 sg13g2_dfrbp_1 _4055_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net201),
    .D(_0155_),
    .Q_N(_1710_),
    .Q(\bitty_inst.d_out[3] ));
 sg13g2_dfrbp_1 _4056_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net193),
    .D(_0156_),
    .Q_N(_1709_),
    .Q(\bitty_inst.d_out[4] ));
 sg13g2_dfrbp_1 _4057_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net185),
    .D(_0157_),
    .Q_N(_1708_),
    .Q(\bitty_inst.d_out[5] ));
 sg13g2_dfrbp_1 _4058_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net177),
    .D(_0158_),
    .Q_N(_1707_),
    .Q(\bitty_inst.d_out[6] ));
 sg13g2_dfrbp_1 _4059_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net169),
    .D(_0159_),
    .Q_N(_1706_),
    .Q(\bitty_inst.d_out[7] ));
 sg13g2_dfrbp_1 _4060_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net161),
    .D(_0160_),
    .Q_N(_1705_),
    .Q(\bitty_inst.d_out[8] ));
 sg13g2_dfrbp_1 _4061_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net153),
    .D(_0161_),
    .Q_N(_1704_),
    .Q(\bitty_inst.d_out[9] ));
 sg13g2_dfrbp_1 _4062_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net145),
    .D(_0162_),
    .Q_N(_1703_),
    .Q(\bitty_inst.d_out[10] ));
 sg13g2_dfrbp_1 _4063_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net137),
    .D(_0163_),
    .Q_N(_1702_),
    .Q(\bitty_inst.d_out[11] ));
 sg13g2_dfrbp_1 _4064_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net129),
    .D(_0164_),
    .Q_N(_1701_),
    .Q(\bitty_inst.d_out[12] ));
 sg13g2_dfrbp_1 _4065_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net121),
    .D(_0165_),
    .Q_N(_1700_),
    .Q(\bitty_inst.d_out[13] ));
 sg13g2_dfrbp_1 _4066_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net97),
    .D(_0166_),
    .Q_N(_1699_),
    .Q(\bitty_inst.d_out[14] ));
 sg13g2_dfrbp_1 _4067_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net89),
    .D(_0167_),
    .Q_N(_1698_),
    .Q(\bitty_inst.d_out[15] ));
 sg13g2_dfrbp_1 _4068_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net81),
    .D(_0168_),
    .Q_N(_0051_),
    .Q(\bitty_inst.alu_inst.in_a[0] ));
 sg13g2_dfrbp_1 _4069_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net67),
    .D(_0169_),
    .Q_N(_0050_),
    .Q(\bitty_inst.alu_inst.in_a[1] ));
 sg13g2_dfrbp_1 _4070_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net59),
    .D(_0170_),
    .Q_N(_0049_),
    .Q(\bitty_inst.alu_inst.in_a[2] ));
 sg13g2_dfrbp_1 _4071_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net51),
    .D(_0171_),
    .Q_N(_0048_),
    .Q(\bitty_inst.alu_inst.in_a[3] ));
 sg13g2_dfrbp_1 _4072_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net294),
    .D(_0172_),
    .Q_N(_0047_),
    .Q(\bitty_inst.alu_inst.in_a[4] ));
 sg13g2_dfrbp_1 _4073_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net286),
    .D(_0173_),
    .Q_N(_0046_),
    .Q(\bitty_inst.alu_inst.in_a[5] ));
 sg13g2_dfrbp_1 _4074_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net278),
    .D(_0174_),
    .Q_N(_0045_),
    .Q(\bitty_inst.alu_inst.in_a[6] ));
 sg13g2_dfrbp_1 _4075_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net266),
    .D(_0175_),
    .Q_N(_0044_),
    .Q(\bitty_inst.alu_inst.in_a[7] ));
 sg13g2_dfrbp_1 _4076_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net237),
    .D(_0176_),
    .Q_N(_0043_),
    .Q(\bitty_inst.alu_inst.in_a[8] ));
 sg13g2_dfrbp_1 _4077_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net221),
    .D(_0177_),
    .Q_N(_0042_),
    .Q(\bitty_inst.alu_inst.in_a[9] ));
 sg13g2_dfrbp_1 _4078_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net205),
    .D(_0178_),
    .Q_N(_0041_),
    .Q(\bitty_inst.alu_inst.in_a[10] ));
 sg13g2_dfrbp_1 _4079_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net189),
    .D(_0179_),
    .Q_N(_0040_),
    .Q(\bitty_inst.alu_inst.in_a[11] ));
 sg13g2_dfrbp_1 _4080_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net173),
    .D(_0180_),
    .Q_N(_0039_),
    .Q(\bitty_inst.alu_inst.in_a[12] ));
 sg13g2_dfrbp_1 _4081_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net157),
    .D(_0181_),
    .Q_N(_0038_),
    .Q(\bitty_inst.alu_inst.in_a[13] ));
 sg13g2_dfrbp_1 _4082_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net141),
    .D(_0182_),
    .Q_N(_0037_),
    .Q(\bitty_inst.alu_inst.in_a[14] ));
 sg13g2_dfrbp_1 _4083_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net125),
    .D(_0183_),
    .Q_N(_0036_),
    .Q(\bitty_inst.alu_inst.in_a[15] ));
 sg13g2_dfrbp_1 _4084_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net93),
    .D(_0184_),
    .Q_N(_1697_),
    .Q(\bitty_inst.cpu_inst.d_inst[0] ));
 sg13g2_dfrbp_1 _4085_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net71),
    .D(_0185_),
    .Q_N(_1696_),
    .Q(\bitty_inst.cpu_inst.d_inst[1] ));
 sg13g2_dfrbp_1 _4086_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net55),
    .D(_0186_),
    .Q_N(_0035_),
    .Q(\bitty_inst.cpu_inst.d_inst[2] ));
 sg13g2_dfrbp_1 _4087_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net290),
    .D(_0187_),
    .Q_N(_1695_),
    .Q(\bitty_inst.cpu_inst.d_inst[3] ));
 sg13g2_dfrbp_1 _4088_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net274),
    .D(_0188_),
    .Q_N(_1694_),
    .Q(\bitty_inst.cpu_inst.d_inst[4] ));
 sg13g2_dfrbp_1 _4089_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net229),
    .D(_0189_),
    .Q_N(_1693_),
    .Q(\bitty_inst.cpu_inst.d_inst[5] ));
 sg13g2_dfrbp_1 _4090_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net197),
    .D(_0190_),
    .Q_N(_1692_),
    .Q(\bitty_inst.cpu_inst.d_inst[6] ));
 sg13g2_dfrbp_1 _4091_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net165),
    .D(_0191_),
    .Q_N(_1691_),
    .Q(\bitty_inst.cpu_inst.d_inst[7] ));
 sg13g2_dfrbp_1 _4092_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net133),
    .D(net403),
    .Q_N(_1690_),
    .Q(\bitty_inst.cpu_inst.d_inst[8] ));
 sg13g2_dfrbp_1 _4093_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net85),
    .D(_0193_),
    .Q_N(_1689_),
    .Q(\bitty_inst.cpu_inst.d_inst[9] ));
 sg13g2_dfrbp_1 _4094_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net47),
    .D(net440),
    .Q_N(_1688_),
    .Q(\bitty_inst.cpu_inst.d_inst[10] ));
 sg13g2_dfrbp_1 _4095_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net245),
    .D(_0195_),
    .Q_N(_0034_),
    .Q(\bitty_inst.cpu_inst.d_inst[11] ));
 sg13g2_dfrbp_1 _4096_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net181),
    .D(_0196_),
    .Q_N(_0033_),
    .Q(\bitty_inst.cpu_inst.d_inst[12] ));
 sg13g2_dfrbp_1 _4097_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net101),
    .D(_0197_),
    .Q_N(_1687_),
    .Q(\bitty_inst.cpu_inst.d_inst[13] ));
 sg13g2_dfrbp_1 _4098_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net282),
    .D(_0198_),
    .Q_N(_1686_),
    .Q(\bitty_inst.cpu_inst.d_inst[14] ));
 sg13g2_dfrbp_1 _4099_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net149),
    .D(_0199_),
    .Q_N(_1685_),
    .Q(\bitty_inst.cpu_inst.d_inst[15] ));
 sg13g2_dllrq_1 _4100_ (.D(\bitty_inst.lsu_inst.rx_data[0] ),
    .GATE_N(_0030_),
    .RESET_B(net296),
    .Q(\bitty_inst.data_to_ld[8] ));
 sg13g2_dllrq_1 _4101_ (.D(\bitty_inst.lsu_inst.rx_data[1] ),
    .GATE_N(_0030_),
    .RESET_B(net297),
    .Q(\bitty_inst.data_to_ld[9] ));
 sg13g2_dllrq_1 _4102_ (.D(\bitty_inst.lsu_inst.rx_data[2] ),
    .GATE_N(_0030_),
    .RESET_B(net298),
    .Q(\bitty_inst.data_to_ld[10] ));
 sg13g2_dllrq_1 _4103_ (.D(\bitty_inst.lsu_inst.rx_data[3] ),
    .GATE_N(_0030_),
    .RESET_B(net299),
    .Q(\bitty_inst.data_to_ld[11] ));
 sg13g2_dllrq_1 _4104_ (.D(\bitty_inst.lsu_inst.rx_data[4] ),
    .GATE_N(_0030_),
    .RESET_B(net300),
    .Q(\bitty_inst.data_to_ld[12] ));
 sg13g2_dllrq_1 _4105_ (.D(\bitty_inst.lsu_inst.rx_data[5] ),
    .GATE_N(_0030_),
    .RESET_B(net301),
    .Q(\bitty_inst.data_to_ld[13] ));
 sg13g2_dllrq_1 _4106_ (.D(\bitty_inst.lsu_inst.rx_data[6] ),
    .GATE_N(_0030_),
    .RESET_B(net302),
    .Q(\bitty_inst.data_to_ld[14] ));
 sg13g2_dllrq_1 _4107_ (.D(\bitty_inst.lsu_inst.rx_data[7] ),
    .GATE_N(_0030_),
    .RESET_B(net303),
    .Q(\bitty_inst.data_to_ld[15] ));
 sg13g2_dllrq_1 _4108_ (.D(\bitty_inst.lsu_inst.rx_data[0] ),
    .GATE_N(net781),
    .RESET_B(net304),
    .Q(\bitty_inst.data_to_ld[0] ));
 sg13g2_dllrq_1 _4109_ (.D(\bitty_inst.lsu_inst.rx_data[1] ),
    .GATE_N(net781),
    .RESET_B(net305),
    .Q(\bitty_inst.data_to_ld[1] ));
 sg13g2_dllrq_1 _4110_ (.D(\bitty_inst.lsu_inst.rx_data[2] ),
    .GATE_N(net781),
    .RESET_B(net306),
    .Q(\bitty_inst.data_to_ld[2] ));
 sg13g2_dllrq_1 _4111_ (.D(\bitty_inst.lsu_inst.rx_data[3] ),
    .GATE_N(net781),
    .RESET_B(net307),
    .Q(\bitty_inst.data_to_ld[3] ));
 sg13g2_dllrq_1 _4112_ (.D(\bitty_inst.lsu_inst.rx_data[4] ),
    .GATE_N(net781),
    .RESET_B(net308),
    .Q(\bitty_inst.data_to_ld[4] ));
 sg13g2_dllrq_1 _4113_ (.D(\bitty_inst.lsu_inst.rx_data[5] ),
    .GATE_N(net781),
    .RESET_B(net309),
    .Q(\bitty_inst.data_to_ld[5] ));
 sg13g2_dllrq_1 _4114_ (.D(\bitty_inst.lsu_inst.rx_data[6] ),
    .GATE_N(net781),
    .RESET_B(net310),
    .Q(\bitty_inst.data_to_ld[6] ));
 sg13g2_dllrq_1 _4115_ (.D(\bitty_inst.lsu_inst.rx_data[7] ),
    .GATE_N(net781),
    .RESET_B(net311),
    .Q(\bitty_inst.data_to_ld[7] ));
 sg13g2_dllrq_1 _4116_ (.D(_0304_),
    .GATE_N(_0028_),
    .RESET_B(net312),
    .Q(\bitty_inst.lsu_inst.next_state[0] ));
 sg13g2_dllrq_1 _4117_ (.D(_0305_),
    .GATE_N(_0028_),
    .RESET_B(net313),
    .Q(\bitty_inst.lsu_inst.next_state[1] ));
 sg13g2_dllrq_1 _4118_ (.D(_0306_),
    .GATE_N(_0028_),
    .RESET_B(net314),
    .Q(\bitty_inst.lsu_inst.next_state[2] ));
 sg13g2_dfrbp_1 _4119_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net213),
    .D(_0200_),
    .Q_N(_1684_),
    .Q(tx_data_bit));
 sg13g2_tiehi _3834__26 (.L_HI(net26));
 sg13g2_tiehi _3829__27 (.L_HI(net27));
 sg13g2_tiehi _3830__28 (.L_HI(net28));
 sg13g2_tiehi _3831__29 (.L_HI(net29));
 sg13g2_tiehi _3832__30 (.L_HI(net30));
 sg13g2_tiehi _3835__31 (.L_HI(net31));
 sg13g2_tiehi _3836__32 (.L_HI(net32));
 sg13g2_tiehi _3837__33 (.L_HI(net33));
 sg13g2_tiehi _3838__34 (.L_HI(net34));
 sg13g2_tiehi _3839__35 (.L_HI(net35));
 sg13g2_tiehi _3840__36 (.L_HI(net36));
 sg13g2_tiehi _3841__37 (.L_HI(net37));
 sg13g2_tiehi _3842__38 (.L_HI(net38));
 sg13g2_tiehi _3843__39 (.L_HI(net39));
 sg13g2_tiehi _3844__40 (.L_HI(net40));
 sg13g2_tiehi _3845__41 (.L_HI(net41));
 sg13g2_tiehi _3846__42 (.L_HI(net42));
 sg13g2_tiehi _3847__43 (.L_HI(net43));
 sg13g2_tiehi _3848__44 (.L_HI(net44));
 sg13g2_tiehi _3849__45 (.L_HI(net45));
 sg13g2_tiehi _3850__46 (.L_HI(net46));
 sg13g2_tiehi _4094__47 (.L_HI(net47));
 sg13g2_tiehi _3981__48 (.L_HI(net48));
 sg13g2_tiehi _4041__49 (.L_HI(net49));
 sg13g2_tiehi _3980__50 (.L_HI(net50));
 sg13g2_tiehi _4071__51 (.L_HI(net51));
 sg13g2_tiehi _3979__52 (.L_HI(net52));
 sg13g2_tiehi _4040__53 (.L_HI(net53));
 sg13g2_tiehi _3978__54 (.L_HI(net54));
 sg13g2_tiehi _4086__55 (.L_HI(net55));
 sg13g2_tiehi _3977__56 (.L_HI(net56));
 sg13g2_tiehi _4039__57 (.L_HI(net57));
 sg13g2_tiehi _3976__58 (.L_HI(net58));
 sg13g2_tiehi _4070__59 (.L_HI(net59));
 sg13g2_tiehi _3975__60 (.L_HI(net60));
 sg13g2_tiehi _4038__61 (.L_HI(net61));
 sg13g2_tiehi _3974__62 (.L_HI(net62));
 sg13g2_tiehi _3922__63 (.L_HI(net63));
 sg13g2_tiehi _3973__64 (.L_HI(net64));
 sg13g2_tiehi _4037__65 (.L_HI(net65));
 sg13g2_tiehi _3972__66 (.L_HI(net66));
 sg13g2_tiehi _4069__67 (.L_HI(net67));
 sg13g2_tiehi _3971__68 (.L_HI(net68));
 sg13g2_tiehi _4036__69 (.L_HI(net69));
 sg13g2_tiehi _3970__70 (.L_HI(net70));
 sg13g2_tiehi _4085__71 (.L_HI(net71));
 sg13g2_tiehi _3969__72 (.L_HI(net72));
 sg13g2_tiehi _4035__73 (.L_HI(net73));
 sg13g2_tiehi _3833__74 (.L_HI(net74));
 sg13g2_tiehi _3877__75 (.L_HI(net75));
 sg13g2_tiehi _3878__76 (.L_HI(net76));
 sg13g2_tiehi _3879__77 (.L_HI(net77));
 sg13g2_tiehi _3880__78 (.L_HI(net78));
 sg13g2_tiehi _3881__79 (.L_HI(net79));
 sg13g2_tiehi _3968__80 (.L_HI(net80));
 sg13g2_tiehi _4068__81 (.L_HI(net81));
 sg13g2_tiehi _3967__82 (.L_HI(net82));
 sg13g2_tiehi _4034__83 (.L_HI(net83));
 sg13g2_tiehi _3966__84 (.L_HI(net84));
 sg13g2_tiehi _4093__85 (.L_HI(net85));
 sg13g2_tiehi _3965__86 (.L_HI(net86));
 sg13g2_tiehi _4033__87 (.L_HI(net87));
 sg13g2_tiehi _3964__88 (.L_HI(net88));
 sg13g2_tiehi _4067__89 (.L_HI(net89));
 sg13g2_tiehi _3963__90 (.L_HI(net90));
 sg13g2_tiehi _4032__91 (.L_HI(net91));
 sg13g2_tiehi _3962__92 (.L_HI(net92));
 sg13g2_tiehi _4084__93 (.L_HI(net93));
 sg13g2_tiehi _3961__94 (.L_HI(net94));
 sg13g2_tiehi _4031__95 (.L_HI(net95));
 sg13g2_tiehi _3960__96 (.L_HI(net96));
 sg13g2_tiehi _4066__97 (.L_HI(net97));
 sg13g2_tiehi _3959__98 (.L_HI(net98));
 sg13g2_tiehi _4030__99 (.L_HI(net99));
 sg13g2_tiehi _3958__100 (.L_HI(net100));
 sg13g2_tiehi _4097__101 (.L_HI(net101));
 sg13g2_tiehi _3957__102 (.L_HI(net102));
 sg13g2_tiehi _4029__103 (.L_HI(net103));
 sg13g2_tiehi _3882__104 (.L_HI(net104));
 sg13g2_tiehi _3907__105 (.L_HI(net105));
 sg13g2_tiehi _3908__106 (.L_HI(net106));
 sg13g2_tiehi _3909__107 (.L_HI(net107));
 sg13g2_tiehi _3910__108 (.L_HI(net108));
 sg13g2_tiehi _3911__109 (.L_HI(net109));
 sg13g2_tiehi _3912__110 (.L_HI(net110));
 sg13g2_tiehi _3913__111 (.L_HI(net111));
 sg13g2_tiehi _3914__112 (.L_HI(net112));
 sg13g2_tiehi _3915__113 (.L_HI(net113));
 sg13g2_tiehi _3916__114 (.L_HI(net114));
 sg13g2_tiehi _3917__115 (.L_HI(net115));
 sg13g2_tiehi _3918__116 (.L_HI(net116));
 sg13g2_tiehi _3919__117 (.L_HI(net117));
 sg13g2_tiehi _3920__118 (.L_HI(net118));
 sg13g2_tiehi _3921__119 (.L_HI(net119));
 sg13g2_tiehi _3956__120 (.L_HI(net120));
 sg13g2_tiehi _4065__121 (.L_HI(net121));
 sg13g2_tiehi _3955__122 (.L_HI(net122));
 sg13g2_tiehi _4028__123 (.L_HI(net123));
 sg13g2_tiehi _3954__124 (.L_HI(net124));
 sg13g2_tiehi _4083__125 (.L_HI(net125));
 sg13g2_tiehi _3953__126 (.L_HI(net126));
 sg13g2_tiehi _4027__127 (.L_HI(net127));
 sg13g2_tiehi _3952__128 (.L_HI(net128));
 sg13g2_tiehi _4064__129 (.L_HI(net129));
 sg13g2_tiehi _3951__130 (.L_HI(net130));
 sg13g2_tiehi _4026__131 (.L_HI(net131));
 sg13g2_tiehi _3950__132 (.L_HI(net132));
 sg13g2_tiehi _4092__133 (.L_HI(net133));
 sg13g2_tiehi _3949__134 (.L_HI(net134));
 sg13g2_tiehi _4025__135 (.L_HI(net135));
 sg13g2_tiehi _3948__136 (.L_HI(net136));
 sg13g2_tiehi _4063__137 (.L_HI(net137));
 sg13g2_tiehi _3947__138 (.L_HI(net138));
 sg13g2_tiehi _4024__139 (.L_HI(net139));
 sg13g2_tiehi _3946__140 (.L_HI(net140));
 sg13g2_tiehi _4082__141 (.L_HI(net141));
 sg13g2_tiehi _3945__142 (.L_HI(net142));
 sg13g2_tiehi _4023__143 (.L_HI(net143));
 sg13g2_tiehi _3944__144 (.L_HI(net144));
 sg13g2_tiehi _4062__145 (.L_HI(net145));
 sg13g2_tiehi _3943__146 (.L_HI(net146));
 sg13g2_tiehi _4022__147 (.L_HI(net147));
 sg13g2_tiehi _3942__148 (.L_HI(net148));
 sg13g2_tiehi _4099__149 (.L_HI(net149));
 sg13g2_tiehi _3941__150 (.L_HI(net150));
 sg13g2_tiehi _4021__151 (.L_HI(net151));
 sg13g2_tiehi _3940__152 (.L_HI(net152));
 sg13g2_tiehi _4061__153 (.L_HI(net153));
 sg13g2_tiehi _3939__154 (.L_HI(net154));
 sg13g2_tiehi _4020__155 (.L_HI(net155));
 sg13g2_tiehi _3938__156 (.L_HI(net156));
 sg13g2_tiehi _4081__157 (.L_HI(net157));
 sg13g2_tiehi _3937__158 (.L_HI(net158));
 sg13g2_tiehi _4019__159 (.L_HI(net159));
 sg13g2_tiehi _3936__160 (.L_HI(net160));
 sg13g2_tiehi _4060__161 (.L_HI(net161));
 sg13g2_tiehi _3935__162 (.L_HI(net162));
 sg13g2_tiehi _4018__163 (.L_HI(net163));
 sg13g2_tiehi _3934__164 (.L_HI(net164));
 sg13g2_tiehi _4091__165 (.L_HI(net165));
 sg13g2_tiehi _3933__166 (.L_HI(net166));
 sg13g2_tiehi _4017__167 (.L_HI(net167));
 sg13g2_tiehi _3932__168 (.L_HI(net168));
 sg13g2_tiehi _4059__169 (.L_HI(net169));
 sg13g2_tiehi _3931__170 (.L_HI(net170));
 sg13g2_tiehi _4016__171 (.L_HI(net171));
 sg13g2_tiehi _3930__172 (.L_HI(net172));
 sg13g2_tiehi _4080__173 (.L_HI(net173));
 sg13g2_tiehi _3929__174 (.L_HI(net174));
 sg13g2_tiehi _4015__175 (.L_HI(net175));
 sg13g2_tiehi _3928__176 (.L_HI(net176));
 sg13g2_tiehi _4058__177 (.L_HI(net177));
 sg13g2_tiehi _3927__178 (.L_HI(net178));
 sg13g2_tiehi _4014__179 (.L_HI(net179));
 sg13g2_tiehi _3926__180 (.L_HI(net180));
 sg13g2_tiehi _4096__181 (.L_HI(net181));
 sg13g2_tiehi _3925__182 (.L_HI(net182));
 sg13g2_tiehi _4013__183 (.L_HI(net183));
 sg13g2_tiehi _3924__184 (.L_HI(net184));
 sg13g2_tiehi _4057__185 (.L_HI(net185));
 sg13g2_tiehi _3923__186 (.L_HI(net186));
 sg13g2_tiehi _4012__187 (.L_HI(net187));
 sg13g2_tiehi _3906__188 (.L_HI(net188));
 sg13g2_tiehi _4079__189 (.L_HI(net189));
 sg13g2_tiehi _3905__190 (.L_HI(net190));
 sg13g2_tiehi _4011__191 (.L_HI(net191));
 sg13g2_tiehi _3904__192 (.L_HI(net192));
 sg13g2_tiehi _4056__193 (.L_HI(net193));
 sg13g2_tiehi _3903__194 (.L_HI(net194));
 sg13g2_tiehi _4010__195 (.L_HI(net195));
 sg13g2_tiehi _3902__196 (.L_HI(net196));
 sg13g2_tiehi _4090__197 (.L_HI(net197));
 sg13g2_tiehi _3901__198 (.L_HI(net198));
 sg13g2_tiehi _4009__199 (.L_HI(net199));
 sg13g2_tiehi _3900__200 (.L_HI(net200));
 sg13g2_tiehi _4055__201 (.L_HI(net201));
 sg13g2_tiehi _3899__202 (.L_HI(net202));
 sg13g2_tiehi _4008__203 (.L_HI(net203));
 sg13g2_tiehi _3898__204 (.L_HI(net204));
 sg13g2_tiehi _4078__205 (.L_HI(net205));
 sg13g2_tiehi _3897__206 (.L_HI(net206));
 sg13g2_tiehi _4007__207 (.L_HI(net207));
 sg13g2_tiehi _3896__208 (.L_HI(net208));
 sg13g2_tiehi _4054__209 (.L_HI(net209));
 sg13g2_tiehi _3895__210 (.L_HI(net210));
 sg13g2_tiehi _4006__211 (.L_HI(net211));
 sg13g2_tiehi _3894__212 (.L_HI(net212));
 sg13g2_tiehi _4119__213 (.L_HI(net213));
 sg13g2_tiehi _3893__214 (.L_HI(net214));
 sg13g2_tiehi _4005__215 (.L_HI(net215));
 sg13g2_tiehi _3892__216 (.L_HI(net216));
 sg13g2_tiehi _4053__217 (.L_HI(net217));
 sg13g2_tiehi _3891__218 (.L_HI(net218));
 sg13g2_tiehi _4004__219 (.L_HI(net219));
 sg13g2_tiehi _3890__220 (.L_HI(net220));
 sg13g2_tiehi _4077__221 (.L_HI(net221));
 sg13g2_tiehi _3889__222 (.L_HI(net222));
 sg13g2_tiehi _4003__223 (.L_HI(net223));
 sg13g2_tiehi _3888__224 (.L_HI(net224));
 sg13g2_tiehi _4052__225 (.L_HI(net225));
 sg13g2_tiehi _3887__226 (.L_HI(net226));
 sg13g2_tiehi _4002__227 (.L_HI(net227));
 sg13g2_tiehi _3886__228 (.L_HI(net228));
 sg13g2_tiehi _4089__229 (.L_HI(net229));
 sg13g2_tiehi _3885__230 (.L_HI(net230));
 sg13g2_tiehi _4001__231 (.L_HI(net231));
 sg13g2_tiehi _3884__232 (.L_HI(net232));
 sg13g2_tiehi _4051__233 (.L_HI(net233));
 sg13g2_tiehi _3883__234 (.L_HI(net234));
 sg13g2_tiehi _4000__235 (.L_HI(net235));
 sg13g2_tiehi _3876__236 (.L_HI(net236));
 sg13g2_tiehi _4076__237 (.L_HI(net237));
 sg13g2_tiehi _3875__238 (.L_HI(net238));
 sg13g2_tiehi _3999__239 (.L_HI(net239));
 sg13g2_tiehi _3874__240 (.L_HI(net240));
 sg13g2_tiehi _4050__241 (.L_HI(net241));
 sg13g2_tiehi _3873__242 (.L_HI(net242));
 sg13g2_tiehi _3998__243 (.L_HI(net243));
 sg13g2_tiehi _3872__244 (.L_HI(net244));
 sg13g2_tiehi _4095__245 (.L_HI(net245));
 sg13g2_tiehi _3871__246 (.L_HI(net246));
 sg13g2_tiehi _3997__247 (.L_HI(net247));
 sg13g2_tiehi _3870__248 (.L_HI(net248));
 sg13g2_tiehi _3869__249 (.L_HI(net249));
 sg13g2_tiehi _3868__250 (.L_HI(net250));
 sg13g2_tiehi _3867__251 (.L_HI(net251));
 sg13g2_tiehi _3866__252 (.L_HI(net252));
 sg13g2_tiehi _3865__253 (.L_HI(net253));
 sg13g2_tiehi _3864__254 (.L_HI(net254));
 sg13g2_tiehi _3863__255 (.L_HI(net255));
 sg13g2_tiehi _3862__256 (.L_HI(net256));
 sg13g2_tiehi _3861__257 (.L_HI(net257));
 sg13g2_tiehi _3860__258 (.L_HI(net258));
 sg13g2_tiehi _3859__259 (.L_HI(net259));
 sg13g2_tiehi _3858__260 (.L_HI(net260));
 sg13g2_tiehi _3857__261 (.L_HI(net261));
 sg13g2_tiehi _4049__262 (.L_HI(net262));
 sg13g2_tiehi _3856__263 (.L_HI(net263));
 sg13g2_tiehi _3996__264 (.L_HI(net264));
 sg13g2_tiehi _3855__265 (.L_HI(net265));
 sg13g2_tiehi _4075__266 (.L_HI(net266));
 sg13g2_tiehi _3854__267 (.L_HI(net267));
 sg13g2_tiehi _3853__268 (.L_HI(net268));
 sg13g2_tiehi _3852__269 (.L_HI(net269));
 sg13g2_tiehi _3851__270 (.L_HI(net270));
 sg13g2_tiehi _3995__271 (.L_HI(net271));
 sg13g2_tiehi _4048__272 (.L_HI(net272));
 sg13g2_tiehi _3994__273 (.L_HI(net273));
 sg13g2_tiehi _4088__274 (.L_HI(net274));
 sg13g2_tiehi _3993__275 (.L_HI(net275));
 sg13g2_tiehi _4047__276 (.L_HI(net276));
 sg13g2_tiehi _3992__277 (.L_HI(net277));
 sg13g2_tiehi _4074__278 (.L_HI(net278));
 sg13g2_tiehi _3991__279 (.L_HI(net279));
 sg13g2_tiehi _4046__280 (.L_HI(net280));
 sg13g2_tiehi _3990__281 (.L_HI(net281));
 sg13g2_tiehi _4098__282 (.L_HI(net282));
 sg13g2_tiehi _3989__283 (.L_HI(net283));
 sg13g2_tiehi _4045__284 (.L_HI(net284));
 sg13g2_tiehi _3988__285 (.L_HI(net285));
 sg13g2_tiehi _4073__286 (.L_HI(net286));
 sg13g2_tiehi _3987__287 (.L_HI(net287));
 sg13g2_tiehi _4044__288 (.L_HI(net288));
 sg13g2_tiehi _3986__289 (.L_HI(net289));
 sg13g2_tiehi _4087__290 (.L_HI(net290));
 sg13g2_tiehi _3985__291 (.L_HI(net291));
 sg13g2_tiehi _4043__292 (.L_HI(net292));
 sg13g2_tiehi _3984__293 (.L_HI(net293));
 sg13g2_tiehi _4072__294 (.L_HI(net294));
 sg13g2_tiehi _3983__295 (.L_HI(net295));
 sg13g2_tiehi _4100__296 (.L_HI(net296));
 sg13g2_tiehi _4101__297 (.L_HI(net297));
 sg13g2_tiehi _4102__298 (.L_HI(net298));
 sg13g2_tiehi _4103__299 (.L_HI(net299));
 sg13g2_tiehi _4104__300 (.L_HI(net300));
 sg13g2_tiehi _4105__301 (.L_HI(net301));
 sg13g2_tiehi _4106__302 (.L_HI(net302));
 sg13g2_tiehi _4107__303 (.L_HI(net303));
 sg13g2_tiehi _4108__304 (.L_HI(net304));
 sg13g2_tiehi _4109__305 (.L_HI(net305));
 sg13g2_tiehi _4110__306 (.L_HI(net306));
 sg13g2_tiehi _4111__307 (.L_HI(net307));
 sg13g2_tiehi _4112__308 (.L_HI(net308));
 sg13g2_tiehi _4113__309 (.L_HI(net309));
 sg13g2_tiehi _4114__310 (.L_HI(net310));
 sg13g2_tiehi _4115__311 (.L_HI(net311));
 sg13g2_tiehi _4116__312 (.L_HI(net312));
 sg13g2_tiehi _4117__313 (.L_HI(net313));
 sg13g2_tiehi _4118__314 (.L_HI(net314));
 sg13g2_tiehi _4042__315 (.L_HI(net315));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_bitty_3 (.L_LO(net3));
 sg13g2_tielo tt_um_bitty_4 (.L_LO(net4));
 sg13g2_tielo tt_um_bitty_5 (.L_LO(net5));
 sg13g2_tielo tt_um_bitty_6 (.L_LO(net6));
 sg13g2_tielo tt_um_bitty_7 (.L_LO(net7));
 sg13g2_tielo tt_um_bitty_8 (.L_LO(net8));
 sg13g2_tielo tt_um_bitty_9 (.L_LO(net9));
 sg13g2_tielo tt_um_bitty_10 (.L_LO(net10));
 sg13g2_tielo tt_um_bitty_11 (.L_LO(net11));
 sg13g2_tielo tt_um_bitty_12 (.L_LO(net12));
 sg13g2_tielo tt_um_bitty_13 (.L_LO(net13));
 sg13g2_tielo tt_um_bitty_14 (.L_LO(net14));
 sg13g2_tielo tt_um_bitty_15 (.L_LO(net15));
 sg13g2_tielo tt_um_bitty_16 (.L_LO(net16));
 sg13g2_tielo tt_um_bitty_17 (.L_LO(net17));
 sg13g2_tielo tt_um_bitty_18 (.L_LO(net18));
 sg13g2_tielo tt_um_bitty_19 (.L_LO(net19));
 sg13g2_tielo tt_um_bitty_20 (.L_LO(net20));
 sg13g2_tielo tt_um_bitty_21 (.L_LO(net21));
 sg13g2_tielo tt_um_bitty_22 (.L_LO(net22));
 sg13g2_tielo tt_um_bitty_23 (.L_LO(net23));
 sg13g2_tielo tt_um_bitty_24 (.L_LO(net24));
 sg13g2_tiehi _3982__25 (.L_HI(net25));
 sg13g2_buf_1 _4434_ (.A(tx_data_bit),
    .X(uo_out[0]));
 sg13g2_buf_2 fanout652 (.A(_0318_),
    .X(net652));
 sg13g2_buf_4 fanout653 (.X(net653),
    .A(_1652_));
 sg13g2_buf_2 fanout654 (.A(_1652_),
    .X(net654));
 sg13g2_buf_4 fanout655 (.X(net655),
    .A(_1584_));
 sg13g2_buf_2 fanout656 (.A(_0980_),
    .X(net656));
 sg13g2_buf_1 fanout657 (.A(_0980_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_0734_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_0734_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_0725_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_0725_),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(_0681_),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(_0672_),
    .X(net663));
 sg13g2_buf_4 fanout664 (.X(net664),
    .A(net666));
 sg13g2_buf_4 fanout665 (.X(net665),
    .A(_0788_));
 sg13g2_buf_2 fanout666 (.A(_0788_),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(net668),
    .X(net667));
 sg13g2_buf_1 fanout668 (.A(_0787_),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(net672),
    .X(net669));
 sg13g2_buf_1 fanout670 (.A(net672),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_1 fanout672 (.A(net673),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(_0787_),
    .X(net673));
 sg13g2_buf_4 fanout674 (.X(net674),
    .A(net675));
 sg13g2_buf_4 fanout675 (.X(net675),
    .A(net676));
 sg13g2_buf_4 fanout676 (.X(net676),
    .A(_0776_));
 sg13g2_buf_2 fanout677 (.A(net678),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(_0775_),
    .X(net678));
 sg13g2_buf_4 fanout679 (.X(net679),
    .A(net681));
 sg13g2_buf_4 fanout680 (.X(net680),
    .A(net681));
 sg13g2_buf_2 fanout681 (.A(net682),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(_0775_),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(net685),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(net685),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(net686),
    .X(net685));
 sg13g2_buf_4 fanout686 (.X(net686),
    .A(_0762_));
 sg13g2_buf_4 fanout687 (.X(net687),
    .A(net688));
 sg13g2_buf_2 fanout688 (.A(_0761_),
    .X(net688));
 sg13g2_buf_4 fanout689 (.X(net689),
    .A(_0761_));
 sg13g2_buf_4 fanout690 (.X(net690),
    .A(net692));
 sg13g2_buf_1 fanout691 (.A(net692),
    .X(net691));
 sg13g2_buf_4 fanout692 (.X(net692),
    .A(_0747_));
 sg13g2_buf_4 fanout693 (.X(net693),
    .A(_0746_));
 sg13g2_buf_2 fanout694 (.A(_0715_),
    .X(net694));
 sg13g2_buf_1 fanout695 (.A(_0715_),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(_0416_),
    .X(net696));
 sg13g2_buf_4 fanout697 (.X(net697),
    .A(_0908_));
 sg13g2_buf_1 fanout698 (.A(_0908_),
    .X(net698));
 sg13g2_buf_4 fanout699 (.X(net699),
    .A(_0849_));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(_0849_));
 sg13g2_buf_2 fanout701 (.A(_0844_),
    .X(net701));
 sg13g2_buf_4 fanout702 (.X(net702),
    .A(_0841_));
 sg13g2_buf_2 fanout703 (.A(_0841_),
    .X(net703));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(_0625_));
 sg13g2_buf_4 fanout705 (.X(net705),
    .A(_0625_));
 sg13g2_buf_4 fanout706 (.X(net706),
    .A(_0624_));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(_0624_));
 sg13g2_buf_4 fanout708 (.X(net708),
    .A(_0623_));
 sg13g2_buf_2 fanout709 (.A(_0623_),
    .X(net709));
 sg13g2_buf_4 fanout710 (.X(net710),
    .A(_0622_));
 sg13g2_buf_2 fanout711 (.A(_0622_),
    .X(net711));
 sg13g2_buf_4 fanout712 (.X(net712),
    .A(_0617_));
 sg13g2_buf_4 fanout713 (.X(net713),
    .A(_0617_));
 sg13g2_buf_4 fanout714 (.X(net714),
    .A(_0616_));
 sg13g2_buf_2 fanout715 (.A(_0616_),
    .X(net715));
 sg13g2_buf_4 fanout716 (.X(net716),
    .A(_0613_));
 sg13g2_buf_4 fanout717 (.X(net717),
    .A(_0612_));
 sg13g2_buf_4 fanout718 (.X(net718),
    .A(_0612_));
 sg13g2_buf_4 fanout719 (.X(net719),
    .A(net723));
 sg13g2_buf_2 fanout720 (.A(net723),
    .X(net720));
 sg13g2_buf_4 fanout721 (.X(net721),
    .A(net722));
 sg13g2_buf_4 fanout722 (.X(net722),
    .A(net723));
 sg13g2_buf_4 fanout723 (.X(net723),
    .A(_0541_));
 sg13g2_buf_2 fanout724 (.A(net726),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(net726),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(_0524_),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(net728),
    .X(net727));
 sg13g2_buf_4 fanout728 (.X(net728),
    .A(_0524_));
 sg13g2_buf_2 fanout729 (.A(_1622_),
    .X(net729));
 sg13g2_buf_4 fanout730 (.X(net730),
    .A(_0848_));
 sg13g2_buf_2 fanout731 (.A(_0848_),
    .X(net731));
 sg13g2_buf_4 fanout732 (.X(net732),
    .A(_0847_));
 sg13g2_buf_4 fanout733 (.X(net733),
    .A(_0847_));
 sg13g2_buf_2 fanout734 (.A(_0614_),
    .X(net734));
 sg13g2_buf_4 fanout735 (.X(net735),
    .A(_0611_));
 sg13g2_buf_2 fanout736 (.A(_0610_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(_0610_),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_0607_),
    .X(net738));
 sg13g2_buf_4 fanout739 (.X(net739),
    .A(_0607_));
 sg13g2_buf_2 fanout740 (.A(net742),
    .X(net740));
 sg13g2_buf_1 fanout741 (.A(net742),
    .X(net741));
 sg13g2_buf_4 fanout742 (.X(net742),
    .A(_0606_));
 sg13g2_buf_4 fanout743 (.X(net743),
    .A(_0603_));
 sg13g2_buf_2 fanout744 (.A(_0602_),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(net749),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(net749),
    .X(net746));
 sg13g2_buf_4 fanout747 (.X(net747),
    .A(net748));
 sg13g2_buf_4 fanout748 (.X(net748),
    .A(net749));
 sg13g2_buf_2 fanout749 (.A(_0575_),
    .X(net749));
 sg13g2_buf_4 fanout750 (.X(net750),
    .A(net752));
 sg13g2_buf_1 fanout751 (.A(net752),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(_0558_),
    .X(net752));
 sg13g2_buf_4 fanout753 (.X(net753),
    .A(net754));
 sg13g2_buf_2 fanout754 (.A(_0558_),
    .X(net754));
 sg13g2_buf_4 fanout755 (.X(net755),
    .A(net756));
 sg13g2_buf_4 fanout756 (.X(net756),
    .A(net759));
 sg13g2_buf_2 fanout757 (.A(net758),
    .X(net757));
 sg13g2_buf_4 fanout758 (.X(net758),
    .A(net759));
 sg13g2_buf_2 fanout759 (.A(_0507_),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(net762),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(net762),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(_0490_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(net764),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(_0490_),
    .X(net764));
 sg13g2_buf_4 fanout765 (.X(net765),
    .A(net767));
 sg13g2_buf_2 fanout766 (.A(net767),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(_0472_),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(net769),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(_0472_),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(net771),
    .X(net770));
 sg13g2_buf_4 fanout771 (.X(net771),
    .A(net774));
 sg13g2_buf_4 fanout772 (.X(net772),
    .A(net773));
 sg13g2_buf_4 fanout773 (.X(net773),
    .A(net774));
 sg13g2_buf_4 fanout774 (.X(net774),
    .A(_0455_));
 sg13g2_buf_2 fanout775 (.A(_1273_),
    .X(net775));
 sg13g2_buf_4 fanout776 (.X(net776),
    .A(_0867_));
 sg13g2_buf_2 fanout777 (.A(_0866_),
    .X(net777));
 sg13g2_buf_1 fanout778 (.A(_0866_),
    .X(net778));
 sg13g2_buf_4 fanout779 (.X(net779),
    .A(net780));
 sg13g2_buf_2 fanout780 (.A(_0866_),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(_0029_),
    .X(net781));
 sg13g2_buf_4 fanout782 (.X(net782),
    .A(net783));
 sg13g2_buf_2 fanout783 (.A(net787),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(net787),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(net787),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(net787),
    .X(net786));
 sg13g2_buf_4 fanout787 (.X(net787),
    .A(_1597_));
 sg13g2_buf_2 fanout788 (.A(_1522_),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(_1520_),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(net791),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(net792),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(_1272_),
    .X(net792));
 sg13g2_buf_2 fanout793 (.A(_1596_),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(_1480_),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(_1475_),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(_1434_),
    .X(net796));
 sg13g2_buf_2 fanout797 (.A(net798),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(net800),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(net800),
    .X(net799));
 sg13g2_buf_4 fanout800 (.X(net800),
    .A(_1367_));
 sg13g2_buf_4 fanout801 (.X(net801),
    .A(net943));
 sg13g2_buf_4 fanout802 (.X(net802),
    .A(_0037_));
 sg13g2_buf_4 fanout803 (.X(net803),
    .A(_0038_));
 sg13g2_buf_4 fanout804 (.X(net804),
    .A(_0039_));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(_0040_));
 sg13g2_buf_4 fanout806 (.X(net806),
    .A(_0041_));
 sg13g2_buf_2 fanout807 (.A(net809),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(net809),
    .X(net808));
 sg13g2_buf_4 fanout809 (.X(net809),
    .A(net546));
 sg13g2_buf_2 fanout810 (.A(net811),
    .X(net810));
 sg13g2_buf_1 fanout811 (.A(net812),
    .X(net811));
 sg13g2_buf_1 fanout812 (.A(\cur_state[7] ),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(net814),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(net894),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(\uart_inst.T0.bit_counter[0] ),
    .X(net815));
 sg13g2_buf_1 fanout816 (.A(\uart_inst.T0.bit_counter[0] ),
    .X(net816));
 sg13g2_buf_4 fanout817 (.X(net817),
    .A(_1473_));
 sg13g2_buf_2 fanout818 (.A(_1469_),
    .X(net818));
 sg13g2_buf_4 fanout819 (.X(net819),
    .A(net822));
 sg13g2_buf_4 fanout820 (.X(net820),
    .A(net821));
 sg13g2_buf_4 fanout821 (.X(net821),
    .A(net822));
 sg13g2_buf_4 fanout822 (.X(net822),
    .A(_1439_));
 sg13g2_buf_2 fanout823 (.A(net824),
    .X(net823));
 sg13g2_buf_2 fanout824 (.A(ui_in[2]),
    .X(net824));
 sg13g2_buf_4 fanout825 (.X(net825),
    .A(net1));
 sg13g2_buf_2 fanout826 (.A(net827),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(ui_in[0]),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(net829),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(net830),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(net862),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(net832),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(net833),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(net862),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(net837),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(net837),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(net837),
    .X(net836));
 sg13g2_buf_1 fanout837 (.A(net844),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(net844),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(net844),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(net841),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(net842),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(net843),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(net844),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(net862),
    .X(net844));
 sg13g2_buf_4 fanout845 (.X(net845),
    .A(net846));
 sg13g2_buf_2 fanout846 (.A(net848),
    .X(net846));
 sg13g2_buf_4 fanout847 (.X(net847),
    .A(net848));
 sg13g2_buf_2 fanout848 (.A(net862),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(net850),
    .X(net849));
 sg13g2_buf_1 fanout850 (.A(net853),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(net853),
    .X(net851));
 sg13g2_buf_1 fanout852 (.A(net853),
    .X(net852));
 sg13g2_buf_4 fanout853 (.X(net853),
    .A(net862));
 sg13g2_buf_2 fanout854 (.A(net856),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(net856),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(net861),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(net861),
    .X(net857));
 sg13g2_buf_4 fanout858 (.X(net858),
    .A(net860));
 sg13g2_buf_2 fanout859 (.A(net860),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(net861),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(net862),
    .X(net861));
 sg13g2_buf_8 fanout862 (.A(rst_n),
    .X(net862));
 sg13g2_buf_2 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_tielo tt_um_bitty_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_33_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_20_clk));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_9_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_10_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_5_clk));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_19_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0070_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold2 (.A(\cur_state[4] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold3 (.A(\fi_inst.state[0] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold4 (.A(_1466_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0073_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0005_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold7 (.A(\bitty_inst.cpu_inst.d_inst[12] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold8 (.A(\bitty_inst.gen_dff[5].reg_out.mux_out[13] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0297_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold10 (.A(\cur_state[0] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0002_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold12 (.A(\bitty_inst.gen_dff[5].reg_out.mux_out[7] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0291_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold14 (.A(\bitty_inst.gen_dff[7].reg_out.mux_out[14] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0266_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold16 (.A(\bitty_inst.gen_dff[6].reg_out.mux_out[9] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0277_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold18 (.A(\bitty_inst.gen_dff[6].reg_out.mux_out[3] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0271_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold20 (.A(\bitty_inst.gen_dff[5].reg_out.mux_out[3] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0287_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold22 (.A(\bitty_inst.gen_dff[5].reg_out.mux_out[5] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0289_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold24 (.A(\bitty_inst.gen_dff[7].reg_out.mux_out[5] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0257_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold26 (.A(\bitty_inst.gen_dff[6].reg_out.mux_out[13] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0281_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold28 (.A(\bitty_inst.gen_dff[5].reg_out.mux_out[9] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0293_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold30 (.A(\bitty_inst.gen_dff[7].reg_out.mux_out[9] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0261_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold32 (.A(\bitty_inst.gen_dff[6].reg_out.mux_out[10] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0278_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold34 (.A(\bitty_inst.gen_dff[5].reg_out.mux_out[2] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0286_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold36 (.A(\bitty_inst.gen_dff[5].reg_out.mux_out[8] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0292_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold38 (.A(\bitty_inst.gen_dff[7].reg_out.mux_out[15] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0267_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold40 (.A(\bitty_inst.cpu_inst.d_inst[6] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold41 (.A(\bitty_inst.gen_dff[5].reg_out.mux_out[14] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0298_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold43 (.A(\bitty_inst.gen_dff[6].reg_out.mux_out[7] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0275_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold45 (.A(\bitty_inst.gen_dff[7].reg_out.mux_out[8] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0260_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold47 (.A(\bitty_inst.gen_dff[5].reg_out.mux_out[6] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0290_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold49 (.A(\bitty_inst.gen_dff[7].reg_out.mux_out[2] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0254_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold51 (.A(\bitty_inst.gen_dff[7].reg_out.mux_out[11] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0263_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold53 (.A(\bitty_inst.gen_dff[6].reg_out.mux_out[15] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0283_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold55 (.A(\bitty_inst.gen_dff[6].reg_out.mux_out[2] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0270_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold57 (.A(\bitty_inst.gen_dff[6].reg_out.mux_out[5] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0273_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold59 (.A(\bitty_inst.gen_dff[5].reg_out.mux_out[10] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0294_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold61 (.A(\bitty_inst.gen_dff[5].reg_out.mux_out[11] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0295_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold63 (.A(\bitty_inst.gen_dff[6].reg_out.mux_out[14] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0282_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold65 (.A(\bitty_inst.gen_dff[5].reg_out.mux_out[12] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0296_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold67 (.A(\bitty_inst.gen_dff[7].reg_out.mux_out[12] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0264_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold69 (.A(\bitty_inst.gen_dff[5].reg_out.mux_out[15] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0299_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold71 (.A(\bitty_inst.gen_dff[7].reg_out.mux_out[6] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0258_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold73 (.A(\bitty_inst.gen_dff[7].reg_out.mux_out[7] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0259_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold75 (.A(\bitty_inst.gen_dff[6].reg_out.mux_out[6] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0274_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold77 (.A(\bitty_inst.gen_dff[6].reg_out.mux_out[12] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0280_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold79 (.A(\bitty_inst.gen_dff[6].reg_out.mux_out[11] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0279_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold81 (.A(\bitty_inst.gen_dff[6].reg_out.mux_out[4] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0272_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold83 (.A(\bitty_inst.gen_dff[7].reg_out.mux_out[3] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0255_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold85 (.A(\bitty_inst.gen_dff[7].reg_out.mux_out[13] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0265_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold87 (.A(\bitty_inst.cpu_inst.d_inst[8] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0192_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold89 (.A(\bitty_inst.gen_dff[6].reg_out.mux_out[8] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0276_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold91 (.A(\bitty_inst.gen_dff[7].reg_out.mux_out[4] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0256_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold93 (.A(\bitty_inst.gen_dff[6].reg_out.mux_out[0] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0268_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold95 (.A(\bitty_inst.gen_dff[7].reg_out.mux_out[0] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0252_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold97 (.A(\uart_inst.T0.clk_counter[4] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold98 (.A(_1659_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold99 (.A(\bitty_inst.gen_dff[5].reg_out.mux_out[1] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0285_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold101 (.A(\bitty_inst.gen_dff[6].reg_out.mux_out[1] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0269_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold103 (.A(\uart_inst.T0.clk_counter[2] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold104 (.A(_1655_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0209_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold106 (.A(\uart_inst.T0.PS[4] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0027_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold108 (.A(\uart_inst.T0.clk_counter[6] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold109 (.A(_1663_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0213_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold111 (.A(\bitty_inst.gen_dff[7].reg_out.mux_out[1] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0253_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold113 (.A(\bitty_inst.gen_dff[5].reg_out.mux_out[4] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0288_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold115 (.A(\uart_inst.R0.clk_counter[4] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0379_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold117 (.A(\bitty_inst.gen_dff[5].reg_out.mux_out[0] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0284_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold119 (.A(\cur_state[3] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold120 (.A(_1463_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0012_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold122 (.A(\bitty_inst.gen_dff[7].reg_out.mux_out[10] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0262_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold124 (.A(\bitty_inst.cpu_inst.d_inst[10] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0194_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold126 (.A(\fi_inst.state[5] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold127 (.A(_1533_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0075_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold129 (.A(_1461_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold130 (.A(\uart_inst.R0.clk_counter[2] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0372_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold132 (.A(\cur_state[1] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold133 (.A(_1626_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold134 (.A(\bitty_inst.cpu_inst.d_inst[2] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold135 (.A(\bitty_inst.gen_dff[0].reg_out.mux_out[13] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0149_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold137 (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[12] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0084_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold139 (.A(\uart_inst.T0.clk_counter[8] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold140 (.A(_1667_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold141 (.A(\bitty_inst.gen_dff[1].reg_out.mux_out[15] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0135_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold143 (.A(\bitty_inst.cpu_inst.d_inst[11] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold144 (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[10] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0082_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold146 (.A(\uart_inst.R0.clk_counter[5] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0382_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold148 (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[14] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0086_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold150 (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[0] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0300_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold152 (.A(\bitty_inst.gen_dff[1].reg_out.mux_out[7] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0127_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold154 (.A(\bitty_inst.gen_dff[2].reg_out.mux_out[12] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0116_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold156 (.A(\uart_inst.T0.PS[0] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0024_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold158 (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[12] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0100_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold160 (.A(\bitty_inst.gen_dff[2].reg_out.mux_out[4] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0108_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold162 (.A(\bitty_inst.gen_dff[0].reg_out.mux_out[15] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0151_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold164 (.A(\bitty_inst.gen_dff[0].reg_out.mux_out[11] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0147_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold166 (.A(\bitty_inst.gen_dff[2].reg_out.mux_out[2] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0106_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold168 (.A(\bitty_inst.cpu_inst.cur_state[1] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold169 (.A(_1528_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0011_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold171 (.A(\bitty_inst.gen_dff[2].reg_out.mux_out[3] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0107_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold173 (.A(\bitty_inst.gen_dff[1].reg_out.mux_out[5] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0125_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold175 (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[15] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0087_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0055_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold178 (.A(\bitty_inst.gen_dff[0].reg_out.mux_out[7] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0143_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold180 (.A(\bitty_inst.gen_dff[1].reg_out.mux_out[3] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0123_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold182 (.A(\fi_inst.state[4] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold183 (.A(_1505_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold184 (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[3] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0303_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold186 (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[6] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0094_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold188 (.A(\bitty_inst.cpu_inst.run ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0008_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold190 (.A(\bitty_inst.gen_dff[0].reg_out.mux_out[6] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0142_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold192 (.A(\bitty_inst.gen_dff[2].reg_out.mux_out[13] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0117_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold194 (.A(\bitty_inst.gen_dff[1].reg_out.mux_out[6] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0126_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold196 (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[8] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0096_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold198 (.A(\bitty_inst.gen_dff[1].reg_out.mux_out[2] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0122_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold200 (.A(\bitty_inst.gen_dff[0].reg_out.mux_out[2] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0138_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold202 (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[15] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0103_),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold204 (.A(\bitty_inst.gen_dff[2].reg_out.mux_out[0] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0104_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold206 (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[2] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0302_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold208 (.A(\bitty_inst.gen_dff[0].reg_out.mux_out[1] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0137_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold210 (.A(\bitty_inst.gen_dff[2].reg_out.mux_out[10] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0114_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold212 (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[14] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0102_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold214 (.A(\bitty_inst.gen_dff[2].reg_out.mux_out[14] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0118_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold216 (.A(\bitty_inst.gen_dff[2].reg_out.mux_out[1] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0105_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0069_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold219 (.A(\bitty_inst.gen_dff[0].reg_out.mux_out[4] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0140_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold221 (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[2] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0090_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold223 (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[11] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0083_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold225 (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[13] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0085_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold227 (.A(\bitty_inst.gen_dff[0].reg_out.mux_out[3] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0139_),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold229 (.A(\bitty_inst.gen_dff[1].reg_out.mux_out[0] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0120_),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold231 (.A(\bitty_inst.cpu_inst.cur_state[2] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold232 (.A(\bitty_inst.gen_dff[2].reg_out.mux_out[15] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0119_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold234 (.A(\bitty_inst.gen_dff[1].reg_out.mux_out[10] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0130_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold236 (.A(\bitty_inst.gen_dff[1].reg_out.mux_out[14] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0134_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold238 (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[6] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0078_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold240 (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[10] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0098_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold242 (.A(\bitty_inst.gen_dff[1].reg_out.mux_out[13] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0133_),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold244 (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[9] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold245 (.A(\bitty_inst.gen_dff[2].reg_out.mux_out[5] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0109_),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold247 (.A(\bitty_inst.cpu_inst.d_inst[3] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold248 (.A(\bitty_inst.gen_dff[0].reg_out.mux_out[14] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0150_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold250 (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[4] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0092_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold252 (.A(\bitty_inst.gen_dff[2].reg_out.mux_out[11] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0115_),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold254 (.A(\uart_inst.T0.PS[2] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold255 (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[11] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0099_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold257 (.A(\bitty_inst.gen_dff[0].reg_out.mux_out[5] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0141_),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold259 (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[3] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0091_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold261 (.A(\bitty_inst.gen_dff[1].reg_out.mux_out[9] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold262 (.A(\bitty_inst.gen_dff[1].reg_out.mux_out[4] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0124_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold264 (.A(\bitty_inst.gen_dff[0].reg_out.mux_out[8] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0144_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold266 (.A(\uart_inst.R0.clk_counter[8] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0391_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold268 (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[8] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0080_),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold270 (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[7] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0079_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold272 (.A(\bitty_inst.gen_dff[1].reg_out.mux_out[8] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0128_),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold274 (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[5] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0077_),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold276 (.A(\bitty_inst.alu_inst.in_a[3] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold277 (.A(\bitty_inst.gen_dff[0].reg_out.mux_out[0] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0136_),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold279 (.A(\bitty_inst.gen_dff[0].reg_out.mux_out[12] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0148_),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold281 (.A(\uart_inst.R0.PS[0] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold282 (.A(_1586_),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold283 (.A(\bitty_inst.gen_dff[1].reg_out.mux_out[11] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0131_),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold285 (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[0] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0088_),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0064_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0362_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0228_),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold290 (.A(\bitty_inst.alu_inst.in_a[14] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold291 (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[1] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0089_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold293 (.A(\bitty_inst.gen_dff[2].reg_out.mux_out[9] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold294 (.A(\cur_state[7] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold295 (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[7] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0095_),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold297 (.A(\bitty_inst.gen_dff[2].reg_out.mux_out[6] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0110_),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold299 (.A(\bitty_inst.gen_dff[1].reg_out.mux_out[12] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0132_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold301 (.A(\bitty_inst.gen_dff[0].reg_out.mux_out[9] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold302 (.A(\uart_inst.R0.PS[5] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold303 (.A(\uart_inst.R0.clk_counter[9] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0393_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold305 (.A(\bitty_inst.gen_dff[0].reg_out.mux_out[10] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0146_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold307 (.A(\bitty_inst.cpu_inst.d_inst[5] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold308 (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[4] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0076_),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold310 (.A(\bitty_inst.gen_dff[2].reg_out.mux_out[8] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0112_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold312 (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[9] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold313 (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[5] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0093_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold315 (.A(\bitty_inst.cpu_inst.d_inst[7] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold316 (.A(\bitty_inst.gen_dff[2].reg_out.mux_out[7] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0111_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold318 (.A(\bitty_inst.gen_dff[1].reg_out.mux_out[1] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0121_),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold320 (.A(\uart_inst.R0.clk_counter[6] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0386_),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold322 (.A(_0066_),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold323 (.A(_1670_),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold324 (.A(\bitty_inst.cpu_inst.cur_state[0] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold325 (.A(_0009_),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold326 (.A(\bitty_inst.cpu_inst.d_inst[9] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold327 (.A(\bitty_inst.alu_inst.in_a[11] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold328 (.A(\uart_inst.R0.PS[3] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0243_),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold330 (.A(fetch_done),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold331 (.A(\bitty_inst.gen_dff[4].reg_out.mux_out[1] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0301_),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0071_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold334 (.A(_1651_),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0206_),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0065_),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold337 (.A(_1673_),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold338 (.A(_1674_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold339 (.A(\bitty_inst.alu_inst.in_a[10] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold340 (.A(\bitty_inst.alu_inst.in_a[1] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold341 (.A(\bitty_inst.alu_inst.in_a[13] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold342 (.A(\uart_inst.R0.clk_counter[7] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0235_),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold344 (.A(\bitty_inst.gen_dff[3].reg_out.mux_out[13] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0101_),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold346 (.A(\bitty_inst.alu_inst.in_a[8] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold347 (.A(\uart_inst.T0.clk_counter[0] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold348 (.A(_1653_),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold349 (.A(\uart_inst.R0.clk_counter[3] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold350 (.A(_0375_),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold351 (.A(\uart_inst.T0.clk_counter[10] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold352 (.A(_1672_),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold353 (.A(\bitty_inst.alu_inst.in_a[12] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold354 (.A(\uart_inst.T0.clk_counter[7] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold355 (.A(_1665_),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold356 (.A(\uart_inst.R0.bit_counter[0] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0403_),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold358 (.A(_0242_),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold359 (.A(\bitty_inst.alu_inst.in_a[6] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold360 (.A(\uart_inst.R0.PS[1] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold361 (.A(\uart_inst.T0.bit_counter[1] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold362 (.A(_1646_),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold363 (.A(_0205_),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold364 (.A(\uart_inst.T0.clk_counter[12] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold365 (.A(_1676_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold366 (.A(\bitty_inst.alu_inst.in_a[15] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold367 (.A(\bitty_inst.d_out[7] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold368 (.A(\cur_state[2] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold369 (.A(\addr[0] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0244_),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold371 (.A(\bitty_inst.d_out[15] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold372 (.A(\uart_inst.R0.clk_counter[1] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0368_),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold374 (.A(\bitty_inst.alu_inst.in_a[4] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold375 (.A(\bitty_inst.alu_inst.in_a[7] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold376 (.A(\bitty_inst.d_out[13] ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold377 (.A(\bitty_inst.cpu_inst.d_inst[13] ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold378 (.A(\bitty_inst.cpu_inst.d_inst[4] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold379 (.A(\bitty_inst.alu_inst.in_a[9] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold380 (.A(\uart_inst.R0.clk_counter[10] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold381 (.A(_0396_),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold382 (.A(\addr[1] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold383 (.A(\bitty_inst.alu_inst.in_a[0] ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold384 (.A(\uart_inst.R0.PS[2] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold385 (.A(_0324_),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold386 (.A(\uart_inst.T0.clk_counter[3] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold387 (.A(_1657_),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold388 (.A(\addr[2] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold389 (.A(\bitty_inst.alu_inst.in_a[5] ),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold390 (.A(\bitty_inst.cpu_inst.d_inst[14] ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold391 (.A(\uart_inst.T0.clk_counter[5] ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold392 (.A(_1661_),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold393 (.A(\bitty_inst.d_out[0] ),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold394 (.A(\uart_inst.T0.PS[1] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold395 (.A(_1644_),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0204_),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold397 (.A(\bitty_inst.alu_inst.in_a[2] ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold398 (.A(\bitty_inst.lsu_inst.rx_data[2] ),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0222_),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold400 (.A(\addr[4] ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0248_),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold402 (.A(\bitty_inst.lsu_inst.rx_data[1] ),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold403 (.A(_0221_),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold404 (.A(\addr[5] ),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold405 (.A(_0249_),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold406 (.A(\addr[7] ),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0251_),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold408 (.A(\uart_inst.T0.PS[1] ),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold409 (.A(\bitty_inst.d_out[5] ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0065_),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold411 (.A(\addr[6] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0250_),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold413 (.A(\bitty_inst.d_out[3] ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold414 (.A(\bitty_inst.cpu_inst.d_inst[0] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold415 (.A(\bitty_inst.d_out[9] ),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold416 (.A(\addr[3] ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold417 (.A(\bitty_inst.cpu_inst.d_inst[1] ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold418 (.A(\bitty_inst.lsu_inst.rx_data[6] ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold419 (.A(\bitty_inst.lsu_inst.rx_data[4] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold420 (.A(_0224_),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold421 (.A(\bitty_inst.d_out[10] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold422 (.A(\uart_inst.R0.PS[1] ),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0241_),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold424 (.A(\bitty_inst.d_out[4] ),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold425 (.A(\bitty_inst.d_out[12] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold426 (.A(\bitty_inst.d_out[1] ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold427 (.A(\bitty_inst.lsu_inst.rx_data[3] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold428 (.A(\bitty_inst.d_out[11] ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold429 (.A(\uart_inst.R0.clk_counter[11] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0239_),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold431 (.A(\bitty_inst.d_out[14] ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold432 (.A(\bitty_inst.lsu_inst.rx_data[7] ),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold433 (.A(\bitty_inst.lsu_inst.rx_data[5] ),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold434 (.A(\bitty_inst.d_out[8] ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold435 (.A(\bitty_inst.d_out[2] ),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold436 (.A(\bitty_inst.cpu_inst.d_inst[15] ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold437 (.A(\bitty_inst.d_out[6] ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold438 (.A(\uart_inst.T0.clk_counter[3] ),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold439 (.A(\uart_inst.R0.clk_counter[10] ),
    .X(net965));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_fill_1 FILLER_0_245 ();
 sg13g2_fill_1 FILLER_0_312 ();
 sg13g2_fill_1 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_365 ();
 sg13g2_decap_8 FILLER_0_372 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_4 FILLER_1_231 ();
 sg13g2_fill_2 FILLER_1_296 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_4 FILLER_2_210 ();
 sg13g2_fill_2 FILLER_2_214 ();
 sg13g2_fill_1 FILLER_2_294 ();
 sg13g2_fill_2 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_4 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_4 FILLER_3_210 ();
 sg13g2_fill_1 FILLER_3_214 ();
 sg13g2_fill_1 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_362 ();
 sg13g2_decap_8 FILLER_3_369 ();
 sg13g2_decap_8 FILLER_3_376 ();
 sg13g2_decap_8 FILLER_3_383 ();
 sg13g2_decap_8 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_207 ();
 sg13g2_fill_1 FILLER_4_214 ();
 sg13g2_fill_1 FILLER_4_238 ();
 sg13g2_fill_1 FILLER_4_275 ();
 sg13g2_fill_1 FILLER_4_291 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_4 FILLER_4_403 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_fill_2 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_171 ();
 sg13g2_decap_4 FILLER_5_178 ();
 sg13g2_fill_1 FILLER_5_182 ();
 sg13g2_fill_2 FILLER_5_187 ();
 sg13g2_fill_1 FILLER_5_218 ();
 sg13g2_fill_1 FILLER_5_273 ();
 sg13g2_fill_1 FILLER_5_304 ();
 sg13g2_decap_8 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_374 ();
 sg13g2_decap_8 FILLER_5_381 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_4 FILLER_6_140 ();
 sg13g2_fill_1 FILLER_6_144 ();
 sg13g2_fill_2 FILLER_6_183 ();
 sg13g2_fill_2 FILLER_6_208 ();
 sg13g2_fill_2 FILLER_6_227 ();
 sg13g2_fill_1 FILLER_6_243 ();
 sg13g2_fill_1 FILLER_6_294 ();
 sg13g2_fill_2 FILLER_6_309 ();
 sg13g2_decap_8 FILLER_6_377 ();
 sg13g2_decap_8 FILLER_6_384 ();
 sg13g2_decap_8 FILLER_6_391 ();
 sg13g2_decap_8 FILLER_6_398 ();
 sg13g2_decap_4 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_fill_2 FILLER_7_133 ();
 sg13g2_fill_1 FILLER_7_161 ();
 sg13g2_fill_2 FILLER_7_192 ();
 sg13g2_fill_2 FILLER_7_253 ();
 sg13g2_fill_1 FILLER_7_270 ();
 sg13g2_fill_1 FILLER_7_302 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_fill_1 FILLER_9_192 ();
 sg13g2_fill_2 FILLER_9_211 ();
 sg13g2_fill_1 FILLER_9_213 ();
 sg13g2_fill_2 FILLER_9_230 ();
 sg13g2_fill_1 FILLER_9_232 ();
 sg13g2_fill_1 FILLER_9_251 ();
 sg13g2_decap_8 FILLER_9_380 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_fill_2 FILLER_10_112 ();
 sg13g2_fill_2 FILLER_10_238 ();
 sg13g2_fill_1 FILLER_10_240 ();
 sg13g2_fill_1 FILLER_10_256 ();
 sg13g2_fill_2 FILLER_10_288 ();
 sg13g2_fill_1 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_381 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_395 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_fill_2 FILLER_11_105 ();
 sg13g2_fill_1 FILLER_11_107 ();
 sg13g2_fill_2 FILLER_11_126 ();
 sg13g2_fill_1 FILLER_11_128 ();
 sg13g2_fill_1 FILLER_11_185 ();
 sg13g2_fill_2 FILLER_11_206 ();
 sg13g2_decap_4 FILLER_11_232 ();
 sg13g2_fill_2 FILLER_11_236 ();
 sg13g2_fill_1 FILLER_11_300 ();
 sg13g2_fill_2 FILLER_11_306 ();
 sg13g2_fill_1 FILLER_11_334 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_fill_1 FILLER_12_112 ();
 sg13g2_fill_2 FILLER_12_125 ();
 sg13g2_fill_2 FILLER_12_179 ();
 sg13g2_fill_2 FILLER_12_191 ();
 sg13g2_fill_1 FILLER_12_193 ();
 sg13g2_fill_2 FILLER_12_244 ();
 sg13g2_fill_2 FILLER_12_277 ();
 sg13g2_fill_2 FILLER_12_315 ();
 sg13g2_fill_2 FILLER_12_348 ();
 sg13g2_fill_1 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_4 FILLER_13_119 ();
 sg13g2_fill_2 FILLER_13_123 ();
 sg13g2_fill_1 FILLER_13_133 ();
 sg13g2_fill_2 FILLER_13_241 ();
 sg13g2_fill_1 FILLER_13_309 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_4 FILLER_14_140 ();
 sg13g2_fill_1 FILLER_14_144 ();
 sg13g2_fill_1 FILLER_14_153 ();
 sg13g2_fill_2 FILLER_14_187 ();
 sg13g2_fill_1 FILLER_14_189 ();
 sg13g2_fill_1 FILLER_14_205 ();
 sg13g2_decap_4 FILLER_14_214 ();
 sg13g2_decap_4 FILLER_14_227 ();
 sg13g2_fill_2 FILLER_14_231 ();
 sg13g2_decap_4 FILLER_14_242 ();
 sg13g2_fill_2 FILLER_14_246 ();
 sg13g2_fill_1 FILLER_14_264 ();
 sg13g2_fill_2 FILLER_14_286 ();
 sg13g2_fill_1 FILLER_14_324 ();
 sg13g2_fill_2 FILLER_14_346 ();
 sg13g2_decap_8 FILLER_14_393 ();
 sg13g2_decap_8 FILLER_14_400 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_4 FILLER_15_133 ();
 sg13g2_fill_2 FILLER_15_137 ();
 sg13g2_decap_4 FILLER_15_170 ();
 sg13g2_fill_1 FILLER_15_174 ();
 sg13g2_decap_4 FILLER_15_191 ();
 sg13g2_decap_4 FILLER_15_221 ();
 sg13g2_fill_2 FILLER_15_225 ();
 sg13g2_fill_2 FILLER_15_236 ();
 sg13g2_fill_1 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_264 ();
 sg13g2_decap_4 FILLER_15_271 ();
 sg13g2_fill_1 FILLER_15_282 ();
 sg13g2_fill_1 FILLER_15_301 ();
 sg13g2_fill_2 FILLER_15_307 ();
 sg13g2_fill_1 FILLER_15_314 ();
 sg13g2_fill_2 FILLER_15_330 ();
 sg13g2_fill_1 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_4 FILLER_16_119 ();
 sg13g2_fill_1 FILLER_16_123 ();
 sg13g2_decap_4 FILLER_16_160 ();
 sg13g2_fill_1 FILLER_16_164 ();
 sg13g2_fill_1 FILLER_16_174 ();
 sg13g2_fill_1 FILLER_16_191 ();
 sg13g2_decap_4 FILLER_16_201 ();
 sg13g2_fill_2 FILLER_16_224 ();
 sg13g2_fill_1 FILLER_16_226 ();
 sg13g2_fill_2 FILLER_16_239 ();
 sg13g2_fill_1 FILLER_16_280 ();
 sg13g2_fill_1 FILLER_16_286 ();
 sg13g2_fill_2 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_decap_8 FILLER_16_397 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_4 FILLER_17_105 ();
 sg13g2_fill_1 FILLER_17_109 ();
 sg13g2_decap_4 FILLER_17_150 ();
 sg13g2_fill_2 FILLER_17_154 ();
 sg13g2_fill_1 FILLER_17_187 ();
 sg13g2_fill_2 FILLER_17_206 ();
 sg13g2_fill_1 FILLER_17_213 ();
 sg13g2_fill_2 FILLER_17_226 ();
 sg13g2_fill_1 FILLER_17_228 ();
 sg13g2_fill_2 FILLER_17_257 ();
 sg13g2_fill_2 FILLER_17_302 ();
 sg13g2_fill_1 FILLER_17_304 ();
 sg13g2_fill_1 FILLER_17_335 ();
 sg13g2_fill_2 FILLER_17_364 ();
 sg13g2_fill_1 FILLER_17_366 ();
 sg13g2_decap_8 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_fill_2 FILLER_18_112 ();
 sg13g2_decap_4 FILLER_18_137 ();
 sg13g2_fill_2 FILLER_18_141 ();
 sg13g2_fill_2 FILLER_18_149 ();
 sg13g2_fill_1 FILLER_18_151 ();
 sg13g2_fill_2 FILLER_18_161 ();
 sg13g2_fill_2 FILLER_18_198 ();
 sg13g2_fill_2 FILLER_18_205 ();
 sg13g2_fill_1 FILLER_18_207 ();
 sg13g2_fill_1 FILLER_18_276 ();
 sg13g2_fill_1 FILLER_18_309 ();
 sg13g2_fill_2 FILLER_18_320 ();
 sg13g2_fill_1 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_fill_2 FILLER_19_119 ();
 sg13g2_fill_1 FILLER_19_121 ();
 sg13g2_fill_2 FILLER_19_144 ();
 sg13g2_fill_2 FILLER_19_198 ();
 sg13g2_fill_2 FILLER_19_226 ();
 sg13g2_fill_1 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_305 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_4 FILLER_20_112 ();
 sg13g2_fill_1 FILLER_20_116 ();
 sg13g2_fill_1 FILLER_20_133 ();
 sg13g2_fill_1 FILLER_20_191 ();
 sg13g2_decap_8 FILLER_20_220 ();
 sg13g2_fill_2 FILLER_20_227 ();
 sg13g2_fill_1 FILLER_20_229 ();
 sg13g2_fill_2 FILLER_20_244 ();
 sg13g2_fill_1 FILLER_20_246 ();
 sg13g2_fill_2 FILLER_20_269 ();
 sg13g2_fill_1 FILLER_20_301 ();
 sg13g2_fill_2 FILLER_20_306 ();
 sg13g2_fill_2 FILLER_20_339 ();
 sg13g2_fill_2 FILLER_20_348 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_4 FILLER_21_105 ();
 sg13g2_fill_2 FILLER_21_176 ();
 sg13g2_fill_1 FILLER_21_178 ();
 sg13g2_fill_2 FILLER_21_184 ();
 sg13g2_fill_1 FILLER_21_186 ();
 sg13g2_fill_1 FILLER_21_208 ();
 sg13g2_decap_8 FILLER_21_213 ();
 sg13g2_fill_1 FILLER_21_220 ();
 sg13g2_fill_1 FILLER_21_309 ();
 sg13g2_fill_1 FILLER_21_320 ();
 sg13g2_fill_1 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_112 ();
 sg13g2_fill_2 FILLER_22_131 ();
 sg13g2_fill_2 FILLER_22_141 ();
 sg13g2_fill_1 FILLER_22_183 ();
 sg13g2_fill_2 FILLER_22_188 ();
 sg13g2_fill_1 FILLER_22_195 ();
 sg13g2_fill_2 FILLER_22_204 ();
 sg13g2_fill_1 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_219 ();
 sg13g2_decap_4 FILLER_22_230 ();
 sg13g2_fill_1 FILLER_22_256 ();
 sg13g2_fill_1 FILLER_22_301 ();
 sg13g2_fill_2 FILLER_22_331 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_4 FILLER_23_105 ();
 sg13g2_fill_1 FILLER_23_109 ();
 sg13g2_fill_2 FILLER_23_166 ();
 sg13g2_fill_1 FILLER_23_168 ();
 sg13g2_fill_2 FILLER_23_185 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_fill_2 FILLER_23_240 ();
 sg13g2_fill_1 FILLER_23_242 ();
 sg13g2_fill_2 FILLER_23_281 ();
 sg13g2_fill_2 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_fill_2 FILLER_24_158 ();
 sg13g2_fill_2 FILLER_24_165 ();
 sg13g2_fill_2 FILLER_24_254 ();
 sg13g2_fill_1 FILLER_24_256 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_fill_2 FILLER_25_128 ();
 sg13g2_fill_1 FILLER_25_130 ();
 sg13g2_fill_2 FILLER_25_165 ();
 sg13g2_decap_8 FILLER_25_172 ();
 sg13g2_fill_2 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_181 ();
 sg13g2_decap_8 FILLER_25_225 ();
 sg13g2_decap_4 FILLER_25_232 ();
 sg13g2_fill_2 FILLER_25_236 ();
 sg13g2_fill_2 FILLER_25_242 ();
 sg13g2_fill_1 FILLER_25_244 ();
 sg13g2_fill_2 FILLER_25_249 ();
 sg13g2_fill_1 FILLER_25_251 ();
 sg13g2_fill_1 FILLER_25_258 ();
 sg13g2_fill_2 FILLER_25_282 ();
 sg13g2_fill_2 FILLER_25_306 ();
 sg13g2_fill_2 FILLER_25_313 ();
 sg13g2_fill_1 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_fill_2 FILLER_26_119 ();
 sg13g2_fill_1 FILLER_26_121 ();
 sg13g2_decap_4 FILLER_26_161 ();
 sg13g2_fill_2 FILLER_26_186 ();
 sg13g2_fill_1 FILLER_26_196 ();
 sg13g2_fill_1 FILLER_26_201 ();
 sg13g2_decap_4 FILLER_26_205 ();
 sg13g2_fill_2 FILLER_26_217 ();
 sg13g2_fill_1 FILLER_26_219 ();
 sg13g2_decap_4 FILLER_26_255 ();
 sg13g2_fill_1 FILLER_26_295 ();
 sg13g2_fill_1 FILLER_26_326 ();
 sg13g2_fill_2 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_4 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_116 ();
 sg13g2_fill_1 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_202 ();
 sg13g2_fill_1 FILLER_27_209 ();
 sg13g2_decap_4 FILLER_27_213 ();
 sg13g2_decap_4 FILLER_27_222 ();
 sg13g2_fill_1 FILLER_27_226 ();
 sg13g2_fill_1 FILLER_27_236 ();
 sg13g2_decap_8 FILLER_27_241 ();
 sg13g2_decap_8 FILLER_27_248 ();
 sg13g2_fill_1 FILLER_27_255 ();
 sg13g2_fill_1 FILLER_27_277 ();
 sg13g2_fill_2 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_397 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_4 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_102 ();
 sg13g2_fill_2 FILLER_28_171 ();
 sg13g2_fill_1 FILLER_28_209 ();
 sg13g2_fill_2 FILLER_28_223 ();
 sg13g2_fill_1 FILLER_28_225 ();
 sg13g2_fill_2 FILLER_28_309 ();
 sg13g2_fill_1 FILLER_28_354 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_fill_2 FILLER_29_91 ();
 sg13g2_fill_1 FILLER_29_93 ();
 sg13g2_fill_2 FILLER_29_124 ();
 sg13g2_fill_1 FILLER_29_145 ();
 sg13g2_fill_2 FILLER_29_151 ();
 sg13g2_decap_4 FILLER_29_172 ();
 sg13g2_fill_1 FILLER_29_176 ();
 sg13g2_fill_1 FILLER_29_185 ();
 sg13g2_fill_2 FILLER_29_206 ();
 sg13g2_fill_1 FILLER_29_231 ();
 sg13g2_decap_4 FILLER_29_258 ();
 sg13g2_fill_2 FILLER_29_262 ();
 sg13g2_fill_1 FILLER_29_319 ();
 sg13g2_fill_1 FILLER_29_325 ();
 sg13g2_fill_1 FILLER_29_352 ();
 sg13g2_decap_8 FILLER_29_391 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_152 ();
 sg13g2_decap_4 FILLER_30_159 ();
 sg13g2_fill_1 FILLER_30_163 ();
 sg13g2_decap_4 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_208 ();
 sg13g2_decap_4 FILLER_30_222 ();
 sg13g2_fill_2 FILLER_30_234 ();
 sg13g2_fill_1 FILLER_30_236 ();
 sg13g2_fill_2 FILLER_30_358 ();
 sg13g2_decap_8 FILLER_30_394 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_fill_2 FILLER_31_84 ();
 sg13g2_fill_2 FILLER_31_108 ();
 sg13g2_decap_8 FILLER_31_143 ();
 sg13g2_fill_2 FILLER_31_157 ();
 sg13g2_decap_4 FILLER_31_172 ();
 sg13g2_fill_1 FILLER_31_176 ();
 sg13g2_decap_8 FILLER_31_181 ();
 sg13g2_decap_8 FILLER_31_188 ();
 sg13g2_decap_8 FILLER_31_195 ();
 sg13g2_decap_4 FILLER_31_202 ();
 sg13g2_fill_2 FILLER_31_206 ();
 sg13g2_fill_2 FILLER_31_212 ();
 sg13g2_fill_2 FILLER_31_219 ();
 sg13g2_decap_8 FILLER_31_232 ();
 sg13g2_decap_8 FILLER_31_239 ();
 sg13g2_decap_8 FILLER_31_246 ();
 sg13g2_decap_4 FILLER_31_253 ();
 sg13g2_fill_1 FILLER_31_257 ();
 sg13g2_fill_1 FILLER_31_270 ();
 sg13g2_fill_2 FILLER_31_358 ();
 sg13g2_decap_8 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_fill_2 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_118 ();
 sg13g2_fill_2 FILLER_32_192 ();
 sg13g2_fill_2 FILLER_32_207 ();
 sg13g2_fill_2 FILLER_32_228 ();
 sg13g2_fill_2 FILLER_32_256 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_fill_2 FILLER_32_268 ();
 sg13g2_fill_1 FILLER_32_353 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_fill_1 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_141 ();
 sg13g2_decap_8 FILLER_33_199 ();
 sg13g2_fill_1 FILLER_33_206 ();
 sg13g2_decap_8 FILLER_33_220 ();
 sg13g2_fill_2 FILLER_33_253 ();
 sg13g2_fill_1 FILLER_33_255 ();
 sg13g2_fill_1 FILLER_33_327 ();
 sg13g2_fill_1 FILLER_33_372 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_fill_2 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_106 ();
 sg13g2_fill_2 FILLER_34_150 ();
 sg13g2_fill_2 FILLER_34_267 ();
 sg13g2_fill_2 FILLER_34_278 ();
 sg13g2_fill_1 FILLER_34_280 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_91 ();
 sg13g2_fill_2 FILLER_35_109 ();
 sg13g2_fill_2 FILLER_35_144 ();
 sg13g2_fill_1 FILLER_35_146 ();
 sg13g2_fill_2 FILLER_35_188 ();
 sg13g2_fill_1 FILLER_35_190 ();
 sg13g2_fill_2 FILLER_35_218 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_fill_1 FILLER_35_238 ();
 sg13g2_fill_2 FILLER_35_271 ();
 sg13g2_fill_1 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_284 ();
 sg13g2_fill_2 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_351 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_fill_2 FILLER_36_98 ();
 sg13g2_fill_1 FILLER_36_100 ();
 sg13g2_fill_1 FILLER_36_127 ();
 sg13g2_fill_2 FILLER_36_155 ();
 sg13g2_decap_4 FILLER_36_166 ();
 sg13g2_fill_2 FILLER_36_170 ();
 sg13g2_decap_4 FILLER_36_180 ();
 sg13g2_decap_8 FILLER_36_228 ();
 sg13g2_fill_1 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_244 ();
 sg13g2_fill_2 FILLER_36_250 ();
 sg13g2_decap_8 FILLER_36_271 ();
 sg13g2_decap_8 FILLER_36_278 ();
 sg13g2_fill_2 FILLER_36_313 ();
 sg13g2_fill_2 FILLER_36_324 ();
 sg13g2_fill_1 FILLER_36_375 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_fill_2 FILLER_37_105 ();
 sg13g2_fill_1 FILLER_37_124 ();
 sg13g2_decap_8 FILLER_37_151 ();
 sg13g2_decap_8 FILLER_37_158 ();
 sg13g2_decap_8 FILLER_37_165 ();
 sg13g2_decap_8 FILLER_37_172 ();
 sg13g2_decap_4 FILLER_37_179 ();
 sg13g2_decap_4 FILLER_37_186 ();
 sg13g2_fill_1 FILLER_37_190 ();
 sg13g2_decap_4 FILLER_37_194 ();
 sg13g2_fill_1 FILLER_37_198 ();
 sg13g2_fill_1 FILLER_37_213 ();
 sg13g2_fill_2 FILLER_37_228 ();
 sg13g2_fill_1 FILLER_37_230 ();
 sg13g2_fill_2 FILLER_37_235 ();
 sg13g2_fill_2 FILLER_37_258 ();
 sg13g2_decap_4 FILLER_37_282 ();
 sg13g2_fill_1 FILLER_37_286 ();
 sg13g2_fill_2 FILLER_37_292 ();
 sg13g2_fill_2 FILLER_37_302 ();
 sg13g2_fill_1 FILLER_37_383 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_91 ();
 sg13g2_fill_1 FILLER_38_93 ();
 sg13g2_fill_2 FILLER_38_125 ();
 sg13g2_decap_8 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_143 ();
 sg13g2_fill_1 FILLER_38_147 ();
 sg13g2_fill_2 FILLER_38_160 ();
 sg13g2_fill_1 FILLER_38_162 ();
 sg13g2_fill_2 FILLER_38_183 ();
 sg13g2_fill_2 FILLER_38_189 ();
 sg13g2_decap_4 FILLER_38_201 ();
 sg13g2_fill_2 FILLER_38_205 ();
 sg13g2_decap_8 FILLER_38_221 ();
 sg13g2_fill_2 FILLER_38_228 ();
 sg13g2_decap_8 FILLER_38_284 ();
 sg13g2_decap_4 FILLER_38_291 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_decap_4 FILLER_38_330 ();
 sg13g2_fill_2 FILLER_38_334 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_decap_4 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_fill_1 FILLER_39_91 ();
 sg13g2_fill_2 FILLER_39_108 ();
 sg13g2_decap_8 FILLER_39_118 ();
 sg13g2_decap_4 FILLER_39_125 ();
 sg13g2_fill_1 FILLER_39_129 ();
 sg13g2_decap_4 FILLER_39_154 ();
 sg13g2_fill_1 FILLER_39_158 ();
 sg13g2_fill_2 FILLER_39_207 ();
 sg13g2_fill_1 FILLER_39_209 ();
 sg13g2_fill_1 FILLER_39_232 ();
 sg13g2_fill_1 FILLER_39_239 ();
 sg13g2_fill_2 FILLER_39_249 ();
 sg13g2_fill_2 FILLER_39_256 ();
 sg13g2_fill_2 FILLER_39_268 ();
 sg13g2_fill_1 FILLER_39_270 ();
 sg13g2_decap_8 FILLER_39_309 ();
 sg13g2_decap_4 FILLER_39_316 ();
 sg13g2_fill_2 FILLER_39_320 ();
 sg13g2_decap_8 FILLER_39_330 ();
 sg13g2_decap_4 FILLER_39_337 ();
 sg13g2_fill_2 FILLER_39_341 ();
 sg13g2_decap_8 FILLER_39_402 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_fill_1 FILLER_40_107 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_fill_1 FILLER_40_119 ();
 sg13g2_decap_4 FILLER_40_158 ();
 sg13g2_fill_2 FILLER_40_207 ();
 sg13g2_decap_8 FILLER_40_234 ();
 sg13g2_decap_8 FILLER_40_241 ();
 sg13g2_decap_8 FILLER_40_248 ();
 sg13g2_decap_4 FILLER_40_255 ();
 sg13g2_fill_2 FILLER_40_319 ();
 sg13g2_fill_1 FILLER_40_337 ();
 sg13g2_decap_4 FILLER_40_346 ();
 sg13g2_fill_2 FILLER_40_350 ();
 sg13g2_fill_1 FILLER_40_360 ();
 sg13g2_fill_2 FILLER_40_367 ();
 sg13g2_decap_4 FILLER_40_404 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_fill_2 FILLER_41_108 ();
 sg13g2_fill_1 FILLER_41_110 ();
 sg13g2_fill_1 FILLER_41_158 ();
 sg13g2_fill_1 FILLER_41_178 ();
 sg13g2_decap_8 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_230 ();
 sg13g2_fill_1 FILLER_41_237 ();
 sg13g2_decap_4 FILLER_41_258 ();
 sg13g2_fill_2 FILLER_41_268 ();
 sg13g2_fill_1 FILLER_41_270 ();
 sg13g2_decap_4 FILLER_41_289 ();
 sg13g2_fill_2 FILLER_41_293 ();
 sg13g2_fill_2 FILLER_41_308 ();
 sg13g2_fill_1 FILLER_41_310 ();
 sg13g2_fill_2 FILLER_41_335 ();
 sg13g2_fill_1 FILLER_41_363 ();
 sg13g2_decap_4 FILLER_41_369 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_fill_2 FILLER_41_406 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_4 FILLER_42_77 ();
 sg13g2_fill_2 FILLER_42_81 ();
 sg13g2_fill_2 FILLER_42_129 ();
 sg13g2_fill_1 FILLER_42_131 ();
 sg13g2_fill_1 FILLER_42_152 ();
 sg13g2_fill_2 FILLER_42_168 ();
 sg13g2_fill_1 FILLER_42_170 ();
 sg13g2_fill_2 FILLER_42_186 ();
 sg13g2_decap_8 FILLER_42_193 ();
 sg13g2_decap_8 FILLER_42_200 ();
 sg13g2_decap_8 FILLER_42_207 ();
 sg13g2_decap_4 FILLER_42_214 ();
 sg13g2_decap_8 FILLER_42_222 ();
 sg13g2_fill_1 FILLER_42_229 ();
 sg13g2_decap_4 FILLER_42_258 ();
 sg13g2_fill_2 FILLER_42_262 ();
 sg13g2_decap_8 FILLER_42_272 ();
 sg13g2_decap_4 FILLER_42_279 ();
 sg13g2_decap_8 FILLER_42_288 ();
 sg13g2_decap_4 FILLER_42_295 ();
 sg13g2_decap_8 FILLER_42_304 ();
 sg13g2_decap_8 FILLER_42_324 ();
 sg13g2_fill_2 FILLER_42_331 ();
 sg13g2_fill_2 FILLER_42_351 ();
 sg13g2_fill_1 FILLER_42_353 ();
 sg13g2_fill_2 FILLER_42_369 ();
 sg13g2_fill_1 FILLER_42_371 ();
 sg13g2_fill_1 FILLER_42_381 ();
 sg13g2_decap_8 FILLER_42_395 ();
 sg13g2_decap_8 FILLER_42_402 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_fill_2 FILLER_43_70 ();
 sg13g2_fill_1 FILLER_43_72 ();
 sg13g2_fill_1 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_83 ();
 sg13g2_decap_8 FILLER_43_90 ();
 sg13g2_decap_4 FILLER_43_97 ();
 sg13g2_fill_2 FILLER_43_101 ();
 sg13g2_fill_1 FILLER_43_112 ();
 sg13g2_fill_1 FILLER_43_117 ();
 sg13g2_fill_2 FILLER_43_161 ();
 sg13g2_fill_1 FILLER_43_163 ();
 sg13g2_decap_8 FILLER_43_184 ();
 sg13g2_decap_4 FILLER_43_191 ();
 sg13g2_fill_1 FILLER_43_195 ();
 sg13g2_fill_1 FILLER_43_201 ();
 sg13g2_fill_2 FILLER_43_219 ();
 sg13g2_fill_2 FILLER_43_251 ();
 sg13g2_decap_4 FILLER_43_269 ();
 sg13g2_decap_4 FILLER_43_277 ();
 sg13g2_fill_2 FILLER_43_281 ();
 sg13g2_decap_8 FILLER_43_287 ();
 sg13g2_decap_8 FILLER_43_294 ();
 sg13g2_fill_2 FILLER_43_301 ();
 sg13g2_fill_1 FILLER_43_343 ();
 sg13g2_decap_4 FILLER_43_405 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_94 ();
 sg13g2_fill_1 FILLER_44_101 ();
 sg13g2_fill_1 FILLER_44_150 ();
 sg13g2_decap_4 FILLER_44_156 ();
 sg13g2_decap_8 FILLER_44_163 ();
 sg13g2_fill_2 FILLER_44_170 ();
 sg13g2_decap_4 FILLER_44_182 ();
 sg13g2_fill_1 FILLER_44_204 ();
 sg13g2_decap_4 FILLER_44_215 ();
 sg13g2_fill_2 FILLER_44_219 ();
 sg13g2_decap_4 FILLER_44_225 ();
 sg13g2_fill_2 FILLER_44_229 ();
 sg13g2_fill_2 FILLER_44_241 ();
 sg13g2_decap_8 FILLER_44_257 ();
 sg13g2_decap_8 FILLER_44_288 ();
 sg13g2_fill_2 FILLER_44_295 ();
 sg13g2_fill_1 FILLER_44_297 ();
 sg13g2_fill_1 FILLER_44_358 ();
 sg13g2_fill_1 FILLER_44_374 ();
 sg13g2_decap_8 FILLER_44_401 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_fill_1 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_100 ();
 sg13g2_decap_8 FILLER_45_107 ();
 sg13g2_decap_8 FILLER_45_114 ();
 sg13g2_decap_8 FILLER_45_121 ();
 sg13g2_decap_8 FILLER_45_128 ();
 sg13g2_decap_4 FILLER_45_135 ();
 sg13g2_fill_1 FILLER_45_139 ();
 sg13g2_decap_4 FILLER_45_149 ();
 sg13g2_fill_1 FILLER_45_153 ();
 sg13g2_decap_8 FILLER_45_163 ();
 sg13g2_fill_1 FILLER_45_170 ();
 sg13g2_fill_2 FILLER_45_177 ();
 sg13g2_fill_2 FILLER_45_197 ();
 sg13g2_decap_4 FILLER_45_231 ();
 sg13g2_fill_1 FILLER_45_235 ();
 sg13g2_decap_8 FILLER_45_248 ();
 sg13g2_fill_1 FILLER_45_255 ();
 sg13g2_decap_4 FILLER_45_288 ();
 sg13g2_fill_1 FILLER_45_292 ();
 sg13g2_decap_4 FILLER_45_301 ();
 sg13g2_fill_2 FILLER_45_314 ();
 sg13g2_fill_1 FILLER_45_364 ();
 sg13g2_decap_8 FILLER_45_401 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_fill_1 FILLER_46_70 ();
 sg13g2_fill_2 FILLER_46_107 ();
 sg13g2_decap_8 FILLER_46_113 ();
 sg13g2_decap_8 FILLER_46_120 ();
 sg13g2_decap_8 FILLER_46_127 ();
 sg13g2_fill_1 FILLER_46_138 ();
 sg13g2_fill_2 FILLER_46_144 ();
 sg13g2_fill_1 FILLER_46_146 ();
 sg13g2_fill_2 FILLER_46_180 ();
 sg13g2_fill_1 FILLER_46_182 ();
 sg13g2_fill_2 FILLER_46_195 ();
 sg13g2_decap_8 FILLER_46_212 ();
 sg13g2_decap_4 FILLER_46_219 ();
 sg13g2_fill_2 FILLER_46_223 ();
 sg13g2_decap_4 FILLER_46_234 ();
 sg13g2_fill_2 FILLER_46_248 ();
 sg13g2_fill_2 FILLER_46_258 ();
 sg13g2_fill_2 FILLER_46_265 ();
 sg13g2_fill_2 FILLER_46_298 ();
 sg13g2_fill_1 FILLER_46_300 ();
 sg13g2_decap_4 FILLER_46_309 ();
 sg13g2_decap_8 FILLER_46_396 ();
 sg13g2_decap_4 FILLER_46_403 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_4 FILLER_47_56 ();
 sg13g2_fill_2 FILLER_47_64 ();
 sg13g2_fill_1 FILLER_47_149 ();
 sg13g2_fill_1 FILLER_47_179 ();
 sg13g2_fill_2 FILLER_47_211 ();
 sg13g2_fill_1 FILLER_47_213 ();
 sg13g2_fill_1 FILLER_47_219 ();
 sg13g2_fill_1 FILLER_47_224 ();
 sg13g2_fill_1 FILLER_47_234 ();
 sg13g2_fill_1 FILLER_47_256 ();
 sg13g2_fill_2 FILLER_47_262 ();
 sg13g2_fill_1 FILLER_47_270 ();
 sg13g2_fill_1 FILLER_47_297 ();
 sg13g2_fill_2 FILLER_47_320 ();
 sg13g2_fill_2 FILLER_47_336 ();
 sg13g2_fill_2 FILLER_47_357 ();
 sg13g2_fill_1 FILLER_47_365 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_fill_2 FILLER_47_406 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_fill_2 FILLER_48_75 ();
 sg13g2_decap_8 FILLER_48_139 ();
 sg13g2_fill_1 FILLER_48_146 ();
 sg13g2_decap_8 FILLER_48_162 ();
 sg13g2_fill_2 FILLER_48_169 ();
 sg13g2_fill_1 FILLER_48_171 ();
 sg13g2_decap_4 FILLER_48_185 ();
 sg13g2_fill_1 FILLER_48_189 ();
 sg13g2_fill_1 FILLER_48_195 ();
 sg13g2_fill_2 FILLER_48_206 ();
 sg13g2_fill_1 FILLER_48_208 ();
 sg13g2_decap_4 FILLER_48_226 ();
 sg13g2_fill_2 FILLER_48_240 ();
 sg13g2_fill_1 FILLER_48_242 ();
 sg13g2_fill_2 FILLER_48_262 ();
 sg13g2_fill_2 FILLER_48_287 ();
 sg13g2_fill_2 FILLER_48_297 ();
 sg13g2_fill_1 FILLER_48_313 ();
 sg13g2_fill_2 FILLER_48_318 ();
 sg13g2_fill_2 FILLER_48_327 ();
 sg13g2_fill_1 FILLER_48_335 ();
 sg13g2_fill_1 FILLER_48_349 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_fill_2 FILLER_48_406 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_4 FILLER_49_49 ();
 sg13g2_fill_2 FILLER_49_53 ();
 sg13g2_fill_1 FILLER_49_103 ();
 sg13g2_fill_1 FILLER_49_114 ();
 sg13g2_decap_8 FILLER_49_144 ();
 sg13g2_decap_8 FILLER_49_151 ();
 sg13g2_decap_8 FILLER_49_158 ();
 sg13g2_decap_4 FILLER_49_165 ();
 sg13g2_fill_2 FILLER_49_179 ();
 sg13g2_fill_2 FILLER_49_200 ();
 sg13g2_fill_1 FILLER_49_202 ();
 sg13g2_fill_2 FILLER_49_209 ();
 sg13g2_fill_2 FILLER_49_219 ();
 sg13g2_fill_1 FILLER_49_221 ();
 sg13g2_fill_2 FILLER_49_227 ();
 sg13g2_fill_1 FILLER_49_229 ();
 sg13g2_decap_8 FILLER_49_235 ();
 sg13g2_fill_2 FILLER_49_242 ();
 sg13g2_fill_1 FILLER_49_244 ();
 sg13g2_decap_8 FILLER_49_250 ();
 sg13g2_fill_1 FILLER_49_257 ();
 sg13g2_fill_1 FILLER_49_267 ();
 sg13g2_decap_4 FILLER_49_273 ();
 sg13g2_fill_1 FILLER_49_277 ();
 sg13g2_fill_2 FILLER_49_291 ();
 sg13g2_fill_1 FILLER_49_302 ();
 sg13g2_decap_8 FILLER_49_398 ();
 sg13g2_decap_4 FILLER_49_405 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_4 FILLER_50_56 ();
 sg13g2_fill_2 FILLER_50_60 ();
 sg13g2_fill_1 FILLER_50_83 ();
 sg13g2_fill_2 FILLER_50_110 ();
 sg13g2_fill_1 FILLER_50_128 ();
 sg13g2_decap_4 FILLER_50_151 ();
 sg13g2_fill_1 FILLER_50_155 ();
 sg13g2_fill_1 FILLER_50_197 ();
 sg13g2_fill_2 FILLER_50_208 ();
 sg13g2_fill_2 FILLER_50_220 ();
 sg13g2_fill_1 FILLER_50_222 ();
 sg13g2_fill_2 FILLER_50_245 ();
 sg13g2_decap_8 FILLER_50_260 ();
 sg13g2_fill_1 FILLER_50_272 ();
 sg13g2_fill_1 FILLER_50_276 ();
 sg13g2_fill_1 FILLER_50_307 ();
 sg13g2_fill_2 FILLER_50_322 ();
 sg13g2_fill_2 FILLER_50_330 ();
 sg13g2_fill_2 FILLER_50_377 ();
 sg13g2_decap_8 FILLER_50_397 ();
 sg13g2_decap_4 FILLER_50_404 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_4 FILLER_51_42 ();
 sg13g2_fill_2 FILLER_51_46 ();
 sg13g2_fill_2 FILLER_51_99 ();
 sg13g2_fill_1 FILLER_51_101 ();
 sg13g2_fill_1 FILLER_51_123 ();
 sg13g2_fill_1 FILLER_51_150 ();
 sg13g2_decap_8 FILLER_51_171 ();
 sg13g2_decap_4 FILLER_51_178 ();
 sg13g2_fill_2 FILLER_51_224 ();
 sg13g2_fill_2 FILLER_51_236 ();
 sg13g2_fill_1 FILLER_51_251 ();
 sg13g2_fill_1 FILLER_51_286 ();
 sg13g2_fill_2 FILLER_51_333 ();
 sg13g2_fill_1 FILLER_51_367 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_fill_2 FILLER_52_42 ();
 sg13g2_fill_1 FILLER_52_77 ();
 sg13g2_fill_2 FILLER_52_87 ();
 sg13g2_fill_1 FILLER_52_181 ();
 sg13g2_fill_2 FILLER_52_257 ();
 sg13g2_fill_1 FILLER_52_259 ();
 sg13g2_fill_1 FILLER_52_293 ();
 sg13g2_fill_1 FILLER_52_358 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_4 FILLER_53_35 ();
 sg13g2_fill_2 FILLER_53_73 ();
 sg13g2_fill_1 FILLER_53_75 ();
 sg13g2_fill_2 FILLER_53_113 ();
 sg13g2_decap_8 FILLER_53_151 ();
 sg13g2_fill_2 FILLER_53_158 ();
 sg13g2_fill_1 FILLER_53_160 ();
 sg13g2_decap_8 FILLER_53_186 ();
 sg13g2_fill_1 FILLER_53_216 ();
 sg13g2_fill_2 FILLER_53_225 ();
 sg13g2_fill_2 FILLER_53_236 ();
 sg13g2_fill_2 FILLER_53_297 ();
 sg13g2_fill_1 FILLER_53_366 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_fill_1 FILLER_54_35 ();
 sg13g2_fill_2 FILLER_54_71 ();
 sg13g2_fill_1 FILLER_54_79 ();
 sg13g2_fill_1 FILLER_54_94 ();
 sg13g2_fill_1 FILLER_54_110 ();
 sg13g2_fill_2 FILLER_54_144 ();
 sg13g2_fill_1 FILLER_54_146 ();
 sg13g2_fill_2 FILLER_54_198 ();
 sg13g2_decap_4 FILLER_54_217 ();
 sg13g2_fill_2 FILLER_54_221 ();
 sg13g2_decap_4 FILLER_54_235 ();
 sg13g2_fill_1 FILLER_54_250 ();
 sg13g2_decap_8 FILLER_54_256 ();
 sg13g2_fill_1 FILLER_54_263 ();
 sg13g2_decap_8 FILLER_54_269 ();
 sg13g2_decap_4 FILLER_54_284 ();
 sg13g2_decap_4 FILLER_54_292 ();
 sg13g2_fill_1 FILLER_54_308 ();
 sg13g2_fill_2 FILLER_54_350 ();
 sg13g2_fill_2 FILLER_54_384 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_4 FILLER_55_35 ();
 sg13g2_fill_2 FILLER_55_39 ();
 sg13g2_fill_1 FILLER_55_140 ();
 sg13g2_fill_1 FILLER_55_154 ();
 sg13g2_decap_4 FILLER_55_160 ();
 sg13g2_fill_1 FILLER_55_164 ();
 sg13g2_decap_4 FILLER_55_169 ();
 sg13g2_fill_1 FILLER_55_173 ();
 sg13g2_decap_8 FILLER_55_178 ();
 sg13g2_fill_2 FILLER_55_185 ();
 sg13g2_fill_1 FILLER_55_187 ();
 sg13g2_decap_4 FILLER_55_201 ();
 sg13g2_fill_2 FILLER_55_224 ();
 sg13g2_decap_4 FILLER_55_265 ();
 sg13g2_fill_1 FILLER_55_329 ();
 sg13g2_decap_8 FILLER_55_401 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_4 FILLER_56_35 ();
 sg13g2_fill_1 FILLER_56_39 ();
 sg13g2_decap_4 FILLER_56_157 ();
 sg13g2_decap_8 FILLER_56_177 ();
 sg13g2_decap_4 FILLER_56_184 ();
 sg13g2_fill_1 FILLER_56_188 ();
 sg13g2_decap_8 FILLER_56_199 ();
 sg13g2_decap_8 FILLER_56_206 ();
 sg13g2_decap_4 FILLER_56_213 ();
 sg13g2_fill_2 FILLER_56_221 ();
 sg13g2_fill_2 FILLER_56_243 ();
 sg13g2_fill_1 FILLER_56_245 ();
 sg13g2_decap_8 FILLER_56_256 ();
 sg13g2_fill_1 FILLER_56_367 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_4 FILLER_57_42 ();
 sg13g2_fill_1 FILLER_57_46 ();
 sg13g2_decap_8 FILLER_57_167 ();
 sg13g2_fill_2 FILLER_57_205 ();
 sg13g2_fill_1 FILLER_57_221 ();
 sg13g2_fill_1 FILLER_57_242 ();
 sg13g2_decap_8 FILLER_57_276 ();
 sg13g2_decap_4 FILLER_57_283 ();
 sg13g2_decap_4 FILLER_57_291 ();
 sg13g2_fill_2 FILLER_57_295 ();
 sg13g2_fill_2 FILLER_57_323 ();
 sg13g2_fill_1 FILLER_57_385 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_4 FILLER_58_42 ();
 sg13g2_decap_4 FILLER_58_83 ();
 sg13g2_fill_2 FILLER_58_87 ();
 sg13g2_fill_2 FILLER_58_101 ();
 sg13g2_fill_1 FILLER_58_112 ();
 sg13g2_fill_1 FILLER_58_125 ();
 sg13g2_fill_1 FILLER_58_153 ();
 sg13g2_fill_1 FILLER_58_180 ();
 sg13g2_fill_2 FILLER_58_195 ();
 sg13g2_fill_1 FILLER_58_197 ();
 sg13g2_fill_2 FILLER_58_208 ();
 sg13g2_fill_2 FILLER_58_214 ();
 sg13g2_fill_2 FILLER_58_272 ();
 sg13g2_fill_1 FILLER_58_274 ();
 sg13g2_decap_8 FILLER_58_279 ();
 sg13g2_fill_2 FILLER_58_286 ();
 sg13g2_decap_4 FILLER_58_292 ();
 sg13g2_fill_1 FILLER_58_296 ();
 sg13g2_fill_1 FILLER_58_332 ();
 sg13g2_decap_4 FILLER_58_403 ();
 sg13g2_fill_2 FILLER_58_407 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_fill_2 FILLER_59_62 ();
 sg13g2_fill_1 FILLER_59_64 ();
 sg13g2_decap_4 FILLER_59_81 ();
 sg13g2_fill_1 FILLER_59_85 ();
 sg13g2_decap_4 FILLER_59_91 ();
 sg13g2_fill_1 FILLER_59_95 ();
 sg13g2_decap_8 FILLER_59_104 ();
 sg13g2_fill_2 FILLER_59_111 ();
 sg13g2_fill_1 FILLER_59_113 ();
 sg13g2_fill_1 FILLER_59_122 ();
 sg13g2_fill_1 FILLER_59_195 ();
 sg13g2_decap_4 FILLER_59_206 ();
 sg13g2_decap_8 FILLER_59_224 ();
 sg13g2_decap_4 FILLER_59_231 ();
 sg13g2_fill_1 FILLER_59_271 ();
 sg13g2_fill_1 FILLER_59_349 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_fill_1 FILLER_60_47 ();
 sg13g2_fill_2 FILLER_60_71 ();
 sg13g2_fill_1 FILLER_60_73 ();
 sg13g2_fill_1 FILLER_60_152 ();
 sg13g2_decap_4 FILLER_60_206 ();
 sg13g2_decap_8 FILLER_60_216 ();
 sg13g2_fill_1 FILLER_60_223 ();
 sg13g2_decap_8 FILLER_60_234 ();
 sg13g2_decap_4 FILLER_60_241 ();
 sg13g2_fill_2 FILLER_60_245 ();
 sg13g2_decap_8 FILLER_60_259 ();
 sg13g2_fill_1 FILLER_60_340 ();
 sg13g2_fill_1 FILLER_60_376 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_4 FILLER_61_21 ();
 sg13g2_fill_1 FILLER_61_59 ();
 sg13g2_fill_2 FILLER_61_92 ();
 sg13g2_fill_2 FILLER_61_143 ();
 sg13g2_fill_1 FILLER_61_145 ();
 sg13g2_fill_1 FILLER_61_172 ();
 sg13g2_decap_8 FILLER_61_177 ();
 sg13g2_decap_4 FILLER_61_184 ();
 sg13g2_fill_2 FILLER_61_188 ();
 sg13g2_fill_1 FILLER_61_218 ();
 sg13g2_decap_8 FILLER_61_242 ();
 sg13g2_decap_4 FILLER_61_249 ();
 sg13g2_fill_1 FILLER_61_261 ();
 sg13g2_fill_1 FILLER_61_267 ();
 sg13g2_fill_1 FILLER_61_273 ();
 sg13g2_fill_1 FILLER_61_282 ();
 sg13g2_fill_1 FILLER_61_289 ();
 sg13g2_fill_2 FILLER_61_316 ();
 sg13g2_fill_1 FILLER_61_333 ();
 sg13g2_fill_2 FILLER_61_406 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_4 FILLER_62_14 ();
 sg13g2_fill_1 FILLER_62_58 ();
 sg13g2_fill_2 FILLER_62_136 ();
 sg13g2_fill_2 FILLER_62_162 ();
 sg13g2_fill_2 FILLER_62_180 ();
 sg13g2_fill_2 FILLER_62_195 ();
 sg13g2_fill_1 FILLER_62_197 ();
 sg13g2_fill_1 FILLER_62_203 ();
 sg13g2_fill_1 FILLER_62_237 ();
 sg13g2_fill_2 FILLER_62_248 ();
 sg13g2_fill_1 FILLER_62_250 ();
 sg13g2_decap_4 FILLER_62_255 ();
 sg13g2_fill_1 FILLER_62_308 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_fill_2 FILLER_63_21 ();
 sg13g2_fill_2 FILLER_63_49 ();
 sg13g2_fill_1 FILLER_63_51 ();
 sg13g2_fill_1 FILLER_63_84 ();
 sg13g2_fill_2 FILLER_63_111 ();
 sg13g2_fill_1 FILLER_63_122 ();
 sg13g2_fill_1 FILLER_63_136 ();
 sg13g2_fill_1 FILLER_63_162 ();
 sg13g2_fill_2 FILLER_63_223 ();
 sg13g2_fill_1 FILLER_63_225 ();
 sg13g2_fill_1 FILLER_63_254 ();
 sg13g2_fill_2 FILLER_63_299 ();
 sg13g2_fill_2 FILLER_63_334 ();
 sg13g2_fill_2 FILLER_63_356 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_fill_2 FILLER_64_14 ();
 sg13g2_fill_2 FILLER_64_69 ();
 sg13g2_fill_1 FILLER_64_84 ();
 sg13g2_fill_1 FILLER_64_124 ();
 sg13g2_fill_1 FILLER_64_146 ();
 sg13g2_fill_1 FILLER_64_223 ();
 sg13g2_fill_1 FILLER_64_261 ();
 sg13g2_fill_1 FILLER_64_275 ();
 sg13g2_fill_2 FILLER_64_291 ();
 sg13g2_fill_2 FILLER_64_339 ();
 sg13g2_fill_2 FILLER_64_355 ();
 sg13g2_fill_2 FILLER_64_406 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_4 FILLER_65_21 ();
 sg13g2_fill_2 FILLER_65_25 ();
 sg13g2_fill_1 FILLER_65_58 ();
 sg13g2_fill_1 FILLER_65_71 ();
 sg13g2_fill_1 FILLER_65_77 ();
 sg13g2_fill_2 FILLER_65_103 ();
 sg13g2_fill_2 FILLER_65_122 ();
 sg13g2_fill_2 FILLER_65_150 ();
 sg13g2_decap_8 FILLER_65_175 ();
 sg13g2_decap_8 FILLER_65_182 ();
 sg13g2_decap_4 FILLER_65_189 ();
 sg13g2_fill_1 FILLER_65_193 ();
 sg13g2_fill_2 FILLER_65_203 ();
 sg13g2_decap_4 FILLER_65_210 ();
 sg13g2_fill_1 FILLER_65_214 ();
 sg13g2_fill_1 FILLER_65_225 ();
 sg13g2_decap_4 FILLER_65_230 ();
 sg13g2_fill_1 FILLER_65_234 ();
 sg13g2_fill_2 FILLER_65_258 ();
 sg13g2_fill_2 FILLER_65_265 ();
 sg13g2_fill_1 FILLER_65_293 ();
 sg13g2_fill_2 FILLER_65_325 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_fill_1 FILLER_66_28 ();
 sg13g2_fill_2 FILLER_66_46 ();
 sg13g2_fill_1 FILLER_66_48 ();
 sg13g2_fill_1 FILLER_66_57 ();
 sg13g2_fill_2 FILLER_66_162 ();
 sg13g2_fill_1 FILLER_66_164 ();
 sg13g2_decap_4 FILLER_66_211 ();
 sg13g2_fill_2 FILLER_66_215 ();
 sg13g2_fill_1 FILLER_66_231 ();
 sg13g2_decap_4 FILLER_66_250 ();
 sg13g2_fill_1 FILLER_66_254 ();
 sg13g2_fill_2 FILLER_66_269 ();
 sg13g2_fill_1 FILLER_66_271 ();
 sg13g2_fill_2 FILLER_66_319 ();
 sg13g2_decap_8 FILLER_66_399 ();
 sg13g2_fill_2 FILLER_66_406 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_4 FILLER_67_14 ();
 sg13g2_fill_1 FILLER_67_18 ();
 sg13g2_fill_2 FILLER_67_54 ();
 sg13g2_fill_1 FILLER_67_56 ();
 sg13g2_fill_2 FILLER_67_65 ();
 sg13g2_fill_1 FILLER_67_67 ();
 sg13g2_fill_2 FILLER_67_75 ();
 sg13g2_fill_2 FILLER_67_144 ();
 sg13g2_decap_4 FILLER_67_202 ();
 sg13g2_fill_2 FILLER_67_223 ();
 sg13g2_fill_1 FILLER_67_225 ();
 sg13g2_fill_2 FILLER_67_236 ();
 sg13g2_fill_1 FILLER_67_238 ();
 sg13g2_fill_2 FILLER_67_248 ();
 sg13g2_fill_1 FILLER_67_255 ();
 sg13g2_decap_4 FILLER_67_261 ();
 sg13g2_decap_4 FILLER_67_273 ();
 sg13g2_fill_1 FILLER_67_284 ();
 sg13g2_fill_2 FILLER_67_302 ();
 sg13g2_fill_2 FILLER_67_379 ();
 sg13g2_decap_8 FILLER_67_394 ();
 sg13g2_decap_8 FILLER_67_401 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_4 FILLER_68_21 ();
 sg13g2_fill_1 FILLER_68_54 ();
 sg13g2_fill_2 FILLER_68_131 ();
 sg13g2_fill_1 FILLER_68_133 ();
 sg13g2_decap_4 FILLER_68_195 ();
 sg13g2_fill_1 FILLER_68_215 ();
 sg13g2_fill_1 FILLER_68_304 ();
 sg13g2_fill_1 FILLER_68_324 ();
 sg13g2_fill_1 FILLER_68_365 ();
 sg13g2_decap_8 FILLER_68_398 ();
 sg13g2_decap_4 FILLER_68_405 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_fill_2 FILLER_69_35 ();
 sg13g2_fill_1 FILLER_69_54 ();
 sg13g2_fill_1 FILLER_69_61 ();
 sg13g2_fill_1 FILLER_69_96 ();
 sg13g2_fill_2 FILLER_69_114 ();
 sg13g2_fill_1 FILLER_69_121 ();
 sg13g2_fill_2 FILLER_69_129 ();
 sg13g2_fill_1 FILLER_69_141 ();
 sg13g2_decap_4 FILLER_69_161 ();
 sg13g2_decap_8 FILLER_69_169 ();
 sg13g2_decap_4 FILLER_69_176 ();
 sg13g2_fill_1 FILLER_69_180 ();
 sg13g2_fill_2 FILLER_69_185 ();
 sg13g2_fill_1 FILLER_69_196 ();
 sg13g2_decap_8 FILLER_69_200 ();
 sg13g2_fill_2 FILLER_69_207 ();
 sg13g2_decap_8 FILLER_69_236 ();
 sg13g2_fill_2 FILLER_69_243 ();
 sg13g2_fill_1 FILLER_69_245 ();
 sg13g2_fill_2 FILLER_69_252 ();
 sg13g2_decap_8 FILLER_69_261 ();
 sg13g2_decap_8 FILLER_69_268 ();
 sg13g2_fill_1 FILLER_69_275 ();
 sg13g2_fill_1 FILLER_69_286 ();
 sg13g2_fill_2 FILLER_69_330 ();
 sg13g2_decap_8 FILLER_69_395 ();
 sg13g2_decap_8 FILLER_69_402 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_fill_2 FILLER_70_42 ();
 sg13g2_fill_1 FILLER_70_68 ();
 sg13g2_fill_2 FILLER_70_79 ();
 sg13g2_decap_8 FILLER_70_87 ();
 sg13g2_decap_4 FILLER_70_94 ();
 sg13g2_decap_4 FILLER_70_174 ();
 sg13g2_fill_2 FILLER_70_178 ();
 sg13g2_decap_8 FILLER_70_207 ();
 sg13g2_decap_8 FILLER_70_214 ();
 sg13g2_decap_8 FILLER_70_229 ();
 sg13g2_fill_2 FILLER_70_236 ();
 sg13g2_fill_1 FILLER_70_238 ();
 sg13g2_fill_1 FILLER_70_255 ();
 sg13g2_fill_2 FILLER_70_269 ();
 sg13g2_fill_2 FILLER_70_288 ();
 sg13g2_fill_1 FILLER_70_290 ();
 sg13g2_fill_2 FILLER_70_356 ();
 sg13g2_fill_1 FILLER_70_364 ();
 sg13g2_fill_1 FILLER_70_379 ();
 sg13g2_decap_8 FILLER_70_394 ();
 sg13g2_decap_8 FILLER_70_401 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_4 FILLER_71_28 ();
 sg13g2_decap_4 FILLER_71_35 ();
 sg13g2_fill_1 FILLER_71_39 ();
 sg13g2_decap_8 FILLER_71_48 ();
 sg13g2_decap_4 FILLER_71_55 ();
 sg13g2_decap_8 FILLER_71_146 ();
 sg13g2_fill_2 FILLER_71_153 ();
 sg13g2_fill_2 FILLER_71_163 ();
 sg13g2_fill_1 FILLER_71_195 ();
 sg13g2_fill_2 FILLER_71_210 ();
 sg13g2_fill_1 FILLER_71_212 ();
 sg13g2_decap_8 FILLER_71_217 ();
 sg13g2_fill_2 FILLER_71_224 ();
 sg13g2_fill_1 FILLER_71_226 ();
 sg13g2_fill_1 FILLER_71_232 ();
 sg13g2_fill_2 FILLER_71_238 ();
 sg13g2_decap_8 FILLER_71_245 ();
 sg13g2_decap_4 FILLER_71_257 ();
 sg13g2_fill_2 FILLER_71_340 ();
 sg13g2_decap_8 FILLER_71_391 ();
 sg13g2_decap_8 FILLER_71_398 ();
 sg13g2_decap_4 FILLER_71_405 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_4 FILLER_72_21 ();
 sg13g2_fill_2 FILLER_72_117 ();
 sg13g2_fill_2 FILLER_72_146 ();
 sg13g2_fill_2 FILLER_72_155 ();
 sg13g2_fill_2 FILLER_72_183 ();
 sg13g2_fill_2 FILLER_72_194 ();
 sg13g2_fill_1 FILLER_72_196 ();
 sg13g2_fill_1 FILLER_72_209 ();
 sg13g2_fill_1 FILLER_72_216 ();
 sg13g2_decap_8 FILLER_72_231 ();
 sg13g2_decap_8 FILLER_72_238 ();
 sg13g2_fill_2 FILLER_72_299 ();
 sg13g2_fill_1 FILLER_72_301 ();
 sg13g2_fill_2 FILLER_72_311 ();
 sg13g2_fill_1 FILLER_72_313 ();
 sg13g2_decap_8 FILLER_72_402 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_4 FILLER_73_21 ();
 sg13g2_fill_2 FILLER_73_25 ();
 sg13g2_fill_2 FILLER_73_55 ();
 sg13g2_fill_1 FILLER_73_70 ();
 sg13g2_fill_1 FILLER_73_89 ();
 sg13g2_fill_1 FILLER_73_95 ();
 sg13g2_fill_2 FILLER_73_104 ();
 sg13g2_fill_1 FILLER_73_106 ();
 sg13g2_fill_1 FILLER_73_122 ();
 sg13g2_fill_1 FILLER_73_195 ();
 sg13g2_fill_1 FILLER_73_242 ();
 sg13g2_fill_2 FILLER_73_255 ();
 sg13g2_fill_2 FILLER_73_286 ();
 sg13g2_fill_1 FILLER_73_288 ();
 sg13g2_decap_8 FILLER_73_397 ();
 sg13g2_decap_4 FILLER_73_404 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_4 FILLER_74_28 ();
 sg13g2_fill_1 FILLER_74_49 ();
 sg13g2_fill_2 FILLER_74_63 ();
 sg13g2_fill_1 FILLER_74_78 ();
 sg13g2_fill_2 FILLER_74_119 ();
 sg13g2_fill_1 FILLER_74_121 ();
 sg13g2_fill_2 FILLER_74_138 ();
 sg13g2_fill_1 FILLER_74_140 ();
 sg13g2_fill_2 FILLER_74_165 ();
 sg13g2_fill_1 FILLER_74_167 ();
 sg13g2_fill_1 FILLER_74_207 ();
 sg13g2_fill_1 FILLER_74_233 ();
 sg13g2_fill_2 FILLER_74_283 ();
 sg13g2_fill_1 FILLER_74_285 ();
 sg13g2_fill_2 FILLER_74_329 ();
 sg13g2_fill_1 FILLER_74_331 ();
 sg13g2_fill_1 FILLER_74_357 ();
 sg13g2_decap_4 FILLER_74_403 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_fill_2 FILLER_75_28 ();
 sg13g2_decap_4 FILLER_75_56 ();
 sg13g2_fill_1 FILLER_75_69 ();
 sg13g2_fill_1 FILLER_75_84 ();
 sg13g2_fill_1 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_172 ();
 sg13g2_fill_1 FILLER_75_179 ();
 sg13g2_fill_2 FILLER_75_193 ();
 sg13g2_fill_1 FILLER_75_205 ();
 sg13g2_fill_1 FILLER_75_209 ();
 sg13g2_decap_8 FILLER_75_219 ();
 sg13g2_fill_1 FILLER_75_226 ();
 sg13g2_fill_1 FILLER_75_242 ();
 sg13g2_fill_1 FILLER_75_273 ();
 sg13g2_fill_1 FILLER_75_287 ();
 sg13g2_fill_1 FILLER_75_315 ();
 sg13g2_fill_2 FILLER_75_330 ();
 sg13g2_decap_8 FILLER_75_396 ();
 sg13g2_decap_4 FILLER_75_403 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_fill_2 FILLER_76_57 ();
 sg13g2_fill_1 FILLER_76_59 ();
 sg13g2_fill_2 FILLER_76_86 ();
 sg13g2_fill_1 FILLER_76_102 ();
 sg13g2_fill_1 FILLER_76_147 ();
 sg13g2_fill_2 FILLER_76_174 ();
 sg13g2_fill_1 FILLER_76_199 ();
 sg13g2_fill_2 FILLER_76_205 ();
 sg13g2_fill_1 FILLER_76_243 ();
 sg13g2_fill_1 FILLER_76_256 ();
 sg13g2_fill_2 FILLER_76_262 ();
 sg13g2_fill_1 FILLER_76_273 ();
 sg13g2_fill_1 FILLER_76_326 ();
 sg13g2_fill_2 FILLER_76_336 ();
 sg13g2_fill_2 FILLER_76_352 ();
 sg13g2_decap_8 FILLER_76_401 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_fill_1 FILLER_77_21 ();
 sg13g2_fill_1 FILLER_77_46 ();
 sg13g2_fill_2 FILLER_77_113 ();
 sg13g2_fill_2 FILLER_77_158 ();
 sg13g2_decap_4 FILLER_77_244 ();
 sg13g2_fill_2 FILLER_77_271 ();
 sg13g2_decap_8 FILLER_77_391 ();
 sg13g2_decap_8 FILLER_77_398 ();
 sg13g2_decap_4 FILLER_77_405 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_fill_2 FILLER_78_28 ();
 sg13g2_fill_1 FILLER_78_60 ();
 sg13g2_fill_1 FILLER_78_79 ();
 sg13g2_fill_2 FILLER_78_89 ();
 sg13g2_fill_1 FILLER_78_91 ();
 sg13g2_fill_1 FILLER_78_174 ();
 sg13g2_fill_1 FILLER_78_179 ();
 sg13g2_fill_2 FILLER_78_203 ();
 sg13g2_decap_4 FILLER_78_236 ();
 sg13g2_fill_2 FILLER_78_240 ();
 sg13g2_fill_1 FILLER_78_268 ();
 sg13g2_fill_1 FILLER_78_309 ();
 sg13g2_decap_8 FILLER_78_384 ();
 sg13g2_decap_8 FILLER_78_391 ();
 sg13g2_decap_8 FILLER_78_398 ();
 sg13g2_decap_4 FILLER_78_405 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_fill_1 FILLER_79_28 ();
 sg13g2_fill_2 FILLER_79_85 ();
 sg13g2_fill_2 FILLER_79_143 ();
 sg13g2_fill_1 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_218 ();
 sg13g2_decap_8 FILLER_79_229 ();
 sg13g2_decap_4 FILLER_79_236 ();
 sg13g2_fill_2 FILLER_79_240 ();
 sg13g2_decap_8 FILLER_79_273 ();
 sg13g2_fill_2 FILLER_79_284 ();
 sg13g2_fill_2 FILLER_79_329 ();
 sg13g2_fill_2 FILLER_79_345 ();
 sg13g2_decap_8 FILLER_79_377 ();
 sg13g2_decap_8 FILLER_79_384 ();
 sg13g2_decap_8 FILLER_79_391 ();
 sg13g2_decap_8 FILLER_79_398 ();
 sg13g2_decap_4 FILLER_79_405 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_4 FILLER_80_21 ();
 sg13g2_fill_2 FILLER_80_66 ();
 sg13g2_fill_1 FILLER_80_68 ();
 sg13g2_fill_2 FILLER_80_74 ();
 sg13g2_fill_1 FILLER_80_76 ();
 sg13g2_fill_1 FILLER_80_101 ();
 sg13g2_fill_1 FILLER_80_115 ();
 sg13g2_fill_2 FILLER_80_142 ();
 sg13g2_fill_2 FILLER_80_157 ();
 sg13g2_fill_1 FILLER_80_159 ();
 sg13g2_decap_4 FILLER_80_180 ();
 sg13g2_fill_2 FILLER_80_188 ();
 sg13g2_fill_2 FILLER_80_198 ();
 sg13g2_decap_4 FILLER_80_204 ();
 sg13g2_decap_4 FILLER_80_220 ();
 sg13g2_decap_4 FILLER_80_228 ();
 sg13g2_decap_8 FILLER_80_236 ();
 sg13g2_decap_8 FILLER_80_243 ();
 sg13g2_fill_2 FILLER_80_250 ();
 sg13g2_fill_1 FILLER_80_252 ();
 sg13g2_fill_2 FILLER_80_266 ();
 sg13g2_decap_8 FILLER_80_277 ();
 sg13g2_decap_8 FILLER_80_284 ();
 sg13g2_fill_1 FILLER_80_318 ();
 sg13g2_fill_2 FILLER_80_328 ();
 sg13g2_fill_2 FILLER_80_335 ();
 sg13g2_fill_1 FILLER_80_346 ();
 sg13g2_decap_8 FILLER_80_374 ();
 sg13g2_decap_8 FILLER_80_381 ();
 sg13g2_decap_8 FILLER_80_388 ();
 sg13g2_decap_8 FILLER_80_395 ();
 sg13g2_decap_8 FILLER_80_402 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
 assign uo_out[1] = net18;
 assign uo_out[2] = net19;
 assign uo_out[3] = net20;
 assign uo_out[4] = net21;
 assign uo_out[5] = net22;
 assign uo_out[6] = net23;
 assign uo_out[7] = net24;
endmodule

module tt_um_rejunity_e2m0_x_i8_matmul (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire clknet_leaf_0_clk;
 wire net32;
 wire \systolic_array.arg_left_div2_next[0] ;
 wire \systolic_array.arg_left_div2_next[1] ;
 wire \systolic_array.arg_left_div2_next[3] ;
 wire \systolic_array.arg_left_div2_next[4] ;
 wire \systolic_array.arg_left_mul2_next[0] ;
 wire \systolic_array.arg_left_mul2_next[1] ;
 wire \systolic_array.arg_left_mul2_next[2] ;
 wire \systolic_array.arg_left_mul2_next[3] ;
 wire \systolic_array.arg_left_mul2_next[4] ;
 wire \systolic_array.arg_left_mul2_next[5] ;
 wire \systolic_array.arg_left_sign_next[0] ;
 wire \systolic_array.arg_left_sign_next[1] ;
 wire \systolic_array.arg_left_sign_next[2] ;
 wire \systolic_array.arg_left_sign_next[3] ;
 wire \systolic_array.arg_left_sign_next[4] ;
 wire \systolic_array.arg_left_sign_next[5] ;
 wire \systolic_array.arg_left_zero_next[0] ;
 wire \systolic_array.arg_left_zero_next[1] ;
 wire \systolic_array.arg_left_zero_next[2] ;
 wire \systolic_array.arg_left_zero_next[3] ;
 wire \systolic_array.arg_left_zero_next[4] ;
 wire \systolic_array.arg_left_zero_next[5] ;
 wire \systolic_array.arg_top_curr[0] ;
 wire \systolic_array.arg_top_curr[10] ;
 wire \systolic_array.arg_top_curr[11] ;
 wire \systolic_array.arg_top_curr[12] ;
 wire \systolic_array.arg_top_curr[13] ;
 wire \systolic_array.arg_top_curr[14] ;
 wire \systolic_array.arg_top_curr[15] ;
 wire \systolic_array.arg_top_curr[1] ;
 wire \systolic_array.arg_top_curr[2] ;
 wire \systolic_array.arg_top_curr[3] ;
 wire \systolic_array.arg_top_curr[4] ;
 wire \systolic_array.arg_top_curr[5] ;
 wire \systolic_array.arg_top_curr[6] ;
 wire \systolic_array.arg_top_curr[7] ;
 wire \systolic_array.arg_top_curr[8] ;
 wire \systolic_array.arg_top_curr[9] ;
 wire \systolic_array.arg_top_next[0] ;
 wire \systolic_array.arg_top_next[10] ;
 wire \systolic_array.arg_top_next[11] ;
 wire \systolic_array.arg_top_next[12] ;
 wire \systolic_array.arg_top_next[13] ;
 wire \systolic_array.arg_top_next[14] ;
 wire \systolic_array.arg_top_next[15] ;
 wire \systolic_array.arg_top_next[1] ;
 wire \systolic_array.arg_top_next[2] ;
 wire \systolic_array.arg_top_next[3] ;
 wire \systolic_array.arg_top_next[4] ;
 wire \systolic_array.arg_top_next[5] ;
 wire \systolic_array.arg_top_next[6] ;
 wire \systolic_array.arg_top_next[7] ;
 wire \systolic_array.arg_top_next[8] ;
 wire \systolic_array.arg_top_next[9] ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[0].A ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[10].A ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[11].A ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[12].A ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[13].A ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[14].A ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[15].A ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[16].A ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[1].A ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[2].A ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[3].A ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[4].A ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[5].A ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[6].A ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[7].A ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[8].A ;
 wire \systolic_array.genblk1[0].accumulators_dlygate[9].A ;
 wire \systolic_array.genblk1[0].out_queue_dlygate[10].A ;
 wire \systolic_array.genblk1[0].out_queue_dlygate[11].A ;
 wire \systolic_array.genblk1[0].out_queue_dlygate[12].A ;
 wire \systolic_array.genblk1[0].out_queue_dlygate[13].A ;
 wire \systolic_array.genblk1[0].out_queue_dlygate[14].A ;
 wire \systolic_array.genblk1[0].out_queue_dlygate[15].A ;
 wire \systolic_array.genblk1[0].out_queue_dlygate[16].A ;
 wire \systolic_array.genblk1[0].out_queue_dlygate[9].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[0].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[10].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[11].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[12].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[13].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[14].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[15].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[16].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[1].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[2].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[3].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[4].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[5].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[6].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[7].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[8].A ;
 wire \systolic_array.genblk1[10].accumulators_dlygate[9].A ;
 wire \systolic_array.genblk1[10].out_queue_dlygate[10].A ;
 wire \systolic_array.genblk1[10].out_queue_dlygate[11].A ;
 wire \systolic_array.genblk1[10].out_queue_dlygate[12].A ;
 wire \systolic_array.genblk1[10].out_queue_dlygate[13].A ;
 wire \systolic_array.genblk1[10].out_queue_dlygate[14].A ;
 wire \systolic_array.genblk1[10].out_queue_dlygate[15].A ;
 wire \systolic_array.genblk1[10].out_queue_dlygate[16].A ;
 wire \systolic_array.genblk1[10].out_queue_dlygate[9].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[0].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[10].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[11].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[12].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[13].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[14].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[15].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[16].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[1].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[2].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[3].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[4].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[5].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[6].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[7].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[8].A ;
 wire \systolic_array.genblk1[11].accumulators_dlygate[9].A ;
 wire \systolic_array.genblk1[11].out_queue_dlygate[10].A ;
 wire \systolic_array.genblk1[11].out_queue_dlygate[11].A ;
 wire \systolic_array.genblk1[11].out_queue_dlygate[12].A ;
 wire \systolic_array.genblk1[11].out_queue_dlygate[13].A ;
 wire \systolic_array.genblk1[11].out_queue_dlygate[14].A ;
 wire \systolic_array.genblk1[11].out_queue_dlygate[15].A ;
 wire \systolic_array.genblk1[11].out_queue_dlygate[16].A ;
 wire \systolic_array.genblk1[11].out_queue_dlygate[9].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[0].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[10].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[11].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[12].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[13].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[14].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[15].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[16].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[1].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[2].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[3].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[4].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[5].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[6].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[7].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[8].A ;
 wire \systolic_array.genblk1[1].accumulators_dlygate[9].A ;
 wire \systolic_array.genblk1[1].out_queue_dlygate[10].A ;
 wire \systolic_array.genblk1[1].out_queue_dlygate[11].A ;
 wire \systolic_array.genblk1[1].out_queue_dlygate[12].A ;
 wire \systolic_array.genblk1[1].out_queue_dlygate[13].A ;
 wire \systolic_array.genblk1[1].out_queue_dlygate[14].A ;
 wire \systolic_array.genblk1[1].out_queue_dlygate[15].A ;
 wire \systolic_array.genblk1[1].out_queue_dlygate[16].A ;
 wire \systolic_array.genblk1[1].out_queue_dlygate[9].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[0].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[10].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[11].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[12].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[13].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[14].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[15].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[16].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[1].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[2].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[3].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[4].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[5].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[6].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[7].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[8].A ;
 wire \systolic_array.genblk1[2].accumulators_dlygate[9].A ;
 wire \systolic_array.genblk1[2].out_queue_dlygate[10].A ;
 wire \systolic_array.genblk1[2].out_queue_dlygate[11].A ;
 wire \systolic_array.genblk1[2].out_queue_dlygate[12].A ;
 wire \systolic_array.genblk1[2].out_queue_dlygate[13].A ;
 wire \systolic_array.genblk1[2].out_queue_dlygate[14].A ;
 wire \systolic_array.genblk1[2].out_queue_dlygate[15].A ;
 wire \systolic_array.genblk1[2].out_queue_dlygate[16].A ;
 wire \systolic_array.genblk1[2].out_queue_dlygate[9].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[0].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[10].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[11].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[12].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[13].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[14].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[15].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[16].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[1].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[2].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[3].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[4].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[5].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[6].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[7].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[8].A ;
 wire \systolic_array.genblk1[3].accumulators_dlygate[9].A ;
 wire \systolic_array.genblk1[3].out_queue_dlygate[10].A ;
 wire \systolic_array.genblk1[3].out_queue_dlygate[11].A ;
 wire \systolic_array.genblk1[3].out_queue_dlygate[12].A ;
 wire \systolic_array.genblk1[3].out_queue_dlygate[13].A ;
 wire \systolic_array.genblk1[3].out_queue_dlygate[14].A ;
 wire \systolic_array.genblk1[3].out_queue_dlygate[15].A ;
 wire \systolic_array.genblk1[3].out_queue_dlygate[16].A ;
 wire \systolic_array.genblk1[3].out_queue_dlygate[9].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[0].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[10].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[11].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[12].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[13].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[14].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[15].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[16].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[1].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[2].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[3].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[4].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[5].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[6].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[7].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[8].A ;
 wire \systolic_array.genblk1[4].accumulators_dlygate[9].A ;
 wire \systolic_array.genblk1[4].out_queue_dlygate[10].A ;
 wire \systolic_array.genblk1[4].out_queue_dlygate[11].A ;
 wire \systolic_array.genblk1[4].out_queue_dlygate[12].A ;
 wire \systolic_array.genblk1[4].out_queue_dlygate[13].A ;
 wire \systolic_array.genblk1[4].out_queue_dlygate[14].A ;
 wire \systolic_array.genblk1[4].out_queue_dlygate[15].A ;
 wire \systolic_array.genblk1[4].out_queue_dlygate[16].A ;
 wire \systolic_array.genblk1[4].out_queue_dlygate[9].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[0].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[10].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[11].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[12].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[13].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[14].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[15].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[16].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[1].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[2].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[3].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[4].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[5].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[6].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[7].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[8].A ;
 wire \systolic_array.genblk1[5].accumulators_dlygate[9].A ;
 wire \systolic_array.genblk1[5].out_queue_dlygate[10].A ;
 wire \systolic_array.genblk1[5].out_queue_dlygate[11].A ;
 wire \systolic_array.genblk1[5].out_queue_dlygate[12].A ;
 wire \systolic_array.genblk1[5].out_queue_dlygate[13].A ;
 wire \systolic_array.genblk1[5].out_queue_dlygate[14].A ;
 wire \systolic_array.genblk1[5].out_queue_dlygate[15].A ;
 wire \systolic_array.genblk1[5].out_queue_dlygate[16].A ;
 wire \systolic_array.genblk1[5].out_queue_dlygate[9].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[0].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[10].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[11].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[12].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[13].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[14].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[15].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[16].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[1].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[2].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[3].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[4].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[5].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[6].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[7].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[8].A ;
 wire \systolic_array.genblk1[6].accumulators_dlygate[9].A ;
 wire \systolic_array.genblk1[6].out_queue_dlygate[10].A ;
 wire \systolic_array.genblk1[6].out_queue_dlygate[11].A ;
 wire \systolic_array.genblk1[6].out_queue_dlygate[12].A ;
 wire \systolic_array.genblk1[6].out_queue_dlygate[13].A ;
 wire \systolic_array.genblk1[6].out_queue_dlygate[14].A ;
 wire \systolic_array.genblk1[6].out_queue_dlygate[15].A ;
 wire \systolic_array.genblk1[6].out_queue_dlygate[16].A ;
 wire \systolic_array.genblk1[6].out_queue_dlygate[9].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[0].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[10].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[11].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[12].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[13].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[14].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[15].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[16].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[1].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[2].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[3].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[4].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[5].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[6].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[7].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[8].A ;
 wire \systolic_array.genblk1[7].accumulators_dlygate[9].A ;
 wire \systolic_array.genblk1[7].out_queue_dlygate[10].A ;
 wire \systolic_array.genblk1[7].out_queue_dlygate[11].A ;
 wire \systolic_array.genblk1[7].out_queue_dlygate[12].A ;
 wire \systolic_array.genblk1[7].out_queue_dlygate[13].A ;
 wire \systolic_array.genblk1[7].out_queue_dlygate[14].A ;
 wire \systolic_array.genblk1[7].out_queue_dlygate[15].A ;
 wire \systolic_array.genblk1[7].out_queue_dlygate[16].A ;
 wire \systolic_array.genblk1[7].out_queue_dlygate[9].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[0].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[10].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[11].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[12].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[13].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[14].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[15].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[16].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[1].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[2].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[3].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[4].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[5].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[6].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[7].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[8].A ;
 wire \systolic_array.genblk1[8].accumulators_dlygate[9].A ;
 wire \systolic_array.genblk1[8].out_queue_dlygate[10].A ;
 wire \systolic_array.genblk1[8].out_queue_dlygate[11].A ;
 wire \systolic_array.genblk1[8].out_queue_dlygate[12].A ;
 wire \systolic_array.genblk1[8].out_queue_dlygate[13].A ;
 wire \systolic_array.genblk1[8].out_queue_dlygate[14].A ;
 wire \systolic_array.genblk1[8].out_queue_dlygate[15].A ;
 wire \systolic_array.genblk1[8].out_queue_dlygate[16].A ;
 wire \systolic_array.genblk1[8].out_queue_dlygate[9].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[0].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[10].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[11].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[12].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[13].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[14].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[15].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[16].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[1].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[2].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[3].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[4].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[5].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[6].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[7].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[8].A ;
 wire \systolic_array.genblk1[9].accumulators_dlygate[9].A ;
 wire \systolic_array.genblk1[9].out_queue_dlygate[10].A ;
 wire \systolic_array.genblk1[9].out_queue_dlygate[11].A ;
 wire \systolic_array.genblk1[9].out_queue_dlygate[12].A ;
 wire \systolic_array.genblk1[9].out_queue_dlygate[13].A ;
 wire \systolic_array.genblk1[9].out_queue_dlygate[14].A ;
 wire \systolic_array.genblk1[9].out_queue_dlygate[15].A ;
 wire \systolic_array.genblk1[9].out_queue_dlygate[16].A ;
 wire \systolic_array.genblk1[9].out_queue_dlygate[9].A ;
 wire \systolic_array.genblk2[0].mac[0].div2 ;
 wire \systolic_array.genblk2[0].mac[0].mul2 ;
 wire \systolic_array.genblk2[0].mac[0].sign ;
 wire \systolic_array.genblk2[0].mac[0].zero ;
 wire \systolic_array.genblk2[0].mac[1].div2 ;
 wire \systolic_array.genblk2[0].mac[1].mul2 ;
 wire \systolic_array.genblk2[0].mac[1].sign ;
 wire \systolic_array.genblk2[0].mac[1].zero ;
 wire \systolic_array.genblk2[0].mac[2].mul2 ;
 wire \systolic_array.genblk2[0].mac[2].sign ;
 wire \systolic_array.genblk2[0].mac[2].zero ;
 wire \systolic_array.genblk2[0].mac[3].div2 ;
 wire \systolic_array.genblk2[0].mac[3].mul2 ;
 wire \systolic_array.genblk2[0].mac[3].sign ;
 wire \systolic_array.genblk2[0].mac[3].zero ;
 wire \systolic_array.genblk2[0].mac[4].div2 ;
 wire \systolic_array.genblk2[0].mac[4].mul2 ;
 wire \systolic_array.genblk2[0].mac[4].sign ;
 wire \systolic_array.genblk2[0].mac[4].zero ;
 wire \systolic_array.genblk2[0].mac[5].mul2 ;
 wire \systolic_array.genblk2[0].mac[5].sign ;
 wire \systolic_array.genblk2[0].mac[5].zero ;
 wire \systolic_array.slice_counter ;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;

 sg13g2_inv_2 _2395_ (.Y(_1460_),
    .A(net719));
 sg13g2_inv_1 _2396_ (.Y(_1461_),
    .A(net697));
 sg13g2_inv_1 _2397_ (.Y(_1462_),
    .A(net701));
 sg13g2_inv_4 _2398_ (.A(net5),
    .Y(_1463_));
 sg13g2_inv_1 _2399_ (.Y(_1464_),
    .A(net698));
 sg13g2_inv_4 _2400_ (.A(net678),
    .Y(_1465_));
 sg13g2_inv_2 _2401_ (.Y(_1466_),
    .A(\systolic_array.arg_top_curr[6] ));
 sg13g2_inv_4 _2402_ (.A(_0115_),
    .Y(_1467_));
 sg13g2_inv_2 _2403_ (.Y(_1468_),
    .A(net680));
 sg13g2_inv_2 _2404_ (.Y(_1469_),
    .A(\systolic_array.arg_top_curr[4] ));
 sg13g2_inv_1 _2405_ (.Y(_1470_),
    .A(\systolic_array.arg_top_curr[0] ));
 sg13g2_inv_2 _2406_ (.Y(_1471_),
    .A(\systolic_array.genblk2[0].mac[0].sign ));
 sg13g2_inv_1 _2407_ (.Y(_1472_),
    .A(net836));
 sg13g2_inv_1 _2408_ (.Y(_1473_),
    .A(\systolic_array.genblk1[0].accumulators_dlygate[7].A ));
 sg13g2_inv_1 _2409_ (.Y(_1474_),
    .A(\systolic_array.genblk1[0].accumulators_dlygate[5].A ));
 sg13g2_inv_1 _2410_ (.Y(_1475_),
    .A(net902));
 sg13g2_inv_1 _2411_ (.Y(_1476_),
    .A(net879));
 sg13g2_inv_1 _2412_ (.Y(_1477_),
    .A(net659));
 sg13g2_inv_1 _2413_ (.Y(_1478_),
    .A(net992));
 sg13g2_inv_1 _2414_ (.Y(_1479_),
    .A(_0118_));
 sg13g2_inv_1 _2415_ (.Y(_1480_),
    .A(net673));
 sg13g2_inv_1 _2416_ (.Y(_1481_),
    .A(net635));
 sg13g2_inv_2 _2417_ (.Y(_1482_),
    .A(net662));
 sg13g2_inv_1 _2418_ (.Y(_1483_),
    .A(_0119_));
 sg13g2_inv_1 _2419_ (.Y(_1484_),
    .A(\systolic_array.genblk1[2].accumulators_dlygate[7].A ));
 sg13g2_inv_1 _2420_ (.Y(_1485_),
    .A(net896));
 sg13g2_inv_1 _2421_ (.Y(_1486_),
    .A(net963));
 sg13g2_inv_1 _2422_ (.Y(_1487_),
    .A(net849));
 sg13g2_inv_1 _2423_ (.Y(_1488_),
    .A(net887));
 sg13g2_inv_1 _2424_ (.Y(_1489_),
    .A(net656));
 sg13g2_inv_1 _2425_ (.Y(_1490_),
    .A(_0096_));
 sg13g2_inv_1 _2426_ (.Y(_1491_),
    .A(_0097_));
 sg13g2_inv_1 _2427_ (.Y(_1492_),
    .A(net964));
 sg13g2_inv_2 _2428_ (.Y(_1493_),
    .A(\systolic_array.genblk2[0].mac[2].sign ));
 sg13g2_inv_1 _2429_ (.Y(_1494_),
    .A(_0098_));
 sg13g2_inv_1 _2430_ (.Y(_1495_),
    .A(net874));
 sg13g2_inv_1 _2431_ (.Y(_1496_),
    .A(net854));
 sg13g2_inv_1 _2432_ (.Y(_1497_),
    .A(net845));
 sg13g2_inv_1 _2433_ (.Y(_1498_),
    .A(net654));
 sg13g2_inv_1 _2434_ (.Y(_1499_),
    .A(_0103_));
 sg13g2_inv_2 _2435_ (.Y(_1500_),
    .A(net668));
 sg13g2_inv_1 _2436_ (.Y(_1501_),
    .A(net633));
 sg13g2_inv_2 _2437_ (.Y(_1502_),
    .A(net951));
 sg13g2_inv_1 _2438_ (.Y(_1503_),
    .A(net923));
 sg13g2_inv_1 _2439_ (.Y(_1504_),
    .A(net881));
 sg13g2_inv_1 _2440_ (.Y(_1505_),
    .A(\systolic_array.genblk1[6].accumulators_dlygate[3].A ));
 sg13g2_inv_1 _2441_ (.Y(_1506_),
    .A(net652));
 sg13g2_inv_1 _2442_ (.Y(_1507_),
    .A(_0106_));
 sg13g2_inv_1 _2443_ (.Y(_1508_),
    .A(_0107_));
 sg13g2_inv_2 _2444_ (.Y(_1509_),
    .A(net665));
 sg13g2_inv_2 _2445_ (.Y(_1510_),
    .A(net980));
 sg13g2_inv_1 _2446_ (.Y(_1511_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[6].A ));
 sg13g2_inv_1 _2447_ (.Y(_1512_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[4].A ));
 sg13g2_inv_1 _2448_ (.Y(_1513_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[3].A ));
 sg13g2_inv_1 _2449_ (.Y(_1514_),
    .A(net974));
 sg13g2_inv_1 _2450_ (.Y(_1515_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[10].A ));
 sg13g2_inv_1 _2451_ (.Y(_1516_),
    .A(_0110_));
 sg13g2_inv_1 _2452_ (.Y(_1517_),
    .A(\systolic_array.genblk2[0].mac[5].sign ));
 sg13g2_inv_1 _2453_ (.Y(_1518_),
    .A(_0111_));
 sg13g2_inv_1 _2454_ (.Y(_1519_),
    .A(\systolic_array.genblk1[10].accumulators_dlygate[6].A ));
 sg13g2_inv_1 _2455_ (.Y(_1520_),
    .A(net858));
 sg13g2_inv_1 _2456_ (.Y(_1521_),
    .A(net649));
 sg13g2_inv_1 _2457_ (.Y(_1522_),
    .A(_0113_));
 sg13g2_inv_1 _2458_ (.Y(_1523_),
    .A(net782));
 sg13g2_inv_1 _2459_ (.Y(_1524_),
    .A(net525));
 sg13g2_inv_1 _2460_ (.Y(_1525_),
    .A(net531));
 sg13g2_inv_1 _2461_ (.Y(_1526_),
    .A(net532));
 sg13g2_inv_1 _2462_ (.Y(_1527_),
    .A(net759));
 sg13g2_inv_1 _2463_ (.Y(_1528_),
    .A(net756));
 sg13g2_inv_1 _2464_ (.Y(_1529_),
    .A(net517));
 sg13g2_inv_1 _2465_ (.Y(_1530_),
    .A(net535));
 sg13g2_inv_1 _2466_ (.Y(_1531_),
    .A(net408));
 sg13g2_nand2_2 _2467_ (.Y(_1532_),
    .A(net709),
    .B(net711));
 sg13g2_and2_1 _2468_ (.A(net712),
    .B(net711),
    .X(_1533_));
 sg13g2_nand2_1 _2469_ (.Y(_1534_),
    .A(net712),
    .B(net3));
 sg13g2_and2_1 _2470_ (.A(net709),
    .B(_1533_),
    .X(_1535_));
 sg13g2_nor2_2 _2471_ (.A(net696),
    .B(_1463_),
    .Y(_1536_));
 sg13g2_nand2_1 _2472_ (.Y(_1537_),
    .A(net702),
    .B(net707));
 sg13g2_nor2_1 _2473_ (.A(_1461_),
    .B(net694),
    .Y(_1538_));
 sg13g2_nand2_1 _2474_ (.Y(_1539_),
    .A(net712),
    .B(net714));
 sg13g2_nand4_1 _2475_ (.B(_1535_),
    .C(_1536_),
    .A(net714),
    .Y(_1540_),
    .D(_1538_));
 sg13g2_and2_1 _2476_ (.A(net1),
    .B(_1540_),
    .X(_1541_));
 sg13g2_nand2_2 _2477_ (.Y(_1542_),
    .A(net1),
    .B(_1540_));
 sg13g2_nand2b_1 _2478_ (.Y(_1543_),
    .B(net674),
    .A_N(net681));
 sg13g2_mux2_1 _2479_ (.A0(net680),
    .A1(\systolic_array.arg_top_curr[6] ),
    .S(net636),
    .X(_1544_));
 sg13g2_o21ai_1 _2480_ (.B1(_1543_),
    .Y(_1545_),
    .A1(net676),
    .A2(_1544_));
 sg13g2_nand2b_1 _2481_ (.Y(_1546_),
    .B(net674),
    .A_N(net687));
 sg13g2_mux2_1 _2482_ (.A0(net683),
    .A1(net681),
    .S(net636),
    .X(_1547_));
 sg13g2_o21ai_1 _2483_ (.B1(_1546_),
    .Y(_1548_),
    .A1(net675),
    .A2(_1547_));
 sg13g2_nor2b_1 _2484_ (.A(net690),
    .B_N(\systolic_array.genblk2[0].mac[0].div2 ),
    .Y(_1549_));
 sg13g2_nor2_1 _2485_ (.A(net636),
    .B(net692),
    .Y(_1550_));
 sg13g2_or3_2 _2486_ (.A(net675),
    .B(_1549_),
    .C(_1550_),
    .X(_1551_));
 sg13g2_nand2b_1 _2487_ (.Y(_1552_),
    .B(net674),
    .A_N(net692));
 sg13g2_mux2_1 _2488_ (.A0(net690),
    .A1(net686),
    .S(net636),
    .X(_1553_));
 sg13g2_o21ai_1 _2489_ (.B1(_1552_),
    .Y(_1554_),
    .A1(net674),
    .A2(_1553_));
 sg13g2_nand2b_1 _2490_ (.Y(_1555_),
    .B(net674),
    .A_N(net690));
 sg13g2_mux2_1 _2491_ (.A0(net686),
    .A1(net683),
    .S(net636),
    .X(_1556_));
 sg13g2_o21ai_1 _2492_ (.B1(_1555_),
    .Y(_1557_),
    .A1(net675),
    .A2(_1556_));
 sg13g2_nand3_1 _2493_ (.B(_1554_),
    .C(_1557_),
    .A(_1551_),
    .Y(_1558_));
 sg13g2_and4_1 _2494_ (.A(_1548_),
    .B(_1551_),
    .C(_1554_),
    .D(_1557_),
    .X(_1559_));
 sg13g2_nand4_1 _2495_ (.B(_1551_),
    .C(_1554_),
    .A(_1548_),
    .Y(_1560_),
    .D(_1557_));
 sg13g2_nand2b_1 _2496_ (.Y(_1561_),
    .B(net674),
    .A_N(net684));
 sg13g2_mux2_1 _2497_ (.A0(net681),
    .A1(net680),
    .S(net636),
    .X(_1562_));
 sg13g2_o21ai_1 _2498_ (.B1(_1561_),
    .Y(_1563_),
    .A1(net675),
    .A2(_1562_));
 sg13g2_and2_1 _2499_ (.A(_1545_),
    .B(_1563_),
    .X(_1564_));
 sg13g2_nand2b_1 _2500_ (.Y(_1565_),
    .B(\systolic_array.arg_top_curr[6] ),
    .A_N(net636));
 sg13g2_a21oi_1 _2501_ (.A1(net678),
    .A2(net636),
    .Y(_1566_),
    .B1(net674));
 sg13g2_a22oi_1 _2502_ (.Y(_1567_),
    .B1(_1565_),
    .B2(_1566_),
    .A2(_1468_),
    .A1(net674));
 sg13g2_inv_1 _2503_ (.Y(_1568_),
    .A(_1567_));
 sg13g2_nand3_1 _2504_ (.B(_1564_),
    .C(_1568_),
    .A(_1559_),
    .Y(_1569_));
 sg13g2_nand2_1 _2505_ (.Y(_1570_),
    .A(_0116_),
    .B(net676));
 sg13g2_o21ai_1 _2506_ (.B1(_1570_),
    .Y(_1571_),
    .A1(_1467_),
    .A2(net676));
 sg13g2_nand4_1 _2507_ (.B(_1564_),
    .C(_1568_),
    .A(_1559_),
    .Y(_1572_),
    .D(_1571_));
 sg13g2_nor2_1 _2508_ (.A(net678),
    .B(\systolic_array.genblk2[0].mac[0].sign ),
    .Y(_1573_));
 sg13g2_a22oi_1 _2509_ (.Y(_1574_),
    .B1(_1572_),
    .B2(_1573_),
    .A2(\systolic_array.genblk2[0].mac[0].sign ),
    .A1(_1467_));
 sg13g2_nand2b_1 _2510_ (.Y(_1575_),
    .B(net559),
    .A_N(_0114_));
 sg13g2_xor2_1 _2511_ (.B(net559),
    .A(_0114_),
    .X(_1576_));
 sg13g2_or3_2 _2512_ (.A(_1465_),
    .B(\systolic_array.genblk2[0].mac[0].sign ),
    .C(_1572_),
    .X(_1577_));
 sg13g2_nand3_1 _2513_ (.B(net559),
    .C(_1577_),
    .A(\systolic_array.genblk1[0].accumulators_dlygate[8].A ),
    .Y(_1578_));
 sg13g2_a21oi_1 _2514_ (.A1(_1559_),
    .A2(_1563_),
    .Y(_1579_),
    .B1(\systolic_array.genblk2[0].mac[0].sign ));
 sg13g2_xnor2_1 _2515_ (.Y(_1580_),
    .A(_1545_),
    .B(_1579_));
 sg13g2_nand2_1 _2516_ (.Y(_1581_),
    .A(_1474_),
    .B(_1580_));
 sg13g2_xnor2_1 _2517_ (.Y(_1582_),
    .A(_1474_),
    .B(_1580_));
 sg13g2_nand2_1 _2518_ (.Y(_1583_),
    .A(_1471_),
    .B(_1558_));
 sg13g2_xnor2_1 _2519_ (.Y(_1584_),
    .A(_1548_),
    .B(_1583_));
 sg13g2_nor2_1 _2520_ (.A(\systolic_array.genblk1[0].accumulators_dlygate[3].A ),
    .B(_1584_),
    .Y(_1585_));
 sg13g2_a21oi_1 _2521_ (.A1(_1551_),
    .A2(_1554_),
    .Y(_1586_),
    .B1(\systolic_array.genblk2[0].mac[0].sign ));
 sg13g2_xor2_1 _2522_ (.B(_1586_),
    .A(_1557_),
    .X(_1587_));
 sg13g2_and2_1 _2523_ (.A(\systolic_array.genblk1[0].accumulators_dlygate[2].A ),
    .B(_1587_),
    .X(_1588_));
 sg13g2_or4_1 _2524_ (.A(net676),
    .B(\systolic_array.genblk2[0].mac[0].sign ),
    .C(_1549_),
    .D(_1550_),
    .X(_1589_));
 sg13g2_xor2_1 _2525_ (.B(_1589_),
    .A(_1554_),
    .X(_1590_));
 sg13g2_nand2b_1 _2526_ (.Y(_1591_),
    .B(\systolic_array.genblk1[0].accumulators_dlygate[1].A ),
    .A_N(_1590_));
 sg13g2_nor2_1 _2527_ (.A(\systolic_array.genblk1[0].accumulators_dlygate[0].A ),
    .B(_1551_),
    .Y(_1592_));
 sg13g2_and2_1 _2528_ (.A(_1476_),
    .B(_1590_),
    .X(_1593_));
 sg13g2_xnor2_1 _2529_ (.Y(_1594_),
    .A(\systolic_array.genblk1[0].accumulators_dlygate[1].A ),
    .B(_1590_));
 sg13g2_o21ai_1 _2530_ (.B1(_1591_),
    .Y(_1595_),
    .A1(_1592_),
    .A2(_1593_));
 sg13g2_or2_1 _2531_ (.X(_1596_),
    .B(_1587_),
    .A(\systolic_array.genblk1[0].accumulators_dlygate[2].A ));
 sg13g2_nand2b_1 _2532_ (.Y(_1597_),
    .B(_1596_),
    .A_N(_1588_));
 sg13g2_a21oi_1 _2533_ (.A1(_1595_),
    .A2(_1596_),
    .Y(_1598_),
    .B1(_1588_));
 sg13g2_a221oi_1 _2534_ (.B2(_1596_),
    .C1(_1588_),
    .B1(_1595_),
    .A1(\systolic_array.genblk1[0].accumulators_dlygate[3].A ),
    .Y(_1599_),
    .A2(_1584_));
 sg13g2_nor2_1 _2535_ (.A(_1585_),
    .B(_1599_),
    .Y(_1600_));
 sg13g2_nand3_1 _2536_ (.B(_1560_),
    .C(_1563_),
    .A(_1471_),
    .Y(_1601_));
 sg13g2_a21o_1 _2537_ (.A2(_1560_),
    .A1(_1471_),
    .B1(_1563_),
    .X(_1602_));
 sg13g2_nand2_1 _2538_ (.Y(_1603_),
    .A(_1601_),
    .B(_1602_));
 sg13g2_nor2_1 _2539_ (.A(_1475_),
    .B(_1603_),
    .Y(_1604_));
 sg13g2_nand3_1 _2540_ (.B(_1601_),
    .C(_1602_),
    .A(\systolic_array.genblk1[0].accumulators_dlygate[4].A ),
    .Y(_1605_));
 sg13g2_nand2_1 _2541_ (.Y(_1606_),
    .A(_1475_),
    .B(_1603_));
 sg13g2_xnor2_1 _2542_ (.Y(_1607_),
    .A(_1475_),
    .B(_1603_));
 sg13g2_or4_1 _2543_ (.A(_1582_),
    .B(_1585_),
    .C(_1599_),
    .D(_1607_),
    .X(_1608_));
 sg13g2_and3_1 _2544_ (.X(_1609_),
    .A(_1471_),
    .B(_1569_),
    .C(_1571_));
 sg13g2_a21oi_1 _2545_ (.A1(_1471_),
    .A2(_1569_),
    .Y(_1610_),
    .B1(_1571_));
 sg13g2_nor2_1 _2546_ (.A(_1609_),
    .B(_1610_),
    .Y(_1611_));
 sg13g2_nor2_1 _2547_ (.A(\systolic_array.genblk1[0].accumulators_dlygate[7].A ),
    .B(_1611_),
    .Y(_1612_));
 sg13g2_o21ai_1 _2548_ (.B1(_1473_),
    .Y(_1613_),
    .A1(_1609_),
    .A2(_1610_));
 sg13g2_a21oi_1 _2549_ (.A1(_1559_),
    .A2(_1564_),
    .Y(_1614_),
    .B1(\systolic_array.genblk2[0].mac[0].sign ));
 sg13g2_xnor2_1 _2550_ (.Y(_1615_),
    .A(_1567_),
    .B(_1614_));
 sg13g2_and2_1 _2551_ (.A(\systolic_array.genblk1[0].accumulators_dlygate[6].A ),
    .B(_1615_),
    .X(_1616_));
 sg13g2_o21ai_1 _2552_ (.B1(_1605_),
    .Y(_1617_),
    .A1(_1474_),
    .A2(_1580_));
 sg13g2_nand2_1 _2553_ (.Y(_1618_),
    .A(_1581_),
    .B(_1617_));
 sg13g2_nor3_1 _2554_ (.A(_1473_),
    .B(_1609_),
    .C(_1610_),
    .Y(_1619_));
 sg13g2_nand2_1 _2555_ (.Y(_1620_),
    .A(\systolic_array.genblk1[0].accumulators_dlygate[7].A ),
    .B(_1611_));
 sg13g2_a221oi_1 _2556_ (.B2(_1581_),
    .C1(_1619_),
    .B1(_1617_),
    .A1(_1613_),
    .Y(_1621_),
    .A2(_1616_));
 sg13g2_nor2_1 _2557_ (.A(\systolic_array.genblk1[0].accumulators_dlygate[6].A ),
    .B(_1615_),
    .Y(_1622_));
 sg13g2_a221oi_1 _2558_ (.B2(_1620_),
    .C1(_1612_),
    .B1(_1622_),
    .A1(_1608_),
    .Y(_1623_),
    .A2(_1621_));
 sg13g2_inv_1 _2559_ (.Y(_1624_),
    .A(_1623_));
 sg13g2_a21o_1 _2560_ (.A2(_1577_),
    .A1(net559),
    .B1(\systolic_array.genblk1[0].accumulators_dlygate[8].A ),
    .X(_1625_));
 sg13g2_nand2_2 _2561_ (.Y(_1626_),
    .A(_1578_),
    .B(_1625_));
 sg13g2_o21ai_1 _2562_ (.B1(_1578_),
    .Y(_1627_),
    .A1(_1624_),
    .A2(_1626_));
 sg13g2_xnor2_1 _2563_ (.Y(_1628_),
    .A(_1576_),
    .B(_1627_));
 sg13g2_mux2_1 _2564_ (.A0(net952),
    .A1(_1628_),
    .S(net630),
    .X(_1629_));
 sg13g2_mux2_1 _2565_ (.A0(net521),
    .A1(_1629_),
    .S(net603),
    .X(_0015_));
 sg13g2_nor2_1 _2566_ (.A(net732),
    .B(net603),
    .Y(_1630_));
 sg13g2_and2_1 _2567_ (.A(_1575_),
    .B(_1578_),
    .X(_1631_));
 sg13g2_inv_1 _2568_ (.Y(_1632_),
    .A(_1631_));
 sg13g2_nor2_1 _2569_ (.A(_1576_),
    .B(_1626_),
    .Y(_1633_));
 sg13g2_a21oi_1 _2570_ (.A1(_1623_),
    .A2(_1633_),
    .Y(_1634_),
    .B1(_1632_));
 sg13g2_nand2_1 _2571_ (.Y(_1635_),
    .A(\systolic_array.genblk1[0].accumulators_dlygate[10].A ),
    .B(_1574_));
 sg13g2_xnor2_1 _2572_ (.Y(_1636_),
    .A(\systolic_array.genblk1[0].accumulators_dlygate[10].A ),
    .B(_1574_));
 sg13g2_or2_1 _2573_ (.X(_1637_),
    .B(_1636_),
    .A(_1634_));
 sg13g2_a21oi_1 _2574_ (.A1(_1634_),
    .A2(_1636_),
    .Y(_1638_),
    .B1(net660));
 sg13g2_a22oi_1 _2575_ (.Y(_1639_),
    .B1(_1637_),
    .B2(_1638_),
    .A2(net979),
    .A1(net660));
 sg13g2_a21oi_1 _2576_ (.A1(net603),
    .A2(_1639_),
    .Y(_0008_),
    .B1(_1630_));
 sg13g2_nand2b_1 _2577_ (.Y(_1640_),
    .B(_1574_),
    .A_N(_0117_));
 sg13g2_xor2_1 _2578_ (.B(net559),
    .A(_0117_),
    .X(_1641_));
 sg13g2_o21ai_1 _2579_ (.B1(_1635_),
    .Y(_1642_),
    .A1(_1634_),
    .A2(_1636_));
 sg13g2_xnor2_1 _2580_ (.Y(_1643_),
    .A(_1641_),
    .B(_1642_));
 sg13g2_mux2_1 _2581_ (.A0(net962),
    .A1(_1643_),
    .S(net630),
    .X(_1644_));
 sg13g2_mux2_1 _2582_ (.A0(net523),
    .A1(_1644_),
    .S(net603),
    .X(_0009_));
 sg13g2_nand3_1 _2583_ (.B(_1635_),
    .C(_1640_),
    .A(_1631_),
    .Y(_1645_));
 sg13g2_nor4_2 _2584_ (.A(_1576_),
    .B(_1626_),
    .C(_1636_),
    .Y(_1646_),
    .D(_1641_));
 sg13g2_nand2_1 _2585_ (.Y(_1647_),
    .A(_1623_),
    .B(_1646_));
 sg13g2_a21oi_2 _2586_ (.B1(_1645_),
    .Y(_1648_),
    .A2(_1646_),
    .A1(_1623_));
 sg13g2_nand2_1 _2587_ (.Y(_1649_),
    .A(\systolic_array.genblk1[0].accumulators_dlygate[12].A ),
    .B(net559));
 sg13g2_xnor2_1 _2588_ (.Y(_1650_),
    .A(\systolic_array.genblk1[0].accumulators_dlygate[12].A ),
    .B(net558));
 sg13g2_a21oi_1 _2589_ (.A1(_1648_),
    .A2(_1650_),
    .Y(_1651_),
    .B1(net659));
 sg13g2_o21ai_1 _2590_ (.B1(_1651_),
    .Y(_1652_),
    .A1(_1648_),
    .A2(_1650_));
 sg13g2_o21ai_1 _2591_ (.B1(_1652_),
    .Y(_1653_),
    .A1(net630),
    .A2(_1478_));
 sg13g2_mux2_1 _2592_ (.A0(net526),
    .A1(_1653_),
    .S(net605),
    .X(_0010_));
 sg13g2_xnor2_1 _2593_ (.Y(_1654_),
    .A(_0118_),
    .B(net559));
 sg13g2_o21ai_1 _2594_ (.B1(_1649_),
    .Y(_1655_),
    .A1(_1648_),
    .A2(_1650_));
 sg13g2_xor2_1 _2595_ (.B(_1655_),
    .A(_1654_),
    .X(_1656_));
 sg13g2_mux2_1 _2596_ (.A0(net981),
    .A1(_1656_),
    .S(net630),
    .X(_1657_));
 sg13g2_mux2_1 _2597_ (.A0(net734),
    .A1(_1657_),
    .S(net605),
    .X(_0011_));
 sg13g2_nor2_1 _2598_ (.A(net528),
    .B(net603),
    .Y(_1658_));
 sg13g2_o21ai_1 _2599_ (.B1(net558),
    .Y(_1659_),
    .A1(\systolic_array.genblk1[0].accumulators_dlygate[12].A ),
    .A2(_1479_));
 sg13g2_nand2b_1 _2600_ (.Y(_1660_),
    .B(_1654_),
    .A_N(_1650_));
 sg13g2_o21ai_1 _2601_ (.B1(_1659_),
    .Y(_1661_),
    .A1(_1648_),
    .A2(_1660_));
 sg13g2_xnor2_1 _2602_ (.Y(_1662_),
    .A(\systolic_array.genblk1[0].accumulators_dlygate[14].A ),
    .B(net558));
 sg13g2_nor2b_1 _2603_ (.A(_1662_),
    .B_N(_1661_),
    .Y(_1663_));
 sg13g2_nor2b_1 _2604_ (.A(_1661_),
    .B_N(_1662_),
    .Y(_1664_));
 sg13g2_nor3_1 _2605_ (.A(net659),
    .B(_1663_),
    .C(_1664_),
    .Y(_0401_));
 sg13g2_a21oi_1 _2606_ (.A1(net659),
    .A2(net984),
    .Y(_0402_),
    .B1(_0401_));
 sg13g2_a21oi_1 _2607_ (.A1(net603),
    .A2(_0402_),
    .Y(_0012_),
    .B1(_1658_));
 sg13g2_nand2b_1 _2608_ (.Y(_0403_),
    .B(net659),
    .A_N(net987));
 sg13g2_xnor2_1 _2609_ (.Y(_0404_),
    .A(\systolic_array.genblk1[0].accumulators_dlygate[15].A ),
    .B(net558));
 sg13g2_a21o_1 _2610_ (.A2(net558),
    .A1(\systolic_array.genblk1[0].accumulators_dlygate[14].A ),
    .B1(_1663_),
    .X(_0405_));
 sg13g2_xnor2_1 _2611_ (.Y(_0406_),
    .A(_0404_),
    .B(_0405_));
 sg13g2_o21ai_1 _2612_ (.B1(_0403_),
    .Y(_0407_),
    .A1(net659),
    .A2(_0406_));
 sg13g2_nor2_1 _2613_ (.A(net842),
    .B(net604),
    .Y(_0408_));
 sg13g2_a21oi_1 _2614_ (.A1(net603),
    .A2(_0407_),
    .Y(_0013_),
    .B1(_0408_));
 sg13g2_nor2_1 _2615_ (.A(net785),
    .B(net604),
    .Y(_0409_));
 sg13g2_nor4_1 _2616_ (.A(_1647_),
    .B(_1660_),
    .C(_1662_),
    .D(_0404_),
    .Y(_0410_));
 sg13g2_o21ai_1 _2617_ (.B1(net558),
    .Y(_0411_),
    .A1(\systolic_array.genblk1[0].accumulators_dlygate[14].A ),
    .A2(\systolic_array.genblk1[0].accumulators_dlygate[15].A ));
 sg13g2_nand2_1 _2618_ (.Y(_0412_),
    .A(_1659_),
    .B(_0411_));
 sg13g2_nor3_1 _2619_ (.A(_1645_),
    .B(_0410_),
    .C(_0412_),
    .Y(_0413_));
 sg13g2_nor2b_1 _2620_ (.A(net558),
    .B_N(_0413_),
    .Y(_0414_));
 sg13g2_nor2b_1 _2621_ (.A(_0413_),
    .B_N(net558),
    .Y(_0415_));
 sg13g2_nor3_1 _2622_ (.A(net659),
    .B(_0414_),
    .C(_0415_),
    .Y(_0416_));
 sg13g2_xnor2_1 _2623_ (.Y(_0417_),
    .A(net895),
    .B(_0416_));
 sg13g2_a21oi_1 _2624_ (.A1(net604),
    .A2(_0417_),
    .Y(_0014_),
    .B1(_0409_));
 sg13g2_mux2_1 _2625_ (.A0(net508),
    .A1(net847),
    .S(net615),
    .X(_0031_));
 sg13g2_mux2_1 _2626_ (.A0(net481),
    .A1(net813),
    .S(net615),
    .X(_0024_));
 sg13g2_mux2_1 _2627_ (.A0(net484),
    .A1(net834),
    .S(net615),
    .X(_0025_));
 sg13g2_mux2_1 _2628_ (.A0(net440),
    .A1(net776),
    .S(net613),
    .X(_0026_));
 sg13g2_mux2_1 _2629_ (.A0(net447),
    .A1(net850),
    .S(net615),
    .X(_0027_));
 sg13g2_mux2_1 _2630_ (.A0(net478),
    .A1(net805),
    .S(net613),
    .X(_0028_));
 sg13g2_mux2_1 _2631_ (.A0(net439),
    .A1(net790),
    .S(net613),
    .X(_0029_));
 sg13g2_mux2_1 _2632_ (.A0(net510),
    .A1(net811),
    .S(net613),
    .X(_0030_));
 sg13g2_nand2b_1 _2633_ (.Y(_0418_),
    .B(net671),
    .A_N(net686));
 sg13g2_mux2_1 _2634_ (.A0(net683),
    .A1(net681),
    .S(net634),
    .X(_0419_));
 sg13g2_o21ai_1 _2635_ (.B1(_0418_),
    .Y(_0420_),
    .A1(net671),
    .A2(_0419_));
 sg13g2_nor2b_1 _2636_ (.A(net689),
    .B_N(net634),
    .Y(_0421_));
 sg13g2_nor2_1 _2637_ (.A(net692),
    .B(net634),
    .Y(_0422_));
 sg13g2_or3_2 _2638_ (.A(net672),
    .B(_0421_),
    .C(_0422_),
    .X(_0423_));
 sg13g2_nand2b_1 _2639_ (.Y(_0424_),
    .B(net671),
    .A_N(net692));
 sg13g2_mux2_1 _2640_ (.A0(net689),
    .A1(net686),
    .S(net634),
    .X(_0425_));
 sg13g2_o21ai_1 _2641_ (.B1(_0424_),
    .Y(_0426_),
    .A1(net671),
    .A2(_0425_));
 sg13g2_nand2b_1 _2642_ (.Y(_0427_),
    .B(net671),
    .A_N(net689));
 sg13g2_mux2_1 _2643_ (.A0(net686),
    .A1(net683),
    .S(net634),
    .X(_0428_));
 sg13g2_o21ai_1 _2644_ (.B1(_0427_),
    .Y(_0429_),
    .A1(net671),
    .A2(_0428_));
 sg13g2_nand3_1 _2645_ (.B(_0426_),
    .C(_0429_),
    .A(_0423_),
    .Y(_0430_));
 sg13g2_and4_1 _2646_ (.A(_0420_),
    .B(_0423_),
    .C(_0426_),
    .D(_0429_),
    .X(_0431_));
 sg13g2_nand4_1 _2647_ (.B(_0423_),
    .C(_0426_),
    .A(_0420_),
    .Y(_0432_),
    .D(_0429_));
 sg13g2_nand2b_1 _2648_ (.Y(_0433_),
    .B(net673),
    .A_N(net683));
 sg13g2_nand2_1 _2649_ (.Y(_0434_),
    .A(net679),
    .B(net635));
 sg13g2_o21ai_1 _2650_ (.B1(_0434_),
    .Y(_0435_),
    .A1(_1469_),
    .A2(net635));
 sg13g2_o21ai_1 _2651_ (.B1(_0433_),
    .Y(_0436_),
    .A1(net673),
    .A2(_0435_));
 sg13g2_mux2_1 _2652_ (.A0(net683),
    .A1(_0435_),
    .S(_1480_),
    .X(_0437_));
 sg13g2_nand2b_1 _2653_ (.Y(_0438_),
    .B(net679),
    .A_N(net634));
 sg13g2_a21oi_1 _2654_ (.A1(\systolic_array.arg_top_curr[6] ),
    .A2(net634),
    .Y(_0439_),
    .B1(net672));
 sg13g2_a22oi_1 _2655_ (.Y(_0440_),
    .B1(_0438_),
    .B2(_0439_),
    .A2(net671),
    .A1(_1469_));
 sg13g2_inv_1 _2656_ (.Y(_0441_),
    .A(_0440_));
 sg13g2_nor3_1 _2657_ (.A(_0432_),
    .B(_0437_),
    .C(_0440_),
    .Y(_0442_));
 sg13g2_nand2_1 _2658_ (.Y(_0443_),
    .A(_1465_),
    .B(net634));
 sg13g2_a21oi_1 _2659_ (.A1(_1466_),
    .A2(_1481_),
    .Y(_0444_),
    .B1(net671));
 sg13g2_a22oi_1 _2660_ (.Y(_0445_),
    .B1(_0443_),
    .B2(_0444_),
    .A2(net672),
    .A1(net679));
 sg13g2_and4_1 _2661_ (.A(_0431_),
    .B(_0436_),
    .C(_0441_),
    .D(_0445_),
    .X(_0446_));
 sg13g2_nand4_1 _2662_ (.B(_0436_),
    .C(_0441_),
    .A(_0431_),
    .Y(_0447_),
    .D(_0445_));
 sg13g2_nor2_1 _2663_ (.A(_0115_),
    .B(net673),
    .Y(_0448_));
 sg13g2_nand2b_1 _2664_ (.Y(_0449_),
    .B(net673),
    .A_N(_0116_));
 sg13g2_nor2b_1 _2665_ (.A(_0448_),
    .B_N(_0449_),
    .Y(_0450_));
 sg13g2_nand2b_1 _2666_ (.Y(_0451_),
    .B(_0449_),
    .A_N(_0448_));
 sg13g2_nor2_1 _2667_ (.A(net678),
    .B(\systolic_array.genblk2[0].mac[1].sign ),
    .Y(_0452_));
 sg13g2_o21ai_1 _2668_ (.B1(_0452_),
    .Y(_0453_),
    .A1(_0447_),
    .A2(_0451_));
 sg13g2_nand2_1 _2669_ (.Y(_0454_),
    .A(_1467_),
    .B(\systolic_array.genblk2[0].mac[1].sign ));
 sg13g2_and2_1 _2670_ (.A(_0453_),
    .B(_0454_),
    .X(_0455_));
 sg13g2_xnor2_1 _2671_ (.Y(_0456_),
    .A(_1483_),
    .B(_0455_));
 sg13g2_nand4_1 _2672_ (.B(_1482_),
    .C(_0446_),
    .A(net677),
    .Y(_0457_),
    .D(_0450_));
 sg13g2_nand3_1 _2673_ (.B(_0454_),
    .C(_0457_),
    .A(_0453_),
    .Y(_0458_));
 sg13g2_and4_1 _2674_ (.A(\systolic_array.genblk1[2].accumulators_dlygate[8].A ),
    .B(_0453_),
    .C(_0454_),
    .D(_0457_),
    .X(_0459_));
 sg13g2_a21oi_1 _2675_ (.A1(_0431_),
    .A2(_0436_),
    .Y(_0460_),
    .B1(net662));
 sg13g2_xnor2_1 _2676_ (.Y(_0461_),
    .A(_0441_),
    .B(_0460_));
 sg13g2_nand2_1 _2677_ (.Y(_0462_),
    .A(_1486_),
    .B(_0461_));
 sg13g2_xnor2_1 _2678_ (.Y(_0463_),
    .A(_1486_),
    .B(_0461_));
 sg13g2_nand2_1 _2679_ (.Y(_0464_),
    .A(_1482_),
    .B(_0430_));
 sg13g2_xnor2_1 _2680_ (.Y(_0465_),
    .A(_0420_),
    .B(_0464_));
 sg13g2_nor2_1 _2681_ (.A(\systolic_array.genblk1[2].accumulators_dlygate[3].A ),
    .B(_0465_),
    .Y(_0466_));
 sg13g2_a21oi_1 _2682_ (.A1(_0423_),
    .A2(_0426_),
    .Y(_0467_),
    .B1(net662));
 sg13g2_xor2_1 _2683_ (.B(_0467_),
    .A(_0429_),
    .X(_0468_));
 sg13g2_and2_1 _2684_ (.A(\systolic_array.genblk1[2].accumulators_dlygate[2].A ),
    .B(_0468_),
    .X(_0469_));
 sg13g2_or4_1 _2685_ (.A(net672),
    .B(net662),
    .C(_0421_),
    .D(_0422_),
    .X(_0470_));
 sg13g2_xnor2_1 _2686_ (.Y(_0471_),
    .A(_0426_),
    .B(_0470_));
 sg13g2_nand2_1 _2687_ (.Y(_0472_),
    .A(\systolic_array.genblk1[2].accumulators_dlygate[1].A ),
    .B(_0471_));
 sg13g2_nor2_1 _2688_ (.A(\systolic_array.genblk1[2].accumulators_dlygate[0].A ),
    .B(_0423_),
    .Y(_0473_));
 sg13g2_nor2_1 _2689_ (.A(\systolic_array.genblk1[2].accumulators_dlygate[1].A ),
    .B(_0471_),
    .Y(_0474_));
 sg13g2_xnor2_1 _2690_ (.Y(_0475_),
    .A(_1488_),
    .B(_0471_));
 sg13g2_o21ai_1 _2691_ (.B1(_0472_),
    .Y(_0476_),
    .A1(_0473_),
    .A2(_0474_));
 sg13g2_or2_1 _2692_ (.X(_0477_),
    .B(_0468_),
    .A(\systolic_array.genblk1[2].accumulators_dlygate[2].A ));
 sg13g2_nand2b_1 _2693_ (.Y(_0478_),
    .B(_0477_),
    .A_N(_0469_));
 sg13g2_a21oi_1 _2694_ (.A1(_0476_),
    .A2(_0477_),
    .Y(_0479_),
    .B1(_0469_));
 sg13g2_a221oi_1 _2695_ (.B2(_0477_),
    .C1(_0469_),
    .B1(_0476_),
    .A1(\systolic_array.genblk1[2].accumulators_dlygate[3].A ),
    .Y(_0480_),
    .A2(_0465_));
 sg13g2_nand3_1 _2696_ (.B(_0432_),
    .C(_0436_),
    .A(_1482_),
    .Y(_0481_));
 sg13g2_o21ai_1 _2697_ (.B1(_0437_),
    .Y(_0482_),
    .A1(net662),
    .A2(_0431_));
 sg13g2_nand2_1 _2698_ (.Y(_0483_),
    .A(_0481_),
    .B(_0482_));
 sg13g2_nor2_1 _2699_ (.A(_1487_),
    .B(_0483_),
    .Y(_0484_));
 sg13g2_nand3_1 _2700_ (.B(_0481_),
    .C(_0482_),
    .A(\systolic_array.genblk1[2].accumulators_dlygate[4].A ),
    .Y(_0485_));
 sg13g2_xnor2_1 _2701_ (.Y(_0486_),
    .A(_1487_),
    .B(_0483_));
 sg13g2_nor3_2 _2702_ (.A(_0466_),
    .B(_0480_),
    .C(_0486_),
    .Y(_0487_));
 sg13g2_nor2b_1 _2703_ (.A(_0463_),
    .B_N(_0487_),
    .Y(_0488_));
 sg13g2_or4_1 _2704_ (.A(_0463_),
    .B(_0466_),
    .C(_0480_),
    .D(_0486_),
    .X(_0489_));
 sg13g2_nor3_1 _2705_ (.A(net662),
    .B(_0446_),
    .C(_0451_),
    .Y(_0490_));
 sg13g2_a21oi_1 _2706_ (.A1(_1482_),
    .A2(_0447_),
    .Y(_0491_),
    .B1(_0450_));
 sg13g2_o21ai_1 _2707_ (.B1(_1484_),
    .Y(_0492_),
    .A1(_0490_),
    .A2(_0491_));
 sg13g2_or3_1 _2708_ (.A(net662),
    .B(_0442_),
    .C(_0445_),
    .X(_0493_));
 sg13g2_o21ai_1 _2709_ (.B1(_0445_),
    .Y(_0494_),
    .A1(net662),
    .A2(_0442_));
 sg13g2_nand2_1 _2710_ (.Y(_0495_),
    .A(_0493_),
    .B(_0494_));
 sg13g2_a21oi_1 _2711_ (.A1(_0493_),
    .A2(_0494_),
    .Y(_0496_),
    .B1(_1485_));
 sg13g2_nor3_1 _2712_ (.A(_1484_),
    .B(_0490_),
    .C(_0491_),
    .Y(_0497_));
 sg13g2_or3_1 _2713_ (.A(_1484_),
    .B(_0490_),
    .C(_0491_),
    .X(_0498_));
 sg13g2_o21ai_1 _2714_ (.B1(_0485_),
    .Y(_0499_),
    .A1(_1486_),
    .A2(_0461_));
 sg13g2_and2_1 _2715_ (.A(_0462_),
    .B(_0499_),
    .X(_0500_));
 sg13g2_a221oi_1 _2716_ (.B2(_0462_),
    .C1(_0497_),
    .B1(_0499_),
    .A1(_0492_),
    .Y(_0501_),
    .A2(_0496_));
 sg13g2_o21ai_1 _2717_ (.B1(_0492_),
    .Y(_0502_),
    .A1(\systolic_array.genblk1[2].accumulators_dlygate[6].A ),
    .A2(_0495_));
 sg13g2_a22oi_1 _2718_ (.Y(_0503_),
    .B1(_0502_),
    .B2(_0498_),
    .A2(_0501_),
    .A1(_0489_));
 sg13g2_xor2_1 _2719_ (.B(_0458_),
    .A(\systolic_array.genblk1[2].accumulators_dlygate[8].A ),
    .X(_0504_));
 sg13g2_inv_1 _2720_ (.Y(_0505_),
    .A(_0504_));
 sg13g2_a21oi_1 _2721_ (.A1(_0503_),
    .A2(_0505_),
    .Y(_0506_),
    .B1(_0459_));
 sg13g2_xor2_1 _2722_ (.B(_0506_),
    .A(_0456_),
    .X(_0507_));
 sg13g2_mux2_1 _2723_ (.A0(net953),
    .A1(_0507_),
    .S(net627),
    .X(_0508_));
 sg13g2_mux2_1 _2724_ (.A0(net802),
    .A1(_0508_),
    .S(net602),
    .X(_0039_));
 sg13g2_a21oi_2 _2725_ (.B1(_0459_),
    .Y(_0509_),
    .A2(net551),
    .A1(_1483_));
 sg13g2_nand3b_1 _2726_ (.B(_0503_),
    .C(_0505_),
    .Y(_0510_),
    .A_N(_0456_));
 sg13g2_xnor2_1 _2727_ (.Y(_0511_),
    .A(\systolic_array.genblk1[2].accumulators_dlygate[10].A ),
    .B(net551));
 sg13g2_a21oi_1 _2728_ (.A1(_0509_),
    .A2(_0510_),
    .Y(_0512_),
    .B1(_0511_));
 sg13g2_nand3_1 _2729_ (.B(_0510_),
    .C(_0511_),
    .A(_0509_),
    .Y(_0513_));
 sg13g2_nand2_1 _2730_ (.Y(_0514_),
    .A(net658),
    .B(net990));
 sg13g2_nand2_1 _2731_ (.Y(_0515_),
    .A(net627),
    .B(_0513_));
 sg13g2_o21ai_1 _2732_ (.B1(net991),
    .Y(_0516_),
    .A1(_0512_),
    .A2(_0515_));
 sg13g2_mux2_1 _2733_ (.A0(net765),
    .A1(_0516_),
    .S(net602),
    .X(_0032_));
 sg13g2_xnor2_1 _2734_ (.Y(_0517_),
    .A(_1490_),
    .B(net551));
 sg13g2_a21oi_1 _2735_ (.A1(\systolic_array.genblk1[2].accumulators_dlygate[10].A ),
    .A2(net551),
    .Y(_0518_),
    .B1(_0512_));
 sg13g2_nor2_1 _2736_ (.A(net627),
    .B(net946),
    .Y(_0519_));
 sg13g2_xnor2_1 _2737_ (.Y(_0520_),
    .A(_0517_),
    .B(_0518_));
 sg13g2_a21oi_1 _2738_ (.A1(net627),
    .A2(_0520_),
    .Y(_0521_),
    .B1(_0519_));
 sg13g2_mux2_1 _2739_ (.A0(net722),
    .A1(_0521_),
    .S(net603),
    .X(_0033_));
 sg13g2_nor4_2 _2740_ (.A(_0456_),
    .B(_0504_),
    .C(_0511_),
    .Y(_0522_),
    .D(_0517_));
 sg13g2_nand2_1 _2741_ (.Y(_0523_),
    .A(_0503_),
    .B(_0522_));
 sg13g2_o21ai_1 _2742_ (.B1(net551),
    .Y(_0524_),
    .A1(\systolic_array.genblk1[2].accumulators_dlygate[10].A ),
    .A2(_1490_));
 sg13g2_nand2_1 _2743_ (.Y(_0525_),
    .A(_0509_),
    .B(_0524_));
 sg13g2_a21oi_2 _2744_ (.B1(_0525_),
    .Y(_0526_),
    .A2(_0522_),
    .A1(_0503_));
 sg13g2_xnor2_1 _2745_ (.Y(_0527_),
    .A(\systolic_array.genblk1[2].accumulators_dlygate[12].A ),
    .B(net551));
 sg13g2_nor2_1 _2746_ (.A(_0526_),
    .B(_0527_),
    .Y(_0528_));
 sg13g2_nand2_1 _2747_ (.Y(_0529_),
    .A(net656),
    .B(net994));
 sg13g2_a21o_1 _2748_ (.A2(_0527_),
    .A1(_0526_),
    .B1(net656),
    .X(_0530_));
 sg13g2_o21ai_1 _2749_ (.B1(_0529_),
    .Y(_0531_),
    .A1(_0528_),
    .A2(_0530_));
 sg13g2_mux2_1 _2750_ (.A0(net808),
    .A1(_0531_),
    .S(net604),
    .X(_0034_));
 sg13g2_xnor2_1 _2751_ (.Y(_0532_),
    .A(_0097_),
    .B(net551));
 sg13g2_a21oi_1 _2752_ (.A1(\systolic_array.genblk1[2].accumulators_dlygate[12].A ),
    .A2(net550),
    .Y(_0533_),
    .B1(_0528_));
 sg13g2_xnor2_1 _2753_ (.Y(_0534_),
    .A(_0532_),
    .B(_0533_));
 sg13g2_mux2_1 _2754_ (.A0(net965),
    .A1(_0534_),
    .S(net627),
    .X(_0535_));
 sg13g2_mux2_1 _2755_ (.A0(net763),
    .A1(_0535_),
    .S(net604),
    .X(_0035_));
 sg13g2_nor2_1 _2756_ (.A(net863),
    .B(net601),
    .Y(_0536_));
 sg13g2_and2_1 _2757_ (.A(\systolic_array.genblk1[2].accumulators_dlygate[14].A ),
    .B(net550),
    .X(_0537_));
 sg13g2_xnor2_1 _2758_ (.Y(_0538_),
    .A(\systolic_array.genblk1[2].accumulators_dlygate[14].A ),
    .B(net550));
 sg13g2_inv_1 _2759_ (.Y(_0539_),
    .A(_0538_));
 sg13g2_o21ai_1 _2760_ (.B1(net550),
    .Y(_0540_),
    .A1(\systolic_array.genblk1[2].accumulators_dlygate[12].A ),
    .A2(_1491_));
 sg13g2_nand2b_1 _2761_ (.Y(_0541_),
    .B(_0532_),
    .A_N(_0527_));
 sg13g2_o21ai_1 _2762_ (.B1(_0540_),
    .Y(_0542_),
    .A1(_0526_),
    .A2(_0541_));
 sg13g2_nand2_1 _2763_ (.Y(_0543_),
    .A(_0539_),
    .B(_0542_));
 sg13g2_nor2_1 _2764_ (.A(_0539_),
    .B(_0542_),
    .Y(_0544_));
 sg13g2_nor2_1 _2765_ (.A(net656),
    .B(_0544_),
    .Y(_0545_));
 sg13g2_a22oi_1 _2766_ (.Y(_0546_),
    .B1(_0543_),
    .B2(_0545_),
    .A2(net967),
    .A1(net656));
 sg13g2_a21oi_1 _2767_ (.A1(net602),
    .A2(_0546_),
    .Y(_0036_),
    .B1(_0536_));
 sg13g2_xnor2_1 _2768_ (.Y(_0547_),
    .A(\systolic_array.genblk1[2].accumulators_dlygate[15].A ),
    .B(net550));
 sg13g2_a21oi_1 _2769_ (.A1(_0539_),
    .A2(_0542_),
    .Y(_0548_),
    .B1(_0537_));
 sg13g2_xnor2_1 _2770_ (.Y(_0549_),
    .A(_0547_),
    .B(_0548_));
 sg13g2_nor2_1 _2771_ (.A(net656),
    .B(_0549_),
    .Y(_0550_));
 sg13g2_a21oi_1 _2772_ (.A1(net656),
    .A2(net948),
    .Y(_0551_),
    .B1(_0550_));
 sg13g2_nor2_1 _2773_ (.A(net861),
    .B(net601),
    .Y(_0552_));
 sg13g2_a21oi_1 _2774_ (.A1(net601),
    .A2(_0551_),
    .Y(_0037_),
    .B1(_0552_));
 sg13g2_nor2_1 _2775_ (.A(net744),
    .B(net604),
    .Y(_0553_));
 sg13g2_nor4_1 _2776_ (.A(_0523_),
    .B(_0538_),
    .C(_0541_),
    .D(_0547_),
    .Y(_0554_));
 sg13g2_o21ai_1 _2777_ (.B1(net550),
    .Y(_0555_),
    .A1(\systolic_array.genblk1[2].accumulators_dlygate[14].A ),
    .A2(\systolic_array.genblk1[2].accumulators_dlygate[15].A ));
 sg13g2_nand4_1 _2778_ (.B(_0524_),
    .C(_0540_),
    .A(_0509_),
    .Y(_0556_),
    .D(_0555_));
 sg13g2_nor2_1 _2779_ (.A(_0554_),
    .B(_0556_),
    .Y(_0557_));
 sg13g2_nor3_1 _2780_ (.A(net550),
    .B(_0554_),
    .C(_0556_),
    .Y(_0558_));
 sg13g2_nor2b_1 _2781_ (.A(_0557_),
    .B_N(net550),
    .Y(_0559_));
 sg13g2_nor3_2 _2782_ (.A(net656),
    .B(_0558_),
    .C(_0559_),
    .Y(_0560_));
 sg13g2_xnor2_1 _2783_ (.Y(_0561_),
    .A(net901),
    .B(_0560_));
 sg13g2_a21oi_1 _2784_ (.A1(net604),
    .A2(_0561_),
    .Y(_0038_),
    .B1(_0553_));
 sg13g2_mux2_1 _2785_ (.A0(net498),
    .A1(net801),
    .S(net614),
    .X(_0047_));
 sg13g2_mux2_1 _2786_ (.A0(net456),
    .A1(net789),
    .S(net614),
    .X(_0040_));
 sg13g2_mux2_1 _2787_ (.A0(net467),
    .A1(net812),
    .S(net613),
    .X(_0041_));
 sg13g2_mux2_1 _2788_ (.A0(net488),
    .A1(net867),
    .S(net613),
    .X(_0042_));
 sg13g2_mux2_1 _2789_ (.A0(net490),
    .A1(net784),
    .S(net613),
    .X(_0043_));
 sg13g2_mux2_1 _2790_ (.A0(net469),
    .A1(net795),
    .S(net614),
    .X(_0044_));
 sg13g2_mux2_1 _2791_ (.A0(net492),
    .A1(net815),
    .S(net614),
    .X(_0045_));
 sg13g2_mux2_1 _2792_ (.A0(net479),
    .A1(net783),
    .S(net613),
    .X(_0046_));
 sg13g2_nor2_1 _2793_ (.A(_1467_),
    .B(_1493_),
    .Y(_0562_));
 sg13g2_nand2b_1 _2794_ (.Y(_0563_),
    .B(net689),
    .A_N(net670));
 sg13g2_nor2b_1 _2795_ (.A(net670),
    .B_N(net686),
    .Y(_0564_));
 sg13g2_a21o_1 _2796_ (.A2(net669),
    .A1(net689),
    .B1(_0564_),
    .X(_0565_));
 sg13g2_nor3_1 _2797_ (.A(net689),
    .B(net692),
    .C(_0564_),
    .Y(_0566_));
 sg13g2_nor2b_1 _2798_ (.A(net670),
    .B_N(net683),
    .Y(_0567_));
 sg13g2_a21oi_1 _2799_ (.A1(net686),
    .A2(net670),
    .Y(_0568_),
    .B1(_0567_));
 sg13g2_nor4_2 _2800_ (.A(net686),
    .B(net689),
    .C(net692),
    .Y(_0569_),
    .D(_0567_));
 sg13g2_nand2b_1 _2801_ (.Y(_0570_),
    .B(net669),
    .A_N(net683));
 sg13g2_o21ai_1 _2802_ (.B1(_0570_),
    .Y(_0571_),
    .A1(\systolic_array.arg_top_curr[4] ),
    .A2(net669));
 sg13g2_mux2_1 _2803_ (.A0(net680),
    .A1(\systolic_array.arg_top_curr[4] ),
    .S(net669),
    .X(_0572_));
 sg13g2_inv_1 _2804_ (.Y(_0573_),
    .A(_0572_));
 sg13g2_nand3_1 _2805_ (.B(_0571_),
    .C(_0573_),
    .A(_0569_),
    .Y(_0574_));
 sg13g2_mux2_1 _2806_ (.A0(_0116_),
    .A1(_0099_),
    .S(net669),
    .X(_0575_));
 sg13g2_nand4_1 _2807_ (.B(_0571_),
    .C(_0573_),
    .A(_0569_),
    .Y(_0576_),
    .D(_0575_));
 sg13g2_nor2_1 _2808_ (.A(net678),
    .B(net669),
    .Y(_0577_));
 sg13g2_a21oi_2 _2809_ (.B1(_0577_),
    .Y(_0578_),
    .A2(net669),
    .A1(_1466_));
 sg13g2_o21ai_1 _2810_ (.B1(_1465_),
    .Y(_0579_),
    .A1(_0576_),
    .A2(_0578_));
 sg13g2_a21o_1 _2811_ (.A2(_0579_),
    .A1(_1493_),
    .B1(_0562_),
    .X(_0580_));
 sg13g2_or4_2 _2812_ (.A(_1465_),
    .B(_0562_),
    .C(_0576_),
    .D(_0578_),
    .X(_0581_));
 sg13g2_and3_1 _2813_ (.X(_0582_),
    .A(\systolic_array.genblk1[4].accumulators_dlygate[8].A ),
    .B(net557),
    .C(_0581_));
 sg13g2_and3_1 _2814_ (.X(_0583_),
    .A(_1493_),
    .B(_0576_),
    .C(_0578_));
 sg13g2_a21oi_1 _2815_ (.A1(_1493_),
    .A2(_0576_),
    .Y(_0584_),
    .B1(_0578_));
 sg13g2_or3_1 _2816_ (.A(\systolic_array.genblk1[4].accumulators_dlygate[7].A ),
    .B(_0583_),
    .C(_0584_),
    .X(_0585_));
 sg13g2_o21ai_1 _2817_ (.B1(\systolic_array.genblk1[4].accumulators_dlygate[7].A ),
    .Y(_0586_),
    .A1(_0583_),
    .A2(_0584_));
 sg13g2_nand2_1 _2818_ (.Y(_0587_),
    .A(_1493_),
    .B(_0574_));
 sg13g2_xor2_1 _2819_ (.B(_0587_),
    .A(_0575_),
    .X(_0588_));
 sg13g2_nand2_1 _2820_ (.Y(_0589_),
    .A(_1495_),
    .B(_0588_));
 sg13g2_inv_1 _2821_ (.Y(_0590_),
    .A(_0589_));
 sg13g2_nand2_1 _2822_ (.Y(_0591_),
    .A(_0585_),
    .B(_0589_));
 sg13g2_or2_1 _2823_ (.X(_0592_),
    .B(_0588_),
    .A(_1495_));
 sg13g2_o21ai_1 _2824_ (.B1(_0586_),
    .Y(_0593_),
    .A1(_1495_),
    .A2(_0588_));
 sg13g2_a21oi_1 _2825_ (.A1(_0569_),
    .A2(_0571_),
    .Y(_0594_),
    .B1(\systolic_array.genblk2[0].mac[2].sign ));
 sg13g2_xnor2_1 _2826_ (.Y(_0595_),
    .A(_0572_),
    .B(_0594_));
 sg13g2_nor2_1 _2827_ (.A(\systolic_array.genblk1[4].accumulators_dlygate[5].A ),
    .B(_0595_),
    .Y(_0596_));
 sg13g2_nor2_1 _2828_ (.A(\systolic_array.genblk2[0].mac[2].sign ),
    .B(_0566_),
    .Y(_0597_));
 sg13g2_xor2_1 _2829_ (.B(_0597_),
    .A(_0568_),
    .X(_0598_));
 sg13g2_nand2_1 _2830_ (.Y(_0599_),
    .A(\systolic_array.genblk1[4].accumulators_dlygate[3].A ),
    .B(_0598_));
 sg13g2_a21oi_1 _2831_ (.A1(_1470_),
    .A2(_0563_),
    .Y(_0600_),
    .B1(\systolic_array.genblk2[0].mac[2].sign ));
 sg13g2_xnor2_1 _2832_ (.Y(_0601_),
    .A(_0565_),
    .B(_0600_));
 sg13g2_and2_1 _2833_ (.A(net854),
    .B(_0601_),
    .X(_0602_));
 sg13g2_nor2b_1 _2834_ (.A(net669),
    .B_N(\systolic_array.arg_top_curr[0] ),
    .Y(_0603_));
 sg13g2_a221oi_1 _2835_ (.B2(net689),
    .C1(\systolic_array.genblk2[0].mac[2].sign ),
    .B1(_0603_),
    .A1(_1470_),
    .Y(_0604_),
    .A2(_0563_));
 sg13g2_and2_1 _2836_ (.A(net670),
    .B(_0100_),
    .X(_0605_));
 sg13g2_nor2b_1 _2837_ (.A(net670),
    .B_N(_0101_),
    .Y(_0606_));
 sg13g2_nor3_1 _2838_ (.A(_1493_),
    .B(_0605_),
    .C(_0606_),
    .Y(_0607_));
 sg13g2_nor3_1 _2839_ (.A(_1497_),
    .B(_0604_),
    .C(_0607_),
    .Y(_0608_));
 sg13g2_nand2b_1 _2840_ (.Y(_0609_),
    .B(_0603_),
    .A_N(\systolic_array.genblk1[4].accumulators_dlygate[0].A ));
 sg13g2_o21ai_1 _2841_ (.B1(_1497_),
    .Y(_0610_),
    .A1(_0604_),
    .A2(_0607_));
 sg13g2_nand2b_1 _2842_ (.Y(_0611_),
    .B(_0610_),
    .A_N(_0608_));
 sg13g2_a21o_1 _2843_ (.A2(_0610_),
    .A1(_0609_),
    .B1(_0608_),
    .X(_0612_));
 sg13g2_xnor2_1 _2844_ (.Y(_0613_),
    .A(_1496_),
    .B(_0601_));
 sg13g2_a21oi_1 _2845_ (.A1(_0612_),
    .A2(_0613_),
    .Y(_0614_),
    .B1(_0602_));
 sg13g2_xnor2_1 _2846_ (.Y(_0615_),
    .A(net916),
    .B(_0598_));
 sg13g2_o21ai_1 _2847_ (.B1(_0599_),
    .Y(_0616_),
    .A1(_0614_),
    .A2(_0615_));
 sg13g2_nor2_1 _2848_ (.A(\systolic_array.genblk2[0].mac[2].sign ),
    .B(_0569_),
    .Y(_0617_));
 sg13g2_xor2_1 _2849_ (.B(_0617_),
    .A(_0571_),
    .X(_0618_));
 sg13g2_and2_1 _2850_ (.A(\systolic_array.genblk1[4].accumulators_dlygate[4].A ),
    .B(_0618_),
    .X(_0619_));
 sg13g2_nand2_1 _2851_ (.Y(_0620_),
    .A(\systolic_array.genblk1[4].accumulators_dlygate[4].A ),
    .B(_0618_));
 sg13g2_xor2_1 _2852_ (.B(_0618_),
    .A(\systolic_array.genblk1[4].accumulators_dlygate[4].A ),
    .X(_0621_));
 sg13g2_nand2_1 _2853_ (.Y(_0622_),
    .A(\systolic_array.genblk1[4].accumulators_dlygate[5].A ),
    .B(_0595_));
 sg13g2_nor2b_1 _2854_ (.A(_0596_),
    .B_N(_0622_),
    .Y(_0623_));
 sg13g2_nand3_1 _2855_ (.B(_0621_),
    .C(_0623_),
    .A(_0616_),
    .Y(_0624_));
 sg13g2_o21ai_1 _2856_ (.B1(_0622_),
    .Y(_0625_),
    .A1(_0596_),
    .A2(_0620_));
 sg13g2_nor2b_1 _2857_ (.A(_0625_),
    .B_N(_0624_),
    .Y(_0626_));
 sg13g2_a21oi_1 _2858_ (.A1(_0585_),
    .A2(_0593_),
    .Y(_0627_),
    .B1(_0625_));
 sg13g2_a22oi_1 _2859_ (.Y(_0628_),
    .B1(_0624_),
    .B2(_0627_),
    .A2(_0591_),
    .A1(_0586_));
 sg13g2_a21oi_1 _2860_ (.A1(net557),
    .A2(_0581_),
    .Y(_0629_),
    .B1(\systolic_array.genblk1[4].accumulators_dlygate[8].A ));
 sg13g2_or2_1 _2861_ (.X(_0630_),
    .B(_0629_),
    .A(_0582_));
 sg13g2_inv_1 _2862_ (.Y(_0631_),
    .A(_0630_));
 sg13g2_a21oi_1 _2863_ (.A1(_0628_),
    .A2(_0631_),
    .Y(_0632_),
    .B1(_0582_));
 sg13g2_xnor2_1 _2864_ (.Y(_0633_),
    .A(_1494_),
    .B(net557));
 sg13g2_a21oi_1 _2865_ (.A1(_0632_),
    .A2(_0633_),
    .Y(_0634_),
    .B1(net653));
 sg13g2_o21ai_1 _2866_ (.B1(_0634_),
    .Y(_0635_),
    .A1(_0632_),
    .A2(_0633_));
 sg13g2_o21ai_1 _2867_ (.B1(_0635_),
    .Y(_0636_),
    .A1(_1492_),
    .A2(net626));
 sg13g2_mux2_1 _2868_ (.A0(net806),
    .A1(_0636_),
    .S(net602),
    .X(_0055_));
 sg13g2_a21oi_1 _2869_ (.A1(_1494_),
    .A2(net557),
    .Y(_0637_),
    .B1(_0582_));
 sg13g2_nor2_1 _2870_ (.A(_0630_),
    .B(_0633_),
    .Y(_0638_));
 sg13g2_nand2_1 _2871_ (.Y(_0639_),
    .A(_0628_),
    .B(_0638_));
 sg13g2_nand2_1 _2872_ (.Y(_0640_),
    .A(\systolic_array.genblk1[4].accumulators_dlygate[10].A ),
    .B(net557));
 sg13g2_xnor2_1 _2873_ (.Y(_0641_),
    .A(\systolic_array.genblk1[4].accumulators_dlygate[10].A ),
    .B(net557));
 sg13g2_a21o_1 _2874_ (.A2(_0639_),
    .A1(_0637_),
    .B1(_0641_),
    .X(_0642_));
 sg13g2_nand3_1 _2875_ (.B(_0639_),
    .C(_0641_),
    .A(_0637_),
    .Y(_0643_));
 sg13g2_and2_1 _2876_ (.A(net626),
    .B(_0643_),
    .X(_0644_));
 sg13g2_a22oi_1 _2877_ (.Y(_0645_),
    .B1(_0642_),
    .B2(_0644_),
    .A2(net978),
    .A1(net654));
 sg13g2_nor2_1 _2878_ (.A(net828),
    .B(net598),
    .Y(_0646_));
 sg13g2_a21oi_1 _2879_ (.A1(net602),
    .A2(_0645_),
    .Y(_0048_),
    .B1(_0646_));
 sg13g2_nand2b_1 _2880_ (.Y(_0647_),
    .B(net556),
    .A_N(_0102_));
 sg13g2_xor2_1 _2881_ (.B(net557),
    .A(_0102_),
    .X(_0648_));
 sg13g2_a21oi_1 _2882_ (.A1(_0640_),
    .A2(_0642_),
    .Y(_0649_),
    .B1(_0648_));
 sg13g2_and3_1 _2883_ (.X(_0650_),
    .A(_0640_),
    .B(_0642_),
    .C(_0648_));
 sg13g2_nor3_1 _2884_ (.A(net653),
    .B(_0649_),
    .C(_0650_),
    .Y(_0651_));
 sg13g2_a21oi_1 _2885_ (.A1(net654),
    .A2(net928),
    .Y(_0652_),
    .B1(_0651_));
 sg13g2_nor2_1 _2886_ (.A(net767),
    .B(net602),
    .Y(_0653_));
 sg13g2_a21oi_1 _2887_ (.A1(net602),
    .A2(_0652_),
    .Y(_0049_),
    .B1(_0653_));
 sg13g2_nand3_1 _2888_ (.B(_0640_),
    .C(_0647_),
    .A(_0637_),
    .Y(_0654_));
 sg13g2_nor4_1 _2889_ (.A(_0630_),
    .B(_0633_),
    .C(_0641_),
    .D(_0648_),
    .Y(_0655_));
 sg13g2_and2_1 _2890_ (.A(_0628_),
    .B(_0655_),
    .X(_0656_));
 sg13g2_a21o_1 _2891_ (.A2(_0655_),
    .A1(_0628_),
    .B1(_0654_),
    .X(_0657_));
 sg13g2_and2_1 _2892_ (.A(\systolic_array.genblk1[4].accumulators_dlygate[12].A ),
    .B(net555),
    .X(_0658_));
 sg13g2_xor2_1 _2893_ (.B(net556),
    .A(\systolic_array.genblk1[4].accumulators_dlygate[12].A ),
    .X(_0659_));
 sg13g2_o21ai_1 _2894_ (.B1(net626),
    .Y(_0660_),
    .A1(_0657_),
    .A2(_0659_));
 sg13g2_a21oi_1 _2895_ (.A1(_0657_),
    .A2(_0659_),
    .Y(_0661_),
    .B1(_0660_));
 sg13g2_a21o_1 _2896_ (.A2(net993),
    .A1(net653),
    .B1(_0661_),
    .X(_0662_));
 sg13g2_mux2_1 _2897_ (.A0(net892),
    .A1(_0662_),
    .S(net598),
    .X(_0050_));
 sg13g2_nor2_1 _2898_ (.A(net930),
    .B(net598),
    .Y(_0663_));
 sg13g2_xnor2_1 _2899_ (.Y(_0664_),
    .A(_0103_),
    .B(net555));
 sg13g2_a21oi_1 _2900_ (.A1(_0657_),
    .A2(_0659_),
    .Y(_0665_),
    .B1(_0658_));
 sg13g2_nand2b_1 _2901_ (.Y(_0666_),
    .B(net653),
    .A_N(net969));
 sg13g2_xnor2_1 _2902_ (.Y(_0667_),
    .A(_0664_),
    .B(_0665_));
 sg13g2_o21ai_1 _2903_ (.B1(_0666_),
    .Y(_0668_),
    .A1(net653),
    .A2(_0667_));
 sg13g2_a21oi_2 _2904_ (.B1(_0663_),
    .Y(_0051_),
    .A2(_0668_),
    .A1(net601));
 sg13g2_xor2_1 _2905_ (.B(net555),
    .A(\systolic_array.genblk1[4].accumulators_dlygate[14].A ),
    .X(_0669_));
 sg13g2_o21ai_1 _2906_ (.B1(net555),
    .Y(_0670_),
    .A1(\systolic_array.genblk1[4].accumulators_dlygate[12].A ),
    .A2(_1499_));
 sg13g2_inv_1 _2907_ (.Y(_0671_),
    .A(_0670_));
 sg13g2_and2_1 _2908_ (.A(_0659_),
    .B(_0664_),
    .X(_0672_));
 sg13g2_a21o_1 _2909_ (.A2(_0672_),
    .A1(_0657_),
    .B1(_0671_),
    .X(_0673_));
 sg13g2_and2_1 _2910_ (.A(_0669_),
    .B(_0673_),
    .X(_0674_));
 sg13g2_nand2_1 _2911_ (.Y(_0675_),
    .A(net653),
    .B(net995));
 sg13g2_o21ai_1 _2912_ (.B1(net626),
    .Y(_0676_),
    .A1(_0669_),
    .A2(_0673_));
 sg13g2_o21ai_1 _2913_ (.B1(_0675_),
    .Y(_0677_),
    .A1(_0674_),
    .A2(_0676_));
 sg13g2_mux2_1 _2914_ (.A0(net541),
    .A1(_0677_),
    .S(net601),
    .X(_0052_));
 sg13g2_nand2_1 _2915_ (.Y(_0678_),
    .A(net653),
    .B(net989));
 sg13g2_xor2_1 _2916_ (.B(net556),
    .A(\systolic_array.genblk1[4].accumulators_dlygate[15].A ),
    .X(_0679_));
 sg13g2_a21oi_1 _2917_ (.A1(\systolic_array.genblk1[4].accumulators_dlygate[14].A ),
    .A2(net555),
    .Y(_0680_),
    .B1(_0674_));
 sg13g2_xor2_1 _2918_ (.B(_0680_),
    .A(_0679_),
    .X(_0681_));
 sg13g2_o21ai_1 _2919_ (.B1(_0678_),
    .Y(_0682_),
    .A1(net653),
    .A2(_0681_));
 sg13g2_mux2_1 _2920_ (.A0(net853),
    .A1(_0682_),
    .S(net601),
    .X(_0053_));
 sg13g2_nor2_1 _2921_ (.A(net876),
    .B(net601),
    .Y(_0683_));
 sg13g2_nand4_1 _2922_ (.B(_0669_),
    .C(_0672_),
    .A(_0656_),
    .Y(_0684_),
    .D(_0679_));
 sg13g2_o21ai_1 _2923_ (.B1(net555),
    .Y(_0685_),
    .A1(\systolic_array.genblk1[4].accumulators_dlygate[14].A ),
    .A2(\systolic_array.genblk1[4].accumulators_dlygate[15].A ));
 sg13g2_and2_1 _2924_ (.A(_0670_),
    .B(_0685_),
    .X(_0686_));
 sg13g2_nand3b_1 _2925_ (.B(_0684_),
    .C(_0686_),
    .Y(_0687_),
    .A_N(_0654_));
 sg13g2_o21ai_1 _2926_ (.B1(net626),
    .Y(_0688_),
    .A1(net555),
    .A2(_0687_));
 sg13g2_a21oi_1 _2927_ (.A1(net555),
    .A2(_0687_),
    .Y(_0689_),
    .B1(_0688_));
 sg13g2_xnor2_1 _2928_ (.Y(_0690_),
    .A(net918),
    .B(_0689_));
 sg13g2_a21oi_1 _2929_ (.A1(net601),
    .A2(_0690_),
    .Y(_0054_),
    .B1(_0683_));
 sg13g2_mux2_1 _2930_ (.A0(net509),
    .A1(net792),
    .S(net615),
    .X(_0063_));
 sg13g2_mux2_1 _2931_ (.A0(net418),
    .A1(net820),
    .S(net611),
    .X(_0056_));
 sg13g2_mux2_1 _2932_ (.A0(net493),
    .A1(net810),
    .S(net614),
    .X(_0057_));
 sg13g2_mux2_1 _2933_ (.A0(net448),
    .A1(net791),
    .S(net610),
    .X(_0058_));
 sg13g2_mux2_1 _2934_ (.A0(net496),
    .A1(net797),
    .S(net610),
    .X(_0059_));
 sg13g2_mux2_1 _2935_ (.A0(net454),
    .A1(net817),
    .S(net614),
    .X(_0060_));
 sg13g2_mux2_1 _2936_ (.A0(net499),
    .A1(net821),
    .S(net610),
    .X(_0061_));
 sg13g2_mux2_1 _2937_ (.A0(net474),
    .A1(net819),
    .S(net614),
    .X(_0062_));
 sg13g2_mux2_1 _2938_ (.A0(net682),
    .A1(net681),
    .S(net633),
    .X(_0691_));
 sg13g2_mux2_1 _2939_ (.A0(net685),
    .A1(_0691_),
    .S(_1500_),
    .X(_0692_));
 sg13g2_nor2b_1 _2940_ (.A(net688),
    .B_N(\systolic_array.genblk2[0].mac[3].div2 ),
    .Y(_0693_));
 sg13g2_nor2_1 _2941_ (.A(net691),
    .B(\systolic_array.genblk2[0].mac[3].div2 ),
    .Y(_0694_));
 sg13g2_nor3_2 _2942_ (.A(net668),
    .B(_0693_),
    .C(_0694_),
    .Y(_0695_));
 sg13g2_or3_1 _2943_ (.A(net668),
    .B(_0693_),
    .C(_0694_),
    .X(_0696_));
 sg13g2_nand2b_1 _2944_ (.Y(_0697_),
    .B(net668),
    .A_N(net691));
 sg13g2_mux2_1 _2945_ (.A0(net688),
    .A1(net685),
    .S(\systolic_array.genblk2[0].mac[3].div2 ),
    .X(_0698_));
 sg13g2_o21ai_1 _2946_ (.B1(_0697_),
    .Y(_0699_),
    .A1(net668),
    .A2(_0698_));
 sg13g2_mux2_1 _2947_ (.A0(net691),
    .A1(_0698_),
    .S(_1500_),
    .X(_0700_));
 sg13g2_mux2_1 _2948_ (.A0(net685),
    .A1(net682),
    .S(net633),
    .X(_0701_));
 sg13g2_mux2_1 _2949_ (.A0(net688),
    .A1(_0701_),
    .S(_1500_),
    .X(_0702_));
 sg13g2_nand3b_1 _2950_ (.B(_0696_),
    .C(_0699_),
    .Y(_0703_),
    .A_N(_0702_));
 sg13g2_nor4_2 _2951_ (.A(_0692_),
    .B(_0695_),
    .C(_0700_),
    .Y(_0704_),
    .D(_0702_));
 sg13g2_nand2_1 _2952_ (.Y(_0705_),
    .A(_1468_),
    .B(net633));
 sg13g2_a21oi_1 _2953_ (.A1(_1469_),
    .A2(_1501_),
    .Y(_0706_),
    .B1(net667));
 sg13g2_a22oi_1 _2954_ (.Y(_0707_),
    .B1(_0705_),
    .B2(_0706_),
    .A2(net667),
    .A1(net682));
 sg13g2_nand2b_1 _2955_ (.Y(_0708_),
    .B(net679),
    .A_N(net633));
 sg13g2_a21oi_1 _2956_ (.A1(\systolic_array.arg_top_curr[6] ),
    .A2(net633),
    .Y(_0709_),
    .B1(net667));
 sg13g2_a22oi_1 _2957_ (.Y(_0710_),
    .B1(_0708_),
    .B2(_0709_),
    .A2(net667),
    .A1(_1469_));
 sg13g2_inv_1 _2958_ (.Y(_0711_),
    .A(_0710_));
 sg13g2_nand3_1 _2959_ (.B(_0707_),
    .C(_0711_),
    .A(_0704_),
    .Y(_0712_));
 sg13g2_nand2_1 _2960_ (.Y(_0713_),
    .A(_1465_),
    .B(net633));
 sg13g2_a21oi_1 _2961_ (.A1(_1466_),
    .A2(_1501_),
    .Y(_0714_),
    .B1(net667));
 sg13g2_a22oi_1 _2962_ (.Y(_0715_),
    .B1(_0713_),
    .B2(_0714_),
    .A2(net667),
    .A1(net679));
 sg13g2_and4_1 _2963_ (.A(_0704_),
    .B(_0707_),
    .C(_0711_),
    .D(_0715_),
    .X(_0716_));
 sg13g2_nand2_1 _2964_ (.Y(_0717_),
    .A(_0116_),
    .B(net667));
 sg13g2_o21ai_1 _2965_ (.B1(_0717_),
    .Y(_0718_),
    .A1(_1467_),
    .A2(net667));
 sg13g2_nand2_1 _2966_ (.Y(_0719_),
    .A(_0716_),
    .B(_0718_));
 sg13g2_nor2_1 _2967_ (.A(net677),
    .B(\systolic_array.genblk2[0].mac[3].sign ),
    .Y(_0720_));
 sg13g2_a22oi_1 _2968_ (.Y(_0721_),
    .B1(_0719_),
    .B2(_0720_),
    .A2(\systolic_array.genblk2[0].mac[3].sign ),
    .A1(_1467_));
 sg13g2_inv_1 _2969_ (.Y(_0722_),
    .A(net548));
 sg13g2_xor2_1 _2970_ (.B(net549),
    .A(_0104_),
    .X(_0723_));
 sg13g2_nand4_1 _2971_ (.B(_1502_),
    .C(_0716_),
    .A(net677),
    .Y(_0724_),
    .D(_0718_));
 sg13g2_nand3_1 _2972_ (.B(net549),
    .C(_0724_),
    .A(\systolic_array.genblk1[6].accumulators_dlygate[8].A ),
    .Y(_0725_));
 sg13g2_a21oi_1 _2973_ (.A1(_0696_),
    .A2(_0699_),
    .Y(_0726_),
    .B1(\systolic_array.genblk2[0].mac[3].sign ));
 sg13g2_nand2_1 _2974_ (.Y(_0727_),
    .A(_0695_),
    .B(_0700_));
 sg13g2_mux2_1 _2975_ (.A0(_0101_),
    .A1(_0105_),
    .S(net633),
    .X(_0728_));
 sg13g2_nand2_1 _2976_ (.Y(_0729_),
    .A(_0100_),
    .B(net668));
 sg13g2_a21oi_1 _2977_ (.A1(_1500_),
    .A2(_0728_),
    .Y(_0730_),
    .B1(_1502_));
 sg13g2_a22oi_1 _2978_ (.Y(_0731_),
    .B1(_0729_),
    .B2(_0730_),
    .A2(_0727_),
    .A1(_0726_));
 sg13g2_and2_1 _2979_ (.A(\systolic_array.genblk1[6].accumulators_dlygate[1].A ),
    .B(_0731_),
    .X(_0732_));
 sg13g2_nand2b_1 _2980_ (.Y(_0733_),
    .B(_0695_),
    .A_N(\systolic_array.genblk1[6].accumulators_dlygate[0].A ));
 sg13g2_xor2_1 _2981_ (.B(_0731_),
    .A(net914),
    .X(_0734_));
 sg13g2_a21oi_1 _2982_ (.A1(_0733_),
    .A2(_0734_),
    .Y(_0735_),
    .B1(_0732_));
 sg13g2_a21o_1 _2983_ (.A2(_0734_),
    .A1(_0733_),
    .B1(_0732_),
    .X(_0736_));
 sg13g2_nand3_1 _2984_ (.B(_0692_),
    .C(_0703_),
    .A(_1502_),
    .Y(_0737_));
 sg13g2_a21o_1 _2985_ (.A2(_0703_),
    .A1(_1502_),
    .B1(_0692_),
    .X(_0738_));
 sg13g2_nand3_1 _2986_ (.B(_0737_),
    .C(_0738_),
    .A(_1505_),
    .Y(_0739_));
 sg13g2_a21oi_1 _2987_ (.A1(_0737_),
    .A2(_0738_),
    .Y(_0740_),
    .B1(_1505_));
 sg13g2_a21o_1 _2988_ (.A2(_0738_),
    .A1(_0737_),
    .B1(_1505_),
    .X(_0741_));
 sg13g2_nand2_1 _2989_ (.Y(_0742_),
    .A(_0739_),
    .B(_0741_));
 sg13g2_xnor2_1 _2990_ (.Y(_0743_),
    .A(_0702_),
    .B(_0726_));
 sg13g2_and2_1 _2991_ (.A(\systolic_array.genblk1[6].accumulators_dlygate[2].A ),
    .B(_0743_),
    .X(_0744_));
 sg13g2_xor2_1 _2992_ (.B(_0743_),
    .A(\systolic_array.genblk1[6].accumulators_dlygate[2].A ),
    .X(_0745_));
 sg13g2_nand3_1 _2993_ (.B(_0741_),
    .C(_0745_),
    .A(_0739_),
    .Y(_0746_));
 sg13g2_a21oi_1 _2994_ (.A1(_0739_),
    .A2(_0744_),
    .Y(_0747_),
    .B1(_0740_));
 sg13g2_o21ai_1 _2995_ (.B1(_0747_),
    .Y(_0748_),
    .A1(_0735_),
    .A2(_0746_));
 sg13g2_a21oi_1 _2996_ (.A1(_0704_),
    .A2(_0707_),
    .Y(_0749_),
    .B1(\systolic_array.genblk2[0].mac[3].sign ));
 sg13g2_xnor2_1 _2997_ (.Y(_0750_),
    .A(_0710_),
    .B(_0749_));
 sg13g2_nor2_1 _2998_ (.A(\systolic_array.genblk1[6].accumulators_dlygate[5].A ),
    .B(_0750_),
    .Y(_0751_));
 sg13g2_xor2_1 _2999_ (.B(_0750_),
    .A(\systolic_array.genblk1[6].accumulators_dlygate[5].A ),
    .X(_0752_));
 sg13g2_nor2_1 _3000_ (.A(\systolic_array.genblk2[0].mac[3].sign ),
    .B(_0704_),
    .Y(_0753_));
 sg13g2_xnor2_1 _3001_ (.Y(_0754_),
    .A(_0707_),
    .B(_0753_));
 sg13g2_nand2b_1 _3002_ (.Y(_0755_),
    .B(\systolic_array.genblk1[6].accumulators_dlygate[4].A ),
    .A_N(_0754_));
 sg13g2_xnor2_1 _3003_ (.Y(_0756_),
    .A(\systolic_array.genblk1[6].accumulators_dlygate[4].A ),
    .B(_0754_));
 sg13g2_and2_1 _3004_ (.A(_0752_),
    .B(_0756_),
    .X(_0757_));
 sg13g2_nor2_1 _3005_ (.A(_0751_),
    .B(_0755_),
    .Y(_0758_));
 sg13g2_a221oi_1 _3006_ (.B2(_0748_),
    .C1(_0758_),
    .B1(_0757_),
    .A1(\systolic_array.genblk1[6].accumulators_dlygate[5].A ),
    .Y(_0759_),
    .A2(_0750_));
 sg13g2_nor2_1 _3007_ (.A(\systolic_array.genblk2[0].mac[3].sign ),
    .B(_0716_),
    .Y(_0760_));
 sg13g2_xnor2_1 _3008_ (.Y(_0761_),
    .A(_0718_),
    .B(_0760_));
 sg13g2_nand2_1 _3009_ (.Y(_0762_),
    .A(_1503_),
    .B(_0761_));
 sg13g2_nand2_1 _3010_ (.Y(_0763_),
    .A(_1502_),
    .B(_0712_));
 sg13g2_xor2_1 _3011_ (.B(_0763_),
    .A(_0715_),
    .X(_0764_));
 sg13g2_nor2_1 _3012_ (.A(_1504_),
    .B(_0764_),
    .Y(_0765_));
 sg13g2_nor2_1 _3013_ (.A(_1503_),
    .B(_0761_),
    .Y(_0766_));
 sg13g2_a21oi_1 _3014_ (.A1(_0762_),
    .A2(_0765_),
    .Y(_0767_),
    .B1(_0766_));
 sg13g2_nand2_1 _3015_ (.Y(_0768_),
    .A(_1504_),
    .B(_0764_));
 sg13g2_a21oi_1 _3016_ (.A1(_0762_),
    .A2(_0768_),
    .Y(_0769_),
    .B1(_0766_));
 sg13g2_a21o_2 _3017_ (.A2(_0767_),
    .A1(_0759_),
    .B1(_0769_),
    .X(_0770_));
 sg13g2_a21o_1 _3018_ (.A2(_0724_),
    .A1(net549),
    .B1(\systolic_array.genblk1[6].accumulators_dlygate[8].A ),
    .X(_0771_));
 sg13g2_nand2_2 _3019_ (.Y(_0772_),
    .A(_0725_),
    .B(_0771_));
 sg13g2_o21ai_1 _3020_ (.B1(_0725_),
    .Y(_0773_),
    .A1(_0770_),
    .A2(_0772_));
 sg13g2_xnor2_1 _3021_ (.Y(_0774_),
    .A(_0723_),
    .B(_0773_));
 sg13g2_mux2_1 _3022_ (.A0(net958),
    .A1(_0774_),
    .S(net624),
    .X(_0775_));
 sg13g2_mux2_1 _3023_ (.A0(net904),
    .A1(_0775_),
    .S(net600),
    .X(_0071_));
 sg13g2_nor2_1 _3024_ (.A(net869),
    .B(net600),
    .Y(_0776_));
 sg13g2_o21ai_1 _3025_ (.B1(_0725_),
    .Y(_0777_),
    .A1(_0104_),
    .A2(_0722_));
 sg13g2_nor3_1 _3026_ (.A(_0723_),
    .B(_0770_),
    .C(_0772_),
    .Y(_0778_));
 sg13g2_nor2_1 _3027_ (.A(_0777_),
    .B(_0778_),
    .Y(_0779_));
 sg13g2_nand2_1 _3028_ (.Y(_0780_),
    .A(\systolic_array.genblk1[6].accumulators_dlygate[10].A ),
    .B(net548));
 sg13g2_xnor2_1 _3029_ (.Y(_0781_),
    .A(\systolic_array.genblk1[6].accumulators_dlygate[10].A ),
    .B(net548));
 sg13g2_or2_1 _3030_ (.X(_0782_),
    .B(_0781_),
    .A(_0779_));
 sg13g2_a21oi_1 _3031_ (.A1(_0779_),
    .A2(_0781_),
    .Y(_0783_),
    .B1(net651));
 sg13g2_a22oi_1 _3032_ (.Y(_0784_),
    .B1(_0782_),
    .B2(_0783_),
    .A2(net960),
    .A1(net651));
 sg13g2_a21oi_1 _3033_ (.A1(net596),
    .A2(_0784_),
    .Y(_0064_),
    .B1(_0776_));
 sg13g2_xnor2_1 _3034_ (.Y(_0785_),
    .A(_1507_),
    .B(net548));
 sg13g2_o21ai_1 _3035_ (.B1(_0780_),
    .Y(_0786_),
    .A1(_0779_),
    .A2(_0781_));
 sg13g2_nor2_1 _3036_ (.A(net624),
    .B(net973),
    .Y(_0787_));
 sg13g2_xor2_1 _3037_ (.B(_0786_),
    .A(_0785_),
    .X(_0788_));
 sg13g2_a21oi_1 _3038_ (.A1(net624),
    .A2(_0788_),
    .Y(_0789_),
    .B1(_0787_));
 sg13g2_mux2_1 _3039_ (.A0(net909),
    .A1(_0789_),
    .S(net597),
    .X(_0065_));
 sg13g2_or4_1 _3040_ (.A(_0723_),
    .B(_0772_),
    .C(_0781_),
    .D(_0785_),
    .X(_0790_));
 sg13g2_nor2_1 _3041_ (.A(_0770_),
    .B(_0790_),
    .Y(_0791_));
 sg13g2_o21ai_1 _3042_ (.B1(net548),
    .Y(_0792_),
    .A1(\systolic_array.genblk1[6].accumulators_dlygate[10].A ),
    .A2(_1507_));
 sg13g2_nor2b_1 _3043_ (.A(_0777_),
    .B_N(_0792_),
    .Y(_0793_));
 sg13g2_o21ai_1 _3044_ (.B1(_0793_),
    .Y(_0794_),
    .A1(_0770_),
    .A2(_0790_));
 sg13g2_xnor2_1 _3045_ (.Y(_0795_),
    .A(\systolic_array.genblk1[6].accumulators_dlygate[12].A ),
    .B(net547));
 sg13g2_nor2b_1 _3046_ (.A(_0795_),
    .B_N(_0794_),
    .Y(_0796_));
 sg13g2_xnor2_1 _3047_ (.Y(_0797_),
    .A(_0794_),
    .B(_0795_));
 sg13g2_nand2b_1 _3048_ (.Y(_0798_),
    .B(net651),
    .A_N(net999));
 sg13g2_o21ai_1 _3049_ (.B1(_0798_),
    .Y(_0799_),
    .A1(net651),
    .A2(_0797_));
 sg13g2_nor2_1 _3050_ (.A(net835),
    .B(net596),
    .Y(_0800_));
 sg13g2_a21oi_1 _3051_ (.A1(net599),
    .A2(_0799_),
    .Y(_0066_),
    .B1(_0800_));
 sg13g2_xnor2_1 _3052_ (.Y(_0801_),
    .A(_0107_),
    .B(net547));
 sg13g2_a21oi_1 _3053_ (.A1(\systolic_array.genblk1[6].accumulators_dlygate[12].A ),
    .A2(net547),
    .Y(_0802_),
    .B1(_0796_));
 sg13g2_xnor2_1 _3054_ (.Y(_0803_),
    .A(_0801_),
    .B(_0802_));
 sg13g2_mux2_1 _3055_ (.A0(net966),
    .A1(_0803_),
    .S(net624),
    .X(_0804_));
 sg13g2_mux2_1 _3056_ (.A0(net838),
    .A1(_0804_),
    .S(net599),
    .X(_0067_));
 sg13g2_o21ai_1 _3057_ (.B1(net547),
    .Y(_0805_),
    .A1(\systolic_array.genblk1[6].accumulators_dlygate[12].A ),
    .A2(_1508_));
 sg13g2_inv_1 _3058_ (.Y(_0806_),
    .A(_0805_));
 sg13g2_nor2b_1 _3059_ (.A(_0795_),
    .B_N(_0801_),
    .Y(_0807_));
 sg13g2_inv_1 _3060_ (.Y(_0808_),
    .A(_0807_));
 sg13g2_a21oi_1 _3061_ (.A1(_0794_),
    .A2(_0807_),
    .Y(_0809_),
    .B1(_0806_));
 sg13g2_nand2_1 _3062_ (.Y(_0810_),
    .A(\systolic_array.genblk1[6].accumulators_dlygate[14].A ),
    .B(net547));
 sg13g2_xnor2_1 _3063_ (.Y(_0811_),
    .A(\systolic_array.genblk1[6].accumulators_dlygate[14].A ),
    .B(net547));
 sg13g2_or2_1 _3064_ (.X(_0812_),
    .B(_0811_),
    .A(_0809_));
 sg13g2_a21oi_1 _3065_ (.A1(_0809_),
    .A2(_0811_),
    .Y(_0813_),
    .B1(net651));
 sg13g2_a22oi_1 _3066_ (.Y(_0814_),
    .B1(_0812_),
    .B2(_0813_),
    .A2(net985),
    .A1(net651));
 sg13g2_nor2_1 _3067_ (.A(net736),
    .B(net599),
    .Y(_0815_));
 sg13g2_a21oi_1 _3068_ (.A1(net598),
    .A2(_0814_),
    .Y(_0068_),
    .B1(_0815_));
 sg13g2_nand2b_1 _3069_ (.Y(_0816_),
    .B(net651),
    .A_N(net998));
 sg13g2_xnor2_1 _3070_ (.Y(_0817_),
    .A(\systolic_array.genblk1[6].accumulators_dlygate[15].A ),
    .B(net547));
 sg13g2_o21ai_1 _3071_ (.B1(_0810_),
    .Y(_0818_),
    .A1(_0809_),
    .A2(_0811_));
 sg13g2_xnor2_1 _3072_ (.Y(_0819_),
    .A(_0817_),
    .B(_0818_));
 sg13g2_o21ai_1 _3073_ (.B1(_0816_),
    .Y(_0820_),
    .A1(net651),
    .A2(_0819_));
 sg13g2_nor2_1 _3074_ (.A(net848),
    .B(net599),
    .Y(_0821_));
 sg13g2_a21oi_2 _3075_ (.B1(_0821_),
    .Y(_0069_),
    .A2(_0820_),
    .A1(net599));
 sg13g2_nor2_1 _3076_ (.A(net724),
    .B(net598),
    .Y(_0822_));
 sg13g2_nor3_1 _3077_ (.A(_0808_),
    .B(_0811_),
    .C(_0817_),
    .Y(_0823_));
 sg13g2_o21ai_1 _3078_ (.B1(net547),
    .Y(_0824_),
    .A1(\systolic_array.genblk1[6].accumulators_dlygate[14].A ),
    .A2(\systolic_array.genblk1[6].accumulators_dlygate[15].A ));
 sg13g2_nand3_1 _3079_ (.B(_0805_),
    .C(_0824_),
    .A(_0793_),
    .Y(_0825_));
 sg13g2_a21oi_1 _3080_ (.A1(_0791_),
    .A2(_0823_),
    .Y(_0826_),
    .B1(_0825_));
 sg13g2_o21ai_1 _3081_ (.B1(net624),
    .Y(_0827_),
    .A1(_0722_),
    .A2(_0826_));
 sg13g2_a21oi_2 _3082_ (.B1(_0827_),
    .Y(_0828_),
    .A2(_0826_),
    .A1(_0722_));
 sg13g2_xnor2_1 _3083_ (.Y(_0829_),
    .A(net921),
    .B(_0828_));
 sg13g2_a21oi_1 _3084_ (.A1(net598),
    .A2(_0829_),
    .Y(_0070_),
    .B1(_0822_));
 sg13g2_mux2_1 _3085_ (.A0(net446),
    .A1(net809),
    .S(net612),
    .X(_0079_));
 sg13g2_mux2_1 _3086_ (.A0(net451),
    .A1(net775),
    .S(net612),
    .X(_0072_));
 sg13g2_mux2_1 _3087_ (.A0(net453),
    .A1(net781),
    .S(net612),
    .X(_0073_));
 sg13g2_mux2_1 _3088_ (.A0(net486),
    .A1(net844),
    .S(net608),
    .X(_0074_));
 sg13g2_mux2_1 _3089_ (.A0(net466),
    .A1(net825),
    .S(net611),
    .X(_0075_));
 sg13g2_mux2_1 _3090_ (.A0(net443),
    .A1(net796),
    .S(net611),
    .X(_0076_));
 sg13g2_mux2_1 _3091_ (.A0(net435),
    .A1(net830),
    .S(net611),
    .X(_0077_));
 sg13g2_mux2_1 _3092_ (.A0(net491),
    .A1(net818),
    .S(net610),
    .X(_0078_));
 sg13g2_mux2_1 _3093_ (.A0(net682),
    .A1(net681),
    .S(net632),
    .X(_0830_));
 sg13g2_mux2_2 _3094_ (.A0(net685),
    .A1(_0830_),
    .S(_1509_),
    .X(_0831_));
 sg13g2_nor2b_1 _3095_ (.A(net688),
    .B_N(net631),
    .Y(_0832_));
 sg13g2_nor2_1 _3096_ (.A(net691),
    .B(net631),
    .Y(_0833_));
 sg13g2_nor3_2 _3097_ (.A(net666),
    .B(_0832_),
    .C(_0833_),
    .Y(_0834_));
 sg13g2_or3_1 _3098_ (.A(net666),
    .B(_0832_),
    .C(_0833_),
    .X(_0835_));
 sg13g2_nand2b_1 _3099_ (.Y(_0836_),
    .B(net666),
    .A_N(net691));
 sg13g2_mux2_1 _3100_ (.A0(net688),
    .A1(net685),
    .S(net631),
    .X(_0837_));
 sg13g2_o21ai_1 _3101_ (.B1(_0836_),
    .Y(_0838_),
    .A1(net666),
    .A2(_0837_));
 sg13g2_mux2_1 _3102_ (.A0(net691),
    .A1(_0837_),
    .S(_1509_),
    .X(_0839_));
 sg13g2_mux2_1 _3103_ (.A0(net685),
    .A1(net682),
    .S(net631),
    .X(_0840_));
 sg13g2_mux2_2 _3104_ (.A0(net688),
    .A1(_0840_),
    .S(_1509_),
    .X(_0841_));
 sg13g2_nand3b_1 _3105_ (.B(_0835_),
    .C(_0838_),
    .Y(_0842_),
    .A_N(_0841_));
 sg13g2_nor4_2 _3106_ (.A(_0831_),
    .B(_0834_),
    .C(_0839_),
    .Y(_0843_),
    .D(_0841_));
 sg13g2_or4_1 _3107_ (.A(_0831_),
    .B(_0834_),
    .C(_0839_),
    .D(_0841_),
    .X(_0844_));
 sg13g2_nand2b_1 _3108_ (.Y(_0845_),
    .B(net665),
    .A_N(net682));
 sg13g2_nand2_1 _3109_ (.Y(_0846_),
    .A(net679),
    .B(net631));
 sg13g2_o21ai_1 _3110_ (.B1(_0846_),
    .Y(_0847_),
    .A1(_1469_),
    .A2(net632));
 sg13g2_o21ai_1 _3111_ (.B1(_0845_),
    .Y(_0848_),
    .A1(net665),
    .A2(_0847_));
 sg13g2_mux2_2 _3112_ (.A0(net682),
    .A1(_0847_),
    .S(_1509_),
    .X(_0849_));
 sg13g2_nand2b_1 _3113_ (.Y(_0850_),
    .B(net679),
    .A_N(net631));
 sg13g2_a21oi_1 _3114_ (.A1(\systolic_array.arg_top_curr[6] ),
    .A2(net631),
    .Y(_0851_),
    .B1(net666));
 sg13g2_a22oi_1 _3115_ (.Y(_0852_),
    .B1(_0850_),
    .B2(_0851_),
    .A2(net665),
    .A1(_1469_));
 sg13g2_nor3_1 _3116_ (.A(_0844_),
    .B(_0849_),
    .C(_0852_),
    .Y(_0853_));
 sg13g2_mux2_1 _3117_ (.A0(\systolic_array.arg_top_curr[6] ),
    .A1(net677),
    .S(net631),
    .X(_0854_));
 sg13g2_nor2_1 _3118_ (.A(net665),
    .B(_0854_),
    .Y(_0855_));
 sg13g2_a21oi_2 _3119_ (.B1(_0855_),
    .Y(_0856_),
    .A2(net665),
    .A1(_1468_));
 sg13g2_nor4_1 _3120_ (.A(_0844_),
    .B(_0849_),
    .C(_0852_),
    .D(_0856_),
    .Y(_0857_));
 sg13g2_or4_1 _3121_ (.A(_0844_),
    .B(_0849_),
    .C(_0852_),
    .D(_0856_),
    .X(_0858_));
 sg13g2_nand2_1 _3122_ (.Y(_0859_),
    .A(_0116_),
    .B(net665));
 sg13g2_o21ai_1 _3123_ (.B1(_0859_),
    .Y(_0860_),
    .A1(_1467_),
    .A2(net665));
 sg13g2_inv_1 _3124_ (.Y(_0861_),
    .A(_0860_));
 sg13g2_nor2_1 _3125_ (.A(net677),
    .B(\systolic_array.genblk2[0].mac[4].sign ),
    .Y(_0862_));
 sg13g2_o21ai_1 _3126_ (.B1(_0862_),
    .Y(_0863_),
    .A1(_0858_),
    .A2(_0861_));
 sg13g2_nand2_2 _3127_ (.Y(_0864_),
    .A(_1467_),
    .B(\systolic_array.genblk2[0].mac[4].sign ));
 sg13g2_and2_1 _3128_ (.A(_0863_),
    .B(_0864_),
    .X(_0865_));
 sg13g2_nand2_2 _3129_ (.Y(_0866_),
    .A(_0863_),
    .B(_0864_));
 sg13g2_xnor2_1 _3130_ (.Y(_0867_),
    .A(_0108_),
    .B(_0866_));
 sg13g2_nand4_1 _3131_ (.B(_1510_),
    .C(_0857_),
    .A(net677),
    .Y(_0868_),
    .D(_0860_));
 sg13g2_nand3_1 _3132_ (.B(_0864_),
    .C(_0868_),
    .A(_0863_),
    .Y(_0869_));
 sg13g2_nand3_1 _3133_ (.B(net546),
    .C(_0868_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[8].A ),
    .Y(_0870_));
 sg13g2_nand3_1 _3134_ (.B(_0858_),
    .C(_0860_),
    .A(_1510_),
    .Y(_0871_));
 sg13g2_o21ai_1 _3135_ (.B1(_0861_),
    .Y(_0872_),
    .A1(\systolic_array.genblk2[0].mac[4].sign ),
    .A2(_0857_));
 sg13g2_nand2_1 _3136_ (.Y(_0873_),
    .A(_0871_),
    .B(_0872_));
 sg13g2_nand2b_1 _3137_ (.Y(_0874_),
    .B(_0873_),
    .A_N(\systolic_array.genblk1[8].accumulators_dlygate[7].A ));
 sg13g2_and3_1 _3138_ (.X(_0875_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[7].A ),
    .B(_0871_),
    .C(_0872_));
 sg13g2_nor2_1 _3139_ (.A(\systolic_array.genblk2[0].mac[4].sign ),
    .B(_0853_),
    .Y(_0876_));
 sg13g2_xor2_1 _3140_ (.B(_0876_),
    .A(_0856_),
    .X(_0877_));
 sg13g2_nand2_1 _3141_ (.Y(_0878_),
    .A(_1511_),
    .B(_0877_));
 sg13g2_a21oi_1 _3142_ (.A1(_0874_),
    .A2(_0878_),
    .Y(_0879_),
    .B1(_0875_));
 sg13g2_a21oi_1 _3143_ (.A1(_0835_),
    .A2(_0838_),
    .Y(_0880_),
    .B1(\systolic_array.genblk2[0].mac[4].sign ));
 sg13g2_nand2_1 _3144_ (.Y(_0881_),
    .A(_0834_),
    .B(_0839_));
 sg13g2_mux2_1 _3145_ (.A0(_0101_),
    .A1(_0105_),
    .S(net632),
    .X(_0882_));
 sg13g2_nand2_1 _3146_ (.Y(_0883_),
    .A(_0100_),
    .B(net666));
 sg13g2_a21oi_1 _3147_ (.A1(_1509_),
    .A2(_0882_),
    .Y(_0884_),
    .B1(_1510_));
 sg13g2_a22oi_1 _3148_ (.Y(_0885_),
    .B1(_0883_),
    .B2(_0884_),
    .A2(_0881_),
    .A1(_0880_));
 sg13g2_and2_1 _3149_ (.A(\systolic_array.genblk1[8].accumulators_dlygate[1].A ),
    .B(_0885_),
    .X(_0886_));
 sg13g2_nand2b_2 _3150_ (.Y(_0887_),
    .B(_0834_),
    .A_N(net851));
 sg13g2_xor2_1 _3151_ (.B(_0885_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[1].A ),
    .X(_0888_));
 sg13g2_a21oi_1 _3152_ (.A1(_0887_),
    .A2(_0888_),
    .Y(_0889_),
    .B1(_0886_));
 sg13g2_a21o_1 _3153_ (.A2(_0888_),
    .A1(_0887_),
    .B1(_0886_),
    .X(_0890_));
 sg13g2_nand3_1 _3154_ (.B(_0831_),
    .C(_0842_),
    .A(_1510_),
    .Y(_0891_));
 sg13g2_a21o_1 _3155_ (.A2(_0842_),
    .A1(_1510_),
    .B1(_0831_),
    .X(_0892_));
 sg13g2_nand3_1 _3156_ (.B(_0891_),
    .C(_0892_),
    .A(_1513_),
    .Y(_0893_));
 sg13g2_a21oi_1 _3157_ (.A1(_0891_),
    .A2(_0892_),
    .Y(_0894_),
    .B1(_1513_));
 sg13g2_a21o_1 _3158_ (.A2(_0892_),
    .A1(_0891_),
    .B1(_1513_),
    .X(_0895_));
 sg13g2_nand2_1 _3159_ (.Y(_0896_),
    .A(_0893_),
    .B(_0895_));
 sg13g2_xnor2_1 _3160_ (.Y(_0897_),
    .A(_0841_),
    .B(_0880_));
 sg13g2_and2_1 _3161_ (.A(\systolic_array.genblk1[8].accumulators_dlygate[2].A ),
    .B(_0897_),
    .X(_0898_));
 sg13g2_xor2_1 _3162_ (.B(_0897_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[2].A ),
    .X(_0899_));
 sg13g2_nand3_1 _3163_ (.B(_0895_),
    .C(_0899_),
    .A(_0893_),
    .Y(_0900_));
 sg13g2_a21oi_1 _3164_ (.A1(_0893_),
    .A2(_0898_),
    .Y(_0901_),
    .B1(_0894_));
 sg13g2_o21ai_1 _3165_ (.B1(_0901_),
    .Y(_0902_),
    .A1(_0889_),
    .A2(_0900_));
 sg13g2_a21oi_1 _3166_ (.A1(_0843_),
    .A2(_0848_),
    .Y(_0903_),
    .B1(\systolic_array.genblk2[0].mac[4].sign ));
 sg13g2_xnor2_1 _3167_ (.Y(_0904_),
    .A(_0852_),
    .B(_0903_));
 sg13g2_nand2_1 _3168_ (.Y(_0905_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[5].A ),
    .B(_0904_));
 sg13g2_xor2_1 _3169_ (.B(_0904_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[5].A ),
    .X(_0906_));
 sg13g2_nor3_2 _3170_ (.A(\systolic_array.genblk2[0].mac[4].sign ),
    .B(_0843_),
    .C(_0849_),
    .Y(_0907_));
 sg13g2_a21oi_1 _3171_ (.A1(_1510_),
    .A2(_0844_),
    .Y(_0908_),
    .B1(_0848_));
 sg13g2_nor3_1 _3172_ (.A(_1512_),
    .B(_0907_),
    .C(_0908_),
    .Y(_0909_));
 sg13g2_o21ai_1 _3173_ (.B1(_1512_),
    .Y(_0910_),
    .A1(_0907_),
    .A2(_0908_));
 sg13g2_nor2b_1 _3174_ (.A(_0909_),
    .B_N(_0910_),
    .Y(_0911_));
 sg13g2_and2_1 _3175_ (.A(_0906_),
    .B(_0911_),
    .X(_0912_));
 sg13g2_nand2_1 _3176_ (.Y(_0913_),
    .A(_0902_),
    .B(_0912_));
 sg13g2_o21ai_1 _3177_ (.B1(_0909_),
    .Y(_0914_),
    .A1(\systolic_array.genblk1[8].accumulators_dlygate[5].A ),
    .A2(_0904_));
 sg13g2_nand3_1 _3178_ (.B(_0913_),
    .C(_0914_),
    .A(_0905_),
    .Y(_0915_));
 sg13g2_nor2_1 _3179_ (.A(_1511_),
    .B(_0877_),
    .Y(_0916_));
 sg13g2_nand3b_1 _3180_ (.B(_0905_),
    .C(_0914_),
    .Y(_0917_),
    .A_N(_0875_));
 sg13g2_a221oi_1 _3181_ (.B2(_0874_),
    .C1(_0917_),
    .B1(_0916_),
    .A1(_0902_),
    .Y(_0918_),
    .A2(_0912_));
 sg13g2_or2_1 _3182_ (.X(_0919_),
    .B(_0918_),
    .A(_0879_));
 sg13g2_xor2_1 _3183_ (.B(_0869_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[8].A ),
    .X(_0920_));
 sg13g2_o21ai_1 _3184_ (.B1(_0870_),
    .Y(_0921_),
    .A1(_0919_),
    .A2(_0920_));
 sg13g2_xnor2_1 _3185_ (.Y(_0922_),
    .A(_0867_),
    .B(_0921_));
 sg13g2_mux2_1 _3186_ (.A0(net983),
    .A1(_0922_),
    .S(net621),
    .X(_0923_));
 sg13g2_mux2_1 _3187_ (.A0(net748),
    .A1(_0923_),
    .S(net600),
    .X(_0087_));
 sg13g2_o21ai_1 _3188_ (.B1(_0870_),
    .Y(_0924_),
    .A1(_0108_),
    .A2(_0866_));
 sg13g2_or2_1 _3189_ (.X(_0925_),
    .B(_0920_),
    .A(_0867_));
 sg13g2_nor3_1 _3190_ (.A(_0879_),
    .B(_0918_),
    .C(_0925_),
    .Y(_0926_));
 sg13g2_nor2_1 _3191_ (.A(_0924_),
    .B(_0926_),
    .Y(_0927_));
 sg13g2_nand2_1 _3192_ (.Y(_0928_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[10].A ),
    .B(net546));
 sg13g2_xnor2_1 _3193_ (.Y(_0929_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[10].A ),
    .B(net546));
 sg13g2_xnor2_1 _3194_ (.Y(_0930_),
    .A(_0927_),
    .B(_0929_));
 sg13g2_nand2_1 _3195_ (.Y(_0931_),
    .A(net621),
    .B(_0930_));
 sg13g2_o21ai_1 _3196_ (.B1(_0931_),
    .Y(_0932_),
    .A1(net621),
    .A2(net988));
 sg13g2_nor2_1 _3197_ (.A(net539),
    .B(net600),
    .Y(_0933_));
 sg13g2_a21oi_1 _3198_ (.A1(net600),
    .A2(_0932_),
    .Y(_0080_),
    .B1(_0933_));
 sg13g2_xnor2_1 _3199_ (.Y(_0934_),
    .A(_0109_),
    .B(net546));
 sg13g2_o21ai_1 _3200_ (.B1(_0928_),
    .Y(_0935_),
    .A1(_0927_),
    .A2(_0929_));
 sg13g2_o21ai_1 _3201_ (.B1(net621),
    .Y(_0936_),
    .A1(_0934_),
    .A2(_0935_));
 sg13g2_a21oi_1 _3202_ (.A1(_0934_),
    .A2(_0935_),
    .Y(_0937_),
    .B1(_0936_));
 sg13g2_a21o_1 _3203_ (.A2(net982),
    .A1(net650),
    .B1(_0937_),
    .X(_0938_));
 sg13g2_mux2_1 _3204_ (.A0(net726),
    .A1(_0938_),
    .S(net596),
    .X(_0081_));
 sg13g2_nand2b_1 _3205_ (.Y(_0939_),
    .B(_0934_),
    .A_N(_0929_));
 sg13g2_nor4_1 _3206_ (.A(_0879_),
    .B(_0918_),
    .C(_0925_),
    .D(_0939_),
    .Y(_0940_));
 sg13g2_a21oi_1 _3207_ (.A1(_1515_),
    .A2(_0109_),
    .Y(_0941_),
    .B1(_0866_));
 sg13g2_nor2_1 _3208_ (.A(_0924_),
    .B(_0941_),
    .Y(_0942_));
 sg13g2_nand2b_1 _3209_ (.Y(_0943_),
    .B(_0942_),
    .A_N(_0940_));
 sg13g2_xnor2_1 _3210_ (.Y(_0944_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[12].A ),
    .B(net545));
 sg13g2_nor2b_1 _3211_ (.A(_0944_),
    .B_N(_0943_),
    .Y(_0945_));
 sg13g2_xnor2_1 _3212_ (.Y(_0946_),
    .A(_0943_),
    .B(_0944_));
 sg13g2_nand2b_1 _3213_ (.Y(_0947_),
    .B(net650),
    .A_N(net997));
 sg13g2_o21ai_1 _3214_ (.B1(_0947_),
    .Y(_0948_),
    .A1(net650),
    .A2(_0946_));
 sg13g2_nor2_1 _3215_ (.A(net754),
    .B(net596),
    .Y(_0949_));
 sg13g2_a21oi_1 _3216_ (.A1(net596),
    .A2(_0948_),
    .Y(_0082_),
    .B1(_0949_));
 sg13g2_xnor2_1 _3217_ (.Y(_0950_),
    .A(_0110_),
    .B(net545));
 sg13g2_a21oi_1 _3218_ (.A1(\systolic_array.genblk1[8].accumulators_dlygate[12].A ),
    .A2(net545),
    .Y(_0951_),
    .B1(_0945_));
 sg13g2_xnor2_1 _3219_ (.Y(_0952_),
    .A(_0950_),
    .B(_0951_));
 sg13g2_mux2_1 _3220_ (.A0(net968),
    .A1(_0952_),
    .S(net621),
    .X(_0953_));
 sg13g2_mux2_1 _3221_ (.A0(net769),
    .A1(_0953_),
    .S(net596),
    .X(_0083_));
 sg13g2_nor2_1 _3222_ (.A(net856),
    .B(net596),
    .Y(_0954_));
 sg13g2_o21ai_1 _3223_ (.B1(net545),
    .Y(_0955_),
    .A1(\systolic_array.genblk1[8].accumulators_dlygate[12].A ),
    .A2(_1516_));
 sg13g2_inv_1 _3224_ (.Y(_0956_),
    .A(_0955_));
 sg13g2_nor2b_1 _3225_ (.A(_0944_),
    .B_N(_0950_),
    .Y(_0957_));
 sg13g2_a21oi_1 _3226_ (.A1(_0943_),
    .A2(_0957_),
    .Y(_0958_),
    .B1(_0956_));
 sg13g2_nand2_1 _3227_ (.Y(_0959_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[14].A ),
    .B(net545));
 sg13g2_xnor2_1 _3228_ (.Y(_0960_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[14].A ),
    .B(net545));
 sg13g2_or2_1 _3229_ (.X(_0961_),
    .B(_0960_),
    .A(_0958_));
 sg13g2_a21oi_1 _3230_ (.A1(_0958_),
    .A2(_0960_),
    .Y(_0962_),
    .B1(net650));
 sg13g2_a22oi_1 _3231_ (.Y(_0963_),
    .B1(_0961_),
    .B2(_0962_),
    .A2(net975),
    .A1(net650));
 sg13g2_a21oi_1 _3232_ (.A1(net596),
    .A2(_0963_),
    .Y(_0084_),
    .B1(_0954_));
 sg13g2_nand2b_1 _3233_ (.Y(_0964_),
    .B(net650),
    .A_N(net996));
 sg13g2_xnor2_1 _3234_ (.Y(_0965_),
    .A(\systolic_array.genblk1[8].accumulators_dlygate[15].A ),
    .B(net545));
 sg13g2_o21ai_1 _3235_ (.B1(_0959_),
    .Y(_0966_),
    .A1(_0958_),
    .A2(_0960_));
 sg13g2_xnor2_1 _3236_ (.Y(_0967_),
    .A(_0965_),
    .B(_0966_));
 sg13g2_o21ai_1 _3237_ (.B1(_0964_),
    .Y(_0968_),
    .A1(net650),
    .A2(_0967_));
 sg13g2_nor2_1 _3238_ (.A(net728),
    .B(net597),
    .Y(_0969_));
 sg13g2_a21oi_1 _3239_ (.A1(net597),
    .A2(_0968_),
    .Y(_0085_),
    .B1(_0969_));
 sg13g2_nor2_1 _3240_ (.A(net787),
    .B(net598),
    .Y(_0970_));
 sg13g2_nor2_1 _3241_ (.A(_0960_),
    .B(_0965_),
    .Y(_0971_));
 sg13g2_nand3_1 _3242_ (.B(_0957_),
    .C(_0971_),
    .A(_0940_),
    .Y(_0972_));
 sg13g2_o21ai_1 _3243_ (.B1(net545),
    .Y(_0973_),
    .A1(\systolic_array.genblk1[8].accumulators_dlygate[14].A ),
    .A2(\systolic_array.genblk1[8].accumulators_dlygate[15].A ));
 sg13g2_and4_1 _3244_ (.A(_0942_),
    .B(_0955_),
    .C(_0972_),
    .D(_0973_),
    .X(_0974_));
 sg13g2_o21ai_1 _3245_ (.B1(net621),
    .Y(_0975_),
    .A1(_0866_),
    .A2(_0974_));
 sg13g2_a21oi_2 _3246_ (.B1(_0975_),
    .Y(_0976_),
    .A2(_0974_),
    .A1(_0866_));
 sg13g2_xnor2_1 _3247_ (.Y(_0977_),
    .A(net944),
    .B(_0976_));
 sg13g2_a21oi_1 _3248_ (.A1(net598),
    .A2(_0977_),
    .Y(_0086_),
    .B1(_0970_));
 sg13g2_mux2_1 _3249_ (.A0(net410),
    .A1(net740),
    .S(net612),
    .X(_0095_));
 sg13g2_mux2_1 _3250_ (.A0(net487),
    .A1(net814),
    .S(net608),
    .X(_0088_));
 sg13g2_mux2_1 _3251_ (.A0(net503),
    .A1(net779),
    .S(net608),
    .X(_0089_));
 sg13g2_mux2_1 _3252_ (.A0(net470),
    .A1(net824),
    .S(net608),
    .X(_0090_));
 sg13g2_mux2_1 _3253_ (.A0(net507),
    .A1(net831),
    .S(net608),
    .X(_0091_));
 sg13g2_mux2_1 _3254_ (.A0(net502),
    .A1(net816),
    .S(net607),
    .X(_0092_));
 sg13g2_mux2_1 _3255_ (.A0(net489),
    .A1(net826),
    .S(net609),
    .X(_0093_));
 sg13g2_mux2_1 _3256_ (.A0(net424),
    .A1(net771),
    .S(net610),
    .X(_0094_));
 sg13g2_nand2_1 _3257_ (.Y(_0978_),
    .A(net742),
    .B(net608));
 sg13g2_nand2_1 _3258_ (.Y(_0979_),
    .A(_0115_),
    .B(net661));
 sg13g2_nand2b_1 _3259_ (.Y(_0980_),
    .B(net690),
    .A_N(net664));
 sg13g2_nor2b_1 _3260_ (.A(net664),
    .B_N(net687),
    .Y(_0981_));
 sg13g2_a21o_1 _3261_ (.A2(net664),
    .A1(net690),
    .B1(_0981_),
    .X(_0982_));
 sg13g2_nor3_1 _3262_ (.A(net690),
    .B(net692),
    .C(_0981_),
    .Y(_0983_));
 sg13g2_nor2b_1 _3263_ (.A(net663),
    .B_N(net684),
    .Y(_0984_));
 sg13g2_a21oi_1 _3264_ (.A1(net685),
    .A2(net663),
    .Y(_0985_),
    .B1(_0984_));
 sg13g2_nor4_2 _3265_ (.A(net685),
    .B(net688),
    .C(net691),
    .Y(_0986_),
    .D(_0984_));
 sg13g2_nor2_1 _3266_ (.A(net681),
    .B(net663),
    .Y(_0987_));
 sg13g2_nand2b_1 _3267_ (.Y(_0988_),
    .B(net663),
    .A_N(net682));
 sg13g2_nor2b_1 _3268_ (.A(_0987_),
    .B_N(_0988_),
    .Y(_0989_));
 sg13g2_nand2b_1 _3269_ (.Y(_0990_),
    .B(_0988_),
    .A_N(_0987_));
 sg13g2_and2_1 _3270_ (.A(_0986_),
    .B(_0990_),
    .X(_0991_));
 sg13g2_mux2_1 _3271_ (.A0(net679),
    .A1(net681),
    .S(net663),
    .X(_0992_));
 sg13g2_inv_1 _3272_ (.Y(_0993_),
    .A(_0992_));
 sg13g2_mux2_1 _3273_ (.A0(_0116_),
    .A1(_0099_),
    .S(net663),
    .X(_0994_));
 sg13g2_and4_1 _3274_ (.A(_0986_),
    .B(_0990_),
    .C(_0993_),
    .D(_0994_),
    .X(_0995_));
 sg13g2_nand2_1 _3275_ (.Y(_0996_),
    .A(\systolic_array.arg_top_curr[6] ),
    .B(net663));
 sg13g2_o21ai_1 _3276_ (.B1(_0996_),
    .Y(_0997_),
    .A1(_1465_),
    .A2(net663));
 sg13g2_inv_1 _3277_ (.Y(_0998_),
    .A(_0997_));
 sg13g2_a21oi_1 _3278_ (.A1(_0995_),
    .A2(_0998_),
    .Y(_0999_),
    .B1(net677));
 sg13g2_o21ai_1 _3279_ (.B1(_0979_),
    .Y(_1000_),
    .A1(net661),
    .A2(_0999_));
 sg13g2_and4_1 _3280_ (.A(net677),
    .B(_0979_),
    .C(_0995_),
    .D(_0998_),
    .X(_1001_));
 sg13g2_inv_1 _3281_ (.Y(_1002_),
    .A(_1001_));
 sg13g2_and3_1 _3282_ (.X(_1003_),
    .A(\systolic_array.genblk1[10].accumulators_dlygate[8].A ),
    .B(net554),
    .C(_1002_));
 sg13g2_a21oi_1 _3283_ (.A1(_0986_),
    .A2(_0990_),
    .Y(_1004_),
    .B1(net661));
 sg13g2_xnor2_1 _3284_ (.Y(_1005_),
    .A(_0992_),
    .B(_1004_));
 sg13g2_nor2_1 _3285_ (.A(\systolic_array.genblk1[10].accumulators_dlygate[5].A ),
    .B(_1005_),
    .Y(_1006_));
 sg13g2_nand2_1 _3286_ (.Y(_1007_),
    .A(\systolic_array.genblk1[10].accumulators_dlygate[5].A ),
    .B(_1005_));
 sg13g2_nand2b_1 _3287_ (.Y(_1008_),
    .B(_1007_),
    .A_N(_1006_));
 sg13g2_nor2_1 _3288_ (.A(\systolic_array.genblk2[0].mac[5].sign ),
    .B(_0983_),
    .Y(_1009_));
 sg13g2_xor2_1 _3289_ (.B(_1009_),
    .A(_0985_),
    .X(_1010_));
 sg13g2_and2_1 _3290_ (.A(\systolic_array.genblk1[10].accumulators_dlygate[3].A ),
    .B(_1010_),
    .X(_1011_));
 sg13g2_a21oi_1 _3291_ (.A1(_1470_),
    .A2(_0980_),
    .Y(_1012_),
    .B1(\systolic_array.genblk2[0].mac[5].sign ));
 sg13g2_xnor2_1 _3292_ (.Y(_1013_),
    .A(_0982_),
    .B(_1012_));
 sg13g2_nand2_1 _3293_ (.Y(_1014_),
    .A(\systolic_array.genblk1[10].accumulators_dlygate[2].A ),
    .B(_1013_));
 sg13g2_nor2b_1 _3294_ (.A(net664),
    .B_N(net691),
    .Y(_1015_));
 sg13g2_a221oi_1 _3295_ (.B2(net688),
    .C1(net661),
    .B1(_1015_),
    .A1(_1470_),
    .Y(_1016_),
    .A2(_0980_));
 sg13g2_and2_1 _3296_ (.A(_0100_),
    .B(net664),
    .X(_1017_));
 sg13g2_nor2b_1 _3297_ (.A(net664),
    .B_N(_0101_),
    .Y(_1018_));
 sg13g2_nor3_1 _3298_ (.A(_1517_),
    .B(_1017_),
    .C(_1018_),
    .Y(_1019_));
 sg13g2_nor3_1 _3299_ (.A(_1520_),
    .B(_1016_),
    .C(_1019_),
    .Y(_1020_));
 sg13g2_nand2b_1 _3300_ (.Y(_1021_),
    .B(_1015_),
    .A_N(\systolic_array.genblk1[10].accumulators_dlygate[0].A ));
 sg13g2_o21ai_1 _3301_ (.B1(_1520_),
    .Y(_1022_),
    .A1(_1016_),
    .A2(_1019_));
 sg13g2_nand2b_1 _3302_ (.Y(_1023_),
    .B(_1022_),
    .A_N(_1020_));
 sg13g2_a21oi_1 _3303_ (.A1(_1021_),
    .A2(_1022_),
    .Y(_1024_),
    .B1(_1020_));
 sg13g2_xnor2_1 _3304_ (.Y(_1025_),
    .A(\systolic_array.genblk1[10].accumulators_dlygate[2].A ),
    .B(_1013_));
 sg13g2_o21ai_1 _3305_ (.B1(_1014_),
    .Y(_1026_),
    .A1(_1024_),
    .A2(_1025_));
 sg13g2_xor2_1 _3306_ (.B(_1010_),
    .A(net927),
    .X(_1027_));
 sg13g2_a21oi_2 _3307_ (.B1(_1011_),
    .Y(_1028_),
    .A2(_1027_),
    .A1(_1026_));
 sg13g2_nor2_1 _3308_ (.A(net661),
    .B(_0986_),
    .Y(_1029_));
 sg13g2_xnor2_1 _3309_ (.Y(_1030_),
    .A(_0989_),
    .B(_1029_));
 sg13g2_nand2_1 _3310_ (.Y(_1031_),
    .A(\systolic_array.genblk1[10].accumulators_dlygate[4].A ),
    .B(_1030_));
 sg13g2_xnor2_1 _3311_ (.Y(_1032_),
    .A(\systolic_array.genblk1[10].accumulators_dlygate[4].A ),
    .B(_1030_));
 sg13g2_nor3_2 _3312_ (.A(_1008_),
    .B(_1028_),
    .C(_1032_),
    .Y(_1033_));
 sg13g2_or3_1 _3313_ (.A(net661),
    .B(_0995_),
    .C(_0997_),
    .X(_1034_));
 sg13g2_o21ai_1 _3314_ (.B1(_0997_),
    .Y(_1035_),
    .A1(net661),
    .A2(_0995_));
 sg13g2_and2_1 _3315_ (.A(_1034_),
    .B(_1035_),
    .X(_1036_));
 sg13g2_a21oi_1 _3316_ (.A1(_1034_),
    .A2(_1035_),
    .Y(_1037_),
    .B1(\systolic_array.genblk1[10].accumulators_dlygate[7].A ));
 sg13g2_a21oi_1 _3317_ (.A1(_0991_),
    .A2(_0993_),
    .Y(_1038_),
    .B1(net661));
 sg13g2_xnor2_1 _3318_ (.Y(_1039_),
    .A(_0994_),
    .B(_1038_));
 sg13g2_nor3_1 _3319_ (.A(_1519_),
    .B(_1037_),
    .C(_1039_),
    .Y(_1040_));
 sg13g2_and2_1 _3320_ (.A(\systolic_array.genblk1[10].accumulators_dlygate[7].A ),
    .B(_1036_),
    .X(_1041_));
 sg13g2_nand2_1 _3321_ (.Y(_1042_),
    .A(\systolic_array.genblk1[10].accumulators_dlygate[7].A ),
    .B(_1036_));
 sg13g2_o21ai_1 _3322_ (.B1(_1007_),
    .Y(_1043_),
    .A1(_1006_),
    .A2(_1031_));
 sg13g2_or3_1 _3323_ (.A(_1040_),
    .B(_1041_),
    .C(_1043_),
    .X(_1044_));
 sg13g2_and2_1 _3324_ (.A(_1519_),
    .B(_1039_),
    .X(_1045_));
 sg13g2_o21ai_1 _3325_ (.B1(_1042_),
    .Y(_1046_),
    .A1(_1037_),
    .A2(_1045_));
 sg13g2_o21ai_1 _3326_ (.B1(_1046_),
    .Y(_1047_),
    .A1(_1033_),
    .A2(_1044_));
 sg13g2_a21oi_1 _3327_ (.A1(net554),
    .A2(_1002_),
    .Y(_1048_),
    .B1(\systolic_array.genblk1[10].accumulators_dlygate[8].A ));
 sg13g2_or2_1 _3328_ (.X(_1049_),
    .B(_1048_),
    .A(_1003_));
 sg13g2_nor2_1 _3329_ (.A(_1047_),
    .B(_1049_),
    .Y(_1050_));
 sg13g2_nor2_1 _3330_ (.A(_1003_),
    .B(_1050_),
    .Y(_1051_));
 sg13g2_xnor2_1 _3331_ (.Y(_1052_),
    .A(_1518_),
    .B(net554));
 sg13g2_nand2b_1 _3332_ (.Y(_1053_),
    .B(net648),
    .A_N(net827));
 sg13g2_xor2_1 _3333_ (.B(_1052_),
    .A(_1051_),
    .X(_1054_));
 sg13g2_o21ai_1 _3334_ (.B1(_1053_),
    .Y(_1055_),
    .A1(net648),
    .A2(_1054_));
 sg13g2_o21ai_1 _3335_ (.B1(_0978_),
    .Y(_0023_),
    .A1(net609),
    .A2(_1055_));
 sg13g2_nand2_1 _3336_ (.Y(_1056_),
    .A(net746),
    .B(net608));
 sg13g2_a21oi_2 _3337_ (.B1(_1003_),
    .Y(_1057_),
    .A2(net554),
    .A1(_1518_));
 sg13g2_nor2_1 _3338_ (.A(_1049_),
    .B(_1052_),
    .Y(_1058_));
 sg13g2_nand2b_1 _3339_ (.Y(_1059_),
    .B(_1058_),
    .A_N(_1047_));
 sg13g2_nand2_1 _3340_ (.Y(_1060_),
    .A(\systolic_array.genblk1[10].accumulators_dlygate[10].A ),
    .B(net553));
 sg13g2_xnor2_1 _3341_ (.Y(_1061_),
    .A(\systolic_array.genblk1[10].accumulators_dlygate[10].A ),
    .B(net553));
 sg13g2_a21o_1 _3342_ (.A2(_1059_),
    .A1(_1057_),
    .B1(_1061_),
    .X(_1062_));
 sg13g2_and3_1 _3343_ (.X(_1063_),
    .A(_1057_),
    .B(_1059_),
    .C(_1061_));
 sg13g2_nor2_1 _3344_ (.A(net647),
    .B(_1063_),
    .Y(_1064_));
 sg13g2_a22oi_1 _3345_ (.Y(_1065_),
    .B1(_1062_),
    .B2(_1064_),
    .A2(net976),
    .A1(net648));
 sg13g2_o21ai_1 _3346_ (.B1(_1056_),
    .Y(_0016_),
    .A1(net608),
    .A2(_1065_));
 sg13g2_nand2_1 _3347_ (.Y(_1066_),
    .A(net761),
    .B(net607));
 sg13g2_nand2b_1 _3348_ (.Y(_1067_),
    .B(net552),
    .A_N(_0112_));
 sg13g2_xor2_1 _3349_ (.B(net553),
    .A(_0112_),
    .X(_1068_));
 sg13g2_a21oi_1 _3350_ (.A1(_1060_),
    .A2(_1062_),
    .Y(_1069_),
    .B1(_1068_));
 sg13g2_and3_1 _3351_ (.X(_1070_),
    .A(_1060_),
    .B(_1062_),
    .C(_1068_));
 sg13g2_nor3_1 _3352_ (.A(net647),
    .B(_1069_),
    .C(_1070_),
    .Y(_1071_));
 sg13g2_a21oi_2 _3353_ (.B1(_1071_),
    .Y(_1072_),
    .A2(net893),
    .A1(net647));
 sg13g2_o21ai_1 _3354_ (.B1(_1066_),
    .Y(_0017_),
    .A1(net606),
    .A2(_1072_));
 sg13g2_nand2_1 _3355_ (.Y(_1073_),
    .A(net757),
    .B(net606));
 sg13g2_nand3_1 _3356_ (.B(_1060_),
    .C(_1067_),
    .A(_1057_),
    .Y(_1074_));
 sg13g2_inv_1 _3357_ (.Y(_1075_),
    .A(_1074_));
 sg13g2_nor2_1 _3358_ (.A(_1061_),
    .B(_1068_),
    .Y(_1076_));
 sg13g2_nand3b_1 _3359_ (.B(_1058_),
    .C(_1076_),
    .Y(_1077_),
    .A_N(_1047_));
 sg13g2_nand2_1 _3360_ (.Y(_1078_),
    .A(_1075_),
    .B(_1077_));
 sg13g2_and2_1 _3361_ (.A(\systolic_array.genblk1[10].accumulators_dlygate[12].A ),
    .B(net552),
    .X(_1079_));
 sg13g2_xor2_1 _3362_ (.B(net552),
    .A(\systolic_array.genblk1[10].accumulators_dlygate[12].A ),
    .X(_1080_));
 sg13g2_o21ai_1 _3363_ (.B1(net618),
    .Y(_1081_),
    .A1(_1078_),
    .A2(_1080_));
 sg13g2_a21oi_1 _3364_ (.A1(_1078_),
    .A2(_1080_),
    .Y(_1082_),
    .B1(_1081_));
 sg13g2_a21oi_1 _3365_ (.A1(net647),
    .A2(net986),
    .Y(_1083_),
    .B1(_1082_));
 sg13g2_o21ai_1 _3366_ (.B1(_1073_),
    .Y(_0018_),
    .A1(net606),
    .A2(_1083_));
 sg13g2_nand2_1 _3367_ (.Y(_1084_),
    .A(net738),
    .B(net606));
 sg13g2_xnor2_1 _3368_ (.Y(_1085_),
    .A(_0113_),
    .B(net552));
 sg13g2_a21oi_1 _3369_ (.A1(_1078_),
    .A2(_1080_),
    .Y(_1086_),
    .B1(_1079_));
 sg13g2_nand2b_1 _3370_ (.Y(_1087_),
    .B(net647),
    .A_N(net741));
 sg13g2_xnor2_1 _3371_ (.Y(_1088_),
    .A(_1085_),
    .B(_1086_));
 sg13g2_o21ai_1 _3372_ (.B1(_1087_),
    .Y(_1089_),
    .A1(net647),
    .A2(_1088_));
 sg13g2_o21ai_1 _3373_ (.B1(_1084_),
    .Y(_0019_),
    .A1(net606),
    .A2(_1089_));
 sg13g2_nand2_1 _3374_ (.Y(_1090_),
    .A(net533),
    .B(net607));
 sg13g2_nand2_1 _3375_ (.Y(_1091_),
    .A(\systolic_array.genblk1[10].accumulators_dlygate[14].A ),
    .B(net552));
 sg13g2_xor2_1 _3376_ (.B(net552),
    .A(\systolic_array.genblk1[10].accumulators_dlygate[14].A ),
    .X(_1092_));
 sg13g2_o21ai_1 _3377_ (.B1(net552),
    .Y(_1093_),
    .A1(\systolic_array.genblk1[10].accumulators_dlygate[12].A ),
    .A2(_1522_));
 sg13g2_inv_1 _3378_ (.Y(_1094_),
    .A(_1093_));
 sg13g2_nand2_1 _3379_ (.Y(_1095_),
    .A(_1080_),
    .B(_1085_));
 sg13g2_a21oi_1 _3380_ (.A1(_1075_),
    .A2(_1077_),
    .Y(_1096_),
    .B1(_1095_));
 sg13g2_o21ai_1 _3381_ (.B1(_1092_),
    .Y(_1097_),
    .A1(_1094_),
    .A2(_1096_));
 sg13g2_nor3_1 _3382_ (.A(_1092_),
    .B(_1094_),
    .C(_1096_),
    .Y(_1098_));
 sg13g2_nor2_1 _3383_ (.A(net647),
    .B(_1098_),
    .Y(_1099_));
 sg13g2_a22oi_1 _3384_ (.Y(_1100_),
    .B1(_1097_),
    .B2(_1099_),
    .A2(net959),
    .A1(net647));
 sg13g2_o21ai_1 _3385_ (.B1(_1090_),
    .Y(_0020_),
    .A1(net607),
    .A2(_1100_));
 sg13g2_nand2_1 _3386_ (.Y(_1101_),
    .A(net730),
    .B(net607));
 sg13g2_nand2b_1 _3387_ (.Y(_1102_),
    .B(net648),
    .A_N(net954));
 sg13g2_xor2_1 _3388_ (.B(net553),
    .A(\systolic_array.genblk1[10].accumulators_dlygate[15].A ),
    .X(_1103_));
 sg13g2_nand2_1 _3389_ (.Y(_1104_),
    .A(_1091_),
    .B(_1097_));
 sg13g2_xor2_1 _3390_ (.B(_1104_),
    .A(_1103_),
    .X(_1105_));
 sg13g2_o21ai_1 _3391_ (.B1(_1102_),
    .Y(_1106_),
    .A1(net648),
    .A2(_1105_));
 sg13g2_o21ai_1 _3392_ (.B1(_1101_),
    .Y(_0021_),
    .A1(net609),
    .A2(_1106_));
 sg13g2_nand2_1 _3393_ (.Y(_1107_),
    .A(net760),
    .B(net610));
 sg13g2_nand2_1 _3394_ (.Y(_1108_),
    .A(_1092_),
    .B(_1103_));
 sg13g2_or3_1 _3395_ (.A(_1077_),
    .B(_1095_),
    .C(_1108_),
    .X(_1109_));
 sg13g2_o21ai_1 _3396_ (.B1(net552),
    .Y(_1110_),
    .A1(\systolic_array.genblk1[10].accumulators_dlygate[14].A ),
    .A2(\systolic_array.genblk1[10].accumulators_dlygate[15].A ));
 sg13g2_nand4_1 _3397_ (.B(_1093_),
    .C(_1109_),
    .A(_1075_),
    .Y(_1111_),
    .D(_1110_));
 sg13g2_a21oi_1 _3398_ (.A1(net554),
    .A2(_1111_),
    .Y(_1112_),
    .B1(net648));
 sg13g2_o21ai_1 _3399_ (.B1(_1112_),
    .Y(_1113_),
    .A1(net554),
    .A2(_1111_));
 sg13g2_xor2_1 _3400_ (.B(_1113_),
    .A(net778),
    .X(_1114_));
 sg13g2_o21ai_1 _3401_ (.B1(_1107_),
    .Y(_0022_),
    .A1(net610),
    .A2(_1114_));
 sg13g2_mux2_1 _3402_ (.A0(net530),
    .A1(net919),
    .S(net641),
    .X(_0000_));
 sg13g2_mux2_1 _3403_ (.A0(net494),
    .A1(net860),
    .S(net641),
    .X(_0001_));
 sg13g2_mux2_1 _3404_ (.A0(net774),
    .A1(net878),
    .S(net641),
    .X(_0002_));
 sg13g2_mux2_1 _3405_ (.A0(net433),
    .A1(net721),
    .S(net645),
    .X(_0003_));
 sg13g2_mux2_1 _3406_ (.A0(net483),
    .A1(net804),
    .S(net644),
    .X(_0004_));
 sg13g2_mux2_2 _3407_ (.A0(net514),
    .A1(net955),
    .S(net643),
    .X(_0005_));
 sg13g2_mux2_2 _3408_ (.A0(net520),
    .A1(net912),
    .S(net643),
    .X(_0006_));
 sg13g2_mux2_2 _3409_ (.A0(net497),
    .A1(net929),
    .S(net643),
    .X(_0007_));
 sg13g2_nand2_2 _3410_ (.Y(_1115_),
    .A(net719),
    .B(net697));
 sg13g2_nor2_1 _3411_ (.A(net712),
    .B(net714),
    .Y(_1116_));
 sg13g2_o21ai_1 _3412_ (.B1(net711),
    .Y(_1117_),
    .A1(net712),
    .A2(net714));
 sg13g2_nor2b_2 _3413_ (.A(net710),
    .B_N(_1117_),
    .Y(_1118_));
 sg13g2_nand2b_1 _3414_ (.Y(_1119_),
    .B(_1117_),
    .A_N(net708));
 sg13g2_nand3_1 _3415_ (.B(net704),
    .C(_1119_),
    .A(net701),
    .Y(_1120_));
 sg13g2_and2_1 _3416_ (.A(net698),
    .B(_1120_),
    .X(_1121_));
 sg13g2_nand2_1 _3417_ (.Y(_1122_),
    .A(net698),
    .B(_1120_));
 sg13g2_nor2_2 _3418_ (.A(net702),
    .B(net707),
    .Y(_1123_));
 sg13g2_nand2_1 _3419_ (.Y(_1124_),
    .A(_1532_),
    .B(_1123_));
 sg13g2_nand2_1 _3420_ (.Y(_1125_),
    .A(net694),
    .B(_1124_));
 sg13g2_a21oi_1 _3421_ (.A1(_1122_),
    .A2(_1125_),
    .Y(_0120_),
    .B1(_1115_));
 sg13g2_o21ai_1 _3422_ (.B1(_0978_),
    .Y(_0121_),
    .A1(_1523_),
    .A2(net609));
 sg13g2_o21ai_1 _3423_ (.B1(_1056_),
    .Y(_0122_),
    .A1(_1524_),
    .A2(net606));
 sg13g2_o21ai_1 _3424_ (.B1(_1066_),
    .Y(_0123_),
    .A1(_1525_),
    .A2(net607));
 sg13g2_o21ai_1 _3425_ (.B1(_1073_),
    .Y(_0124_),
    .A1(_1526_),
    .A2(net606));
 sg13g2_o21ai_1 _3426_ (.B1(_1084_),
    .Y(_0125_),
    .A1(_1527_),
    .A2(net606));
 sg13g2_o21ai_1 _3427_ (.B1(_1090_),
    .Y(_0126_),
    .A1(_1528_),
    .A2(net609));
 sg13g2_o21ai_1 _3428_ (.B1(_1101_),
    .Y(_0127_),
    .A1(_1529_),
    .A2(net607));
 sg13g2_o21ai_1 _3429_ (.B1(_1107_),
    .Y(_0128_),
    .A1(_1530_),
    .A2(net610));
 sg13g2_and2_1 _3430_ (.A(net715),
    .B(net530),
    .X(_0129_));
 sg13g2_and2_1 _3431_ (.A(net715),
    .B(net494),
    .X(_0130_));
 sg13g2_and2_1 _3432_ (.A(net715),
    .B(net774),
    .X(_0131_));
 sg13g2_and2_1 _3433_ (.A(net720),
    .B(net433),
    .X(_0132_));
 sg13g2_and2_1 _3434_ (.A(net718),
    .B(net483),
    .X(_0133_));
 sg13g2_and2_1 _3435_ (.A(net717),
    .B(net514),
    .X(_0134_));
 sg13g2_and2_1 _3436_ (.A(net717),
    .B(net520),
    .X(_0135_));
 sg13g2_and2_1 _3437_ (.A(net717),
    .B(net497),
    .X(_0136_));
 sg13g2_and2_1 _3438_ (.A(net720),
    .B(net7),
    .X(_0137_));
 sg13g2_and2_1 _3439_ (.A(net720),
    .B(net8),
    .X(_0138_));
 sg13g2_and2_1 _3440_ (.A(net718),
    .B(net9),
    .X(_0139_));
 sg13g2_and2_1 _3441_ (.A(net717),
    .B(net10),
    .X(_0140_));
 sg13g2_and2_1 _3442_ (.A(net717),
    .B(net11),
    .X(_0141_));
 sg13g2_and2_1 _3443_ (.A(net717),
    .B(net12),
    .X(_0142_));
 sg13g2_and2_1 _3444_ (.A(net717),
    .B(net13),
    .X(_0143_));
 sg13g2_and2_1 _3445_ (.A(net717),
    .B(net14),
    .X(_0144_));
 sg13g2_and2_1 _3446_ (.A(net715),
    .B(net945),
    .X(_0145_));
 sg13g2_and2_1 _3447_ (.A(net715),
    .B(net970),
    .X(_0146_));
 sg13g2_and2_1 _3448_ (.A(net716),
    .B(net822),
    .X(_0147_));
 sg13g2_and2_1 _3449_ (.A(net718),
    .B(net780),
    .X(_0148_));
 sg13g2_and2_1 _3450_ (.A(net715),
    .B(net908),
    .X(_0149_));
 sg13g2_and2_1 _3451_ (.A(net716),
    .B(net832),
    .X(_0150_));
 sg13g2_nor2b_1 _3452_ (.A(net641),
    .B_N(net482),
    .Y(_0151_));
 sg13g2_nor2b_1 _3453_ (.A(net640),
    .B_N(net477),
    .Y(_0152_));
 sg13g2_nor2b_1 _3454_ (.A(net640),
    .B_N(net500),
    .Y(_0153_));
 sg13g2_nor2b_1 _3455_ (.A(net645),
    .B_N(net512),
    .Y(_0154_));
 sg13g2_nor2b_1 _3456_ (.A(net643),
    .B_N(net471),
    .Y(_0155_));
 sg13g2_nor2b_1 _3457_ (.A(net643),
    .B_N(net442),
    .Y(_0156_));
 sg13g2_nor2b_1 _3458_ (.A(net643),
    .B_N(net461),
    .Y(_0157_));
 sg13g2_nor2b_1 _3459_ (.A(net643),
    .B_N(net473),
    .Y(_0158_));
 sg13g2_and2_1 _3460_ (.A(net716),
    .B(net920),
    .X(_0159_));
 sg13g2_and2_1 _3461_ (.A(net715),
    .B(net800),
    .X(_0160_));
 sg13g2_mux2_1 _3462_ (.A0(net752),
    .A1(\systolic_array.genblk2[0].mac[0].mul2 ),
    .S(net640),
    .X(_0161_));
 sg13g2_nor2_1 _3463_ (.A(net639),
    .B(net543),
    .Y(_1126_));
 sg13g2_a21oi_1 _3464_ (.A1(net639),
    .A2(_1480_),
    .Y(_0162_),
    .B1(_1126_));
 sg13g2_mux2_1 _3465_ (.A0(net750),
    .A1(net670),
    .S(net640),
    .X(_0163_));
 sg13g2_nor2_1 _3466_ (.A(net638),
    .B(net890),
    .Y(_1127_));
 sg13g2_a21oi_1 _3467_ (.A1(net638),
    .A2(_1500_),
    .Y(_0164_),
    .B1(_1127_));
 sg13g2_nor2_1 _3468_ (.A(net637),
    .B(net977),
    .Y(_1128_));
 sg13g2_a21oi_1 _3469_ (.A1(net637),
    .A2(_1509_),
    .Y(_0165_),
    .B1(_1128_));
 sg13g2_mux2_1 _3470_ (.A0(net866),
    .A1(net664),
    .S(net638),
    .X(_0166_));
 sg13g2_nor2_1 _3471_ (.A(net644),
    .B(net793),
    .Y(_1129_));
 sg13g2_a21oi_1 _3472_ (.A1(net644),
    .A2(_1471_),
    .Y(_0167_),
    .B1(_1129_));
 sg13g2_nor2_1 _3473_ (.A(net639),
    .B(net772),
    .Y(_1130_));
 sg13g2_a21oi_1 _3474_ (.A1(net639),
    .A2(_1482_),
    .Y(_0168_),
    .B1(_1130_));
 sg13g2_nor2_1 _3475_ (.A(net640),
    .B(net536),
    .Y(_1131_));
 sg13g2_a21oi_1 _3476_ (.A1(net640),
    .A2(_1493_),
    .Y(_0169_),
    .B1(_1131_));
 sg13g2_nor2_1 _3477_ (.A(net637),
    .B(net945),
    .Y(_1132_));
 sg13g2_a21oi_1 _3478_ (.A1(net637),
    .A2(_1502_),
    .Y(_0170_),
    .B1(_1132_));
 sg13g2_nor2_1 _3479_ (.A(net637),
    .B(net970),
    .Y(_1133_));
 sg13g2_a21oi_1 _3480_ (.A1(net637),
    .A2(_1510_),
    .Y(_0171_),
    .B1(_1133_));
 sg13g2_nor2_1 _3481_ (.A(net638),
    .B(net822),
    .Y(_1134_));
 sg13g2_a21oi_1 _3482_ (.A1(net646),
    .A2(_1517_),
    .Y(_0172_),
    .B1(_1134_));
 sg13g2_nor2_1 _3483_ (.A(net644),
    .B(net777),
    .Y(_1135_));
 sg13g2_a21oi_1 _3484_ (.A1(net643),
    .A2(net630),
    .Y(_0173_),
    .B1(_1135_));
 sg13g2_nor2_1 _3485_ (.A(net642),
    .B(net833),
    .Y(_1136_));
 sg13g2_a21oi_1 _3486_ (.A1(net639),
    .A2(net628),
    .Y(_0174_),
    .B1(_1136_));
 sg13g2_nor2_1 _3487_ (.A(net640),
    .B(net538),
    .Y(_1137_));
 sg13g2_a21oi_1 _3488_ (.A1(net640),
    .A2(net625),
    .Y(_0175_),
    .B1(_1137_));
 sg13g2_nor2_2 _3489_ (.A(net645),
    .B(net780),
    .Y(_1138_));
 sg13g2_a21oi_1 _3490_ (.A1(net637),
    .A2(net623),
    .Y(_0176_),
    .B1(_1138_));
 sg13g2_nor2_2 _3491_ (.A(net642),
    .B(net908),
    .Y(_1139_));
 sg13g2_a21oi_1 _3492_ (.A1(net637),
    .A2(_1514_),
    .Y(_0177_),
    .B1(_1139_));
 sg13g2_nor2_1 _3493_ (.A(net646),
    .B(net832),
    .Y(_1140_));
 sg13g2_a21oi_1 _3494_ (.A1(net638),
    .A2(net616),
    .Y(_0178_),
    .B1(_1140_));
 sg13g2_and2_1 _3495_ (.A(net716),
    .B(net890),
    .X(_0179_));
 sg13g2_and2_1 _3496_ (.A(net715),
    .B(net977),
    .X(_0180_));
 sg13g2_and2_1 _3497_ (.A(net716),
    .B(net866),
    .X(_0181_));
 sg13g2_nor2_1 _3498_ (.A(net709),
    .B(net711),
    .Y(_1141_));
 sg13g2_a21oi_2 _3499_ (.B1(net711),
    .Y(_1142_),
    .A2(net713),
    .A1(net712));
 sg13g2_and2_1 _3500_ (.A(_1539_),
    .B(_1141_),
    .X(_1143_));
 sg13g2_nor2_1 _3501_ (.A(net709),
    .B(net704),
    .Y(_1144_));
 sg13g2_a21oi_2 _3502_ (.B1(net695),
    .Y(_1145_),
    .A2(_1144_),
    .A1(_1142_));
 sg13g2_or3_1 _3503_ (.A(net697),
    .B(net698),
    .C(_1145_),
    .X(_1146_));
 sg13g2_nand2_1 _3504_ (.Y(_1147_),
    .A(_1538_),
    .B(_1122_));
 sg13g2_a21oi_1 _3505_ (.A1(_1146_),
    .A2(_1147_),
    .Y(_0182_),
    .B1(_1460_));
 sg13g2_nand2_1 _3506_ (.Y(_1148_),
    .A(net713),
    .B(_1533_));
 sg13g2_a21oi_2 _3507_ (.B1(net709),
    .Y(_1149_),
    .A2(_1533_),
    .A1(net714));
 sg13g2_or2_1 _3508_ (.X(_1150_),
    .B(net711),
    .A(net712));
 sg13g2_inv_1 _3509_ (.Y(_1151_),
    .A(_1150_));
 sg13g2_nand3_1 _3510_ (.B(_1149_),
    .C(net693),
    .A(net704),
    .Y(_1152_));
 sg13g2_o21ai_1 _3511_ (.B1(_1121_),
    .Y(_1153_),
    .A1(net701),
    .A2(_1152_));
 sg13g2_o21ai_1 _3512_ (.B1(net704),
    .Y(_1154_),
    .A1(net708),
    .A2(net711));
 sg13g2_o21ai_1 _3513_ (.B1(_1463_),
    .Y(_1155_),
    .A1(_1532_),
    .A2(_1539_));
 sg13g2_nand2_1 _3514_ (.Y(_1156_),
    .A(net701),
    .B(_1155_));
 sg13g2_nand3_1 _3515_ (.B(_1154_),
    .C(_1155_),
    .A(net703),
    .Y(_1157_));
 sg13g2_nor2_1 _3516_ (.A(net695),
    .B(net698),
    .Y(_1158_));
 sg13g2_a21oi_1 _3517_ (.A1(_1463_),
    .A2(_1532_),
    .Y(_1159_),
    .B1(net701));
 sg13g2_nor2_1 _3518_ (.A(net698),
    .B(_1159_),
    .Y(_1160_));
 sg13g2_nor2_2 _3519_ (.A(net713),
    .B(net693),
    .Y(_1161_));
 sg13g2_nand2_1 _3520_ (.Y(_1162_),
    .A(net705),
    .B(net694));
 sg13g2_a21oi_1 _3521_ (.A1(_1116_),
    .A2(_1141_),
    .Y(_1163_),
    .B1(_1162_));
 sg13g2_o21ai_1 _3522_ (.B1(_1157_),
    .Y(_1164_),
    .A1(_1160_),
    .A2(_1163_));
 sg13g2_and3_1 _3523_ (.X(_1165_),
    .A(net697),
    .B(_1153_),
    .C(_1164_));
 sg13g2_nor2_2 _3524_ (.A(_1460_),
    .B(net697),
    .Y(_1166_));
 sg13g2_nor2b_2 _3525_ (.A(_1161_),
    .B_N(net710),
    .Y(_1167_));
 sg13g2_and2_1 _3526_ (.A(_1534_),
    .B(_1167_),
    .X(_1168_));
 sg13g2_nor2_2 _3527_ (.A(net695),
    .B(net705),
    .Y(_1169_));
 sg13g2_nand2_1 _3528_ (.Y(_1170_),
    .A(net702),
    .B(_1463_));
 sg13g2_nor2b_2 _3529_ (.A(_1142_),
    .B_N(net708),
    .Y(_1171_));
 sg13g2_nor2_2 _3530_ (.A(net708),
    .B(_1533_),
    .Y(_1172_));
 sg13g2_or3_1 _3531_ (.A(net704),
    .B(_1171_),
    .C(_1172_),
    .X(_1173_));
 sg13g2_nand2b_1 _3532_ (.Y(_1174_),
    .B(net695),
    .A_N(_1173_));
 sg13g2_nor2b_1 _3533_ (.A(_1142_),
    .B_N(_1144_),
    .Y(_1175_));
 sg13g2_a22oi_1 _3534_ (.Y(_1176_),
    .B1(_1175_),
    .B2(net703),
    .A2(_1123_),
    .A1(_1118_));
 sg13g2_a21oi_1 _3535_ (.A1(_1168_),
    .A2(_1169_),
    .Y(_1177_),
    .B1(net694));
 sg13g2_a221oi_1 _3536_ (.B2(_1174_),
    .C1(net697),
    .B1(_1177_),
    .A1(_1464_),
    .Y(_1178_),
    .A2(_1176_));
 sg13g2_o21ai_1 _3537_ (.B1(net719),
    .Y(_1179_),
    .A1(_1165_),
    .A2(_1178_));
 sg13g2_inv_1 _3538_ (.Y(_0183_),
    .A(_1179_));
 sg13g2_nor2b_2 _3539_ (.A(net713),
    .B_N(net3),
    .Y(_1180_));
 sg13g2_nand2b_2 _3540_ (.Y(_1181_),
    .B(net3),
    .A_N(net713));
 sg13g2_nand2b_2 _3541_ (.Y(_1182_),
    .B(net713),
    .A_N(net711));
 sg13g2_nor2b_2 _3542_ (.A(net710),
    .B_N(net712),
    .Y(_1183_));
 sg13g2_nor2_1 _3543_ (.A(_1182_),
    .B(_1183_),
    .Y(_1184_));
 sg13g2_nand2_1 _3544_ (.Y(_1185_),
    .A(_1181_),
    .B(_1183_));
 sg13g2_nand2_1 _3545_ (.Y(_1186_),
    .A(_1181_),
    .B(_1182_));
 sg13g2_nor2_1 _3546_ (.A(_1180_),
    .B(_1184_),
    .Y(_1187_));
 sg13g2_nor2b_2 _3547_ (.A(net2),
    .B_N(net710),
    .Y(_1188_));
 sg13g2_a21oi_1 _3548_ (.A1(_1182_),
    .A2(_1188_),
    .Y(_1189_),
    .B1(net707));
 sg13g2_and2_1 _3549_ (.A(_1182_),
    .B(_1183_),
    .X(_1190_));
 sg13g2_nor3_1 _3550_ (.A(_1180_),
    .B(_1184_),
    .C(_1190_),
    .Y(_1191_));
 sg13g2_nor2_1 _3551_ (.A(_1189_),
    .B(_1191_),
    .Y(_1192_));
 sg13g2_a21oi_1 _3552_ (.A1(_1182_),
    .A2(_1188_),
    .Y(_1193_),
    .B1(_1187_));
 sg13g2_a21oi_1 _3553_ (.A1(_1463_),
    .A2(_1187_),
    .Y(_1194_),
    .B1(_1192_));
 sg13g2_nor2_1 _3554_ (.A(_1180_),
    .B(_1188_),
    .Y(_1195_));
 sg13g2_o21ai_1 _3555_ (.B1(_1185_),
    .Y(_1196_),
    .A1(_1183_),
    .A2(_1195_));
 sg13g2_xnor2_1 _3556_ (.Y(_1197_),
    .A(net702),
    .B(_1196_));
 sg13g2_and2_1 _3557_ (.A(_1194_),
    .B(_1197_),
    .X(_1198_));
 sg13g2_nor2_1 _3558_ (.A(net700),
    .B(_1198_),
    .Y(_1199_));
 sg13g2_nand2b_1 _3559_ (.Y(_1200_),
    .B(_1184_),
    .A_N(_1188_));
 sg13g2_nand2_1 _3560_ (.Y(_1201_),
    .A(_1180_),
    .B(_1188_));
 sg13g2_nand3b_1 _3561_ (.B(_1200_),
    .C(_1201_),
    .Y(_1202_),
    .A_N(_1190_));
 sg13g2_inv_1 _3562_ (.Y(_1203_),
    .A(_1202_));
 sg13g2_a22oi_1 _3563_ (.Y(_1204_),
    .B1(_1203_),
    .B2(net707),
    .A2(_1189_),
    .A1(_1185_));
 sg13g2_nand2_1 _3564_ (.Y(_1205_),
    .A(_1181_),
    .B(_1188_));
 sg13g2_and2_1 _3565_ (.A(_1182_),
    .B(_1205_),
    .X(_1206_));
 sg13g2_and2_1 _3566_ (.A(net708),
    .B(net693),
    .X(_1207_));
 sg13g2_o21ai_1 _3567_ (.B1(_1206_),
    .Y(_1208_),
    .A1(_1181_),
    .A2(_1188_));
 sg13g2_nand2_1 _3568_ (.Y(_1209_),
    .A(net707),
    .B(_1193_));
 sg13g2_o21ai_1 _3569_ (.B1(_1209_),
    .Y(_1210_),
    .A1(net707),
    .A2(_1208_));
 sg13g2_nor2_1 _3570_ (.A(net707),
    .B(_1202_),
    .Y(_1211_));
 sg13g2_a21oi_1 _3571_ (.A1(net707),
    .A2(_1196_),
    .Y(_1212_),
    .B1(_1211_));
 sg13g2_nor3_1 _3572_ (.A(net702),
    .B(_1204_),
    .C(_1212_),
    .Y(_1213_));
 sg13g2_a21oi_1 _3573_ (.A1(net702),
    .A2(_1204_),
    .Y(_1214_),
    .B1(_1213_));
 sg13g2_nor2_2 _3574_ (.A(net702),
    .B(_1463_),
    .Y(_1215_));
 sg13g2_o21ai_1 _3575_ (.B1(_1182_),
    .Y(_1216_),
    .A1(net713),
    .A2(_1534_));
 sg13g2_nor2_1 _3576_ (.A(net710),
    .B(_1216_),
    .Y(_1217_));
 sg13g2_o21ai_1 _3577_ (.B1(_1217_),
    .Y(_1218_),
    .A1(net2),
    .A2(_1180_));
 sg13g2_nand3_1 _3578_ (.B(_1539_),
    .C(_1186_),
    .A(net710),
    .Y(_1219_));
 sg13g2_nand2_1 _3579_ (.Y(_1220_),
    .A(_1218_),
    .B(_1219_));
 sg13g2_nand3_1 _3580_ (.B(_1534_),
    .C(net693),
    .A(net713),
    .Y(_1221_));
 sg13g2_o21ai_1 _3581_ (.B1(_1169_),
    .Y(_1222_),
    .A1(net4),
    .A2(_1216_));
 sg13g2_a21oi_1 _3582_ (.A1(_1167_),
    .A2(_1221_),
    .Y(_1223_),
    .B1(_1222_));
 sg13g2_a221oi_1 _3583_ (.B2(_1220_),
    .C1(_1223_),
    .B1(_1215_),
    .A1(_1123_),
    .Y(_1224_),
    .A2(_1191_));
 sg13g2_o21ai_1 _3584_ (.B1(_1224_),
    .Y(_1225_),
    .A1(_1537_),
    .A2(_1208_));
 sg13g2_and2_1 _3585_ (.A(net694),
    .B(_1225_),
    .X(_1226_));
 sg13g2_nand2b_1 _3586_ (.Y(_1227_),
    .B(_1226_),
    .A_N(_1214_));
 sg13g2_a21oi_1 _3587_ (.A1(net700),
    .A2(_1198_),
    .Y(_1228_),
    .B1(net6));
 sg13g2_a21oi_1 _3588_ (.A1(_1180_),
    .A2(_1183_),
    .Y(_1229_),
    .B1(_1170_));
 sg13g2_o21ai_1 _3589_ (.B1(_1123_),
    .Y(_1230_),
    .A1(_1184_),
    .A2(_1206_));
 sg13g2_nor2_1 _3590_ (.A(_1537_),
    .B(_1161_),
    .Y(_1231_));
 sg13g2_nand2_1 _3591_ (.Y(_1232_),
    .A(_1181_),
    .B(_1190_));
 sg13g2_nand3_1 _3592_ (.B(_1215_),
    .C(_1232_),
    .A(_1201_),
    .Y(_1233_));
 sg13g2_nand2_1 _3593_ (.Y(_1234_),
    .A(_1230_),
    .B(_1233_));
 sg13g2_a221oi_1 _3594_ (.B2(_1118_),
    .C1(_1234_),
    .B1(_1231_),
    .A1(_1200_),
    .Y(_1235_),
    .A2(_1229_));
 sg13g2_nor2_1 _3595_ (.A(net694),
    .B(_1235_),
    .Y(_1236_));
 sg13g2_xnor2_1 _3596_ (.Y(_1237_),
    .A(net696),
    .B(_1202_));
 sg13g2_a21oi_1 _3597_ (.A1(_1210_),
    .A2(_1237_),
    .Y(_1238_),
    .B1(net700));
 sg13g2_o21ai_1 _3598_ (.B1(net697),
    .Y(_1239_),
    .A1(_1236_),
    .A2(_1238_));
 sg13g2_nand2_1 _3599_ (.Y(_1240_),
    .A(net719),
    .B(_1239_));
 sg13g2_a21oi_1 _3600_ (.A1(_1227_),
    .A2(_1228_),
    .Y(_0184_),
    .B1(_1240_));
 sg13g2_or2_1 _3601_ (.X(_1241_),
    .B(_1143_),
    .A(net704));
 sg13g2_nor2_1 _3602_ (.A(net708),
    .B(net693),
    .Y(_1242_));
 sg13g2_a21oi_1 _3603_ (.A1(net704),
    .A2(_1242_),
    .Y(_1243_),
    .B1(net703));
 sg13g2_a22oi_1 _3604_ (.Y(_1244_),
    .B1(_1241_),
    .B2(_1243_),
    .A2(_1172_),
    .A1(_1169_));
 sg13g2_a22oi_1 _3605_ (.Y(_1245_),
    .B1(_1244_),
    .B2(_1121_),
    .A2(_1160_),
    .A1(_1156_));
 sg13g2_nor2_2 _3606_ (.A(_1532_),
    .B(_1116_),
    .Y(_1246_));
 sg13g2_nor3_1 _3607_ (.A(net706),
    .B(_1168_),
    .C(_1246_),
    .Y(_1247_));
 sg13g2_nand2_1 _3608_ (.Y(_1248_),
    .A(net701),
    .B(_1247_));
 sg13g2_nand2_1 _3609_ (.Y(_1249_),
    .A(_1123_),
    .B(_1172_));
 sg13g2_a22oi_1 _3610_ (.Y(_1250_),
    .B1(_1246_),
    .B2(_1536_),
    .A2(_1215_),
    .A1(_1207_));
 sg13g2_nand4_1 _3611_ (.B(_1248_),
    .C(_1249_),
    .A(net698),
    .Y(_1251_),
    .D(_1250_));
 sg13g2_a22oi_1 _3612_ (.Y(_1252_),
    .B1(_1154_),
    .B2(net696),
    .A2(_1149_),
    .A1(_1145_));
 sg13g2_a21o_1 _3613_ (.A2(_1252_),
    .A1(_1241_),
    .B1(net698),
    .X(_1253_));
 sg13g2_nand3_1 _3614_ (.B(_1251_),
    .C(_1253_),
    .A(_1166_),
    .Y(_1254_));
 sg13g2_o21ai_1 _3615_ (.B1(_1254_),
    .Y(_0185_),
    .A1(_1115_),
    .A2(_1245_));
 sg13g2_xor2_1 _3616_ (.B(_1226_),
    .A(_1214_),
    .X(_1255_));
 sg13g2_o21ai_1 _3617_ (.B1(net719),
    .Y(_1256_),
    .A1(_1461_),
    .A2(_1255_));
 sg13g2_a21oi_1 _3618_ (.A1(_1239_),
    .A2(_1255_),
    .Y(_0186_),
    .B1(_1256_));
 sg13g2_nor2_1 _3619_ (.A(net695),
    .B(net694),
    .Y(_1257_));
 sg13g2_nand2_1 _3620_ (.Y(_1258_),
    .A(net719),
    .B(_1257_));
 sg13g2_o21ai_1 _3621_ (.B1(_1115_),
    .Y(_1259_),
    .A1(_1247_),
    .A2(_1258_));
 sg13g2_a21oi_1 _3622_ (.A1(net706),
    .A2(_1119_),
    .Y(_1260_),
    .B1(net701));
 sg13g2_nand2_1 _3623_ (.Y(_1261_),
    .A(_1152_),
    .B(_1260_));
 sg13g2_o21ai_1 _3624_ (.B1(_1261_),
    .Y(_1262_),
    .A1(_1461_),
    .A2(_1121_));
 sg13g2_o21ai_1 _3625_ (.B1(_1262_),
    .Y(_1263_),
    .A1(net700),
    .A2(_1124_));
 sg13g2_and2_1 _3626_ (.A(_1259_),
    .B(_1263_),
    .X(_0187_));
 sg13g2_o21ai_1 _3627_ (.B1(_1155_),
    .Y(_1264_),
    .A1(_1535_),
    .A2(_1154_));
 sg13g2_a22oi_1 _3628_ (.Y(_1265_),
    .B1(_1264_),
    .B2(net695),
    .A2(_1152_),
    .A1(_1145_));
 sg13g2_or2_1 _3629_ (.X(_1266_),
    .B(_1265_),
    .A(net699));
 sg13g2_a21oi_1 _3630_ (.A1(net709),
    .A2(net693),
    .Y(_1267_),
    .B1(_1118_));
 sg13g2_or3_1 _3631_ (.A(_1141_),
    .B(_1167_),
    .C(_1170_),
    .X(_1268_));
 sg13g2_nor2b_1 _3632_ (.A(_1161_),
    .B_N(_1172_),
    .Y(_1269_));
 sg13g2_nand2b_1 _3633_ (.Y(_1270_),
    .B(_1172_),
    .A_N(_1161_));
 sg13g2_nand3_1 _3634_ (.B(_1536_),
    .C(_1117_),
    .A(net708),
    .Y(_1271_));
 sg13g2_a22oi_1 _3635_ (.Y(_1272_),
    .B1(_1269_),
    .B2(_1123_),
    .A2(_1267_),
    .A1(_1215_));
 sg13g2_nand4_1 _3636_ (.B(_1268_),
    .C(_1271_),
    .A(net699),
    .Y(_1273_),
    .D(_1272_));
 sg13g2_nand3_1 _3637_ (.B(_1266_),
    .C(_1273_),
    .A(_1166_),
    .Y(_1274_));
 sg13g2_nand4_1 _3638_ (.B(_1148_),
    .C(net693),
    .A(net708),
    .Y(_1275_),
    .D(_1169_));
 sg13g2_o21ai_1 _3639_ (.B1(_1275_),
    .Y(_1276_),
    .A1(_1124_),
    .A2(_1149_));
 sg13g2_a221oi_1 _3640_ (.B2(_1215_),
    .C1(_1276_),
    .B1(_1171_),
    .A1(_1535_),
    .Y(_1277_),
    .A2(_1536_));
 sg13g2_nor2_1 _3641_ (.A(net699),
    .B(_1277_),
    .Y(_1278_));
 sg13g2_o21ai_1 _3642_ (.B1(_1463_),
    .Y(_1279_),
    .A1(_1143_),
    .A2(_1246_));
 sg13g2_a221oi_1 _3643_ (.B2(_1243_),
    .C1(_1122_),
    .B1(_1279_),
    .A1(_1169_),
    .Y(_1280_),
    .A2(_1270_));
 sg13g2_nor2_1 _3644_ (.A(_1278_),
    .B(_1280_),
    .Y(_1281_));
 sg13g2_o21ai_1 _3645_ (.B1(_1274_),
    .Y(_0188_),
    .A1(_1115_),
    .A2(_1281_));
 sg13g2_o21ai_1 _3646_ (.B1(_1461_),
    .Y(_1282_),
    .A1(_1199_),
    .A2(_1225_));
 sg13g2_nor2_1 _3647_ (.A(_1226_),
    .B(_1282_),
    .Y(_1283_));
 sg13g2_nand2_1 _3648_ (.Y(_1284_),
    .A(net702),
    .B(_1212_));
 sg13g2_xnor2_1 _3649_ (.Y(_1285_),
    .A(_1194_),
    .B(_1284_));
 sg13g2_nor2_1 _3650_ (.A(_1236_),
    .B(_1285_),
    .Y(_1286_));
 sg13g2_a21oi_1 _3651_ (.A1(net700),
    .A2(_1285_),
    .Y(_1287_),
    .B1(_1286_));
 sg13g2_a21oi_1 _3652_ (.A1(net6),
    .A2(_1287_),
    .Y(_1288_),
    .B1(_1283_));
 sg13g2_nor2_1 _3653_ (.A(_1460_),
    .B(_1288_),
    .Y(_0189_));
 sg13g2_nand2b_1 _3654_ (.Y(_1289_),
    .B(_1156_),
    .A_N(_1125_));
 sg13g2_nand2_1 _3655_ (.Y(_1290_),
    .A(net719),
    .B(_1146_));
 sg13g2_a221oi_1 _3656_ (.B2(net697),
    .C1(_1290_),
    .B1(_1289_),
    .A1(net700),
    .Y(_0190_),
    .A2(_1249_));
 sg13g2_nand3b_1 _3657_ (.B(net705),
    .C(_1532_),
    .Y(_1291_),
    .A_N(_1149_));
 sg13g2_nand3_1 _3658_ (.B(_1463_),
    .C(_1117_),
    .A(net709),
    .Y(_1292_));
 sg13g2_a21oi_1 _3659_ (.A1(_1291_),
    .A2(_1292_),
    .Y(_1293_),
    .B1(net695));
 sg13g2_nor2_1 _3660_ (.A(_1154_),
    .B(_1167_),
    .Y(_1294_));
 sg13g2_a221oi_1 _3661_ (.B2(net695),
    .C1(net699),
    .B1(_1294_),
    .A1(_1123_),
    .Y(_1295_),
    .A2(_1267_));
 sg13g2_nand2b_1 _3662_ (.Y(_1296_),
    .B(_1295_),
    .A_N(_1293_));
 sg13g2_a22oi_1 _3663_ (.Y(_1297_),
    .B1(_1171_),
    .B2(_1123_),
    .A2(_1169_),
    .A1(_1535_));
 sg13g2_o21ai_1 _3664_ (.B1(_1536_),
    .Y(_1298_),
    .A1(_1143_),
    .A2(_1246_));
 sg13g2_nand4_1 _3665_ (.B(_1148_),
    .C(net693),
    .A(net710),
    .Y(_1299_),
    .D(_1215_));
 sg13g2_nand4_1 _3666_ (.B(_1297_),
    .C(_1298_),
    .A(net699),
    .Y(_1300_),
    .D(_1299_));
 sg13g2_nand3_1 _3667_ (.B(_1296_),
    .C(_1300_),
    .A(_1166_),
    .Y(_1301_));
 sg13g2_a221oi_1 _3668_ (.B2(net705),
    .C1(net699),
    .B1(_1269_),
    .A1(_1144_),
    .Y(_1302_),
    .A2(_1151_));
 sg13g2_nor2_1 _3669_ (.A(net694),
    .B(_1175_),
    .Y(_1303_));
 sg13g2_a21oi_1 _3670_ (.A1(_1291_),
    .A2(_1303_),
    .Y(_1304_),
    .B1(_1302_));
 sg13g2_nor2_1 _3671_ (.A(net701),
    .B(_1304_),
    .Y(_1305_));
 sg13g2_o21ai_1 _3672_ (.B1(_1158_),
    .Y(_1306_),
    .A1(net704),
    .A2(_1119_));
 sg13g2_a21oi_1 _3673_ (.A1(_1173_),
    .A2(_1257_),
    .Y(_1307_),
    .B1(_1115_));
 sg13g2_o21ai_1 _3674_ (.B1(_1307_),
    .Y(_1308_),
    .A1(_1294_),
    .A2(_1306_));
 sg13g2_o21ai_1 _3675_ (.B1(_1301_),
    .Y(_0191_),
    .A1(_1305_),
    .A2(_1308_));
 sg13g2_nor2_1 _3676_ (.A(_1460_),
    .B(_1542_),
    .Y(_1309_));
 sg13g2_nand2_1 _3677_ (.Y(_1310_),
    .A(net719),
    .B(net615));
 sg13g2_nor3_1 _3678_ (.A(net644),
    .B(_1531_),
    .C(net566),
    .Y(_0192_));
 sg13g2_and2_1 _3679_ (.A(net444),
    .B(net595),
    .X(_0193_));
 sg13g2_and2_1 _3680_ (.A(net427),
    .B(net594),
    .X(_0194_));
 sg13g2_and2_1 _3681_ (.A(net429),
    .B(net594),
    .X(_0195_));
 sg13g2_and2_1 _3682_ (.A(net515),
    .B(net589),
    .X(_0196_));
 sg13g2_and2_1 _3683_ (.A(net501),
    .B(net594),
    .X(_0197_));
 sg13g2_and2_1 _3684_ (.A(net455),
    .B(net588),
    .X(_0198_));
 sg13g2_and2_1 _3685_ (.A(net459),
    .B(net588),
    .X(_0199_));
 sg13g2_and2_1 _3686_ (.A(net437),
    .B(net588),
    .X(_0200_));
 sg13g2_and2_1 _3687_ (.A(net415),
    .B(net588),
    .X(_0201_));
 sg13g2_and2_1 _3688_ (.A(net508),
    .B(net589),
    .X(_0202_));
 sg13g2_and2_1 _3689_ (.A(net481),
    .B(net588),
    .X(_0203_));
 sg13g2_and2_1 _3690_ (.A(net484),
    .B(net589),
    .X(_0204_));
 sg13g2_and2_1 _3691_ (.A(net440),
    .B(net587),
    .X(_0205_));
 sg13g2_and2_1 _3692_ (.A(net447),
    .B(net587),
    .X(_0206_));
 sg13g2_and2_1 _3693_ (.A(net478),
    .B(net587),
    .X(_0207_));
 sg13g2_and2_1 _3694_ (.A(net439),
    .B(net587),
    .X(_0208_));
 sg13g2_and2_1 _3695_ (.A(net510),
    .B(net587),
    .X(_0209_));
 sg13g2_nor2_1 _3696_ (.A(\systolic_array.genblk2[0].mac[0].zero ),
    .B(_1551_),
    .Y(_1311_));
 sg13g2_xnor2_1 _3697_ (.Y(_1312_),
    .A(net884),
    .B(_1311_));
 sg13g2_nor2_1 _3698_ (.A(net566),
    .B(net885),
    .Y(_0210_));
 sg13g2_xnor2_1 _3699_ (.Y(_1313_),
    .A(_1592_),
    .B(_1594_));
 sg13g2_o21ai_1 _3700_ (.B1(net595),
    .Y(_1314_),
    .A1(net660),
    .A2(_1313_));
 sg13g2_a21oi_1 _3701_ (.A1(_1476_),
    .A2(net660),
    .Y(_0211_),
    .B1(_1314_));
 sg13g2_xor2_1 _3702_ (.B(_1597_),
    .A(_1595_),
    .X(_1315_));
 sg13g2_o21ai_1 _3703_ (.B1(net594),
    .Y(_1316_),
    .A1(net907),
    .A2(net630));
 sg13g2_a21oi_1 _3704_ (.A1(net629),
    .A2(_1315_),
    .Y(_0212_),
    .B1(_1316_));
 sg13g2_xnor2_1 _3705_ (.Y(_1317_),
    .A(net917),
    .B(_1584_));
 sg13g2_xnor2_1 _3706_ (.Y(_1318_),
    .A(_1598_),
    .B(_1317_));
 sg13g2_o21ai_1 _3707_ (.B1(net594),
    .Y(_1319_),
    .A1(net917),
    .A2(net629));
 sg13g2_a21oi_1 _3708_ (.A1(net630),
    .A2(_1318_),
    .Y(_0213_),
    .B1(_1319_));
 sg13g2_xnor2_1 _3709_ (.Y(_1320_),
    .A(_1600_),
    .B(_1607_));
 sg13g2_o21ai_1 _3710_ (.B1(net595),
    .Y(_1321_),
    .A1(net660),
    .A2(_1320_));
 sg13g2_a21oi_1 _3711_ (.A1(_1475_),
    .A2(net660),
    .Y(_0214_),
    .B1(_1321_));
 sg13g2_a21oi_1 _3712_ (.A1(_1600_),
    .A2(_1606_),
    .Y(_1322_),
    .B1(_1604_));
 sg13g2_xnor2_1 _3713_ (.Y(_1323_),
    .A(_1582_),
    .B(_1322_));
 sg13g2_o21ai_1 _3714_ (.B1(net588),
    .Y(_1324_),
    .A1(net871),
    .A2(net629));
 sg13g2_a21oi_1 _3715_ (.A1(net629),
    .A2(_1323_),
    .Y(_0215_),
    .B1(_1324_));
 sg13g2_nor2_1 _3716_ (.A(_1616_),
    .B(_1622_),
    .Y(_1325_));
 sg13g2_nand2_1 _3717_ (.Y(_1326_),
    .A(_1608_),
    .B(_1618_));
 sg13g2_xnor2_1 _3718_ (.Y(_1327_),
    .A(_1325_),
    .B(_1326_));
 sg13g2_o21ai_1 _3719_ (.B1(net588),
    .Y(_1328_),
    .A1(net922),
    .A2(net629));
 sg13g2_a21oi_1 _3720_ (.A1(net629),
    .A2(_1327_),
    .Y(_0216_),
    .B1(_1328_));
 sg13g2_nor2_1 _3721_ (.A(_1612_),
    .B(_1619_),
    .Y(_1329_));
 sg13g2_a21o_1 _3722_ (.A2(_1326_),
    .A1(_1325_),
    .B1(_1616_),
    .X(_1330_));
 sg13g2_xnor2_1 _3723_ (.Y(_1331_),
    .A(_1329_),
    .B(_1330_));
 sg13g2_o21ai_1 _3724_ (.B1(net588),
    .Y(_1332_),
    .A1(net956),
    .A2(net629));
 sg13g2_a21oi_1 _3725_ (.A1(net629),
    .A2(_1331_),
    .Y(_0217_),
    .B1(_1332_));
 sg13g2_xnor2_1 _3726_ (.Y(_1333_),
    .A(_1623_),
    .B(_1626_));
 sg13g2_o21ai_1 _3727_ (.B1(net589),
    .Y(_1334_),
    .A1(net659),
    .A2(_1333_));
 sg13g2_a21oi_1 _3728_ (.A1(_1472_),
    .A2(net660),
    .Y(_0218_),
    .B1(_1334_));
 sg13g2_and2_1 _3729_ (.A(_1629_),
    .B(net589),
    .X(_0219_));
 sg13g2_nor2_1 _3730_ (.A(_1639_),
    .B(net565),
    .Y(_0220_));
 sg13g2_and2_1 _3731_ (.A(_1644_),
    .B(net589),
    .X(_0221_));
 sg13g2_and2_1 _3732_ (.A(_1653_),
    .B(net587),
    .X(_0222_));
 sg13g2_and2_1 _3733_ (.A(_1657_),
    .B(net586),
    .X(_0223_));
 sg13g2_nor2_1 _3734_ (.A(_0402_),
    .B(net566),
    .Y(_0224_));
 sg13g2_nor2_1 _3735_ (.A(_0407_),
    .B(net565),
    .Y(_0225_));
 sg13g2_nor2_1 _3736_ (.A(_0417_),
    .B(net566),
    .Y(_0226_));
 sg13g2_and2_1 _3737_ (.A(net414),
    .B(net576),
    .X(_0227_));
 sg13g2_and2_1 _3738_ (.A(net516),
    .B(net593),
    .X(_0228_));
 sg13g2_and2_1 _3739_ (.A(net436),
    .B(net593),
    .X(_0229_));
 sg13g2_and2_1 _3740_ (.A(net511),
    .B(net583),
    .X(_0230_));
 sg13g2_and2_1 _3741_ (.A(net518),
    .B(net593),
    .X(_0231_));
 sg13g2_and2_1 _3742_ (.A(net422),
    .B(net593),
    .X(_0232_));
 sg13g2_and2_1 _3743_ (.A(net416),
    .B(net583),
    .X(_0233_));
 sg13g2_and2_1 _3744_ (.A(net419),
    .B(net584),
    .X(_0234_));
 sg13g2_and2_1 _3745_ (.A(net438),
    .B(net584),
    .X(_0235_));
 sg13g2_and2_1 _3746_ (.A(net498),
    .B(net584),
    .X(_0236_));
 sg13g2_and2_1 _3747_ (.A(net456),
    .B(net585),
    .X(_0237_));
 sg13g2_and2_1 _3748_ (.A(net467),
    .B(net586),
    .X(_0238_));
 sg13g2_and2_1 _3749_ (.A(net488),
    .B(net586),
    .X(_0239_));
 sg13g2_and2_1 _3750_ (.A(net490),
    .B(net586),
    .X(_0240_));
 sg13g2_and2_1 _3751_ (.A(net469),
    .B(net585),
    .X(_0241_));
 sg13g2_and2_1 _3752_ (.A(net492),
    .B(net582),
    .X(_0242_));
 sg13g2_and2_1 _3753_ (.A(net479),
    .B(net586),
    .X(_0243_));
 sg13g2_nor2_1 _3754_ (.A(net657),
    .B(_0423_),
    .Y(_1335_));
 sg13g2_xnor2_1 _3755_ (.Y(_1336_),
    .A(net889),
    .B(_1335_));
 sg13g2_nor2_1 _3756_ (.A(net564),
    .B(_1336_),
    .Y(_0244_));
 sg13g2_xnor2_1 _3757_ (.Y(_1337_),
    .A(_0473_),
    .B(_0475_));
 sg13g2_o21ai_1 _3758_ (.B1(net593),
    .Y(_1338_),
    .A1(net657),
    .A2(_1337_));
 sg13g2_a21oi_1 _3759_ (.A1(_1488_),
    .A2(net657),
    .Y(_0245_),
    .B1(_1338_));
 sg13g2_xor2_1 _3760_ (.B(_0478_),
    .A(_0476_),
    .X(_1339_));
 sg13g2_o21ai_1 _3761_ (.B1(net593),
    .Y(_1340_),
    .A1(net900),
    .A2(net628));
 sg13g2_a21oi_1 _3762_ (.A1(net628),
    .A2(_1339_),
    .Y(_0246_),
    .B1(_1340_));
 sg13g2_xnor2_1 _3763_ (.Y(_1341_),
    .A(net936),
    .B(_0465_));
 sg13g2_xnor2_1 _3764_ (.Y(_1342_),
    .A(_0479_),
    .B(_1341_));
 sg13g2_o21ai_1 _3765_ (.B1(net583),
    .Y(_1343_),
    .A1(net936),
    .A2(net628));
 sg13g2_a21oi_1 _3766_ (.A1(net628),
    .A2(_1342_),
    .Y(_0247_),
    .B1(_1343_));
 sg13g2_o21ai_1 _3767_ (.B1(_0486_),
    .Y(_1344_),
    .A1(_0466_),
    .A2(_0480_));
 sg13g2_nor2b_1 _3768_ (.A(_0487_),
    .B_N(_1344_),
    .Y(_1345_));
 sg13g2_o21ai_1 _3769_ (.B1(net593),
    .Y(_1346_),
    .A1(net657),
    .A2(_1345_));
 sg13g2_a21oi_1 _3770_ (.A1(_1487_),
    .A2(net657),
    .Y(_0248_),
    .B1(_1346_));
 sg13g2_nor3_1 _3771_ (.A(_0463_),
    .B(_0484_),
    .C(_0487_),
    .Y(_1347_));
 sg13g2_o21ai_1 _3772_ (.B1(_0463_),
    .Y(_1348_),
    .A1(_0484_),
    .A2(_0487_));
 sg13g2_nor2_1 _3773_ (.A(net657),
    .B(_1347_),
    .Y(_1349_));
 sg13g2_a221oi_1 _3774_ (.B2(_1349_),
    .C1(net566),
    .B1(_1348_),
    .A1(_1486_),
    .Y(_0249_),
    .A2(net657));
 sg13g2_xnor2_1 _3775_ (.Y(_1350_),
    .A(_1485_),
    .B(_0495_));
 sg13g2_o21ai_1 _3776_ (.B1(_1350_),
    .Y(_1351_),
    .A1(_0488_),
    .A2(_0500_));
 sg13g2_or3_1 _3777_ (.A(_0488_),
    .B(_0500_),
    .C(_1350_),
    .X(_1352_));
 sg13g2_and2_1 _3778_ (.A(_1351_),
    .B(_1352_),
    .X(_1353_));
 sg13g2_o21ai_1 _3779_ (.B1(net584),
    .Y(_1354_),
    .A1(net658),
    .A2(_1353_));
 sg13g2_a21oi_1 _3780_ (.A1(_1485_),
    .A2(net657),
    .Y(_0250_),
    .B1(_1354_));
 sg13g2_nand2_1 _3781_ (.Y(_1355_),
    .A(_0492_),
    .B(_0498_));
 sg13g2_nor2b_1 _3782_ (.A(_0496_),
    .B_N(_1351_),
    .Y(_1356_));
 sg13g2_xnor2_1 _3783_ (.Y(_1357_),
    .A(_1355_),
    .B(_1356_));
 sg13g2_o21ai_1 _3784_ (.B1(net584),
    .Y(_1358_),
    .A1(net872),
    .A2(net628));
 sg13g2_a21oi_1 _3785_ (.A1(net627),
    .A2(_1357_),
    .Y(_0251_),
    .B1(_1358_));
 sg13g2_xnor2_1 _3786_ (.Y(_1359_),
    .A(_0503_),
    .B(_0505_));
 sg13g2_o21ai_1 _3787_ (.B1(net583),
    .Y(_1360_),
    .A1(net913),
    .A2(net627));
 sg13g2_a21oi_1 _3788_ (.A1(net627),
    .A2(_1359_),
    .Y(_0252_),
    .B1(_1360_));
 sg13g2_and2_1 _3789_ (.A(_0508_),
    .B(net584),
    .X(_0253_));
 sg13g2_and2_1 _3790_ (.A(_0516_),
    .B(net585),
    .X(_0254_));
 sg13g2_and2_1 _3791_ (.A(_0521_),
    .B(net586),
    .X(_0255_));
 sg13g2_and2_1 _3792_ (.A(_0531_),
    .B(net586),
    .X(_0256_));
 sg13g2_and2_1 _3793_ (.A(_0535_),
    .B(net586),
    .X(_0257_));
 sg13g2_nor2_1 _3794_ (.A(_0546_),
    .B(net565),
    .Y(_0258_));
 sg13g2_nor2_1 _3795_ (.A(_0551_),
    .B(net565),
    .Y(_0259_));
 sg13g2_nor2_1 _3796_ (.A(_0561_),
    .B(net566),
    .Y(_0260_));
 sg13g2_and2_1 _3797_ (.A(net428),
    .B(net592),
    .X(_0261_));
 sg13g2_and2_1 _3798_ (.A(net458),
    .B(net593),
    .X(_0262_));
 sg13g2_and2_1 _3799_ (.A(net463),
    .B(net594),
    .X(_0263_));
 sg13g2_and2_1 _3800_ (.A(net464),
    .B(net591),
    .X(_0264_));
 sg13g2_and2_1 _3801_ (.A(net475),
    .B(net591),
    .X(_0265_));
 sg13g2_and2_1 _3802_ (.A(net417),
    .B(net579),
    .X(_0266_));
 sg13g2_and2_1 _3803_ (.A(net468),
    .B(net591),
    .X(_0267_));
 sg13g2_and2_1 _3804_ (.A(net434),
    .B(net578),
    .X(_0268_));
 sg13g2_and2_1 _3805_ (.A(net432),
    .B(net583),
    .X(_0269_));
 sg13g2_and2_1 _3806_ (.A(net509),
    .B(net583),
    .X(_0270_));
 sg13g2_and2_1 _3807_ (.A(net418),
    .B(net570),
    .X(_0271_));
 sg13g2_and2_1 _3808_ (.A(net493),
    .B(net582),
    .X(_0272_));
 sg13g2_and2_1 _3809_ (.A(net448),
    .B(net570),
    .X(_0273_));
 sg13g2_and2_1 _3810_ (.A(net496),
    .B(net582),
    .X(_0274_));
 sg13g2_and2_1 _3811_ (.A(net454),
    .B(net582),
    .X(_0275_));
 sg13g2_and2_1 _3812_ (.A(net499),
    .B(net582),
    .X(_0276_));
 sg13g2_and2_1 _3813_ (.A(net474),
    .B(net582),
    .X(_0277_));
 sg13g2_and2_1 _3814_ (.A(net625),
    .B(_0603_),
    .X(_1361_));
 sg13g2_xnor2_1 _3815_ (.Y(_1362_),
    .A(net865),
    .B(_1361_));
 sg13g2_nor2_1 _3816_ (.A(net566),
    .B(_1362_),
    .Y(_0278_));
 sg13g2_xnor2_1 _3817_ (.Y(_1363_),
    .A(_0609_),
    .B(_0611_));
 sg13g2_o21ai_1 _3818_ (.B1(net592),
    .Y(_1364_),
    .A1(net655),
    .A2(_1363_));
 sg13g2_a21oi_1 _3819_ (.A1(_1497_),
    .A2(net655),
    .Y(_0279_),
    .B1(_1364_));
 sg13g2_xor2_1 _3820_ (.B(_0613_),
    .A(_0612_),
    .X(_1365_));
 sg13g2_o21ai_1 _3821_ (.B1(net591),
    .Y(_1366_),
    .A1(net655),
    .A2(_1365_));
 sg13g2_a21oi_1 _3822_ (.A1(_1496_),
    .A2(net655),
    .Y(_0280_),
    .B1(_1366_));
 sg13g2_xnor2_1 _3823_ (.Y(_1367_),
    .A(_0614_),
    .B(_0615_));
 sg13g2_o21ai_1 _3824_ (.B1(net592),
    .Y(_1368_),
    .A1(net916),
    .A2(_1498_));
 sg13g2_a21oi_1 _3825_ (.A1(net625),
    .A2(_1367_),
    .Y(_0281_),
    .B1(_1368_));
 sg13g2_xnor2_1 _3826_ (.Y(_1369_),
    .A(_0616_),
    .B(_0621_));
 sg13g2_o21ai_1 _3827_ (.B1(net591),
    .Y(_1370_),
    .A1(net957),
    .A2(net625));
 sg13g2_a21oi_1 _3828_ (.A1(net625),
    .A2(_1369_),
    .Y(_0282_),
    .B1(_1370_));
 sg13g2_a21oi_1 _3829_ (.A1(_0616_),
    .A2(_0621_),
    .Y(_1371_),
    .B1(_0619_));
 sg13g2_xor2_1 _3830_ (.B(_1371_),
    .A(_0623_),
    .X(_1372_));
 sg13g2_o21ai_1 _3831_ (.B1(net591),
    .Y(_1373_),
    .A1(net932),
    .A2(net625));
 sg13g2_a21oi_1 _3832_ (.A1(net625),
    .A2(_1372_),
    .Y(_0283_),
    .B1(_1373_));
 sg13g2_and2_1 _3833_ (.A(_0589_),
    .B(_0592_),
    .X(_1374_));
 sg13g2_xnor2_1 _3834_ (.Y(_1375_),
    .A(_0626_),
    .B(_1374_));
 sg13g2_o21ai_1 _3835_ (.B1(net591),
    .Y(_1376_),
    .A1(net655),
    .A2(_1375_));
 sg13g2_a21oi_1 _3836_ (.A1(_1495_),
    .A2(net655),
    .Y(_0284_),
    .B1(_1376_));
 sg13g2_nand2_1 _3837_ (.Y(_1377_),
    .A(_0585_),
    .B(_0586_));
 sg13g2_o21ai_1 _3838_ (.B1(_0592_),
    .Y(_1378_),
    .A1(_0590_),
    .A2(_0626_));
 sg13g2_or2_1 _3839_ (.X(_1379_),
    .B(_1378_),
    .A(_1377_));
 sg13g2_a21oi_1 _3840_ (.A1(_1377_),
    .A2(_1378_),
    .Y(_1380_),
    .B1(net655));
 sg13g2_o21ai_1 _3841_ (.B1(net591),
    .Y(_1381_),
    .A1(net933),
    .A2(net625));
 sg13g2_a21oi_1 _3842_ (.A1(_1379_),
    .A2(_1380_),
    .Y(_0285_),
    .B1(_1381_));
 sg13g2_xnor2_1 _3843_ (.Y(_1382_),
    .A(_0628_),
    .B(_0631_));
 sg13g2_o21ai_1 _3844_ (.B1(net583),
    .Y(_1383_),
    .A1(net911),
    .A2(net626));
 sg13g2_a21oi_1 _3845_ (.A1(net626),
    .A2(_1382_),
    .Y(_0286_),
    .B1(_1383_));
 sg13g2_and2_1 _3846_ (.A(_0636_),
    .B(net583),
    .X(_0287_));
 sg13g2_nor2_1 _3847_ (.A(_0645_),
    .B(net565),
    .Y(_0288_));
 sg13g2_nor2_1 _3848_ (.A(_0652_),
    .B(net565),
    .Y(_0289_));
 sg13g2_and2_1 _3849_ (.A(_0662_),
    .B(net570),
    .X(_0290_));
 sg13g2_nor2_1 _3850_ (.A(_0668_),
    .B(net565),
    .Y(_0291_));
 sg13g2_and2_1 _3851_ (.A(_0677_),
    .B(net582),
    .X(_0292_));
 sg13g2_and2_1 _3852_ (.A(_0682_),
    .B(net582),
    .X(_0293_));
 sg13g2_nor2_1 _3853_ (.A(_0690_),
    .B(net565),
    .Y(_0294_));
 sg13g2_and2_1 _3854_ (.A(net457),
    .B(net574),
    .X(_0295_));
 sg13g2_and2_1 _3855_ (.A(net485),
    .B(net578),
    .X(_0296_));
 sg13g2_and2_1 _3856_ (.A(net413),
    .B(net578),
    .X(_0297_));
 sg13g2_and2_1 _3857_ (.A(net426),
    .B(net578),
    .X(_0298_));
 sg13g2_and2_1 _3858_ (.A(net445),
    .B(net575),
    .X(_0299_));
 sg13g2_and2_1 _3859_ (.A(net430),
    .B(net575),
    .X(_0300_));
 sg13g2_and2_1 _3860_ (.A(net431),
    .B(net574),
    .X(_0301_));
 sg13g2_and2_1 _3861_ (.A(net480),
    .B(net575),
    .X(_0302_));
 sg13g2_and2_1 _3862_ (.A(net519),
    .B(net573),
    .X(_0303_));
 sg13g2_and2_1 _3863_ (.A(net446),
    .B(net568),
    .X(_0304_));
 sg13g2_and2_1 _3864_ (.A(net451),
    .B(net568),
    .X(_0305_));
 sg13g2_and2_1 _3865_ (.A(net453),
    .B(net568),
    .X(_0306_));
 sg13g2_and2_1 _3866_ (.A(net486),
    .B(net571),
    .X(_0307_));
 sg13g2_and2_1 _3867_ (.A(net466),
    .B(net571),
    .X(_0308_));
 sg13g2_and2_1 _3868_ (.A(net443),
    .B(net570),
    .X(_0309_));
 sg13g2_and2_1 _3869_ (.A(net435),
    .B(net571),
    .X(_0310_));
 sg13g2_and2_1 _3870_ (.A(net491),
    .B(net570),
    .X(_0311_));
 sg13g2_nor2_1 _3871_ (.A(net652),
    .B(_0696_),
    .Y(_1384_));
 sg13g2_xnor2_1 _3872_ (.Y(_1385_),
    .A(net915),
    .B(_1384_));
 sg13g2_nor2_1 _3873_ (.A(net564),
    .B(_1385_),
    .Y(_0312_));
 sg13g2_xnor2_1 _3874_ (.Y(_1386_),
    .A(_0733_),
    .B(_0734_));
 sg13g2_o21ai_1 _3875_ (.B1(net578),
    .Y(_1387_),
    .A1(net914),
    .A2(net622));
 sg13g2_a21oi_1 _3876_ (.A1(net622),
    .A2(_1386_),
    .Y(_0313_),
    .B1(_1387_));
 sg13g2_xnor2_1 _3877_ (.Y(_1388_),
    .A(_0736_),
    .B(_0745_));
 sg13g2_o21ai_1 _3878_ (.B1(net578),
    .Y(_1389_),
    .A1(net926),
    .A2(net623));
 sg13g2_a21oi_1 _3879_ (.A1(net623),
    .A2(_1388_),
    .Y(_0314_),
    .B1(_1389_));
 sg13g2_a21oi_1 _3880_ (.A1(_0736_),
    .A2(_0745_),
    .Y(_1390_),
    .B1(_0744_));
 sg13g2_xnor2_1 _3881_ (.Y(_1391_),
    .A(_0742_),
    .B(_1390_));
 sg13g2_o21ai_1 _3882_ (.B1(net578),
    .Y(_1392_),
    .A1(net873),
    .A2(net622));
 sg13g2_a21oi_1 _3883_ (.A1(net622),
    .A2(_1391_),
    .Y(_0315_),
    .B1(_1392_));
 sg13g2_nand2_1 _3884_ (.Y(_1393_),
    .A(_0748_),
    .B(_0756_));
 sg13g2_xnor2_1 _3885_ (.Y(_1394_),
    .A(_0748_),
    .B(_0756_));
 sg13g2_o21ai_1 _3886_ (.B1(net575),
    .Y(_1395_),
    .A1(net937),
    .A2(net622));
 sg13g2_a21oi_1 _3887_ (.A1(net622),
    .A2(_1394_),
    .Y(_0316_),
    .B1(_1395_));
 sg13g2_nand2_1 _3888_ (.Y(_1396_),
    .A(_0755_),
    .B(_1393_));
 sg13g2_xnor2_1 _3889_ (.Y(_1397_),
    .A(_0752_),
    .B(_1396_));
 sg13g2_o21ai_1 _3890_ (.B1(net575),
    .Y(_1398_),
    .A1(net961),
    .A2(net622));
 sg13g2_a21oi_1 _3891_ (.A1(net622),
    .A2(_1397_),
    .Y(_0317_),
    .B1(_1398_));
 sg13g2_nand2b_1 _3892_ (.Y(_1399_),
    .B(_0768_),
    .A_N(_0765_));
 sg13g2_nor2_1 _3893_ (.A(_0759_),
    .B(_1399_),
    .Y(_1400_));
 sg13g2_xor2_1 _3894_ (.B(_1399_),
    .A(_0759_),
    .X(_1401_));
 sg13g2_o21ai_1 _3895_ (.B1(net575),
    .Y(_1402_),
    .A1(net652),
    .A2(_1401_));
 sg13g2_a21oi_1 _3896_ (.A1(_1504_),
    .A2(net652),
    .Y(_0318_),
    .B1(_1402_));
 sg13g2_xnor2_1 _3897_ (.Y(_1403_),
    .A(_1503_),
    .B(_0761_));
 sg13g2_o21ai_1 _3898_ (.B1(_1403_),
    .Y(_1404_),
    .A1(_0765_),
    .A2(_1400_));
 sg13g2_nor3_1 _3899_ (.A(_0765_),
    .B(_1400_),
    .C(_1403_),
    .Y(_1405_));
 sg13g2_nor2_1 _3900_ (.A(net652),
    .B(_1405_),
    .Y(_1406_));
 sg13g2_a221oi_1 _3901_ (.B2(_1406_),
    .C1(net564),
    .B1(_1404_),
    .A1(_1503_),
    .Y(_0319_),
    .A2(net652));
 sg13g2_xnor2_1 _3902_ (.Y(_1407_),
    .A(_0770_),
    .B(_0772_));
 sg13g2_o21ai_1 _3903_ (.B1(net576),
    .Y(_1408_),
    .A1(net888),
    .A2(net624));
 sg13g2_a21oi_1 _3904_ (.A1(net624),
    .A2(_1407_),
    .Y(_0320_),
    .B1(_1408_));
 sg13g2_and2_1 _3905_ (.A(_0775_),
    .B(net567),
    .X(_0321_));
 sg13g2_nor2_1 _3906_ (.A(_0784_),
    .B(net564),
    .Y(_0322_));
 sg13g2_and2_1 _3907_ (.A(_0789_),
    .B(net568),
    .X(_0323_));
 sg13g2_nor2_1 _3908_ (.A(_0799_),
    .B(net563),
    .Y(_0324_));
 sg13g2_and2_1 _3909_ (.A(_0804_),
    .B(net571),
    .X(_0325_));
 sg13g2_nor2_1 _3910_ (.A(_0814_),
    .B(net563),
    .Y(_0326_));
 sg13g2_nor2_1 _3911_ (.A(_0820_),
    .B(net563),
    .Y(_0327_));
 sg13g2_nor2_1 _3912_ (.A(_0829_),
    .B(net563),
    .Y(_0328_));
 sg13g2_and2_1 _3913_ (.A(net412),
    .B(net572),
    .X(_0329_));
 sg13g2_and2_1 _3914_ (.A(net465),
    .B(net574),
    .X(_0330_));
 sg13g2_and2_1 _3915_ (.A(net421),
    .B(net574),
    .X(_0331_));
 sg13g2_and2_1 _3916_ (.A(net425),
    .B(net574),
    .X(_0332_));
 sg13g2_and2_1 _3917_ (.A(net462),
    .B(net573),
    .X(_0333_));
 sg13g2_and2_1 _3918_ (.A(net409),
    .B(net573),
    .X(_0334_));
 sg13g2_and2_1 _3919_ (.A(net460),
    .B(net572),
    .X(_0335_));
 sg13g2_and2_1 _3920_ (.A(net476),
    .B(net572),
    .X(_0336_));
 sg13g2_and2_1 _3921_ (.A(net411),
    .B(net572),
    .X(_0337_));
 sg13g2_and2_1 _3922_ (.A(net410),
    .B(net567),
    .X(_0338_));
 sg13g2_and2_1 _3923_ (.A(net487),
    .B(net567),
    .X(_0339_));
 sg13g2_and2_1 _3924_ (.A(net503),
    .B(net567),
    .X(_0340_));
 sg13g2_and2_1 _3925_ (.A(net470),
    .B(net569),
    .X(_0341_));
 sg13g2_and2_1 _3926_ (.A(net507),
    .B(net567),
    .X(_0342_));
 sg13g2_and2_1 _3927_ (.A(net502),
    .B(net569),
    .X(_0343_));
 sg13g2_and2_1 _3928_ (.A(net489),
    .B(net569),
    .X(_0344_));
 sg13g2_and2_1 _3929_ (.A(net424),
    .B(net570),
    .X(_0345_));
 sg13g2_nor2_1 _3930_ (.A(\systolic_array.genblk2[0].mac[4].zero ),
    .B(_0835_),
    .Y(_1409_));
 sg13g2_xnor2_1 _3931_ (.Y(_1410_),
    .A(net851),
    .B(_1409_));
 sg13g2_nor2_1 _3932_ (.A(net564),
    .B(net852),
    .Y(_0346_));
 sg13g2_xnor2_1 _3933_ (.Y(_1411_),
    .A(_0887_),
    .B(_0888_));
 sg13g2_o21ai_1 _3934_ (.B1(net574),
    .Y(_1412_),
    .A1(net938),
    .A2(net619));
 sg13g2_a21oi_1 _3935_ (.A1(net620),
    .A2(_1411_),
    .Y(_0347_),
    .B1(_1412_));
 sg13g2_xnor2_1 _3936_ (.Y(_1413_),
    .A(_0890_),
    .B(_0899_));
 sg13g2_o21ai_1 _3937_ (.B1(net574),
    .Y(_1414_),
    .A1(net925),
    .A2(net620));
 sg13g2_a21oi_1 _3938_ (.A1(net620),
    .A2(_1413_),
    .Y(_0348_),
    .B1(_1414_));
 sg13g2_a21oi_1 _3939_ (.A1(_0890_),
    .A2(_0899_),
    .Y(_1415_),
    .B1(_0898_));
 sg13g2_xnor2_1 _3940_ (.Y(_1416_),
    .A(_0896_),
    .B(_1415_));
 sg13g2_o21ai_1 _3941_ (.B1(net574),
    .Y(_1417_),
    .A1(net883),
    .A2(net619));
 sg13g2_a21oi_1 _3942_ (.A1(net619),
    .A2(_1416_),
    .Y(_0349_),
    .B1(_1417_));
 sg13g2_xnor2_1 _3943_ (.Y(_1418_),
    .A(_0902_),
    .B(_0911_));
 sg13g2_o21ai_1 _3944_ (.B1(net573),
    .Y(_1419_),
    .A1(net868),
    .A2(net620));
 sg13g2_a21oi_1 _3945_ (.A1(net620),
    .A2(_1418_),
    .Y(_0350_),
    .B1(_1419_));
 sg13g2_a21oi_1 _3946_ (.A1(_0902_),
    .A2(_0911_),
    .Y(_1420_),
    .B1(_0909_));
 sg13g2_xnor2_1 _3947_ (.Y(_1421_),
    .A(_0906_),
    .B(_1420_));
 sg13g2_nor2_1 _3948_ (.A(net650),
    .B(_1421_),
    .Y(_1422_));
 sg13g2_o21ai_1 _3949_ (.B1(net572),
    .Y(_1423_),
    .A1(net971),
    .A2(net619));
 sg13g2_nor2_1 _3950_ (.A(_1422_),
    .B(_1423_),
    .Y(_0351_));
 sg13g2_xnor2_1 _3951_ (.Y(_1424_),
    .A(net941),
    .B(_0877_));
 sg13g2_xnor2_1 _3952_ (.Y(_1425_),
    .A(_0915_),
    .B(_1424_));
 sg13g2_o21ai_1 _3953_ (.B1(net572),
    .Y(_1426_),
    .A1(net941),
    .A2(net619));
 sg13g2_a21oi_1 _3954_ (.A1(net619),
    .A2(_1425_),
    .Y(_0352_),
    .B1(_1426_));
 sg13g2_xor2_1 _3955_ (.B(_0873_),
    .A(net943),
    .X(_1427_));
 sg13g2_a21oi_1 _3956_ (.A1(_0878_),
    .A2(_0915_),
    .Y(_1428_),
    .B1(_0916_));
 sg13g2_xnor2_1 _3957_ (.Y(_1429_),
    .A(_1427_),
    .B(_1428_));
 sg13g2_o21ai_1 _3958_ (.B1(net572),
    .Y(_1430_),
    .A1(net943),
    .A2(net619));
 sg13g2_a21oi_1 _3959_ (.A1(net619),
    .A2(_1429_),
    .Y(_0353_),
    .B1(_1430_));
 sg13g2_xnor2_1 _3960_ (.Y(_1431_),
    .A(_0919_),
    .B(_0920_));
 sg13g2_o21ai_1 _3961_ (.B1(net572),
    .Y(_1432_),
    .A1(net935),
    .A2(net621));
 sg13g2_a21oi_1 _3962_ (.A1(net621),
    .A2(_1431_),
    .Y(_0354_),
    .B1(_1432_));
 sg13g2_and2_1 _3963_ (.A(_0923_),
    .B(net567),
    .X(_0355_));
 sg13g2_nor2_1 _3964_ (.A(_0932_),
    .B(net564),
    .Y(_0356_));
 sg13g2_and2_1 _3965_ (.A(_0938_),
    .B(net567),
    .X(_0357_));
 sg13g2_nor2_1 _3966_ (.A(_0948_),
    .B(net562),
    .Y(_0358_));
 sg13g2_and2_1 _3967_ (.A(_0953_),
    .B(net567),
    .X(_0359_));
 sg13g2_nor2_1 _3968_ (.A(_0963_),
    .B(net562),
    .Y(_0360_));
 sg13g2_nor2_1 _3969_ (.A(_0968_),
    .B(net562),
    .Y(_0361_));
 sg13g2_nor2_1 _3970_ (.A(_0977_),
    .B(net563),
    .Y(_0362_));
 sg13g2_mux2_1 _3971_ (.A0(net798),
    .A1(\systolic_array.genblk2[0].mac[0].div2 ),
    .S(net639),
    .X(_0363_));
 sg13g2_mux2_1 _3972_ (.A0(net504),
    .A1(net635),
    .S(net639),
    .X(_0364_));
 sg13g2_nor2_1 _3973_ (.A(net638),
    .B(net920),
    .Y(_1433_));
 sg13g2_a21oi_1 _3974_ (.A1(net638),
    .A2(_1501_),
    .Y(_0365_),
    .B1(_1433_));
 sg13g2_mux2_1 _3975_ (.A0(net800),
    .A1(net906),
    .S(net639),
    .X(_0366_));
 sg13g2_and2_1 _3976_ (.A(net617),
    .B(_1015_),
    .X(_1434_));
 sg13g2_xnor2_1 _3977_ (.Y(_1435_),
    .A(net840),
    .B(_1434_));
 sg13g2_nor2_1 _3978_ (.A(net564),
    .B(_1435_),
    .Y(_0367_));
 sg13g2_xnor2_1 _3979_ (.Y(_1436_),
    .A(_1021_),
    .B(_1023_));
 sg13g2_o21ai_1 _3980_ (.B1(net578),
    .Y(_1437_),
    .A1(net649),
    .A2(_1436_));
 sg13g2_a21oi_1 _3981_ (.A1(_1520_),
    .A2(net649),
    .Y(_0368_),
    .B1(_1437_));
 sg13g2_xnor2_1 _3982_ (.Y(_1438_),
    .A(_1024_),
    .B(_1025_));
 sg13g2_o21ai_1 _3983_ (.B1(net577),
    .Y(_1439_),
    .A1(net949),
    .A2(net617));
 sg13g2_a21oi_1 _3984_ (.A1(net617),
    .A2(_1438_),
    .Y(_0369_),
    .B1(_1439_));
 sg13g2_xnor2_1 _3985_ (.Y(_1440_),
    .A(_1026_),
    .B(_1027_));
 sg13g2_o21ai_1 _3986_ (.B1(net576),
    .Y(_1441_),
    .A1(net927),
    .A2(net617));
 sg13g2_a21oi_1 _3987_ (.A1(net616),
    .A2(_1440_),
    .Y(_0370_),
    .B1(_1441_));
 sg13g2_xnor2_1 _3988_ (.Y(_1442_),
    .A(_1028_),
    .B(_1032_));
 sg13g2_o21ai_1 _3989_ (.B1(net576),
    .Y(_1443_),
    .A1(net940),
    .A2(net617));
 sg13g2_a21oi_1 _3990_ (.A1(net616),
    .A2(_1442_),
    .Y(_0371_),
    .B1(_1443_));
 sg13g2_o21ai_1 _3991_ (.B1(_1031_),
    .Y(_1444_),
    .A1(_1028_),
    .A2(_1032_));
 sg13g2_nor2_1 _3992_ (.A(_1008_),
    .B(_1444_),
    .Y(_1445_));
 sg13g2_nand2_1 _3993_ (.Y(_1446_),
    .A(_1008_),
    .B(_1444_));
 sg13g2_nor2_1 _3994_ (.A(net649),
    .B(_1445_),
    .Y(_1447_));
 sg13g2_o21ai_1 _3995_ (.B1(net577),
    .Y(_1448_),
    .A1(net898),
    .A2(net616));
 sg13g2_a21oi_1 _3996_ (.A1(_1446_),
    .A2(_1447_),
    .Y(_0372_),
    .B1(_1448_));
 sg13g2_xnor2_1 _3997_ (.Y(_1449_),
    .A(\systolic_array.genblk1[10].accumulators_dlygate[6].A ),
    .B(_1039_));
 sg13g2_nor2_1 _3998_ (.A(_1033_),
    .B(_1043_),
    .Y(_1450_));
 sg13g2_o21ai_1 _3999_ (.B1(_1449_),
    .Y(_1451_),
    .A1(_1033_),
    .A2(_1043_));
 sg13g2_xor2_1 _4000_ (.B(_1450_),
    .A(_1449_),
    .X(_1452_));
 sg13g2_o21ai_1 _4001_ (.B1(net576),
    .Y(_1453_),
    .A1(net942),
    .A2(net616));
 sg13g2_a21oi_1 _4002_ (.A1(net616),
    .A2(_1452_),
    .Y(_0373_),
    .B1(_1453_));
 sg13g2_nor2_1 _4003_ (.A(_1037_),
    .B(_1041_),
    .Y(_1454_));
 sg13g2_o21ai_1 _4004_ (.B1(_1451_),
    .Y(_1455_),
    .A1(_1519_),
    .A2(_1039_));
 sg13g2_xnor2_1 _4005_ (.Y(_1456_),
    .A(_1454_),
    .B(_1455_));
 sg13g2_o21ai_1 _4006_ (.B1(net577),
    .Y(_1457_),
    .A1(net947),
    .A2(net616));
 sg13g2_a21oi_1 _4007_ (.A1(net616),
    .A2(_1456_),
    .Y(_0374_),
    .B1(_1457_));
 sg13g2_xnor2_1 _4008_ (.Y(_1458_),
    .A(_1047_),
    .B(_1049_));
 sg13g2_o21ai_1 _4009_ (.B1(net570),
    .Y(_1459_),
    .A1(net894),
    .A2(net618));
 sg13g2_a21oi_1 _4010_ (.A1(net618),
    .A2(_1458_),
    .Y(_0375_),
    .B1(_1459_));
 sg13g2_nor2_1 _4011_ (.A(_1055_),
    .B(net562),
    .Y(_0376_));
 sg13g2_nor2_1 _4012_ (.A(_1065_),
    .B(net560),
    .Y(_0377_));
 sg13g2_nor2_1 _4013_ (.A(_1072_),
    .B(net560),
    .Y(_0378_));
 sg13g2_nor2_1 _4014_ (.A(_1083_),
    .B(net560),
    .Y(_0379_));
 sg13g2_nor2_1 _4015_ (.A(_1089_),
    .B(net560),
    .Y(_0380_));
 sg13g2_nor2_1 _4016_ (.A(_1100_),
    .B(net561),
    .Y(_0381_));
 sg13g2_nor2_1 _4017_ (.A(_1106_),
    .B(net561),
    .Y(_0382_));
 sg13g2_nor2_1 _4018_ (.A(_1114_),
    .B(net563),
    .Y(_0383_));
 sg13g2_and2_1 _4019_ (.A(net452),
    .B(net579),
    .X(_0384_));
 sg13g2_and2_1 _4020_ (.A(net423),
    .B(net579),
    .X(_0385_));
 sg13g2_and2_1 _4021_ (.A(net472),
    .B(net577),
    .X(_0386_));
 sg13g2_and2_1 _4022_ (.A(net506),
    .B(net576),
    .X(_0387_));
 sg13g2_and2_1 _4023_ (.A(net449),
    .B(net576),
    .X(_0388_));
 sg13g2_and2_1 _4024_ (.A(net441),
    .B(net577),
    .X(_0389_));
 sg13g2_and2_1 _4025_ (.A(net450),
    .B(net576),
    .X(_0390_));
 sg13g2_and2_1 _4026_ (.A(net420),
    .B(net577),
    .X(_0391_));
 sg13g2_and2_1 _4027_ (.A(net495),
    .B(net570),
    .X(_0392_));
 sg13g2_nor2_1 _4028_ (.A(_1523_),
    .B(net561),
    .Y(_0393_));
 sg13g2_nor2_1 _4029_ (.A(_1524_),
    .B(net560),
    .Y(_0394_));
 sg13g2_nor2_1 _4030_ (.A(_1525_),
    .B(net560),
    .Y(_0395_));
 sg13g2_nor2_1 _4031_ (.A(_1526_),
    .B(net560),
    .Y(_0396_));
 sg13g2_nor2_1 _4032_ (.A(_1527_),
    .B(net560),
    .Y(_0397_));
 sg13g2_nor2_1 _4033_ (.A(_1528_),
    .B(net561),
    .Y(_0398_));
 sg13g2_nor2_1 _4034_ (.A(_1529_),
    .B(net561),
    .Y(_0399_));
 sg13g2_nor2_1 _4035_ (.A(_1530_),
    .B(net563),
    .Y(_0400_));
 sg13g2_dfrbp_1 _4036_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net79),
    .D(_0120_),
    .Q_N(_1927_),
    .Q(\systolic_array.arg_left_sign_next[3] ));
 sg13g2_dfrbp_1 _4037_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net80),
    .D(_0000_),
    .Q_N(_0100_),
    .Q(\systolic_array.arg_top_curr[0] ));
 sg13g2_dfrbp_1 _4038_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net81),
    .D(_0001_),
    .Q_N(_0101_),
    .Q(\systolic_array.arg_top_curr[1] ));
 sg13g2_dfrbp_1 _4039_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net82),
    .D(_0002_),
    .Q_N(_0105_),
    .Q(\systolic_array.arg_top_curr[2] ));
 sg13g2_dfrbp_1 _4040_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net83),
    .D(_0003_),
    .Q_N(_1928_),
    .Q(\systolic_array.arg_top_curr[3] ));
 sg13g2_dfrbp_1 _4041_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net84),
    .D(_0004_),
    .Q_N(_1929_),
    .Q(\systolic_array.arg_top_curr[4] ));
 sg13g2_dfrbp_1 _4042_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net85),
    .D(_0005_),
    .Q_N(_0099_),
    .Q(\systolic_array.arg_top_curr[5] ));
 sg13g2_dfrbp_1 _4043_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net332),
    .D(_0006_),
    .Q_N(_0116_),
    .Q(\systolic_array.arg_top_curr[6] ));
 sg13g2_dfrbp_1 _4044_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net78),
    .D(_0007_),
    .Q_N(_0115_),
    .Q(\systolic_array.arg_top_curr[7] ));
 sg13g2_dfrbp_1 _4045_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net60),
    .D(net743),
    .Q_N(_1926_),
    .Q(\systolic_array.genblk1[11].out_queue_dlygate[9].A ));
 sg13g2_dfrbp_1 _4046_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net356),
    .D(_0122_),
    .Q_N(_1925_),
    .Q(\systolic_array.genblk1[11].out_queue_dlygate[10].A ));
 sg13g2_dfrbp_1 _4047_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net355),
    .D(_0123_),
    .Q_N(_1924_),
    .Q(\systolic_array.genblk1[11].out_queue_dlygate[11].A ));
 sg13g2_dfrbp_1 _4048_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net354),
    .D(_0124_),
    .Q_N(_1923_),
    .Q(\systolic_array.genblk1[11].out_queue_dlygate[12].A ));
 sg13g2_dfrbp_1 _4049_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net353),
    .D(net739),
    .Q_N(_1922_),
    .Q(\systolic_array.genblk1[11].out_queue_dlygate[13].A ));
 sg13g2_dfrbp_1 _4050_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net352),
    .D(_0126_),
    .Q_N(_1921_),
    .Q(\systolic_array.genblk1[11].out_queue_dlygate[14].A ));
 sg13g2_dfrbp_1 _4051_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net351),
    .D(_0127_),
    .Q_N(_1920_),
    .Q(\systolic_array.genblk1[11].out_queue_dlygate[15].A ));
 sg13g2_dfrbp_1 _4052_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net350),
    .D(_0128_),
    .Q_N(_1919_),
    .Q(\systolic_array.genblk1[11].out_queue_dlygate[16].A ));
 sg13g2_dfrbp_1 _4053_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net349),
    .D(_0129_),
    .Q_N(_1918_),
    .Q(\systolic_array.arg_top_next[0] ));
 sg13g2_dfrbp_1 _4054_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net348),
    .D(_0130_),
    .Q_N(_1917_),
    .Q(\systolic_array.arg_top_next[1] ));
 sg13g2_dfrbp_1 _4055_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net347),
    .D(_0131_),
    .Q_N(_1916_),
    .Q(\systolic_array.arg_top_next[2] ));
 sg13g2_dfrbp_1 _4056_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net346),
    .D(_0132_),
    .Q_N(_1915_),
    .Q(\systolic_array.arg_top_next[3] ));
 sg13g2_dfrbp_1 _4057_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net345),
    .D(_0133_),
    .Q_N(_1914_),
    .Q(\systolic_array.arg_top_next[4] ));
 sg13g2_dfrbp_1 _4058_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net344),
    .D(_0134_),
    .Q_N(_1913_),
    .Q(\systolic_array.arg_top_next[5] ));
 sg13g2_dfrbp_1 _4059_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net343),
    .D(_0135_),
    .Q_N(_1912_),
    .Q(\systolic_array.arg_top_next[6] ));
 sg13g2_dfrbp_1 _4060_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net342),
    .D(_0136_),
    .Q_N(_1911_),
    .Q(\systolic_array.arg_top_next[7] ));
 sg13g2_dfrbp_1 _4061_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net341),
    .D(_0137_),
    .Q_N(_1910_),
    .Q(\systolic_array.arg_top_next[8] ));
 sg13g2_dfrbp_1 _4062_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net340),
    .D(_0138_),
    .Q_N(_1909_),
    .Q(\systolic_array.arg_top_next[9] ));
 sg13g2_dfrbp_1 _4063_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net331),
    .D(_0139_),
    .Q_N(_1908_),
    .Q(\systolic_array.arg_top_next[10] ));
 sg13g2_dfrbp_1 _4064_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net330),
    .D(_0140_),
    .Q_N(_1907_),
    .Q(\systolic_array.arg_top_next[11] ));
 sg13g2_dfrbp_1 _4065_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net329),
    .D(_0141_),
    .Q_N(_1906_),
    .Q(\systolic_array.arg_top_next[12] ));
 sg13g2_dfrbp_1 _4066_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net328),
    .D(_0142_),
    .Q_N(_1905_),
    .Q(\systolic_array.arg_top_next[13] ));
 sg13g2_dfrbp_1 _4067_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net327),
    .D(_0143_),
    .Q_N(_1904_),
    .Q(\systolic_array.arg_top_next[14] ));
 sg13g2_dfrbp_1 _4068_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net326),
    .D(_0144_),
    .Q_N(_1903_),
    .Q(\systolic_array.arg_top_next[15] ));
 sg13g2_dfrbp_1 _4069_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net325),
    .D(_0145_),
    .Q_N(_1902_),
    .Q(\systolic_array.arg_left_sign_next[0] ));
 sg13g2_dfrbp_1 _4070_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net324),
    .D(_0146_),
    .Q_N(_1901_),
    .Q(\systolic_array.arg_left_sign_next[1] ));
 sg13g2_dfrbp_1 _4071_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net323),
    .D(_0147_),
    .Q_N(_1900_),
    .Q(\systolic_array.arg_left_sign_next[2] ));
 sg13g2_dfrbp_1 _4072_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net322),
    .D(_0148_),
    .Q_N(_1899_),
    .Q(\systolic_array.arg_left_zero_next[0] ));
 sg13g2_dfrbp_1 _4073_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net321),
    .D(_0149_),
    .Q_N(_1898_),
    .Q(\systolic_array.arg_left_zero_next[1] ));
 sg13g2_dfrbp_1 _4074_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net320),
    .D(_0150_),
    .Q_N(_1897_),
    .Q(\systolic_array.arg_left_zero_next[2] ));
 sg13g2_dfrbp_1 _4075_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net319),
    .D(_0151_),
    .Q_N(_1896_),
    .Q(\systolic_array.arg_top_curr[8] ));
 sg13g2_dfrbp_1 _4076_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net318),
    .D(_0152_),
    .Q_N(_1895_),
    .Q(\systolic_array.arg_top_curr[9] ));
 sg13g2_dfrbp_1 _4077_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net317),
    .D(_0153_),
    .Q_N(_1894_),
    .Q(\systolic_array.arg_top_curr[10] ));
 sg13g2_dfrbp_1 _4078_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net316),
    .D(net513),
    .Q_N(_1893_),
    .Q(\systolic_array.arg_top_curr[11] ));
 sg13g2_dfrbp_1 _4079_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net315),
    .D(_0155_),
    .Q_N(_1892_),
    .Q(\systolic_array.arg_top_curr[12] ));
 sg13g2_dfrbp_1 _4080_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net314),
    .D(_0156_),
    .Q_N(_1891_),
    .Q(\systolic_array.arg_top_curr[13] ));
 sg13g2_dfrbp_1 _4081_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net313),
    .D(_0157_),
    .Q_N(_1890_),
    .Q(\systolic_array.arg_top_curr[14] ));
 sg13g2_dfrbp_1 _4082_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net312),
    .D(_0158_),
    .Q_N(_1889_),
    .Q(\systolic_array.arg_top_curr[15] ));
 sg13g2_dfrbp_1 _4083_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net311),
    .D(_0159_),
    .Q_N(_1888_),
    .Q(\systolic_array.arg_left_div2_next[0] ));
 sg13g2_dfrbp_1 _4084_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net310),
    .D(_0160_),
    .Q_N(_1887_),
    .Q(\systolic_array.arg_left_div2_next[1] ));
 sg13g2_dfrbp_1 _4085_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net309),
    .D(net753),
    .Q_N(_1886_),
    .Q(\systolic_array.genblk2[0].mac[0].mul2 ));
 sg13g2_dfrbp_1 _4086_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net308),
    .D(net544),
    .Q_N(_1885_),
    .Q(\systolic_array.genblk2[0].mac[1].mul2 ));
 sg13g2_dfrbp_1 _4087_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net307),
    .D(net751),
    .Q_N(_1884_),
    .Q(\systolic_array.genblk2[0].mac[2].mul2 ));
 sg13g2_dfrbp_1 _4088_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net306),
    .D(net891),
    .Q_N(_1883_),
    .Q(\systolic_array.genblk2[0].mac[3].mul2 ));
 sg13g2_dfrbp_1 _4089_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net305),
    .D(_0165_),
    .Q_N(_1882_),
    .Q(\systolic_array.genblk2[0].mac[4].mul2 ));
 sg13g2_dfrbp_1 _4090_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net304),
    .D(_0166_),
    .Q_N(_1881_),
    .Q(\systolic_array.genblk2[0].mac[5].mul2 ));
 sg13g2_dfrbp_1 _4091_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net303),
    .D(net794),
    .Q_N(_1880_),
    .Q(\systolic_array.genblk2[0].mac[0].sign ));
 sg13g2_dfrbp_1 _4092_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net302),
    .D(net773),
    .Q_N(_1879_),
    .Q(\systolic_array.genblk2[0].mac[1].sign ));
 sg13g2_dfrbp_1 _4093_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net301),
    .D(net537),
    .Q_N(_1878_),
    .Q(\systolic_array.genblk2[0].mac[2].sign ));
 sg13g2_dfrbp_1 _4094_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net300),
    .D(_0170_),
    .Q_N(_1877_),
    .Q(\systolic_array.genblk2[0].mac[3].sign ));
 sg13g2_dfrbp_1 _4095_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net299),
    .D(_0171_),
    .Q_N(_1876_),
    .Q(\systolic_array.genblk2[0].mac[4].sign ));
 sg13g2_dfrbp_1 _4096_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net298),
    .D(net823),
    .Q_N(_1875_),
    .Q(\systolic_array.genblk2[0].mac[5].sign ));
 sg13g2_dfrbp_1 _4097_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net297),
    .D(_0173_),
    .Q_N(_1874_),
    .Q(\systolic_array.genblk2[0].mac[0].zero ));
 sg13g2_dfrbp_1 _4098_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net296),
    .D(_0174_),
    .Q_N(_1873_),
    .Q(\systolic_array.genblk2[0].mac[1].zero ));
 sg13g2_dfrbp_1 _4099_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net295),
    .D(_0175_),
    .Q_N(_1872_),
    .Q(\systolic_array.genblk2[0].mac[2].zero ));
 sg13g2_dfrbp_1 _4100_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net294),
    .D(_0176_),
    .Q_N(_1871_),
    .Q(\systolic_array.genblk2[0].mac[3].zero ));
 sg13g2_dfrbp_1 _4101_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net293),
    .D(_0177_),
    .Q_N(_1870_),
    .Q(\systolic_array.genblk2[0].mac[4].zero ));
 sg13g2_dfrbp_1 _4102_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net292),
    .D(_0178_),
    .Q_N(_1869_),
    .Q(\systolic_array.genblk2[0].mac[5].zero ));
 sg13g2_dfrbp_1 _4103_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net291),
    .D(_0179_),
    .Q_N(_1868_),
    .Q(\systolic_array.arg_left_mul2_next[0] ));
 sg13g2_dfrbp_1 _4104_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net290),
    .D(_0180_),
    .Q_N(_1867_),
    .Q(\systolic_array.arg_left_mul2_next[1] ));
 sg13g2_dfrbp_1 _4105_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net289),
    .D(_0181_),
    .Q_N(_1866_),
    .Q(\systolic_array.arg_left_mul2_next[2] ));
 sg13g2_dfrbp_1 _4106_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net288),
    .D(_0182_),
    .Q_N(_1865_),
    .Q(\systolic_array.arg_left_zero_next[3] ));
 sg13g2_dfrbp_1 _4107_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net287),
    .D(_0183_),
    .Q_N(_1864_),
    .Q(\systolic_array.arg_left_zero_next[4] ));
 sg13g2_dfrbp_1 _4108_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net286),
    .D(_0184_),
    .Q_N(_1863_),
    .Q(\systolic_array.arg_left_zero_next[5] ));
 sg13g2_dfrbp_1 _4109_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net285),
    .D(_0185_),
    .Q_N(_1862_),
    .Q(\systolic_array.arg_left_sign_next[4] ));
 sg13g2_dfrbp_1 _4110_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net284),
    .D(_0186_),
    .Q_N(_1861_),
    .Q(\systolic_array.arg_left_sign_next[5] ));
 sg13g2_dfrbp_1 _4111_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net283),
    .D(_0187_),
    .Q_N(_1860_),
    .Q(\systolic_array.arg_left_mul2_next[3] ));
 sg13g2_dfrbp_1 _4112_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net282),
    .D(_0188_),
    .Q_N(_1859_),
    .Q(\systolic_array.arg_left_mul2_next[4] ));
 sg13g2_dfrbp_1 _4113_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net281),
    .D(_0189_),
    .Q_N(_1858_),
    .Q(\systolic_array.arg_left_mul2_next[5] ));
 sg13g2_dfrbp_1 _4114_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net280),
    .D(_0190_),
    .Q_N(_1857_),
    .Q(\systolic_array.arg_left_div2_next[3] ));
 sg13g2_dfrbp_1 _4115_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net279),
    .D(_0191_),
    .Q_N(_1856_),
    .Q(\systolic_array.arg_left_div2_next[4] ));
 sg13g2_dfrbp_1 _4116_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net278),
    .D(_0192_),
    .Q_N(_1665_),
    .Q(\systolic_array.slice_counter ));
 sg13g2_dfrbp_1 _4117_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net277),
    .D(_0193_),
    .Q_N(_1855_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[0].A ));
 sg13g2_dfrbp_1 _4118_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net276),
    .D(_0194_),
    .Q_N(_1854_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[1].A ));
 sg13g2_dfrbp_1 _4119_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net275),
    .D(_0195_),
    .Q_N(_1853_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[2].A ));
 sg13g2_dfrbp_1 _4120_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net274),
    .D(_0196_),
    .Q_N(_1852_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[3].A ));
 sg13g2_dfrbp_1 _4121_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net273),
    .D(_0197_),
    .Q_N(_1851_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[4].A ));
 sg13g2_dfrbp_1 _4122_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net272),
    .D(_0198_),
    .Q_N(_1850_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[5].A ));
 sg13g2_dfrbp_1 _4123_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net271),
    .D(_0199_),
    .Q_N(_1849_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[6].A ));
 sg13g2_dfrbp_1 _4124_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net270),
    .D(_0200_),
    .Q_N(_1848_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[7].A ));
 sg13g2_dfrbp_1 _4125_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net269),
    .D(_0201_),
    .Q_N(_1847_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[8].A ));
 sg13g2_dfrbp_1 _4126_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net268),
    .D(_0202_),
    .Q_N(_0114_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[9].A ));
 sg13g2_dfrbp_1 _4127_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net267),
    .D(_0203_),
    .Q_N(_1846_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[10].A ));
 sg13g2_dfrbp_1 _4128_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net266),
    .D(_0204_),
    .Q_N(_0117_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[11].A ));
 sg13g2_dfrbp_1 _4129_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net265),
    .D(_0205_),
    .Q_N(_1845_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[12].A ));
 sg13g2_dfrbp_1 _4130_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net264),
    .D(_0206_),
    .Q_N(_0118_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[13].A ));
 sg13g2_dfrbp_1 _4131_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net263),
    .D(_0207_),
    .Q_N(_1844_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[14].A ));
 sg13g2_dfrbp_1 _4132_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net262),
    .D(_0208_),
    .Q_N(_1843_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[15].A ));
 sg13g2_dfrbp_1 _4133_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net261),
    .D(_0209_),
    .Q_N(_1842_),
    .Q(\systolic_array.genblk1[0].accumulators_dlygate[16].A ));
 sg13g2_dfrbp_1 _4134_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net260),
    .D(_0210_),
    .Q_N(_1841_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[0].A ));
 sg13g2_dfrbp_1 _4135_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net259),
    .D(net880),
    .Q_N(_1840_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[1].A ));
 sg13g2_dfrbp_1 _4136_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net258),
    .D(_0212_),
    .Q_N(_1839_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[2].A ));
 sg13g2_dfrbp_1 _4137_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net257),
    .D(_0213_),
    .Q_N(_1838_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[3].A ));
 sg13g2_dfrbp_1 _4138_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net256),
    .D(net903),
    .Q_N(_1837_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[4].A ));
 sg13g2_dfrbp_1 _4139_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net255),
    .D(_0215_),
    .Q_N(_1836_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[5].A ));
 sg13g2_dfrbp_1 _4140_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net254),
    .D(_0216_),
    .Q_N(_1835_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[6].A ));
 sg13g2_dfrbp_1 _4141_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net253),
    .D(_0217_),
    .Q_N(_1834_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[7].A ));
 sg13g2_dfrbp_1 _4142_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net252),
    .D(net837),
    .Q_N(_1833_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[8].A ));
 sg13g2_dfrbp_1 _4143_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net251),
    .D(_0219_),
    .Q_N(_1832_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[9].A ));
 sg13g2_dfrbp_1 _4144_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net250),
    .D(_0220_),
    .Q_N(_1831_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[10].A ));
 sg13g2_dfrbp_1 _4145_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net249),
    .D(_0221_),
    .Q_N(_1830_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[11].A ));
 sg13g2_dfrbp_1 _4146_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net248),
    .D(_0222_),
    .Q_N(_1829_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[12].A ));
 sg13g2_dfrbp_1 _4147_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net247),
    .D(_0223_),
    .Q_N(_1828_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[13].A ));
 sg13g2_dfrbp_1 _4148_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net246),
    .D(_0224_),
    .Q_N(_1827_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[14].A ));
 sg13g2_dfrbp_1 _4149_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net245),
    .D(_0225_),
    .Q_N(_1826_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[15].A ));
 sg13g2_dfrbp_1 _4150_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net244),
    .D(_0226_),
    .Q_N(_1825_),
    .Q(\systolic_array.genblk1[1].accumulators_dlygate[16].A ));
 sg13g2_dfrbp_1 _4151_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net243),
    .D(_0227_),
    .Q_N(_1824_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[0].A ));
 sg13g2_dfrbp_1 _4152_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net242),
    .D(_0228_),
    .Q_N(_1823_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[1].A ));
 sg13g2_dfrbp_1 _4153_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net241),
    .D(_0229_),
    .Q_N(_1822_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[2].A ));
 sg13g2_dfrbp_1 _4154_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net240),
    .D(_0230_),
    .Q_N(_1821_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[3].A ));
 sg13g2_dfrbp_1 _4155_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net239),
    .D(_0231_),
    .Q_N(_1820_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[4].A ));
 sg13g2_dfrbp_1 _4156_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net238),
    .D(_0232_),
    .Q_N(_1819_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[5].A ));
 sg13g2_dfrbp_1 _4157_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net237),
    .D(_0233_),
    .Q_N(_1818_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[6].A ));
 sg13g2_dfrbp_1 _4158_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net236),
    .D(_0234_),
    .Q_N(_1817_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[7].A ));
 sg13g2_dfrbp_1 _4159_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net235),
    .D(_0235_),
    .Q_N(_1816_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[8].A ));
 sg13g2_dfrbp_1 _4160_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net234),
    .D(_0236_),
    .Q_N(_0119_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[9].A ));
 sg13g2_dfrbp_1 _4161_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net233),
    .D(_0237_),
    .Q_N(_1815_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[10].A ));
 sg13g2_dfrbp_1 _4162_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net232),
    .D(_0238_),
    .Q_N(_0096_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[11].A ));
 sg13g2_dfrbp_1 _4163_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net231),
    .D(_0239_),
    .Q_N(_1814_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[12].A ));
 sg13g2_dfrbp_1 _4164_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net230),
    .D(_0240_),
    .Q_N(_0097_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[13].A ));
 sg13g2_dfrbp_1 _4165_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net229),
    .D(_0241_),
    .Q_N(_1813_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[14].A ));
 sg13g2_dfrbp_1 _4166_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net228),
    .D(_0242_),
    .Q_N(_1812_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[15].A ));
 sg13g2_dfrbp_1 _4167_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net227),
    .D(_0243_),
    .Q_N(_1811_),
    .Q(\systolic_array.genblk1[2].accumulators_dlygate[16].A ));
 sg13g2_dfrbp_1 _4168_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net226),
    .D(_0244_),
    .Q_N(_1810_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[0].A ));
 sg13g2_dfrbp_1 _4169_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net225),
    .D(_0245_),
    .Q_N(_1809_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[1].A ));
 sg13g2_dfrbp_1 _4170_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net224),
    .D(_0246_),
    .Q_N(_1808_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[2].A ));
 sg13g2_dfrbp_1 _4171_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net223),
    .D(_0247_),
    .Q_N(_1807_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[3].A ));
 sg13g2_dfrbp_1 _4172_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net222),
    .D(_0248_),
    .Q_N(_1806_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[4].A ));
 sg13g2_dfrbp_1 _4173_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net221),
    .D(_0249_),
    .Q_N(_1805_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[5].A ));
 sg13g2_dfrbp_1 _4174_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net220),
    .D(net897),
    .Q_N(_1804_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[6].A ));
 sg13g2_dfrbp_1 _4175_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net219),
    .D(_0251_),
    .Q_N(_1803_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[7].A ));
 sg13g2_dfrbp_1 _4176_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net218),
    .D(_0252_),
    .Q_N(_1802_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[8].A ));
 sg13g2_dfrbp_1 _4177_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net217),
    .D(_0253_),
    .Q_N(_1801_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[9].A ));
 sg13g2_dfrbp_1 _4178_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net216),
    .D(_0254_),
    .Q_N(_1800_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[10].A ));
 sg13g2_dfrbp_1 _4179_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net215),
    .D(_0255_),
    .Q_N(_1799_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[11].A ));
 sg13g2_dfrbp_1 _4180_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net214),
    .D(_0256_),
    .Q_N(_1798_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[12].A ));
 sg13g2_dfrbp_1 _4181_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net213),
    .D(_0257_),
    .Q_N(_1797_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[13].A ));
 sg13g2_dfrbp_1 _4182_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net212),
    .D(_0258_),
    .Q_N(_1796_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[14].A ));
 sg13g2_dfrbp_1 _4183_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net211),
    .D(_0259_),
    .Q_N(_1795_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[15].A ));
 sg13g2_dfrbp_1 _4184_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net210),
    .D(_0260_),
    .Q_N(_1794_),
    .Q(\systolic_array.genblk1[3].accumulators_dlygate[16].A ));
 sg13g2_dfrbp_1 _4185_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net209),
    .D(_0261_),
    .Q_N(_1793_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[0].A ));
 sg13g2_dfrbp_1 _4186_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net208),
    .D(_0262_),
    .Q_N(_1792_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[1].A ));
 sg13g2_dfrbp_1 _4187_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net207),
    .D(_0263_),
    .Q_N(_1791_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[2].A ));
 sg13g2_dfrbp_1 _4188_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net206),
    .D(_0264_),
    .Q_N(_1790_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[3].A ));
 sg13g2_dfrbp_1 _4189_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net205),
    .D(_0265_),
    .Q_N(_1789_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[4].A ));
 sg13g2_dfrbp_1 _4190_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net204),
    .D(_0266_),
    .Q_N(_1788_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[5].A ));
 sg13g2_dfrbp_1 _4191_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net203),
    .D(_0267_),
    .Q_N(_1787_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[6].A ));
 sg13g2_dfrbp_1 _4192_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net202),
    .D(_0268_),
    .Q_N(_1786_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[7].A ));
 sg13g2_dfrbp_1 _4193_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net201),
    .D(_0269_),
    .Q_N(_1785_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[8].A ));
 sg13g2_dfrbp_1 _4194_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net200),
    .D(_0270_),
    .Q_N(_0098_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[9].A ));
 sg13g2_dfrbp_1 _4195_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net199),
    .D(_0271_),
    .Q_N(_1784_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[10].A ));
 sg13g2_dfrbp_1 _4196_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net198),
    .D(_0272_),
    .Q_N(_0102_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[11].A ));
 sg13g2_dfrbp_1 _4197_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net197),
    .D(_0273_),
    .Q_N(_1783_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[12].A ));
 sg13g2_dfrbp_1 _4198_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net196),
    .D(_0274_),
    .Q_N(_0103_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[13].A ));
 sg13g2_dfrbp_1 _4199_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net195),
    .D(_0275_),
    .Q_N(_1782_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[14].A ));
 sg13g2_dfrbp_1 _4200_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net194),
    .D(_0276_),
    .Q_N(_1781_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[15].A ));
 sg13g2_dfrbp_1 _4201_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net193),
    .D(_0277_),
    .Q_N(_1780_),
    .Q(\systolic_array.genblk1[4].accumulators_dlygate[16].A ));
 sg13g2_dfrbp_1 _4202_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net192),
    .D(_0278_),
    .Q_N(_1779_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[0].A ));
 sg13g2_dfrbp_1 _4203_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net191),
    .D(net846),
    .Q_N(_1778_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[1].A ));
 sg13g2_dfrbp_1 _4204_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net190),
    .D(net855),
    .Q_N(_1777_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[2].A ));
 sg13g2_dfrbp_1 _4205_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net189),
    .D(_0281_),
    .Q_N(_1776_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[3].A ));
 sg13g2_dfrbp_1 _4206_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net188),
    .D(_0282_),
    .Q_N(_1775_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[4].A ));
 sg13g2_dfrbp_1 _4207_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net187),
    .D(_0283_),
    .Q_N(_1774_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[5].A ));
 sg13g2_dfrbp_1 _4208_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net186),
    .D(net875),
    .Q_N(_1773_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[6].A ));
 sg13g2_dfrbp_1 _4209_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net185),
    .D(net934),
    .Q_N(_1772_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[7].A ));
 sg13g2_dfrbp_1 _4210_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net184),
    .D(_0286_),
    .Q_N(_1771_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[8].A ));
 sg13g2_dfrbp_1 _4211_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net183),
    .D(_0287_),
    .Q_N(_1770_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[9].A ));
 sg13g2_dfrbp_1 _4212_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net182),
    .D(_0288_),
    .Q_N(_1769_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[10].A ));
 sg13g2_dfrbp_1 _4213_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net181),
    .D(_0289_),
    .Q_N(_1768_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[11].A ));
 sg13g2_dfrbp_1 _4214_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net180),
    .D(_0290_),
    .Q_N(_1767_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[12].A ));
 sg13g2_dfrbp_1 _4215_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net179),
    .D(_0291_),
    .Q_N(_1766_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[13].A ));
 sg13g2_dfrbp_1 _4216_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net178),
    .D(_0292_),
    .Q_N(_1765_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[14].A ));
 sg13g2_dfrbp_1 _4217_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net177),
    .D(_0293_),
    .Q_N(_1764_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[15].A ));
 sg13g2_dfrbp_1 _4218_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net176),
    .D(_0294_),
    .Q_N(_1763_),
    .Q(\systolic_array.genblk1[5].accumulators_dlygate[16].A ));
 sg13g2_dfrbp_1 _4219_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net175),
    .D(_0295_),
    .Q_N(_1762_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[0].A ));
 sg13g2_dfrbp_1 _4220_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net174),
    .D(_0296_),
    .Q_N(_1761_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[1].A ));
 sg13g2_dfrbp_1 _4221_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net173),
    .D(_0297_),
    .Q_N(_1760_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[2].A ));
 sg13g2_dfrbp_1 _4222_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net172),
    .D(_0298_),
    .Q_N(_1759_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[3].A ));
 sg13g2_dfrbp_1 _4223_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net171),
    .D(_0299_),
    .Q_N(_1758_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[4].A ));
 sg13g2_dfrbp_1 _4224_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net170),
    .D(_0300_),
    .Q_N(_1757_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[5].A ));
 sg13g2_dfrbp_1 _4225_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net169),
    .D(_0301_),
    .Q_N(_1756_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[6].A ));
 sg13g2_dfrbp_1 _4226_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net168),
    .D(_0302_),
    .Q_N(_1755_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[7].A ));
 sg13g2_dfrbp_1 _4227_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net167),
    .D(_0303_),
    .Q_N(_1754_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[8].A ));
 sg13g2_dfrbp_1 _4228_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net166),
    .D(_0304_),
    .Q_N(_0104_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[9].A ));
 sg13g2_dfrbp_1 _4229_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net165),
    .D(_0305_),
    .Q_N(_1753_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[10].A ));
 sg13g2_dfrbp_1 _4230_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net164),
    .D(_0306_),
    .Q_N(_0106_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[11].A ));
 sg13g2_dfrbp_1 _4231_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net163),
    .D(_0307_),
    .Q_N(_1752_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[12].A ));
 sg13g2_dfrbp_1 _4232_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net162),
    .D(_0308_),
    .Q_N(_0107_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[13].A ));
 sg13g2_dfrbp_1 _4233_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net161),
    .D(_0309_),
    .Q_N(_1751_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[14].A ));
 sg13g2_dfrbp_1 _4234_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net160),
    .D(_0310_),
    .Q_N(_1750_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[15].A ));
 sg13g2_dfrbp_1 _4235_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net159),
    .D(_0311_),
    .Q_N(_1749_),
    .Q(\systolic_array.genblk1[6].accumulators_dlygate[16].A ));
 sg13g2_dfrbp_1 _4236_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net158),
    .D(_0312_),
    .Q_N(_1748_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[0].A ));
 sg13g2_dfrbp_1 _4237_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net157),
    .D(_0313_),
    .Q_N(_1747_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[1].A ));
 sg13g2_dfrbp_1 _4238_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net156),
    .D(_0314_),
    .Q_N(_1746_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[2].A ));
 sg13g2_dfrbp_1 _4239_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net155),
    .D(_0315_),
    .Q_N(_1745_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[3].A ));
 sg13g2_dfrbp_1 _4240_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net154),
    .D(_0316_),
    .Q_N(_1744_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[4].A ));
 sg13g2_dfrbp_1 _4241_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net153),
    .D(_0317_),
    .Q_N(_1743_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[5].A ));
 sg13g2_dfrbp_1 _4242_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net152),
    .D(net882),
    .Q_N(_1742_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[6].A ));
 sg13g2_dfrbp_1 _4243_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net151),
    .D(net924),
    .Q_N(_1741_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[7].A ));
 sg13g2_dfrbp_1 _4244_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net150),
    .D(_0320_),
    .Q_N(_1740_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[8].A ));
 sg13g2_dfrbp_1 _4245_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net149),
    .D(_0321_),
    .Q_N(_1739_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[9].A ));
 sg13g2_dfrbp_1 _4246_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net148),
    .D(_0322_),
    .Q_N(_1738_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[10].A ));
 sg13g2_dfrbp_1 _4247_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net147),
    .D(_0323_),
    .Q_N(_1737_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[11].A ));
 sg13g2_dfrbp_1 _4248_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net146),
    .D(_0324_),
    .Q_N(_1736_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[12].A ));
 sg13g2_dfrbp_1 _4249_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net145),
    .D(_0325_),
    .Q_N(_1735_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[13].A ));
 sg13g2_dfrbp_1 _4250_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net144),
    .D(_0326_),
    .Q_N(_1734_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[14].A ));
 sg13g2_dfrbp_1 _4251_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net143),
    .D(_0327_),
    .Q_N(_1733_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[15].A ));
 sg13g2_dfrbp_1 _4252_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net142),
    .D(_0328_),
    .Q_N(_1732_),
    .Q(\systolic_array.genblk1[7].accumulators_dlygate[16].A ));
 sg13g2_dfrbp_1 _4253_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net141),
    .D(_0329_),
    .Q_N(_1731_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[0].A ));
 sg13g2_dfrbp_1 _4254_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net140),
    .D(_0330_),
    .Q_N(_1730_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[1].A ));
 sg13g2_dfrbp_1 _4255_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net139),
    .D(_0331_),
    .Q_N(_1729_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[2].A ));
 sg13g2_dfrbp_1 _4256_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net138),
    .D(_0332_),
    .Q_N(_1728_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[3].A ));
 sg13g2_dfrbp_1 _4257_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net137),
    .D(_0333_),
    .Q_N(_1727_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[4].A ));
 sg13g2_dfrbp_1 _4258_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net136),
    .D(_0334_),
    .Q_N(_1726_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[5].A ));
 sg13g2_dfrbp_1 _4259_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net135),
    .D(_0335_),
    .Q_N(_1725_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[6].A ));
 sg13g2_dfrbp_1 _4260_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net134),
    .D(_0336_),
    .Q_N(_1724_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[7].A ));
 sg13g2_dfrbp_1 _4261_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net133),
    .D(_0337_),
    .Q_N(_1723_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[8].A ));
 sg13g2_dfrbp_1 _4262_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net132),
    .D(_0338_),
    .Q_N(_0108_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[9].A ));
 sg13g2_dfrbp_1 _4263_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net131),
    .D(_0339_),
    .Q_N(_1722_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[10].A ));
 sg13g2_dfrbp_1 _4264_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net130),
    .D(_0340_),
    .Q_N(_0109_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[11].A ));
 sg13g2_dfrbp_1 _4265_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net129),
    .D(_0341_),
    .Q_N(_1721_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[12].A ));
 sg13g2_dfrbp_1 _4266_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net128),
    .D(_0342_),
    .Q_N(_0110_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[13].A ));
 sg13g2_dfrbp_1 _4267_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net127),
    .D(_0343_),
    .Q_N(_1720_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[14].A ));
 sg13g2_dfrbp_1 _4268_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net126),
    .D(_0344_),
    .Q_N(_1719_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[15].A ));
 sg13g2_dfrbp_1 _4269_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net125),
    .D(_0345_),
    .Q_N(_1718_),
    .Q(\systolic_array.genblk1[8].accumulators_dlygate[16].A ));
 sg13g2_dfrbp_1 _4270_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net124),
    .D(_0346_),
    .Q_N(_1717_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[0].A ));
 sg13g2_dfrbp_1 _4271_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net123),
    .D(net939),
    .Q_N(_1716_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[1].A ));
 sg13g2_dfrbp_1 _4272_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net122),
    .D(_0348_),
    .Q_N(_1715_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[2].A ));
 sg13g2_dfrbp_1 _4273_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net121),
    .D(_0349_),
    .Q_N(_1714_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[3].A ));
 sg13g2_dfrbp_1 _4274_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net120),
    .D(_0350_),
    .Q_N(_1713_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[4].A ));
 sg13g2_dfrbp_1 _4275_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net119),
    .D(net972),
    .Q_N(_1712_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[5].A ));
 sg13g2_dfrbp_1 _4276_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net118),
    .D(_0352_),
    .Q_N(_1711_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[6].A ));
 sg13g2_dfrbp_1 _4277_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net117),
    .D(_0353_),
    .Q_N(_1710_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[7].A ));
 sg13g2_dfrbp_1 _4278_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net116),
    .D(_0354_),
    .Q_N(_1709_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[8].A ));
 sg13g2_dfrbp_1 _4279_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net115),
    .D(_0355_),
    .Q_N(_1708_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[9].A ));
 sg13g2_dfrbp_1 _4280_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net114),
    .D(_0356_),
    .Q_N(_1707_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[10].A ));
 sg13g2_dfrbp_1 _4281_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net113),
    .D(_0357_),
    .Q_N(_1706_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[11].A ));
 sg13g2_dfrbp_1 _4282_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net112),
    .D(_0358_),
    .Q_N(_1705_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[12].A ));
 sg13g2_dfrbp_1 _4283_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net111),
    .D(_0359_),
    .Q_N(_1704_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[13].A ));
 sg13g2_dfrbp_1 _4284_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net110),
    .D(_0360_),
    .Q_N(_1703_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[14].A ));
 sg13g2_dfrbp_1 _4285_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net109),
    .D(_0361_),
    .Q_N(_1702_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[15].A ));
 sg13g2_dfrbp_1 _4286_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net108),
    .D(_0362_),
    .Q_N(_1701_),
    .Q(\systolic_array.genblk1[9].accumulators_dlygate[16].A ));
 sg13g2_dfrbp_1 _4287_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net107),
    .D(net799),
    .Q_N(_1700_),
    .Q(\systolic_array.genblk2[0].mac[0].div2 ));
 sg13g2_dfrbp_1 _4288_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net106),
    .D(net505),
    .Q_N(_1699_),
    .Q(\systolic_array.genblk2[0].mac[1].div2 ));
 sg13g2_dfrbp_1 _4289_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net105),
    .D(_0365_),
    .Q_N(_1698_),
    .Q(\systolic_array.genblk2[0].mac[3].div2 ));
 sg13g2_dfrbp_1 _4290_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net333),
    .D(_0366_),
    .Q_N(_1930_),
    .Q(\systolic_array.genblk2[0].mac[4].div2 ));
 sg13g2_dfrbp_1 _4291_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net334),
    .D(_0023_),
    .Q_N(_1931_),
    .Q(\systolic_array.genblk1[10].out_queue_dlygate[9].A ));
 sg13g2_dfrbp_1 _4292_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net335),
    .D(net747),
    .Q_N(_1932_),
    .Q(\systolic_array.genblk1[10].out_queue_dlygate[10].A ));
 sg13g2_dfrbp_1 _4293_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net336),
    .D(net762),
    .Q_N(_1933_),
    .Q(\systolic_array.genblk1[10].out_queue_dlygate[11].A ));
 sg13g2_dfrbp_1 _4294_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net337),
    .D(net758),
    .Q_N(_1934_),
    .Q(\systolic_array.genblk1[10].out_queue_dlygate[12].A ));
 sg13g2_dfrbp_1 _4295_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net338),
    .D(_0019_),
    .Q_N(_1935_),
    .Q(\systolic_array.genblk1[10].out_queue_dlygate[13].A ));
 sg13g2_dfrbp_1 _4296_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net339),
    .D(net534),
    .Q_N(_1936_),
    .Q(\systolic_array.genblk1[10].out_queue_dlygate[14].A ));
 sg13g2_dfrbp_1 _4297_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net357),
    .D(net731),
    .Q_N(_1937_),
    .Q(\systolic_array.genblk1[10].out_queue_dlygate[15].A ));
 sg13g2_dfrbp_1 _4298_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net104),
    .D(_0022_),
    .Q_N(_1697_),
    .Q(\systolic_array.genblk1[10].out_queue_dlygate[16].A ));
 sg13g2_dfrbp_1 _4299_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net103),
    .D(_0367_),
    .Q_N(_1696_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[0].A ));
 sg13g2_dfrbp_1 _4300_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net102),
    .D(net859),
    .Q_N(_1695_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[1].A ));
 sg13g2_dfrbp_1 _4301_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net101),
    .D(net950),
    .Q_N(_1694_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[2].A ));
 sg13g2_dfrbp_1 _4302_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net100),
    .D(_0370_),
    .Q_N(_1693_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[3].A ));
 sg13g2_dfrbp_1 _4303_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net99),
    .D(_0371_),
    .Q_N(_1692_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[4].A ));
 sg13g2_dfrbp_1 _4304_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net98),
    .D(net899),
    .Q_N(_1691_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[5].A ));
 sg13g2_dfrbp_1 _4305_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net97),
    .D(_0373_),
    .Q_N(_1690_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[6].A ));
 sg13g2_dfrbp_1 _4306_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net96),
    .D(_0374_),
    .Q_N(_1689_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[7].A ));
 sg13g2_dfrbp_1 _4307_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net95),
    .D(_0375_),
    .Q_N(_1688_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[8].A ));
 sg13g2_dfrbp_1 _4308_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net94),
    .D(_0376_),
    .Q_N(_1687_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[9].A ));
 sg13g2_dfrbp_1 _4309_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net93),
    .D(_0377_),
    .Q_N(_1686_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[10].A ));
 sg13g2_dfrbp_1 _4310_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net92),
    .D(_0378_),
    .Q_N(_1685_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[11].A ));
 sg13g2_dfrbp_1 _4311_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net91),
    .D(_0379_),
    .Q_N(_1684_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[12].A ));
 sg13g2_dfrbp_1 _4312_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net90),
    .D(_0380_),
    .Q_N(_1683_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[13].A ));
 sg13g2_dfrbp_1 _4313_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net89),
    .D(_0381_),
    .Q_N(_1682_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[14].A ));
 sg13g2_dfrbp_1 _4314_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net88),
    .D(_0382_),
    .Q_N(_1681_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[15].A ));
 sg13g2_dfrbp_1 _4315_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net358),
    .D(_0383_),
    .Q_N(_1938_),
    .Q(\systolic_array.genblk1[11].accumulators_dlygate[16].A ));
 sg13g2_dfrbp_1 _4316_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net359),
    .D(net749),
    .Q_N(_1939_),
    .Q(\systolic_array.genblk1[8].out_queue_dlygate[9].A ));
 sg13g2_dfrbp_1 _4317_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net360),
    .D(net540),
    .Q_N(_1940_),
    .Q(\systolic_array.genblk1[8].out_queue_dlygate[10].A ));
 sg13g2_dfrbp_1 _4318_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net361),
    .D(net727),
    .Q_N(_1941_),
    .Q(\systolic_array.genblk1[8].out_queue_dlygate[11].A ));
 sg13g2_dfrbp_1 _4319_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net362),
    .D(net755),
    .Q_N(_1942_),
    .Q(\systolic_array.genblk1[8].out_queue_dlygate[12].A ));
 sg13g2_dfrbp_1 _4320_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net363),
    .D(net770),
    .Q_N(_1943_),
    .Q(\systolic_array.genblk1[8].out_queue_dlygate[13].A ));
 sg13g2_dfrbp_1 _4321_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net364),
    .D(net857),
    .Q_N(_1944_),
    .Q(\systolic_array.genblk1[8].out_queue_dlygate[14].A ));
 sg13g2_dfrbp_1 _4322_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net365),
    .D(net729),
    .Q_N(_1945_),
    .Q(\systolic_array.genblk1[8].out_queue_dlygate[15].A ));
 sg13g2_dfrbp_1 _4323_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net366),
    .D(net788),
    .Q_N(_1946_),
    .Q(\systolic_array.genblk1[8].out_queue_dlygate[16].A ));
 sg13g2_dfrbp_1 _4324_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net367),
    .D(_0095_),
    .Q_N(_1947_),
    .Q(\systolic_array.genblk1[9].out_queue_dlygate[9].A ));
 sg13g2_dfrbp_1 _4325_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net368),
    .D(_0088_),
    .Q_N(_1948_),
    .Q(\systolic_array.genblk1[9].out_queue_dlygate[10].A ));
 sg13g2_dfrbp_1 _4326_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net369),
    .D(_0089_),
    .Q_N(_1949_),
    .Q(\systolic_array.genblk1[9].out_queue_dlygate[11].A ));
 sg13g2_dfrbp_1 _4327_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net370),
    .D(_0090_),
    .Q_N(_1950_),
    .Q(\systolic_array.genblk1[9].out_queue_dlygate[12].A ));
 sg13g2_dfrbp_1 _4328_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net371),
    .D(_0091_),
    .Q_N(_1951_),
    .Q(\systolic_array.genblk1[9].out_queue_dlygate[13].A ));
 sg13g2_dfrbp_1 _4329_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net372),
    .D(_0092_),
    .Q_N(_1952_),
    .Q(\systolic_array.genblk1[9].out_queue_dlygate[14].A ));
 sg13g2_dfrbp_1 _4330_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net373),
    .D(_0093_),
    .Q_N(_1953_),
    .Q(\systolic_array.genblk1[9].out_queue_dlygate[15].A ));
 sg13g2_dfrbp_1 _4331_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net374),
    .D(_0094_),
    .Q_N(_1954_),
    .Q(\systolic_array.genblk1[9].out_queue_dlygate[16].A ));
 sg13g2_dfrbp_1 _4332_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net375),
    .D(net905),
    .Q_N(_1955_),
    .Q(\systolic_array.genblk1[6].out_queue_dlygate[9].A ));
 sg13g2_dfrbp_1 _4333_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net376),
    .D(net870),
    .Q_N(_1956_),
    .Q(\systolic_array.genblk1[6].out_queue_dlygate[10].A ));
 sg13g2_dfrbp_1 _4334_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net377),
    .D(net910),
    .Q_N(_1957_),
    .Q(\systolic_array.genblk1[6].out_queue_dlygate[11].A ));
 sg13g2_dfrbp_1 _4335_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net378),
    .D(_0066_),
    .Q_N(_1958_),
    .Q(\systolic_array.genblk1[6].out_queue_dlygate[12].A ));
 sg13g2_dfrbp_1 _4336_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net379),
    .D(net839),
    .Q_N(_1959_),
    .Q(\systolic_array.genblk1[6].out_queue_dlygate[13].A ));
 sg13g2_dfrbp_1 _4337_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net380),
    .D(net737),
    .Q_N(_1960_),
    .Q(\systolic_array.genblk1[6].out_queue_dlygate[14].A ));
 sg13g2_dfrbp_1 _4338_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net381),
    .D(_0069_),
    .Q_N(_1961_),
    .Q(\systolic_array.genblk1[6].out_queue_dlygate[15].A ));
 sg13g2_dfrbp_1 _4339_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net382),
    .D(net725),
    .Q_N(_1962_),
    .Q(\systolic_array.genblk1[6].out_queue_dlygate[16].A ));
 sg13g2_dfrbp_1 _4340_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net383),
    .D(_0079_),
    .Q_N(_1963_),
    .Q(\systolic_array.genblk1[7].out_queue_dlygate[9].A ));
 sg13g2_dfrbp_1 _4341_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net384),
    .D(_0072_),
    .Q_N(_1964_),
    .Q(\systolic_array.genblk1[7].out_queue_dlygate[10].A ));
 sg13g2_dfrbp_1 _4342_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net385),
    .D(_0073_),
    .Q_N(_1965_),
    .Q(\systolic_array.genblk1[7].out_queue_dlygate[11].A ));
 sg13g2_dfrbp_1 _4343_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net386),
    .D(_0074_),
    .Q_N(_1966_),
    .Q(\systolic_array.genblk1[7].out_queue_dlygate[12].A ));
 sg13g2_dfrbp_1 _4344_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net387),
    .D(_0075_),
    .Q_N(_1967_),
    .Q(\systolic_array.genblk1[7].out_queue_dlygate[13].A ));
 sg13g2_dfrbp_1 _4345_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net388),
    .D(_0076_),
    .Q_N(_1968_),
    .Q(\systolic_array.genblk1[7].out_queue_dlygate[14].A ));
 sg13g2_dfrbp_1 _4346_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net389),
    .D(_0077_),
    .Q_N(_1969_),
    .Q(\systolic_array.genblk1[7].out_queue_dlygate[15].A ));
 sg13g2_dfrbp_1 _4347_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net390),
    .D(_0078_),
    .Q_N(_1970_),
    .Q(\systolic_array.genblk1[7].out_queue_dlygate[16].A ));
 sg13g2_dfrbp_1 _4348_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net391),
    .D(net807),
    .Q_N(_1971_),
    .Q(\systolic_array.genblk1[4].out_queue_dlygate[9].A ));
 sg13g2_dfrbp_1 _4349_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net392),
    .D(net829),
    .Q_N(_1972_),
    .Q(\systolic_array.genblk1[4].out_queue_dlygate[10].A ));
 sg13g2_dfrbp_1 _4350_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net393),
    .D(net768),
    .Q_N(_1973_),
    .Q(\systolic_array.genblk1[4].out_queue_dlygate[11].A ));
 sg13g2_dfrbp_1 _4351_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net394),
    .D(_0050_),
    .Q_N(_1974_),
    .Q(\systolic_array.genblk1[4].out_queue_dlygate[12].A ));
 sg13g2_dfrbp_1 _4352_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net395),
    .D(net931),
    .Q_N(_1975_),
    .Q(\systolic_array.genblk1[4].out_queue_dlygate[13].A ));
 sg13g2_dfrbp_1 _4353_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net396),
    .D(net542),
    .Q_N(_1976_),
    .Q(\systolic_array.genblk1[4].out_queue_dlygate[14].A ));
 sg13g2_dfrbp_1 _4354_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net397),
    .D(_0053_),
    .Q_N(_1977_),
    .Q(\systolic_array.genblk1[4].out_queue_dlygate[15].A ));
 sg13g2_dfrbp_1 _4355_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net398),
    .D(net877),
    .Q_N(_1978_),
    .Q(\systolic_array.genblk1[4].out_queue_dlygate[16].A ));
 sg13g2_dfrbp_1 _4356_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net399),
    .D(_0063_),
    .Q_N(_1979_),
    .Q(\systolic_array.genblk1[5].out_queue_dlygate[9].A ));
 sg13g2_dfrbp_1 _4357_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net400),
    .D(_0056_),
    .Q_N(_1980_),
    .Q(\systolic_array.genblk1[5].out_queue_dlygate[10].A ));
 sg13g2_dfrbp_1 _4358_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net401),
    .D(_0057_),
    .Q_N(_1981_),
    .Q(\systolic_array.genblk1[5].out_queue_dlygate[11].A ));
 sg13g2_dfrbp_1 _4359_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net402),
    .D(_0058_),
    .Q_N(_1982_),
    .Q(\systolic_array.genblk1[5].out_queue_dlygate[12].A ));
 sg13g2_dfrbp_1 _4360_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net403),
    .D(_0059_),
    .Q_N(_1983_),
    .Q(\systolic_array.genblk1[5].out_queue_dlygate[13].A ));
 sg13g2_dfrbp_1 _4361_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net404),
    .D(_0060_),
    .Q_N(_1984_),
    .Q(\systolic_array.genblk1[5].out_queue_dlygate[14].A ));
 sg13g2_dfrbp_1 _4362_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net405),
    .D(_0061_),
    .Q_N(_1985_),
    .Q(\systolic_array.genblk1[5].out_queue_dlygate[15].A ));
 sg13g2_dfrbp_1 _4363_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net406),
    .D(_0062_),
    .Q_N(_1986_),
    .Q(\systolic_array.genblk1[5].out_queue_dlygate[16].A ));
 sg13g2_dfrbp_1 _4364_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net407),
    .D(net803),
    .Q_N(_1987_),
    .Q(\systolic_array.genblk1[2].out_queue_dlygate[9].A ));
 sg13g2_dfrbp_1 _4365_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net31),
    .D(net766),
    .Q_N(_1988_),
    .Q(\systolic_array.genblk1[2].out_queue_dlygate[10].A ));
 sg13g2_dfrbp_1 _4366_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net32),
    .D(net723),
    .Q_N(_1989_),
    .Q(\systolic_array.genblk1[2].out_queue_dlygate[11].A ));
 sg13g2_dfrbp_1 _4367_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net33),
    .D(_0034_),
    .Q_N(_1990_),
    .Q(\systolic_array.genblk1[2].out_queue_dlygate[12].A ));
 sg13g2_dfrbp_1 _4368_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net34),
    .D(net764),
    .Q_N(_1991_),
    .Q(\systolic_array.genblk1[2].out_queue_dlygate[13].A ));
 sg13g2_dfrbp_1 _4369_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net35),
    .D(net864),
    .Q_N(_1992_),
    .Q(\systolic_array.genblk1[2].out_queue_dlygate[14].A ));
 sg13g2_dfrbp_1 _4370_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net36),
    .D(net862),
    .Q_N(_1993_),
    .Q(\systolic_array.genblk1[2].out_queue_dlygate[15].A ));
 sg13g2_dfrbp_1 _4371_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net37),
    .D(net745),
    .Q_N(_1994_),
    .Q(\systolic_array.genblk1[2].out_queue_dlygate[16].A ));
 sg13g2_dfrbp_1 _4372_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net38),
    .D(_0047_),
    .Q_N(_1995_),
    .Q(\systolic_array.genblk1[3].out_queue_dlygate[9].A ));
 sg13g2_dfrbp_1 _4373_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net39),
    .D(_0040_),
    .Q_N(_1996_),
    .Q(\systolic_array.genblk1[3].out_queue_dlygate[10].A ));
 sg13g2_dfrbp_1 _4374_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net40),
    .D(_0041_),
    .Q_N(_1997_),
    .Q(\systolic_array.genblk1[3].out_queue_dlygate[11].A ));
 sg13g2_dfrbp_1 _4375_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net41),
    .D(_0042_),
    .Q_N(_1998_),
    .Q(\systolic_array.genblk1[3].out_queue_dlygate[12].A ));
 sg13g2_dfrbp_1 _4376_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net42),
    .D(_0043_),
    .Q_N(_1999_),
    .Q(\systolic_array.genblk1[3].out_queue_dlygate[13].A ));
 sg13g2_dfrbp_1 _4377_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net43),
    .D(_0044_),
    .Q_N(_2000_),
    .Q(\systolic_array.genblk1[3].out_queue_dlygate[14].A ));
 sg13g2_dfrbp_1 _4378_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net44),
    .D(_0045_),
    .Q_N(_2001_),
    .Q(\systolic_array.genblk1[3].out_queue_dlygate[15].A ));
 sg13g2_dfrbp_1 _4379_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net45),
    .D(_0046_),
    .Q_N(_2002_),
    .Q(\systolic_array.genblk1[3].out_queue_dlygate[16].A ));
 sg13g2_dfrbp_1 _4380_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net46),
    .D(net522),
    .Q_N(_2003_),
    .Q(\systolic_array.genblk1[0].out_queue_dlygate[9].A ));
 sg13g2_dfrbp_1 _4381_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net47),
    .D(net733),
    .Q_N(_2004_),
    .Q(\systolic_array.genblk1[0].out_queue_dlygate[10].A ));
 sg13g2_dfrbp_1 _4382_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net48),
    .D(net524),
    .Q_N(_2005_),
    .Q(\systolic_array.genblk1[0].out_queue_dlygate[11].A ));
 sg13g2_dfrbp_1 _4383_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net49),
    .D(net527),
    .Q_N(_2006_),
    .Q(\systolic_array.genblk1[0].out_queue_dlygate[12].A ));
 sg13g2_dfrbp_1 _4384_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net50),
    .D(net735),
    .Q_N(_2007_),
    .Q(\systolic_array.genblk1[0].out_queue_dlygate[13].A ));
 sg13g2_dfrbp_1 _4385_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net51),
    .D(net529),
    .Q_N(_2008_),
    .Q(\systolic_array.genblk1[0].out_queue_dlygate[14].A ));
 sg13g2_dfrbp_1 _4386_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net52),
    .D(net843),
    .Q_N(_2009_),
    .Q(\systolic_array.genblk1[0].out_queue_dlygate[15].A ));
 sg13g2_dfrbp_1 _4387_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net53),
    .D(net786),
    .Q_N(_2010_),
    .Q(\systolic_array.genblk1[0].out_queue_dlygate[16].A ));
 sg13g2_dfrbp_1 _4388_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net54),
    .D(_0031_),
    .Q_N(_2011_),
    .Q(\systolic_array.genblk1[1].out_queue_dlygate[9].A ));
 sg13g2_dfrbp_1 _4389_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net55),
    .D(_0024_),
    .Q_N(_2012_),
    .Q(\systolic_array.genblk1[1].out_queue_dlygate[10].A ));
 sg13g2_dfrbp_1 _4390_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net56),
    .D(_0025_),
    .Q_N(_2013_),
    .Q(\systolic_array.genblk1[1].out_queue_dlygate[11].A ));
 sg13g2_dfrbp_1 _4391_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net57),
    .D(_0026_),
    .Q_N(_2014_),
    .Q(\systolic_array.genblk1[1].out_queue_dlygate[12].A ));
 sg13g2_dfrbp_1 _4392_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net58),
    .D(_0027_),
    .Q_N(_2015_),
    .Q(\systolic_array.genblk1[1].out_queue_dlygate[13].A ));
 sg13g2_dfrbp_1 _4393_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net59),
    .D(_0028_),
    .Q_N(_2016_),
    .Q(\systolic_array.genblk1[1].out_queue_dlygate[14].A ));
 sg13g2_dfrbp_1 _4394_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net61),
    .D(_0029_),
    .Q_N(_2017_),
    .Q(\systolic_array.genblk1[1].out_queue_dlygate[15].A ));
 sg13g2_dfrbp_1 _4395_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net87),
    .D(_0030_),
    .Q_N(_1680_),
    .Q(\systolic_array.genblk1[1].out_queue_dlygate[16].A ));
 sg13g2_dfrbp_1 _4396_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net86),
    .D(_0384_),
    .Q_N(_1679_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[0].A ));
 sg13g2_dfrbp_1 _4397_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net77),
    .D(_0385_),
    .Q_N(_1678_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[1].A ));
 sg13g2_dfrbp_1 _4398_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net76),
    .D(_0386_),
    .Q_N(_1677_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[2].A ));
 sg13g2_dfrbp_1 _4399_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net75),
    .D(_0387_),
    .Q_N(_1676_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[3].A ));
 sg13g2_dfrbp_1 _4400_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net74),
    .D(_0388_),
    .Q_N(_1675_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[4].A ));
 sg13g2_dfrbp_1 _4401_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net73),
    .D(_0389_),
    .Q_N(_1674_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[5].A ));
 sg13g2_dfrbp_1 _4402_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net72),
    .D(_0390_),
    .Q_N(_1673_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[6].A ));
 sg13g2_dfrbp_1 _4403_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net71),
    .D(_0391_),
    .Q_N(_1672_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[7].A ));
 sg13g2_dfrbp_1 _4404_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net70),
    .D(_0392_),
    .Q_N(_1671_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[8].A ));
 sg13g2_dfrbp_1 _4405_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net69),
    .D(_0393_),
    .Q_N(_0111_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[9].A ));
 sg13g2_dfrbp_1 _4406_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net68),
    .D(_0394_),
    .Q_N(_1670_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[10].A ));
 sg13g2_dfrbp_1 _4407_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net67),
    .D(_0395_),
    .Q_N(_0112_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[11].A ));
 sg13g2_dfrbp_1 _4408_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net66),
    .D(_0396_),
    .Q_N(_1669_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[12].A ));
 sg13g2_dfrbp_1 _4409_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net65),
    .D(_0397_),
    .Q_N(_0113_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[13].A ));
 sg13g2_dfrbp_1 _4410_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net64),
    .D(_0398_),
    .Q_N(_1668_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[14].A ));
 sg13g2_dfrbp_1 _4411_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net63),
    .D(_0399_),
    .Q_N(_1667_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[15].A ));
 sg13g2_dfrbp_1 _4412_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net62),
    .D(_0400_),
    .Q_N(_1666_),
    .Q(\systolic_array.genblk1[10].accumulators_dlygate[16].A ));
 sg13g2_tiehi _4366__32 (.L_HI(net32));
 sg13g2_tiehi _4367__33 (.L_HI(net33));
 sg13g2_tiehi _4368__34 (.L_HI(net34));
 sg13g2_tiehi _4369__35 (.L_HI(net35));
 sg13g2_tiehi _4370__36 (.L_HI(net36));
 sg13g2_tiehi _4371__37 (.L_HI(net37));
 sg13g2_tiehi _4372__38 (.L_HI(net38));
 sg13g2_tiehi _4373__39 (.L_HI(net39));
 sg13g2_tiehi _4374__40 (.L_HI(net40));
 sg13g2_tiehi _4375__41 (.L_HI(net41));
 sg13g2_tiehi _4376__42 (.L_HI(net42));
 sg13g2_tiehi _4377__43 (.L_HI(net43));
 sg13g2_tiehi _4378__44 (.L_HI(net44));
 sg13g2_tiehi _4379__45 (.L_HI(net45));
 sg13g2_tiehi _4380__46 (.L_HI(net46));
 sg13g2_tiehi _4381__47 (.L_HI(net47));
 sg13g2_tiehi _4382__48 (.L_HI(net48));
 sg13g2_tiehi _4383__49 (.L_HI(net49));
 sg13g2_tiehi _4384__50 (.L_HI(net50));
 sg13g2_tiehi _4385__51 (.L_HI(net51));
 sg13g2_tiehi _4386__52 (.L_HI(net52));
 sg13g2_tiehi _4387__53 (.L_HI(net53));
 sg13g2_tiehi _4388__54 (.L_HI(net54));
 sg13g2_tiehi _4389__55 (.L_HI(net55));
 sg13g2_tiehi _4390__56 (.L_HI(net56));
 sg13g2_tiehi _4391__57 (.L_HI(net57));
 sg13g2_tiehi _4392__58 (.L_HI(net58));
 sg13g2_tiehi _4393__59 (.L_HI(net59));
 sg13g2_tiehi _4045__60 (.L_HI(net60));
 sg13g2_tiehi _4394__61 (.L_HI(net61));
 sg13g2_tiehi _4412__62 (.L_HI(net62));
 sg13g2_tiehi _4411__63 (.L_HI(net63));
 sg13g2_tiehi _4410__64 (.L_HI(net64));
 sg13g2_tiehi _4409__65 (.L_HI(net65));
 sg13g2_tiehi _4408__66 (.L_HI(net66));
 sg13g2_tiehi _4407__67 (.L_HI(net67));
 sg13g2_tiehi _4406__68 (.L_HI(net68));
 sg13g2_tiehi _4405__69 (.L_HI(net69));
 sg13g2_tiehi _4404__70 (.L_HI(net70));
 sg13g2_tiehi _4403__71 (.L_HI(net71));
 sg13g2_tiehi _4402__72 (.L_HI(net72));
 sg13g2_tiehi _4401__73 (.L_HI(net73));
 sg13g2_tiehi _4400__74 (.L_HI(net74));
 sg13g2_tiehi _4399__75 (.L_HI(net75));
 sg13g2_tiehi _4398__76 (.L_HI(net76));
 sg13g2_tiehi _4397__77 (.L_HI(net77));
 sg13g2_tiehi _4044__78 (.L_HI(net78));
 sg13g2_tiehi _4036__79 (.L_HI(net79));
 sg13g2_tiehi _4037__80 (.L_HI(net80));
 sg13g2_tiehi _4038__81 (.L_HI(net81));
 sg13g2_tiehi _4039__82 (.L_HI(net82));
 sg13g2_tiehi _4040__83 (.L_HI(net83));
 sg13g2_tiehi _4041__84 (.L_HI(net84));
 sg13g2_tiehi _4042__85 (.L_HI(net85));
 sg13g2_tiehi _4396__86 (.L_HI(net86));
 sg13g2_tiehi _4395__87 (.L_HI(net87));
 sg13g2_tiehi _4314__88 (.L_HI(net88));
 sg13g2_tiehi _4313__89 (.L_HI(net89));
 sg13g2_tiehi _4312__90 (.L_HI(net90));
 sg13g2_tiehi _4311__91 (.L_HI(net91));
 sg13g2_tiehi _4310__92 (.L_HI(net92));
 sg13g2_tiehi _4309__93 (.L_HI(net93));
 sg13g2_tiehi _4308__94 (.L_HI(net94));
 sg13g2_tiehi _4307__95 (.L_HI(net95));
 sg13g2_tiehi _4306__96 (.L_HI(net96));
 sg13g2_tiehi _4305__97 (.L_HI(net97));
 sg13g2_tiehi _4304__98 (.L_HI(net98));
 sg13g2_tiehi _4303__99 (.L_HI(net99));
 sg13g2_tiehi _4302__100 (.L_HI(net100));
 sg13g2_tiehi _4301__101 (.L_HI(net101));
 sg13g2_tiehi _4300__102 (.L_HI(net102));
 sg13g2_tiehi _4299__103 (.L_HI(net103));
 sg13g2_tiehi _4298__104 (.L_HI(net104));
 sg13g2_tiehi _4289__105 (.L_HI(net105));
 sg13g2_tiehi _4288__106 (.L_HI(net106));
 sg13g2_tiehi _4287__107 (.L_HI(net107));
 sg13g2_tiehi _4286__108 (.L_HI(net108));
 sg13g2_tiehi _4285__109 (.L_HI(net109));
 sg13g2_tiehi _4284__110 (.L_HI(net110));
 sg13g2_tiehi _4283__111 (.L_HI(net111));
 sg13g2_tiehi _4282__112 (.L_HI(net112));
 sg13g2_tiehi _4281__113 (.L_HI(net113));
 sg13g2_tiehi _4280__114 (.L_HI(net114));
 sg13g2_tiehi _4279__115 (.L_HI(net115));
 sg13g2_tiehi _4278__116 (.L_HI(net116));
 sg13g2_tiehi _4277__117 (.L_HI(net117));
 sg13g2_tiehi _4276__118 (.L_HI(net118));
 sg13g2_tiehi _4275__119 (.L_HI(net119));
 sg13g2_tiehi _4274__120 (.L_HI(net120));
 sg13g2_tiehi _4273__121 (.L_HI(net121));
 sg13g2_tiehi _4272__122 (.L_HI(net122));
 sg13g2_tiehi _4271__123 (.L_HI(net123));
 sg13g2_tiehi _4270__124 (.L_HI(net124));
 sg13g2_tiehi _4269__125 (.L_HI(net125));
 sg13g2_tiehi _4268__126 (.L_HI(net126));
 sg13g2_tiehi _4267__127 (.L_HI(net127));
 sg13g2_tiehi _4266__128 (.L_HI(net128));
 sg13g2_tiehi _4265__129 (.L_HI(net129));
 sg13g2_tiehi _4264__130 (.L_HI(net130));
 sg13g2_tiehi _4263__131 (.L_HI(net131));
 sg13g2_tiehi _4262__132 (.L_HI(net132));
 sg13g2_tiehi _4261__133 (.L_HI(net133));
 sg13g2_tiehi _4260__134 (.L_HI(net134));
 sg13g2_tiehi _4259__135 (.L_HI(net135));
 sg13g2_tiehi _4258__136 (.L_HI(net136));
 sg13g2_tiehi _4257__137 (.L_HI(net137));
 sg13g2_tiehi _4256__138 (.L_HI(net138));
 sg13g2_tiehi _4255__139 (.L_HI(net139));
 sg13g2_tiehi _4254__140 (.L_HI(net140));
 sg13g2_tiehi _4253__141 (.L_HI(net141));
 sg13g2_tiehi _4252__142 (.L_HI(net142));
 sg13g2_tiehi _4251__143 (.L_HI(net143));
 sg13g2_tiehi _4250__144 (.L_HI(net144));
 sg13g2_tiehi _4249__145 (.L_HI(net145));
 sg13g2_tiehi _4248__146 (.L_HI(net146));
 sg13g2_tiehi _4247__147 (.L_HI(net147));
 sg13g2_tiehi _4246__148 (.L_HI(net148));
 sg13g2_tiehi _4245__149 (.L_HI(net149));
 sg13g2_tiehi _4244__150 (.L_HI(net150));
 sg13g2_tiehi _4243__151 (.L_HI(net151));
 sg13g2_tiehi _4242__152 (.L_HI(net152));
 sg13g2_tiehi _4241__153 (.L_HI(net153));
 sg13g2_tiehi _4240__154 (.L_HI(net154));
 sg13g2_tiehi _4239__155 (.L_HI(net155));
 sg13g2_tiehi _4238__156 (.L_HI(net156));
 sg13g2_tiehi _4237__157 (.L_HI(net157));
 sg13g2_tiehi _4236__158 (.L_HI(net158));
 sg13g2_tiehi _4235__159 (.L_HI(net159));
 sg13g2_tiehi _4234__160 (.L_HI(net160));
 sg13g2_tiehi _4233__161 (.L_HI(net161));
 sg13g2_tiehi _4232__162 (.L_HI(net162));
 sg13g2_tiehi _4231__163 (.L_HI(net163));
 sg13g2_tiehi _4230__164 (.L_HI(net164));
 sg13g2_tiehi _4229__165 (.L_HI(net165));
 sg13g2_tiehi _4228__166 (.L_HI(net166));
 sg13g2_tiehi _4227__167 (.L_HI(net167));
 sg13g2_tiehi _4226__168 (.L_HI(net168));
 sg13g2_tiehi _4225__169 (.L_HI(net169));
 sg13g2_tiehi _4224__170 (.L_HI(net170));
 sg13g2_tiehi _4223__171 (.L_HI(net171));
 sg13g2_tiehi _4222__172 (.L_HI(net172));
 sg13g2_tiehi _4221__173 (.L_HI(net173));
 sg13g2_tiehi _4220__174 (.L_HI(net174));
 sg13g2_tiehi _4219__175 (.L_HI(net175));
 sg13g2_tiehi _4218__176 (.L_HI(net176));
 sg13g2_tiehi _4217__177 (.L_HI(net177));
 sg13g2_tiehi _4216__178 (.L_HI(net178));
 sg13g2_tiehi _4215__179 (.L_HI(net179));
 sg13g2_tiehi _4214__180 (.L_HI(net180));
 sg13g2_tiehi _4213__181 (.L_HI(net181));
 sg13g2_tiehi _4212__182 (.L_HI(net182));
 sg13g2_tiehi _4211__183 (.L_HI(net183));
 sg13g2_tiehi _4210__184 (.L_HI(net184));
 sg13g2_tiehi _4209__185 (.L_HI(net185));
 sg13g2_tiehi _4208__186 (.L_HI(net186));
 sg13g2_tiehi _4207__187 (.L_HI(net187));
 sg13g2_tiehi _4206__188 (.L_HI(net188));
 sg13g2_tiehi _4205__189 (.L_HI(net189));
 sg13g2_tiehi _4204__190 (.L_HI(net190));
 sg13g2_tiehi _4203__191 (.L_HI(net191));
 sg13g2_tiehi _4202__192 (.L_HI(net192));
 sg13g2_tiehi _4201__193 (.L_HI(net193));
 sg13g2_tiehi _4200__194 (.L_HI(net194));
 sg13g2_tiehi _4199__195 (.L_HI(net195));
 sg13g2_tiehi _4198__196 (.L_HI(net196));
 sg13g2_tiehi _4197__197 (.L_HI(net197));
 sg13g2_tiehi _4196__198 (.L_HI(net198));
 sg13g2_tiehi _4195__199 (.L_HI(net199));
 sg13g2_tiehi _4194__200 (.L_HI(net200));
 sg13g2_tiehi _4193__201 (.L_HI(net201));
 sg13g2_tiehi _4192__202 (.L_HI(net202));
 sg13g2_tiehi _4191__203 (.L_HI(net203));
 sg13g2_tiehi _4190__204 (.L_HI(net204));
 sg13g2_tiehi _4189__205 (.L_HI(net205));
 sg13g2_tiehi _4188__206 (.L_HI(net206));
 sg13g2_tiehi _4187__207 (.L_HI(net207));
 sg13g2_tiehi _4186__208 (.L_HI(net208));
 sg13g2_tiehi _4185__209 (.L_HI(net209));
 sg13g2_tiehi _4184__210 (.L_HI(net210));
 sg13g2_tiehi _4183__211 (.L_HI(net211));
 sg13g2_tiehi _4182__212 (.L_HI(net212));
 sg13g2_tiehi _4181__213 (.L_HI(net213));
 sg13g2_tiehi _4180__214 (.L_HI(net214));
 sg13g2_tiehi _4179__215 (.L_HI(net215));
 sg13g2_tiehi _4178__216 (.L_HI(net216));
 sg13g2_tiehi _4177__217 (.L_HI(net217));
 sg13g2_tiehi _4176__218 (.L_HI(net218));
 sg13g2_tiehi _4175__219 (.L_HI(net219));
 sg13g2_tiehi _4174__220 (.L_HI(net220));
 sg13g2_tiehi _4173__221 (.L_HI(net221));
 sg13g2_tiehi _4172__222 (.L_HI(net222));
 sg13g2_tiehi _4171__223 (.L_HI(net223));
 sg13g2_tiehi _4170__224 (.L_HI(net224));
 sg13g2_tiehi _4169__225 (.L_HI(net225));
 sg13g2_tiehi _4168__226 (.L_HI(net226));
 sg13g2_tiehi _4167__227 (.L_HI(net227));
 sg13g2_tiehi _4166__228 (.L_HI(net228));
 sg13g2_tiehi _4165__229 (.L_HI(net229));
 sg13g2_tiehi _4164__230 (.L_HI(net230));
 sg13g2_tiehi _4163__231 (.L_HI(net231));
 sg13g2_tiehi _4162__232 (.L_HI(net232));
 sg13g2_tiehi _4161__233 (.L_HI(net233));
 sg13g2_tiehi _4160__234 (.L_HI(net234));
 sg13g2_tiehi _4159__235 (.L_HI(net235));
 sg13g2_tiehi _4158__236 (.L_HI(net236));
 sg13g2_tiehi _4157__237 (.L_HI(net237));
 sg13g2_tiehi _4156__238 (.L_HI(net238));
 sg13g2_tiehi _4155__239 (.L_HI(net239));
 sg13g2_tiehi _4154__240 (.L_HI(net240));
 sg13g2_tiehi _4153__241 (.L_HI(net241));
 sg13g2_tiehi _4152__242 (.L_HI(net242));
 sg13g2_tiehi _4151__243 (.L_HI(net243));
 sg13g2_tiehi _4150__244 (.L_HI(net244));
 sg13g2_tiehi _4149__245 (.L_HI(net245));
 sg13g2_tiehi _4148__246 (.L_HI(net246));
 sg13g2_tiehi _4147__247 (.L_HI(net247));
 sg13g2_tiehi _4146__248 (.L_HI(net248));
 sg13g2_tiehi _4145__249 (.L_HI(net249));
 sg13g2_tiehi _4144__250 (.L_HI(net250));
 sg13g2_tiehi _4143__251 (.L_HI(net251));
 sg13g2_tiehi _4142__252 (.L_HI(net252));
 sg13g2_tiehi _4141__253 (.L_HI(net253));
 sg13g2_tiehi _4140__254 (.L_HI(net254));
 sg13g2_tiehi _4139__255 (.L_HI(net255));
 sg13g2_tiehi _4138__256 (.L_HI(net256));
 sg13g2_tiehi _4137__257 (.L_HI(net257));
 sg13g2_tiehi _4136__258 (.L_HI(net258));
 sg13g2_tiehi _4135__259 (.L_HI(net259));
 sg13g2_tiehi _4134__260 (.L_HI(net260));
 sg13g2_tiehi _4133__261 (.L_HI(net261));
 sg13g2_tiehi _4132__262 (.L_HI(net262));
 sg13g2_tiehi _4131__263 (.L_HI(net263));
 sg13g2_tiehi _4130__264 (.L_HI(net264));
 sg13g2_tiehi _4129__265 (.L_HI(net265));
 sg13g2_tiehi _4128__266 (.L_HI(net266));
 sg13g2_tiehi _4127__267 (.L_HI(net267));
 sg13g2_tiehi _4126__268 (.L_HI(net268));
 sg13g2_tiehi _4125__269 (.L_HI(net269));
 sg13g2_tiehi _4124__270 (.L_HI(net270));
 sg13g2_tiehi _4123__271 (.L_HI(net271));
 sg13g2_tiehi _4122__272 (.L_HI(net272));
 sg13g2_tiehi _4121__273 (.L_HI(net273));
 sg13g2_tiehi _4120__274 (.L_HI(net274));
 sg13g2_tiehi _4119__275 (.L_HI(net275));
 sg13g2_tiehi _4118__276 (.L_HI(net276));
 sg13g2_tiehi _4117__277 (.L_HI(net277));
 sg13g2_tiehi _4116__278 (.L_HI(net278));
 sg13g2_tiehi _4115__279 (.L_HI(net279));
 sg13g2_tiehi _4114__280 (.L_HI(net280));
 sg13g2_tiehi _4113__281 (.L_HI(net281));
 sg13g2_tiehi _4112__282 (.L_HI(net282));
 sg13g2_tiehi _4111__283 (.L_HI(net283));
 sg13g2_tiehi _4110__284 (.L_HI(net284));
 sg13g2_tiehi _4109__285 (.L_HI(net285));
 sg13g2_tiehi _4108__286 (.L_HI(net286));
 sg13g2_tiehi _4107__287 (.L_HI(net287));
 sg13g2_tiehi _4106__288 (.L_HI(net288));
 sg13g2_tiehi _4105__289 (.L_HI(net289));
 sg13g2_tiehi _4104__290 (.L_HI(net290));
 sg13g2_tiehi _4103__291 (.L_HI(net291));
 sg13g2_tiehi _4102__292 (.L_HI(net292));
 sg13g2_tiehi _4101__293 (.L_HI(net293));
 sg13g2_tiehi _4100__294 (.L_HI(net294));
 sg13g2_tiehi _4099__295 (.L_HI(net295));
 sg13g2_tiehi _4098__296 (.L_HI(net296));
 sg13g2_tiehi _4097__297 (.L_HI(net297));
 sg13g2_tiehi _4096__298 (.L_HI(net298));
 sg13g2_tiehi _4095__299 (.L_HI(net299));
 sg13g2_tiehi _4094__300 (.L_HI(net300));
 sg13g2_tiehi _4093__301 (.L_HI(net301));
 sg13g2_tiehi _4092__302 (.L_HI(net302));
 sg13g2_tiehi _4091__303 (.L_HI(net303));
 sg13g2_tiehi _4090__304 (.L_HI(net304));
 sg13g2_tiehi _4089__305 (.L_HI(net305));
 sg13g2_tiehi _4088__306 (.L_HI(net306));
 sg13g2_tiehi _4087__307 (.L_HI(net307));
 sg13g2_tiehi _4086__308 (.L_HI(net308));
 sg13g2_tiehi _4085__309 (.L_HI(net309));
 sg13g2_tiehi _4084__310 (.L_HI(net310));
 sg13g2_tiehi _4083__311 (.L_HI(net311));
 sg13g2_tiehi _4082__312 (.L_HI(net312));
 sg13g2_tiehi _4081__313 (.L_HI(net313));
 sg13g2_tiehi _4080__314 (.L_HI(net314));
 sg13g2_tiehi _4079__315 (.L_HI(net315));
 sg13g2_tiehi _4078__316 (.L_HI(net316));
 sg13g2_tiehi _4077__317 (.L_HI(net317));
 sg13g2_tiehi _4076__318 (.L_HI(net318));
 sg13g2_tiehi _4075__319 (.L_HI(net319));
 sg13g2_tiehi _4074__320 (.L_HI(net320));
 sg13g2_tiehi _4073__321 (.L_HI(net321));
 sg13g2_tiehi _4072__322 (.L_HI(net322));
 sg13g2_tiehi _4071__323 (.L_HI(net323));
 sg13g2_tiehi _4070__324 (.L_HI(net324));
 sg13g2_tiehi _4069__325 (.L_HI(net325));
 sg13g2_tiehi _4068__326 (.L_HI(net326));
 sg13g2_tiehi _4067__327 (.L_HI(net327));
 sg13g2_tiehi _4066__328 (.L_HI(net328));
 sg13g2_tiehi _4065__329 (.L_HI(net329));
 sg13g2_tiehi _4064__330 (.L_HI(net330));
 sg13g2_tiehi _4063__331 (.L_HI(net331));
 sg13g2_tiehi _4043__332 (.L_HI(net332));
 sg13g2_tiehi _4290__333 (.L_HI(net333));
 sg13g2_tiehi _4291__334 (.L_HI(net334));
 sg13g2_tiehi _4292__335 (.L_HI(net335));
 sg13g2_tiehi _4293__336 (.L_HI(net336));
 sg13g2_tiehi _4294__337 (.L_HI(net337));
 sg13g2_tiehi _4295__338 (.L_HI(net338));
 sg13g2_tiehi _4296__339 (.L_HI(net339));
 sg13g2_tiehi _4062__340 (.L_HI(net340));
 sg13g2_tiehi _4061__341 (.L_HI(net341));
 sg13g2_tiehi _4060__342 (.L_HI(net342));
 sg13g2_tiehi _4059__343 (.L_HI(net343));
 sg13g2_tiehi _4058__344 (.L_HI(net344));
 sg13g2_tiehi _4057__345 (.L_HI(net345));
 sg13g2_tiehi _4056__346 (.L_HI(net346));
 sg13g2_tiehi _4055__347 (.L_HI(net347));
 sg13g2_tiehi _4054__348 (.L_HI(net348));
 sg13g2_tiehi _4053__349 (.L_HI(net349));
 sg13g2_tiehi _4052__350 (.L_HI(net350));
 sg13g2_tiehi _4051__351 (.L_HI(net351));
 sg13g2_tiehi _4050__352 (.L_HI(net352));
 sg13g2_tiehi _4049__353 (.L_HI(net353));
 sg13g2_tiehi _4048__354 (.L_HI(net354));
 sg13g2_tiehi _4047__355 (.L_HI(net355));
 sg13g2_tiehi _4046__356 (.L_HI(net356));
 sg13g2_tiehi _4297__357 (.L_HI(net357));
 sg13g2_tiehi _4315__358 (.L_HI(net358));
 sg13g2_tiehi _4316__359 (.L_HI(net359));
 sg13g2_tiehi _4317__360 (.L_HI(net360));
 sg13g2_tiehi _4318__361 (.L_HI(net361));
 sg13g2_tiehi _4319__362 (.L_HI(net362));
 sg13g2_tiehi _4320__363 (.L_HI(net363));
 sg13g2_tiehi _4321__364 (.L_HI(net364));
 sg13g2_tiehi _4322__365 (.L_HI(net365));
 sg13g2_tiehi _4323__366 (.L_HI(net366));
 sg13g2_tiehi _4324__367 (.L_HI(net367));
 sg13g2_tiehi _4325__368 (.L_HI(net368));
 sg13g2_tiehi _4326__369 (.L_HI(net369));
 sg13g2_tiehi _4327__370 (.L_HI(net370));
 sg13g2_tiehi _4328__371 (.L_HI(net371));
 sg13g2_tiehi _4329__372 (.L_HI(net372));
 sg13g2_tiehi _4330__373 (.L_HI(net373));
 sg13g2_tiehi _4331__374 (.L_HI(net374));
 sg13g2_tiehi _4332__375 (.L_HI(net375));
 sg13g2_tiehi _4333__376 (.L_HI(net376));
 sg13g2_tiehi _4334__377 (.L_HI(net377));
 sg13g2_tiehi _4335__378 (.L_HI(net378));
 sg13g2_tiehi _4336__379 (.L_HI(net379));
 sg13g2_tiehi _4337__380 (.L_HI(net380));
 sg13g2_tiehi _4338__381 (.L_HI(net381));
 sg13g2_tiehi _4339__382 (.L_HI(net382));
 sg13g2_tiehi _4340__383 (.L_HI(net383));
 sg13g2_tiehi _4341__384 (.L_HI(net384));
 sg13g2_tiehi _4342__385 (.L_HI(net385));
 sg13g2_tiehi _4343__386 (.L_HI(net386));
 sg13g2_tiehi _4344__387 (.L_HI(net387));
 sg13g2_tiehi _4345__388 (.L_HI(net388));
 sg13g2_tiehi _4346__389 (.L_HI(net389));
 sg13g2_tiehi _4347__390 (.L_HI(net390));
 sg13g2_tiehi _4348__391 (.L_HI(net391));
 sg13g2_tiehi _4349__392 (.L_HI(net392));
 sg13g2_tiehi _4350__393 (.L_HI(net393));
 sg13g2_tiehi _4351__394 (.L_HI(net394));
 sg13g2_tiehi _4352__395 (.L_HI(net395));
 sg13g2_tiehi _4353__396 (.L_HI(net396));
 sg13g2_tiehi _4354__397 (.L_HI(net397));
 sg13g2_tiehi _4355__398 (.L_HI(net398));
 sg13g2_tiehi _4356__399 (.L_HI(net399));
 sg13g2_tiehi _4357__400 (.L_HI(net400));
 sg13g2_tiehi _4358__401 (.L_HI(net401));
 sg13g2_tiehi _4359__402 (.L_HI(net402));
 sg13g2_tiehi _4360__403 (.L_HI(net403));
 sg13g2_tiehi _4361__404 (.L_HI(net404));
 sg13g2_tiehi _4362__405 (.L_HI(net405));
 sg13g2_tiehi _4363__406 (.L_HI(net406));
 sg13g2_tiehi _4364__407 (.L_HI(net407));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_rejunity_e2m0_x_i8_matmul_16 (.L_LO(net16));
 sg13g2_tielo tt_um_rejunity_e2m0_x_i8_matmul_17 (.L_LO(net17));
 sg13g2_tielo tt_um_rejunity_e2m0_x_i8_matmul_18 (.L_LO(net18));
 sg13g2_tielo tt_um_rejunity_e2m0_x_i8_matmul_19 (.L_LO(net19));
 sg13g2_tielo tt_um_rejunity_e2m0_x_i8_matmul_20 (.L_LO(net20));
 sg13g2_tielo tt_um_rejunity_e2m0_x_i8_matmul_21 (.L_LO(net21));
 sg13g2_tielo tt_um_rejunity_e2m0_x_i8_matmul_22 (.L_LO(net22));
 sg13g2_tielo tt_um_rejunity_e2m0_x_i8_matmul_23 (.L_LO(net23));
 sg13g2_tielo tt_um_rejunity_e2m0_x_i8_matmul_24 (.L_LO(net24));
 sg13g2_tielo tt_um_rejunity_e2m0_x_i8_matmul_25 (.L_LO(net25));
 sg13g2_tielo tt_um_rejunity_e2m0_x_i8_matmul_26 (.L_LO(net26));
 sg13g2_tielo tt_um_rejunity_e2m0_x_i8_matmul_27 (.L_LO(net27));
 sg13g2_tielo tt_um_rejunity_e2m0_x_i8_matmul_28 (.L_LO(net28));
 sg13g2_tielo tt_um_rejunity_e2m0_x_i8_matmul_29 (.L_LO(net29));
 sg13g2_tielo tt_um_rejunity_e2m0_x_i8_matmul_30 (.L_LO(net30));
 sg13g2_tiehi _4365__31 (.L_HI(net31));
 sg13g2_buf_1 _4806_ (.A(\systolic_array.genblk1[0].out_queue_dlygate[9].A ),
    .X(uo_out[0]));
 sg13g2_buf_2 _4807_ (.A(\systolic_array.genblk1[0].out_queue_dlygate[10].A ),
    .X(uo_out[1]));
 sg13g2_buf_1 _4808_ (.A(\systolic_array.genblk1[0].out_queue_dlygate[11].A ),
    .X(uo_out[2]));
 sg13g2_buf_1 _4809_ (.A(\systolic_array.genblk1[0].out_queue_dlygate[12].A ),
    .X(uo_out[3]));
 sg13g2_buf_1 _4810_ (.A(\systolic_array.genblk1[0].out_queue_dlygate[13].A ),
    .X(uo_out[4]));
 sg13g2_buf_1 _4811_ (.A(\systolic_array.genblk1[0].out_queue_dlygate[14].A ),
    .X(uo_out[5]));
 sg13g2_buf_1 _4812_ (.A(\systolic_array.genblk1[0].out_queue_dlygate[15].A ),
    .X(uo_out[6]));
 sg13g2_buf_1 _4813_ (.A(\systolic_array.genblk1[0].out_queue_dlygate[16].A ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout545 (.A(_0865_),
    .X(net545));
 sg13g2_buf_1 fanout546 (.A(_0865_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(net548),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(net549),
    .X(net548));
 sg13g2_buf_1 fanout549 (.A(_0721_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(net551),
    .X(net550));
 sg13g2_buf_4 fanout551 (.X(net551),
    .A(_0455_));
 sg13g2_buf_2 fanout552 (.A(net553),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(net554),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(_1000_),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(net556),
    .X(net555));
 sg13g2_buf_1 fanout556 (.A(net557),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_0580_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(net559),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_1574_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(net562),
    .X(net560));
 sg13g2_buf_1 fanout561 (.A(net562),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(net563),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(net564),
    .X(net563));
 sg13g2_buf_8 fanout564 (.A(_1310_),
    .X(net564));
 sg13g2_buf_4 fanout565 (.X(net565),
    .A(net566));
 sg13g2_buf_4 fanout566 (.X(net566),
    .A(_1310_));
 sg13g2_buf_2 fanout567 (.A(net569),
    .X(net567));
 sg13g2_buf_1 fanout568 (.A(net569),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(net581),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(net581),
    .X(net570));
 sg13g2_buf_1 fanout571 (.A(net581),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(net573),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(net580),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(net580),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(net580),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(net579),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(net579),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(net579),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(net580),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(net581),
    .X(net580));
 sg13g2_buf_4 fanout581 (.X(net581),
    .A(_1309_));
 sg13g2_buf_2 fanout582 (.A(net585),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(net585),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(net585),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(net595),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(net590),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(net590),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(net590),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(net590),
    .X(net589));
 sg13g2_buf_1 fanout590 (.A(net595),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(net592),
    .X(net591));
 sg13g2_buf_1 fanout592 (.A(net594),
    .X(net592));
 sg13g2_buf_4 fanout593 (.X(net593),
    .A(net594));
 sg13g2_buf_4 fanout594 (.X(net594),
    .A(net595));
 sg13g2_buf_2 fanout595 (.A(_1309_),
    .X(net595));
 sg13g2_buf_4 fanout596 (.X(net596),
    .A(net597));
 sg13g2_buf_2 fanout597 (.A(net600),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(net600),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(net600),
    .X(net599));
 sg13g2_buf_4 fanout600 (.X(net600),
    .A(_1542_));
 sg13g2_buf_4 fanout601 (.X(net601),
    .A(net602));
 sg13g2_buf_4 fanout602 (.X(net602),
    .A(net605));
 sg13g2_buf_4 fanout603 (.X(net603),
    .A(net604));
 sg13g2_buf_4 fanout604 (.X(net604),
    .A(net605));
 sg13g2_buf_2 fanout605 (.A(_1542_),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(net607),
    .X(net606));
 sg13g2_buf_4 fanout607 (.X(net607),
    .A(net609));
 sg13g2_buf_4 fanout608 (.X(net608),
    .A(net609));
 sg13g2_buf_2 fanout609 (.A(net612),
    .X(net609));
 sg13g2_buf_4 fanout610 (.X(net610),
    .A(net612));
 sg13g2_buf_2 fanout611 (.A(net612),
    .X(net611));
 sg13g2_buf_4 fanout612 (.X(net612),
    .A(_1541_));
 sg13g2_buf_4 fanout613 (.X(net613),
    .A(net614));
 sg13g2_buf_4 fanout614 (.X(net614),
    .A(net615));
 sg13g2_buf_4 fanout615 (.X(net615),
    .A(_1541_));
 sg13g2_buf_2 fanout616 (.A(net618),
    .X(net616));
 sg13g2_buf_1 fanout617 (.A(net618),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_1521_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_1514_),
    .X(net619));
 sg13g2_buf_1 fanout620 (.A(_1514_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_1514_),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(net623),
    .X(net622));
 sg13g2_buf_1 fanout623 (.A(net624),
    .X(net623));
 sg13g2_buf_4 fanout624 (.X(net624),
    .A(_1506_));
 sg13g2_buf_2 fanout625 (.A(net626),
    .X(net625));
 sg13g2_buf_4 fanout626 (.X(net626),
    .A(_1498_));
 sg13g2_buf_4 fanout627 (.X(net627),
    .A(_1489_));
 sg13g2_buf_2 fanout628 (.A(_1489_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(net630),
    .X(net629));
 sg13g2_buf_4 fanout630 (.X(net630),
    .A(_1477_));
 sg13g2_buf_2 fanout631 (.A(net632),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(\systolic_array.genblk2[0].mac[4].div2 ),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(\systolic_array.genblk2[0].mac[3].div2 ),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(net635),
    .X(net634));
 sg13g2_buf_1 fanout635 (.A(\systolic_array.genblk2[0].mac[1].div2 ),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(\systolic_array.genblk2[0].mac[0].div2 ),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(net638),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(net646),
    .X(net638));
 sg13g2_buf_4 fanout639 (.X(net639),
    .A(net642));
 sg13g2_buf_2 fanout640 (.A(net642),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(net642),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(net646),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(net644),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(net645),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(net646),
    .X(net645));
 sg13g2_buf_4 fanout646 (.X(net646),
    .A(net841));
 sg13g2_buf_2 fanout647 (.A(net648),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(net649),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(\systolic_array.genblk2[0].mac[5].zero ),
    .X(net649));
 sg13g2_buf_4 fanout650 (.X(net650),
    .A(\systolic_array.genblk2[0].mac[4].zero ));
 sg13g2_buf_2 fanout651 (.A(net652),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(\systolic_array.genblk2[0].mac[3].zero ),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(net654),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(net655),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(\systolic_array.genblk2[0].mac[2].zero ),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(net658),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(net658),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(\systolic_array.genblk2[0].mac[1].zero ),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(net660),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(\systolic_array.genblk2[0].mac[0].zero ),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(\systolic_array.genblk2[0].mac[5].sign ),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(\systolic_array.genblk2[0].mac[1].sign ),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(\systolic_array.genblk2[0].mac[5].mul2 ),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(net886),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(net666),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(\systolic_array.genblk2[0].mac[4].mul2 ),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(\systolic_array.genblk2[0].mac[3].mul2 ),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(\systolic_array.genblk2[0].mac[3].mul2 ),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(net670),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(\systolic_array.genblk2[0].mac[2].mul2 ),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_1 fanout672 (.A(net673),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(\systolic_array.genblk2[0].mac[1].mul2 ),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(net676),
    .X(net674));
 sg13g2_buf_1 fanout675 (.A(net676),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(\systolic_array.genblk2[0].mac[0].mul2 ),
    .X(net676));
 sg13g2_buf_4 fanout677 (.X(net677),
    .A(\systolic_array.arg_top_curr[7] ));
 sg13g2_buf_2 fanout678 (.A(\systolic_array.arg_top_curr[7] ),
    .X(net678));
 sg13g2_buf_4 fanout679 (.X(net679),
    .A(\systolic_array.arg_top_curr[5] ));
 sg13g2_buf_2 fanout680 (.A(\systolic_array.arg_top_curr[5] ),
    .X(net680));
 sg13g2_buf_4 fanout681 (.X(net681),
    .A(\systolic_array.arg_top_curr[4] ));
 sg13g2_buf_2 fanout682 (.A(net684),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(net684),
    .X(net683));
 sg13g2_buf_4 fanout684 (.X(net684),
    .A(\systolic_array.arg_top_curr[3] ));
 sg13g2_buf_2 fanout685 (.A(net687),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(\systolic_array.arg_top_curr[2] ),
    .X(net687));
 sg13g2_buf_4 fanout688 (.X(net688),
    .A(net690));
 sg13g2_buf_2 fanout689 (.A(net690),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(\systolic_array.arg_top_curr[1] ),
    .X(net690));
 sg13g2_buf_4 fanout691 (.X(net691),
    .A(net692));
 sg13g2_buf_4 fanout692 (.X(net692),
    .A(\systolic_array.arg_top_curr[0] ));
 sg13g2_buf_2 fanout693 (.A(_1150_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_1464_),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(_1462_),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(net6),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(net699),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(net700),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(ui_in[6]),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(net703),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(net703),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(ui_in[5]),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(net706),
    .X(net704));
 sg13g2_buf_1 fanout705 (.A(net706),
    .X(net705));
 sg13g2_buf_1 fanout706 (.A(net5),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(net5),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(net709),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(net710),
    .X(net709));
 sg13g2_buf_2 fanout710 (.A(net4),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(net3),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(net2),
    .X(net712));
 sg13g2_buf_4 fanout713 (.X(net713),
    .A(net714));
 sg13g2_buf_2 fanout714 (.A(ui_in[0]),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(rst_n),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(rst_n),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(net718),
    .X(net717));
 sg13g2_buf_1 fanout718 (.A(net720),
    .X(net718));
 sg13g2_buf_4 fanout719 (.X(net719),
    .A(net720));
 sg13g2_buf_2 fanout720 (.A(rst_n),
    .X(net720));
 sg13g2_buf_4 input1 (.X(net1),
    .A(ena));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[7]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[0]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[1]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[4]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[5]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[6]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[7]),
    .X(net14));
 sg13g2_tielo tt_um_rejunity_e2m0_x_i8_matmul_15 (.L_LO(net15));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_48_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_34_clk));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_35_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_38_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_31_clk));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_11_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_15_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_29_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_30_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_1665_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold2 (.A(\systolic_array.genblk1[9].accumulators_dlygate[5].A ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold3 (.A(\systolic_array.genblk1[9].accumulators_dlygate[9].A ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold4 (.A(\systolic_array.genblk1[9].accumulators_dlygate[8].A ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold5 (.A(\systolic_array.genblk1[9].accumulators_dlygate[0].A ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold6 (.A(\systolic_array.genblk1[7].accumulators_dlygate[2].A ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold7 (.A(\systolic_array.genblk1[3].accumulators_dlygate[0].A ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold8 (.A(\systolic_array.genblk1[1].accumulators_dlygate[8].A ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold9 (.A(\systolic_array.genblk1[3].accumulators_dlygate[6].A ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold10 (.A(\systolic_array.genblk1[5].accumulators_dlygate[5].A ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold11 (.A(\systolic_array.genblk1[5].accumulators_dlygate[10].A ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold12 (.A(\systolic_array.genblk1[3].accumulators_dlygate[7].A ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold13 (.A(\systolic_array.genblk1[11].accumulators_dlygate[7].A ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold14 (.A(\systolic_array.genblk1[9].accumulators_dlygate[2].A ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold15 (.A(\systolic_array.genblk1[3].accumulators_dlygate[5].A ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold16 (.A(\systolic_array.genblk1[11].accumulators_dlygate[1].A ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold17 (.A(\systolic_array.genblk1[9].accumulators_dlygate[16].A ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold18 (.A(\systolic_array.genblk1[9].accumulators_dlygate[3].A ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold19 (.A(\systolic_array.genblk1[7].accumulators_dlygate[3].A ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold20 (.A(\systolic_array.genblk1[1].accumulators_dlygate[1].A ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold21 (.A(\systolic_array.genblk1[5].accumulators_dlygate[0].A ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold22 (.A(\systolic_array.genblk1[1].accumulators_dlygate[2].A ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold23 (.A(\systolic_array.genblk1[7].accumulators_dlygate[5].A ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold24 (.A(\systolic_array.genblk1[7].accumulators_dlygate[6].A ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold25 (.A(\systolic_array.genblk1[5].accumulators_dlygate[8].A ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold26 (.A(\systolic_array.arg_top_next[11] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold27 (.A(\systolic_array.genblk1[5].accumulators_dlygate[7].A ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold28 (.A(\systolic_array.genblk1[7].accumulators_dlygate[15].A ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold29 (.A(\systolic_array.genblk1[3].accumulators_dlygate[2].A ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold30 (.A(\systolic_array.genblk1[1].accumulators_dlygate[7].A ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold31 (.A(\systolic_array.genblk1[3].accumulators_dlygate[8].A ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold32 (.A(\systolic_array.genblk1[1].accumulators_dlygate[15].A ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold33 (.A(\systolic_array.genblk1[1].accumulators_dlygate[12].A ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold34 (.A(\systolic_array.genblk1[11].accumulators_dlygate[5].A ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold35 (.A(\systolic_array.arg_top_next[5] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold36 (.A(\systolic_array.genblk1[7].accumulators_dlygate[14].A ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold37 (.A(\systolic_array.genblk1[1].accumulators_dlygate[0].A ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold38 (.A(\systolic_array.genblk1[7].accumulators_dlygate[4].A ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold39 (.A(\systolic_array.genblk1[7].accumulators_dlygate[9].A ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold40 (.A(\systolic_array.genblk1[1].accumulators_dlygate[13].A ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold41 (.A(\systolic_array.genblk1[5].accumulators_dlygate[12].A ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold42 (.A(\systolic_array.genblk1[11].accumulators_dlygate[4].A ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold43 (.A(\systolic_array.genblk1[11].accumulators_dlygate[6].A ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold44 (.A(\systolic_array.genblk1[7].accumulators_dlygate[10].A ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold45 (.A(\systolic_array.genblk1[11].accumulators_dlygate[0].A ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold46 (.A(\systolic_array.genblk1[7].accumulators_dlygate[11].A ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold47 (.A(\systolic_array.genblk1[5].accumulators_dlygate[14].A ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold48 (.A(\systolic_array.genblk1[1].accumulators_dlygate[5].A ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold49 (.A(\systolic_array.genblk1[3].accumulators_dlygate[10].A ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold50 (.A(\systolic_array.genblk1[7].accumulators_dlygate[0].A ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold51 (.A(\systolic_array.genblk1[5].accumulators_dlygate[1].A ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold52 (.A(\systolic_array.genblk1[1].accumulators_dlygate[6].A ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold53 (.A(\systolic_array.genblk1[9].accumulators_dlygate[6].A ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold54 (.A(\systolic_array.arg_top_next[6] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold55 (.A(\systolic_array.genblk1[9].accumulators_dlygate[4].A ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold56 (.A(\systolic_array.genblk1[5].accumulators_dlygate[2].A ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold57 (.A(\systolic_array.genblk1[5].accumulators_dlygate[3].A ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold58 (.A(\systolic_array.genblk1[9].accumulators_dlygate[1].A ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold59 (.A(\systolic_array.genblk1[7].accumulators_dlygate[13].A ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold60 (.A(\systolic_array.genblk1[3].accumulators_dlygate[11].A ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold61 (.A(\systolic_array.genblk1[5].accumulators_dlygate[6].A ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold62 (.A(\systolic_array.genblk1[3].accumulators_dlygate[14].A ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold63 (.A(\systolic_array.genblk1[9].accumulators_dlygate[12].A ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold64 (.A(\systolic_array.arg_top_next[4] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold65 (.A(\systolic_array.genblk1[11].accumulators_dlygate[2].A ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold66 (.A(\systolic_array.arg_top_next[7] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold67 (.A(\systolic_array.genblk1[5].accumulators_dlygate[16].A ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold68 (.A(\systolic_array.genblk1[5].accumulators_dlygate[4].A ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold69 (.A(\systolic_array.genblk1[9].accumulators_dlygate[7].A ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold70 (.A(\systolic_array.arg_top_next[1] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold71 (.A(\systolic_array.genblk1[1].accumulators_dlygate[14].A ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold72 (.A(\systolic_array.genblk1[3].accumulators_dlygate[16].A ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold73 (.A(\systolic_array.genblk1[7].accumulators_dlygate[7].A ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold74 (.A(\systolic_array.genblk1[1].accumulators_dlygate[10].A ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold75 (.A(\systolic_array.arg_top_next[0] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold76 (.A(\systolic_array.arg_top_next[12] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold77 (.A(\systolic_array.genblk1[1].accumulators_dlygate[11].A ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold78 (.A(\systolic_array.genblk1[7].accumulators_dlygate[1].A ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold79 (.A(\systolic_array.genblk1[7].accumulators_dlygate[12].A ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold80 (.A(\systolic_array.genblk1[9].accumulators_dlygate[10].A ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold81 (.A(\systolic_array.genblk1[3].accumulators_dlygate[12].A ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold82 (.A(\systolic_array.genblk1[9].accumulators_dlygate[15].A ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold83 (.A(\systolic_array.genblk1[3].accumulators_dlygate[13].A ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold84 (.A(\systolic_array.genblk1[7].accumulators_dlygate[16].A ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold85 (.A(\systolic_array.genblk1[3].accumulators_dlygate[15].A ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold86 (.A(\systolic_array.genblk1[5].accumulators_dlygate[11].A ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold87 (.A(\systolic_array.arg_top_next[9] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold88 (.A(\systolic_array.genblk1[11].accumulators_dlygate[8].A ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold89 (.A(\systolic_array.genblk1[5].accumulators_dlygate[13].A ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold90 (.A(\systolic_array.arg_top_next[15] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold91 (.A(\systolic_array.genblk1[3].accumulators_dlygate[9].A ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold92 (.A(\systolic_array.genblk1[5].accumulators_dlygate[15].A ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold93 (.A(\systolic_array.arg_top_next[2] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold94 (.A(\systolic_array.genblk1[1].accumulators_dlygate[4].A ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold95 (.A(\systolic_array.genblk1[9].accumulators_dlygate[14].A ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold96 (.A(\systolic_array.genblk1[9].accumulators_dlygate[11].A ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold97 (.A(\systolic_array.arg_left_div2_next[1] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0364_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold99 (.A(\systolic_array.genblk1[11].accumulators_dlygate[3].A ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold100 (.A(\systolic_array.genblk1[9].accumulators_dlygate[13].A ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold101 (.A(\systolic_array.genblk1[1].accumulators_dlygate[9].A ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold102 (.A(\systolic_array.genblk1[5].accumulators_dlygate[9].A ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold103 (.A(\systolic_array.genblk1[1].accumulators_dlygate[16].A ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold104 (.A(\systolic_array.genblk1[3].accumulators_dlygate[3].A ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold105 (.A(\systolic_array.arg_top_next[3] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0154_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold107 (.A(\systolic_array.arg_top_next[13] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold108 (.A(\systolic_array.genblk1[1].accumulators_dlygate[3].A ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold109 (.A(\systolic_array.genblk1[3].accumulators_dlygate[1].A ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold110 (.A(\systolic_array.genblk1[11].accumulators_dlygate[15].A ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold111 (.A(\systolic_array.genblk1[3].accumulators_dlygate[4].A ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold112 (.A(\systolic_array.genblk1[7].accumulators_dlygate[8].A ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold113 (.A(\systolic_array.arg_top_next[14] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold114 (.A(\systolic_array.genblk1[1].out_queue_dlygate[9].A ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0015_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold116 (.A(\systolic_array.genblk1[1].out_queue_dlygate[11].A ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0009_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold118 (.A(\systolic_array.genblk1[11].accumulators_dlygate[10].A ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold119 (.A(\systolic_array.genblk1[1].out_queue_dlygate[12].A ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0010_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold121 (.A(\systolic_array.genblk1[1].out_queue_dlygate[14].A ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0012_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold123 (.A(\systolic_array.arg_top_next[8] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold124 (.A(\systolic_array.genblk1[11].accumulators_dlygate[11].A ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold125 (.A(\systolic_array.genblk1[11].accumulators_dlygate[12].A ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold126 (.A(\systolic_array.genblk1[11].out_queue_dlygate[14].A ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0020_),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold128 (.A(\systolic_array.genblk1[11].accumulators_dlygate[16].A ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold129 (.A(\systolic_array.arg_left_sign_next[2] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0169_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold131 (.A(\systolic_array.arg_left_zero_next[2] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold132 (.A(\systolic_array.genblk1[9].out_queue_dlygate[10].A ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0080_),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold134 (.A(\systolic_array.genblk1[5].out_queue_dlygate[14].A ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0052_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold136 (.A(\systolic_array.arg_left_mul2_next[1] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0162_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold138 (.A(\systolic_array.arg_top_curr[11] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold139 (.A(\systolic_array.genblk1[3].out_queue_dlygate[11].A ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0033_),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold141 (.A(\systolic_array.genblk1[7].out_queue_dlygate[16].A ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0070_),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold143 (.A(\systolic_array.genblk1[9].out_queue_dlygate[11].A ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0081_),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold145 (.A(\systolic_array.genblk1[9].out_queue_dlygate[15].A ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0085_),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold147 (.A(\systolic_array.genblk1[11].out_queue_dlygate[15].A ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0021_),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold149 (.A(\systolic_array.genblk1[1].out_queue_dlygate[10].A ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0008_),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold151 (.A(\systolic_array.genblk1[1].out_queue_dlygate[13].A ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0011_),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold153 (.A(\systolic_array.genblk1[7].out_queue_dlygate[14].A ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0068_),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold155 (.A(\systolic_array.genblk1[11].out_queue_dlygate[13].A ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0125_),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold157 (.A(\systolic_array.genblk1[10].out_queue_dlygate[9].A ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold158 (.A(\systolic_array.genblk1[10].accumulators_dlygate[13].A ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold159 (.A(\systolic_array.genblk1[11].out_queue_dlygate[9].A ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0121_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold161 (.A(\systolic_array.genblk1[3].out_queue_dlygate[16].A ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0038_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold163 (.A(\systolic_array.genblk1[11].out_queue_dlygate[10].A ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0016_),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold165 (.A(\systolic_array.genblk1[9].out_queue_dlygate[9].A ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0087_),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold167 (.A(\systolic_array.arg_left_mul2_next[2] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0163_),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold169 (.A(\systolic_array.arg_left_mul2_next[0] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0161_),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold171 (.A(\systolic_array.genblk1[9].out_queue_dlygate[12].A ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0082_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold173 (.A(\systolic_array.genblk1[11].accumulators_dlygate[14].A ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold174 (.A(\systolic_array.genblk1[11].out_queue_dlygate[12].A ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0018_),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold176 (.A(\systolic_array.genblk1[11].accumulators_dlygate[13].A ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold177 (.A(\systolic_array.genblk1[11].out_queue_dlygate[16].A ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold178 (.A(\systolic_array.genblk1[11].out_queue_dlygate[11].A ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0017_),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold180 (.A(\systolic_array.genblk1[3].out_queue_dlygate[13].A ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0035_),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold182 (.A(\systolic_array.genblk1[3].out_queue_dlygate[10].A ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0032_),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold184 (.A(\systolic_array.genblk1[5].out_queue_dlygate[11].A ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0049_),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold186 (.A(\systolic_array.genblk1[9].out_queue_dlygate[13].A ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0083_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold188 (.A(\systolic_array.genblk1[10].out_queue_dlygate[16].A ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold189 (.A(\systolic_array.arg_left_sign_next[1] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0168_),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold191 (.A(\systolic_array.arg_top_next[10] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold192 (.A(\systolic_array.genblk1[8].out_queue_dlygate[10].A ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold193 (.A(\systolic_array.genblk1[2].out_queue_dlygate[12].A ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold194 (.A(\systolic_array.arg_left_zero_next[0] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold195 (.A(\systolic_array.genblk1[10].accumulators_dlygate[16].A ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold196 (.A(\systolic_array.genblk1[10].out_queue_dlygate[11].A ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold197 (.A(\systolic_array.arg_left_zero_next[3] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold198 (.A(\systolic_array.genblk1[8].out_queue_dlygate[11].A ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold199 (.A(\systolic_array.genblk1[11].accumulators_dlygate[9].A ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold200 (.A(\systolic_array.genblk1[4].out_queue_dlygate[16].A ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold201 (.A(\systolic_array.genblk1[4].out_queue_dlygate[13].A ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold202 (.A(\systolic_array.genblk1[1].out_queue_dlygate[16].A ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0014_),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold204 (.A(\systolic_array.genblk1[9].out_queue_dlygate[16].A ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0086_),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold206 (.A(\systolic_array.genblk1[4].out_queue_dlygate[10].A ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold207 (.A(\systolic_array.genblk1[2].out_queue_dlygate[15].A ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold208 (.A(\systolic_array.genblk1[6].out_queue_dlygate[12].A ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold209 (.A(\systolic_array.genblk1[6].out_queue_dlygate[9].A ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold210 (.A(\systolic_array.arg_left_sign_next[0] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0167_),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold212 (.A(\systolic_array.genblk1[4].out_queue_dlygate[14].A ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold213 (.A(\systolic_array.genblk1[8].out_queue_dlygate[14].A ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold214 (.A(\systolic_array.genblk1[6].out_queue_dlygate[13].A ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold215 (.A(\systolic_array.arg_left_div2_next[0] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0363_),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold217 (.A(\systolic_array.arg_left_div2_next[4] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold218 (.A(\systolic_array.genblk1[4].out_queue_dlygate[9].A ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold219 (.A(\systolic_array.genblk1[3].out_queue_dlygate[9].A ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0039_),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold221 (.A(\systolic_array.arg_top_curr[12] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold222 (.A(\systolic_array.genblk1[2].out_queue_dlygate[14].A ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold223 (.A(\systolic_array.genblk1[5].out_queue_dlygate[9].A ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0055_),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold225 (.A(\systolic_array.genblk1[3].out_queue_dlygate[12].A ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold226 (.A(\systolic_array.genblk1[8].out_queue_dlygate[9].A ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold227 (.A(\systolic_array.genblk1[6].out_queue_dlygate[11].A ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold228 (.A(\systolic_array.genblk1[2].out_queue_dlygate[16].A ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold229 (.A(\systolic_array.genblk1[4].out_queue_dlygate[11].A ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold230 (.A(\systolic_array.genblk1[2].out_queue_dlygate[10].A ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold231 (.A(\systolic_array.genblk1[10].out_queue_dlygate[10].A ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold232 (.A(\systolic_array.genblk1[4].out_queue_dlygate[15].A ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold233 (.A(\systolic_array.genblk1[10].out_queue_dlygate[14].A ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold234 (.A(\systolic_array.genblk1[6].out_queue_dlygate[14].A ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold235 (.A(\systolic_array.genblk1[8].out_queue_dlygate[16].A ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold236 (.A(\systolic_array.genblk1[6].out_queue_dlygate[16].A ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold237 (.A(\systolic_array.genblk1[6].out_queue_dlygate[10].A ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold238 (.A(\systolic_array.genblk1[6].out_queue_dlygate[15].A ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold239 (.A(\systolic_array.arg_left_sign_next[5] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0172_),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold241 (.A(\systolic_array.genblk1[10].out_queue_dlygate[12].A ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold242 (.A(\systolic_array.genblk1[8].out_queue_dlygate[13].A ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold243 (.A(\systolic_array.genblk1[10].out_queue_dlygate[15].A ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold244 (.A(\systolic_array.genblk1[10].accumulators_dlygate[9].A ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold245 (.A(\systolic_array.genblk1[5].out_queue_dlygate[10].A ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0048_),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold247 (.A(\systolic_array.genblk1[8].out_queue_dlygate[15].A ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold248 (.A(\systolic_array.genblk1[10].out_queue_dlygate[13].A ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold249 (.A(\systolic_array.arg_left_zero_next[5] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold250 (.A(\systolic_array.arg_left_zero_next[1] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold251 (.A(\systolic_array.genblk1[2].out_queue_dlygate[11].A ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold252 (.A(\systolic_array.genblk1[7].out_queue_dlygate[12].A ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold253 (.A(\systolic_array.genblk1[0].accumulators_dlygate[8].A ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0218_),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold255 (.A(\systolic_array.genblk1[7].out_queue_dlygate[13].A ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0067_),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold257 (.A(\systolic_array.genblk1[10].accumulators_dlygate[0].A ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold258 (.A(\systolic_array.slice_counter ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold259 (.A(\systolic_array.genblk1[1].out_queue_dlygate[15].A ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0013_),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold261 (.A(\systolic_array.genblk1[8].out_queue_dlygate[12].A ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold262 (.A(\systolic_array.genblk1[4].accumulators_dlygate[1].A ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0279_),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold264 (.A(\systolic_array.genblk1[2].out_queue_dlygate[9].A ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold265 (.A(\systolic_array.genblk1[7].out_queue_dlygate[15].A ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold266 (.A(\systolic_array.genblk1[2].accumulators_dlygate[4].A ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold267 (.A(\systolic_array.genblk1[2].out_queue_dlygate[13].A ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold268 (.A(\systolic_array.genblk1[8].accumulators_dlygate[0].A ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold269 (.A(_1410_),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold270 (.A(\systolic_array.genblk1[5].out_queue_dlygate[15].A ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold271 (.A(\systolic_array.genblk1[4].accumulators_dlygate[2].A ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0280_),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold273 (.A(\systolic_array.genblk1[9].out_queue_dlygate[14].A ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0084_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold275 (.A(\systolic_array.genblk1[10].accumulators_dlygate[1].A ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0368_),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold277 (.A(\systolic_array.arg_top_curr[9] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold278 (.A(\systolic_array.genblk1[3].out_queue_dlygate[15].A ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0037_),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold280 (.A(\systolic_array.genblk1[3].out_queue_dlygate[14].A ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0036_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold282 (.A(\systolic_array.genblk1[4].accumulators_dlygate[0].A ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold283 (.A(\systolic_array.arg_left_mul2_next[5] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold284 (.A(\systolic_array.genblk1[4].out_queue_dlygate[12].A ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold285 (.A(\systolic_array.genblk1[8].accumulators_dlygate[4].A ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold286 (.A(\systolic_array.genblk1[7].out_queue_dlygate[10].A ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0064_),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold288 (.A(\systolic_array.genblk1[0].accumulators_dlygate[5].A ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold289 (.A(\systolic_array.genblk1[2].accumulators_dlygate[7].A ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold290 (.A(\systolic_array.genblk1[6].accumulators_dlygate[3].A ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold291 (.A(\systolic_array.genblk1[4].accumulators_dlygate[6].A ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0284_),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold293 (.A(\systolic_array.genblk1[5].out_queue_dlygate[16].A ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold294 (.A(_0054_),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold295 (.A(\systolic_array.arg_top_curr[10] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold296 (.A(\systolic_array.genblk1[0].accumulators_dlygate[1].A ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0211_),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold298 (.A(\systolic_array.genblk1[6].accumulators_dlygate[6].A ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0318_),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold300 (.A(\systolic_array.genblk1[8].accumulators_dlygate[3].A ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold301 (.A(\systolic_array.genblk1[0].accumulators_dlygate[0].A ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold302 (.A(_1312_),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold303 (.A(\systolic_array.genblk2[0].mac[5].mul2 ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold304 (.A(\systolic_array.genblk1[2].accumulators_dlygate[1].A ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold305 (.A(\systolic_array.genblk1[6].accumulators_dlygate[8].A ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold306 (.A(\systolic_array.genblk1[2].accumulators_dlygate[0].A ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold307 (.A(\systolic_array.arg_left_mul2_next[3] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0164_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold309 (.A(\systolic_array.genblk1[5].out_queue_dlygate[12].A ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold310 (.A(\systolic_array.genblk1[10].accumulators_dlygate[11].A ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold311 (.A(\systolic_array.genblk1[10].accumulators_dlygate[8].A ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold312 (.A(\systolic_array.genblk1[0].accumulators_dlygate[16].A ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold313 (.A(\systolic_array.genblk1[2].accumulators_dlygate[6].A ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0250_),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold315 (.A(\systolic_array.genblk1[10].accumulators_dlygate[5].A ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0372_),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold317 (.A(\systolic_array.genblk1[2].accumulators_dlygate[2].A ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold318 (.A(\systolic_array.genblk1[2].accumulators_dlygate[16].A ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold319 (.A(\systolic_array.genblk1[0].accumulators_dlygate[4].A ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0214_),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold321 (.A(\systolic_array.genblk1[7].out_queue_dlygate[9].A ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold322 (.A(_0071_),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold323 (.A(\systolic_array.genblk2[0].mac[4].div2 ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold324 (.A(\systolic_array.genblk1[0].accumulators_dlygate[2].A ),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold325 (.A(\systolic_array.arg_left_zero_next[4] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold326 (.A(\systolic_array.genblk1[7].out_queue_dlygate[11].A ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold327 (.A(_0065_),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold328 (.A(\systolic_array.genblk1[4].accumulators_dlygate[8].A ),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold329 (.A(\systolic_array.arg_top_curr[14] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold330 (.A(\systolic_array.genblk1[2].accumulators_dlygate[8].A ),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold331 (.A(\systolic_array.genblk1[6].accumulators_dlygate[1].A ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold332 (.A(\systolic_array.genblk1[6].accumulators_dlygate[0].A ),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold333 (.A(\systolic_array.genblk1[4].accumulators_dlygate[3].A ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold334 (.A(\systolic_array.genblk1[0].accumulators_dlygate[3].A ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold335 (.A(\systolic_array.genblk1[4].accumulators_dlygate[16].A ),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold336 (.A(\systolic_array.arg_top_curr[8] ),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold337 (.A(\systolic_array.arg_left_div2_next[3] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold338 (.A(\systolic_array.genblk1[6].accumulators_dlygate[16].A ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold339 (.A(\systolic_array.genblk1[0].accumulators_dlygate[6].A ),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold340 (.A(\systolic_array.genblk1[6].accumulators_dlygate[7].A ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0319_),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold342 (.A(\systolic_array.genblk1[8].accumulators_dlygate[2].A ),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold343 (.A(\systolic_array.genblk1[6].accumulators_dlygate[2].A ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold344 (.A(\systolic_array.genblk1[10].accumulators_dlygate[3].A ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold345 (.A(\systolic_array.genblk1[4].accumulators_dlygate[11].A ),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold346 (.A(\systolic_array.arg_top_curr[15] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold347 (.A(\systolic_array.genblk1[5].out_queue_dlygate[13].A ),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0051_),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold349 (.A(\systolic_array.genblk1[4].accumulators_dlygate[5].A ),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold350 (.A(\systolic_array.genblk1[4].accumulators_dlygate[7].A ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0285_),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold352 (.A(\systolic_array.genblk1[8].accumulators_dlygate[8].A ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold353 (.A(\systolic_array.genblk1[2].accumulators_dlygate[3].A ),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold354 (.A(\systolic_array.genblk1[6].accumulators_dlygate[4].A ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold355 (.A(\systolic_array.genblk1[8].accumulators_dlygate[1].A ),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0347_),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold357 (.A(\systolic_array.genblk1[10].accumulators_dlygate[4].A ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold358 (.A(\systolic_array.genblk1[8].accumulators_dlygate[6].A ),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold359 (.A(\systolic_array.genblk1[10].accumulators_dlygate[6].A ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold360 (.A(\systolic_array.genblk1[8].accumulators_dlygate[7].A ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold361 (.A(\systolic_array.genblk1[8].accumulators_dlygate[16].A ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold362 (.A(\systolic_array.arg_left_sign_next[3] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold363 (.A(\systolic_array.genblk1[2].accumulators_dlygate[11].A ),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold364 (.A(\systolic_array.genblk1[10].accumulators_dlygate[7].A ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold365 (.A(\systolic_array.genblk1[2].accumulators_dlygate[15].A ),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold366 (.A(\systolic_array.genblk1[10].accumulators_dlygate[2].A ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0369_),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold368 (.A(\systolic_array.genblk2[0].mac[3].sign ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold369 (.A(\systolic_array.genblk1[0].accumulators_dlygate[9].A ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold370 (.A(\systolic_array.genblk1[2].accumulators_dlygate[9].A ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold371 (.A(\systolic_array.genblk1[10].accumulators_dlygate[15].A ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold372 (.A(\systolic_array.arg_top_curr[13] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold373 (.A(\systolic_array.genblk1[0].accumulators_dlygate[7].A ),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold374 (.A(\systolic_array.genblk1[4].accumulators_dlygate[4].A ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold375 (.A(\systolic_array.genblk1[6].accumulators_dlygate[9].A ),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold376 (.A(\systolic_array.genblk1[10].accumulators_dlygate[14].A ),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold377 (.A(\systolic_array.genblk1[6].accumulators_dlygate[10].A ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold378 (.A(\systolic_array.genblk1[6].accumulators_dlygate[5].A ),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold379 (.A(\systolic_array.genblk1[0].accumulators_dlygate[11].A ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold380 (.A(\systolic_array.genblk1[2].accumulators_dlygate[5].A ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold381 (.A(\systolic_array.genblk1[4].accumulators_dlygate[9].A ),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold382 (.A(\systolic_array.genblk1[2].accumulators_dlygate[13].A ),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold383 (.A(\systolic_array.genblk1[6].accumulators_dlygate[13].A ),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold384 (.A(\systolic_array.genblk1[2].accumulators_dlygate[14].A ),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold385 (.A(\systolic_array.genblk1[8].accumulators_dlygate[13].A ),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold386 (.A(\systolic_array.genblk1[4].accumulators_dlygate[13].A ),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold387 (.A(\systolic_array.arg_left_sign_next[4] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold388 (.A(\systolic_array.genblk1[8].accumulators_dlygate[5].A ),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0351_),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold390 (.A(\systolic_array.genblk1[6].accumulators_dlygate[11].A ),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold391 (.A(\systolic_array.genblk2[0].mac[4].zero ),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold392 (.A(\systolic_array.genblk1[8].accumulators_dlygate[14].A ),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold393 (.A(\systolic_array.genblk1[10].accumulators_dlygate[10].A ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold394 (.A(\systolic_array.arg_left_mul2_next[4] ),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold395 (.A(\systolic_array.genblk1[4].accumulators_dlygate[10].A ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold396 (.A(\systolic_array.genblk1[0].accumulators_dlygate[10].A ),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold397 (.A(\systolic_array.genblk2[0].mac[4].sign ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold398 (.A(\systolic_array.genblk1[0].accumulators_dlygate[13].A ),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold399 (.A(\systolic_array.genblk1[8].accumulators_dlygate[11].A ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold400 (.A(\systolic_array.genblk1[8].accumulators_dlygate[9].A ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold401 (.A(\systolic_array.genblk1[0].accumulators_dlygate[14].A ),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold402 (.A(\systolic_array.genblk1[6].accumulators_dlygate[14].A ),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold403 (.A(\systolic_array.genblk1[10].accumulators_dlygate[12].A ),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold404 (.A(\systolic_array.genblk1[0].accumulators_dlygate[15].A ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold405 (.A(\systolic_array.genblk1[8].accumulators_dlygate[10].A ),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold406 (.A(\systolic_array.genblk1[4].accumulators_dlygate[15].A ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold407 (.A(\systolic_array.genblk1[2].accumulators_dlygate[10].A ),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold408 (.A(_0514_),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold409 (.A(\systolic_array.genblk1[0].accumulators_dlygate[12].A ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold410 (.A(\systolic_array.genblk1[4].accumulators_dlygate[12].A ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold411 (.A(\systolic_array.genblk1[2].accumulators_dlygate[12].A ),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold412 (.A(\systolic_array.genblk1[4].accumulators_dlygate[14].A ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold413 (.A(\systolic_array.genblk1[8].accumulators_dlygate[15].A ),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold414 (.A(\systolic_array.genblk1[8].accumulators_dlygate[12].A ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold415 (.A(\systolic_array.genblk1[6].accumulators_dlygate[15].A ),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold416 (.A(\systolic_array.genblk1[6].accumulators_dlygate[12].A ),
    .X(net999));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_4 FILLER_0_28 ();
 sg13g2_decap_4 FILLER_0_36 ();
 sg13g2_fill_1 FILLER_0_66 ();
 sg13g2_fill_2 FILLER_0_90 ();
 sg13g2_fill_1 FILLER_0_92 ();
 sg13g2_fill_2 FILLER_0_103 ();
 sg13g2_fill_1 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_124 ();
 sg13g2_decap_8 FILLER_0_131 ();
 sg13g2_decap_4 FILLER_0_138 ();
 sg13g2_decap_8 FILLER_0_150 ();
 sg13g2_decap_8 FILLER_0_157 ();
 sg13g2_decap_8 FILLER_0_164 ();
 sg13g2_decap_8 FILLER_0_171 ();
 sg13g2_decap_8 FILLER_0_178 ();
 sg13g2_decap_8 FILLER_0_185 ();
 sg13g2_decap_8 FILLER_0_192 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_decap_8 FILLER_0_206 ();
 sg13g2_decap_8 FILLER_0_213 ();
 sg13g2_decap_8 FILLER_0_220 ();
 sg13g2_decap_4 FILLER_0_231 ();
 sg13g2_fill_2 FILLER_0_235 ();
 sg13g2_decap_4 FILLER_0_241 ();
 sg13g2_fill_1 FILLER_0_245 ();
 sg13g2_fill_2 FILLER_0_250 ();
 sg13g2_fill_2 FILLER_0_260 ();
 sg13g2_fill_1 FILLER_0_262 ();
 sg13g2_fill_2 FILLER_0_268 ();
 sg13g2_fill_1 FILLER_0_270 ();
 sg13g2_fill_2 FILLER_0_276 ();
 sg13g2_fill_1 FILLER_0_278 ();
 sg13g2_decap_4 FILLER_0_283 ();
 sg13g2_decap_8 FILLER_0_292 ();
 sg13g2_decap_8 FILLER_0_299 ();
 sg13g2_fill_2 FILLER_0_306 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_4 FILLER_1_14 ();
 sg13g2_fill_2 FILLER_1_18 ();
 sg13g2_fill_2 FILLER_1_34 ();
 sg13g2_fill_1 FILLER_1_67 ();
 sg13g2_fill_2 FILLER_1_94 ();
 sg13g2_fill_2 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_180 ();
 sg13g2_decap_4 FILLER_1_187 ();
 sg13g2_fill_1 FILLER_1_191 ();
 sg13g2_fill_1 FILLER_1_244 ();
 sg13g2_fill_2 FILLER_1_280 ();
 sg13g2_fill_2 FILLER_1_287 ();
 sg13g2_fill_1 FILLER_1_289 ();
 sg13g2_fill_2 FILLER_1_299 ();
 sg13g2_decap_8 FILLER_1_335 ();
 sg13g2_decap_8 FILLER_1_342 ();
 sg13g2_decap_8 FILLER_1_349 ();
 sg13g2_decap_8 FILLER_1_356 ();
 sg13g2_decap_8 FILLER_1_363 ();
 sg13g2_decap_8 FILLER_1_370 ();
 sg13g2_decap_8 FILLER_1_377 ();
 sg13g2_decap_8 FILLER_1_384 ();
 sg13g2_decap_8 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_398 ();
 sg13g2_decap_4 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_fill_2 FILLER_2_14 ();
 sg13g2_fill_2 FILLER_2_72 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_4 FILLER_2_196 ();
 sg13g2_fill_2 FILLER_2_282 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_4 FILLER_3_14 ();
 sg13g2_fill_1 FILLER_3_22 ();
 sg13g2_fill_1 FILLER_3_49 ();
 sg13g2_fill_2 FILLER_3_90 ();
 sg13g2_fill_2 FILLER_3_106 ();
 sg13g2_fill_2 FILLER_3_150 ();
 sg13g2_fill_1 FILLER_3_171 ();
 sg13g2_fill_1 FILLER_3_179 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_fill_1 FILLER_3_196 ();
 sg13g2_fill_2 FILLER_3_214 ();
 sg13g2_fill_1 FILLER_3_216 ();
 sg13g2_fill_2 FILLER_3_226 ();
 sg13g2_fill_1 FILLER_3_228 ();
 sg13g2_fill_2 FILLER_3_248 ();
 sg13g2_fill_1 FILLER_3_307 ();
 sg13g2_decap_8 FILLER_3_334 ();
 sg13g2_decap_8 FILLER_3_341 ();
 sg13g2_decap_8 FILLER_3_348 ();
 sg13g2_decap_8 FILLER_3_355 ();
 sg13g2_decap_8 FILLER_3_362 ();
 sg13g2_decap_8 FILLER_3_369 ();
 sg13g2_decap_8 FILLER_3_376 ();
 sg13g2_decap_8 FILLER_3_383 ();
 sg13g2_decap_8 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_103 ();
 sg13g2_fill_2 FILLER_4_114 ();
 sg13g2_fill_1 FILLER_4_116 ();
 sg13g2_fill_2 FILLER_4_261 ();
 sg13g2_fill_1 FILLER_4_288 ();
 sg13g2_fill_1 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_339 ();
 sg13g2_decap_8 FILLER_4_346 ();
 sg13g2_decap_8 FILLER_4_353 ();
 sg13g2_decap_8 FILLER_4_360 ();
 sg13g2_decap_8 FILLER_4_367 ();
 sg13g2_decap_8 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_fill_2 FILLER_5_14 ();
 sg13g2_fill_1 FILLER_5_16 ();
 sg13g2_fill_1 FILLER_5_98 ();
 sg13g2_fill_2 FILLER_5_133 ();
 sg13g2_fill_1 FILLER_5_176 ();
 sg13g2_fill_2 FILLER_5_186 ();
 sg13g2_fill_2 FILLER_5_253 ();
 sg13g2_fill_2 FILLER_5_280 ();
 sg13g2_fill_1 FILLER_5_282 ();
 sg13g2_fill_2 FILLER_5_297 ();
 sg13g2_fill_1 FILLER_5_299 ();
 sg13g2_fill_1 FILLER_5_309 ();
 sg13g2_decap_4 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_4 FILLER_6_21 ();
 sg13g2_fill_1 FILLER_6_38 ();
 sg13g2_decap_4 FILLER_6_96 ();
 sg13g2_fill_1 FILLER_6_145 ();
 sg13g2_fill_2 FILLER_6_172 ();
 sg13g2_fill_1 FILLER_6_218 ();
 sg13g2_fill_2 FILLER_6_256 ();
 sg13g2_decap_4 FILLER_6_310 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_4 FILLER_6_403 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_fill_1 FILLER_7_66 ();
 sg13g2_fill_2 FILLER_7_71 ();
 sg13g2_fill_1 FILLER_7_73 ();
 sg13g2_fill_2 FILLER_7_104 ();
 sg13g2_fill_1 FILLER_7_119 ();
 sg13g2_fill_1 FILLER_7_151 ();
 sg13g2_fill_1 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_194 ();
 sg13g2_decap_8 FILLER_7_201 ();
 sg13g2_decap_8 FILLER_7_208 ();
 sg13g2_fill_2 FILLER_7_243 ();
 sg13g2_fill_1 FILLER_7_245 ();
 sg13g2_decap_4 FILLER_7_250 ();
 sg13g2_fill_2 FILLER_7_254 ();
 sg13g2_fill_1 FILLER_7_274 ();
 sg13g2_decap_8 FILLER_7_363 ();
 sg13g2_decap_8 FILLER_7_370 ();
 sg13g2_decap_8 FILLER_7_377 ();
 sg13g2_decap_8 FILLER_7_384 ();
 sg13g2_decap_8 FILLER_7_391 ();
 sg13g2_decap_8 FILLER_7_398 ();
 sg13g2_decap_4 FILLER_7_405 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_28 ();
 sg13g2_fill_1 FILLER_8_82 ();
 sg13g2_fill_1 FILLER_8_175 ();
 sg13g2_fill_1 FILLER_8_185 ();
 sg13g2_decap_4 FILLER_8_191 ();
 sg13g2_fill_2 FILLER_8_195 ();
 sg13g2_fill_1 FILLER_8_201 ();
 sg13g2_fill_1 FILLER_8_221 ();
 sg13g2_fill_1 FILLER_8_235 ();
 sg13g2_decap_4 FILLER_8_262 ();
 sg13g2_fill_1 FILLER_8_266 ();
 sg13g2_fill_2 FILLER_8_298 ();
 sg13g2_fill_1 FILLER_8_300 ();
 sg13g2_fill_1 FILLER_8_310 ();
 sg13g2_decap_8 FILLER_8_360 ();
 sg13g2_decap_8 FILLER_8_367 ();
 sg13g2_decap_8 FILLER_8_374 ();
 sg13g2_decap_8 FILLER_8_381 ();
 sg13g2_decap_8 FILLER_8_388 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_4 ();
 sg13g2_fill_1 FILLER_9_55 ();
 sg13g2_fill_1 FILLER_9_80 ();
 sg13g2_fill_1 FILLER_9_133 ();
 sg13g2_fill_2 FILLER_9_153 ();
 sg13g2_fill_1 FILLER_9_170 ();
 sg13g2_fill_2 FILLER_9_217 ();
 sg13g2_fill_1 FILLER_9_229 ();
 sg13g2_fill_2 FILLER_9_261 ();
 sg13g2_decap_8 FILLER_9_275 ();
 sg13g2_decap_8 FILLER_9_282 ();
 sg13g2_decap_8 FILLER_9_289 ();
 sg13g2_fill_1 FILLER_9_305 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_fill_1 FILLER_9_344 ();
 sg13g2_decap_8 FILLER_9_390 ();
 sg13g2_decap_8 FILLER_9_397 ();
 sg13g2_decap_4 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_fill_1 FILLER_10_14 ();
 sg13g2_fill_2 FILLER_10_41 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_fill_2 FILLER_10_95 ();
 sg13g2_fill_2 FILLER_10_127 ();
 sg13g2_fill_1 FILLER_10_221 ();
 sg13g2_decap_8 FILLER_10_227 ();
 sg13g2_fill_2 FILLER_10_247 ();
 sg13g2_decap_8 FILLER_10_275 ();
 sg13g2_decap_4 FILLER_10_282 ();
 sg13g2_decap_8 FILLER_10_290 ();
 sg13g2_decap_4 FILLER_10_297 ();
 sg13g2_fill_1 FILLER_10_301 ();
 sg13g2_decap_4 FILLER_10_306 ();
 sg13g2_fill_2 FILLER_10_310 ();
 sg13g2_decap_8 FILLER_10_320 ();
 sg13g2_fill_1 FILLER_10_327 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_4 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_39 ();
 sg13g2_fill_1 FILLER_11_41 ();
 sg13g2_fill_2 FILLER_11_61 ();
 sg13g2_fill_1 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_73 ();
 sg13g2_decap_4 FILLER_11_80 ();
 sg13g2_fill_1 FILLER_11_84 ();
 sg13g2_fill_2 FILLER_11_89 ();
 sg13g2_decap_4 FILLER_11_99 ();
 sg13g2_decap_4 FILLER_11_120 ();
 sg13g2_fill_2 FILLER_11_124 ();
 sg13g2_fill_2 FILLER_11_152 ();
 sg13g2_fill_1 FILLER_11_154 ();
 sg13g2_fill_1 FILLER_11_164 ();
 sg13g2_fill_2 FILLER_11_186 ();
 sg13g2_fill_1 FILLER_11_201 ();
 sg13g2_fill_1 FILLER_11_216 ();
 sg13g2_fill_2 FILLER_11_222 ();
 sg13g2_fill_1 FILLER_11_224 ();
 sg13g2_decap_4 FILLER_11_238 ();
 sg13g2_fill_1 FILLER_11_242 ();
 sg13g2_fill_2 FILLER_11_265 ();
 sg13g2_fill_1 FILLER_11_267 ();
 sg13g2_fill_1 FILLER_11_275 ();
 sg13g2_decap_8 FILLER_11_302 ();
 sg13g2_decap_8 FILLER_11_309 ();
 sg13g2_decap_8 FILLER_11_316 ();
 sg13g2_fill_2 FILLER_11_323 ();
 sg13g2_fill_1 FILLER_11_325 ();
 sg13g2_fill_1 FILLER_11_347 ();
 sg13g2_fill_2 FILLER_11_362 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_17 ();
 sg13g2_fill_2 FILLER_12_21 ();
 sg13g2_fill_2 FILLER_12_57 ();
 sg13g2_fill_1 FILLER_12_59 ();
 sg13g2_fill_2 FILLER_12_78 ();
 sg13g2_fill_1 FILLER_12_80 ();
 sg13g2_fill_2 FILLER_12_141 ();
 sg13g2_fill_1 FILLER_12_143 ();
 sg13g2_fill_2 FILLER_12_160 ();
 sg13g2_fill_1 FILLER_12_162 ();
 sg13g2_fill_2 FILLER_12_171 ();
 sg13g2_fill_2 FILLER_12_183 ();
 sg13g2_fill_2 FILLER_12_225 ();
 sg13g2_fill_1 FILLER_12_243 ();
 sg13g2_fill_1 FILLER_12_252 ();
 sg13g2_fill_2 FILLER_12_329 ();
 sg13g2_fill_1 FILLER_12_331 ();
 sg13g2_fill_1 FILLER_12_341 ();
 sg13g2_decap_4 FILLER_12_355 ();
 sg13g2_fill_1 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_4 FILLER_13_28 ();
 sg13g2_fill_1 FILLER_13_32 ();
 sg13g2_fill_1 FILLER_13_44 ();
 sg13g2_fill_1 FILLER_13_86 ();
 sg13g2_fill_2 FILLER_13_113 ();
 sg13g2_fill_2 FILLER_13_141 ();
 sg13g2_fill_2 FILLER_13_152 ();
 sg13g2_fill_1 FILLER_13_154 ();
 sg13g2_fill_2 FILLER_13_181 ();
 sg13g2_fill_1 FILLER_13_306 ();
 sg13g2_decap_8 FILLER_13_328 ();
 sg13g2_decap_4 FILLER_13_335 ();
 sg13g2_fill_1 FILLER_13_339 ();
 sg13g2_decap_4 FILLER_13_348 ();
 sg13g2_fill_1 FILLER_13_352 ();
 sg13g2_decap_4 FILLER_13_358 ();
 sg13g2_fill_2 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_fill_1 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_32 ();
 sg13g2_fill_2 FILLER_14_39 ();
 sg13g2_fill_1 FILLER_14_57 ();
 sg13g2_fill_2 FILLER_14_149 ();
 sg13g2_fill_1 FILLER_14_151 ();
 sg13g2_fill_2 FILLER_14_166 ();
 sg13g2_fill_2 FILLER_14_177 ();
 sg13g2_decap_8 FILLER_14_188 ();
 sg13g2_fill_2 FILLER_14_195 ();
 sg13g2_fill_1 FILLER_14_197 ();
 sg13g2_fill_1 FILLER_14_235 ();
 sg13g2_fill_1 FILLER_14_241 ();
 sg13g2_fill_2 FILLER_14_267 ();
 sg13g2_fill_1 FILLER_14_269 ();
 sg13g2_decap_4 FILLER_14_334 ();
 sg13g2_fill_1 FILLER_14_338 ();
 sg13g2_fill_2 FILLER_14_362 ();
 sg13g2_fill_1 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_12 ();
 sg13g2_decap_4 FILLER_15_19 ();
 sg13g2_fill_2 FILLER_15_46 ();
 sg13g2_fill_1 FILLER_15_53 ();
 sg13g2_fill_1 FILLER_15_58 ();
 sg13g2_decap_4 FILLER_15_84 ();
 sg13g2_fill_2 FILLER_15_131 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_fill_2 FILLER_15_210 ();
 sg13g2_fill_1 FILLER_15_212 ();
 sg13g2_fill_2 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_fill_2 FILLER_15_231 ();
 sg13g2_fill_2 FILLER_15_259 ();
 sg13g2_fill_2 FILLER_15_290 ();
 sg13g2_fill_1 FILLER_15_297 ();
 sg13g2_fill_2 FILLER_15_306 ();
 sg13g2_fill_2 FILLER_15_317 ();
 sg13g2_fill_1 FILLER_15_319 ();
 sg13g2_fill_2 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_2 ();
 sg13g2_decap_4 FILLER_16_76 ();
 sg13g2_fill_2 FILLER_16_80 ();
 sg13g2_fill_2 FILLER_16_121 ();
 sg13g2_fill_1 FILLER_16_123 ();
 sg13g2_decap_8 FILLER_16_199 ();
 sg13g2_decap_8 FILLER_16_206 ();
 sg13g2_fill_1 FILLER_16_213 ();
 sg13g2_decap_8 FILLER_16_218 ();
 sg13g2_decap_8 FILLER_16_225 ();
 sg13g2_decap_8 FILLER_16_232 ();
 sg13g2_decap_4 FILLER_16_239 ();
 sg13g2_fill_1 FILLER_16_243 ();
 sg13g2_decap_8 FILLER_16_248 ();
 sg13g2_decap_8 FILLER_16_255 ();
 sg13g2_decap_4 FILLER_16_266 ();
 sg13g2_fill_2 FILLER_16_270 ();
 sg13g2_fill_1 FILLER_16_296 ();
 sg13g2_fill_1 FILLER_16_305 ();
 sg13g2_fill_2 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_2 ();
 sg13g2_fill_2 FILLER_17_64 ();
 sg13g2_fill_1 FILLER_17_120 ();
 sg13g2_decap_4 FILLER_17_199 ();
 sg13g2_decap_4 FILLER_17_234 ();
 sg13g2_fill_2 FILLER_17_238 ();
 sg13g2_fill_1 FILLER_17_246 ();
 sg13g2_fill_2 FILLER_17_256 ();
 sg13g2_fill_2 FILLER_17_269 ();
 sg13g2_fill_1 FILLER_17_271 ();
 sg13g2_fill_2 FILLER_17_288 ();
 sg13g2_fill_2 FILLER_17_306 ();
 sg13g2_fill_1 FILLER_17_308 ();
 sg13g2_fill_2 FILLER_17_319 ();
 sg13g2_decap_4 FILLER_17_364 ();
 sg13g2_fill_2 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_fill_1 FILLER_18_26 ();
 sg13g2_fill_2 FILLER_18_101 ();
 sg13g2_fill_1 FILLER_18_103 ();
 sg13g2_fill_2 FILLER_18_207 ();
 sg13g2_fill_1 FILLER_18_214 ();
 sg13g2_fill_1 FILLER_18_272 ();
 sg13g2_decap_4 FILLER_18_289 ();
 sg13g2_fill_1 FILLER_18_293 ();
 sg13g2_fill_2 FILLER_18_298 ();
 sg13g2_decap_4 FILLER_18_304 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_41 ();
 sg13g2_fill_2 FILLER_19_51 ();
 sg13g2_fill_1 FILLER_19_53 ();
 sg13g2_fill_2 FILLER_19_64 ();
 sg13g2_fill_2 FILLER_19_105 ();
 sg13g2_fill_1 FILLER_19_107 ();
 sg13g2_fill_2 FILLER_19_144 ();
 sg13g2_fill_1 FILLER_19_146 ();
 sg13g2_fill_2 FILLER_19_152 ();
 sg13g2_fill_1 FILLER_19_154 ();
 sg13g2_fill_1 FILLER_19_164 ();
 sg13g2_fill_2 FILLER_19_179 ();
 sg13g2_fill_2 FILLER_19_216 ();
 sg13g2_fill_2 FILLER_19_240 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_fill_1 FILLER_19_252 ();
 sg13g2_fill_1 FILLER_19_285 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_4 FILLER_19_336 ();
 sg13g2_fill_2 FILLER_19_340 ();
 sg13g2_fill_1 FILLER_19_358 ();
 sg13g2_fill_1 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_fill_2 FILLER_20_37 ();
 sg13g2_fill_2 FILLER_20_109 ();
 sg13g2_fill_1 FILLER_20_111 ();
 sg13g2_fill_2 FILLER_20_135 ();
 sg13g2_fill_2 FILLER_20_146 ();
 sg13g2_fill_1 FILLER_20_148 ();
 sg13g2_fill_1 FILLER_20_159 ();
 sg13g2_decap_4 FILLER_20_169 ();
 sg13g2_fill_2 FILLER_20_173 ();
 sg13g2_fill_2 FILLER_20_183 ();
 sg13g2_fill_2 FILLER_20_190 ();
 sg13g2_fill_1 FILLER_20_192 ();
 sg13g2_fill_2 FILLER_20_201 ();
 sg13g2_decap_8 FILLER_20_235 ();
 sg13g2_decap_4 FILLER_20_242 ();
 sg13g2_fill_2 FILLER_20_246 ();
 sg13g2_decap_4 FILLER_20_252 ();
 sg13g2_fill_2 FILLER_20_256 ();
 sg13g2_fill_2 FILLER_20_272 ();
 sg13g2_decap_8 FILLER_20_283 ();
 sg13g2_fill_2 FILLER_20_290 ();
 sg13g2_fill_1 FILLER_20_292 ();
 sg13g2_decap_4 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_307 ();
 sg13g2_decap_4 FILLER_20_313 ();
 sg13g2_decap_8 FILLER_20_331 ();
 sg13g2_decap_4 FILLER_20_338 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_63 ();
 sg13g2_fill_1 FILLER_21_85 ();
 sg13g2_fill_2 FILLER_21_214 ();
 sg13g2_fill_1 FILLER_21_216 ();
 sg13g2_fill_2 FILLER_21_226 ();
 sg13g2_fill_1 FILLER_21_228 ();
 sg13g2_fill_1 FILLER_21_233 ();
 sg13g2_fill_2 FILLER_21_257 ();
 sg13g2_fill_2 FILLER_21_325 ();
 sg13g2_fill_1 FILLER_21_327 ();
 sg13g2_decap_8 FILLER_21_384 ();
 sg13g2_decap_8 FILLER_21_391 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_4 FILLER_22_14 ();
 sg13g2_fill_2 FILLER_22_18 ();
 sg13g2_fill_2 FILLER_22_98 ();
 sg13g2_fill_1 FILLER_22_100 ();
 sg13g2_fill_2 FILLER_22_153 ();
 sg13g2_fill_1 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_279 ();
 sg13g2_fill_2 FILLER_22_286 ();
 sg13g2_fill_2 FILLER_22_317 ();
 sg13g2_fill_1 FILLER_22_319 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_4 FILLER_22_357 ();
 sg13g2_decap_4 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_383 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_fill_2 FILLER_23_31 ();
 sg13g2_fill_2 FILLER_23_37 ();
 sg13g2_fill_2 FILLER_23_43 ();
 sg13g2_fill_1 FILLER_23_45 ();
 sg13g2_fill_1 FILLER_23_55 ();
 sg13g2_fill_1 FILLER_23_90 ();
 sg13g2_fill_2 FILLER_23_149 ();
 sg13g2_fill_1 FILLER_23_160 ();
 sg13g2_fill_1 FILLER_23_169 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_decap_8 FILLER_23_278 ();
 sg13g2_fill_2 FILLER_23_285 ();
 sg13g2_fill_2 FILLER_23_296 ();
 sg13g2_decap_4 FILLER_23_303 ();
 sg13g2_fill_2 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_354 ();
 sg13g2_decap_4 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_27 ();
 sg13g2_decap_8 FILLER_24_34 ();
 sg13g2_decap_8 FILLER_24_41 ();
 sg13g2_fill_1 FILLER_24_48 ();
 sg13g2_decap_8 FILLER_24_58 ();
 sg13g2_decap_8 FILLER_24_65 ();
 sg13g2_fill_2 FILLER_24_72 ();
 sg13g2_decap_4 FILLER_24_78 ();
 sg13g2_fill_2 FILLER_24_82 ();
 sg13g2_fill_2 FILLER_24_128 ();
 sg13g2_fill_1 FILLER_24_130 ();
 sg13g2_fill_2 FILLER_24_148 ();
 sg13g2_decap_8 FILLER_24_159 ();
 sg13g2_decap_4 FILLER_24_166 ();
 sg13g2_fill_2 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_fill_2 FILLER_24_320 ();
 sg13g2_fill_2 FILLER_24_330 ();
 sg13g2_fill_1 FILLER_24_332 ();
 sg13g2_decap_4 FILLER_24_337 ();
 sg13g2_fill_2 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_11 ();
 sg13g2_fill_2 FILLER_25_55 ();
 sg13g2_fill_1 FILLER_25_57 ();
 sg13g2_decap_8 FILLER_25_66 ();
 sg13g2_decap_4 FILLER_25_73 ();
 sg13g2_fill_1 FILLER_25_77 ();
 sg13g2_fill_2 FILLER_25_87 ();
 sg13g2_fill_1 FILLER_25_89 ();
 sg13g2_fill_2 FILLER_25_116 ();
 sg13g2_fill_1 FILLER_25_118 ();
 sg13g2_fill_2 FILLER_25_124 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_fill_2 FILLER_25_153 ();
 sg13g2_fill_1 FILLER_25_155 ();
 sg13g2_decap_4 FILLER_25_171 ();
 sg13g2_decap_4 FILLER_25_188 ();
 sg13g2_decap_4 FILLER_25_218 ();
 sg13g2_decap_4 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_313 ();
 sg13g2_decap_8 FILLER_25_320 ();
 sg13g2_decap_4 FILLER_25_327 ();
 sg13g2_fill_1 FILLER_25_331 ();
 sg13g2_fill_2 FILLER_25_368 ();
 sg13g2_fill_1 FILLER_25_370 ();
 sg13g2_fill_2 FILLER_25_388 ();
 sg13g2_fill_1 FILLER_25_390 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_11 ();
 sg13g2_fill_2 FILLER_26_96 ();
 sg13g2_fill_2 FILLER_26_107 ();
 sg13g2_fill_2 FILLER_26_117 ();
 sg13g2_fill_1 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_207 ();
 sg13g2_fill_2 FILLER_26_249 ();
 sg13g2_fill_2 FILLER_26_265 ();
 sg13g2_fill_1 FILLER_26_324 ();
 sg13g2_decap_8 FILLER_26_381 ();
 sg13g2_decap_8 FILLER_26_388 ();
 sg13g2_decap_8 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_4 ();
 sg13g2_fill_2 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_54 ();
 sg13g2_fill_2 FILLER_27_86 ();
 sg13g2_fill_2 FILLER_27_93 ();
 sg13g2_fill_1 FILLER_27_95 ();
 sg13g2_fill_1 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_111 ();
 sg13g2_fill_1 FILLER_27_138 ();
 sg13g2_fill_1 FILLER_27_165 ();
 sg13g2_fill_2 FILLER_27_184 ();
 sg13g2_fill_2 FILLER_27_194 ();
 sg13g2_fill_2 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_267 ();
 sg13g2_decap_8 FILLER_27_290 ();
 sg13g2_fill_2 FILLER_27_340 ();
 sg13g2_fill_2 FILLER_27_374 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_97 ();
 sg13g2_decap_4 FILLER_28_200 ();
 sg13g2_fill_2 FILLER_28_204 ();
 sg13g2_fill_2 FILLER_28_210 ();
 sg13g2_fill_1 FILLER_28_272 ();
 sg13g2_fill_2 FILLER_28_326 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_fill_2 FILLER_29_59 ();
 sg13g2_fill_1 FILLER_29_151 ();
 sg13g2_fill_1 FILLER_29_173 ();
 sg13g2_decap_8 FILLER_29_190 ();
 sg13g2_decap_8 FILLER_29_197 ();
 sg13g2_decap_8 FILLER_29_204 ();
 sg13g2_decap_4 FILLER_29_211 ();
 sg13g2_fill_1 FILLER_29_215 ();
 sg13g2_fill_1 FILLER_29_230 ();
 sg13g2_fill_1 FILLER_29_264 ();
 sg13g2_decap_8 FILLER_29_278 ();
 sg13g2_decap_4 FILLER_29_285 ();
 sg13g2_fill_1 FILLER_29_289 ();
 sg13g2_fill_2 FILLER_29_308 ();
 sg13g2_fill_1 FILLER_29_310 ();
 sg13g2_decap_8 FILLER_29_349 ();
 sg13g2_decap_8 FILLER_29_356 ();
 sg13g2_fill_1 FILLER_29_363 ();
 sg13g2_fill_1 FILLER_29_372 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_fill_2 FILLER_30_35 ();
 sg13g2_fill_1 FILLER_30_37 ();
 sg13g2_fill_2 FILLER_30_81 ();
 sg13g2_fill_1 FILLER_30_83 ();
 sg13g2_fill_1 FILLER_30_110 ();
 sg13g2_fill_2 FILLER_30_121 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_fill_2 FILLER_30_133 ();
 sg13g2_fill_2 FILLER_30_161 ();
 sg13g2_fill_1 FILLER_30_163 ();
 sg13g2_fill_2 FILLER_30_186 ();
 sg13g2_fill_1 FILLER_30_188 ();
 sg13g2_fill_1 FILLER_30_215 ();
 sg13g2_fill_2 FILLER_30_220 ();
 sg13g2_fill_1 FILLER_30_222 ();
 sg13g2_decap_4 FILLER_30_227 ();
 sg13g2_fill_1 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_235 ();
 sg13g2_fill_1 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_285 ();
 sg13g2_decap_8 FILLER_30_292 ();
 sg13g2_decap_4 FILLER_30_299 ();
 sg13g2_fill_1 FILLER_30_320 ();
 sg13g2_fill_1 FILLER_30_325 ();
 sg13g2_decap_8 FILLER_30_334 ();
 sg13g2_decap_8 FILLER_30_341 ();
 sg13g2_decap_8 FILLER_30_348 ();
 sg13g2_decap_8 FILLER_30_355 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_15 ();
 sg13g2_fill_1 FILLER_31_70 ();
 sg13g2_fill_1 FILLER_31_84 ();
 sg13g2_fill_1 FILLER_31_145 ();
 sg13g2_decap_8 FILLER_31_150 ();
 sg13g2_decap_8 FILLER_31_157 ();
 sg13g2_fill_1 FILLER_31_164 ();
 sg13g2_decap_8 FILLER_31_181 ();
 sg13g2_decap_8 FILLER_31_188 ();
 sg13g2_decap_4 FILLER_31_195 ();
 sg13g2_fill_1 FILLER_31_199 ();
 sg13g2_fill_1 FILLER_31_204 ();
 sg13g2_fill_2 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_344 ();
 sg13g2_decap_4 FILLER_31_351 ();
 sg13g2_fill_1 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_4 FILLER_32_14 ();
 sg13g2_fill_2 FILLER_32_18 ();
 sg13g2_fill_2 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_109 ();
 sg13g2_fill_1 FILLER_32_150 ();
 sg13g2_decap_4 FILLER_32_200 ();
 sg13g2_fill_2 FILLER_32_249 ();
 sg13g2_fill_1 FILLER_32_251 ();
 sg13g2_fill_2 FILLER_32_308 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_4 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_25 ();
 sg13g2_fill_2 FILLER_33_30 ();
 sg13g2_fill_1 FILLER_33_40 ();
 sg13g2_fill_2 FILLER_33_71 ();
 sg13g2_fill_1 FILLER_33_73 ();
 sg13g2_fill_1 FILLER_33_105 ();
 sg13g2_fill_2 FILLER_33_160 ();
 sg13g2_decap_8 FILLER_33_166 ();
 sg13g2_decap_4 FILLER_33_173 ();
 sg13g2_fill_1 FILLER_33_177 ();
 sg13g2_decap_4 FILLER_33_204 ();
 sg13g2_fill_2 FILLER_33_222 ();
 sg13g2_decap_4 FILLER_33_237 ();
 sg13g2_fill_2 FILLER_33_250 ();
 sg13g2_fill_2 FILLER_33_267 ();
 sg13g2_fill_1 FILLER_33_269 ();
 sg13g2_fill_1 FILLER_33_279 ();
 sg13g2_decap_4 FILLER_33_288 ();
 sg13g2_fill_1 FILLER_33_305 ();
 sg13g2_fill_2 FILLER_33_338 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_14 ();
 sg13g2_fill_2 FILLER_34_42 ();
 sg13g2_fill_1 FILLER_34_44 ();
 sg13g2_fill_1 FILLER_34_59 ();
 sg13g2_fill_2 FILLER_34_83 ();
 sg13g2_fill_2 FILLER_34_93 ();
 sg13g2_fill_2 FILLER_34_121 ();
 sg13g2_fill_1 FILLER_34_123 ();
 sg13g2_fill_1 FILLER_34_148 ();
 sg13g2_decap_8 FILLER_34_170 ();
 sg13g2_decap_8 FILLER_34_177 ();
 sg13g2_decap_8 FILLER_34_270 ();
 sg13g2_decap_8 FILLER_34_277 ();
 sg13g2_decap_8 FILLER_34_284 ();
 sg13g2_decap_8 FILLER_34_291 ();
 sg13g2_fill_2 FILLER_34_351 ();
 sg13g2_fill_1 FILLER_34_353 ();
 sg13g2_fill_2 FILLER_34_359 ();
 sg13g2_fill_1 FILLER_34_361 ();
 sg13g2_fill_2 FILLER_34_385 ();
 sg13g2_fill_2 FILLER_34_397 ();
 sg13g2_fill_1 FILLER_34_399 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_fill_1 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_38 ();
 sg13g2_fill_1 FILLER_35_45 ();
 sg13g2_decap_8 FILLER_35_87 ();
 sg13g2_decap_8 FILLER_35_94 ();
 sg13g2_decap_8 FILLER_35_101 ();
 sg13g2_fill_1 FILLER_35_117 ();
 sg13g2_fill_2 FILLER_35_123 ();
 sg13g2_fill_1 FILLER_35_125 ();
 sg13g2_fill_1 FILLER_35_131 ();
 sg13g2_fill_2 FILLER_35_146 ();
 sg13g2_fill_2 FILLER_35_152 ();
 sg13g2_decap_8 FILLER_35_180 ();
 sg13g2_fill_2 FILLER_35_219 ();
 sg13g2_decap_4 FILLER_35_243 ();
 sg13g2_decap_8 FILLER_35_251 ();
 sg13g2_decap_8 FILLER_35_258 ();
 sg13g2_decap_8 FILLER_35_265 ();
 sg13g2_decap_8 FILLER_35_272 ();
 sg13g2_decap_8 FILLER_35_279 ();
 sg13g2_fill_1 FILLER_35_286 ();
 sg13g2_fill_1 FILLER_35_295 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_4 FILLER_35_308 ();
 sg13g2_fill_1 FILLER_35_312 ();
 sg13g2_decap_8 FILLER_35_317 ();
 sg13g2_decap_8 FILLER_35_328 ();
 sg13g2_fill_2 FILLER_35_343 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_fill_2 FILLER_35_350 ();
 sg13g2_fill_1 FILLER_35_352 ();
 sg13g2_fill_2 FILLER_35_377 ();
 sg13g2_decap_8 FILLER_36_30 ();
 sg13g2_decap_8 FILLER_36_151 ();
 sg13g2_decap_8 FILLER_36_158 ();
 sg13g2_decap_4 FILLER_36_196 ();
 sg13g2_decap_4 FILLER_36_223 ();
 sg13g2_fill_1 FILLER_36_227 ();
 sg13g2_fill_1 FILLER_36_232 ();
 sg13g2_decap_8 FILLER_36_237 ();
 sg13g2_decap_8 FILLER_36_244 ();
 sg13g2_decap_8 FILLER_36_251 ();
 sg13g2_decap_4 FILLER_36_258 ();
 sg13g2_fill_1 FILLER_36_262 ();
 sg13g2_fill_2 FILLER_36_273 ();
 sg13g2_fill_1 FILLER_36_275 ();
 sg13g2_decap_8 FILLER_36_310 ();
 sg13g2_decap_8 FILLER_36_317 ();
 sg13g2_decap_4 FILLER_36_324 ();
 sg13g2_fill_1 FILLER_36_328 ();
 sg13g2_fill_2 FILLER_36_377 ();
 sg13g2_fill_1 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_37 ();
 sg13g2_fill_1 FILLER_37_39 ();
 sg13g2_fill_2 FILLER_37_44 ();
 sg13g2_decap_8 FILLER_37_129 ();
 sg13g2_decap_4 FILLER_37_136 ();
 sg13g2_fill_1 FILLER_37_140 ();
 sg13g2_fill_1 FILLER_37_167 ();
 sg13g2_decap_8 FILLER_37_220 ();
 sg13g2_decap_8 FILLER_37_227 ();
 sg13g2_fill_2 FILLER_37_234 ();
 sg13g2_fill_1 FILLER_37_236 ();
 sg13g2_fill_2 FILLER_37_253 ();
 sg13g2_decap_4 FILLER_37_290 ();
 sg13g2_decap_4 FILLER_37_304 ();
 sg13g2_fill_1 FILLER_37_318 ();
 sg13g2_fill_2 FILLER_37_327 ();
 sg13g2_fill_2 FILLER_37_378 ();
 sg13g2_fill_1 FILLER_37_380 ();
 sg13g2_fill_2 FILLER_37_395 ();
 sg13g2_fill_1 FILLER_37_397 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_7 ();
 sg13g2_fill_2 FILLER_38_88 ();
 sg13g2_fill_1 FILLER_38_90 ();
 sg13g2_fill_1 FILLER_38_125 ();
 sg13g2_fill_1 FILLER_38_191 ();
 sg13g2_fill_1 FILLER_38_197 ();
 sg13g2_fill_2 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_4 FILLER_38_224 ();
 sg13g2_fill_1 FILLER_38_315 ();
 sg13g2_fill_2 FILLER_38_326 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_fill_1 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_365 ();
 sg13g2_fill_2 FILLER_38_381 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_4 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_30 ();
 sg13g2_decap_4 FILLER_39_37 ();
 sg13g2_fill_1 FILLER_39_41 ();
 sg13g2_fill_1 FILLER_39_89 ();
 sg13g2_decap_8 FILLER_39_96 ();
 sg13g2_fill_2 FILLER_39_103 ();
 sg13g2_fill_1 FILLER_39_105 ();
 sg13g2_decap_4 FILLER_39_111 ();
 sg13g2_fill_2 FILLER_39_115 ();
 sg13g2_fill_1 FILLER_39_133 ();
 sg13g2_fill_2 FILLER_39_154 ();
 sg13g2_decap_4 FILLER_39_186 ();
 sg13g2_fill_1 FILLER_39_203 ();
 sg13g2_fill_2 FILLER_39_250 ();
 sg13g2_fill_2 FILLER_39_260 ();
 sg13g2_decap_4 FILLER_39_307 ();
 sg13g2_fill_2 FILLER_39_311 ();
 sg13g2_decap_8 FILLER_39_321 ();
 sg13g2_decap_8 FILLER_39_328 ();
 sg13g2_decap_8 FILLER_39_354 ();
 sg13g2_fill_2 FILLER_39_361 ();
 sg13g2_fill_1 FILLER_39_363 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_fill_2 FILLER_40_52 ();
 sg13g2_fill_1 FILLER_40_54 ();
 sg13g2_fill_1 FILLER_40_127 ();
 sg13g2_fill_2 FILLER_40_165 ();
 sg13g2_fill_2 FILLER_40_172 ();
 sg13g2_fill_1 FILLER_40_174 ();
 sg13g2_fill_2 FILLER_40_210 ();
 sg13g2_fill_2 FILLER_40_234 ();
 sg13g2_fill_1 FILLER_40_236 ();
 sg13g2_decap_8 FILLER_40_249 ();
 sg13g2_decap_4 FILLER_40_256 ();
 sg13g2_fill_2 FILLER_40_270 ();
 sg13g2_fill_1 FILLER_40_272 ();
 sg13g2_fill_1 FILLER_40_287 ();
 sg13g2_decap_8 FILLER_40_292 ();
 sg13g2_decap_4 FILLER_40_299 ();
 sg13g2_fill_1 FILLER_40_334 ();
 sg13g2_decap_4 FILLER_40_376 ();
 sg13g2_fill_1 FILLER_40_389 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_4 FILLER_41_14 ();
 sg13g2_fill_2 FILLER_41_18 ();
 sg13g2_fill_1 FILLER_41_92 ();
 sg13g2_fill_1 FILLER_41_100 ();
 sg13g2_fill_1 FILLER_41_119 ();
 sg13g2_fill_2 FILLER_41_177 ();
 sg13g2_decap_8 FILLER_41_187 ();
 sg13g2_decap_4 FILLER_41_194 ();
 sg13g2_fill_2 FILLER_41_206 ();
 sg13g2_decap_4 FILLER_41_259 ();
 sg13g2_decap_8 FILLER_41_272 ();
 sg13g2_decap_4 FILLER_41_279 ();
 sg13g2_decap_4 FILLER_41_289 ();
 sg13g2_fill_2 FILLER_41_355 ();
 sg13g2_fill_1 FILLER_41_369 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_7 ();
 sg13g2_fill_1 FILLER_42_9 ();
 sg13g2_fill_1 FILLER_42_45 ();
 sg13g2_fill_1 FILLER_42_63 ();
 sg13g2_fill_2 FILLER_42_80 ();
 sg13g2_fill_2 FILLER_42_89 ();
 sg13g2_fill_2 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_198 ();
 sg13g2_decap_8 FILLER_42_205 ();
 sg13g2_fill_2 FILLER_42_212 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_fill_2 FILLER_42_231 ();
 sg13g2_fill_1 FILLER_42_259 ();
 sg13g2_decap_8 FILLER_42_281 ();
 sg13g2_fill_1 FILLER_42_318 ();
 sg13g2_fill_2 FILLER_42_328 ();
 sg13g2_fill_1 FILLER_42_343 ();
 sg13g2_fill_1 FILLER_42_360 ();
 sg13g2_fill_1 FILLER_42_382 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_34 ();
 sg13g2_fill_2 FILLER_43_89 ();
 sg13g2_fill_1 FILLER_43_91 ();
 sg13g2_fill_2 FILLER_43_97 ();
 sg13g2_fill_1 FILLER_43_99 ();
 sg13g2_fill_2 FILLER_43_136 ();
 sg13g2_fill_1 FILLER_43_138 ();
 sg13g2_decap_4 FILLER_43_208 ();
 sg13g2_fill_2 FILLER_43_221 ();
 sg13g2_decap_4 FILLER_43_236 ();
 sg13g2_fill_2 FILLER_43_252 ();
 sg13g2_fill_1 FILLER_43_286 ();
 sg13g2_fill_1 FILLER_43_315 ();
 sg13g2_fill_2 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_356 ();
 sg13g2_fill_2 FILLER_43_363 ();
 sg13g2_fill_2 FILLER_43_375 ();
 sg13g2_fill_1 FILLER_43_377 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_fill_2 FILLER_44_14 ();
 sg13g2_fill_1 FILLER_44_29 ();
 sg13g2_fill_2 FILLER_44_54 ();
 sg13g2_fill_1 FILLER_44_56 ();
 sg13g2_fill_1 FILLER_44_92 ();
 sg13g2_fill_2 FILLER_44_102 ();
 sg13g2_fill_1 FILLER_44_104 ();
 sg13g2_fill_2 FILLER_44_114 ();
 sg13g2_fill_2 FILLER_44_121 ();
 sg13g2_fill_1 FILLER_44_123 ();
 sg13g2_fill_2 FILLER_44_132 ();
 sg13g2_decap_8 FILLER_44_155 ();
 sg13g2_fill_2 FILLER_44_180 ();
 sg13g2_decap_4 FILLER_44_221 ();
 sg13g2_fill_2 FILLER_44_251 ();
 sg13g2_fill_1 FILLER_44_253 ();
 sg13g2_fill_2 FILLER_44_320 ();
 sg13g2_fill_1 FILLER_44_322 ();
 sg13g2_fill_2 FILLER_44_332 ();
 sg13g2_fill_1 FILLER_44_349 ();
 sg13g2_fill_2 FILLER_44_363 ();
 sg13g2_fill_1 FILLER_44_373 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_fill_1 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_54 ();
 sg13g2_fill_2 FILLER_45_61 ();
 sg13g2_decap_8 FILLER_45_165 ();
 sg13g2_fill_1 FILLER_45_176 ();
 sg13g2_fill_2 FILLER_45_190 ();
 sg13g2_fill_1 FILLER_45_225 ();
 sg13g2_decap_8 FILLER_45_248 ();
 sg13g2_fill_1 FILLER_45_255 ();
 sg13g2_decap_4 FILLER_45_269 ();
 sg13g2_fill_2 FILLER_45_278 ();
 sg13g2_fill_1 FILLER_45_280 ();
 sg13g2_decap_8 FILLER_45_285 ();
 sg13g2_decap_4 FILLER_45_292 ();
 sg13g2_decap_8 FILLER_45_331 ();
 sg13g2_fill_1 FILLER_45_338 ();
 sg13g2_fill_1 FILLER_45_343 ();
 sg13g2_fill_2 FILLER_45_380 ();
 sg13g2_fill_1 FILLER_45_382 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_4 FILLER_46_21 ();
 sg13g2_fill_2 FILLER_46_101 ();
 sg13g2_fill_1 FILLER_46_103 ();
 sg13g2_fill_2 FILLER_46_130 ();
 sg13g2_fill_1 FILLER_46_132 ();
 sg13g2_fill_1 FILLER_46_173 ();
 sg13g2_decap_8 FILLER_46_263 ();
 sg13g2_decap_4 FILLER_46_270 ();
 sg13g2_fill_2 FILLER_46_274 ();
 sg13g2_decap_8 FILLER_46_281 ();
 sg13g2_fill_1 FILLER_46_288 ();
 sg13g2_decap_4 FILLER_46_294 ();
 sg13g2_fill_1 FILLER_46_298 ();
 sg13g2_fill_1 FILLER_46_307 ();
 sg13g2_fill_2 FILLER_46_360 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_fill_2 FILLER_47_21 ();
 sg13g2_fill_1 FILLER_47_23 ();
 sg13g2_fill_2 FILLER_47_74 ();
 sg13g2_fill_2 FILLER_47_88 ();
 sg13g2_fill_2 FILLER_47_100 ();
 sg13g2_fill_1 FILLER_47_102 ();
 sg13g2_fill_2 FILLER_47_155 ();
 sg13g2_fill_1 FILLER_47_212 ();
 sg13g2_decap_8 FILLER_47_234 ();
 sg13g2_decap_4 FILLER_47_241 ();
 sg13g2_decap_4 FILLER_47_259 ();
 sg13g2_fill_2 FILLER_47_276 ();
 sg13g2_fill_1 FILLER_47_288 ();
 sg13g2_decap_4 FILLER_47_299 ();
 sg13g2_decap_8 FILLER_47_312 ();
 sg13g2_decap_8 FILLER_47_355 ();
 sg13g2_fill_2 FILLER_47_362 ();
 sg13g2_fill_1 FILLER_47_364 ();
 sg13g2_fill_2 FILLER_47_369 ();
 sg13g2_fill_1 FILLER_47_371 ();
 sg13g2_fill_2 FILLER_47_407 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_4 FILLER_48_21 ();
 sg13g2_fill_1 FILLER_48_51 ();
 sg13g2_decap_8 FILLER_48_83 ();
 sg13g2_decap_8 FILLER_48_90 ();
 sg13g2_decap_4 FILLER_48_97 ();
 sg13g2_fill_2 FILLER_48_105 ();
 sg13g2_fill_1 FILLER_48_138 ();
 sg13g2_fill_2 FILLER_48_183 ();
 sg13g2_fill_1 FILLER_48_185 ();
 sg13g2_fill_2 FILLER_48_191 ();
 sg13g2_fill_1 FILLER_48_193 ();
 sg13g2_fill_2 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_219 ();
 sg13g2_fill_1 FILLER_48_226 ();
 sg13g2_decap_4 FILLER_48_239 ();
 sg13g2_fill_2 FILLER_48_269 ();
 sg13g2_fill_1 FILLER_48_271 ();
 sg13g2_decap_4 FILLER_48_278 ();
 sg13g2_fill_2 FILLER_48_302 ();
 sg13g2_fill_2 FILLER_48_363 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_4 FILLER_49_28 ();
 sg13g2_fill_2 FILLER_49_32 ();
 sg13g2_fill_1 FILLER_49_43 ();
 sg13g2_fill_2 FILLER_49_70 ();
 sg13g2_decap_4 FILLER_49_91 ();
 sg13g2_fill_2 FILLER_49_95 ();
 sg13g2_fill_2 FILLER_49_105 ();
 sg13g2_fill_1 FILLER_49_107 ();
 sg13g2_fill_2 FILLER_49_138 ();
 sg13g2_decap_8 FILLER_49_144 ();
 sg13g2_fill_2 FILLER_49_151 ();
 sg13g2_fill_1 FILLER_49_153 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_4 FILLER_49_196 ();
 sg13g2_fill_1 FILLER_49_200 ();
 sg13g2_fill_2 FILLER_49_227 ();
 sg13g2_fill_2 FILLER_49_238 ();
 sg13g2_fill_1 FILLER_49_240 ();
 sg13g2_decap_4 FILLER_49_250 ();
 sg13g2_decap_8 FILLER_49_258 ();
 sg13g2_decap_4 FILLER_49_265 ();
 sg13g2_fill_1 FILLER_49_269 ();
 sg13g2_fill_1 FILLER_49_305 ();
 sg13g2_fill_2 FILLER_49_398 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_4 FILLER_50_21 ();
 sg13g2_fill_2 FILLER_50_25 ();
 sg13g2_fill_2 FILLER_50_36 ();
 sg13g2_fill_1 FILLER_50_38 ();
 sg13g2_fill_1 FILLER_50_73 ();
 sg13g2_fill_2 FILLER_50_113 ();
 sg13g2_fill_2 FILLER_50_215 ();
 sg13g2_fill_1 FILLER_50_217 ();
 sg13g2_fill_1 FILLER_50_248 ();
 sg13g2_fill_2 FILLER_50_275 ();
 sg13g2_decap_8 FILLER_50_306 ();
 sg13g2_decap_8 FILLER_50_313 ();
 sg13g2_fill_2 FILLER_50_320 ();
 sg13g2_fill_1 FILLER_50_322 ();
 sg13g2_fill_2 FILLER_50_372 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_4 FILLER_51_14 ();
 sg13g2_fill_2 FILLER_51_54 ();
 sg13g2_fill_1 FILLER_51_56 ();
 sg13g2_fill_2 FILLER_51_109 ();
 sg13g2_fill_1 FILLER_51_111 ();
 sg13g2_fill_1 FILLER_51_175 ();
 sg13g2_decap_4 FILLER_51_226 ();
 sg13g2_fill_2 FILLER_51_230 ();
 sg13g2_fill_2 FILLER_51_258 ();
 sg13g2_decap_8 FILLER_51_264 ();
 sg13g2_decap_4 FILLER_51_271 ();
 sg13g2_fill_1 FILLER_51_275 ();
 sg13g2_decap_4 FILLER_51_295 ();
 sg13g2_fill_2 FILLER_51_299 ();
 sg13g2_fill_1 FILLER_51_321 ();
 sg13g2_decap_8 FILLER_51_332 ();
 sg13g2_fill_1 FILLER_51_343 ();
 sg13g2_fill_1 FILLER_51_378 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_fill_1 FILLER_52_28 ();
 sg13g2_fill_1 FILLER_52_33 ();
 sg13g2_fill_1 FILLER_52_81 ();
 sg13g2_fill_1 FILLER_52_96 ();
 sg13g2_fill_2 FILLER_52_117 ();
 sg13g2_fill_1 FILLER_52_119 ();
 sg13g2_fill_2 FILLER_52_134 ();
 sg13g2_fill_1 FILLER_52_136 ();
 sg13g2_fill_1 FILLER_52_181 ();
 sg13g2_decap_8 FILLER_52_230 ();
 sg13g2_fill_2 FILLER_52_255 ();
 sg13g2_decap_4 FILLER_52_277 ();
 sg13g2_fill_1 FILLER_52_281 ();
 sg13g2_fill_2 FILLER_52_347 ();
 sg13g2_fill_1 FILLER_52_354 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_4 FILLER_53_35 ();
 sg13g2_fill_1 FILLER_53_116 ();
 sg13g2_fill_2 FILLER_53_138 ();
 sg13g2_fill_2 FILLER_53_176 ();
 sg13g2_fill_1 FILLER_53_178 ();
 sg13g2_decap_4 FILLER_53_191 ();
 sg13g2_fill_1 FILLER_53_212 ();
 sg13g2_fill_2 FILLER_53_222 ();
 sg13g2_fill_1 FILLER_53_224 ();
 sg13g2_decap_8 FILLER_53_287 ();
 sg13g2_fill_2 FILLER_53_294 ();
 sg13g2_fill_1 FILLER_53_322 ();
 sg13g2_fill_1 FILLER_53_332 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_4 FILLER_54_42 ();
 sg13g2_fill_2 FILLER_54_46 ();
 sg13g2_fill_2 FILLER_54_62 ();
 sg13g2_fill_1 FILLER_54_64 ();
 sg13g2_fill_2 FILLER_54_91 ();
 sg13g2_fill_2 FILLER_54_125 ();
 sg13g2_fill_1 FILLER_54_127 ();
 sg13g2_fill_2 FILLER_54_146 ();
 sg13g2_fill_1 FILLER_54_175 ();
 sg13g2_decap_8 FILLER_54_186 ();
 sg13g2_fill_2 FILLER_54_193 ();
 sg13g2_decap_8 FILLER_54_204 ();
 sg13g2_decap_8 FILLER_54_211 ();
 sg13g2_decap_8 FILLER_54_218 ();
 sg13g2_decap_8 FILLER_54_225 ();
 sg13g2_fill_2 FILLER_54_232 ();
 sg13g2_fill_1 FILLER_54_234 ();
 sg13g2_decap_8 FILLER_54_248 ();
 sg13g2_decap_4 FILLER_54_255 ();
 sg13g2_fill_2 FILLER_54_259 ();
 sg13g2_fill_2 FILLER_54_285 ();
 sg13g2_fill_1 FILLER_54_295 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_fill_2 FILLER_55_42 ();
 sg13g2_fill_1 FILLER_55_44 ();
 sg13g2_fill_1 FILLER_55_106 ();
 sg13g2_fill_2 FILLER_55_127 ();
 sg13g2_decap_4 FILLER_55_158 ();
 sg13g2_fill_2 FILLER_55_162 ();
 sg13g2_fill_2 FILLER_55_169 ();
 sg13g2_decap_8 FILLER_55_201 ();
 sg13g2_decap_4 FILLER_55_208 ();
 sg13g2_fill_2 FILLER_55_212 ();
 sg13g2_fill_1 FILLER_55_228 ();
 sg13g2_fill_2 FILLER_55_238 ();
 sg13g2_decap_4 FILLER_55_245 ();
 sg13g2_fill_1 FILLER_55_249 ();
 sg13g2_decap_8 FILLER_55_257 ();
 sg13g2_decap_4 FILLER_55_264 ();
 sg13g2_decap_4 FILLER_55_282 ();
 sg13g2_fill_1 FILLER_55_349 ();
 sg13g2_fill_2 FILLER_55_380 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_fill_2 FILLER_56_87 ();
 sg13g2_fill_2 FILLER_56_108 ();
 sg13g2_fill_2 FILLER_56_133 ();
 sg13g2_decap_4 FILLER_56_149 ();
 sg13g2_fill_1 FILLER_56_153 ();
 sg13g2_fill_1 FILLER_56_272 ();
 sg13g2_decap_4 FILLER_56_290 ();
 sg13g2_fill_1 FILLER_56_294 ();
 sg13g2_decap_4 FILLER_56_308 ();
 sg13g2_fill_2 FILLER_56_327 ();
 sg13g2_fill_1 FILLER_56_355 ();
 sg13g2_decap_4 FILLER_56_373 ();
 sg13g2_fill_1 FILLER_56_377 ();
 sg13g2_decap_8 FILLER_56_382 ();
 sg13g2_fill_2 FILLER_56_389 ();
 sg13g2_fill_1 FILLER_56_391 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_fill_2 FILLER_57_60 ();
 sg13g2_fill_1 FILLER_57_62 ();
 sg13g2_fill_2 FILLER_57_72 ();
 sg13g2_fill_2 FILLER_57_82 ();
 sg13g2_fill_1 FILLER_57_136 ();
 sg13g2_fill_2 FILLER_57_141 ();
 sg13g2_fill_1 FILLER_57_143 ();
 sg13g2_decap_4 FILLER_57_160 ();
 sg13g2_fill_1 FILLER_57_164 ();
 sg13g2_fill_2 FILLER_57_169 ();
 sg13g2_fill_1 FILLER_57_223 ();
 sg13g2_fill_1 FILLER_57_307 ();
 sg13g2_fill_1 FILLER_57_339 ();
 sg13g2_fill_2 FILLER_57_344 ();
 sg13g2_decap_8 FILLER_57_372 ();
 sg13g2_decap_8 FILLER_57_379 ();
 sg13g2_decap_8 FILLER_57_386 ();
 sg13g2_fill_2 FILLER_57_393 ();
 sg13g2_decap_8 FILLER_57_399 ();
 sg13g2_fill_2 FILLER_57_406 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_fill_1 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_68 ();
 sg13g2_decap_4 FILLER_58_75 ();
 sg13g2_fill_2 FILLER_58_91 ();
 sg13g2_fill_1 FILLER_58_157 ();
 sg13g2_fill_2 FILLER_58_214 ();
 sg13g2_fill_1 FILLER_58_216 ();
 sg13g2_fill_2 FILLER_58_270 ();
 sg13g2_fill_2 FILLER_58_290 ();
 sg13g2_fill_2 FILLER_58_296 ();
 sg13g2_decap_4 FILLER_58_334 ();
 sg13g2_decap_8 FILLER_58_352 ();
 sg13g2_decap_8 FILLER_58_359 ();
 sg13g2_decap_4 FILLER_58_366 ();
 sg13g2_fill_1 FILLER_58_370 ();
 sg13g2_fill_2 FILLER_58_381 ();
 sg13g2_fill_2 FILLER_58_406 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_fill_1 FILLER_59_132 ();
 sg13g2_decap_4 FILLER_59_163 ();
 sg13g2_fill_2 FILLER_59_167 ();
 sg13g2_fill_2 FILLER_59_173 ();
 sg13g2_fill_1 FILLER_59_193 ();
 sg13g2_decap_4 FILLER_59_234 ();
 sg13g2_fill_2 FILLER_59_265 ();
 sg13g2_fill_2 FILLER_59_272 ();
 sg13g2_decap_4 FILLER_59_282 ();
 sg13g2_fill_1 FILLER_59_286 ();
 sg13g2_fill_1 FILLER_59_292 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_4 FILLER_60_49 ();
 sg13g2_decap_4 FILLER_60_112 ();
 sg13g2_fill_2 FILLER_60_142 ();
 sg13g2_fill_2 FILLER_60_148 ();
 sg13g2_decap_8 FILLER_60_169 ();
 sg13g2_decap_4 FILLER_60_176 ();
 sg13g2_decap_8 FILLER_60_224 ();
 sg13g2_decap_8 FILLER_60_231 ();
 sg13g2_decap_8 FILLER_60_242 ();
 sg13g2_decap_4 FILLER_60_249 ();
 sg13g2_fill_2 FILLER_60_253 ();
 sg13g2_fill_2 FILLER_60_267 ();
 sg13g2_decap_4 FILLER_60_282 ();
 sg13g2_fill_1 FILLER_60_346 ();
 sg13g2_fill_1 FILLER_60_366 ();
 sg13g2_fill_2 FILLER_60_388 ();
 sg13g2_fill_1 FILLER_60_390 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_4 FILLER_61_49 ();
 sg13g2_fill_1 FILLER_61_53 ();
 sg13g2_fill_2 FILLER_61_116 ();
 sg13g2_fill_1 FILLER_61_118 ();
 sg13g2_decap_8 FILLER_61_123 ();
 sg13g2_decap_4 FILLER_61_130 ();
 sg13g2_fill_2 FILLER_61_134 ();
 sg13g2_decap_4 FILLER_61_145 ();
 sg13g2_decap_8 FILLER_61_184 ();
 sg13g2_decap_4 FILLER_61_195 ();
 sg13g2_fill_2 FILLER_61_199 ();
 sg13g2_fill_1 FILLER_61_227 ();
 sg13g2_fill_1 FILLER_61_242 ();
 sg13g2_fill_2 FILLER_61_248 ();
 sg13g2_fill_1 FILLER_61_250 ();
 sg13g2_decap_4 FILLER_61_254 ();
 sg13g2_fill_1 FILLER_61_258 ();
 sg13g2_fill_1 FILLER_61_294 ();
 sg13g2_decap_8 FILLER_61_330 ();
 sg13g2_decap_4 FILLER_61_337 ();
 sg13g2_fill_2 FILLER_61_368 ();
 sg13g2_fill_2 FILLER_61_380 ();
 sg13g2_fill_1 FILLER_61_387 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_4 FILLER_62_56 ();
 sg13g2_fill_2 FILLER_62_87 ();
 sg13g2_fill_2 FILLER_62_98 ();
 sg13g2_fill_1 FILLER_62_139 ();
 sg13g2_fill_1 FILLER_62_149 ();
 sg13g2_fill_2 FILLER_62_306 ();
 sg13g2_fill_1 FILLER_62_308 ();
 sg13g2_fill_2 FILLER_62_314 ();
 sg13g2_decap_8 FILLER_62_342 ();
 sg13g2_fill_1 FILLER_62_386 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_fill_2 FILLER_63_101 ();
 sg13g2_fill_1 FILLER_63_103 ();
 sg13g2_fill_2 FILLER_63_156 ();
 sg13g2_fill_1 FILLER_63_158 ();
 sg13g2_fill_2 FILLER_63_173 ();
 sg13g2_fill_1 FILLER_63_225 ();
 sg13g2_fill_2 FILLER_63_300 ();
 sg13g2_fill_2 FILLER_63_319 ();
 sg13g2_decap_8 FILLER_63_347 ();
 sg13g2_fill_2 FILLER_63_354 ();
 sg13g2_fill_2 FILLER_63_360 ();
 sg13g2_fill_1 FILLER_63_362 ();
 sg13g2_fill_2 FILLER_63_367 ();
 sg13g2_fill_1 FILLER_63_369 ();
 sg13g2_fill_1 FILLER_63_379 ();
 sg13g2_fill_1 FILLER_63_389 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_fill_2 FILLER_64_88 ();
 sg13g2_fill_1 FILLER_64_122 ();
 sg13g2_fill_2 FILLER_64_133 ();
 sg13g2_fill_1 FILLER_64_135 ();
 sg13g2_fill_2 FILLER_64_189 ();
 sg13g2_fill_1 FILLER_64_191 ();
 sg13g2_decap_8 FILLER_64_213 ();
 sg13g2_fill_2 FILLER_64_220 ();
 sg13g2_decap_8 FILLER_64_226 ();
 sg13g2_decap_8 FILLER_64_233 ();
 sg13g2_decap_8 FILLER_64_240 ();
 sg13g2_decap_8 FILLER_64_247 ();
 sg13g2_fill_2 FILLER_64_254 ();
 sg13g2_fill_2 FILLER_64_265 ();
 sg13g2_decap_4 FILLER_64_334 ();
 sg13g2_decap_8 FILLER_64_342 ();
 sg13g2_fill_1 FILLER_64_349 ();
 sg13g2_decap_8 FILLER_64_355 ();
 sg13g2_decap_8 FILLER_64_362 ();
 sg13g2_fill_1 FILLER_64_369 ();
 sg13g2_fill_2 FILLER_64_385 ();
 sg13g2_decap_4 FILLER_64_391 ();
 sg13g2_fill_2 FILLER_64_395 ();
 sg13g2_decap_8 FILLER_64_402 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_4 FILLER_65_56 ();
 sg13g2_fill_2 FILLER_65_60 ();
 sg13g2_fill_2 FILLER_65_129 ();
 sg13g2_fill_1 FILLER_65_141 ();
 sg13g2_fill_1 FILLER_65_175 ();
 sg13g2_fill_1 FILLER_65_209 ();
 sg13g2_fill_1 FILLER_65_225 ();
 sg13g2_decap_8 FILLER_65_239 ();
 sg13g2_fill_2 FILLER_65_246 ();
 sg13g2_fill_1 FILLER_65_253 ();
 sg13g2_fill_1 FILLER_65_270 ();
 sg13g2_fill_2 FILLER_65_324 ();
 sg13g2_fill_1 FILLER_65_326 ();
 sg13g2_decap_4 FILLER_65_356 ();
 sg13g2_decap_8 FILLER_65_378 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_fill_1 FILLER_66_49 ();
 sg13g2_fill_1 FILLER_66_112 ();
 sg13g2_fill_2 FILLER_66_181 ();
 sg13g2_fill_2 FILLER_66_246 ();
 sg13g2_fill_2 FILLER_66_279 ();
 sg13g2_fill_1 FILLER_66_303 ();
 sg13g2_fill_2 FILLER_66_360 ();
 sg13g2_fill_1 FILLER_66_366 ();
 sg13g2_decap_4 FILLER_66_375 ();
 sg13g2_fill_2 FILLER_66_379 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_fill_2 FILLER_67_63 ();
 sg13g2_fill_1 FILLER_67_65 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_4 FILLER_67_94 ();
 sg13g2_fill_1 FILLER_67_98 ();
 sg13g2_fill_2 FILLER_67_129 ();
 sg13g2_fill_1 FILLER_67_166 ();
 sg13g2_fill_1 FILLER_67_190 ();
 sg13g2_fill_2 FILLER_67_208 ();
 sg13g2_fill_1 FILLER_67_250 ();
 sg13g2_fill_1 FILLER_67_275 ();
 sg13g2_decap_8 FILLER_67_336 ();
 sg13g2_decap_4 FILLER_67_343 ();
 sg13g2_fill_2 FILLER_67_347 ();
 sg13g2_fill_2 FILLER_67_371 ();
 sg13g2_decap_8 FILLER_67_382 ();
 sg13g2_fill_2 FILLER_67_389 ();
 sg13g2_fill_1 FILLER_67_391 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_fill_2 FILLER_68_70 ();
 sg13g2_fill_1 FILLER_68_72 ();
 sg13g2_fill_2 FILLER_68_83 ();
 sg13g2_fill_1 FILLER_68_85 ();
 sg13g2_fill_2 FILLER_68_117 ();
 sg13g2_fill_2 FILLER_68_166 ();
 sg13g2_decap_4 FILLER_68_192 ();
 sg13g2_fill_2 FILLER_68_212 ();
 sg13g2_fill_1 FILLER_68_214 ();
 sg13g2_fill_2 FILLER_68_250 ();
 sg13g2_fill_1 FILLER_68_270 ();
 sg13g2_fill_2 FILLER_68_311 ();
 sg13g2_fill_2 FILLER_68_367 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_fill_2 FILLER_69_101 ();
 sg13g2_decap_8 FILLER_69_142 ();
 sg13g2_decap_4 FILLER_69_149 ();
 sg13g2_fill_2 FILLER_69_184 ();
 sg13g2_decap_4 FILLER_69_196 ();
 sg13g2_fill_2 FILLER_69_231 ();
 sg13g2_fill_1 FILLER_69_233 ();
 sg13g2_fill_2 FILLER_69_294 ();
 sg13g2_fill_1 FILLER_69_296 ();
 sg13g2_decap_8 FILLER_69_306 ();
 sg13g2_decap_8 FILLER_69_313 ();
 sg13g2_fill_2 FILLER_69_328 ();
 sg13g2_fill_1 FILLER_69_330 ();
 sg13g2_fill_2 FILLER_69_362 ();
 sg13g2_fill_1 FILLER_69_364 ();
 sg13g2_fill_2 FILLER_69_384 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_fill_2 FILLER_70_76 ();
 sg13g2_fill_1 FILLER_70_104 ();
 sg13g2_fill_1 FILLER_70_131 ();
 sg13g2_fill_1 FILLER_70_151 ();
 sg13g2_fill_2 FILLER_70_194 ();
 sg13g2_fill_1 FILLER_70_196 ();
 sg13g2_decap_4 FILLER_70_202 ();
 sg13g2_fill_1 FILLER_70_206 ();
 sg13g2_fill_2 FILLER_70_215 ();
 sg13g2_decap_8 FILLER_70_226 ();
 sg13g2_decap_8 FILLER_70_233 ();
 sg13g2_decap_4 FILLER_70_240 ();
 sg13g2_fill_2 FILLER_70_244 ();
 sg13g2_fill_1 FILLER_70_260 ();
 sg13g2_fill_2 FILLER_70_271 ();
 sg13g2_fill_1 FILLER_70_273 ();
 sg13g2_fill_2 FILLER_70_367 ();
 sg13g2_fill_1 FILLER_70_369 ();
 sg13g2_fill_2 FILLER_70_407 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_4 FILLER_71_56 ();
 sg13g2_fill_2 FILLER_71_86 ();
 sg13g2_fill_2 FILLER_71_110 ();
 sg13g2_fill_2 FILLER_71_209 ();
 sg13g2_decap_8 FILLER_71_221 ();
 sg13g2_fill_1 FILLER_71_273 ();
 sg13g2_fill_2 FILLER_71_279 ();
 sg13g2_fill_1 FILLER_71_281 ();
 sg13g2_decap_8 FILLER_71_336 ();
 sg13g2_decap_4 FILLER_71_343 ();
 sg13g2_fill_2 FILLER_71_372 ();
 sg13g2_decap_4 FILLER_71_403 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_fill_1 FILLER_72_84 ();
 sg13g2_fill_1 FILLER_72_115 ();
 sg13g2_fill_2 FILLER_72_145 ();
 sg13g2_fill_2 FILLER_72_219 ();
 sg13g2_fill_1 FILLER_72_221 ();
 sg13g2_fill_2 FILLER_72_248 ();
 sg13g2_decap_4 FILLER_72_285 ();
 sg13g2_fill_1 FILLER_72_289 ();
 sg13g2_fill_1 FILLER_72_307 ();
 sg13g2_fill_1 FILLER_72_322 ();
 sg13g2_fill_2 FILLER_72_328 ();
 sg13g2_fill_1 FILLER_72_330 ();
 sg13g2_decap_8 FILLER_72_334 ();
 sg13g2_decap_8 FILLER_72_341 ();
 sg13g2_fill_2 FILLER_72_348 ();
 sg13g2_fill_1 FILLER_72_350 ();
 sg13g2_fill_1 FILLER_72_356 ();
 sg13g2_decap_4 FILLER_72_362 ();
 sg13g2_fill_2 FILLER_72_370 ();
 sg13g2_fill_2 FILLER_72_377 ();
 sg13g2_fill_1 FILLER_72_379 ();
 sg13g2_fill_1 FILLER_72_385 ();
 sg13g2_decap_8 FILLER_72_401 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_fill_2 FILLER_73_91 ();
 sg13g2_fill_1 FILLER_73_93 ();
 sg13g2_fill_1 FILLER_73_103 ();
 sg13g2_fill_1 FILLER_73_139 ();
 sg13g2_fill_1 FILLER_73_189 ();
 sg13g2_fill_1 FILLER_73_208 ();
 sg13g2_fill_2 FILLER_73_275 ();
 sg13g2_fill_1 FILLER_73_277 ();
 sg13g2_fill_2 FILLER_73_283 ();
 sg13g2_fill_1 FILLER_73_285 ();
 sg13g2_fill_2 FILLER_73_300 ();
 sg13g2_decap_8 FILLER_73_341 ();
 sg13g2_decap_8 FILLER_73_355 ();
 sg13g2_fill_1 FILLER_73_362 ();
 sg13g2_decap_4 FILLER_73_368 ();
 sg13g2_fill_2 FILLER_73_382 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_fill_1 FILLER_74_98 ();
 sg13g2_decap_4 FILLER_74_103 ();
 sg13g2_fill_2 FILLER_74_107 ();
 sg13g2_fill_1 FILLER_74_122 ();
 sg13g2_fill_1 FILLER_74_163 ();
 sg13g2_fill_2 FILLER_74_200 ();
 sg13g2_fill_2 FILLER_74_264 ();
 sg13g2_fill_1 FILLER_74_266 ();
 sg13g2_fill_1 FILLER_74_298 ();
 sg13g2_fill_1 FILLER_74_342 ();
 sg13g2_fill_1 FILLER_74_356 ();
 sg13g2_fill_2 FILLER_74_374 ();
 sg13g2_fill_2 FILLER_74_406 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_fill_2 FILLER_75_105 ();
 sg13g2_fill_2 FILLER_75_143 ();
 sg13g2_fill_1 FILLER_75_145 ();
 sg13g2_fill_2 FILLER_75_169 ();
 sg13g2_decap_8 FILLER_75_187 ();
 sg13g2_decap_8 FILLER_75_194 ();
 sg13g2_fill_2 FILLER_75_201 ();
 sg13g2_fill_2 FILLER_75_230 ();
 sg13g2_decap_4 FILLER_75_241 ();
 sg13g2_decap_4 FILLER_75_250 ();
 sg13g2_fill_2 FILLER_75_254 ();
 sg13g2_fill_1 FILLER_75_381 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_fill_1 FILLER_76_98 ();
 sg13g2_fill_1 FILLER_76_107 ();
 sg13g2_fill_1 FILLER_76_148 ();
 sg13g2_fill_1 FILLER_76_162 ();
 sg13g2_decap_4 FILLER_76_181 ();
 sg13g2_fill_2 FILLER_76_185 ();
 sg13g2_fill_2 FILLER_76_274 ();
 sg13g2_fill_1 FILLER_76_276 ();
 sg13g2_fill_2 FILLER_76_291 ();
 sg13g2_fill_2 FILLER_76_303 ();
 sg13g2_fill_2 FILLER_76_388 ();
 sg13g2_fill_2 FILLER_76_396 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_4 FILLER_77_91 ();
 sg13g2_fill_2 FILLER_77_176 ();
 sg13g2_fill_1 FILLER_77_178 ();
 sg13g2_fill_2 FILLER_77_209 ();
 sg13g2_fill_1 FILLER_77_211 ();
 sg13g2_fill_2 FILLER_77_225 ();
 sg13g2_fill_2 FILLER_77_267 ();
 sg13g2_fill_1 FILLER_77_269 ();
 sg13g2_fill_1 FILLER_77_281 ();
 sg13g2_fill_1 FILLER_77_291 ();
 sg13g2_fill_1 FILLER_77_327 ();
 sg13g2_fill_2 FILLER_77_349 ();
 sg13g2_fill_1 FILLER_77_351 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_4 FILLER_78_105 ();
 sg13g2_fill_1 FILLER_78_109 ();
 sg13g2_fill_2 FILLER_78_157 ();
 sg13g2_fill_2 FILLER_78_194 ();
 sg13g2_fill_1 FILLER_78_196 ();
 sg13g2_fill_1 FILLER_78_258 ();
 sg13g2_fill_1 FILLER_78_311 ();
 sg13g2_fill_1 FILLER_78_366 ();
 sg13g2_fill_2 FILLER_78_377 ();
 sg13g2_fill_1 FILLER_78_379 ();
 sg13g2_fill_2 FILLER_78_406 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_4 FILLER_79_98 ();
 sg13g2_fill_2 FILLER_79_102 ();
 sg13g2_fill_1 FILLER_79_108 ();
 sg13g2_fill_2 FILLER_79_126 ();
 sg13g2_fill_1 FILLER_79_128 ();
 sg13g2_fill_2 FILLER_79_194 ();
 sg13g2_fill_1 FILLER_79_196 ();
 sg13g2_fill_1 FILLER_79_231 ();
 sg13g2_fill_1 FILLER_79_237 ();
 sg13g2_fill_2 FILLER_79_369 ();
 sg13g2_fill_1 FILLER_79_371 ();
 sg13g2_fill_1 FILLER_79_381 ();
 sg13g2_fill_1 FILLER_79_392 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_fill_1 FILLER_80_145 ();
 sg13g2_decap_4 FILLER_80_188 ();
 sg13g2_fill_2 FILLER_80_192 ();
 sg13g2_fill_2 FILLER_80_198 ();
 sg13g2_fill_2 FILLER_80_209 ();
 sg13g2_decap_8 FILLER_80_220 ();
 sg13g2_decap_8 FILLER_80_231 ();
 sg13g2_decap_4 FILLER_80_242 ();
 sg13g2_fill_2 FILLER_80_246 ();
 sg13g2_fill_1 FILLER_80_252 ();
 sg13g2_fill_1 FILLER_80_304 ();
 sg13g2_fill_2 FILLER_80_349 ();
 sg13g2_fill_1 FILLER_80_351 ();
 sg13g2_fill_2 FILLER_80_357 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_fill_1 FILLER_80_373 ();
 sg13g2_fill_2 FILLER_80_382 ();
 sg13g2_fill_1 FILLER_80_384 ();
 sg13g2_fill_2 FILLER_80_389 ();
 sg13g2_fill_1 FILLER_80_391 ();
 sg13g2_decap_4 FILLER_80_405 ();
 assign uio_oe[0] = net15;
 assign uio_oe[1] = net16;
 assign uio_oe[2] = net17;
 assign uio_oe[3] = net18;
 assign uio_oe[4] = net19;
 assign uio_oe[5] = net20;
 assign uio_oe[6] = net21;
 assign uio_oe[7] = net22;
 assign uio_out[0] = net23;
 assign uio_out[1] = net24;
 assign uio_out[2] = net25;
 assign uio_out[3] = net26;
 assign uio_out[4] = net27;
 assign uio_out[5] = net28;
 assign uio_out[6] = net29;
 assign uio_out[7] = net30;
endmodule

module tt_um_wokwi_group_11 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire \proj_10.net10 ;
 wire \proj_10.net11 ;
 wire \proj_10.net17 ;
 wire \proj_10.net18 ;
 wire \proj_10.net19 ;
 wire \proj_10.net20 ;
 wire \proj_10.net21 ;
 wire \proj_10.net8 ;
 wire \proj_10.net9 ;
 wire \proj_11.net15 ;
 wire \proj_11.net16 ;
 wire \proj_11.net17 ;
 wire \proj_11.net18 ;
 wire \proj_11.net19 ;
 wire \proj_11.net20 ;
 wire \proj_11.net21 ;
 wire \proj_11.net22 ;
 wire \proj_11.net23 ;
 wire \proj_11.net24 ;
 wire \proj_11.net9 ;
 wire \proj_12.net11 ;
 wire \proj_12.net12 ;
 wire \proj_12.net13 ;
 wire \proj_13.net6 ;
 wire \proj_13.net7 ;
 wire \proj_13.net8 ;
 wire \proj_14.net10 ;
 wire \proj_14.net11 ;
 wire \proj_14.net12 ;
 wire \proj_14.net13 ;
 wire \proj_14.net8 ;
 wire \proj_14.net9 ;
 wire \proj_15.net10 ;
 wire \proj_15.net11 ;
 wire \proj_15.net12 ;
 wire \proj_15.net13 ;
 wire \proj_15.net19 ;
 wire \proj_15.net20 ;
 wire \proj_15.net21 ;
 wire \proj_15.net22 ;
 wire \proj_15.net23 ;
 wire \proj_15.net24 ;
 wire \proj_15.net25 ;
 wire \proj_15.net26 ;
 wire \proj_15.net27 ;
 wire \proj_15.net28 ;
 wire \proj_15.net29 ;
 wire \proj_15.net30 ;
 wire \proj_15.net9 ;
 wire \proj__0.net11 ;
 wire \proj__0.net12 ;
 wire \proj__0.net13 ;
 wire \proj__0.net4 ;
 wire \proj__0.net5 ;
 wire \proj__1.net10 ;
 wire \proj__1.net11 ;
 wire \proj__1.net12 ;
 wire \proj__1.net13 ;
 wire \proj__1.net15 ;
 wire \proj__1.net16 ;
 wire \proj__1.net18 ;
 wire \proj__1.net19 ;
 wire \proj__1.net20 ;
 wire \proj__1.net21 ;
 wire \proj__1.net22 ;
 wire \proj__1.net23 ;
 wire \proj__1.net24 ;
 wire \proj__1.net25 ;
 wire \proj__1.net26 ;
 wire \proj__1.net27 ;
 wire \proj__1.net28 ;
 wire \proj__1.net29 ;
 wire \proj__1.net30 ;
 wire \proj__1.net31 ;
 wire \proj__1.net32 ;
 wire \proj__1.net33 ;
 wire \proj__1.net34 ;
 wire \proj__1.net35 ;
 wire \proj__1.net36 ;
 wire \proj__1.net37 ;
 wire \proj__1.net38 ;
 wire \proj__1.net9 ;
 wire \proj__2.net1 ;
 wire \proj__2.net16 ;
 wire \proj__2.net17 ;
 wire \proj__2.net18 ;
 wire \proj__2.net19 ;
 wire \proj__2.net2 ;
 wire \proj__2.net20 ;
 wire \proj__2.net21 ;
 wire \proj__2.net22 ;
 wire \proj__2.net23 ;
 wire \proj__2.net24 ;
 wire \proj__2.net25 ;
 wire \proj__2.net26 ;
 wire \proj__2.net27 ;
 wire \proj__2.net28 ;
 wire \proj__2.net29 ;
 wire \proj__2.net3 ;
 wire \proj__2.net30 ;
 wire \proj__2.net31 ;
 wire \proj__2.net32 ;
 wire \proj__2.net33 ;
 wire \proj__2.net34 ;
 wire \proj__2.net35 ;
 wire \proj__2.net36 ;
 wire \proj__2.net37 ;
 wire \proj__2.net38 ;
 wire \proj__2.net4 ;
 wire \proj__2.net5 ;
 wire \proj__3.net10 ;
 wire \proj__3.net11 ;
 wire \proj__3.net12 ;
 wire \proj__3.net9 ;
 wire \proj__4.net10 ;
 wire \proj__4.net11 ;
 wire \proj__4.net12 ;
 wire \proj__4.net13 ;
 wire \proj__5.net10 ;
 wire \proj__5.net11 ;
 wire \proj__5.net17 ;
 wire \proj__5.net18 ;
 wire \proj__5.net9 ;
 wire \proj__6.net10 ;
 wire \proj__6.net11 ;
 wire \proj__6.net17 ;
 wire \proj__6.net18 ;
 wire \proj__6.net19 ;
 wire \proj__6.net20 ;
 wire \proj__6.net21 ;
 wire \proj__6.net22 ;
 wire \proj__6.net23 ;
 wire \proj__6.net24 ;
 wire \proj__6.net25 ;
 wire \proj__6.net26 ;
 wire \proj__6.net27 ;
 wire \proj__6.net28 ;
 wire \proj__6.net29 ;
 wire \proj__6.net30 ;
 wire \proj__6.net31 ;
 wire \proj__6.net32 ;
 wire \proj__6.net33 ;
 wire \proj__6.net34 ;
 wire \proj__6.net35 ;
 wire \proj__6.net36 ;
 wire \proj__6.net37 ;
 wire \proj__6.net38 ;
 wire \proj__6.net39 ;
 wire \proj__6.net40 ;
 wire \proj__6.net41 ;
 wire \proj__6.net42 ;
 wire \proj__6.net43 ;
 wire \proj__6.net44 ;
 wire \proj__6.net45 ;
 wire \proj__6.net46 ;
 wire \proj__6.net47 ;
 wire \proj__6.net48 ;
 wire \proj__6.net5 ;
 wire \proj__6.net6 ;
 wire \proj__6.net7 ;
 wire \proj__6.net8 ;
 wire \proj__6.net9 ;
 wire \proj__7.net10 ;
 wire \proj__7.net11 ;
 wire \proj__7.net12 ;
 wire \proj__7.net9 ;
 wire \proj__8.net10 ;
 wire \proj__8.net11 ;
 wire \proj__8.net12 ;
 wire \proj__8.net13 ;
 wire \proj__8.net14 ;
 wire \proj__8.net15 ;
 wire \proj__8.net16 ;
 wire \proj__8.net22 ;
 wire \proj__8.net23 ;
 wire \proj__8.net24 ;
 wire \proj__8.net25 ;
 wire \proj__8.net26 ;
 wire \proj__8.net27 ;
 wire \proj__8.net28 ;
 wire \proj__8.net9 ;
 wire \proj__9.net15 ;
 wire \proj__9.net16 ;
 wire \proj__9.net17 ;
 wire \proj__9.net8 ;
 wire \proj__9.net9 ;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire \proj_13.flop1/notq ;
 wire net34;
 wire net35;
 wire clk_regs;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_1_0__leaf_clk_regs;
 wire clknet_1_1__leaf_clk_regs;

 sg13g2_inv_1 _090_ (.Y(_067_),
    .A(net74));
 sg13g2_and2_2 _091_ (.A(net5),
    .B(net4),
    .X(_068_));
 sg13g2_nand2b_1 _092_ (.Y(_069_),
    .B(_068_),
    .A_N(net7));
 sg13g2_nor2b_2 _093_ (.A(net6),
    .B_N(net7),
    .Y(_070_));
 sg13g2_nor2b_2 _094_ (.A(net5),
    .B_N(net4),
    .Y(_071_));
 sg13g2_and2_1 _095_ (.A(_070_),
    .B(_071_),
    .X(_072_));
 sg13g2_nor2_2 _096_ (.A(net5),
    .B(net4),
    .Y(_073_));
 sg13g2_a22oi_1 _097_ (.Y(_074_),
    .B1(_073_),
    .B2(net6),
    .A2(_071_),
    .A1(_070_));
 sg13g2_and2_1 _098_ (.A(net7),
    .B(net6),
    .X(_075_));
 sg13g2_and2_1 _099_ (.A(_073_),
    .B(_075_),
    .X(_076_));
 sg13g2_nor2b_2 _100_ (.A(net7),
    .B_N(net6),
    .Y(_077_));
 sg13g2_and2_2 _101_ (.A(_073_),
    .B(_077_),
    .X(_078_));
 sg13g2_a21oi_1 _102_ (.A1(_069_),
    .A2(_074_),
    .Y(_079_),
    .B1(_067_));
 sg13g2_and2_2 _103_ (.A(_070_),
    .B(_073_),
    .X(_080_));
 sg13g2_nand3_1 _104_ (.B(_068_),
    .C(_070_),
    .A(\proj_11.net9 ),
    .Y(_081_));
 sg13g2_nor2b_1 _105_ (.A(net4),
    .B_N(net5),
    .Y(_000_));
 sg13g2_and2_2 _106_ (.A(_077_),
    .B(_000_),
    .X(_001_));
 sg13g2_and2_1 _107_ (.A(_070_),
    .B(_000_),
    .X(_002_));
 sg13g2_and2_2 _108_ (.A(_071_),
    .B(_077_),
    .X(_003_));
 sg13g2_nand2_1 _109_ (.Y(_004_),
    .A(_071_),
    .B(_077_));
 sg13g2_and2_2 _110_ (.A(_075_),
    .B(_000_),
    .X(_005_));
 sg13g2_nand2_1 _111_ (.Y(_006_),
    .A(\proj_14.net12 ),
    .B(_005_));
 sg13g2_a22oi_1 _112_ (.Y(_007_),
    .B1(_003_),
    .B2(\proj__5.net11 ),
    .A2(_080_),
    .A1(\proj__8.net15 ));
 sg13g2_a221oi_1 _113_ (.B2(\proj_10.net11 ),
    .C1(_079_),
    .B1(_002_),
    .A1(\proj__6.net11 ),
    .Y(_008_),
    .A2(_001_));
 sg13g2_nand4_1 _114_ (.B(_006_),
    .C(_007_),
    .A(_081_),
    .Y(uo_out[6]),
    .D(_008_));
 sg13g2_nor2_2 _115_ (.A(net7),
    .B(net6),
    .Y(_009_));
 sg13g2_nand2_2 _116_ (.Y(_010_),
    .A(_073_),
    .B(_009_));
 sg13g2_nor2_1 _117_ (.A(\proj__0.net5 ),
    .B(_010_),
    .Y(_011_));
 sg13g2_nand3_1 _118_ (.B(_074_),
    .C(_004_),
    .A(_069_),
    .Y(_012_));
 sg13g2_nand2_1 _119_ (.Y(_013_),
    .A(net72),
    .B(_012_));
 sg13g2_a22oi_1 _120_ (.Y(_014_),
    .B1(_005_),
    .B2(\proj_14.net13 ),
    .A2(_080_),
    .A1(\proj__8.net16 ));
 sg13g2_and2_1 _121_ (.A(_010_),
    .B(_014_),
    .X(_015_));
 sg13g2_a21oi_2 _122_ (.B1(_011_),
    .Y(uo_out[7]),
    .A2(_015_),
    .A1(_013_));
 sg13g2_nor2_1 _123_ (.A(\proj__0.net4 ),
    .B(_010_),
    .Y(_016_));
 sg13g2_and2_1 _124_ (.A(_068_),
    .B(_077_),
    .X(_017_));
 sg13g2_and2_1 _125_ (.A(_081_),
    .B(_010_),
    .X(_018_));
 sg13g2_and2_2 _126_ (.A(_071_),
    .B(_009_),
    .X(_019_));
 sg13g2_a22oi_1 _127_ (.Y(_020_),
    .B1(_019_),
    .B2(\proj__1.net9 ),
    .A2(_076_),
    .A1(\proj_12.net11 ));
 sg13g2_and2_1 _128_ (.A(_071_),
    .B(_075_),
    .X(_021_));
 sg13g2_and2_2 _129_ (.A(_068_),
    .B(_075_),
    .X(_022_));
 sg13g2_and2_2 _130_ (.A(_000_),
    .B(_009_),
    .X(_023_));
 sg13g2_and2_1 _131_ (.A(_068_),
    .B(_009_),
    .X(_024_));
 sg13g2_a22oi_1 _132_ (.Y(_025_),
    .B1(_080_),
    .B2(\proj__8.net9 ),
    .A2(_078_),
    .A1(\proj__4.net10 ));
 sg13g2_a22oi_1 _133_ (.Y(_026_),
    .B1(_002_),
    .B2(\proj_10.net8 ),
    .A2(_001_),
    .A1(\proj__6.net5 ));
 sg13g2_and4_1 _134_ (.A(_018_),
    .B(_020_),
    .C(_025_),
    .D(_026_),
    .X(_027_));
 sg13g2_a22oi_1 _135_ (.Y(_028_),
    .B1(_021_),
    .B2(\proj_13.net6 ),
    .A2(_003_),
    .A1(\proj__5.net9 ));
 sg13g2_a22oi_1 _136_ (.Y(_029_),
    .B1(_023_),
    .B2(\proj__2.net1 ),
    .A2(_072_),
    .A1(\proj__9.net8 ));
 sg13g2_a22oi_1 _137_ (.Y(_030_),
    .B1(_022_),
    .B2(\proj_15.net9 ),
    .A2(_017_),
    .A1(\proj__7.net9 ));
 sg13g2_a22oi_1 _138_ (.Y(_031_),
    .B1(_024_),
    .B2(\proj__3.net9 ),
    .A2(_005_),
    .A1(\proj_14.net8 ));
 sg13g2_and4_1 _139_ (.A(_028_),
    .B(_029_),
    .C(_030_),
    .D(_031_),
    .X(_032_));
 sg13g2_a21oi_1 _140_ (.A1(_027_),
    .A2(_032_),
    .Y(uo_out[0]),
    .B1(_016_));
 sg13g2_nand3_1 _141_ (.B(_068_),
    .C(_009_),
    .A(\proj__3.net10 ),
    .Y(_033_));
 sg13g2_nand2_1 _142_ (.Y(_034_),
    .A(\proj_15.net10 ),
    .B(_022_));
 sg13g2_a22oi_1 _143_ (.Y(_035_),
    .B1(_078_),
    .B2(\proj__4.net11 ),
    .A2(_072_),
    .A1(\proj__9.net9 ));
 sg13g2_a22oi_1 _144_ (.Y(_036_),
    .B1(_003_),
    .B2(net89),
    .A2(_001_),
    .A1(\proj__6.net6 ));
 sg13g2_a22oi_1 _145_ (.Y(_037_),
    .B1(_021_),
    .B2(\proj_13.net7 ),
    .A2(_076_),
    .A1(\proj_12.net12 ));
 sg13g2_a22oi_1 _146_ (.Y(_038_),
    .B1(_005_),
    .B2(\proj_14.net9 ),
    .A2(_080_),
    .A1(\proj__8.net10 ));
 sg13g2_nand4_1 _147_ (.B(_036_),
    .C(_037_),
    .A(_035_),
    .Y(_039_),
    .D(_038_));
 sg13g2_a22oi_1 _148_ (.Y(_040_),
    .B1(_019_),
    .B2(\proj__1.net10 ),
    .A2(_002_),
    .A1(\proj_10.net9 ));
 sg13g2_a22oi_1 _149_ (.Y(_041_),
    .B1(_023_),
    .B2(\proj__2.net2 ),
    .A2(_017_),
    .A1(\proj__7.net10 ));
 sg13g2_nand4_1 _150_ (.B(_034_),
    .C(_040_),
    .A(_033_),
    .Y(_042_),
    .D(_041_));
 sg13g2_or2_2 _151_ (.X(uo_out[1]),
    .B(_042_),
    .A(_039_));
 sg13g2_a22oi_1 _152_ (.Y(_043_),
    .B1(_005_),
    .B2(\proj_14.net9 ),
    .A2(_002_),
    .A1(\proj_10.net10 ));
 sg13g2_a22oi_1 _153_ (.Y(_044_),
    .B1(_078_),
    .B2(\proj__4.net12 ),
    .A2(_076_),
    .A1(\proj_12.net13 ));
 sg13g2_a22oi_1 _154_ (.Y(_045_),
    .B1(_023_),
    .B2(\proj__2.net3 ),
    .A2(_017_),
    .A1(\proj__7.net11 ));
 sg13g2_nand3_1 _155_ (.B(_044_),
    .C(_045_),
    .A(_043_),
    .Y(_046_));
 sg13g2_nand3_1 _156_ (.B(_068_),
    .C(_009_),
    .A(\proj__3.net11 ),
    .Y(_047_));
 sg13g2_a22oi_1 _157_ (.Y(_048_),
    .B1(_022_),
    .B2(\proj_15.net11 ),
    .A2(_001_),
    .A1(\proj__6.net7 ));
 sg13g2_a22oi_1 _158_ (.Y(_049_),
    .B1(_019_),
    .B2(\proj__1.net11 ),
    .A2(_080_),
    .A1(\proj__8.net11 ));
 sg13g2_a22oi_1 _159_ (.Y(_050_),
    .B1(_021_),
    .B2(\proj_13.net8 ),
    .A2(_003_),
    .A1(net86));
 sg13g2_nand4_1 _160_ (.B(_048_),
    .C(_049_),
    .A(_047_),
    .Y(_051_),
    .D(_050_));
 sg13g2_or2_1 _161_ (.X(uo_out[2]),
    .B(_051_),
    .A(_046_));
 sg13g2_nand3_1 _162_ (.B(_068_),
    .C(_009_),
    .A(\proj__3.net12 ),
    .Y(_052_));
 sg13g2_nand2_1 _163_ (.Y(_053_),
    .A(\proj__8.net12 ),
    .B(_080_));
 sg13g2_a22oi_1 _164_ (.Y(_054_),
    .B1(_023_),
    .B2(\proj__2.net4 ),
    .A2(_005_),
    .A1(\proj_14.net10 ));
 sg13g2_a22oi_1 _165_ (.Y(_055_),
    .B1(_022_),
    .B2(\proj_15.net12 ),
    .A2(_017_),
    .A1(\proj__7.net12 ));
 sg13g2_a22oi_1 _166_ (.Y(_056_),
    .B1(_019_),
    .B2(\proj__1.net12 ),
    .A2(_078_),
    .A1(\proj__4.net13 ));
 sg13g2_and4_1 _167_ (.A(_081_),
    .B(_053_),
    .C(_055_),
    .D(_056_),
    .X(_057_));
 sg13g2_a22oi_1 _168_ (.Y(_058_),
    .B1(_003_),
    .B2(\proj__5.net10 ),
    .A2(_001_),
    .A1(\proj__6.net8 ));
 sg13g2_nand4_1 _169_ (.B(_054_),
    .C(_057_),
    .A(_052_),
    .Y(uo_out[3]),
    .D(_058_));
 sg13g2_nand2_1 _170_ (.Y(_059_),
    .A(net79),
    .B(_012_));
 sg13g2_and2_1 _171_ (.A(\proj_15.net13 ),
    .B(_022_),
    .X(_060_));
 sg13g2_nand2_1 _172_ (.Y(_061_),
    .A(\proj_14.net11 ),
    .B(_005_));
 sg13g2_and2_1 _173_ (.A(_081_),
    .B(_061_),
    .X(_062_));
 sg13g2_a22oi_1 _174_ (.Y(_063_),
    .B1(_019_),
    .B2(\proj__1.net13 ),
    .A2(_080_),
    .A1(\proj__8.net13 ));
 sg13g2_a221oi_1 _175_ (.B2(\proj__2.net5 ),
    .C1(_060_),
    .B1(_023_),
    .A1(\proj__6.net9 ),
    .Y(_064_),
    .A2(_001_));
 sg13g2_nand4_1 _176_ (.B(_062_),
    .C(_063_),
    .A(_059_),
    .Y(uo_out[4]),
    .D(_064_));
 sg13g2_nand2_1 _177_ (.Y(_065_),
    .A(net77),
    .B(_012_));
 sg13g2_a22oi_1 _178_ (.Y(_066_),
    .B1(_001_),
    .B2(\proj__6.net10 ),
    .A2(_080_),
    .A1(\proj__8.net14 ));
 sg13g2_nand3_1 _179_ (.B(_065_),
    .C(_066_),
    .A(_062_),
    .Y(uo_out[5]));
 sg13g2_tielo \proj__1.and1/_0__9  (.L_LO(net9));
 sg13g2_tielo \proj__1.and3/_0__10  (.L_LO(net10));
 sg13g2_tielo \proj__1.and3/_0__11  (.L_LO(net11));
 sg13g2_tielo \proj__1.xor2/_0__12  (.L_LO(net12));
 sg13g2_tielo \proj__2.and1/_0__13  (.L_LO(net13));
 sg13g2_tielo \proj__2.and3/_0__14  (.L_LO(net14));
 sg13g2_tielo \proj__2.xor1/_0__15  (.L_LO(net15));
 sg13g2_tielo tt_um_wokwi_group_11_16 (.L_LO(net16));
 sg13g2_tielo tt_um_wokwi_group_11_17 (.L_LO(net17));
 sg13g2_tielo tt_um_wokwi_group_11_18 (.L_LO(net18));
 sg13g2_tielo tt_um_wokwi_group_11_19 (.L_LO(net19));
 sg13g2_tielo tt_um_wokwi_group_11_20 (.L_LO(net20));
 sg13g2_tielo tt_um_wokwi_group_11_21 (.L_LO(net21));
 sg13g2_tielo tt_um_wokwi_group_11_22 (.L_LO(net22));
 sg13g2_tielo tt_um_wokwi_group_11_23 (.L_LO(net23));
 sg13g2_tielo tt_um_wokwi_group_11_24 (.L_LO(net24));
 sg13g2_tielo tt_um_wokwi_group_11_25 (.L_LO(net25));
 sg13g2_tielo tt_um_wokwi_group_11_26 (.L_LO(net26));
 sg13g2_tielo tt_um_wokwi_group_11_27 (.L_LO(net27));
 sg13g2_tielo tt_um_wokwi_group_11_28 (.L_LO(net28));
 sg13g2_tielo tt_um_wokwi_group_11_29 (.L_LO(net29));
 sg13g2_tielo tt_um_wokwi_group_11_30 (.L_LO(net30));
 sg13g2_tielo tt_um_wokwi_group_11_31 (.L_LO(net31));
 sg13g2_tiehi \proj_13.flop1/_1__32  (.L_HI(net32));
 sg13g2_and2_1 \proj_10.and1/_0_  (.A(\proj_10.net17 ),
    .B(\proj_10.net11 ),
    .X(\proj_10.net18 ));
 sg13g2_and2_1 \proj_10.and2/_0_  (.A(net75),
    .B(\proj_10.net11 ),
    .X(\proj_10.net19 ));
 sg13g2_and2_1 \proj_10.and3/_0_  (.A(net74),
    .B(net73),
    .X(\proj_10.net21 ));
 sg13g2_and2_1 \proj_10.and4/_0_  (.A(net84),
    .B(net87),
    .X(\proj_10.net9 ));
 sg13g2_inv_1 \proj_10.not1/_0_  (.Y(\proj_10.net8 ),
    .A(net91));
 sg13g2_inv_1 \proj_10.not5/_0_  (.Y(\proj_10.net17 ),
    .A(net73));
 sg13g2_or2_1 \proj_10.or1/_0_  (.X(\proj_10.net20 ),
    .B(\proj_10.net18 ),
    .A(\proj_10.net19 ));
 sg13g2_or2_1 \proj_10.or2/_0_  (.X(\proj_10.net11 ),
    .B(\proj_10.net20 ),
    .A(\proj_10.net21 ));
 sg13g2_or2_1 \proj_10.or3/_0_  (.X(\proj_10.net10 ),
    .B(net80),
    .A(net78));
 sg13g2_and2_1 \proj_11.and1/_0_  (.A(\proj_11.net15 ),
    .B(net91),
    .X(\proj_11.net16 ));
 sg13g2_and2_1 \proj_11.and2/_0_  (.A(\proj_11.net17 ),
    .B(net83),
    .X(\proj_11.net18 ));
 sg13g2_and2_1 \proj_11.and3/_0_  (.A(\proj_11.net19 ),
    .B(net78),
    .X(\proj_11.net20 ));
 sg13g2_and2_1 \proj_11.and4/_0_  (.A(\proj_11.net21 ),
    .B(net74),
    .X(\proj_11.net22 ));
 sg13g2_and2_1 \proj_11.and5/_0_  (.A(\proj_11.net22 ),
    .B(\proj_11.net16 ),
    .X(\proj_11.net23 ));
 sg13g2_and2_1 \proj_11.and6/_0_  (.A(\proj_11.net20 ),
    .B(\proj_11.net18 ),
    .X(\proj_11.net24 ));
 sg13g2_and2_1 \proj_11.and7/_0_  (.A(\proj_11.net24 ),
    .B(\proj_11.net23 ),
    .X(\proj_11.net9 ));
 sg13g2_inv_1 \proj_11.not1/_0_  (.Y(\proj_11.net15 ),
    .A(net87));
 sg13g2_inv_1 \proj_11.not2/_0_  (.Y(\proj_11.net17 ),
    .A(net80));
 sg13g2_inv_1 \proj_11.not3/_0_  (.Y(\proj_11.net19 ),
    .A(net76));
 sg13g2_inv_1 \proj_11.not4/_0_  (.Y(\proj_11.net21 ),
    .A(net72));
 sg13g2_and2_1 \proj_12.and1/_0_  (.A(net1),
    .B(clknet_1_0__leaf_clk),
    .X(\proj_12.net11 ));
 sg13g2_nand2_1 \proj_12.nand1/_0_  (.Y(\proj_12.net13 ),
    .A(net82),
    .B(net86));
 sg13g2_xor2_1 \proj_12.xor1/_0_  (.B(net93),
    .A(net89),
    .X(\proj_12.net12 ));
 sg13g2_and2_1 \proj_13.and1/_0_  (.A(net86),
    .B(net89),
    .X(\proj_13.net7 ));
 sg13g2_dfrbp_1 \proj_13.flop1/_1_  (.CLK(clknet_1_0__leaf_clk_regs),
    .RESET_B(net32),
    .D(net82),
    .Q_N(\proj_13.flop1/notq ),
    .Q(\proj_13.net8 ));
 sg13g2_tiehi \proj__6.flop1/_1__33  (.L_HI(net33));
 sg13g2_inv_1 \proj_13.not1/_0_  (.Y(\proj_13.net6 ),
    .A(net93));
 sg13g2_and2_1 \proj_14.and1/_0_  (.A(net87),
    .B(net91),
    .X(\proj_14.net10 ));
 sg13g2_nand2_1 \proj_14.nand1/_0_  (.Y(\proj_14.net11 ),
    .A(net76),
    .B(net78));
 sg13g2_inv_1 \proj_14.not1/_0_  (.Y(\proj_14.net8 ),
    .A(\proj_14.net10 ));
 sg13g2_inv_1 \proj_14.not2/_0_  (.Y(\proj_14.net13 ),
    .A(net72));
 sg13g2_inv_1 \proj_14.not3/_0_  (.Y(\proj_14.net12 ),
    .A(net84));
 sg13g2_or2_1 \proj_14.or1/_0_  (.X(\proj_14.net9 ),
    .B(\proj_14.net12 ),
    .A(net82));
 sg13g2_and2_1 \proj_15.and1/_0_  (.A(net89),
    .B(net92),
    .X(\proj_15.net19 ));
 sg13g2_and2_1 \proj_15.and2/_0_  (.A(net81),
    .B(net85),
    .X(\proj_15.net21 ));
 sg13g2_and2_1 \proj_15.and3/_0_  (.A(\proj_15.net19 ),
    .B(\proj_15.net20 ),
    .X(\proj_15.net22 ));
 sg13g2_and2_1 \proj_15.and4/_0_  (.A(net77),
    .B(net79),
    .X(\proj_15.net25 ));
 sg13g2_and2_1 \proj_15.and5/_0_  (.A(\proj_15.net24 ),
    .B(\proj_15.net23 ),
    .X(\proj_15.net26 ));
 sg13g2_and2_1 \proj_15.and6/_0_  (.A(net73),
    .B(net75),
    .X(\proj_15.net29 ));
 sg13g2_and2_1 \proj_15.and7/_0_  (.A(\proj_15.net28 ),
    .B(\proj_15.net27 ),
    .X(\proj_15.net30 ));
 sg13g2_or2_1 \proj_15.or1/_0_  (.X(\proj_15.net23 ),
    .B(\proj_15.net21 ),
    .A(\proj_15.net22 ));
 sg13g2_or2_1 \proj_15.or2/_0_  (.X(\proj_15.net27 ),
    .B(\proj_15.net26 ),
    .A(\proj_15.net25 ));
 sg13g2_or2_1 \proj_15.or3/_0_  (.X(\proj_15.net13 ),
    .B(\proj_15.net30 ),
    .A(\proj_15.net29 ));
 sg13g2_xor2_1 \proj_15.xor1/_0_  (.B(net92),
    .A(net88),
    .X(\proj_15.net9 ));
 sg13g2_xor2_1 \proj_15.xor2/_0_  (.B(net85),
    .A(net81),
    .X(\proj_15.net20 ));
 sg13g2_xor2_1 \proj_15.xor3/_0_  (.B(\proj_15.net20 ),
    .A(\proj_15.net19 ),
    .X(\proj_15.net10 ));
 sg13g2_xor2_1 \proj_15.xor4/_0_  (.B(net79),
    .A(net77),
    .X(\proj_15.net24 ));
 sg13g2_xor2_1 \proj_15.xor5/_0_  (.B(\proj_15.net24 ),
    .A(\proj_15.net23 ),
    .X(\proj_15.net11 ));
 sg13g2_xor2_1 \proj_15.xor6/_0_  (.B(net75),
    .A(net73),
    .X(\proj_15.net28 ));
 sg13g2_xor2_1 \proj_15.xor7/_0_  (.B(\proj_15.net27 ),
    .A(\proj_15.net28 ),
    .X(\proj_15.net12 ));
 sg13g2_and2_1 \proj__0.and1/_0_  (.A(net84),
    .B(\proj__0.net11 ),
    .X(\proj__0.net12 ));
 sg13g2_and2_1 \proj__0.and2/_0_  (.A(net90),
    .B(net94),
    .X(\proj__0.net13 ));
 sg13g2_or2_1 \proj__0.or1/_0_  (.X(\proj__0.net5 ),
    .B(\proj__0.net12 ),
    .A(\proj__0.net13 ));
 sg13g2_xor2_1 \proj__0.xor1/_0_  (.B(net94),
    .A(net90),
    .X(\proj__0.net11 ));
 sg13g2_xor2_1 \proj__0.xor2/_0_  (.B(\proj__0.net11 ),
    .A(net84),
    .X(\proj__0.net4 ));
 sg13g2_and2_1 \proj__1.and1/_0_  (.A(net9),
    .B(net8),
    .X(\proj__1.net18 ));
 sg13g2_and2_1 \proj__1.and10/_0_  (.A(net72),
    .B(net82),
    .X(\proj__1.net35 ));
 sg13g2_and2_1 \proj__1.and11/_0_  (.A(\proj__1.net33 ),
    .B(net80),
    .X(\proj__1.net36 ));
 sg13g2_and2_1 \proj__1.and12/_0_  (.A(\proj__1.net33 ),
    .B(net72),
    .X(\proj__1.net37 ));
 sg13g2_and2_1 \proj__1.and2/_0_  (.A(net78),
    .B(net91),
    .X(\proj__1.net16 ));
 sg13g2_and2_1 \proj__1.and3/_0_  (.A(net11),
    .B(net10),
    .X(\proj__1.net19 ));
 sg13g2_and2_1 \proj__1.and4/_0_  (.A(net76),
    .B(net87),
    .X(\proj__1.net23 ));
 sg13g2_and2_1 \proj__1.and5/_0_  (.A(\proj__1.net21 ),
    .B(net87),
    .X(\proj__1.net24 ));
 sg13g2_and2_1 \proj__1.and6/_0_  (.A(\proj__1.net21 ),
    .B(net76),
    .X(\proj__1.net25 ));
 sg13g2_and2_1 \proj__1.and7/_0_  (.A(net74),
    .B(net80),
    .X(\proj__1.net29 ));
 sg13g2_and2_1 \proj__1.and8/_0_  (.A(\proj__1.net27 ),
    .B(net83),
    .X(\proj__1.net30 ));
 sg13g2_and2_1 \proj__1.and9/_0_  (.A(\proj__1.net27 ),
    .B(net74),
    .X(\proj__1.net31 ));
 sg13g2_or2_1 \proj__1.or1/_0_  (.X(\proj__1.net20 ),
    .B(\proj__1.net16 ),
    .A(\proj__1.net18 ));
 sg13g2_or2_1 \proj__1.or2/_0_  (.X(\proj__1.net21 ),
    .B(\proj__1.net20 ),
    .A(\proj__1.net19 ));
 sg13g2_or2_1 \proj__1.or3/_0_  (.X(\proj__1.net26 ),
    .B(\proj__1.net23 ),
    .A(\proj__1.net24 ));
 sg13g2_or2_1 \proj__1.or4/_0_  (.X(\proj__1.net27 ),
    .B(\proj__1.net26 ),
    .A(\proj__1.net25 ));
 sg13g2_or2_1 \proj__1.or5/_0_  (.X(\proj__1.net32 ),
    .B(\proj__1.net29 ),
    .A(\proj__1.net30 ));
 sg13g2_or2_1 \proj__1.or6/_0_  (.X(\proj__1.net33 ),
    .B(\proj__1.net32 ),
    .A(\proj__1.net31 ));
 sg13g2_or2_1 \proj__1.or7/_0_  (.X(\proj__1.net38 ),
    .B(\proj__1.net35 ),
    .A(\proj__1.net36 ));
 sg13g2_or2_1 \proj__1.or8/_0_  (.X(\proj__1.net13 ),
    .B(\proj__1.net38 ),
    .A(\proj__1.net37 ));
 sg13g2_xor2_1 \proj__1.xor1/_0_  (.B(net93),
    .A(net79),
    .X(\proj__1.net15 ));
 sg13g2_xor2_1 \proj__1.xor2/_0_  (.B(net12),
    .A(\proj__1.net15 ),
    .X(\proj__1.net9 ));
 sg13g2_xor2_1 \proj__1.xor3/_0_  (.B(net87),
    .A(net76),
    .X(\proj__1.net22 ));
 sg13g2_xor2_1 \proj__1.xor4/_0_  (.B(\proj__1.net21 ),
    .A(\proj__1.net22 ),
    .X(\proj__1.net10 ));
 sg13g2_xor2_1 \proj__1.xor5/_0_  (.B(net83),
    .A(net74),
    .X(\proj__1.net28 ));
 sg13g2_xor2_1 \proj__1.xor6/_0_  (.B(\proj__1.net27 ),
    .A(\proj__1.net28 ),
    .X(\proj__1.net11 ));
 sg13g2_xor2_1 \proj__1.xor7/_0_  (.B(net80),
    .A(net72),
    .X(\proj__1.net34 ));
 sg13g2_xor2_1 \proj__1.xor8/_0_  (.B(\proj__1.net33 ),
    .A(\proj__1.net34 ),
    .X(\proj__1.net12 ));
 sg13g2_and2_1 \proj__2.and1/_0_  (.A(net88),
    .B(net13),
    .X(\proj__2.net16 ));
 sg13g2_and2_1 \proj__2.and10/_0_  (.A(net73),
    .B(\proj__2.net32 ),
    .X(\proj__2.net34 ));
 sg13g2_and2_1 \proj__2.and11/_0_  (.A(net75),
    .B(net73),
    .X(\proj__2.net35 ));
 sg13g2_and2_1 \proj__2.and12/_0_  (.A(net2),
    .B(\proj__2.net32 ),
    .X(\proj__2.net36 ));
 sg13g2_and2_1 \proj__2.and2/_0_  (.A(net92),
    .B(net88),
    .X(\proj__2.net17 ));
 sg13g2_and2_1 \proj__2.and3/_0_  (.A(net92),
    .B(net14),
    .X(\proj__2.net18 ));
 sg13g2_and2_1 \proj__2.and4/_0_  (.A(net81),
    .B(\proj__2.net20 ),
    .X(\proj__2.net22 ));
 sg13g2_and2_1 \proj__2.and5/_0_  (.A(net85),
    .B(net81),
    .X(\proj__2.net23 ));
 sg13g2_and2_1 \proj__2.and6/_0_  (.A(net85),
    .B(\proj__2.net20 ),
    .X(\proj__2.net24 ));
 sg13g2_and2_1 \proj__2.and7/_0_  (.A(net77),
    .B(\proj__2.net26 ),
    .X(\proj__2.net28 ));
 sg13g2_and2_1 \proj__2.and8/_0_  (.A(net79),
    .B(net76),
    .X(\proj__2.net29 ));
 sg13g2_and2_1 \proj__2.and9/_0_  (.A(net79),
    .B(\proj__2.net26 ),
    .X(\proj__2.net30 ));
 sg13g2_or2_1 \proj__2.or1/_0_  (.X(\proj__2.net19 ),
    .B(\proj__2.net18 ),
    .A(\proj__2.net16 ));
 sg13g2_or2_1 \proj__2.or2/_0_  (.X(\proj__2.net20 ),
    .B(\proj__2.net19 ),
    .A(\proj__2.net17 ));
 sg13g2_or2_1 \proj__2.or3/_0_  (.X(\proj__2.net25 ),
    .B(\proj__2.net24 ),
    .A(\proj__2.net22 ));
 sg13g2_or2_1 \proj__2.or4/_0_  (.X(\proj__2.net26 ),
    .B(\proj__2.net25 ),
    .A(\proj__2.net23 ));
 sg13g2_or2_1 \proj__2.or5/_0_  (.X(\proj__2.net31 ),
    .B(\proj__2.net30 ),
    .A(\proj__2.net28 ));
 sg13g2_or2_1 \proj__2.or6/_0_  (.X(\proj__2.net32 ),
    .B(\proj__2.net31 ),
    .A(\proj__2.net29 ));
 sg13g2_or2_1 \proj__2.or7/_0_  (.X(\proj__2.net37 ),
    .B(\proj__2.net36 ),
    .A(\proj__2.net34 ));
 sg13g2_or2_1 \proj__2.or8/_0_  (.X(\proj__2.net5 ),
    .B(\proj__2.net37 ),
    .A(\proj__2.net35 ));
 sg13g2_xor2_1 \proj__2.xor1/_0_  (.B(net15),
    .A(net92),
    .X(\proj__2.net21 ));
 sg13g2_xor2_1 \proj__2.xor2/_0_  (.B(\proj__2.net21 ),
    .A(net88),
    .X(\proj__2.net1 ));
 sg13g2_xor2_1 \proj__2.xor3/_0_  (.B(\proj__2.net20 ),
    .A(net85),
    .X(\proj__2.net27 ));
 sg13g2_xor2_1 \proj__2.xor4/_0_  (.B(\proj__2.net27 ),
    .A(net81),
    .X(\proj__2.net2 ));
 sg13g2_xor2_1 \proj__2.xor5/_0_  (.B(\proj__2.net26 ),
    .A(net79),
    .X(\proj__2.net33 ));
 sg13g2_xor2_1 \proj__2.xor6/_0_  (.B(\proj__2.net33 ),
    .A(net77),
    .X(\proj__2.net3 ));
 sg13g2_xor2_1 \proj__2.xor7/_0_  (.B(\proj__2.net32 ),
    .A(net75),
    .X(\proj__2.net38 ));
 sg13g2_xor2_1 \proj__2.xor8/_0_  (.B(\proj__2.net38 ),
    .A(net3),
    .X(\proj__2.net4 ));
 sg13g2_inv_1 \proj__3.not1/_0_  (.Y(\proj__3.net9 ),
    .A(net91));
 sg13g2_inv_1 \proj__3.not2/_0_  (.Y(\proj__3.net10 ),
    .A(net88));
 sg13g2_inv_1 \proj__3.not3/_0_  (.Y(\proj__3.net11 ),
    .A(net86));
 sg13g2_inv_1 \proj__3.not4/_0_  (.Y(\proj__3.net12 ),
    .A(net80));
 sg13g2_and2_1 \proj__4.and1/_0_  (.A(net83),
    .B(net90),
    .X(\proj__4.net13 ));
 sg13g2_inv_1 \proj__4.not2/_0_  (.Y(\proj__4.net12 ),
    .A(net81));
 sg13g2_inv_1 \proj__4.not5/_0_  (.Y(\proj__4.net10 ),
    .A(net91));
 sg13g2_inv_1 \proj__4.not6/_0_  (.Y(\proj__4.net11 ),
    .A(net93));
 sg13g2_and2_1 \proj__5.and1/_0_  (.A(\proj__5.net17 ),
    .B(net74),
    .X(\proj__5.net11 ));
 sg13g2_inv_1 \proj__5.not1/_0_  (.Y(\proj__5.net17 ),
    .A(net72));
 sg13g2_inv_1 \proj__5.not2/_0_  (.Y(\proj__5.net10 ),
    .A(net81));
 sg13g2_inv_1 \proj__5.not3/_0_  (.Y(\proj__5.net18 ),
    .A(net93));
 sg13g2_or2_1 \proj__5.or1/_0_  (.X(\proj__5.net9 ),
    .B(\proj__5.net18 ),
    .A(net73));
 sg13g2_and2_1 \proj__6.and1/_0_  (.A(\proj__6.net19 ),
    .B(\proj__6.net17 ),
    .X(\proj__6.net28 ));
 sg13g2_and2_1 \proj__6.and10/_0_  (.A(\proj__6.net22 ),
    .B(\proj__6.net42 ),
    .X(\proj__6.net41 ));
 sg13g2_and2_1 \proj__6.and11/_0_  (.A(\proj__6.net20 ),
    .B(\proj__6.net18 ),
    .X(\proj__6.net42 ));
 sg13g2_and2_1 \proj__6.and12/_0_  (.A(\proj__6.net22 ),
    .B(\proj__6.net18 ),
    .X(\proj__6.net44 ));
 sg13g2_and2_1 \proj__6.and13/_0_  (.A(\proj__6.net19 ),
    .B(\proj__6.net22 ),
    .X(\proj__6.net46 ));
 sg13g2_and2_1 \proj__6.and14/_0_  (.A(\proj__6.net17 ),
    .B(\proj__6.net46 ),
    .X(\proj__6.net45 ));
 sg13g2_and2_1 \proj__6.and15/_0_  (.A(\proj__6.net19 ),
    .B(\proj__6.net18 ),
    .X(\proj__6.net47 ));
 sg13g2_and2_1 \proj__6.and16/_0_  (.A(\proj__6.net22 ),
    .B(\proj__6.net47 ),
    .X(\proj__6.net48 ));
 sg13g2_and2_1 \proj__6.and2/_0_  (.A(\proj__6.net22 ),
    .B(\proj__6.net28 ),
    .X(\proj__6.net29 ));
 sg13g2_and2_1 \proj__6.and3/_0_  (.A(\proj__6.net21 ),
    .B(\proj__6.net31 ),
    .X(\proj__6.net32 ));
 sg13g2_and2_1 \proj__6.and4/_0_  (.A(\proj__6.net20 ),
    .B(\proj__6.net18 ),
    .X(\proj__6.net33 ));
 sg13g2_and2_1 \proj__6.and5/_0_  (.A(\proj__6.net21 ),
    .B(\proj__6.net34 ),
    .X(\proj__6.net35 ));
 sg13g2_and2_1 \proj__6.and6/_0_  (.A(\proj__6.net19 ),
    .B(\proj__6.net22 ),
    .X(\proj__6.net37 ));
 sg13g2_and2_1 \proj__6.and7/_0_  (.A(\proj__6.net20 ),
    .B(\proj__6.net21 ),
    .X(\proj__6.net39 ));
 sg13g2_and2_1 \proj__6.and8/_0_  (.A(\proj__6.net18 ),
    .B(\proj__6.net39 ),
    .X(\proj__6.net38 ));
 sg13g2_and2_1 \proj__6.and9/_0_  (.A(\proj__6.net19 ),
    .B(\proj__6.net18 ),
    .X(\proj__6.net40 ));
 sg13g2_dfrbp_1 \proj__6.flop1/_1_  (.CLK(clknet_1_1__leaf_clk_regs),
    .RESET_B(net33),
    .D(net93),
    .Q_N(\proj__6.net18 ),
    .Q(\proj__6.net17 ));
 sg13g2_tiehi \proj__6.flop2/_1__34  (.L_HI(net34));
 sg13g2_dfrbp_1 \proj__6.flop2/_1_  (.CLK(clknet_1_0__leaf_clk_regs),
    .RESET_B(net34),
    .D(net89),
    .Q_N(\proj__6.net20 ),
    .Q(\proj__6.net19 ));
 sg13g2_tiehi \proj__6.flop3/_1__35  (.L_HI(net35));
 sg13g2_dfrbp_1 \proj__6.flop3/_1_  (.CLK(clknet_1_1__leaf_clk_regs),
    .RESET_B(net35),
    .D(net86),
    .Q_N(\proj__6.net22 ),
    .Q(\proj__6.net21 ));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_inv_1 \proj__6.not1/_0_  (.Y(\proj__6.net26 ),
    .A(\proj__6.net25 ));
 sg13g2_inv_1 \proj__6.not2/_0_  (.Y(\proj__6.net27 ),
    .A(\proj__6.net24 ));
 sg13g2_inv_1 \proj__6.not3/_0_  (.Y(\proj__6.net6 ),
    .A(\proj__6.net32 ));
 sg13g2_inv_1 \proj__6.not4/_0_  (.Y(\proj__6.net7 ),
    .A(\proj__6.net48 ));
 sg13g2_or2_1 \proj__6.or1/_0_  (.X(\proj__6.net25 ),
    .B(\proj__6.net23 ),
    .A(\proj__6.net24 ));
 sg13g2_or2_1 \proj__6.or2/_0_  (.X(\proj__6.net30 ),
    .B(\proj__6.net26 ),
    .A(\proj__6.net27 ));
 sg13g2_or2_1 \proj__6.or3/_0_  (.X(\proj__6.net5 ),
    .B(\proj__6.net30 ),
    .A(\proj__6.net29 ));
 sg13g2_or2_1 \proj__6.or4/_0_  (.X(\proj__6.net10 ),
    .B(\proj__6.net33 ),
    .A(\proj__6.net35 ));
 sg13g2_or2_1 \proj__6.or5/_0_  (.X(\proj__6.net11 ),
    .B(\proj__6.net35 ),
    .A(\proj__6.net36 ));
 sg13g2_or2_1 \proj__6.or6/_0_  (.X(\proj__6.net36 ),
    .B(\proj__6.net37 ),
    .A(\proj__6.net38 ));
 sg13g2_or2_1 \proj__6.or7/_0_  (.X(\proj__6.net9 ),
    .B(\proj__6.net40 ),
    .A(\proj__6.net41 ));
 sg13g2_or2_1 \proj__6.or8/_0_  (.X(\proj__6.net8 ),
    .B(\proj__6.net35 ),
    .A(\proj__6.net43 ));
 sg13g2_or2_1 \proj__6.or9/_0_  (.X(\proj__6.net43 ),
    .B(\proj__6.net44 ),
    .A(\proj__6.net45 ));
 sg13g2_xor2_1 \proj__6.xor1/_0_  (.B(\proj__6.net17 ),
    .A(\proj__6.net19 ),
    .X(\proj__6.net23 ));
 sg13g2_xor2_1 \proj__6.xor2/_0_  (.B(\proj__6.net17 ),
    .A(\proj__6.net21 ),
    .X(\proj__6.net24 ));
 sg13g2_xor2_1 \proj__6.xor3/_0_  (.B(\proj__6.net17 ),
    .A(\proj__6.net19 ),
    .X(\proj__6.net31 ));
 sg13g2_xor2_1 \proj__6.xor4/_0_  (.B(\proj__6.net17 ),
    .A(\proj__6.net19 ),
    .X(\proj__6.net34 ));
 sg13g2_inv_1 \proj__7.not1/_0_  (.Y(\proj__7.net9 ),
    .A(net92));
 sg13g2_inv_1 \proj__7.not2/_0_  (.Y(\proj__7.net10 ),
    .A(net88));
 sg13g2_inv_1 \proj__7.not3/_0_  (.Y(\proj__7.net11 ),
    .A(net85));
 sg13g2_inv_1 \proj__7.not4/_0_  (.Y(\proj__7.net12 ),
    .A(net81));
 sg13g2_and2_1 \proj__8.and1/_0_  (.A(net83),
    .B(\proj__8.net23 ),
    .X(\proj__8.net11 ));
 sg13g2_and2_1 \proj__8.and2/_0_  (.A(\proj__8.net24 ),
    .B(net91),
    .X(\proj__8.net10 ));
 sg13g2_and2_1 \proj__8.and3/_0_  (.A(net78),
    .B(\proj__8.net25 ),
    .X(\proj__8.net13 ));
 sg13g2_and2_1 \proj__8.and4/_0_  (.A(\proj__8.net26 ),
    .B(net78),
    .X(\proj__8.net14 ));
 sg13g2_and2_1 \proj__8.and5/_0_  (.A(\proj__8.net27 ),
    .B(net83),
    .X(\proj__8.net28 ));
 sg13g2_inv_1 \proj__8.not1/_0_  (.Y(\proj__8.net9 ),
    .A(\proj__8.net22 ));
 sg13g2_inv_1 \proj__8.not2/_0_  (.Y(\proj__8.net12 ),
    .A(\proj__8.net28 ));
 sg13g2_or2_1 \proj__8.or1/_0_  (.X(\proj__8.net16 ),
    .B(net75),
    .A(net72));
 sg13g2_or2_1 \proj__8.or2/_0_  (.X(\proj__8.net15 ),
    .B(net76),
    .A(net74));
 sg13g2_or2_1 \proj__8.or3/_0_  (.X(\proj__8.net22 ),
    .B(net76),
    .A(net75));
 sg13g2_xor2_1 \proj__8.xor1/_0_  (.B(net87),
    .A(net83),
    .X(\proj__8.net23 ));
 sg13g2_xor2_1 \proj__8.xor2/_0_  (.B(net83),
    .A(net80),
    .X(\proj__8.net27 ));
 sg13g2_xor2_1 \proj__8.xor3/_0_  (.B(net80),
    .A(net78),
    .X(\proj__8.net25 ));
 sg13g2_xor2_1 \proj__8.xor4/_0_  (.B(net78),
    .A(net77),
    .X(\proj__8.net26 ));
 sg13g2_xor2_1 \proj__8.xor5/_0_  (.B(net91),
    .A(net87),
    .X(\proj__8.net24 ));
 sg13g2_and2_1 \proj__9.and1/_0_  (.A(net88),
    .B(net92),
    .X(\proj__9.net16 ));
 sg13g2_and2_1 \proj__9.and2/_0_  (.A(net85),
    .B(\proj__9.net15 ),
    .X(\proj__9.net17 ));
 sg13g2_or2_1 \proj__9.or1/_0_  (.X(\proj__9.net9 ),
    .B(\proj__9.net17 ),
    .A(\proj__9.net16 ));
 sg13g2_xor2_1 \proj__9.xor1/_0_  (.B(net92),
    .A(net88),
    .X(\proj__9.net15 ));
 sg13g2_xor2_1 \proj__9.xor2/_0_  (.B(\proj__9.net15 ),
    .A(net85),
    .X(\proj__9.net8 ));
 sg13g2_buf_2 fanout72 (.A(net73),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(net3),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(net75),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(net2),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(net77),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(ui_in[5]),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(net79),
    .X(net78));
 sg13g2_buf_4 fanout79 (.X(net79),
    .A(ui_in[4]));
 sg13g2_buf_2 fanout80 (.A(net82),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(net82),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(ui_in[3]),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(net84),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(ui_in[2]),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(ui_in[2]),
    .X(net85));
 sg13g2_buf_1 fanout86 (.A(ui_in[2]),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(net90),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(net89),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(net90),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(ui_in[1]),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(net94),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(net94),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(net94),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(ui_in[0]),
    .X(net94));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[6]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[7]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[0]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(uio_in[1]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(uio_in[2]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(uio_in[3]),
    .X(net7));
 sg13g2_tielo \proj__1.and1/_0__8  (.L_LO(net8));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_1_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_1_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_1_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_1_1__leaf_clk_regs));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_4 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_177 ();
 sg13g2_decap_8 FILLER_18_184 ();
 sg13g2_decap_8 FILLER_18_191 ();
 sg13g2_decap_8 FILLER_18_198 ();
 sg13g2_decap_8 FILLER_18_205 ();
 sg13g2_decap_8 FILLER_18_212 ();
 sg13g2_decap_8 FILLER_18_219 ();
 sg13g2_decap_8 FILLER_18_226 ();
 sg13g2_decap_8 FILLER_18_233 ();
 sg13g2_decap_8 FILLER_18_240 ();
 sg13g2_decap_8 FILLER_18_247 ();
 sg13g2_decap_8 FILLER_18_254 ();
 sg13g2_decap_8 FILLER_18_261 ();
 sg13g2_decap_8 FILLER_18_268 ();
 sg13g2_decap_8 FILLER_18_275 ();
 sg13g2_decap_8 FILLER_18_282 ();
 sg13g2_decap_8 FILLER_18_289 ();
 sg13g2_decap_8 FILLER_18_296 ();
 sg13g2_decap_8 FILLER_18_303 ();
 sg13g2_decap_8 FILLER_18_310 ();
 sg13g2_decap_8 FILLER_18_317 ();
 sg13g2_decap_8 FILLER_18_324 ();
 sg13g2_decap_8 FILLER_18_331 ();
 sg13g2_decap_8 FILLER_18_338 ();
 sg13g2_decap_8 FILLER_18_345 ();
 sg13g2_decap_8 FILLER_18_352 ();
 sg13g2_decap_8 FILLER_18_359 ();
 sg13g2_decap_8 FILLER_18_366 ();
 sg13g2_decap_8 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_fill_2 FILLER_23_266 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_decap_8 FILLER_23_274 ();
 sg13g2_decap_8 FILLER_23_281 ();
 sg13g2_decap_8 FILLER_23_288 ();
 sg13g2_decap_8 FILLER_23_295 ();
 sg13g2_fill_1 FILLER_23_302 ();
 sg13g2_decap_8 FILLER_23_311 ();
 sg13g2_decap_8 FILLER_23_318 ();
 sg13g2_decap_8 FILLER_23_325 ();
 sg13g2_decap_8 FILLER_23_332 ();
 sg13g2_decap_8 FILLER_23_339 ();
 sg13g2_decap_8 FILLER_23_346 ();
 sg13g2_decap_8 FILLER_23_353 ();
 sg13g2_decap_8 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_374 ();
 sg13g2_decap_8 FILLER_23_381 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_4 FILLER_24_271 ();
 sg13g2_fill_2 FILLER_24_280 ();
 sg13g2_fill_1 FILLER_24_282 ();
 sg13g2_fill_1 FILLER_24_293 ();
 sg13g2_fill_1 FILLER_24_320 ();
 sg13g2_decap_8 FILLER_24_334 ();
 sg13g2_decap_8 FILLER_24_341 ();
 sg13g2_decap_4 FILLER_24_348 ();
 sg13g2_fill_1 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_358 ();
 sg13g2_decap_8 FILLER_24_365 ();
 sg13g2_decap_8 FILLER_24_372 ();
 sg13g2_decap_8 FILLER_24_379 ();
 sg13g2_decap_8 FILLER_24_386 ();
 sg13g2_decap_8 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_fill_2 FILLER_25_245 ();
 sg13g2_decap_4 FILLER_25_252 ();
 sg13g2_fill_2 FILLER_25_266 ();
 sg13g2_fill_1 FILLER_25_268 ();
 sg13g2_fill_1 FILLER_25_295 ();
 sg13g2_decap_4 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_310 ();
 sg13g2_decap_4 FILLER_25_317 ();
 sg13g2_decap_4 FILLER_25_339 ();
 sg13g2_decap_8 FILLER_25_353 ();
 sg13g2_decap_8 FILLER_25_360 ();
 sg13g2_decap_8 FILLER_25_367 ();
 sg13g2_decap_8 FILLER_25_374 ();
 sg13g2_decap_8 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_fill_2 FILLER_26_245 ();
 sg13g2_decap_4 FILLER_26_255 ();
 sg13g2_decap_4 FILLER_26_263 ();
 sg13g2_fill_1 FILLER_26_267 ();
 sg13g2_decap_8 FILLER_26_278 ();
 sg13g2_decap_4 FILLER_26_290 ();
 sg13g2_fill_1 FILLER_26_302 ();
 sg13g2_decap_8 FILLER_26_316 ();
 sg13g2_decap_4 FILLER_26_323 ();
 sg13g2_fill_1 FILLER_26_327 ();
 sg13g2_decap_4 FILLER_26_341 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_4 FILLER_27_175 ();
 sg13g2_fill_2 FILLER_27_179 ();
 sg13g2_decap_8 FILLER_27_185 ();
 sg13g2_decap_4 FILLER_27_201 ();
 sg13g2_fill_1 FILLER_27_208 ();
 sg13g2_decap_4 FILLER_27_214 ();
 sg13g2_fill_1 FILLER_27_218 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_fill_2 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_233 ();
 sg13g2_decap_8 FILLER_27_237 ();
 sg13g2_decap_4 FILLER_27_248 ();
 sg13g2_fill_2 FILLER_27_252 ();
 sg13g2_decap_4 FILLER_27_269 ();
 sg13g2_fill_1 FILLER_27_273 ();
 sg13g2_fill_1 FILLER_27_278 ();
 sg13g2_fill_2 FILLER_27_284 ();
 sg13g2_fill_2 FILLER_27_294 ();
 sg13g2_fill_2 FILLER_27_306 ();
 sg13g2_fill_1 FILLER_27_317 ();
 sg13g2_decap_8 FILLER_27_321 ();
 sg13g2_fill_2 FILLER_27_328 ();
 sg13g2_fill_1 FILLER_27_330 ();
 sg13g2_decap_4 FILLER_27_343 ();
 sg13g2_fill_1 FILLER_27_347 ();
 sg13g2_fill_2 FILLER_27_356 ();
 sg13g2_fill_1 FILLER_27_358 ();
 sg13g2_fill_2 FILLER_27_364 ();
 sg13g2_fill_1 FILLER_27_366 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_decap_8 FILLER_27_387 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_184 ();
 sg13g2_fill_2 FILLER_28_211 ();
 sg13g2_fill_1 FILLER_28_221 ();
 sg13g2_fill_2 FILLER_28_235 ();
 sg13g2_fill_2 FILLER_28_241 ();
 sg13g2_fill_2 FILLER_28_260 ();
 sg13g2_fill_1 FILLER_28_262 ();
 sg13g2_fill_2 FILLER_28_269 ();
 sg13g2_fill_1 FILLER_28_271 ();
 sg13g2_fill_2 FILLER_28_284 ();
 sg13g2_decap_8 FILLER_28_289 ();
 sg13g2_decap_8 FILLER_28_296 ();
 sg13g2_decap_4 FILLER_28_303 ();
 sg13g2_fill_2 FILLER_28_307 ();
 sg13g2_fill_1 FILLER_28_314 ();
 sg13g2_fill_1 FILLER_28_321 ();
 sg13g2_decap_8 FILLER_28_345 ();
 sg13g2_fill_2 FILLER_28_352 ();
 sg13g2_fill_1 FILLER_28_354 ();
 sg13g2_decap_8 FILLER_28_365 ();
 sg13g2_decap_8 FILLER_28_376 ();
 sg13g2_decap_8 FILLER_28_383 ();
 sg13g2_decap_8 FILLER_28_390 ();
 sg13g2_decap_8 FILLER_28_397 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_4 FILLER_29_175 ();
 sg13g2_fill_1 FILLER_29_179 ();
 sg13g2_decap_4 FILLER_29_200 ();
 sg13g2_fill_2 FILLER_29_204 ();
 sg13g2_decap_8 FILLER_29_209 ();
 sg13g2_fill_2 FILLER_29_216 ();
 sg13g2_fill_1 FILLER_29_218 ();
 sg13g2_decap_8 FILLER_29_230 ();
 sg13g2_decap_4 FILLER_29_237 ();
 sg13g2_fill_2 FILLER_29_241 ();
 sg13g2_fill_2 FILLER_29_248 ();
 sg13g2_fill_1 FILLER_29_250 ();
 sg13g2_decap_4 FILLER_29_256 ();
 sg13g2_fill_1 FILLER_29_260 ();
 sg13g2_decap_4 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_268 ();
 sg13g2_fill_1 FILLER_29_280 ();
 sg13g2_fill_1 FILLER_29_292 ();
 sg13g2_fill_2 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_307 ();
 sg13g2_fill_2 FILLER_29_316 ();
 sg13g2_fill_2 FILLER_29_323 ();
 sg13g2_fill_1 FILLER_29_325 ();
 sg13g2_fill_1 FILLER_29_340 ();
 sg13g2_decap_4 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_383 ();
 sg13g2_decap_8 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_4 FILLER_30_175 ();
 sg13g2_fill_2 FILLER_30_179 ();
 sg13g2_decap_8 FILLER_30_201 ();
 sg13g2_fill_2 FILLER_30_221 ();
 sg13g2_fill_1 FILLER_30_223 ();
 sg13g2_fill_2 FILLER_30_230 ();
 sg13g2_fill_2 FILLER_30_237 ();
 sg13g2_fill_1 FILLER_30_239 ();
 sg13g2_decap_4 FILLER_30_260 ();
 sg13g2_fill_1 FILLER_30_264 ();
 sg13g2_decap_4 FILLER_30_275 ();
 sg13g2_fill_2 FILLER_30_279 ();
 sg13g2_fill_1 FILLER_30_284 ();
 sg13g2_decap_4 FILLER_30_314 ();
 sg13g2_fill_2 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_30_342 ();
 sg13g2_decap_4 FILLER_30_349 ();
 sg13g2_fill_1 FILLER_30_353 ();
 sg13g2_decap_8 FILLER_30_372 ();
 sg13g2_decap_8 FILLER_30_379 ();
 sg13g2_decap_8 FILLER_30_386 ();
 sg13g2_decap_8 FILLER_30_393 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_fill_2 FILLER_31_182 ();
 sg13g2_fill_1 FILLER_31_184 ();
 sg13g2_fill_2 FILLER_31_190 ();
 sg13g2_decap_8 FILLER_31_221 ();
 sg13g2_fill_2 FILLER_31_228 ();
 sg13g2_fill_1 FILLER_31_240 ();
 sg13g2_fill_2 FILLER_31_246 ();
 sg13g2_decap_4 FILLER_31_259 ();
 sg13g2_fill_1 FILLER_31_263 ();
 sg13g2_fill_2 FILLER_31_267 ();
 sg13g2_decap_8 FILLER_31_275 ();
 sg13g2_decap_8 FILLER_31_282 ();
 sg13g2_fill_2 FILLER_31_305 ();
 sg13g2_decap_4 FILLER_31_318 ();
 sg13g2_fill_1 FILLER_31_338 ();
 sg13g2_decap_8 FILLER_31_348 ();
 sg13g2_fill_2 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_4 FILLER_32_189 ();
 sg13g2_fill_1 FILLER_32_193 ();
 sg13g2_decap_8 FILLER_32_214 ();
 sg13g2_decap_8 FILLER_32_221 ();
 sg13g2_decap_4 FILLER_32_228 ();
 sg13g2_fill_1 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_242 ();
 sg13g2_fill_2 FILLER_32_248 ();
 sg13g2_fill_1 FILLER_32_250 ();
 sg13g2_fill_1 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_306 ();
 sg13g2_decap_4 FILLER_32_313 ();
 sg13g2_fill_1 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_333 ();
 sg13g2_decap_8 FILLER_32_352 ();
 sg13g2_fill_2 FILLER_32_359 ();
 sg13g2_fill_1 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_32_367 ();
 sg13g2_decap_8 FILLER_32_394 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_4 FILLER_33_189 ();
 sg13g2_fill_2 FILLER_33_193 ();
 sg13g2_fill_1 FILLER_33_211 ();
 sg13g2_decap_8 FILLER_33_220 ();
 sg13g2_decap_4 FILLER_33_227 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_fill_2 FILLER_33_262 ();
 sg13g2_fill_2 FILLER_33_270 ();
 sg13g2_decap_4 FILLER_33_283 ();
 sg13g2_fill_1 FILLER_33_287 ();
 sg13g2_decap_4 FILLER_33_294 ();
 sg13g2_decap_4 FILLER_33_320 ();
 sg13g2_fill_1 FILLER_33_327 ();
 sg13g2_decap_8 FILLER_33_334 ();
 sg13g2_decap_4 FILLER_33_347 ();
 sg13g2_fill_2 FILLER_33_351 ();
 sg13g2_decap_4 FILLER_33_356 ();
 sg13g2_fill_1 FILLER_33_360 ();
 sg13g2_fill_2 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_4 FILLER_34_196 ();
 sg13g2_fill_2 FILLER_34_200 ();
 sg13g2_decap_4 FILLER_34_207 ();
 sg13g2_fill_2 FILLER_34_236 ();
 sg13g2_fill_1 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_253 ();
 sg13g2_fill_1 FILLER_34_260 ();
 sg13g2_fill_1 FILLER_34_266 ();
 sg13g2_decap_4 FILLER_34_280 ();
 sg13g2_fill_2 FILLER_34_284 ();
 sg13g2_decap_8 FILLER_34_292 ();
 sg13g2_decap_4 FILLER_34_299 ();
 sg13g2_fill_2 FILLER_34_320 ();
 sg13g2_fill_2 FILLER_34_335 ();
 sg13g2_fill_1 FILLER_34_337 ();
 sg13g2_decap_8 FILLER_34_397 ();
 sg13g2_decap_4 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_220 ();
 sg13g2_decap_4 FILLER_35_227 ();
 sg13g2_fill_2 FILLER_35_231 ();
 sg13g2_fill_1 FILLER_35_255 ();
 sg13g2_fill_2 FILLER_35_279 ();
 sg13g2_decap_4 FILLER_35_297 ();
 sg13g2_fill_2 FILLER_35_301 ();
 sg13g2_fill_2 FILLER_35_316 ();
 sg13g2_fill_1 FILLER_35_328 ();
 sg13g2_fill_2 FILLER_35_340 ();
 sg13g2_fill_2 FILLER_35_368 ();
 sg13g2_fill_1 FILLER_35_370 ();
 sg13g2_decap_4 FILLER_35_376 ();
 sg13g2_fill_2 FILLER_35_380 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_4 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_219 ();
 sg13g2_decap_4 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_237 ();
 sg13g2_decap_4 FILLER_36_256 ();
 sg13g2_fill_2 FILLER_36_260 ();
 sg13g2_fill_2 FILLER_36_270 ();
 sg13g2_fill_1 FILLER_36_272 ();
 sg13g2_decap_8 FILLER_36_277 ();
 sg13g2_fill_1 FILLER_36_284 ();
 sg13g2_decap_4 FILLER_36_293 ();
 sg13g2_fill_1 FILLER_36_297 ();
 sg13g2_fill_1 FILLER_36_311 ();
 sg13g2_fill_1 FILLER_36_342 ();
 sg13g2_decap_8 FILLER_36_369 ();
 sg13g2_decap_4 FILLER_36_376 ();
 sg13g2_fill_1 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_250 ();
 sg13g2_decap_8 FILLER_37_257 ();
 sg13g2_decap_8 FILLER_37_264 ();
 sg13g2_fill_2 FILLER_37_271 ();
 sg13g2_fill_1 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_279 ();
 sg13g2_decap_8 FILLER_37_286 ();
 sg13g2_decap_8 FILLER_37_293 ();
 sg13g2_decap_8 FILLER_37_300 ();
 sg13g2_fill_1 FILLER_37_307 ();
 sg13g2_fill_2 FILLER_37_312 ();
 sg13g2_decap_8 FILLER_37_328 ();
 sg13g2_decap_8 FILLER_37_335 ();
 sg13g2_decap_8 FILLER_37_342 ();
 sg13g2_decap_4 FILLER_37_349 ();
 sg13g2_fill_1 FILLER_37_353 ();
 sg13g2_decap_8 FILLER_37_362 ();
 sg13g2_decap_8 FILLER_37_369 ();
 sg13g2_decap_8 FILLER_37_376 ();
 sg13g2_decap_8 FILLER_37_383 ();
 sg13g2_decap_8 FILLER_37_390 ();
 sg13g2_decap_8 FILLER_37_397 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_decap_8 FILLER_38_257 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_fill_2 FILLER_38_278 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_fill_2 FILLER_38_293 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_2 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_decap_4 FILLER_38_308 ();
 sg13g2_decap_4 FILLER_38_316 ();
 sg13g2_decap_8 FILLER_38_324 ();
 sg13g2_fill_1 FILLER_38_331 ();
 sg13g2_decap_8 FILLER_38_337 ();
 sg13g2_decap_8 FILLER_38_344 ();
 sg13g2_decap_8 FILLER_38_351 ();
 sg13g2_decap_8 FILLER_38_358 ();
 sg13g2_decap_8 FILLER_38_365 ();
 sg13g2_decap_4 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net16;
 assign uio_oe[1] = net17;
 assign uio_oe[2] = net18;
 assign uio_oe[3] = net19;
 assign uio_oe[4] = net20;
 assign uio_oe[5] = net21;
 assign uio_oe[6] = net22;
 assign uio_oe[7] = net23;
 assign uio_out[0] = net24;
 assign uio_out[1] = net25;
 assign uio_out[2] = net26;
 assign uio_out[3] = net27;
 assign uio_out[4] = net28;
 assign uio_out[5] = net29;
 assign uio_out[6] = net30;
 assign uio_out[7] = net31;
endmodule

module tt_um_rebeccargb_vga_pride (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire clknet_0_clk;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire counter_clk;
 wire \flag.flag_abrosexual_inst.pix_x[0] ;
 wire \flag.flag_abrosexual_inst.pix_x[1] ;
 wire \flag.flag_abrosexual_inst.pix_x[2] ;
 wire \flag.flag_abrosexual_inst.pix_x[3] ;
 wire \flag.flag_abrosexual_inst.pix_x[4] ;
 wire \flag.flag_abrosexual_inst.pix_x[5] ;
 wire \flag.flag_abrosexual_inst.pix_x[6] ;
 wire \flag.flag_abrosexual_inst.pix_x[7] ;
 wire \flag.flag_abrosexual_inst.pix_x[8] ;
 wire \flag.flag_abrosexual_inst.pix_x[9] ;
 wire \flag.flag_abrosexual_inst.pix_y[0] ;
 wire \flag.flag_abrosexual_inst.pix_y[1] ;
 wire \flag.flag_abrosexual_inst.pix_y[2] ;
 wire \flag.flag_abrosexual_inst.pix_y[3] ;
 wire \flag.flag_abrosexual_inst.pix_y[4] ;
 wire \flag.flag_abrosexual_inst.pix_y[5] ;
 wire \flag.flag_abrosexual_inst.pix_y[6] ;
 wire \flag.flag_abrosexual_inst.pix_y[7] ;
 wire \flag.flag_abrosexual_inst.pix_y[8] ;
 wire hsync;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;

 sg13g2_inv_4 _3073_ (.A(_0025_),
    .Y(_0063_));
 sg13g2_inv_1 _3074_ (.Y(_0074_),
    .A(\counter[2] ));
 sg13g2_inv_1 _3075_ (.Y(_0085_),
    .A(\counter[1] ));
 sg13g2_inv_2 _3076_ (.Y(_0096_),
    .A(net861));
 sg13g2_inv_4 _3077_ (.A(net824),
    .Y(_0107_));
 sg13g2_inv_2 _3078_ (.Y(_0118_),
    .A(net860));
 sg13g2_inv_2 _3079_ (.Y(_0129_),
    .A(net839));
 sg13g2_inv_4 _3080_ (.A(net849),
    .Y(_0140_));
 sg13g2_inv_4 _3081_ (.A(net850),
    .Y(_0151_));
 sg13g2_inv_1 _3082_ (.Y(_0162_),
    .A(net833));
 sg13g2_inv_2 _3083_ (.Y(_0173_),
    .A(_0002_));
 sg13g2_inv_2 _3084_ (.Y(_0184_),
    .A(net815));
 sg13g2_inv_1 _3085_ (.Y(_0195_),
    .A(net818));
 sg13g2_inv_2 _3086_ (.Y(_0206_),
    .A(net808));
 sg13g2_inv_4 _3087_ (.A(net812),
    .Y(_0217_));
 sg13g2_inv_2 _3088_ (.Y(_0228_),
    .A(net797));
 sg13g2_inv_1 _3089_ (.Y(_0239_),
    .A(net804));
 sg13g2_inv_1 _3090_ (.Y(_0250_),
    .A(net786));
 sg13g2_inv_1 _3091_ (.Y(_0261_),
    .A(net790));
 sg13g2_inv_4 _3092_ (.A(net783),
    .Y(_0272_));
 sg13g2_inv_1 _3093_ (.Y(_0283_),
    .A(net7));
 sg13g2_inv_2 _3094_ (.Y(_0294_),
    .A(net828));
 sg13g2_inv_2 _3095_ (.Y(_0305_),
    .A(_0013_));
 sg13g2_inv_4 _3096_ (.A(net805),
    .Y(_0316_));
 sg13g2_inv_1 _3097_ (.Y(_0327_),
    .A(_0019_));
 sg13g2_inv_1 _3098_ (.Y(_0338_),
    .A(_0022_));
 sg13g2_inv_2 _3099_ (.Y(_0349_),
    .A(net821));
 sg13g2_nor2_2 _3100_ (.A(net4),
    .B(net5),
    .Y(_0360_));
 sg13g2_nor3_2 _3101_ (.A(net4),
    .B(net3),
    .C(net5),
    .Y(_0371_));
 sg13g2_nand2b_1 _3102_ (.Y(_0382_),
    .B(_0360_),
    .A_N(net3));
 sg13g2_nand2b_2 _3103_ (.Y(counter_clk),
    .B(_0371_),
    .A_N(net6));
 sg13g2_nor2b_2 _3104_ (.A(net856),
    .B_N(net852),
    .Y(_0403_));
 sg13g2_nor2_2 _3105_ (.A(_0096_),
    .B(_0118_),
    .Y(_0414_));
 sg13g2_nand2_2 _3106_ (.Y(_0425_),
    .A(net863),
    .B(net859));
 sg13g2_a21oi_2 _3107_ (.B1(_0002_),
    .Y(_0436_),
    .A2(_0425_),
    .A1(_0403_));
 sg13g2_nand2_1 _3108_ (.Y(_0447_),
    .A(net835),
    .B(_0436_));
 sg13g2_nand2_1 _3109_ (.Y(_0458_),
    .A(net850),
    .B(net834));
 sg13g2_nor2_2 _3110_ (.A(net863),
    .B(_0118_),
    .Y(_0469_));
 sg13g2_nand3_1 _3111_ (.B(_0403_),
    .C(_0469_),
    .A(net835),
    .Y(_0480_));
 sg13g2_inv_1 _3112_ (.Y(_0491_),
    .A(_0480_));
 sg13g2_nand3_1 _3113_ (.B(_0458_),
    .C(_0480_),
    .A(_0447_),
    .Y(_0502_));
 sg13g2_inv_1 _3114_ (.Y(_0513_),
    .A(_0502_));
 sg13g2_and2_1 _3115_ (.A(net853),
    .B(net856),
    .X(_0524_));
 sg13g2_nor2_1 _3116_ (.A(net63),
    .B(_0524_),
    .Y(_0535_));
 sg13g2_nor2_2 _3117_ (.A(_0140_),
    .B(_0535_),
    .Y(_0546_));
 sg13g2_and2_2 _3118_ (.A(net841),
    .B(net838),
    .X(_0557_));
 sg13g2_nand2_2 _3119_ (.Y(_0568_),
    .A(net842),
    .B(net838));
 sg13g2_and2_2 _3120_ (.A(net842),
    .B(net847),
    .X(_0579_));
 sg13g2_nand2_2 _3121_ (.Y(_0590_),
    .A(net841),
    .B(net847));
 sg13g2_nand2_2 _3122_ (.Y(_0601_),
    .A(net846),
    .B(_0557_));
 sg13g2_nor2b_2 _3123_ (.A(net850),
    .B_N(net846),
    .Y(_0612_));
 sg13g2_nand2_1 _3124_ (.Y(_0623_),
    .A(net846),
    .B(_0151_));
 sg13g2_nor4_2 _3125_ (.A(net61),
    .B(_0513_),
    .C(_0546_),
    .Y(_0001_),
    .D(_0601_));
 sg13g2_nor2_1 _3126_ (.A(net788),
    .B(_0272_),
    .Y(_0644_));
 sg13g2_nor2_1 _3127_ (.A(_0206_),
    .B(net776),
    .Y(_0655_));
 sg13g2_nand2_2 _3128_ (.Y(_0666_),
    .A(net807),
    .B(net804));
 sg13g2_nand2_2 _3129_ (.Y(_0677_),
    .A(net797),
    .B(net794));
 sg13g2_or2_1 _3130_ (.X(_0688_),
    .B(_0677_),
    .A(_0666_));
 sg13g2_a21oi_1 _3131_ (.A1(_0644_),
    .A2(_0688_),
    .Y(_0699_),
    .B1(net780));
 sg13g2_a21oi_2 _3132_ (.B1(net788),
    .Y(_0710_),
    .A2(net792),
    .A1(net797));
 sg13g2_nor2_1 _3133_ (.A(net807),
    .B(net803),
    .Y(_0721_));
 sg13g2_or2_2 _3134_ (.X(_0732_),
    .B(net804),
    .A(net807));
 sg13g2_nand2b_2 _3135_ (.Y(_0743_),
    .B(net793),
    .A_N(net797));
 sg13g2_o21ai_1 _3136_ (.B1(_0710_),
    .Y(_0754_),
    .A1(net767),
    .A2(_0743_));
 sg13g2_nand2_1 _3137_ (.Y(_0765_),
    .A(net783),
    .B(_0754_));
 sg13g2_nor2_2 _3138_ (.A(_0699_),
    .B(_0765_),
    .Y(_0000_));
 sg13g2_nor2_1 _3139_ (.A(\counter[6] ),
    .B(net867),
    .Y(_0786_));
 sg13g2_nand2b_1 _3140_ (.Y(_0797_),
    .B(net867),
    .A_N(net13));
 sg13g2_nor2b_2 _3141_ (.A(_0786_),
    .B_N(_0797_),
    .Y(_0808_));
 sg13g2_nand2b_2 _3142_ (.Y(_0819_),
    .B(_0797_),
    .A_N(_0786_));
 sg13g2_mux2_1 _3143_ (.A0(\counter[5] ),
    .A1(net12),
    .S(net867),
    .X(_0830_));
 sg13g2_mux2_2 _3144_ (.A0(\counter[4] ),
    .A1(net11),
    .S(net867),
    .X(_0841_));
 sg13g2_nor2b_1 _3145_ (.A(_0830_),
    .B_N(_0841_),
    .Y(_0852_));
 sg13g2_nand2b_1 _3146_ (.Y(_0863_),
    .B(_0841_),
    .A_N(_0830_));
 sg13g2_nand2_1 _3147_ (.Y(_0874_),
    .A(net9),
    .B(net2));
 sg13g2_o21ai_1 _3148_ (.B1(_0874_),
    .Y(_0885_),
    .A1(_0074_),
    .A2(net2));
 sg13g2_mux2_1 _3149_ (.A0(\counter[3] ),
    .A1(net10),
    .S(net867),
    .X(_0896_));
 sg13g2_nor2_2 _3150_ (.A(_0885_),
    .B(_0896_),
    .Y(_0907_));
 sg13g2_or2_2 _3151_ (.X(_0918_),
    .B(net750),
    .A(_0885_));
 sg13g2_nor2_1 _3152_ (.A(\counter[0] ),
    .B(net867),
    .Y(_0929_));
 sg13g2_a21oi_2 _3153_ (.B1(_0929_),
    .Y(_0940_),
    .A2(net867),
    .A1(_0283_));
 sg13g2_inv_2 _3154_ (.Y(_0951_),
    .A(_0940_));
 sg13g2_nand2_1 _3155_ (.Y(_0962_),
    .A(net8),
    .B(net867));
 sg13g2_o21ai_1 _3156_ (.B1(_0962_),
    .Y(_0973_),
    .A1(_0085_),
    .A2(net2));
 sg13g2_inv_2 _3157_ (.Y(_0984_),
    .A(_0973_));
 sg13g2_nor2_2 _3158_ (.A(_0951_),
    .B(_0973_),
    .Y(_0995_));
 sg13g2_nand2_2 _3159_ (.Y(_1006_),
    .A(_0940_),
    .B(_0984_));
 sg13g2_nor2_1 _3160_ (.A(_0918_),
    .B(_1006_),
    .Y(_1017_));
 sg13g2_nand2_2 _3161_ (.Y(_1028_),
    .A(_0907_),
    .B(_0995_));
 sg13g2_nand3_1 _3162_ (.B(_0852_),
    .C(_1017_),
    .A(_0808_),
    .Y(_1039_));
 sg13g2_nor2_2 _3163_ (.A(_0940_),
    .B(_0973_),
    .Y(_1050_));
 sg13g2_nand2_2 _3164_ (.Y(_1061_),
    .A(_0951_),
    .B(_0984_));
 sg13g2_nor2_2 _3165_ (.A(_0918_),
    .B(_1061_),
    .Y(_1072_));
 sg13g2_nand2_2 _3166_ (.Y(_1083_),
    .A(_0907_),
    .B(_1050_));
 sg13g2_nor3_2 _3167_ (.A(_0819_),
    .B(_0863_),
    .C(_1083_),
    .Y(_1094_));
 sg13g2_nand3_1 _3168_ (.B(_0852_),
    .C(_1072_),
    .A(_0808_),
    .Y(_1105_));
 sg13g2_or2_2 _3169_ (.X(_1116_),
    .B(_0841_),
    .A(_0830_));
 sg13g2_nand4_1 _3170_ (.B(_1039_),
    .C(_1105_),
    .A(_0808_),
    .Y(_1127_),
    .D(_1116_));
 sg13g2_nor2_2 _3171_ (.A(net787),
    .B(net792),
    .Y(_1138_));
 sg13g2_nor2_2 _3172_ (.A(_0129_),
    .B(net779),
    .Y(_1149_));
 sg13g2_nand2_1 _3173_ (.Y(_1160_),
    .A(net837),
    .B(net834));
 sg13g2_a21oi_1 _3174_ (.A1(_0579_),
    .A2(net760),
    .Y(_1171_),
    .B1(\hvsync_gen.vpos[9] ));
 sg13g2_o21ai_1 _3175_ (.B1(_1171_),
    .Y(_1182_),
    .A1(net780),
    .A2(_1138_));
 sg13g2_nand2b_2 _3176_ (.Y(_1193_),
    .B(_1127_),
    .A_N(_1182_));
 sg13g2_nor2_2 _3177_ (.A(_0940_),
    .B(_0984_),
    .Y(_1204_));
 sg13g2_nand2_1 _3178_ (.Y(_1215_),
    .A(_0951_),
    .B(_0973_));
 sg13g2_and2_2 _3179_ (.A(_0885_),
    .B(net750),
    .X(_1226_));
 sg13g2_nand2_2 _3180_ (.Y(_1237_),
    .A(_0885_),
    .B(net750));
 sg13g2_nor2_2 _3181_ (.A(_1215_),
    .B(_1237_),
    .Y(_1248_));
 sg13g2_nand2_2 _3182_ (.Y(_1259_),
    .A(_1204_),
    .B(_1226_));
 sg13g2_and2_1 _3183_ (.A(_0819_),
    .B(_0830_),
    .X(_1270_));
 sg13g2_and2_2 _3184_ (.A(_0841_),
    .B(_1270_),
    .X(_1281_));
 sg13g2_nand2_1 _3185_ (.Y(_1292_),
    .A(_0841_),
    .B(_1270_));
 sg13g2_nor2_2 _3186_ (.A(_1259_),
    .B(net665),
    .Y(_1303_));
 sg13g2_nor2_2 _3187_ (.A(net787),
    .B(net782),
    .Y(_1314_));
 sg13g2_nand2_2 _3188_ (.Y(_1325_),
    .A(net774),
    .B(_0272_));
 sg13g2_nor2_2 _3189_ (.A(net792),
    .B(net759),
    .Y(_1336_));
 sg13g2_nor2_2 _3190_ (.A(net825),
    .B(net818),
    .Y(_1347_));
 sg13g2_nand2_2 _3191_ (.Y(_1358_),
    .A(_0107_),
    .B(_0195_));
 sg13g2_nor2_1 _3192_ (.A(net815),
    .B(net817),
    .Y(_1369_));
 sg13g2_nor2_2 _3193_ (.A(net816),
    .B(_1358_),
    .Y(_1380_));
 sg13g2_nor2_2 _3194_ (.A(net816),
    .B(net812),
    .Y(_1391_));
 sg13g2_nor4_2 _3195_ (.A(net824),
    .B(net814),
    .C(net817),
    .Y(_1402_),
    .D(net811));
 sg13g2_or4_2 _3196_ (.A(net824),
    .B(net815),
    .C(net819),
    .D(net810),
    .X(_1413_));
 sg13g2_nor2_1 _3197_ (.A(net799),
    .B(net803),
    .Y(_1424_));
 sg13g2_nor2_2 _3198_ (.A(net798),
    .B(net794),
    .Y(_1435_));
 sg13g2_or2_2 _3199_ (.X(_1446_),
    .B(net794),
    .A(net799));
 sg13g2_nor2_1 _3200_ (.A(net804),
    .B(_1446_),
    .Y(_1457_));
 sg13g2_nand3_1 _3201_ (.B(net767),
    .C(_1435_),
    .A(_0644_),
    .Y(_1468_));
 sg13g2_o21ai_1 _3202_ (.B1(_0004_),
    .Y(_1479_),
    .A1(_1413_),
    .A2(_1468_));
 sg13g2_nor2b_1 _3203_ (.A(net793),
    .B_N(net788),
    .Y(_1490_));
 sg13g2_nor2b_2 _3204_ (.A(net803),
    .B_N(net797),
    .Y(_1501_));
 sg13g2_a21oi_2 _3205_ (.B1(net784),
    .Y(_1512_),
    .A2(_1501_),
    .A1(_1490_));
 sg13g2_nor2b_2 _3206_ (.A(net793),
    .B_N(net798),
    .Y(_1523_));
 sg13g2_nand2b_2 _3207_ (.Y(_1534_),
    .B(net797),
    .A_N(net794));
 sg13g2_and2_1 _3208_ (.A(net767),
    .B(_1391_),
    .X(_1545_));
 sg13g2_nand2_1 _3209_ (.Y(_1556_),
    .A(net767),
    .B(_1391_));
 sg13g2_nor2_1 _3210_ (.A(_0732_),
    .B(_1413_),
    .Y(_1567_));
 sg13g2_nand3_1 _3211_ (.B(_1402_),
    .C(_1523_),
    .A(net767),
    .Y(_1578_));
 sg13g2_nor2_1 _3212_ (.A(net774),
    .B(_1435_),
    .Y(_1589_));
 sg13g2_nand2_1 _3213_ (.Y(_1600_),
    .A(net787),
    .B(_1446_));
 sg13g2_a221oi_1 _3214_ (.B2(_1589_),
    .C1(net784),
    .B1(_1578_),
    .A1(_1490_),
    .Y(_1611_),
    .A2(_1501_));
 sg13g2_nand2_2 _3215_ (.Y(_1622_),
    .A(_0743_),
    .B(_1534_));
 sg13g2_inv_1 _3216_ (.Y(_1633_),
    .A(_1622_));
 sg13g2_a21oi_1 _3217_ (.A1(_0721_),
    .A2(_1402_),
    .Y(_1644_),
    .B1(_0228_));
 sg13g2_xnor2_1 _3218_ (.Y(_1655_),
    .A(_0014_),
    .B(_1644_));
 sg13g2_mux2_2 _3219_ (.A0(_1633_),
    .A1(_1655_),
    .S(net748),
    .X(_1665_));
 sg13g2_inv_1 _3220_ (.Y(_1676_),
    .A(net725));
 sg13g2_nor2_1 _3221_ (.A(net864),
    .B(net859),
    .Y(_1687_));
 sg13g2_or2_2 _3222_ (.X(_1698_),
    .B(net859),
    .A(net864));
 sg13g2_nor2_2 _3223_ (.A(net853),
    .B(net857),
    .Y(_1709_));
 sg13g2_nor4_2 _3224_ (.A(net863),
    .B(net859),
    .C(net852),
    .Y(_1720_),
    .D(net856));
 sg13g2_or4_2 _3225_ (.A(net863),
    .B(net859),
    .C(net852),
    .D(net856),
    .X(_1731_));
 sg13g2_and2_2 _3226_ (.A(net846),
    .B(net850),
    .X(_1742_));
 sg13g2_nand2_2 _3227_ (.Y(_1753_),
    .A(net848),
    .B(net851));
 sg13g2_nand2_2 _3228_ (.Y(_1764_),
    .A(net838),
    .B(_1742_));
 sg13g2_nand4_1 _3229_ (.B(net839),
    .C(net848),
    .A(net843),
    .Y(_1775_),
    .D(net851));
 sg13g2_a21oi_2 _3230_ (.B1(_1775_),
    .Y(_1786_),
    .A2(_1720_),
    .A1(net836));
 sg13g2_a21o_2 _3231_ (.A2(_1720_),
    .A1(net836),
    .B1(_1775_),
    .X(_1796_));
 sg13g2_nor2_1 _3232_ (.A(net772),
    .B(_1786_),
    .Y(_1807_));
 sg13g2_nand2_1 _3233_ (.Y(_1818_),
    .A(net829),
    .B(_1796_));
 sg13g2_nand2_1 _3234_ (.Y(_1829_),
    .A(net840),
    .B(net851));
 sg13g2_nand2_1 _3235_ (.Y(_1840_),
    .A(net843),
    .B(_1742_));
 sg13g2_xnor2_1 _3236_ (.Y(_1851_),
    .A(_0305_),
    .B(_1840_));
 sg13g2_nor3_1 _3237_ (.A(_0012_),
    .B(_1720_),
    .C(_1753_),
    .Y(_1862_));
 sg13g2_xnor2_1 _3238_ (.Y(_1873_),
    .A(net839),
    .B(_1862_));
 sg13g2_mux2_1 _3239_ (.A0(_1851_),
    .A1(_1873_),
    .S(net744),
    .X(_1884_));
 sg13g2_inv_1 _3240_ (.Y(_1895_),
    .A(net721));
 sg13g2_and4_1 _3241_ (.A(net866),
    .B(net771),
    .C(net725),
    .D(net721),
    .X(_1906_));
 sg13g2_nand4_1 _3242_ (.B(net771),
    .C(net724),
    .A(net861),
    .Y(_1917_),
    .D(net721));
 sg13g2_nand2_1 _3243_ (.Y(_1928_),
    .A(net824),
    .B(net817));
 sg13g2_nor2b_2 _3244_ (.A(_1347_),
    .B_N(net761),
    .Y(_1939_));
 sg13g2_nand2_2 _3245_ (.Y(_1950_),
    .A(_1358_),
    .B(net761));
 sg13g2_mux2_2 _3246_ (.A0(net817),
    .A1(_1939_),
    .S(net749),
    .X(_1961_));
 sg13g2_xnor2_1 _3247_ (.Y(_1972_),
    .A(net796),
    .B(_1567_));
 sg13g2_a21oi_1 _3248_ (.A1(_1512_),
    .A2(_1600_),
    .Y(_1982_),
    .B1(net798));
 sg13g2_a21o_2 _3249_ (.A2(_1972_),
    .A1(net748),
    .B1(_1982_),
    .X(_1993_));
 sg13g2_a21oi_2 _3250_ (.B1(_1982_),
    .Y(_2004_),
    .A2(_1972_),
    .A1(net748));
 sg13g2_nand2_2 _3251_ (.Y(_2015_),
    .A(_1961_),
    .B(_1993_));
 sg13g2_a22oi_1 _3252_ (.Y(_2026_),
    .B1(net721),
    .B2(net861),
    .A2(net724),
    .A1(net771));
 sg13g2_or3_1 _3253_ (.A(_1906_),
    .B(_2015_),
    .C(_2026_),
    .X(_2037_));
 sg13g2_o21ai_1 _3254_ (.B1(_1917_),
    .Y(_2048_),
    .A1(_2015_),
    .A2(_2026_));
 sg13g2_nor2_2 _3255_ (.A(_0096_),
    .B(net859),
    .Y(_2059_));
 sg13g2_nor2_2 _3256_ (.A(_0469_),
    .B(_2059_),
    .Y(_2069_));
 sg13g2_o21ai_1 _3257_ (.B1(_0338_),
    .Y(_2080_),
    .A1(net772),
    .A2(_1786_));
 sg13g2_mux2_2 _3258_ (.A0(_0022_),
    .A1(_2069_),
    .S(net744),
    .X(_2091_));
 sg13g2_o21ai_1 _3259_ (.B1(_2080_),
    .Y(_2102_),
    .A1(net743),
    .A2(_2069_));
 sg13g2_and2_1 _3260_ (.A(net721),
    .B(_2102_),
    .X(_2113_));
 sg13g2_nand2_1 _3261_ (.Y(_2124_),
    .A(net724),
    .B(_1961_));
 sg13g2_nand4_1 _3262_ (.B(net721),
    .C(_1961_),
    .A(net724),
    .Y(_2135_),
    .D(net719));
 sg13g2_xnor2_1 _3263_ (.Y(_2146_),
    .A(_2113_),
    .B(_2124_));
 sg13g2_nand2_1 _3264_ (.Y(_2157_),
    .A(_2048_),
    .B(_2146_));
 sg13g2_xnor2_1 _3265_ (.Y(_2168_),
    .A(_2048_),
    .B(_2146_));
 sg13g2_a21oi_2 _3266_ (.B1(_0151_),
    .Y(_2179_),
    .A2(_1796_),
    .A1(net832));
 sg13g2_o21ai_1 _3267_ (.B1(net851),
    .Y(_2189_),
    .A1(net772),
    .A2(_1786_));
 sg13g2_xnor2_1 _3268_ (.Y(_2200_),
    .A(_0016_),
    .B(_1731_));
 sg13g2_a21oi_2 _3269_ (.B1(_2179_),
    .Y(_2211_),
    .A2(_2200_),
    .A1(net744));
 sg13g2_nand4_1 _3270_ (.B(_1731_),
    .C(_1742_),
    .A(net829),
    .Y(_2222_),
    .D(_1775_));
 sg13g2_o21ai_1 _3271_ (.B1(_2222_),
    .Y(_2233_),
    .A1(net829),
    .A2(_1742_));
 sg13g2_xnor2_1 _3272_ (.Y(_2243_),
    .A(net840),
    .B(_2233_));
 sg13g2_a21oi_1 _3273_ (.A1(net832),
    .A2(_1796_),
    .Y(_2253_),
    .B1(_0173_));
 sg13g2_nand2_2 _3274_ (.Y(_2264_),
    .A(_0019_),
    .B(_1687_));
 sg13g2_xnor2_1 _3275_ (.Y(_2273_),
    .A(net854),
    .B(_2264_));
 sg13g2_a21oi_2 _3276_ (.B1(_2253_),
    .Y(_2283_),
    .A2(_2273_),
    .A1(net744));
 sg13g2_a21o_2 _3277_ (.A2(_2273_),
    .A1(net744),
    .B1(_2253_),
    .X(_2293_));
 sg13g2_nand2_2 _3278_ (.Y(_2303_),
    .A(net715),
    .B(net713));
 sg13g2_a21oi_1 _3279_ (.A1(net829),
    .A2(_1796_),
    .Y(_2313_),
    .B1(_0327_));
 sg13g2_xnor2_1 _3280_ (.Y(_2321_),
    .A(_0019_),
    .B(net762));
 sg13g2_a21oi_1 _3281_ (.A1(net744),
    .A2(_2321_),
    .Y(_2329_),
    .B1(_2313_));
 sg13g2_a21o_2 _3282_ (.A2(_2321_),
    .A1(net745),
    .B1(_2313_),
    .X(_2337_));
 sg13g2_nor2_1 _3283_ (.A(_0151_),
    .B(_1720_),
    .Y(_2342_));
 sg13g2_nor3_1 _3284_ (.A(net772),
    .B(_1786_),
    .C(_2342_),
    .Y(_2349_));
 sg13g2_o21ai_1 _3285_ (.B1(_0140_),
    .Y(_2352_),
    .A1(_2179_),
    .A2(_2349_));
 sg13g2_nand3b_1 _3286_ (.B(net848),
    .C(_2189_),
    .Y(_2353_),
    .A_N(_2349_));
 sg13g2_nand2_2 _3287_ (.Y(_2354_),
    .A(_2352_),
    .B(_2353_));
 sg13g2_and2_1 _3288_ (.A(_2352_),
    .B(_2353_),
    .X(_2355_));
 sg13g2_a21oi_2 _3289_ (.B1(_2337_),
    .Y(_2356_),
    .A2(_2353_),
    .A1(_2352_));
 sg13g2_nand2_1 _3290_ (.Y(_2357_),
    .A(net715),
    .B(net711));
 sg13g2_a21oi_2 _3291_ (.B1(_2293_),
    .Y(_2358_),
    .A2(_2353_),
    .A1(_2352_));
 sg13g2_nor2b_1 _3292_ (.A(_2303_),
    .B_N(_2356_),
    .Y(_2359_));
 sg13g2_xnor2_1 _3293_ (.Y(_2360_),
    .A(_2357_),
    .B(_2358_));
 sg13g2_xnor2_1 _3294_ (.Y(_2361_),
    .A(_2211_),
    .B(_2360_));
 sg13g2_o21ai_1 _3295_ (.B1(_2157_),
    .Y(_2362_),
    .A1(_2168_),
    .A2(_2361_));
 sg13g2_nand2b_1 _3296_ (.Y(_2363_),
    .B(net712),
    .A_N(_2135_));
 sg13g2_nand2_1 _3297_ (.Y(_2364_),
    .A(net721),
    .B(net712));
 sg13g2_mux2_1 _3298_ (.A0(net712),
    .A1(_2364_),
    .S(_2135_),
    .X(_2365_));
 sg13g2_xor2_1 _3299_ (.B(_2365_),
    .A(_2303_),
    .X(_2366_));
 sg13g2_nand2_1 _3300_ (.Y(_2367_),
    .A(_2362_),
    .B(_2366_));
 sg13g2_a21o_1 _3301_ (.A2(_2360_),
    .A1(_2113_),
    .B1(_2359_),
    .X(_2368_));
 sg13g2_a21oi_1 _3302_ (.A1(_2211_),
    .A2(_2360_),
    .Y(_2369_),
    .B1(_2359_));
 sg13g2_nand2_2 _3303_ (.Y(_2370_),
    .A(net722),
    .B(net714));
 sg13g2_nand2_2 _3304_ (.Y(_2371_),
    .A(_2283_),
    .B(net712));
 sg13g2_or2_1 _3305_ (.X(_2372_),
    .B(net678),
    .A(_2370_));
 sg13g2_xnor2_1 _3306_ (.Y(_2373_),
    .A(_2303_),
    .B(_2364_));
 sg13g2_nor2_1 _3307_ (.A(_2369_),
    .B(_2373_),
    .Y(_2374_));
 sg13g2_xor2_1 _3308_ (.B(_2373_),
    .A(_2369_),
    .X(_2375_));
 sg13g2_xnor2_1 _3309_ (.Y(_2376_),
    .A(_2368_),
    .B(_2375_));
 sg13g2_xnor2_1 _3310_ (.Y(_2377_),
    .A(_2362_),
    .B(_2366_));
 sg13g2_o21ai_1 _3311_ (.B1(_2367_),
    .Y(_2378_),
    .A1(_2376_),
    .A2(_2377_));
 sg13g2_nand2_1 _3312_ (.Y(_2379_),
    .A(net722),
    .B(_2283_));
 sg13g2_xnor2_1 _3313_ (.Y(_2380_),
    .A(net679),
    .B(_2379_));
 sg13g2_o21ai_1 _3314_ (.B1(_2363_),
    .Y(_2381_),
    .A1(_2303_),
    .A2(_2365_));
 sg13g2_nor2b_1 _3315_ (.A(_2380_),
    .B_N(_2381_),
    .Y(_2382_));
 sg13g2_nand2b_1 _3316_ (.Y(_2383_),
    .B(_2380_),
    .A_N(_2381_));
 sg13g2_nand2b_1 _3317_ (.Y(_2384_),
    .B(_2383_),
    .A_N(_2382_));
 sg13g2_nand2_2 _3318_ (.Y(_2385_),
    .A(net717),
    .B(_2354_));
 sg13g2_nor2b_1 _3319_ (.A(_2379_),
    .B_N(_2357_),
    .Y(_2386_));
 sg13g2_xnor2_1 _3320_ (.Y(_2387_),
    .A(_2385_),
    .B(_2386_));
 sg13g2_xnor2_1 _3321_ (.Y(_2388_),
    .A(_2384_),
    .B(_2387_));
 sg13g2_nand2_1 _3322_ (.Y(_2389_),
    .A(_2378_),
    .B(_2388_));
 sg13g2_nand2_2 _3323_ (.Y(_2390_),
    .A(_0021_),
    .B(_1347_));
 sg13g2_xnor2_1 _3324_ (.Y(_2391_),
    .A(net811),
    .B(_2390_));
 sg13g2_mux2_1 _3325_ (.A0(net809),
    .A1(_2391_),
    .S(net748),
    .X(_2392_));
 sg13g2_inv_4 _3326_ (.A(net709),
    .Y(_2393_));
 sg13g2_nand3_1 _3327_ (.B(_1512_),
    .C(_1600_),
    .A(_1358_),
    .Y(_2394_));
 sg13g2_xor2_1 _3328_ (.B(_2394_),
    .A(net813),
    .X(_2395_));
 sg13g2_xnor2_1 _3329_ (.Y(_2396_),
    .A(net813),
    .B(_2394_));
 sg13g2_nand2_1 _3330_ (.Y(_2397_),
    .A(net724),
    .B(_2395_));
 sg13g2_inv_1 _3331_ (.Y(_2398_),
    .A(_2397_));
 sg13g2_o21ai_1 _3332_ (.B1(_2397_),
    .Y(_2399_),
    .A1(_2004_),
    .A2(net710));
 sg13g2_nand2_1 _3333_ (.Y(_2400_),
    .A(_2015_),
    .B(_2398_));
 sg13g2_nand2_2 _3334_ (.Y(_2401_),
    .A(_2399_),
    .B(_2400_));
 sg13g2_a21oi_1 _3335_ (.A1(_2368_),
    .A2(_2375_),
    .Y(_2402_),
    .B1(_2374_));
 sg13g2_nor2_1 _3336_ (.A(_0316_),
    .B(_1413_),
    .Y(_2403_));
 sg13g2_xnor2_1 _3337_ (.Y(_2404_),
    .A(net806),
    .B(_1402_));
 sg13g2_mux2_1 _3338_ (.A0(net806),
    .A1(_2404_),
    .S(net748),
    .X(_2405_));
 sg13g2_nor2_1 _3339_ (.A(_1676_),
    .B(net707),
    .Y(_2406_));
 sg13g2_nor2_2 _3340_ (.A(_2004_),
    .B(net707),
    .Y(_2407_));
 sg13g2_nor2_2 _3341_ (.A(_1676_),
    .B(net709),
    .Y(_2408_));
 sg13g2_nand2_1 _3342_ (.Y(_2409_),
    .A(_2407_),
    .B(_2408_));
 sg13g2_xnor2_1 _3343_ (.Y(_2410_),
    .A(_2407_),
    .B(_2408_));
 sg13g2_nor2_2 _3344_ (.A(_2004_),
    .B(_2396_),
    .Y(_2411_));
 sg13g2_nand2_1 _3345_ (.Y(_2412_),
    .A(_2408_),
    .B(_2411_));
 sg13g2_xor2_1 _3346_ (.B(_2412_),
    .A(_2410_),
    .X(_2413_));
 sg13g2_xnor2_1 _3347_ (.Y(_2414_),
    .A(net776),
    .B(_2403_));
 sg13g2_mux2_2 _3348_ (.A0(net801),
    .A1(_2414_),
    .S(net748),
    .X(_2415_));
 sg13g2_inv_1 _3349_ (.Y(_2416_),
    .A(net704));
 sg13g2_nor2_2 _3350_ (.A(net706),
    .B(net704),
    .Y(_2417_));
 sg13g2_xnor2_1 _3351_ (.Y(_2418_),
    .A(_2407_),
    .B(net704));
 sg13g2_xor2_1 _3352_ (.B(_2418_),
    .A(_2408_),
    .X(_2419_));
 sg13g2_nand2_1 _3353_ (.Y(_2420_),
    .A(_2413_),
    .B(_2419_));
 sg13g2_xnor2_1 _3354_ (.Y(_2421_),
    .A(_2413_),
    .B(_2419_));
 sg13g2_or2_1 _3355_ (.X(_2422_),
    .B(_2421_),
    .A(_2402_));
 sg13g2_xor2_1 _3356_ (.B(_2421_),
    .A(_2402_),
    .X(_2423_));
 sg13g2_nand2b_1 _3357_ (.Y(_2424_),
    .B(_2423_),
    .A_N(_2401_));
 sg13g2_xor2_1 _3358_ (.B(_2423_),
    .A(_2401_),
    .X(_2425_));
 sg13g2_xnor2_1 _3359_ (.Y(_2426_),
    .A(_2378_),
    .B(_2388_));
 sg13g2_o21ai_1 _3360_ (.B1(_2389_),
    .Y(_2427_),
    .A1(_2425_),
    .A2(_2426_));
 sg13g2_and2_1 _3361_ (.A(net722),
    .B(net717),
    .X(_2428_));
 sg13g2_o21ai_1 _3362_ (.B1(_2372_),
    .Y(_2429_),
    .A1(_2379_),
    .A2(_2385_));
 sg13g2_nor2b_1 _3363_ (.A(_2409_),
    .B_N(_2429_),
    .Y(_2430_));
 sg13g2_xnor2_1 _3364_ (.Y(_2431_),
    .A(_2409_),
    .B(_2429_));
 sg13g2_o21ai_1 _3365_ (.B1(_2420_),
    .Y(_2432_),
    .A1(_2410_),
    .A2(_2412_));
 sg13g2_xor2_1 _3366_ (.B(_2432_),
    .A(_2431_),
    .X(_2433_));
 sg13g2_and3_1 _3367_ (.X(_2434_),
    .A(net714),
    .B(_2358_),
    .C(_2428_));
 sg13g2_a22oi_1 _3368_ (.Y(_2435_),
    .B1(_2358_),
    .B2(net721),
    .A2(net715),
    .A1(net717));
 sg13g2_nor2_1 _3369_ (.A(_2434_),
    .B(_2435_),
    .Y(_2436_));
 sg13g2_a21o_1 _3370_ (.A2(_2387_),
    .A1(_2383_),
    .B1(_2382_),
    .X(_2437_));
 sg13g2_and2_1 _3371_ (.A(_2436_),
    .B(_2437_),
    .X(_2438_));
 sg13g2_xor2_1 _3372_ (.B(_2437_),
    .A(_2436_),
    .X(_2439_));
 sg13g2_xor2_1 _3373_ (.B(_2439_),
    .A(_2433_),
    .X(_2440_));
 sg13g2_nand2_1 _3374_ (.Y(_2441_),
    .A(_2427_),
    .B(_2440_));
 sg13g2_a22oi_1 _3375_ (.Y(_2442_),
    .B1(_2418_),
    .B2(_2408_),
    .A2(_2417_),
    .A1(_1993_));
 sg13g2_a21oi_2 _3376_ (.B1(_2442_),
    .Y(_2443_),
    .A2(_2424_),
    .A1(_2422_));
 sg13g2_nand3_1 _3377_ (.B(_2424_),
    .C(_2442_),
    .A(_2422_),
    .Y(_2444_));
 sg13g2_nand2b_1 _3378_ (.Y(_2445_),
    .B(_2444_),
    .A_N(_2443_));
 sg13g2_xnor2_1 _3379_ (.Y(_2446_),
    .A(_2427_),
    .B(_2440_));
 sg13g2_o21ai_1 _3380_ (.B1(_2441_),
    .Y(_2447_),
    .A1(_2445_),
    .A2(_2446_));
 sg13g2_nand3_1 _3381_ (.B(_1993_),
    .C(_2417_),
    .A(net725),
    .Y(_2448_));
 sg13g2_a21oi_1 _3382_ (.A1(_2431_),
    .A2(_2432_),
    .Y(_2449_),
    .B1(_2430_));
 sg13g2_nor2_1 _3383_ (.A(_2448_),
    .B(_2449_),
    .Y(_2450_));
 sg13g2_xor2_1 _3384_ (.B(_2449_),
    .A(_2448_),
    .X(_2451_));
 sg13g2_inv_1 _3385_ (.Y(_2452_),
    .A(_2451_));
 sg13g2_a21o_1 _3386_ (.A2(_2439_),
    .A1(_2433_),
    .B1(_2438_),
    .X(_2453_));
 sg13g2_a21oi_1 _3387_ (.A1(net714),
    .A2(net679),
    .Y(_2454_),
    .B1(_2428_));
 sg13g2_nand3_1 _3388_ (.B(net679),
    .C(_2428_),
    .A(net714),
    .Y(_2455_));
 sg13g2_nand2b_1 _3389_ (.Y(_2456_),
    .B(_2455_),
    .A_N(_2454_));
 sg13g2_nor2_1 _3390_ (.A(_2434_),
    .B(_2456_),
    .Y(_2457_));
 sg13g2_o21ai_1 _3391_ (.B1(_1993_),
    .Y(_2458_),
    .A1(_2406_),
    .A2(_2416_));
 sg13g2_o21ai_1 _3392_ (.B1(_2458_),
    .Y(_2459_),
    .A1(_1993_),
    .A2(_2406_));
 sg13g2_inv_1 _3393_ (.Y(_2460_),
    .A(_2459_));
 sg13g2_xor2_1 _3394_ (.B(_2459_),
    .A(_2457_),
    .X(_2461_));
 sg13g2_nand2b_1 _3395_ (.Y(_2462_),
    .B(_2453_),
    .A_N(_2461_));
 sg13g2_xor2_1 _3396_ (.B(_2461_),
    .A(_2453_),
    .X(_2463_));
 sg13g2_xnor2_1 _3397_ (.Y(_2464_),
    .A(_2452_),
    .B(_2463_));
 sg13g2_nor2b_1 _3398_ (.A(_2464_),
    .B_N(_2447_),
    .Y(_2465_));
 sg13g2_xnor2_1 _3399_ (.Y(_2466_),
    .A(_2447_),
    .B(_2464_));
 sg13g2_a21o_1 _3400_ (.A2(_2466_),
    .A1(_2443_),
    .B1(_2465_),
    .X(_2467_));
 sg13g2_o21ai_1 _3401_ (.B1(_2462_),
    .Y(_2468_),
    .A1(_2452_),
    .A2(_2463_));
 sg13g2_a21o_1 _3402_ (.A2(_2417_),
    .A1(net725),
    .B1(_2458_),
    .X(_2469_));
 sg13g2_a21oi_1 _3403_ (.A1(_2457_),
    .A2(_2460_),
    .Y(_2470_),
    .B1(_2434_));
 sg13g2_or3_1 _3404_ (.A(_1676_),
    .B(_2407_),
    .C(net705),
    .X(_2471_));
 sg13g2_nor2_2 _3405_ (.A(net722),
    .B(net714),
    .Y(_2472_));
 sg13g2_nand2_1 _3406_ (.Y(_2473_),
    .A(_2354_),
    .B(_2370_));
 sg13g2_o21ai_1 _3407_ (.B1(_2455_),
    .Y(_2474_),
    .A1(_2472_),
    .A2(_2473_));
 sg13g2_nand2b_1 _3408_ (.Y(_2475_),
    .B(_2474_),
    .A_N(_2471_));
 sg13g2_xor2_1 _3409_ (.B(_2474_),
    .A(_2471_),
    .X(_2476_));
 sg13g2_xor2_1 _3410_ (.B(_2476_),
    .A(_2470_),
    .X(_2477_));
 sg13g2_nand2b_1 _3411_ (.Y(_2478_),
    .B(_2477_),
    .A_N(_2469_));
 sg13g2_xnor2_1 _3412_ (.Y(_2479_),
    .A(_2469_),
    .B(_2477_));
 sg13g2_and2_1 _3413_ (.A(_2468_),
    .B(_2479_),
    .X(_2480_));
 sg13g2_or2_1 _3414_ (.X(_2481_),
    .B(_2479_),
    .A(_2468_));
 sg13g2_nand2b_1 _3415_ (.Y(_2482_),
    .B(_2481_),
    .A_N(_2480_));
 sg13g2_xnor2_1 _3416_ (.Y(_2483_),
    .A(_2450_),
    .B(_2482_));
 sg13g2_nand2_1 _3417_ (.Y(_2484_),
    .A(_2467_),
    .B(_2483_));
 sg13g2_mux2_2 _3418_ (.A0(_0023_),
    .A1(_1950_),
    .S(net748),
    .X(_2485_));
 sg13g2_nor2_1 _3419_ (.A(net704),
    .B(_2485_),
    .Y(_2486_));
 sg13g2_nor2_2 _3420_ (.A(_0107_),
    .B(_2004_),
    .Y(_2487_));
 sg13g2_and2_1 _3421_ (.A(_2486_),
    .B(_2487_),
    .X(_2488_));
 sg13g2_o21ai_1 _3422_ (.B1(_2015_),
    .Y(_2489_),
    .A1(_1906_),
    .A2(_2026_));
 sg13g2_and2_1 _3423_ (.A(_2037_),
    .B(_2489_),
    .X(_2490_));
 sg13g2_and3_1 _3424_ (.X(_2491_),
    .A(_2037_),
    .B(_2488_),
    .C(_2489_));
 sg13g2_nand3_1 _3425_ (.B(_2488_),
    .C(_2489_),
    .A(_2037_),
    .Y(_2492_));
 sg13g2_nand2_1 _3426_ (.Y(_2493_),
    .A(_2102_),
    .B(net716));
 sg13g2_nand2_2 _3427_ (.Y(_2494_),
    .A(net718),
    .B(net713));
 sg13g2_inv_1 _3428_ (.Y(_2495_),
    .A(_2494_));
 sg13g2_nand2_2 _3429_ (.Y(_2496_),
    .A(net718),
    .B(net711));
 sg13g2_nor2_1 _3430_ (.A(_2337_),
    .B(_2494_),
    .Y(_2497_));
 sg13g2_nand2_2 _3431_ (.Y(_2498_),
    .A(_2354_),
    .B(_2497_));
 sg13g2_xor2_1 _3432_ (.B(_2494_),
    .A(_2356_),
    .X(_2499_));
 sg13g2_xor2_1 _3433_ (.B(_2499_),
    .A(_2493_),
    .X(_2500_));
 sg13g2_a21o_1 _3434_ (.A2(_2489_),
    .A1(_2037_),
    .B1(_2488_),
    .X(_2501_));
 sg13g2_nand3_1 _3435_ (.B(_2500_),
    .C(_2501_),
    .A(_2492_),
    .Y(_2502_));
 sg13g2_a21o_1 _3436_ (.A2(_2501_),
    .A1(_2500_),
    .B1(_2491_),
    .X(_2503_));
 sg13g2_xor2_1 _3437_ (.B(_2361_),
    .A(_2168_),
    .X(_2504_));
 sg13g2_nand2_1 _3438_ (.Y(_2505_),
    .A(_2503_),
    .B(_2504_));
 sg13g2_xnor2_1 _3439_ (.Y(_2506_),
    .A(_2113_),
    .B(_2360_));
 sg13g2_xnor2_1 _3440_ (.Y(_2507_),
    .A(_2503_),
    .B(_2504_));
 sg13g2_o21ai_1 _3441_ (.B1(_2505_),
    .Y(_2508_),
    .A1(_2506_),
    .A2(_2507_));
 sg13g2_xor2_1 _3442_ (.B(_2377_),
    .A(_2376_),
    .X(_2509_));
 sg13g2_nand2_1 _3443_ (.Y(_2510_),
    .A(_2508_),
    .B(_2509_));
 sg13g2_xnor2_1 _3444_ (.Y(_2511_),
    .A(_2508_),
    .B(_2509_));
 sg13g2_xnor2_1 _3445_ (.Y(_2512_),
    .A(_2124_),
    .B(_2411_));
 sg13g2_nand2_1 _3446_ (.Y(_2513_),
    .A(_2048_),
    .B(_2512_));
 sg13g2_mux2_2 _3447_ (.A0(_0206_),
    .A1(_2404_),
    .S(net748),
    .X(_2514_));
 sg13g2_xnor2_1 _3448_ (.Y(_2515_),
    .A(_2048_),
    .B(_2512_));
 sg13g2_o21ai_1 _3449_ (.B1(_2513_),
    .Y(_2516_),
    .A1(_2514_),
    .A2(_2515_));
 sg13g2_o21ai_1 _3450_ (.B1(_2498_),
    .Y(_2517_),
    .A1(_2493_),
    .A2(_2499_));
 sg13g2_nand2b_1 _3451_ (.Y(_2518_),
    .B(_2517_),
    .A_N(_2400_));
 sg13g2_xor2_1 _3452_ (.B(_2517_),
    .A(_2400_),
    .X(_2519_));
 sg13g2_nand2b_1 _3453_ (.Y(_2520_),
    .B(_2516_),
    .A_N(_2519_));
 sg13g2_xor2_1 _3454_ (.B(_2519_),
    .A(_2516_),
    .X(_2521_));
 sg13g2_o21ai_1 _3455_ (.B1(_2510_),
    .Y(_2522_),
    .A1(_2511_),
    .A2(_2521_));
 sg13g2_xor2_1 _3456_ (.B(_2426_),
    .A(_2425_),
    .X(_2523_));
 sg13g2_nand2_1 _3457_ (.Y(_2524_),
    .A(_2522_),
    .B(_2523_));
 sg13g2_nand2_2 _3458_ (.Y(_2525_),
    .A(_2518_),
    .B(_2520_));
 sg13g2_nand2_1 _3459_ (.Y(_2526_),
    .A(_2417_),
    .B(_2525_));
 sg13g2_xnor2_1 _3460_ (.Y(_2527_),
    .A(_2417_),
    .B(_2525_));
 sg13g2_xnor2_1 _3461_ (.Y(_2528_),
    .A(_2522_),
    .B(_2523_));
 sg13g2_o21ai_1 _3462_ (.B1(_2524_),
    .Y(_2529_),
    .A1(_2527_),
    .A2(_2528_));
 sg13g2_xor2_1 _3463_ (.B(_2446_),
    .A(_2445_),
    .X(_2530_));
 sg13g2_nand2_1 _3464_ (.Y(_2531_),
    .A(_2529_),
    .B(_2530_));
 sg13g2_xnor2_1 _3465_ (.Y(_2532_),
    .A(_2529_),
    .B(_2530_));
 sg13g2_o21ai_1 _3466_ (.B1(_2531_),
    .Y(_2533_),
    .A1(_2526_),
    .A2(_2532_));
 sg13g2_xnor2_1 _3467_ (.Y(_2534_),
    .A(_2443_),
    .B(_2466_));
 sg13g2_nor2b_1 _3468_ (.A(_2534_),
    .B_N(_2533_),
    .Y(_2535_));
 sg13g2_or2_1 _3469_ (.X(_2536_),
    .B(_2534_),
    .A(_2533_));
 sg13g2_nand2_1 _3470_ (.Y(_2537_),
    .A(_2533_),
    .B(_2534_));
 sg13g2_nand2_1 _3471_ (.Y(_2538_),
    .A(_2536_),
    .B(_2537_));
 sg13g2_xor2_1 _3472_ (.B(_2532_),
    .A(_2526_),
    .X(_2539_));
 sg13g2_nand2_2 _3473_ (.Y(_2540_),
    .A(net862),
    .B(_2354_));
 sg13g2_inv_2 _3474_ (.Y(_2541_),
    .A(_2540_));
 sg13g2_a21oi_1 _3475_ (.A1(_2352_),
    .A2(_2353_),
    .Y(_2542_),
    .B1(_2091_));
 sg13g2_nand2_1 _3476_ (.Y(_2543_),
    .A(net861),
    .B(net716));
 sg13g2_nand3_1 _3477_ (.B(net716),
    .C(_2542_),
    .A(net861),
    .Y(_2544_));
 sg13g2_xor2_1 _3478_ (.B(_2543_),
    .A(net677),
    .X(_2545_));
 sg13g2_xor2_1 _3479_ (.B(_2545_),
    .A(_2496_),
    .X(_2546_));
 sg13g2_nor2_2 _3480_ (.A(net821),
    .B(net706),
    .Y(_2547_));
 sg13g2_nand2b_1 _3481_ (.Y(_2548_),
    .B(_2486_),
    .A_N(_2547_));
 sg13g2_xnor2_1 _3482_ (.Y(_2549_),
    .A(_2487_),
    .B(_2548_));
 sg13g2_nor4_2 _3483_ (.A(net820),
    .B(net706),
    .C(net704),
    .Y(_2550_),
    .D(_2485_));
 sg13g2_nor2b_1 _3484_ (.A(_2487_),
    .B_N(_2550_),
    .Y(_2551_));
 sg13g2_a21o_1 _3485_ (.A2(_2549_),
    .A1(_2546_),
    .B1(_2551_),
    .X(_2552_));
 sg13g2_a21o_1 _3486_ (.A2(_2501_),
    .A1(_2492_),
    .B1(_2500_),
    .X(_2553_));
 sg13g2_and3_1 _3487_ (.X(_2554_),
    .A(_2502_),
    .B(_2552_),
    .C(_2553_));
 sg13g2_nand3_1 _3488_ (.B(_2552_),
    .C(_2553_),
    .A(_2502_),
    .Y(_2555_));
 sg13g2_a21oi_1 _3489_ (.A1(_2502_),
    .A2(_2553_),
    .Y(_2556_),
    .B1(_2552_));
 sg13g2_o21ai_1 _3490_ (.B1(_2544_),
    .Y(_2557_),
    .A1(_2496_),
    .A2(_2545_));
 sg13g2_nand2_1 _3491_ (.Y(_2558_),
    .A(_2500_),
    .B(_2557_));
 sg13g2_xnor2_1 _3492_ (.Y(_2559_),
    .A(_2500_),
    .B(_2557_));
 sg13g2_nand2_1 _3493_ (.Y(_2560_),
    .A(_2293_),
    .B(_2496_));
 sg13g2_o21ai_1 _3494_ (.B1(_2560_),
    .Y(_2561_),
    .A1(_2497_),
    .A2(net677));
 sg13g2_xnor2_1 _3495_ (.Y(_2562_),
    .A(_2559_),
    .B(_2561_));
 sg13g2_or3_1 _3496_ (.A(_2554_),
    .B(_2556_),
    .C(_2562_),
    .X(_2563_));
 sg13g2_o21ai_1 _3497_ (.B1(_2555_),
    .Y(_2564_),
    .A1(_2556_),
    .A2(_2562_));
 sg13g2_xnor2_1 _3498_ (.Y(_2565_),
    .A(_2506_),
    .B(_2507_));
 sg13g2_nand2b_1 _3499_ (.Y(_2566_),
    .B(_2564_),
    .A_N(_2565_));
 sg13g2_xor2_1 _3500_ (.B(_2565_),
    .A(_2564_),
    .X(_2567_));
 sg13g2_nand3_1 _3501_ (.B(net716),
    .C(_2487_),
    .A(net861),
    .Y(_2568_));
 sg13g2_nand4_1 _3502_ (.B(net716),
    .C(_2487_),
    .A(net861),
    .Y(_2569_),
    .D(_2490_));
 sg13g2_nand2_2 _3503_ (.Y(_2570_),
    .A(_2395_),
    .B(_2416_));
 sg13g2_xor2_1 _3504_ (.B(_2568_),
    .A(_2490_),
    .X(_2571_));
 sg13g2_o21ai_1 _3505_ (.B1(_2569_),
    .Y(_2572_),
    .A1(_2570_),
    .A2(_2571_));
 sg13g2_o21ai_1 _3506_ (.B1(_2558_),
    .Y(_2573_),
    .A1(_2559_),
    .A2(_2561_));
 sg13g2_xnor2_1 _3507_ (.Y(_2574_),
    .A(_2514_),
    .B(_2515_));
 sg13g2_nor2b_1 _3508_ (.A(_2574_),
    .B_N(_2573_),
    .Y(_2575_));
 sg13g2_xnor2_1 _3509_ (.Y(_2576_),
    .A(_2573_),
    .B(_2574_));
 sg13g2_xnor2_1 _3510_ (.Y(_2577_),
    .A(_2572_),
    .B(_2576_));
 sg13g2_o21ai_1 _3511_ (.B1(_2566_),
    .Y(_2578_),
    .A1(_2567_),
    .A2(_2577_));
 sg13g2_xor2_1 _3512_ (.B(_2521_),
    .A(_2511_),
    .X(_2579_));
 sg13g2_nand2_1 _3513_ (.Y(_2580_),
    .A(_2578_),
    .B(_2579_));
 sg13g2_xnor2_1 _3514_ (.Y(_2581_),
    .A(_2578_),
    .B(_2579_));
 sg13g2_a21oi_1 _3515_ (.A1(_2572_),
    .A2(_2576_),
    .Y(_2582_),
    .B1(_2575_));
 sg13g2_nor2_1 _3516_ (.A(net709),
    .B(net704),
    .Y(_2583_));
 sg13g2_nor2b_1 _3517_ (.A(_2582_),
    .B_N(_2583_),
    .Y(_2584_));
 sg13g2_xnor2_1 _3518_ (.Y(_2585_),
    .A(_2582_),
    .B(_2583_));
 sg13g2_xnor2_1 _3519_ (.Y(_2586_),
    .A(_2398_),
    .B(_2585_));
 sg13g2_o21ai_1 _3520_ (.B1(_2580_),
    .Y(_2587_),
    .A1(_2581_),
    .A2(_2586_));
 sg13g2_xnor2_1 _3521_ (.Y(_2588_),
    .A(_2527_),
    .B(_2528_));
 sg13g2_nor2b_1 _3522_ (.A(_2588_),
    .B_N(_2587_),
    .Y(_2589_));
 sg13g2_a21oi_2 _3523_ (.B1(_2584_),
    .Y(_2590_),
    .A2(_2585_),
    .A1(_2398_));
 sg13g2_xor2_1 _3524_ (.B(_2588_),
    .A(_2587_),
    .X(_2591_));
 sg13g2_nor2_1 _3525_ (.A(_2590_),
    .B(_2591_),
    .Y(_2592_));
 sg13g2_nor3_2 _3526_ (.A(_2539_),
    .B(_2589_),
    .C(_2592_),
    .Y(_2593_));
 sg13g2_or2_1 _3527_ (.X(_2594_),
    .B(_2485_),
    .A(net706));
 sg13g2_nand2b_1 _3528_ (.Y(_2595_),
    .B(net771),
    .A_N(net704));
 sg13g2_a21oi_2 _3529_ (.B1(_2550_),
    .Y(_2596_),
    .A2(_2595_),
    .A1(_2594_));
 sg13g2_nor2_2 _3530_ (.A(net709),
    .B(_2485_),
    .Y(_2597_));
 sg13g2_nor2_1 _3531_ (.A(net820),
    .B(net709),
    .Y(_2598_));
 sg13g2_and2_1 _3532_ (.A(_2547_),
    .B(_2597_),
    .X(_2599_));
 sg13g2_and2_1 _3533_ (.A(_2596_),
    .B(_2599_),
    .X(_2600_));
 sg13g2_nand2_2 _3534_ (.Y(_2601_),
    .A(net719),
    .B(net718));
 sg13g2_and2_2 _3535_ (.A(net862),
    .B(net718),
    .X(_2602_));
 sg13g2_nand2_2 _3536_ (.Y(_2603_),
    .A(net862),
    .B(net718));
 sg13g2_xor2_1 _3537_ (.B(_2601_),
    .A(_2540_),
    .X(_2604_));
 sg13g2_xor2_1 _3538_ (.B(_2599_),
    .A(_2596_),
    .X(_2605_));
 sg13g2_a21oi_2 _3539_ (.B1(_2600_),
    .Y(_2606_),
    .A2(_2605_),
    .A1(_2604_));
 sg13g2_xnor2_1 _3540_ (.Y(_2607_),
    .A(_2546_),
    .B(_2549_));
 sg13g2_nor2_1 _3541_ (.A(_2606_),
    .B(_2607_),
    .Y(_2608_));
 sg13g2_xnor2_1 _3542_ (.Y(_2609_),
    .A(net713),
    .B(_2496_));
 sg13g2_nand2_1 _3543_ (.Y(_2610_),
    .A(net677),
    .B(_2603_));
 sg13g2_xor2_1 _3544_ (.B(_2610_),
    .A(_2609_),
    .X(_2611_));
 sg13g2_xnor2_1 _3545_ (.Y(_2612_),
    .A(_2371_),
    .B(_2611_));
 sg13g2_inv_1 _3546_ (.Y(_2613_),
    .A(_2612_));
 sg13g2_xor2_1 _3547_ (.B(_2607_),
    .A(_2606_),
    .X(_2614_));
 sg13g2_a21oi_1 _3548_ (.A1(_2613_),
    .A2(_2614_),
    .Y(_2615_),
    .B1(_2608_));
 sg13g2_a21o_1 _3549_ (.A2(_2614_),
    .A1(_2613_),
    .B1(_2608_),
    .X(_2616_));
 sg13g2_o21ai_1 _3550_ (.B1(_2562_),
    .Y(_2617_),
    .A1(_2554_),
    .A2(_2556_));
 sg13g2_nand3_1 _3551_ (.B(_2616_),
    .C(_2617_),
    .A(_2563_),
    .Y(_2618_));
 sg13g2_a21oi_1 _3552_ (.A1(_2563_),
    .A2(_2617_),
    .Y(_2619_),
    .B1(_2616_));
 sg13g2_a21o_1 _3553_ (.A2(_2617_),
    .A1(_2563_),
    .B1(_2615_),
    .X(_2620_));
 sg13g2_nand3b_1 _3554_ (.B(_2617_),
    .C(_2563_),
    .Y(_2621_),
    .A_N(_2616_));
 sg13g2_xor2_1 _3555_ (.B(_2543_),
    .A(_2487_),
    .X(_2622_));
 sg13g2_nor2_1 _3556_ (.A(net708),
    .B(net706),
    .Y(_2623_));
 sg13g2_nor2_2 _3557_ (.A(net708),
    .B(_2485_),
    .Y(_2624_));
 sg13g2_xor2_1 _3558_ (.B(_2623_),
    .A(_2486_),
    .X(_2625_));
 sg13g2_xnor2_1 _3559_ (.Y(_2626_),
    .A(net709),
    .B(_2625_));
 sg13g2_nand2b_1 _3560_ (.Y(_2627_),
    .B(_2626_),
    .A_N(_2622_));
 sg13g2_nand3b_1 _3561_ (.B(_2602_),
    .C(net677),
    .Y(_2628_),
    .A_N(_2609_));
 sg13g2_o21ai_1 _3562_ (.B1(_2628_),
    .Y(_2629_),
    .A1(net678),
    .A2(_2611_));
 sg13g2_xor2_1 _3563_ (.B(_2571_),
    .A(_2570_),
    .X(_2630_));
 sg13g2_nand2_1 _3564_ (.Y(_2631_),
    .A(_2629_),
    .B(_2630_));
 sg13g2_xnor2_1 _3565_ (.Y(_2632_),
    .A(_2629_),
    .B(_2630_));
 sg13g2_xnor2_1 _3566_ (.Y(_2633_),
    .A(_2627_),
    .B(_2632_));
 sg13g2_a21oi_1 _3567_ (.A1(_2620_),
    .A2(_2621_),
    .Y(_2634_),
    .B1(_2633_));
 sg13g2_o21ai_1 _3568_ (.B1(_2618_),
    .Y(_2635_),
    .A1(_2619_),
    .A2(_2633_));
 sg13g2_xor2_1 _3569_ (.B(_2577_),
    .A(_2567_),
    .X(_2636_));
 sg13g2_nand2_1 _3570_ (.Y(_2637_),
    .A(_2635_),
    .B(_2636_));
 sg13g2_xnor2_1 _3571_ (.Y(_2638_),
    .A(_2635_),
    .B(_2636_));
 sg13g2_nor2_1 _3572_ (.A(net709),
    .B(net706),
    .Y(_2639_));
 sg13g2_o21ai_1 _3573_ (.B1(_2631_),
    .Y(_2640_),
    .A1(_2627_),
    .A2(_2632_));
 sg13g2_and2_1 _3574_ (.A(_2639_),
    .B(_2640_),
    .X(_2641_));
 sg13g2_xor2_1 _3575_ (.B(_2640_),
    .A(_2639_),
    .X(_2642_));
 sg13g2_xnor2_1 _3576_ (.Y(_2643_),
    .A(_2411_),
    .B(_2642_));
 sg13g2_o21ai_1 _3577_ (.B1(_2637_),
    .Y(_2644_),
    .A1(_2638_),
    .A2(_2643_));
 sg13g2_xor2_1 _3578_ (.B(_2586_),
    .A(_2581_),
    .X(_2645_));
 sg13g2_nand2_1 _3579_ (.Y(_2646_),
    .A(_2644_),
    .B(_2645_));
 sg13g2_a21o_1 _3580_ (.A2(_2642_),
    .A1(_2411_),
    .B1(_2641_),
    .X(_2647_));
 sg13g2_inv_1 _3581_ (.Y(_2648_),
    .A(_2647_));
 sg13g2_xnor2_1 _3582_ (.Y(_2649_),
    .A(_2644_),
    .B(_2645_));
 sg13g2_o21ai_1 _3583_ (.B1(_2646_),
    .Y(_2650_),
    .A1(_2648_),
    .A2(_2649_));
 sg13g2_xor2_1 _3584_ (.B(_2591_),
    .A(_2590_),
    .X(_2651_));
 sg13g2_nand2_1 _3585_ (.Y(_2652_),
    .A(_2650_),
    .B(_2651_));
 sg13g2_o21ai_1 _3586_ (.B1(_2539_),
    .Y(_2653_),
    .A1(_2589_),
    .A2(_2592_));
 sg13g2_and2_1 _3587_ (.A(_2652_),
    .B(_2653_),
    .X(_2654_));
 sg13g2_nand2_2 _3588_ (.Y(_2655_),
    .A(net719),
    .B(net711));
 sg13g2_nor2_2 _3589_ (.A(net709),
    .B(net708),
    .Y(_2656_));
 sg13g2_xnor2_1 _3590_ (.Y(_2657_),
    .A(_2596_),
    .B(_2656_));
 sg13g2_nor2_1 _3591_ (.A(_2540_),
    .B(_2657_),
    .Y(_2658_));
 sg13g2_xnor2_1 _3592_ (.Y(_2659_),
    .A(_2541_),
    .B(_2657_));
 sg13g2_nand2b_1 _3593_ (.Y(_2660_),
    .B(_2659_),
    .A_N(_2655_));
 sg13g2_nor2_1 _3594_ (.A(_0107_),
    .B(net706),
    .Y(_2661_));
 sg13g2_xor2_1 _3595_ (.B(_2661_),
    .A(_2597_),
    .X(_2662_));
 sg13g2_and2_1 _3596_ (.A(_2602_),
    .B(_2662_),
    .X(_2663_));
 sg13g2_xnor2_1 _3597_ (.Y(_2664_),
    .A(_2655_),
    .B(_2659_));
 sg13g2_nand2_1 _3598_ (.Y(_2665_),
    .A(_2663_),
    .B(_2664_));
 sg13g2_a21oi_1 _3599_ (.A1(_2596_),
    .A2(_2656_),
    .Y(_2666_),
    .B1(_2550_));
 sg13g2_a21oi_1 _3600_ (.A1(_2660_),
    .A2(_2665_),
    .Y(_2667_),
    .B1(_2666_));
 sg13g2_nand3_1 _3601_ (.B(_2665_),
    .C(_2666_),
    .A(_2660_),
    .Y(_2668_));
 sg13g2_nand2b_1 _3602_ (.Y(_2669_),
    .B(_2668_),
    .A_N(_2667_));
 sg13g2_nor3_1 _3603_ (.A(net708),
    .B(net706),
    .C(_2669_),
    .Y(_2670_));
 sg13g2_or2_1 _3604_ (.X(_2671_),
    .B(_2670_),
    .A(_2667_));
 sg13g2_and2_1 _3605_ (.A(_2598_),
    .B(_2624_),
    .X(_2672_));
 sg13g2_xnor2_1 _3606_ (.Y(_2673_),
    .A(_2547_),
    .B(_2597_));
 sg13g2_xnor2_1 _3607_ (.Y(_2674_),
    .A(_2672_),
    .B(_2673_));
 sg13g2_xnor2_1 _3608_ (.Y(_2675_),
    .A(_2602_),
    .B(_2674_));
 sg13g2_xnor2_1 _3609_ (.Y(_2676_),
    .A(_2598_),
    .B(_2624_));
 sg13g2_nand3_1 _3610_ (.B(_1961_),
    .C(_2395_),
    .A(net771),
    .Y(_2677_));
 sg13g2_or2_1 _3611_ (.X(_2678_),
    .B(_2677_),
    .A(_2676_));
 sg13g2_nor2_1 _3612_ (.A(_2675_),
    .B(_2678_),
    .Y(_2679_));
 sg13g2_nor2_1 _3613_ (.A(net719),
    .B(_2337_),
    .Y(_2680_));
 sg13g2_xor2_1 _3614_ (.B(_2678_),
    .A(_2675_),
    .X(_2681_));
 sg13g2_a21oi_1 _3615_ (.A1(_2680_),
    .A2(_2681_),
    .Y(_2682_),
    .B1(_2679_));
 sg13g2_nor2_2 _3616_ (.A(net718),
    .B(net713),
    .Y(_2683_));
 sg13g2_nor3_2 _3617_ (.A(net720),
    .B(_2495_),
    .C(_2683_),
    .Y(_2684_));
 sg13g2_a22oi_1 _3618_ (.Y(_2685_),
    .B1(_2674_),
    .B2(_2602_),
    .A2(_2672_),
    .A1(_2662_));
 sg13g2_xnor2_1 _3619_ (.Y(_2686_),
    .A(_2604_),
    .B(_2605_));
 sg13g2_nor2_1 _3620_ (.A(_2685_),
    .B(_2686_),
    .Y(_2687_));
 sg13g2_xor2_1 _3621_ (.B(_2686_),
    .A(_2685_),
    .X(_2688_));
 sg13g2_xnor2_1 _3622_ (.Y(_2689_),
    .A(_2684_),
    .B(_2688_));
 sg13g2_or2_1 _3623_ (.X(_2690_),
    .B(_2689_),
    .A(_2682_));
 sg13g2_xnor2_1 _3624_ (.Y(_2691_),
    .A(_2682_),
    .B(_2689_));
 sg13g2_xnor2_1 _3625_ (.Y(_2692_),
    .A(_2663_),
    .B(_2664_));
 sg13g2_o21ai_1 _3626_ (.B1(_2690_),
    .Y(_2693_),
    .A1(_2691_),
    .A2(_2692_));
 sg13g2_a21oi_2 _3627_ (.B1(_2687_),
    .Y(_2694_),
    .A2(_2688_),
    .A1(_2684_));
 sg13g2_xnor2_1 _3628_ (.Y(_2695_),
    .A(_2612_),
    .B(_2614_));
 sg13g2_nor2b_1 _3629_ (.A(_2694_),
    .B_N(_2695_),
    .Y(_2696_));
 sg13g2_xnor2_1 _3630_ (.Y(_2697_),
    .A(_2694_),
    .B(_2695_));
 sg13g2_nor2_2 _3631_ (.A(net720),
    .B(_2293_),
    .Y(_2698_));
 sg13g2_nor2_1 _3632_ (.A(_2091_),
    .B(_2494_),
    .Y(_2699_));
 sg13g2_xnor2_1 _3633_ (.Y(_2700_),
    .A(_2622_),
    .B(_2626_));
 sg13g2_nand2_1 _3634_ (.Y(_2701_),
    .A(_2699_),
    .B(_2700_));
 sg13g2_xor2_1 _3635_ (.B(_2700_),
    .A(_2699_),
    .X(_2702_));
 sg13g2_nand2_1 _3636_ (.Y(_2703_),
    .A(_2658_),
    .B(_2702_));
 sg13g2_xor2_1 _3637_ (.B(_2702_),
    .A(_2658_),
    .X(_2704_));
 sg13g2_xnor2_1 _3638_ (.Y(_2705_),
    .A(_2697_),
    .B(_2704_));
 sg13g2_nand2b_1 _3639_ (.Y(_2706_),
    .B(_2693_),
    .A_N(_2705_));
 sg13g2_xor2_1 _3640_ (.B(_2705_),
    .A(_2693_),
    .X(_2707_));
 sg13g2_xor2_1 _3641_ (.B(_2669_),
    .A(_2623_),
    .X(_2708_));
 sg13g2_o21ai_1 _3642_ (.B1(_2706_),
    .Y(_2709_),
    .A1(_2707_),
    .A2(_2708_));
 sg13g2_a21oi_2 _3643_ (.B1(_2696_),
    .Y(_2710_),
    .A2(_2704_),
    .A1(_2697_));
 sg13g2_and3_1 _3644_ (.X(_2711_),
    .A(_2620_),
    .B(_2621_),
    .C(_2633_));
 sg13g2_nor3_1 _3645_ (.A(_2634_),
    .B(_2710_),
    .C(_2711_),
    .Y(_2712_));
 sg13g2_or3_1 _3646_ (.A(_2634_),
    .B(_2710_),
    .C(_2711_),
    .X(_2713_));
 sg13g2_o21ai_1 _3647_ (.B1(_2710_),
    .Y(_2714_),
    .A1(_2634_),
    .A2(_2711_));
 sg13g2_a22oi_1 _3648_ (.Y(_2715_),
    .B1(_2625_),
    .B2(_2393_),
    .A2(_2624_),
    .A1(_2417_));
 sg13g2_a21oi_1 _3649_ (.A1(_2701_),
    .A2(_2703_),
    .Y(_2716_),
    .B1(_2715_));
 sg13g2_nand3_1 _3650_ (.B(_2703_),
    .C(_2715_),
    .A(_2701_),
    .Y(_2717_));
 sg13g2_nand2b_1 _3651_ (.Y(_2718_),
    .B(_2717_),
    .A_N(_2716_));
 sg13g2_nor2_1 _3652_ (.A(_2570_),
    .B(_2718_),
    .Y(_2719_));
 sg13g2_xor2_1 _3653_ (.B(_2718_),
    .A(_2570_),
    .X(_2720_));
 sg13g2_nand3_1 _3654_ (.B(_2714_),
    .C(_2720_),
    .A(_2713_),
    .Y(_2721_));
 sg13g2_a21o_1 _3655_ (.A2(_2714_),
    .A1(_2713_),
    .B1(_2720_),
    .X(_2722_));
 sg13g2_and3_1 _3656_ (.X(_2723_),
    .A(_2709_),
    .B(_2721_),
    .C(_2722_));
 sg13g2_nand3_1 _3657_ (.B(_2721_),
    .C(_2722_),
    .A(_2709_),
    .Y(_2724_));
 sg13g2_a21o_1 _3658_ (.A2(_2722_),
    .A1(_2721_),
    .B1(_2709_),
    .X(_2725_));
 sg13g2_nand3_1 _3659_ (.B(_2724_),
    .C(_2725_),
    .A(_2671_),
    .Y(_2726_));
 sg13g2_a21o_1 _3660_ (.A2(_2725_),
    .A1(_2724_),
    .B1(_2671_),
    .X(_2727_));
 sg13g2_xor2_1 _3661_ (.B(_2677_),
    .A(_2676_),
    .X(_2728_));
 sg13g2_nor2_1 _3662_ (.A(_0107_),
    .B(net708),
    .Y(_2729_));
 sg13g2_nand2_1 _3663_ (.Y(_2730_),
    .A(net822),
    .B(_2395_));
 sg13g2_xnor2_1 _3664_ (.Y(_2731_),
    .A(_1961_),
    .B(_2729_));
 sg13g2_nor3_2 _3665_ (.A(net820),
    .B(_2485_),
    .C(_2731_),
    .Y(_2732_));
 sg13g2_nand2_1 _3666_ (.Y(_2733_),
    .A(_2728_),
    .B(_2732_));
 sg13g2_nor2_1 _3667_ (.A(net720),
    .B(net678),
    .Y(_2734_));
 sg13g2_a221oi_1 _3668_ (.B2(net711),
    .C1(_0025_),
    .B1(_2698_),
    .A1(_2293_),
    .Y(_2735_),
    .A2(_2655_));
 sg13g2_inv_1 _3669_ (.Y(_2736_),
    .A(_2735_));
 sg13g2_xnor2_1 _3670_ (.Y(_2737_),
    .A(_2728_),
    .B(_2732_));
 sg13g2_o21ai_1 _3671_ (.B1(_2733_),
    .Y(_2738_),
    .A1(_2736_),
    .A2(_2737_));
 sg13g2_xor2_1 _3672_ (.B(_2681_),
    .A(_2680_),
    .X(_2739_));
 sg13g2_and2_1 _3673_ (.A(_2738_),
    .B(_2739_),
    .X(_2740_));
 sg13g2_or2_1 _3674_ (.X(_2741_),
    .B(_2739_),
    .A(_2738_));
 sg13g2_xnor2_1 _3675_ (.Y(_2742_),
    .A(_2738_),
    .B(_2739_));
 sg13g2_nand2_2 _3676_ (.Y(_2743_),
    .A(net862),
    .B(net713));
 sg13g2_nand2_1 _3677_ (.Y(_2744_),
    .A(net822),
    .B(_2393_));
 sg13g2_or2_1 _3678_ (.X(_2745_),
    .B(_2744_),
    .A(_2743_));
 sg13g2_nand2_2 _3679_ (.Y(_2746_),
    .A(_0063_),
    .B(net711));
 sg13g2_nor3_2 _3680_ (.A(_0025_),
    .B(net720),
    .C(net678),
    .Y(_2747_));
 sg13g2_xnor2_1 _3681_ (.Y(_2748_),
    .A(_2602_),
    .B(_2673_));
 sg13g2_xor2_1 _3682_ (.B(_2748_),
    .A(_2747_),
    .X(_2749_));
 sg13g2_nor2b_1 _3683_ (.A(_2745_),
    .B_N(_2749_),
    .Y(_2750_));
 sg13g2_xnor2_1 _3684_ (.Y(_2751_),
    .A(_2745_),
    .B(_2749_));
 sg13g2_a21oi_1 _3685_ (.A1(_2741_),
    .A2(_2751_),
    .Y(_2752_),
    .B1(_2740_));
 sg13g2_xnor2_1 _3686_ (.Y(_2753_),
    .A(_2691_),
    .B(_2692_));
 sg13g2_nor2_1 _3687_ (.A(_2752_),
    .B(_2753_),
    .Y(_2754_));
 sg13g2_xor2_1 _3688_ (.B(_2753_),
    .A(_2752_),
    .X(_2755_));
 sg13g2_a21oi_1 _3689_ (.A1(_2747_),
    .A2(_2748_),
    .Y(_2756_),
    .B1(_2750_));
 sg13g2_nand2b_1 _3690_ (.Y(_2757_),
    .B(_2599_),
    .A_N(_2756_));
 sg13g2_xnor2_1 _3691_ (.Y(_2758_),
    .A(_2599_),
    .B(_2756_));
 sg13g2_nand2_1 _3692_ (.Y(_2759_),
    .A(_2656_),
    .B(_2758_));
 sg13g2_xor2_1 _3693_ (.B(_2758_),
    .A(_2656_),
    .X(_2760_));
 sg13g2_a21o_1 _3694_ (.A2(_2760_),
    .A1(_2755_),
    .B1(_2754_),
    .X(_2761_));
 sg13g2_xor2_1 _3695_ (.B(_2708_),
    .A(_2707_),
    .X(_2762_));
 sg13g2_nand2_1 _3696_ (.Y(_2763_),
    .A(_2761_),
    .B(_2762_));
 sg13g2_and2_1 _3697_ (.A(_2757_),
    .B(_2759_),
    .X(_2764_));
 sg13g2_xnor2_1 _3698_ (.Y(_2765_),
    .A(_2761_),
    .B(_2762_));
 sg13g2_o21ai_1 _3699_ (.B1(_2763_),
    .Y(_2766_),
    .A1(_2764_),
    .A2(_2765_));
 sg13g2_nand3_1 _3700_ (.B(_2727_),
    .C(_2766_),
    .A(_2726_),
    .Y(_2767_));
 sg13g2_nor2_1 _3701_ (.A(net825),
    .B(_2485_),
    .Y(_2768_));
 sg13g2_inv_1 _3702_ (.Y(_2769_),
    .A(_2768_));
 sg13g2_xnor2_1 _3703_ (.Y(_2770_),
    .A(net720),
    .B(_2746_));
 sg13g2_a21oi_1 _3704_ (.A1(_2730_),
    .A2(_2769_),
    .Y(_2771_),
    .B1(_2770_));
 sg13g2_inv_1 _3705_ (.Y(_2772_),
    .A(_2771_));
 sg13g2_xnor2_1 _3706_ (.Y(_2773_),
    .A(_2736_),
    .B(_2737_));
 sg13g2_nor2_1 _3707_ (.A(_2772_),
    .B(_2773_),
    .Y(_2774_));
 sg13g2_xor2_1 _3708_ (.B(_2744_),
    .A(_2743_),
    .X(_2775_));
 sg13g2_xnor2_1 _3709_ (.Y(_2776_),
    .A(_2772_),
    .B(_2773_));
 sg13g2_inv_1 _3710_ (.Y(_2777_),
    .A(_2776_));
 sg13g2_a21oi_1 _3711_ (.A1(_2775_),
    .A2(_2777_),
    .Y(_2778_),
    .B1(_2774_));
 sg13g2_xnor2_1 _3712_ (.Y(_2779_),
    .A(_2742_),
    .B(_2751_));
 sg13g2_nand2b_1 _3713_ (.Y(_2780_),
    .B(_2779_),
    .A_N(_2778_));
 sg13g2_xor2_1 _3714_ (.B(_2779_),
    .A(_2778_),
    .X(_2781_));
 sg13g2_o21ai_1 _3715_ (.B1(_2780_),
    .Y(_2782_),
    .A1(net708),
    .A2(_2781_));
 sg13g2_xor2_1 _3716_ (.B(_2760_),
    .A(_2755_),
    .X(_2783_));
 sg13g2_nand2_1 _3717_ (.Y(_2784_),
    .A(_2782_),
    .B(_2783_));
 sg13g2_nor3_1 _3718_ (.A(net720),
    .B(_2729_),
    .C(_2768_),
    .Y(_2785_));
 sg13g2_nor3_1 _3719_ (.A(_2746_),
    .B(_2771_),
    .C(_2785_),
    .Y(_2786_));
 sg13g2_inv_1 _3720_ (.Y(_2787_),
    .A(_2786_));
 sg13g2_xor2_1 _3721_ (.B(_2776_),
    .A(_2775_),
    .X(_2788_));
 sg13g2_nor2_1 _3722_ (.A(_2787_),
    .B(_2788_),
    .Y(_2789_));
 sg13g2_nand2_1 _3723_ (.Y(_2790_),
    .A(_2787_),
    .B(_2788_));
 sg13g2_xnor2_1 _3724_ (.Y(_2791_),
    .A(_2786_),
    .B(_2788_));
 sg13g2_nor2_1 _3725_ (.A(_2729_),
    .B(_2785_),
    .Y(_2792_));
 sg13g2_nor2_2 _3726_ (.A(net862),
    .B(net720),
    .Y(_2793_));
 sg13g2_nor2_1 _3727_ (.A(_2792_),
    .B(_2793_),
    .Y(_2794_));
 sg13g2_o21ai_1 _3728_ (.B1(_2794_),
    .Y(_2795_),
    .A1(_2624_),
    .A2(_2791_));
 sg13g2_xnor2_1 _3729_ (.Y(_2796_),
    .A(_2395_),
    .B(_2781_));
 sg13g2_o21ai_1 _3730_ (.B1(_2790_),
    .Y(_2797_),
    .A1(_2624_),
    .A2(_2789_));
 sg13g2_nor2_1 _3731_ (.A(_2782_),
    .B(_2783_),
    .Y(_2798_));
 sg13g2_nor3_1 _3732_ (.A(_2787_),
    .B(_2788_),
    .C(_2795_),
    .Y(_2799_));
 sg13g2_nand2_1 _3733_ (.Y(_2800_),
    .A(_2795_),
    .B(_2797_));
 sg13g2_o21ai_1 _3734_ (.B1(_2800_),
    .Y(_2801_),
    .A1(_2796_),
    .A2(_2799_));
 sg13g2_a221oi_1 _3735_ (.B2(_2801_),
    .C1(_2798_),
    .B1(_2784_),
    .A1(_2764_),
    .Y(_2802_),
    .A2(_2765_));
 sg13g2_o21ai_1 _3736_ (.B1(_2802_),
    .Y(_2803_),
    .A1(_2764_),
    .A2(_2765_));
 sg13g2_nor2_1 _3737_ (.A(_2716_),
    .B(_2719_),
    .Y(_2804_));
 sg13g2_a21oi_1 _3738_ (.A1(_2714_),
    .A2(_2720_),
    .Y(_2805_),
    .B1(_2712_));
 sg13g2_xor2_1 _3739_ (.B(_2643_),
    .A(_2638_),
    .X(_2806_));
 sg13g2_nand2b_1 _3740_ (.Y(_2807_),
    .B(_2806_),
    .A_N(_2805_));
 sg13g2_xnor2_1 _3741_ (.Y(_2808_),
    .A(_2805_),
    .B(_2806_));
 sg13g2_nand2b_1 _3742_ (.Y(_2809_),
    .B(_2808_),
    .A_N(_2804_));
 sg13g2_xor2_1 _3743_ (.B(_2808_),
    .A(_2804_),
    .X(_2810_));
 sg13g2_a21oi_1 _3744_ (.A1(_2671_),
    .A2(_2725_),
    .Y(_2811_),
    .B1(_2723_));
 sg13g2_a21oi_1 _3745_ (.A1(_2726_),
    .A2(_2727_),
    .Y(_2812_),
    .B1(_2766_));
 sg13g2_a221oi_1 _3746_ (.B2(_2811_),
    .C1(_2812_),
    .B1(_2810_),
    .A1(_2767_),
    .Y(_2813_),
    .A2(_2803_));
 sg13g2_and2_1 _3747_ (.A(_2807_),
    .B(_2809_),
    .X(_2814_));
 sg13g2_xnor2_1 _3748_ (.Y(_2815_),
    .A(_2648_),
    .B(_2649_));
 sg13g2_or2_1 _3749_ (.X(_2816_),
    .B(_2811_),
    .A(_2810_));
 sg13g2_o21ai_1 _3750_ (.B1(_2816_),
    .Y(_2817_),
    .A1(_2814_),
    .A2(_2815_));
 sg13g2_nor2_1 _3751_ (.A(_2650_),
    .B(_2651_),
    .Y(_2818_));
 sg13g2_a21oi_1 _3752_ (.A1(_2814_),
    .A2(_2815_),
    .Y(_2819_),
    .B1(_2818_));
 sg13g2_o21ai_1 _3753_ (.B1(_2819_),
    .Y(_2820_),
    .A1(_2813_),
    .A2(_2817_));
 sg13g2_a21oi_1 _3754_ (.A1(_2654_),
    .A2(_2820_),
    .Y(_2821_),
    .B1(_2593_));
 sg13g2_a221oi_1 _3755_ (.B2(_2820_),
    .C1(_2593_),
    .B1(_2654_),
    .A1(_2536_),
    .Y(_2822_),
    .A2(_2537_));
 sg13g2_xnor2_1 _3756_ (.Y(_2823_),
    .A(_2467_),
    .B(_2483_));
 sg13g2_inv_1 _3757_ (.Y(_2824_),
    .A(_2823_));
 sg13g2_o21ai_1 _3758_ (.B1(_2824_),
    .Y(_2825_),
    .A1(_2535_),
    .A2(_2822_));
 sg13g2_a21oi_1 _3759_ (.A1(_2450_),
    .A2(_2481_),
    .Y(_2826_),
    .B1(_2480_));
 sg13g2_o21ai_1 _3760_ (.B1(_2478_),
    .Y(_2827_),
    .A1(_2470_),
    .A2(_2476_));
 sg13g2_o21ai_1 _3761_ (.B1(_2475_),
    .Y(_2828_),
    .A1(net679),
    .A2(_2370_));
 sg13g2_nor2_1 _3762_ (.A(_1895_),
    .B(net715),
    .Y(_2829_));
 sg13g2_o21ai_1 _3763_ (.B1(net725),
    .Y(_2830_),
    .A1(_2004_),
    .A2(_2417_));
 sg13g2_xnor2_1 _3764_ (.Y(_2831_),
    .A(_2829_),
    .B(_2830_));
 sg13g2_xnor2_1 _3765_ (.Y(_2832_),
    .A(_2828_),
    .B(_2831_));
 sg13g2_xnor2_1 _3766_ (.Y(_2833_),
    .A(_2827_),
    .B(_2832_));
 sg13g2_xnor2_1 _3767_ (.Y(_2834_),
    .A(_2826_),
    .B(_2833_));
 sg13g2_and3_2 _3768_ (.X(_2835_),
    .A(_2484_),
    .B(_2825_),
    .C(_2834_));
 sg13g2_a21oi_2 _3769_ (.B1(_2834_),
    .Y(_2836_),
    .A2(_2825_),
    .A1(_2484_));
 sg13g2_nor2_1 _3770_ (.A(_2835_),
    .B(_2836_),
    .Y(_2837_));
 sg13g2_xnor2_1 _3771_ (.Y(_2838_),
    .A(_2538_),
    .B(_2821_));
 sg13g2_o21ai_1 _3772_ (.B1(_2823_),
    .Y(_2839_),
    .A1(_2535_),
    .A2(_2822_));
 sg13g2_or3_1 _3773_ (.A(_2535_),
    .B(_2822_),
    .C(_2823_),
    .X(_2840_));
 sg13g2_nand3_1 _3774_ (.B(_2839_),
    .C(_2840_),
    .A(_2838_),
    .Y(_2841_));
 sg13g2_inv_1 _3775_ (.Y(_2842_),
    .A(_2841_));
 sg13g2_nor2_1 _3776_ (.A(net717),
    .B(net714),
    .Y(_2843_));
 sg13g2_a21oi_2 _3777_ (.B1(_1895_),
    .Y(_2844_),
    .A2(_2843_),
    .A1(net679));
 sg13g2_nand2_2 _3778_ (.Y(_2845_),
    .A(net707),
    .B(net705));
 sg13g2_o21ai_1 _3779_ (.B1(net725),
    .Y(_2846_),
    .A1(_1993_),
    .A2(_2845_));
 sg13g2_nor2b_2 _3780_ (.A(_2844_),
    .B_N(_2846_),
    .Y(_2847_));
 sg13g2_and4_1 _3781_ (.A(_2838_),
    .B(_2839_),
    .C(_2840_),
    .D(_2847_),
    .X(_2848_));
 sg13g2_o21ai_1 _3782_ (.B1(_2848_),
    .Y(_2849_),
    .A1(_2835_),
    .A2(_2836_));
 sg13g2_nor2_2 _3783_ (.A(_1665_),
    .B(net723),
    .Y(_2850_));
 sg13g2_a21oi_1 _3784_ (.A1(_2837_),
    .A2(_2850_),
    .Y(_2851_),
    .B1(_1325_));
 sg13g2_a21oi_1 _3785_ (.A1(_2849_),
    .A2(_2851_),
    .Y(_2852_),
    .B1(_1479_));
 sg13g2_o21ai_1 _3786_ (.B1(_1303_),
    .Y(_2853_),
    .A1(_1336_),
    .A2(_2852_));
 sg13g2_nand2_2 _3787_ (.Y(_2854_),
    .A(net815),
    .B(net819));
 sg13g2_and3_2 _3788_ (.X(_2855_),
    .A(net822),
    .B(net815),
    .C(net819));
 sg13g2_nor2_2 _3789_ (.A(net811),
    .B(_2855_),
    .Y(_2856_));
 sg13g2_o21ai_1 _3790_ (.B1(_1446_),
    .Y(_2857_),
    .A1(net811),
    .A2(_2855_));
 sg13g2_nor2b_2 _3791_ (.A(net810),
    .B_N(net814),
    .Y(_2858_));
 sg13g2_nand2_1 _3792_ (.Y(_2859_),
    .A(net814),
    .B(_0217_));
 sg13g2_nor2b_1 _3793_ (.A(net824),
    .B_N(net817),
    .Y(_2860_));
 sg13g2_nand2b_2 _3794_ (.Y(_2861_),
    .B(net819),
    .A_N(net822));
 sg13g2_nand4_1 _3795_ (.B(_1523_),
    .C(_2858_),
    .A(net767),
    .Y(_2862_),
    .D(_2860_));
 sg13g2_a21oi_1 _3796_ (.A1(net799),
    .A2(_0732_),
    .Y(_2863_),
    .B1(net794));
 sg13g2_nand4_1 _3797_ (.B(_2857_),
    .C(_2862_),
    .A(net763),
    .Y(_2864_),
    .D(_2863_));
 sg13g2_nor2_2 _3798_ (.A(net808),
    .B(net812),
    .Y(_2865_));
 sg13g2_nand2_2 _3799_ (.Y(_2866_),
    .A(_0206_),
    .B(_0217_));
 sg13g2_nand2_1 _3800_ (.Y(_2867_),
    .A(_2854_),
    .B(_2865_));
 sg13g2_xor2_1 _3801_ (.B(_2867_),
    .A(net801),
    .X(_2868_));
 sg13g2_nor3_1 _3802_ (.A(net811),
    .B(_0316_),
    .C(_2855_),
    .Y(_2869_));
 sg13g2_xnor2_1 _3803_ (.Y(_2870_),
    .A(net804),
    .B(_2869_));
 sg13g2_mux2_2 _3804_ (.A0(_2870_),
    .A1(_2868_),
    .S(_2864_),
    .X(_2871_));
 sg13g2_nor2_1 _3805_ (.A(net809),
    .B(_2854_),
    .Y(_2872_));
 sg13g2_nand2_1 _3806_ (.Y(_2873_),
    .A(net809),
    .B(_2854_));
 sg13g2_xnor2_1 _3807_ (.Y(_2874_),
    .A(net809),
    .B(_2854_));
 sg13g2_inv_1 _3808_ (.Y(_2875_),
    .A(_2874_));
 sg13g2_nor2_1 _3809_ (.A(net813),
    .B(_1928_),
    .Y(_2876_));
 sg13g2_xnor2_1 _3810_ (.Y(_2877_),
    .A(net811),
    .B(_2876_));
 sg13g2_nand2_1 _3811_ (.Y(_2878_),
    .A(_2864_),
    .B(_2874_));
 sg13g2_o21ai_1 _3812_ (.B1(_2878_),
    .Y(_2879_),
    .A1(_2864_),
    .A2(_2877_));
 sg13g2_nand2_1 _3813_ (.Y(_2880_),
    .A(_2871_),
    .B(_2879_));
 sg13g2_nand2_1 _3814_ (.Y(_2881_),
    .A(_2293_),
    .B(net680));
 sg13g2_nand3b_1 _3815_ (.B(_2881_),
    .C(net718),
    .Y(_2882_),
    .A_N(_2358_));
 sg13g2_nor2_1 _3816_ (.A(_2880_),
    .B(_2882_),
    .Y(_2883_));
 sg13g2_xor2_1 _3817_ (.B(_2882_),
    .A(_2880_),
    .X(_2884_));
 sg13g2_mux2_1 _3818_ (.A0(_2856_),
    .A1(_2873_),
    .S(_2864_),
    .X(_2885_));
 sg13g2_xnor2_1 _3819_ (.Y(_2886_),
    .A(net805),
    .B(_2885_));
 sg13g2_xnor2_1 _3820_ (.Y(_2887_),
    .A(_0316_),
    .B(_2885_));
 sg13g2_nor2_1 _3821_ (.A(_2879_),
    .B(_2886_),
    .Y(_2888_));
 sg13g2_a221oi_1 _3822_ (.B2(net711),
    .C1(_2683_),
    .B1(_2495_),
    .A1(net713),
    .Y(_2889_),
    .A2(net680));
 sg13g2_nand2_1 _3823_ (.Y(_2890_),
    .A(_2888_),
    .B(_2889_));
 sg13g2_nand2_1 _3824_ (.Y(_2891_),
    .A(_2498_),
    .B(_2890_));
 sg13g2_nand2_1 _3825_ (.Y(_2892_),
    .A(_2884_),
    .B(_2891_));
 sg13g2_and2_1 _3826_ (.A(_2879_),
    .B(_2887_),
    .X(_2893_));
 sg13g2_nand2b_1 _3827_ (.Y(_2894_),
    .B(_2893_),
    .A_N(_2385_));
 sg13g2_xnor2_1 _3828_ (.Y(_2895_),
    .A(_2385_),
    .B(_2893_));
 sg13g2_xor2_1 _3829_ (.B(_2891_),
    .A(_2884_),
    .X(_2896_));
 sg13g2_nand2_1 _3830_ (.Y(_2897_),
    .A(_2895_),
    .B(_2896_));
 sg13g2_nor2_2 _3831_ (.A(net680),
    .B(_2494_),
    .Y(_2898_));
 sg13g2_nand2_1 _3832_ (.Y(_2899_),
    .A(_2871_),
    .B(_2886_));
 sg13g2_xnor2_1 _3833_ (.Y(_2900_),
    .A(_2898_),
    .B(_2899_));
 sg13g2_nand2_1 _3834_ (.Y(_2901_),
    .A(_2883_),
    .B(_2900_));
 sg13g2_xnor2_1 _3835_ (.Y(_2902_),
    .A(_2883_),
    .B(_2900_));
 sg13g2_xnor2_1 _3836_ (.Y(_2903_),
    .A(net680),
    .B(_2902_));
 sg13g2_a21o_1 _3837_ (.A2(_2897_),
    .A1(_2892_),
    .B1(_2903_),
    .X(_2904_));
 sg13g2_nand3_1 _3838_ (.B(_2897_),
    .C(_2903_),
    .A(_2892_),
    .Y(_2905_));
 sg13g2_nand2_1 _3839_ (.Y(_2906_),
    .A(_2904_),
    .B(_2905_));
 sg13g2_o21ai_1 _3840_ (.B1(_2904_),
    .Y(_2907_),
    .A1(_2894_),
    .A2(_2906_));
 sg13g2_o21ai_1 _3841_ (.B1(_2901_),
    .Y(_2908_),
    .A1(net680),
    .A2(_2902_));
 sg13g2_o21ai_1 _3842_ (.B1(_2871_),
    .Y(_2909_),
    .A1(_2887_),
    .A2(_2898_));
 sg13g2_xnor2_1 _3843_ (.Y(_2910_),
    .A(_2908_),
    .B(_2909_));
 sg13g2_xnor2_1 _3844_ (.Y(_2911_),
    .A(_2907_),
    .B(_2910_));
 sg13g2_o21ai_1 _3845_ (.B1(_2498_),
    .Y(_2912_),
    .A1(_2356_),
    .A2(_2497_));
 sg13g2_nand2_2 _3846_ (.Y(_2913_),
    .A(net823),
    .B(_2871_));
 sg13g2_or2_1 _3847_ (.X(_2914_),
    .B(_2913_),
    .A(_2601_));
 sg13g2_xnor2_1 _3848_ (.Y(_2915_),
    .A(_2601_),
    .B(_2913_));
 sg13g2_o21ai_1 _3849_ (.B1(_2914_),
    .Y(_2916_),
    .A1(net678),
    .A2(_2915_));
 sg13g2_nand2_1 _3850_ (.Y(_2917_),
    .A(_2609_),
    .B(_2916_));
 sg13g2_nand2b_1 _3851_ (.Y(_2918_),
    .B(net677),
    .A_N(_2496_));
 sg13g2_xor2_1 _3852_ (.B(net677),
    .A(_2496_),
    .X(_2919_));
 sg13g2_xnor2_1 _3853_ (.Y(_2920_),
    .A(_2609_),
    .B(_2916_));
 sg13g2_o21ai_1 _3854_ (.B1(_2917_),
    .Y(_2921_),
    .A1(_2919_),
    .A2(_2920_));
 sg13g2_nand2b_1 _3855_ (.Y(_2922_),
    .B(_2921_),
    .A_N(_2912_));
 sg13g2_xor2_1 _3856_ (.B(_2921_),
    .A(_2912_),
    .X(_2923_));
 sg13g2_nand2_1 _3857_ (.Y(_2924_),
    .A(net822),
    .B(_0184_));
 sg13g2_xnor2_1 _3858_ (.Y(_2925_),
    .A(_0184_),
    .B(_1928_));
 sg13g2_inv_1 _3859_ (.Y(_2926_),
    .A(_2925_));
 sg13g2_nor2b_1 _3860_ (.A(_1369_),
    .B_N(_2854_),
    .Y(_2927_));
 sg13g2_nand2b_1 _3861_ (.Y(_2928_),
    .B(_2854_),
    .A_N(_1369_));
 sg13g2_nor2_1 _3862_ (.A(_2864_),
    .B(_2925_),
    .Y(_2929_));
 sg13g2_a21oi_2 _3863_ (.B1(_2929_),
    .Y(_2930_),
    .A2(_2928_),
    .A1(_2864_));
 sg13g2_nand2_2 _3864_ (.Y(_2931_),
    .A(_2871_),
    .B(_2930_));
 sg13g2_nor3_2 _3865_ (.A(_2337_),
    .B(net680),
    .C(_2931_),
    .Y(_2932_));
 sg13g2_or2_1 _3866_ (.X(_2933_),
    .B(_2931_),
    .A(_2918_));
 sg13g2_xnor2_1 _3867_ (.Y(_2934_),
    .A(_2918_),
    .B(_2931_));
 sg13g2_mux2_2 _3868_ (.A0(_1939_),
    .A1(net819),
    .S(_2864_),
    .X(_2935_));
 sg13g2_inv_1 _3869_ (.Y(_2936_),
    .A(_2935_));
 sg13g2_nand2_2 _3870_ (.Y(_2937_),
    .A(_2887_),
    .B(_2936_));
 sg13g2_nand2_1 _3871_ (.Y(_2938_),
    .A(_2887_),
    .B(_2930_));
 sg13g2_nand2_1 _3872_ (.Y(_2939_),
    .A(_2871_),
    .B(_2936_));
 sg13g2_nor2_1 _3873_ (.A(_2931_),
    .B(_2937_),
    .Y(_2940_));
 sg13g2_xor2_1 _3874_ (.B(_2939_),
    .A(_2938_),
    .X(_2941_));
 sg13g2_a21oi_1 _3875_ (.A1(net676),
    .A2(_2941_),
    .Y(_2942_),
    .B1(_2940_));
 sg13g2_xnor2_1 _3876_ (.Y(_2943_),
    .A(_2934_),
    .B(_2942_));
 sg13g2_o21ai_1 _3877_ (.B1(_2922_),
    .Y(_2944_),
    .A1(_2923_),
    .A2(_2943_));
 sg13g2_xnor2_1 _3878_ (.Y(_2945_),
    .A(_2888_),
    .B(_2889_));
 sg13g2_nand2b_1 _3879_ (.Y(_2946_),
    .B(_2944_),
    .A_N(_2945_));
 sg13g2_o21ai_1 _3880_ (.B1(_2933_),
    .Y(_2947_),
    .A1(_2934_),
    .A2(_2942_));
 sg13g2_and2_1 _3881_ (.A(_2358_),
    .B(_2947_),
    .X(_2948_));
 sg13g2_xor2_1 _3882_ (.B(_2947_),
    .A(_2358_),
    .X(_2949_));
 sg13g2_xnor2_1 _3883_ (.Y(_2950_),
    .A(_2932_),
    .B(_2949_));
 sg13g2_xor2_1 _3884_ (.B(_2945_),
    .A(_2944_),
    .X(_2951_));
 sg13g2_o21ai_1 _3885_ (.B1(_2946_),
    .Y(_2952_),
    .A1(_2950_),
    .A2(_2951_));
 sg13g2_inv_1 _3886_ (.Y(_2953_),
    .A(_2952_));
 sg13g2_xnor2_1 _3887_ (.Y(_2954_),
    .A(_2895_),
    .B(_2896_));
 sg13g2_a21o_1 _3888_ (.A2(_2949_),
    .A1(_2932_),
    .B1(_2948_),
    .X(_2955_));
 sg13g2_xor2_1 _3889_ (.B(_2954_),
    .A(_2952_),
    .X(_2956_));
 sg13g2_nand2b_1 _3890_ (.Y(_2957_),
    .B(_2955_),
    .A_N(_2956_));
 sg13g2_o21ai_1 _3891_ (.B1(_2957_),
    .Y(_2958_),
    .A1(_2953_),
    .A2(_2954_));
 sg13g2_xnor2_1 _3892_ (.Y(_2959_),
    .A(_2894_),
    .B(_2906_));
 sg13g2_nand2b_1 _3893_ (.Y(_2960_),
    .B(_2958_),
    .A_N(_2959_));
 sg13g2_xnor2_1 _3894_ (.Y(_2961_),
    .A(_2958_),
    .B(_2959_));
 sg13g2_nor2_1 _3895_ (.A(net820),
    .B(_2886_),
    .Y(_2962_));
 sg13g2_nor3_1 _3896_ (.A(net820),
    .B(_2603_),
    .C(_2886_),
    .Y(_2963_));
 sg13g2_nand3_1 _3897_ (.B(_2602_),
    .C(_2887_),
    .A(net771),
    .Y(_2964_));
 sg13g2_o21ai_1 _3898_ (.B1(_2603_),
    .Y(_2965_),
    .A1(net820),
    .A2(_2886_));
 sg13g2_nand3_1 _3899_ (.B(_2964_),
    .C(_2965_),
    .A(_2698_),
    .Y(_2966_));
 sg13g2_a21oi_2 _3900_ (.B1(_2963_),
    .Y(_2967_),
    .A2(_2965_),
    .A1(_2698_));
 sg13g2_xnor2_1 _3901_ (.Y(_2968_),
    .A(net678),
    .B(_2915_));
 sg13g2_nor2_1 _3902_ (.A(_2967_),
    .B(_2968_),
    .Y(_2969_));
 sg13g2_nor2_1 _3903_ (.A(net678),
    .B(_2601_),
    .Y(_2970_));
 sg13g2_xor2_1 _3904_ (.B(_2601_),
    .A(net678),
    .X(_2971_));
 sg13g2_xnor2_1 _3905_ (.Y(_2972_),
    .A(_2540_),
    .B(_2971_));
 sg13g2_xor2_1 _3906_ (.B(_2968_),
    .A(_2967_),
    .X(_2973_));
 sg13g2_a21oi_1 _3907_ (.A1(_2972_),
    .A2(_2973_),
    .Y(_2974_),
    .B1(_2969_));
 sg13g2_xnor2_1 _3908_ (.Y(_2975_),
    .A(_2919_),
    .B(_2920_));
 sg13g2_nor2_1 _3909_ (.A(_2974_),
    .B(_2975_),
    .Y(_2976_));
 sg13g2_nor2_1 _3910_ (.A(_2913_),
    .B(_2937_),
    .Y(_2977_));
 sg13g2_nand2_1 _3911_ (.Y(_2978_),
    .A(net676),
    .B(_2930_));
 sg13g2_inv_1 _3912_ (.Y(_2979_),
    .A(_2978_));
 sg13g2_xor2_1 _3913_ (.B(_2937_),
    .A(_2913_),
    .X(_2980_));
 sg13g2_a21oi_1 _3914_ (.A1(_2979_),
    .A2(_2980_),
    .Y(_2981_),
    .B1(_2977_));
 sg13g2_a21oi_1 _3915_ (.A1(_2541_),
    .A2(_2971_),
    .Y(_2982_),
    .B1(_2970_));
 sg13g2_xor2_1 _3916_ (.B(_2941_),
    .A(net676),
    .X(_2983_));
 sg13g2_nand2b_1 _3917_ (.Y(_2984_),
    .B(_2983_),
    .A_N(_2982_));
 sg13g2_xor2_1 _3918_ (.B(_2983_),
    .A(_2982_),
    .X(_2985_));
 sg13g2_xor2_1 _3919_ (.B(_2985_),
    .A(_2981_),
    .X(_2986_));
 sg13g2_xor2_1 _3920_ (.B(_2975_),
    .A(_2974_),
    .X(_2987_));
 sg13g2_a21oi_1 _3921_ (.A1(_2986_),
    .A2(_2987_),
    .Y(_2988_),
    .B1(_2976_));
 sg13g2_xor2_1 _3922_ (.B(_2943_),
    .A(_2923_),
    .X(_2989_));
 sg13g2_nor2b_1 _3923_ (.A(_2988_),
    .B_N(_2989_),
    .Y(_2990_));
 sg13g2_o21ai_1 _3924_ (.B1(_2984_),
    .Y(_2991_),
    .A1(_2981_),
    .A2(_2985_));
 sg13g2_xor2_1 _3925_ (.B(_2931_),
    .A(_2356_),
    .X(_2992_));
 sg13g2_nand2b_1 _3926_ (.Y(_2993_),
    .B(_2991_),
    .A_N(_2992_));
 sg13g2_xor2_1 _3927_ (.B(_2992_),
    .A(_2991_),
    .X(_2994_));
 sg13g2_a21oi_2 _3928_ (.B1(_2940_),
    .Y(_2995_),
    .A2(_2941_),
    .A1(net677));
 sg13g2_xor2_1 _3929_ (.B(_2995_),
    .A(_2994_),
    .X(_2996_));
 sg13g2_xnor2_1 _3930_ (.Y(_2997_),
    .A(_2988_),
    .B(_2989_));
 sg13g2_a21oi_1 _3931_ (.A1(_2996_),
    .A2(_2997_),
    .Y(_2998_),
    .B1(_2990_));
 sg13g2_xor2_1 _3932_ (.B(_2951_),
    .A(_2950_),
    .X(_2999_));
 sg13g2_nor2b_1 _3933_ (.A(_2998_),
    .B_N(_2999_),
    .Y(_3000_));
 sg13g2_o21ai_1 _3934_ (.B1(_2993_),
    .Y(_3001_),
    .A1(_2994_),
    .A2(_2995_));
 sg13g2_xnor2_1 _3935_ (.Y(_3002_),
    .A(_2998_),
    .B(_2999_));
 sg13g2_a21oi_1 _3936_ (.A1(_3001_),
    .A2(_3002_),
    .Y(_3003_),
    .B1(_3000_));
 sg13g2_inv_1 _3937_ (.Y(_3004_),
    .A(_3003_));
 sg13g2_xor2_1 _3938_ (.B(_2956_),
    .A(_2955_),
    .X(_3005_));
 sg13g2_inv_1 _3939_ (.Y(_3006_),
    .A(_3005_));
 sg13g2_nand2_1 _3940_ (.Y(_3007_),
    .A(_3003_),
    .B(_3005_));
 sg13g2_nand2_1 _3941_ (.Y(_3008_),
    .A(_3004_),
    .B(_3006_));
 sg13g2_xnor2_1 _3942_ (.Y(_3009_),
    .A(_3001_),
    .B(_3002_));
 sg13g2_nand2_2 _3943_ (.Y(_3010_),
    .A(net823),
    .B(net676));
 sg13g2_nor2_1 _3944_ (.A(_2743_),
    .B(_3010_),
    .Y(_3011_));
 sg13g2_a21o_1 _3945_ (.A2(_2965_),
    .A1(_2964_),
    .B1(_2698_),
    .X(_3012_));
 sg13g2_and3_1 _3946_ (.X(_3013_),
    .A(_2966_),
    .B(_3011_),
    .C(_3012_));
 sg13g2_nand3_1 _3947_ (.B(_3011_),
    .C(_3012_),
    .A(_2966_),
    .Y(_3014_));
 sg13g2_a21o_1 _3948_ (.A2(_3012_),
    .A1(_2966_),
    .B1(_3011_),
    .X(_3015_));
 sg13g2_xnor2_1 _3949_ (.Y(_3016_),
    .A(_2337_),
    .B(_2698_));
 sg13g2_xnor2_1 _3950_ (.Y(_3017_),
    .A(_2603_),
    .B(_3016_));
 sg13g2_nand3_1 _3951_ (.B(_3015_),
    .C(_3017_),
    .A(_3014_),
    .Y(_3018_));
 sg13g2_a21oi_2 _3952_ (.B1(_3013_),
    .Y(_3019_),
    .A2(_3017_),
    .A1(_3015_));
 sg13g2_xnor2_1 _3953_ (.Y(_3020_),
    .A(_2972_),
    .B(_2973_));
 sg13g2_nor2_1 _3954_ (.A(_3019_),
    .B(_3020_),
    .Y(_3021_));
 sg13g2_and2_1 _3955_ (.A(net676),
    .B(_2936_),
    .X(_3022_));
 sg13g2_and2_1 _3956_ (.A(_2962_),
    .B(_3022_),
    .X(_3023_));
 sg13g2_a21oi_2 _3957_ (.B1(_2734_),
    .Y(_3024_),
    .A2(_3016_),
    .A1(_2602_));
 sg13g2_xnor2_1 _3958_ (.Y(_3025_),
    .A(_2979_),
    .B(_2980_));
 sg13g2_nor2_1 _3959_ (.A(_3024_),
    .B(_3025_),
    .Y(_3026_));
 sg13g2_xor2_1 _3960_ (.B(_3025_),
    .A(_3024_),
    .X(_3027_));
 sg13g2_xor2_1 _3961_ (.B(_3027_),
    .A(_3023_),
    .X(_3028_));
 sg13g2_xor2_1 _3962_ (.B(_3020_),
    .A(_3019_),
    .X(_3029_));
 sg13g2_a21oi_1 _3963_ (.A1(_3028_),
    .A2(_3029_),
    .Y(_3030_),
    .B1(_3021_));
 sg13g2_xnor2_1 _3964_ (.Y(_3031_),
    .A(_2986_),
    .B(_2987_));
 sg13g2_nor2_1 _3965_ (.A(_3030_),
    .B(_3031_),
    .Y(_3032_));
 sg13g2_and2_2 _3966_ (.A(_2930_),
    .B(_2936_),
    .X(_3033_));
 sg13g2_nand2_1 _3967_ (.Y(_3034_),
    .A(net676),
    .B(_3033_));
 sg13g2_inv_1 _3968_ (.Y(_3035_),
    .A(_3034_));
 sg13g2_nor2_1 _3969_ (.A(_2886_),
    .B(_3034_),
    .Y(_3036_));
 sg13g2_a21oi_1 _3970_ (.A1(_2937_),
    .A2(_2978_),
    .Y(_3037_),
    .B1(_3036_));
 sg13g2_a21oi_2 _3971_ (.B1(_3036_),
    .Y(_3038_),
    .A2(_3037_),
    .A1(_2541_));
 sg13g2_inv_1 _3972_ (.Y(_0053_),
    .A(_3038_));
 sg13g2_a21oi_2 _3973_ (.B1(_3026_),
    .Y(_0054_),
    .A2(_3027_),
    .A1(_3023_));
 sg13g2_xnor2_1 _3974_ (.Y(_0055_),
    .A(net677),
    .B(_2941_));
 sg13g2_nor2_1 _3975_ (.A(_0054_),
    .B(_0055_),
    .Y(_0056_));
 sg13g2_xor2_1 _3976_ (.B(_0055_),
    .A(_0054_),
    .X(_0057_));
 sg13g2_xnor2_1 _3977_ (.Y(_0058_),
    .A(_3038_),
    .B(_0057_));
 sg13g2_xor2_1 _3978_ (.B(_3031_),
    .A(_3030_),
    .X(_0059_));
 sg13g2_a21oi_1 _3979_ (.A1(_0058_),
    .A2(_0059_),
    .Y(_0060_),
    .B1(_3032_));
 sg13g2_xor2_1 _3980_ (.B(_2997_),
    .A(_2996_),
    .X(_0061_));
 sg13g2_nand2b_1 _3981_ (.Y(_0062_),
    .B(_0061_),
    .A_N(_0060_));
 sg13g2_a21oi_1 _3982_ (.A1(_0053_),
    .A2(_0057_),
    .Y(_0064_),
    .B1(_0056_));
 sg13g2_xnor2_1 _3983_ (.Y(_0065_),
    .A(_0060_),
    .B(_0061_));
 sg13g2_inv_1 _3984_ (.Y(_0066_),
    .A(_0065_));
 sg13g2_o21ai_1 _3985_ (.B1(_0062_),
    .Y(_0067_),
    .A1(_0064_),
    .A2(_0066_));
 sg13g2_nor2b_1 _3986_ (.A(_3009_),
    .B_N(_0067_),
    .Y(_0068_));
 sg13g2_xnor2_1 _3987_ (.Y(_0069_),
    .A(_0064_),
    .B(_0065_));
 sg13g2_a21oi_1 _3988_ (.A1(net823),
    .A2(net676),
    .Y(_0070_),
    .B1(_2743_));
 sg13g2_a21o_1 _3989_ (.A2(_3015_),
    .A1(_3014_),
    .B1(_3017_),
    .X(_0071_));
 sg13g2_and3_1 _3990_ (.X(_0072_),
    .A(_3018_),
    .B(_0070_),
    .C(_0071_));
 sg13g2_nand3_1 _3991_ (.B(_0070_),
    .C(_0071_),
    .A(_3018_),
    .Y(_0073_));
 sg13g2_xnor2_1 _3992_ (.Y(_0075_),
    .A(_2962_),
    .B(_3022_));
 sg13g2_nor2_1 _3993_ (.A(_2655_),
    .B(_0075_),
    .Y(_0076_));
 sg13g2_xnor2_1 _3994_ (.Y(_0077_),
    .A(_2655_),
    .B(_0075_));
 sg13g2_a21oi_1 _3995_ (.A1(_3018_),
    .A2(_0071_),
    .Y(_0078_),
    .B1(_0070_));
 sg13g2_or3_1 _3996_ (.A(_0072_),
    .B(_0077_),
    .C(_0078_),
    .X(_0079_));
 sg13g2_o21ai_1 _3997_ (.B1(_0073_),
    .Y(_0080_),
    .A1(_0077_),
    .A2(_0078_));
 sg13g2_xor2_1 _3998_ (.B(_3029_),
    .A(_3028_),
    .X(_0081_));
 sg13g2_nand2_1 _3999_ (.Y(_0082_),
    .A(_0080_),
    .B(_0081_));
 sg13g2_xnor2_1 _4000_ (.Y(_0083_),
    .A(_2540_),
    .B(_3037_));
 sg13g2_xor2_1 _4001_ (.B(_0083_),
    .A(_0076_),
    .X(_0084_));
 sg13g2_xnor2_1 _4002_ (.Y(_0086_),
    .A(_3035_),
    .B(_0084_));
 sg13g2_xnor2_1 _4003_ (.Y(_0087_),
    .A(_0080_),
    .B(_0081_));
 sg13g2_o21ai_1 _4004_ (.B1(_0082_),
    .Y(_0088_),
    .A1(_0086_),
    .A2(_0087_));
 sg13g2_xnor2_1 _4005_ (.Y(_0089_),
    .A(_0058_),
    .B(_0059_));
 sg13g2_nand2b_1 _4006_ (.Y(_0090_),
    .B(_0088_),
    .A_N(_0089_));
 sg13g2_a22oi_1 _4007_ (.Y(_0091_),
    .B1(_0084_),
    .B2(_3035_),
    .A2(_0083_),
    .A1(_0076_));
 sg13g2_xor2_1 _4008_ (.B(_0089_),
    .A(_0088_),
    .X(_0092_));
 sg13g2_o21ai_1 _4009_ (.B1(_0090_),
    .Y(_0093_),
    .A1(_0091_),
    .A2(_0092_));
 sg13g2_and2_1 _4010_ (.A(_0069_),
    .B(_0093_),
    .X(_0094_));
 sg13g2_or2_1 _4011_ (.X(_0095_),
    .B(_0093_),
    .A(_0069_));
 sg13g2_xnor2_1 _4012_ (.Y(_0097_),
    .A(_0069_),
    .B(_0093_));
 sg13g2_xnor2_1 _4013_ (.Y(_0098_),
    .A(_0091_),
    .B(_0092_));
 sg13g2_nand2_1 _4014_ (.Y(_0099_),
    .A(net823),
    .B(_2930_));
 sg13g2_nand4_1 _4015_ (.B(net719),
    .C(net676),
    .A(net822),
    .Y(_0100_),
    .D(_2930_));
 sg13g2_o21ai_1 _4016_ (.B1(_3010_),
    .Y(_0101_),
    .A1(net720),
    .A2(_0099_));
 sg13g2_nand2_1 _4017_ (.Y(_0102_),
    .A(_0100_),
    .B(_0101_));
 sg13g2_or2_1 _4018_ (.X(_0103_),
    .B(_3010_),
    .A(_2746_));
 sg13g2_xor2_1 _4019_ (.B(_3010_),
    .A(_2746_),
    .X(_0104_));
 sg13g2_nand3_1 _4020_ (.B(_0101_),
    .C(_0104_),
    .A(_0100_),
    .Y(_0105_));
 sg13g2_nand2_1 _4021_ (.Y(_0106_),
    .A(_0100_),
    .B(_0105_));
 sg13g2_o21ai_1 _4022_ (.B1(_0077_),
    .Y(_0108_),
    .A1(_0072_),
    .A2(_0078_));
 sg13g2_and3_1 _4023_ (.X(_0109_),
    .A(_0079_),
    .B(_0106_),
    .C(_0108_));
 sg13g2_nand3_1 _4024_ (.B(_0106_),
    .C(_0108_),
    .A(_0079_),
    .Y(_0110_));
 sg13g2_xnor2_1 _4025_ (.Y(_0111_),
    .A(_2930_),
    .B(_3022_));
 sg13g2_xor2_1 _4026_ (.B(_0111_),
    .A(_0103_),
    .X(_0112_));
 sg13g2_nand2_1 _4027_ (.Y(_0113_),
    .A(_3033_),
    .B(_0112_));
 sg13g2_xnor2_1 _4028_ (.Y(_0114_),
    .A(_3033_),
    .B(_0112_));
 sg13g2_a21oi_1 _4029_ (.A1(_0079_),
    .A2(_0108_),
    .Y(_0115_),
    .B1(_0106_));
 sg13g2_or3_1 _4030_ (.A(_0109_),
    .B(_0114_),
    .C(_0115_),
    .X(_0116_));
 sg13g2_o21ai_1 _4031_ (.B1(_0110_),
    .Y(_0117_),
    .A1(_0114_),
    .A2(_0115_));
 sg13g2_xor2_1 _4032_ (.B(_0087_),
    .A(_0086_),
    .X(_0119_));
 sg13g2_and2_1 _4033_ (.A(_0117_),
    .B(_0119_),
    .X(_0120_));
 sg13g2_o21ai_1 _4034_ (.B1(_0113_),
    .Y(_0121_),
    .A1(_0103_),
    .A2(_0111_));
 sg13g2_xor2_1 _4035_ (.B(_0119_),
    .A(_0117_),
    .X(_0122_));
 sg13g2_a21oi_1 _4036_ (.A1(_0121_),
    .A2(_0122_),
    .Y(_0123_),
    .B1(_0120_));
 sg13g2_o21ai_1 _4037_ (.B1(_0114_),
    .Y(_0124_),
    .A1(_0109_),
    .A2(_0115_));
 sg13g2_nand2_2 _4038_ (.Y(_0125_),
    .A(net866),
    .B(net824));
 sg13g2_xor2_1 _4039_ (.B(_0099_),
    .A(_2793_),
    .X(_0126_));
 sg13g2_o21ai_1 _4040_ (.B1(_0126_),
    .Y(_0127_),
    .A1(_2935_),
    .A2(_0125_));
 sg13g2_nand3_1 _4041_ (.B(net815),
    .C(_2935_),
    .A(net822),
    .Y(_0128_));
 sg13g2_nand3_1 _4042_ (.B(_0127_),
    .C(_0128_),
    .A(_2861_),
    .Y(_0130_));
 sg13g2_o21ai_1 _4043_ (.B1(_0130_),
    .Y(_0131_),
    .A1(_2924_),
    .A2(_2935_));
 sg13g2_xnor2_1 _4044_ (.Y(_0132_),
    .A(_0102_),
    .B(_0104_));
 sg13g2_or2_1 _4045_ (.X(_0133_),
    .B(_0132_),
    .A(_0131_));
 sg13g2_nand3_1 _4046_ (.B(net719),
    .C(_0099_),
    .A(net862),
    .Y(_0134_));
 sg13g2_a22oi_1 _4047_ (.Y(_0135_),
    .B1(_0131_),
    .B2(_0132_),
    .A2(_3033_),
    .A1(net822));
 sg13g2_nand2_1 _4048_ (.Y(_0136_),
    .A(_0134_),
    .B(_0135_));
 sg13g2_and4_1 _4049_ (.A(_0116_),
    .B(_0124_),
    .C(_0133_),
    .D(_0136_),
    .X(_0137_));
 sg13g2_o21ai_1 _4050_ (.B1(_0137_),
    .Y(_0138_),
    .A1(_0121_),
    .A2(_0122_));
 sg13g2_a21oi_1 _4051_ (.A1(_0123_),
    .A2(_0138_),
    .Y(_0139_),
    .B1(_0098_));
 sg13g2_a21o_1 _4052_ (.A2(_0139_),
    .A1(_0095_),
    .B1(_0094_),
    .X(_0141_));
 sg13g2_xnor2_1 _4053_ (.Y(_0142_),
    .A(_3009_),
    .B(_0067_));
 sg13g2_a221oi_1 _4054_ (.B2(_0142_),
    .C1(_0068_),
    .B1(_0141_),
    .A1(_3004_),
    .Y(_0143_),
    .A2(_3006_));
 sg13g2_a21o_1 _4055_ (.A2(_3005_),
    .A1(_3003_),
    .B1(_0143_),
    .X(_0144_));
 sg13g2_nand3b_1 _4056_ (.B(_2961_),
    .C(_3007_),
    .Y(_0145_),
    .A_N(_0143_));
 sg13g2_a21o_1 _4057_ (.A2(_0145_),
    .A1(_2960_),
    .B1(_2911_),
    .X(_0146_));
 sg13g2_nand3_1 _4058_ (.B(_2960_),
    .C(_0145_),
    .A(_2911_),
    .Y(_0147_));
 sg13g2_a221oi_1 _4059_ (.B2(_0142_),
    .C1(_0068_),
    .B1(_0141_),
    .A1(_3007_),
    .Y(_0148_),
    .A2(_3008_));
 sg13g2_xor2_1 _4060_ (.B(_0139_),
    .A(_0097_),
    .X(_0149_));
 sg13g2_a21oi_1 _4061_ (.A1(_0141_),
    .A2(_0142_),
    .Y(_0150_),
    .B1(_0149_));
 sg13g2_o21ai_1 _4062_ (.B1(_0150_),
    .Y(_0152_),
    .A1(_0094_),
    .A2(_0142_));
 sg13g2_nor2_2 _4063_ (.A(net842),
    .B(net847),
    .Y(_0153_));
 sg13g2_nor2_2 _4064_ (.A(_0579_),
    .B(_0153_),
    .Y(_0154_));
 sg13g2_mux2_1 _4065_ (.A0(_0012_),
    .A1(_0154_),
    .S(net743),
    .X(_0155_));
 sg13g2_nand2_1 _4066_ (.Y(_0156_),
    .A(net852),
    .B(net744));
 sg13g2_xnor2_1 _4067_ (.Y(_0157_),
    .A(net855),
    .B(net743));
 sg13g2_xnor2_1 _4068_ (.Y(_0158_),
    .A(net855),
    .B(net747));
 sg13g2_a21oi_2 _4069_ (.B1(_2179_),
    .Y(_0159_),
    .A2(net832),
    .A1(_0151_));
 sg13g2_o21ai_1 _4070_ (.B1(_2189_),
    .Y(_0160_),
    .A1(net851),
    .A2(net772));
 sg13g2_nor2_1 _4071_ (.A(net844),
    .B(_0160_),
    .Y(_0161_));
 sg13g2_xnor2_1 _4072_ (.Y(_0163_),
    .A(net858),
    .B(net747));
 sg13g2_xnor2_1 _4073_ (.Y(_0164_),
    .A(net862),
    .B(net747));
 sg13g2_xnor2_1 _4074_ (.Y(_0165_),
    .A(\flag.flag_abrosexual_inst.pix_y[1] ),
    .B(net747));
 sg13g2_nor3_1 _4075_ (.A(_0163_),
    .B(_0164_),
    .C(_0165_),
    .Y(_0166_));
 sg13g2_nor2_2 _4076_ (.A(net840),
    .B(_0140_),
    .Y(_0167_));
 sg13g2_a22oi_1 _4077_ (.Y(_0168_),
    .B1(_0167_),
    .B2(_0159_),
    .A2(_0166_),
    .A1(_0161_));
 sg13g2_o21ai_1 _4078_ (.B1(net702),
    .Y(_0169_),
    .A1(_0157_),
    .A2(_0168_));
 sg13g2_nor2_1 _4079_ (.A(net839),
    .B(_0579_),
    .Y(_0170_));
 sg13g2_nand2_2 _4080_ (.Y(_0171_),
    .A(_0129_),
    .B(_0590_));
 sg13g2_and2_1 _4081_ (.A(_0601_),
    .B(_0171_),
    .X(_0172_));
 sg13g2_nand2_2 _4082_ (.Y(_0174_),
    .A(_0601_),
    .B(_0171_));
 sg13g2_nor2_2 _4083_ (.A(_0013_),
    .B(net743),
    .Y(_0175_));
 sg13g2_a21oi_1 _4084_ (.A1(net743),
    .A2(_0174_),
    .Y(_0176_),
    .B1(_0175_));
 sg13g2_a21o_2 _4085_ (.A2(_0174_),
    .A1(net743),
    .B1(_0175_),
    .X(_0177_));
 sg13g2_nand3_1 _4086_ (.B(net763),
    .C(_1435_),
    .A(net767),
    .Y(_0178_));
 sg13g2_nand2_1 _4087_ (.Y(_0179_),
    .A(_0169_),
    .B(_0178_));
 sg13g2_nor2_1 _4088_ (.A(net814),
    .B(_0217_),
    .Y(_0180_));
 sg13g2_nor2_2 _4089_ (.A(_2858_),
    .B(_0180_),
    .Y(_0181_));
 sg13g2_xnor2_1 _4090_ (.Y(_0182_),
    .A(net819),
    .B(_0165_));
 sg13g2_o21ai_1 _4091_ (.B1(_0182_),
    .Y(_0183_),
    .A1(net820),
    .A2(_0164_));
 sg13g2_nand2_1 _4092_ (.Y(_0185_),
    .A(_0023_),
    .B(_0165_));
 sg13g2_nand2_1 _4093_ (.Y(_0186_),
    .A(_0183_),
    .B(_0185_));
 sg13g2_nand2_1 _4094_ (.Y(_0187_),
    .A(net816),
    .B(_0163_));
 sg13g2_nor2_1 _4095_ (.A(net816),
    .B(_0163_),
    .Y(_0188_));
 sg13g2_xnor2_1 _4096_ (.Y(_0189_),
    .A(net816),
    .B(_0163_));
 sg13g2_a21oi_1 _4097_ (.A1(_0157_),
    .A2(_0181_),
    .Y(_0190_),
    .B1(_0189_));
 sg13g2_nand2_1 _4098_ (.Y(_0191_),
    .A(net812),
    .B(_0158_));
 sg13g2_xnor2_1 _4099_ (.Y(_0192_),
    .A(net812),
    .B(_0157_));
 sg13g2_nand2_1 _4100_ (.Y(_0193_),
    .A(_0184_),
    .B(_2865_));
 sg13g2_nor2_1 _4101_ (.A(net801),
    .B(_2866_),
    .Y(_0194_));
 sg13g2_a22oi_1 _4102_ (.Y(_0196_),
    .B1(_0194_),
    .B2(_0184_),
    .A2(_0193_),
    .A1(net801));
 sg13g2_inv_1 _4103_ (.Y(_0197_),
    .A(_0196_));
 sg13g2_xor2_1 _4104_ (.B(_0196_),
    .A(net844),
    .X(_0198_));
 sg13g2_xnor2_1 _4105_ (.Y(_0199_),
    .A(net805),
    .B(_1391_));
 sg13g2_nor2_1 _4106_ (.A(net700),
    .B(_0199_),
    .Y(_0200_));
 sg13g2_a22oi_1 _4107_ (.Y(_0201_),
    .B1(_0198_),
    .B2(_0200_),
    .A2(_0197_),
    .A1(net849));
 sg13g2_o21ai_1 _4108_ (.B1(_0201_),
    .Y(_0202_),
    .A1(_0187_),
    .A2(_0192_));
 sg13g2_a21o_1 _4109_ (.A2(_0190_),
    .A1(_0186_),
    .B1(_0202_),
    .X(_0203_));
 sg13g2_a21o_1 _4110_ (.A2(_0164_),
    .A1(net820),
    .B1(_0183_),
    .X(_0204_));
 sg13g2_nand2b_1 _4111_ (.Y(_0205_),
    .B(_0198_),
    .A_N(_0200_));
 sg13g2_a21oi_1 _4112_ (.A1(net700),
    .A2(_0199_),
    .Y(_0207_),
    .B1(_0205_));
 sg13g2_inv_1 _4113_ (.Y(_0208_),
    .A(_0207_));
 sg13g2_nand2_1 _4114_ (.Y(_0209_),
    .A(_0190_),
    .B(_0207_));
 sg13g2_o21ai_1 _4115_ (.B1(_0203_),
    .Y(_0210_),
    .A1(_0204_),
    .A2(_0209_));
 sg13g2_o21ai_1 _4116_ (.B1(_0210_),
    .Y(_0211_),
    .A1(_0157_),
    .A2(_0181_));
 sg13g2_nand2_1 _4117_ (.Y(_0212_),
    .A(net799),
    .B(_1556_));
 sg13g2_xnor2_1 _4118_ (.Y(_0213_),
    .A(net800),
    .B(_1545_));
 sg13g2_a22oi_1 _4119_ (.Y(_0214_),
    .B1(_0213_),
    .B2(net701),
    .A2(_0208_),
    .A1(_0201_));
 sg13g2_or2_1 _4120_ (.X(_0215_),
    .B(_0213_),
    .A(net703));
 sg13g2_xnor2_1 _4121_ (.Y(_0216_),
    .A(_0014_),
    .B(_0212_));
 sg13g2_a22oi_1 _4122_ (.Y(_0218_),
    .B1(_0216_),
    .B2(_0177_),
    .A2(_0214_),
    .A1(_0211_));
 sg13g2_nand2_2 _4123_ (.Y(_0219_),
    .A(net786),
    .B(net791));
 sg13g2_nor2_2 _4124_ (.A(net774),
    .B(_0677_),
    .Y(_0220_));
 sg13g2_nand3_1 _4125_ (.B(_1556_),
    .C(_0220_),
    .A(net785),
    .Y(_0221_));
 sg13g2_o21ai_1 _4126_ (.B1(net775),
    .Y(_0222_),
    .A1(_0677_),
    .A2(_1545_));
 sg13g2_a21oi_1 _4127_ (.A1(_0221_),
    .A2(_0222_),
    .Y(_0223_),
    .B1(net784));
 sg13g2_o21ai_1 _4128_ (.B1(_0223_),
    .Y(_0224_),
    .A1(_0177_),
    .A2(_0216_));
 sg13g2_a21oi_2 _4129_ (.B1(_0224_),
    .Y(_0225_),
    .A2(_0218_),
    .A1(_0215_));
 sg13g2_o21ai_1 _4130_ (.B1(_0225_),
    .Y(_0226_),
    .A1(_0148_),
    .A2(_0152_));
 sg13g2_nor3_1 _4131_ (.A(net675),
    .B(_0179_),
    .C(_0226_),
    .Y(_0227_));
 sg13g2_xor2_1 _4132_ (.B(_0144_),
    .A(_2961_),
    .X(_0229_));
 sg13g2_nand4_1 _4133_ (.B(_0147_),
    .C(_0227_),
    .A(_0146_),
    .Y(_0230_),
    .D(_0229_));
 sg13g2_nor2_2 _4134_ (.A(_0808_),
    .B(_1116_),
    .Y(_0231_));
 sg13g2_nand2b_1 _4135_ (.Y(_0232_),
    .B(_0819_),
    .A_N(_1116_));
 sg13g2_nor2b_2 _4136_ (.A(net750),
    .B_N(_0885_),
    .Y(_0233_));
 sg13g2_nand2b_1 _4137_ (.Y(_0234_),
    .B(_0885_),
    .A_N(net750));
 sg13g2_nand2_2 _4138_ (.Y(_0235_),
    .A(_1204_),
    .B(_0233_));
 sg13g2_nor2_1 _4139_ (.A(net673),
    .B(_0235_),
    .Y(_0236_));
 sg13g2_nand3_1 _4140_ (.B(_0231_),
    .C(_0233_),
    .A(_1204_),
    .Y(_0237_));
 sg13g2_nor2_1 _4141_ (.A(_0158_),
    .B(_0163_),
    .Y(_0238_));
 sg13g2_nor2_2 _4142_ (.A(net849),
    .B(_0159_),
    .Y(_0240_));
 sg13g2_nor2_1 _4143_ (.A(_0158_),
    .B(_0159_),
    .Y(_0241_));
 sg13g2_nand2_1 _4144_ (.Y(_0242_),
    .A(net700),
    .B(_0238_));
 sg13g2_nor2_2 _4145_ (.A(net849),
    .B(_0242_),
    .Y(_0243_));
 sg13g2_nor2_1 _4146_ (.A(net701),
    .B(_0243_),
    .Y(_0244_));
 sg13g2_nor3_2 _4147_ (.A(net701),
    .B(net675),
    .C(_0243_),
    .Y(_0245_));
 sg13g2_nand2_1 _4148_ (.Y(_0246_),
    .A(net785),
    .B(_0245_));
 sg13g2_xnor2_1 _4149_ (.Y(_0247_),
    .A(net675),
    .B(_0244_));
 sg13g2_nand2b_1 _4150_ (.Y(_0248_),
    .B(net790),
    .A_N(_0247_));
 sg13g2_xor2_1 _4151_ (.B(_0242_),
    .A(net844),
    .X(_0249_));
 sg13g2_nor2_2 _4152_ (.A(net769),
    .B(_1709_),
    .Y(_0251_));
 sg13g2_xnor2_1 _4153_ (.Y(_0252_),
    .A(net809),
    .B(_0251_));
 sg13g2_inv_1 _4154_ (.Y(_0253_),
    .A(_0252_));
 sg13g2_a21oi_1 _4155_ (.A1(_0186_),
    .A2(_0187_),
    .Y(_0254_),
    .B1(_0188_));
 sg13g2_inv_1 _4156_ (.Y(_0255_),
    .A(_0254_));
 sg13g2_xnor2_1 _4157_ (.Y(_0256_),
    .A(net700),
    .B(_0238_));
 sg13g2_nand2_1 _4158_ (.Y(_0257_),
    .A(net805),
    .B(_0256_));
 sg13g2_o21ai_1 _4159_ (.B1(_0257_),
    .Y(_0258_),
    .A1(net812),
    .A2(_0251_));
 sg13g2_a21oi_1 _4160_ (.A1(_0252_),
    .A2(_0255_),
    .Y(_0259_),
    .B1(_0258_));
 sg13g2_nand2b_1 _4161_ (.Y(_0260_),
    .B(_0316_),
    .A_N(_0256_));
 sg13g2_xor2_1 _4162_ (.B(_0249_),
    .A(net802),
    .X(_0262_));
 sg13g2_nor2b_1 _4163_ (.A(_0259_),
    .B_N(_0262_),
    .Y(_0263_));
 sg13g2_a22oi_1 _4164_ (.Y(_0264_),
    .B1(_0260_),
    .B2(_0263_),
    .A2(_0249_),
    .A1(net777));
 sg13g2_xnor2_1 _4165_ (.Y(_0265_),
    .A(net796),
    .B(net701));
 sg13g2_nand2_1 _4166_ (.Y(_0266_),
    .A(_0157_),
    .B(_0240_));
 sg13g2_nand2_1 _4167_ (.Y(_0267_),
    .A(net702),
    .B(_0240_));
 sg13g2_nand3_1 _4168_ (.B(_0157_),
    .C(_0240_),
    .A(net702),
    .Y(_0268_));
 sg13g2_xnor2_1 _4169_ (.Y(_0269_),
    .A(net701),
    .B(_0243_));
 sg13g2_xnor2_1 _4170_ (.Y(_0270_),
    .A(_0243_),
    .B(_0265_));
 sg13g2_nand2b_1 _4171_ (.Y(_0271_),
    .B(_0270_),
    .A_N(_0264_));
 sg13g2_o21ai_1 _4172_ (.B1(_0271_),
    .Y(_0273_),
    .A1(net800),
    .A2(_0269_));
 sg13g2_a22oi_1 _4173_ (.Y(_0274_),
    .B1(_0248_),
    .B2(_0273_),
    .A2(_0245_),
    .A1(net785));
 sg13g2_nor2_1 _4174_ (.A(_0189_),
    .B(_0204_),
    .Y(_0275_));
 sg13g2_xnor2_1 _4175_ (.Y(_0276_),
    .A(net775),
    .B(_0245_));
 sg13g2_and2_1 _4176_ (.A(_0252_),
    .B(_0260_),
    .X(_0277_));
 sg13g2_nand4_1 _4177_ (.B(_0257_),
    .C(_0275_),
    .A(_0248_),
    .Y(_0278_),
    .D(_0277_));
 sg13g2_nand2_1 _4178_ (.Y(_0279_),
    .A(_0262_),
    .B(_0270_));
 sg13g2_nor3_1 _4179_ (.A(_0276_),
    .B(_0278_),
    .C(_0279_),
    .Y(_0280_));
 sg13g2_nand2_1 _4180_ (.Y(_0281_),
    .A(net773),
    .B(_0247_));
 sg13g2_o21ai_1 _4181_ (.B1(_0281_),
    .Y(_0282_),
    .A1(_0274_),
    .A2(_0280_));
 sg13g2_nand2_1 _4182_ (.Y(_0284_),
    .A(net781),
    .B(_0282_));
 sg13g2_a21oi_2 _4183_ (.B1(_0284_),
    .Y(_0285_),
    .A2(_0276_),
    .A1(_0246_));
 sg13g2_nand2_1 _4184_ (.Y(_0286_),
    .A(_0140_),
    .B(net803));
 sg13g2_and2_1 _4185_ (.A(_0265_),
    .B(_0286_),
    .X(_0287_));
 sg13g2_a22oi_1 _4186_ (.Y(_0288_),
    .B1(net806),
    .B2(_0159_),
    .A2(net776),
    .A1(net849));
 sg13g2_nand2_1 _4187_ (.Y(_0289_),
    .A(net809),
    .B(_0157_));
 sg13g2_nand2_1 _4188_ (.Y(_0290_),
    .A(_0191_),
    .B(_0289_));
 sg13g2_and2_1 _4189_ (.A(_0186_),
    .B(_0189_),
    .X(_0291_));
 sg13g2_a21o_1 _4190_ (.A2(_0163_),
    .A1(net813),
    .B1(_0291_),
    .X(_0292_));
 sg13g2_a22oi_1 _4191_ (.Y(_0293_),
    .B1(_0290_),
    .B2(_0292_),
    .A2(_0158_),
    .A1(net809));
 sg13g2_nor2b_2 _4192_ (.A(_0204_),
    .B_N(_0189_),
    .Y(_0295_));
 sg13g2_and2_1 _4193_ (.A(_0290_),
    .B(_0295_),
    .X(_0296_));
 sg13g2_nand2_1 _4194_ (.Y(_0297_),
    .A(_0316_),
    .B(net700));
 sg13g2_nor2_1 _4195_ (.A(net791),
    .B(_0176_),
    .Y(_0298_));
 sg13g2_nor2_1 _4196_ (.A(net799),
    .B(net703),
    .Y(_0299_));
 sg13g2_nand3_1 _4197_ (.B(_0296_),
    .C(_0297_),
    .A(_0287_),
    .Y(_0300_));
 sg13g2_nor2_1 _4198_ (.A(_0287_),
    .B(_0299_),
    .Y(_0301_));
 sg13g2_nor2b_1 _4199_ (.A(_0293_),
    .B_N(_0297_),
    .Y(_0302_));
 sg13g2_o21ai_1 _4200_ (.B1(_0300_),
    .Y(_0303_),
    .A1(_0299_),
    .A2(_0302_));
 sg13g2_a21oi_1 _4201_ (.A1(_0288_),
    .A2(_0303_),
    .Y(_0304_),
    .B1(_0301_));
 sg13g2_o21ai_1 _4202_ (.B1(net763),
    .Y(_0306_),
    .A1(_0298_),
    .A2(_0304_));
 sg13g2_a21oi_2 _4203_ (.B1(_0306_),
    .Y(_0307_),
    .A2(net675),
    .A1(net791));
 sg13g2_or2_1 _4204_ (.X(_0308_),
    .B(_0307_),
    .A(_0225_));
 sg13g2_nor2_1 _4205_ (.A(_0285_),
    .B(_0308_),
    .Y(_0309_));
 sg13g2_nor2b_2 _4206_ (.A(net786),
    .B_N(net781),
    .Y(_0310_));
 sg13g2_nand3_1 _4207_ (.B(net675),
    .C(_0240_),
    .A(net703),
    .Y(_0311_));
 sg13g2_nand2_1 _4208_ (.Y(_0312_),
    .A(_0310_),
    .B(_0311_));
 sg13g2_xor2_1 _4209_ (.B(_0311_),
    .A(net785),
    .X(_0313_));
 sg13g2_xnor2_1 _4210_ (.Y(_0314_),
    .A(net675),
    .B(_0267_));
 sg13g2_nand2_1 _4211_ (.Y(_0315_),
    .A(net791),
    .B(_0314_));
 sg13g2_nand3_1 _4212_ (.B(_0313_),
    .C(_0315_),
    .A(net781),
    .Y(_0317_));
 sg13g2_nor2_1 _4213_ (.A(_0161_),
    .B(_0240_),
    .Y(_0318_));
 sg13g2_nor2_1 _4214_ (.A(net803),
    .B(_0318_),
    .Y(_0319_));
 sg13g2_xor2_1 _4215_ (.B(_0318_),
    .A(net801),
    .X(_0320_));
 sg13g2_a21oi_1 _4216_ (.A1(net807),
    .A2(_0159_),
    .Y(_0321_),
    .B1(_0320_));
 sg13g2_nor2_1 _4217_ (.A(net807),
    .B(_0159_),
    .Y(_0322_));
 sg13g2_nand2b_1 _4218_ (.Y(_0323_),
    .B(_0293_),
    .A_N(_0322_));
 sg13g2_a21oi_1 _4219_ (.A1(_0321_),
    .A2(_0323_),
    .Y(_0324_),
    .B1(_0319_));
 sg13g2_xnor2_1 _4220_ (.Y(_0325_),
    .A(_0240_),
    .B(_0265_));
 sg13g2_nor2_1 _4221_ (.A(_0324_),
    .B(_0325_),
    .Y(_0326_));
 sg13g2_or2_1 _4222_ (.X(_0328_),
    .B(_0240_),
    .A(net702));
 sg13g2_a21oi_1 _4223_ (.A1(_0267_),
    .A2(_0328_),
    .Y(_0329_),
    .B1(net800));
 sg13g2_nor2_1 _4224_ (.A(net791),
    .B(_0314_),
    .Y(_0330_));
 sg13g2_nor3_1 _4225_ (.A(_0326_),
    .B(_0329_),
    .C(_0330_),
    .Y(_0331_));
 sg13g2_o21ai_1 _4226_ (.B1(_0312_),
    .Y(_0332_),
    .A1(_0317_),
    .A2(_0331_));
 sg13g2_nor3_1 _4227_ (.A(_0322_),
    .B(_0325_),
    .C(_0330_),
    .Y(_0333_));
 sg13g2_nand3_1 _4228_ (.B(_0321_),
    .C(_0333_),
    .A(_0296_),
    .Y(_0334_));
 sg13g2_o21ai_1 _4229_ (.B1(_0332_),
    .Y(_0335_),
    .A1(_0317_),
    .A2(_0334_));
 sg13g2_nand2_1 _4230_ (.Y(_0336_),
    .A(_0158_),
    .B(_0163_));
 sg13g2_and2_1 _4231_ (.A(_0240_),
    .B(_0336_),
    .X(_0337_));
 sg13g2_o21ai_1 _4232_ (.B1(net675),
    .Y(_0339_),
    .A1(net701),
    .A2(_0337_));
 sg13g2_or3_1 _4233_ (.A(net701),
    .B(net675),
    .C(_0337_),
    .X(_0340_));
 sg13g2_and2_1 _4234_ (.A(_0339_),
    .B(_0340_),
    .X(_0341_));
 sg13g2_o21ai_1 _4235_ (.B1(net781),
    .Y(_0342_),
    .A1(net785),
    .A2(_0339_));
 sg13g2_a221oi_1 _4236_ (.B2(net790),
    .C1(_0342_),
    .B1(_0341_),
    .A1(net785),
    .Y(_0343_),
    .A2(_0339_));
 sg13g2_nand2_1 _4237_ (.Y(_0344_),
    .A(net700),
    .B(_0336_));
 sg13g2_xor2_1 _4238_ (.B(_0344_),
    .A(net844),
    .X(_0345_));
 sg13g2_nand2_1 _4239_ (.Y(_0346_),
    .A(net777),
    .B(_0345_));
 sg13g2_xnor2_1 _4240_ (.Y(_0347_),
    .A(net700),
    .B(_0336_));
 sg13g2_xor2_1 _4241_ (.B(_0345_),
    .A(net802),
    .X(_0348_));
 sg13g2_o21ai_1 _4242_ (.B1(_0348_),
    .Y(_0350_),
    .A1(net805),
    .A2(_0347_));
 sg13g2_nand2_1 _4243_ (.Y(_0351_),
    .A(net805),
    .B(_0347_));
 sg13g2_o21ai_1 _4244_ (.B1(_0351_),
    .Y(_0352_),
    .A1(_0252_),
    .A2(_0254_));
 sg13g2_a21oi_1 _4245_ (.A1(_0217_),
    .A2(_0251_),
    .Y(_0353_),
    .B1(_0352_));
 sg13g2_o21ai_1 _4246_ (.B1(_0346_),
    .Y(_0354_),
    .A1(_0350_),
    .A2(_0353_));
 sg13g2_xor2_1 _4247_ (.B(_0337_),
    .A(net701),
    .X(_0355_));
 sg13g2_xnor2_1 _4248_ (.Y(_0356_),
    .A(_0265_),
    .B(_0337_));
 sg13g2_nand2_1 _4249_ (.Y(_0357_),
    .A(_0354_),
    .B(_0356_));
 sg13g2_nor2_1 _4250_ (.A(net790),
    .B(_0341_),
    .Y(_0358_));
 sg13g2_a21oi_1 _4251_ (.A1(_0228_),
    .A2(_0355_),
    .Y(_0359_),
    .B1(_0358_));
 sg13g2_nand2_1 _4252_ (.Y(_0361_),
    .A(_0357_),
    .B(_0359_));
 sg13g2_a22oi_1 _4253_ (.Y(_0362_),
    .B1(_0343_),
    .B2(_0361_),
    .A2(_0339_),
    .A1(net763));
 sg13g2_nand4_1 _4254_ (.B(_0275_),
    .C(_0351_),
    .A(_0253_),
    .Y(_0363_),
    .D(_0356_));
 sg13g2_nor3_1 _4255_ (.A(_0350_),
    .B(_0358_),
    .C(_0363_),
    .Y(_0364_));
 sg13g2_a21o_2 _4256_ (.A2(_0364_),
    .A1(_0343_),
    .B1(_0362_),
    .X(_0365_));
 sg13g2_and2_1 _4257_ (.A(_0335_),
    .B(_0365_),
    .X(_0366_));
 sg13g2_and2_1 _4258_ (.A(_0177_),
    .B(_0268_),
    .X(_0367_));
 sg13g2_xnor2_1 _4259_ (.Y(_0368_),
    .A(_0177_),
    .B(_0268_));
 sg13g2_nand2_1 _4260_ (.Y(_0369_),
    .A(net790),
    .B(_0368_));
 sg13g2_nand2b_1 _4261_ (.Y(_0370_),
    .B(_0266_),
    .A_N(net702));
 sg13g2_a21o_1 _4262_ (.A2(_0370_),
    .A1(_0268_),
    .B1(net800),
    .X(_0372_));
 sg13g2_xnor2_1 _4263_ (.Y(_0373_),
    .A(net844),
    .B(_0241_));
 sg13g2_nand2_1 _4264_ (.Y(_0374_),
    .A(_0192_),
    .B(_0292_));
 sg13g2_and2_2 _4265_ (.A(net853),
    .B(net850),
    .X(_0375_));
 sg13g2_nand2_2 _4266_ (.Y(_0376_),
    .A(net854),
    .B(net850));
 sg13g2_nor2_2 _4267_ (.A(net853),
    .B(net850),
    .Y(_0377_));
 sg13g2_or2_2 _4268_ (.X(_0378_),
    .B(_0377_),
    .A(_0375_));
 sg13g2_nand2_1 _4269_ (.Y(_0379_),
    .A(net805),
    .B(_0378_));
 sg13g2_nand3_1 _4270_ (.B(_0374_),
    .C(_0379_),
    .A(_0289_),
    .Y(_0380_));
 sg13g2_nor2_1 _4271_ (.A(net805),
    .B(_0378_),
    .Y(_0381_));
 sg13g2_xnor2_1 _4272_ (.Y(_0383_),
    .A(net802),
    .B(_0373_));
 sg13g2_nor2_1 _4273_ (.A(_0381_),
    .B(_0383_),
    .Y(_0384_));
 sg13g2_a22oi_1 _4274_ (.Y(_0385_),
    .B1(_0380_),
    .B2(_0384_),
    .A2(_0373_),
    .A1(net777));
 sg13g2_xor2_1 _4275_ (.B(_0266_),
    .A(_0265_),
    .X(_0386_));
 sg13g2_o21ai_1 _4276_ (.B1(_0372_),
    .Y(_0387_),
    .A1(_0385_),
    .A2(_0386_));
 sg13g2_a22oi_1 _4277_ (.Y(_0388_),
    .B1(_0369_),
    .B2(_0387_),
    .A2(_0367_),
    .A1(net785));
 sg13g2_xnor2_1 _4278_ (.Y(_0389_),
    .A(net786),
    .B(_0367_));
 sg13g2_a21oi_1 _4279_ (.A1(net790),
    .A2(_0368_),
    .Y(_0390_),
    .B1(_0386_));
 sg13g2_and4_1 _4280_ (.A(_0379_),
    .B(_0384_),
    .C(_0389_),
    .D(_0390_),
    .X(_0391_));
 sg13g2_nand3_1 _4281_ (.B(_0295_),
    .C(_0391_),
    .A(_0192_),
    .Y(_0392_));
 sg13g2_nand2b_1 _4282_ (.Y(_0393_),
    .B(_0392_),
    .A_N(_0388_));
 sg13g2_o21ai_1 _4283_ (.B1(_0393_),
    .Y(_0394_),
    .A1(net790),
    .A2(_0368_));
 sg13g2_a21o_1 _4284_ (.A2(_0367_),
    .A1(_0007_),
    .B1(_0389_),
    .X(_0395_));
 sg13g2_nand3_1 _4285_ (.B(_0394_),
    .C(_0395_),
    .A(net781),
    .Y(_0396_));
 sg13g2_nand3_1 _4286_ (.B(_0366_),
    .C(_0396_),
    .A(net747),
    .Y(_0397_));
 sg13g2_a21oi_1 _4287_ (.A1(_0309_),
    .A2(_0397_),
    .Y(_0398_),
    .B1(_0237_));
 sg13g2_nor2_2 _4288_ (.A(_0951_),
    .B(_0984_),
    .Y(_0399_));
 sg13g2_nand2_2 _4289_ (.Y(_0400_),
    .A(_0940_),
    .B(_0973_));
 sg13g2_nor2_2 _4290_ (.A(_0918_),
    .B(_0400_),
    .Y(_0401_));
 sg13g2_nor2b_2 _4291_ (.A(_0841_),
    .B_N(_1270_),
    .Y(_0402_));
 sg13g2_nand2b_1 _4292_ (.Y(_0404_),
    .B(_1270_),
    .A_N(_0841_));
 sg13g2_and2_2 _4293_ (.A(_0401_),
    .B(_0402_),
    .X(_0405_));
 sg13g2_xnor2_1 _4294_ (.Y(_0406_),
    .A(net788),
    .B(net793));
 sg13g2_nor2_1 _4295_ (.A(net797),
    .B(net777),
    .Y(_0407_));
 sg13g2_or2_2 _4296_ (.X(_0408_),
    .B(_0407_),
    .A(_1501_));
 sg13g2_inv_1 _4297_ (.Y(_0409_),
    .A(_0408_));
 sg13g2_nor2_1 _4298_ (.A(_0206_),
    .B(_0217_),
    .Y(_0410_));
 sg13g2_nand2_1 _4299_ (.Y(_0411_),
    .A(net808),
    .B(net810));
 sg13g2_nand2_2 _4300_ (.Y(_0412_),
    .A(_2866_),
    .B(_0411_));
 sg13g2_a21oi_1 _4301_ (.A1(net814),
    .A2(net817),
    .Y(_0413_),
    .B1(net810));
 sg13g2_a21oi_2 _4302_ (.B1(_0413_),
    .Y(_0415_),
    .A2(net761),
    .A1(_0184_));
 sg13g2_a21oi_2 _4303_ (.B1(_0410_),
    .Y(_0416_),
    .A2(_0415_),
    .A1(_2866_));
 sg13g2_a21oi_2 _4304_ (.B1(net767),
    .Y(_0417_),
    .A2(_0416_),
    .A1(_0666_));
 sg13g2_nor2_2 _4305_ (.A(_0228_),
    .B(net776),
    .Y(_0418_));
 sg13g2_a21oi_2 _4306_ (.B1(_0418_),
    .Y(_0419_),
    .A2(_0417_),
    .A1(_0408_));
 sg13g2_a21o_1 _4307_ (.A2(_0419_),
    .A1(_0677_),
    .B1(_1435_),
    .X(_0420_));
 sg13g2_a21oi_2 _4308_ (.B1(_1435_),
    .Y(_0421_),
    .A2(_0419_),
    .A1(_0677_));
 sg13g2_xnor2_1 _4309_ (.Y(_0422_),
    .A(_0406_),
    .B(_0421_));
 sg13g2_nand2_1 _4310_ (.Y(_0423_),
    .A(_0012_),
    .B(_0422_));
 sg13g2_nor2_2 _4311_ (.A(net775),
    .B(net783),
    .Y(_0424_));
 sg13g2_nor2_1 _4312_ (.A(_0644_),
    .B(_0424_),
    .Y(_0426_));
 sg13g2_o21ai_1 _4313_ (.B1(_0219_),
    .Y(_0427_),
    .A1(_0406_),
    .A2(_0420_));
 sg13g2_xor2_1 _4314_ (.B(_0427_),
    .A(_0426_),
    .X(_0428_));
 sg13g2_xnor2_1 _4315_ (.Y(_0429_),
    .A(_0129_),
    .B(_0428_));
 sg13g2_nor2_1 _4316_ (.A(_0423_),
    .B(_0429_),
    .Y(_0430_));
 sg13g2_xnor2_1 _4317_ (.Y(_0431_),
    .A(_0012_),
    .B(_0422_));
 sg13g2_xnor2_1 _4318_ (.Y(_0432_),
    .A(_1622_),
    .B(_0419_));
 sg13g2_inv_1 _4319_ (.Y(_0433_),
    .A(_0432_));
 sg13g2_nand2_1 _4320_ (.Y(_0434_),
    .A(net845),
    .B(_0432_));
 sg13g2_nor2_1 _4321_ (.A(_0431_),
    .B(_0434_),
    .Y(_0435_));
 sg13g2_xor2_1 _4322_ (.B(_0432_),
    .A(net845),
    .X(_0437_));
 sg13g2_xnor2_1 _4323_ (.Y(_0438_),
    .A(_0408_),
    .B(_0417_));
 sg13g2_nor2b_1 _4324_ (.A(_0016_),
    .B_N(_0438_),
    .Y(_0439_));
 sg13g2_nor2b_1 _4325_ (.A(_0439_),
    .B_N(_0437_),
    .Y(_0440_));
 sg13g2_nand2b_2 _4326_ (.Y(_0441_),
    .B(net803),
    .A_N(net807));
 sg13g2_nand2_2 _4327_ (.Y(_0442_),
    .A(net807),
    .B(net776));
 sg13g2_nand2_2 _4328_ (.Y(_0443_),
    .A(_0441_),
    .B(_0442_));
 sg13g2_xor2_1 _4329_ (.B(_0443_),
    .A(_0416_),
    .X(_0444_));
 sg13g2_or2_1 _4330_ (.X(_0445_),
    .B(_0444_),
    .A(_0173_));
 sg13g2_xnor2_1 _4331_ (.Y(_0446_),
    .A(_0151_),
    .B(_0438_));
 sg13g2_xnor2_1 _4332_ (.Y(_0448_),
    .A(_0173_),
    .B(_0444_));
 sg13g2_xnor2_1 _4333_ (.Y(_0449_),
    .A(_0412_),
    .B(_0415_));
 sg13g2_nor2_1 _4334_ (.A(_0019_),
    .B(_0449_),
    .Y(_0450_));
 sg13g2_nor2_1 _4335_ (.A(_0448_),
    .B(_0450_),
    .Y(_0451_));
 sg13g2_nand2_1 _4336_ (.Y(_0452_),
    .A(net761),
    .B(_2854_));
 sg13g2_xnor2_1 _4337_ (.Y(_0453_),
    .A(_0181_),
    .B(_0452_));
 sg13g2_nor2_1 _4338_ (.A(_0022_),
    .B(_0453_),
    .Y(_0454_));
 sg13g2_xnor2_1 _4339_ (.Y(_0455_),
    .A(net857),
    .B(_0449_));
 sg13g2_nor2_1 _4340_ (.A(_0454_),
    .B(_0455_),
    .Y(_0456_));
 sg13g2_xor2_1 _4341_ (.B(_0455_),
    .A(_0454_),
    .X(_0457_));
 sg13g2_a21o_2 _4342_ (.A2(_2927_),
    .A1(net761),
    .B1(_2855_),
    .X(_0459_));
 sg13g2_nor2_1 _4343_ (.A(_0025_),
    .B(_0459_),
    .Y(_0460_));
 sg13g2_xnor2_1 _4344_ (.Y(_0461_),
    .A(net860),
    .B(_0453_));
 sg13g2_nor2_1 _4345_ (.A(_0460_),
    .B(_0461_),
    .Y(_0462_));
 sg13g2_a21oi_1 _4346_ (.A1(_0457_),
    .A2(_0462_),
    .Y(_0463_),
    .B1(_0456_));
 sg13g2_xnor2_1 _4347_ (.Y(_0464_),
    .A(_0448_),
    .B(_0450_));
 sg13g2_nor2_1 _4348_ (.A(_0463_),
    .B(_0464_),
    .Y(_0465_));
 sg13g2_xor2_1 _4349_ (.B(_0446_),
    .A(_0445_),
    .X(_0466_));
 sg13g2_o21ai_1 _4350_ (.B1(_0466_),
    .Y(_0467_),
    .A1(_0451_),
    .A2(_0465_));
 sg13g2_o21ai_1 _4351_ (.B1(_0467_),
    .Y(_0468_),
    .A1(_0445_),
    .A2(_0446_));
 sg13g2_xnor2_1 _4352_ (.Y(_0470_),
    .A(_0437_),
    .B(_0439_));
 sg13g2_a21oi_1 _4353_ (.A1(_0468_),
    .A2(_0470_),
    .Y(_0471_),
    .B1(_0440_));
 sg13g2_inv_1 _4354_ (.Y(_0472_),
    .A(_0471_));
 sg13g2_xor2_1 _4355_ (.B(_0434_),
    .A(_0431_),
    .X(_0473_));
 sg13g2_a21oi_1 _4356_ (.A1(_0472_),
    .A2(_0473_),
    .Y(_0474_),
    .B1(_0435_));
 sg13g2_xor2_1 _4357_ (.B(_0429_),
    .A(_0423_),
    .X(_0475_));
 sg13g2_nor2b_1 _4358_ (.A(_0474_),
    .B_N(_0475_),
    .Y(_0476_));
 sg13g2_nor2_1 _4359_ (.A(_0430_),
    .B(_0476_),
    .Y(_0477_));
 sg13g2_and2_1 _4360_ (.A(_0305_),
    .B(_0428_),
    .X(_0478_));
 sg13g2_nand2_2 _4361_ (.Y(_0479_),
    .A(_0272_),
    .B(_0219_));
 sg13g2_a21oi_1 _4362_ (.A1(_1490_),
    .A2(_0421_),
    .Y(_0481_),
    .B1(_0479_));
 sg13g2_inv_1 _4363_ (.Y(_0482_),
    .A(_0481_));
 sg13g2_a21oi_1 _4364_ (.A1(net793),
    .A2(_0421_),
    .Y(_0483_),
    .B1(net788));
 sg13g2_inv_1 _4365_ (.Y(_0484_),
    .A(_0483_));
 sg13g2_a21oi_1 _4366_ (.A1(net783),
    .A2(_0484_),
    .Y(_0485_),
    .B1(_0481_));
 sg13g2_xnor2_1 _4367_ (.Y(_0486_),
    .A(net828),
    .B(_0485_));
 sg13g2_xor2_1 _4368_ (.B(_0486_),
    .A(_0478_),
    .X(_0487_));
 sg13g2_o21ai_1 _4369_ (.B1(_0487_),
    .Y(_0488_),
    .A1(_0430_),
    .A2(_0476_));
 sg13g2_xnor2_1 _4370_ (.Y(_0489_),
    .A(_0477_),
    .B(_0487_));
 sg13g2_a22oi_1 _4371_ (.Y(_0490_),
    .B1(_0484_),
    .B2(net783),
    .A2(_0482_),
    .A1(net828));
 sg13g2_o21ai_1 _4372_ (.B1(_0488_),
    .Y(_0492_),
    .A1(_0478_),
    .A2(_0486_));
 sg13g2_xor2_1 _4373_ (.B(_0492_),
    .A(_0490_),
    .X(_0493_));
 sg13g2_or2_2 _4374_ (.X(_0494_),
    .B(_0493_),
    .A(_0489_));
 sg13g2_inv_1 _4375_ (.Y(_0495_),
    .A(_0494_));
 sg13g2_xnor2_1 _4376_ (.Y(_0496_),
    .A(_0471_),
    .B(_0473_));
 sg13g2_xor2_1 _4377_ (.B(_0470_),
    .A(_0468_),
    .X(_0497_));
 sg13g2_or3_1 _4378_ (.A(_0451_),
    .B(_0465_),
    .C(_0466_),
    .X(_0498_));
 sg13g2_and2_1 _4379_ (.A(_0467_),
    .B(_0498_),
    .X(_0499_));
 sg13g2_and2_1 _4380_ (.A(_0497_),
    .B(_0499_),
    .X(_0500_));
 sg13g2_xnor2_1 _4381_ (.Y(_0501_),
    .A(_0457_),
    .B(_0462_));
 sg13g2_xnor2_1 _4382_ (.Y(_0503_),
    .A(_0463_),
    .B(_0464_));
 sg13g2_nand2_1 _4383_ (.Y(_0504_),
    .A(_0501_),
    .B(_0503_));
 sg13g2_a21o_1 _4384_ (.A2(_0504_),
    .A1(_0500_),
    .B1(_0496_),
    .X(_0505_));
 sg13g2_xnor2_1 _4385_ (.Y(_0506_),
    .A(_0474_),
    .B(_0475_));
 sg13g2_a21oi_2 _4386_ (.B1(_0494_),
    .Y(_0507_),
    .A2(_0506_),
    .A1(_0505_));
 sg13g2_nand2b_1 _4387_ (.Y(_0508_),
    .B(_0405_),
    .A_N(_0507_));
 sg13g2_nor2b_2 _4388_ (.A(_0885_),
    .B_N(net750),
    .Y(_0509_));
 sg13g2_nand2b_1 _4389_ (.Y(_0510_),
    .B(net750),
    .A_N(_0885_));
 sg13g2_nand2_2 _4390_ (.Y(_0511_),
    .A(_1204_),
    .B(_0509_));
 sg13g2_nor2_1 _4391_ (.A(net673),
    .B(_0511_),
    .Y(_0512_));
 sg13g2_xnor2_1 _4392_ (.Y(_0514_),
    .A(net828),
    .B(_0428_));
 sg13g2_nand2_1 _4393_ (.Y(_0515_),
    .A(net840),
    .B(_0433_));
 sg13g2_xnor2_1 _4394_ (.Y(_0516_),
    .A(net845),
    .B(_0438_));
 sg13g2_nand2b_1 _4395_ (.Y(_0517_),
    .B(_0432_),
    .A_N(net840));
 sg13g2_nand3_1 _4396_ (.B(_0516_),
    .C(_0517_),
    .A(_0515_),
    .Y(_0518_));
 sg13g2_xor2_1 _4397_ (.B(_0444_),
    .A(_0016_),
    .X(_0519_));
 sg13g2_xnor2_1 _4398_ (.Y(_0520_),
    .A(_0173_),
    .B(_0449_));
 sg13g2_nand2b_1 _4399_ (.Y(_0521_),
    .B(_0520_),
    .A_N(_0519_));
 sg13g2_xnor2_1 _4400_ (.Y(_0522_),
    .A(_0338_),
    .B(_0459_));
 sg13g2_nand2b_1 _4401_ (.Y(_0523_),
    .B(_0453_),
    .A_N(net857));
 sg13g2_nand2b_1 _4402_ (.Y(_0525_),
    .B(net857),
    .A_N(_0453_));
 sg13g2_nand3_1 _4403_ (.B(_0523_),
    .C(_0525_),
    .A(_0522_),
    .Y(_0526_));
 sg13g2_nor2_1 _4404_ (.A(_0107_),
    .B(net818),
    .Y(_0527_));
 sg13g2_a21oi_1 _4405_ (.A1(_0025_),
    .A2(net818),
    .Y(_0528_),
    .B1(_0527_));
 sg13g2_nand2b_1 _4406_ (.Y(_0529_),
    .B(_0528_),
    .A_N(_0526_));
 sg13g2_o21ai_1 _4407_ (.B1(_0525_),
    .Y(_0530_),
    .A1(_0118_),
    .A2(_0459_));
 sg13g2_nand2_1 _4408_ (.Y(_0531_),
    .A(_0523_),
    .B(_0530_));
 sg13g2_a21oi_1 _4409_ (.A1(_0529_),
    .A2(_0531_),
    .Y(_0532_),
    .B1(_0521_));
 sg13g2_or3_1 _4410_ (.A(_0002_),
    .B(_0449_),
    .C(_0519_),
    .X(_0533_));
 sg13g2_a21oi_1 _4411_ (.A1(net851),
    .A2(_0444_),
    .Y(_0534_),
    .B1(_0532_));
 sg13g2_a21oi_1 _4412_ (.A1(_0533_),
    .A2(_0534_),
    .Y(_0536_),
    .B1(_0518_));
 sg13g2_nor2_1 _4413_ (.A(_0013_),
    .B(_0422_),
    .Y(_0537_));
 sg13g2_nand3_1 _4414_ (.B(_0438_),
    .C(_0517_),
    .A(net848),
    .Y(_0538_));
 sg13g2_nand2_1 _4415_ (.Y(_0539_),
    .A(_0515_),
    .B(_0538_));
 sg13g2_nor3_1 _4416_ (.A(_0536_),
    .B(_0537_),
    .C(_0539_),
    .Y(_0540_));
 sg13g2_a21oi_1 _4417_ (.A1(_0013_),
    .A2(_0422_),
    .Y(_0541_),
    .B1(_0540_));
 sg13g2_a22oi_1 _4418_ (.Y(_0542_),
    .B1(_0514_),
    .B2(_0541_),
    .A2(_0428_),
    .A1(net833));
 sg13g2_xnor2_1 _4419_ (.Y(_0543_),
    .A(_0063_),
    .B(_1939_));
 sg13g2_nor2_1 _4420_ (.A(_0521_),
    .B(_0526_),
    .Y(_0544_));
 sg13g2_nand3_1 _4421_ (.B(_0543_),
    .C(_0544_),
    .A(net821),
    .Y(_0545_));
 sg13g2_a21oi_1 _4422_ (.A1(_0013_),
    .A2(_0422_),
    .Y(_0547_),
    .B1(_0545_));
 sg13g2_nor2_1 _4423_ (.A(_0518_),
    .B(_0537_),
    .Y(_0548_));
 sg13g2_nand3_1 _4424_ (.B(_0547_),
    .C(_0548_),
    .A(_0514_),
    .Y(_0549_));
 sg13g2_nor2_1 _4425_ (.A(_0482_),
    .B(_0542_),
    .Y(_0550_));
 sg13g2_nand2_1 _4426_ (.Y(_0551_),
    .A(_0004_),
    .B(_0219_));
 sg13g2_xor2_1 _4427_ (.B(_0219_),
    .A(net780),
    .X(_0552_));
 sg13g2_nand2_2 _4428_ (.Y(_0553_),
    .A(net815),
    .B(net810));
 sg13g2_a21oi_2 _4429_ (.B1(net817),
    .Y(_0554_),
    .A2(net814),
    .A1(net824));
 sg13g2_a21oi_1 _4430_ (.A1(_0553_),
    .A2(_0554_),
    .Y(_0555_),
    .B1(_1391_));
 sg13g2_nor2_1 _4431_ (.A(_0412_),
    .B(_0555_),
    .Y(_0556_));
 sg13g2_nor2_2 _4432_ (.A(_2865_),
    .B(_0556_),
    .Y(_0558_));
 sg13g2_a21oi_1 _4433_ (.A1(_0732_),
    .A2(_0558_),
    .Y(_0559_),
    .B1(_0655_));
 sg13g2_a21oi_1 _4434_ (.A1(_0408_),
    .A2(_0559_),
    .Y(_0560_),
    .B1(_1424_));
 sg13g2_o21ai_1 _4435_ (.B1(_0743_),
    .Y(_0561_),
    .A1(_1523_),
    .A2(_0560_));
 sg13g2_nor2_1 _4436_ (.A(net775),
    .B(_0561_),
    .Y(_0562_));
 sg13g2_a21oi_1 _4437_ (.A1(net774),
    .A2(_0014_),
    .Y(_0563_),
    .B1(_0562_));
 sg13g2_xor2_1 _4438_ (.B(_0563_),
    .A(_0552_),
    .X(_0564_));
 sg13g2_nand2_1 _4439_ (.Y(_0565_),
    .A(net833),
    .B(_0564_));
 sg13g2_xnor2_1 _4440_ (.Y(_0566_),
    .A(net788),
    .B(_0561_));
 sg13g2_xnor2_1 _4441_ (.Y(_0567_),
    .A(net828),
    .B(_0564_));
 sg13g2_o21ai_1 _4442_ (.B1(_0567_),
    .Y(_0569_),
    .A1(_0305_),
    .A2(_0566_));
 sg13g2_xnor2_1 _4443_ (.Y(_0570_),
    .A(_1622_),
    .B(_0560_));
 sg13g2_nor2_1 _4444_ (.A(net840),
    .B(_0570_),
    .Y(_0571_));
 sg13g2_xnor2_1 _4445_ (.Y(_0572_),
    .A(_0408_),
    .B(_0559_));
 sg13g2_xor2_1 _4446_ (.B(_0558_),
    .A(_0443_),
    .X(_0573_));
 sg13g2_xor2_1 _4447_ (.B(_0555_),
    .A(_0412_),
    .X(_0574_));
 sg13g2_and2_1 _4448_ (.A(_0002_),
    .B(_0574_),
    .X(_0575_));
 sg13g2_xor2_1 _4449_ (.B(_0573_),
    .A(_0016_),
    .X(_0576_));
 sg13g2_nor2_1 _4450_ (.A(_0002_),
    .B(_0574_),
    .Y(_0577_));
 sg13g2_xor2_1 _4451_ (.B(_0554_),
    .A(_0181_),
    .X(_0578_));
 sg13g2_nand2_1 _4452_ (.Y(_0580_),
    .A(net858),
    .B(_0578_));
 sg13g2_inv_1 _4453_ (.Y(_0581_),
    .A(_0580_));
 sg13g2_nor2_1 _4454_ (.A(net858),
    .B(_0578_),
    .Y(_0582_));
 sg13g2_a21oi_2 _4455_ (.B1(_1380_),
    .Y(_0583_),
    .A2(_2927_),
    .A1(_1358_));
 sg13g2_nand2_1 _4456_ (.Y(_0584_),
    .A(net860),
    .B(_0583_));
 sg13g2_a21oi_1 _4457_ (.A1(_0580_),
    .A2(_0584_),
    .Y(_0585_),
    .B1(_0582_));
 sg13g2_nor2_1 _4458_ (.A(_0025_),
    .B(net818),
    .Y(_0586_));
 sg13g2_a21oi_1 _4459_ (.A1(net818),
    .A2(net771),
    .Y(_0587_),
    .B1(_0586_));
 sg13g2_xnor2_1 _4460_ (.Y(_0588_),
    .A(_0338_),
    .B(_0583_));
 sg13g2_nor4_1 _4461_ (.A(_0576_),
    .B(_0581_),
    .C(_0582_),
    .D(_0588_),
    .Y(_0589_));
 sg13g2_nor4_1 _4462_ (.A(_0581_),
    .B(_0582_),
    .C(_0587_),
    .D(_0588_),
    .Y(_0591_));
 sg13g2_nor3_1 _4463_ (.A(_0577_),
    .B(_0585_),
    .C(_0591_),
    .Y(_0592_));
 sg13g2_nor3_1 _4464_ (.A(_0575_),
    .B(_0576_),
    .C(_0592_),
    .Y(_0593_));
 sg13g2_a21o_1 _4465_ (.A2(_0573_),
    .A1(net851),
    .B1(_0593_),
    .X(_0594_));
 sg13g2_xnor2_1 _4466_ (.Y(_0595_),
    .A(net845),
    .B(_0572_));
 sg13g2_a22oi_1 _4467_ (.Y(_0596_),
    .B1(_0594_),
    .B2(_0595_),
    .A2(_0572_),
    .A1(net848));
 sg13g2_and2_1 _4468_ (.A(_0305_),
    .B(_0566_),
    .X(_0597_));
 sg13g2_nand2_1 _4469_ (.Y(_0598_),
    .A(net840),
    .B(_0570_));
 sg13g2_a21oi_1 _4470_ (.A1(_0596_),
    .A2(_0598_),
    .Y(_0599_),
    .B1(_0571_));
 sg13g2_nor2_1 _4471_ (.A(_0597_),
    .B(_0599_),
    .Y(_0600_));
 sg13g2_o21ai_1 _4472_ (.B1(_0565_),
    .Y(_0602_),
    .A1(_0569_),
    .A2(_0600_));
 sg13g2_nand2_1 _4473_ (.Y(_0603_),
    .A(net827),
    .B(_0543_));
 sg13g2_nor3_1 _4474_ (.A(_0575_),
    .B(_0577_),
    .C(_0603_),
    .Y(_0604_));
 sg13g2_nand4_1 _4475_ (.B(_0595_),
    .C(_0598_),
    .A(_0589_),
    .Y(_0605_),
    .D(_0604_));
 sg13g2_nor4_1 _4476_ (.A(_0569_),
    .B(_0571_),
    .C(_0597_),
    .D(_0605_),
    .Y(_0606_));
 sg13g2_nor2_1 _4477_ (.A(net774),
    .B(_0552_),
    .Y(_0607_));
 sg13g2_o21ai_1 _4478_ (.B1(_0424_),
    .Y(_0608_),
    .A1(net792),
    .A2(net780));
 sg13g2_or3_1 _4479_ (.A(net787),
    .B(net792),
    .C(net780),
    .X(_0609_));
 sg13g2_a221oi_1 _4480_ (.B2(_0609_),
    .C1(_0606_),
    .B1(_0608_),
    .A1(_0561_),
    .Y(_0610_),
    .A2(_0607_));
 sg13g2_a22oi_1 _4481_ (.Y(_0611_),
    .B1(_0602_),
    .B2(_0610_),
    .A2(_0550_),
    .A1(_0549_));
 sg13g2_xnor2_1 _4482_ (.Y(_0613_),
    .A(net745),
    .B(_0611_));
 sg13g2_and2_1 _4483_ (.A(_0512_),
    .B(_0613_),
    .X(_0614_));
 sg13g2_nor2_1 _4484_ (.A(net835),
    .B(_0557_),
    .Y(_0615_));
 sg13g2_nor2_2 _4485_ (.A(net846),
    .B(\flag.flag_abrosexual_inst.pix_y[4] ),
    .Y(_0616_));
 sg13g2_or2_1 _4486_ (.X(_0617_),
    .B(\flag.flag_abrosexual_inst.pix_y[4] ),
    .A(net846));
 sg13g2_nor2_1 _4487_ (.A(net835),
    .B(_0617_),
    .Y(_0618_));
 sg13g2_and2_1 _4488_ (.A(_0403_),
    .B(net762),
    .X(_0619_));
 sg13g2_nand2_1 _4489_ (.Y(_0620_),
    .A(_0403_),
    .B(net762));
 sg13g2_o21ai_1 _4490_ (.B1(net854),
    .Y(_0621_),
    .A1(net856),
    .A2(_1698_));
 sg13g2_a21oi_2 _4491_ (.B1(_0615_),
    .Y(_0622_),
    .A2(_0621_),
    .A1(_0618_));
 sg13g2_nand2_1 _4492_ (.Y(_0624_),
    .A(net832),
    .B(_0616_));
 sg13g2_nor2_1 _4493_ (.A(net768),
    .B(_0624_),
    .Y(_0625_));
 sg13g2_nor3_2 _4494_ (.A(net768),
    .B(_0620_),
    .C(_0624_),
    .Y(_0626_));
 sg13g2_nor2_2 _4495_ (.A(_0622_),
    .B(_0626_),
    .Y(_0627_));
 sg13g2_nor3_2 _4496_ (.A(_1083_),
    .B(_0307_),
    .C(net660),
    .Y(_0628_));
 sg13g2_nor3_2 _4497_ (.A(_1028_),
    .B(_0307_),
    .C(net660),
    .Y(_0629_));
 sg13g2_nor2_2 _4498_ (.A(net842),
    .B(net837),
    .Y(_0630_));
 sg13g2_or2_2 _4499_ (.X(_0631_),
    .B(net837),
    .A(net841));
 sg13g2_nor2_1 _4500_ (.A(net846),
    .B(_0631_),
    .Y(_0632_));
 sg13g2_nor2_2 _4501_ (.A(net778),
    .B(_0632_),
    .Y(_0633_));
 sg13g2_o21ai_1 _4502_ (.B1(net834),
    .Y(_0634_),
    .A1(net847),
    .A2(_0631_));
 sg13g2_a21oi_2 _4503_ (.B1(_0633_),
    .Y(_0635_),
    .A2(_0375_),
    .A1(net834));
 sg13g2_nand2_1 _4504_ (.Y(_0636_),
    .A(_2390_),
    .B(_2393_));
 sg13g2_a21oi_2 _4505_ (.B1(_2845_),
    .Y(_0637_),
    .A2(_2393_),
    .A1(_2390_));
 sg13g2_nor2_1 _4506_ (.A(_2004_),
    .B(_0637_),
    .Y(_0638_));
 sg13g2_nand2_1 _4507_ (.Y(_0639_),
    .A(net724),
    .B(_0638_));
 sg13g2_nor2_1 _4508_ (.A(_0808_),
    .B(_0863_),
    .Y(_0640_));
 sg13g2_nand2_1 _4509_ (.Y(_0641_),
    .A(_0819_),
    .B(_0852_));
 sg13g2_nand2_1 _4510_ (.Y(_0642_),
    .A(_0401_),
    .B(net671));
 sg13g2_o21ai_1 _4511_ (.B1(_1578_),
    .Y(_0643_),
    .A1(net788),
    .A2(_1446_));
 sg13g2_a21oi_1 _4512_ (.A1(net774),
    .A2(_1435_),
    .Y(_0645_),
    .B1(_1512_));
 sg13g2_a22oi_1 _4513_ (.Y(_0646_),
    .B1(_0645_),
    .B2(_1600_),
    .A2(_0643_),
    .A1(_1512_));
 sg13g2_nor4_1 _4514_ (.A(_2004_),
    .B(_2390_),
    .C(net710),
    .D(_2845_),
    .Y(_0647_));
 sg13g2_a21oi_1 _4515_ (.A1(_2355_),
    .A2(_2683_),
    .Y(_0648_),
    .B1(_2370_));
 sg13g2_a21oi_1 _4516_ (.A1(net724),
    .A2(_0647_),
    .Y(_0649_),
    .B1(_0648_));
 sg13g2_nand3_1 _4517_ (.B(_0646_),
    .C(_0649_),
    .A(_0639_),
    .Y(_0650_));
 sg13g2_a21oi_2 _4518_ (.B1(net717),
    .Y(_0651_),
    .A2(net713),
    .A1(_2264_));
 sg13g2_nand2_1 _4519_ (.Y(_0652_),
    .A(net680),
    .B(_0651_));
 sg13g2_xnor2_1 _4520_ (.Y(_0653_),
    .A(_2354_),
    .B(_0651_));
 sg13g2_nand3_1 _4521_ (.B(_2264_),
    .C(net713),
    .A(net717),
    .Y(_0654_));
 sg13g2_nor2b_1 _4522_ (.A(_0651_),
    .B_N(_0654_),
    .Y(_0656_));
 sg13g2_xnor2_1 _4523_ (.Y(_0657_),
    .A(_0173_),
    .B(_2264_));
 sg13g2_inv_1 _4524_ (.Y(_0658_),
    .A(_0657_));
 sg13g2_o21ai_1 _4525_ (.B1(_0156_),
    .Y(_0659_),
    .A1(net744),
    .A2(_0657_));
 sg13g2_nand3_1 _4526_ (.B(_1698_),
    .C(net711),
    .A(net826),
    .Y(_0660_));
 sg13g2_nor3_1 _4527_ (.A(net826),
    .B(_0327_),
    .C(net821),
    .Y(_0661_));
 sg13g2_o21ai_1 _4528_ (.B1(net762),
    .Y(_0662_),
    .A1(_0019_),
    .A2(_0349_));
 sg13g2_o21ai_1 _4529_ (.B1(_0660_),
    .Y(_0663_),
    .A1(_0661_),
    .A2(_0662_));
 sg13g2_a21o_1 _4530_ (.A2(_0659_),
    .A1(_1961_),
    .B1(_0663_),
    .X(_0664_));
 sg13g2_o21ai_1 _4531_ (.B1(_0664_),
    .Y(_0665_),
    .A1(_1961_),
    .A2(_0659_));
 sg13g2_a21oi_1 _4532_ (.A1(net708),
    .A2(_0656_),
    .Y(_0667_),
    .B1(_0665_));
 sg13g2_xnor2_1 _4533_ (.Y(_0668_),
    .A(net714),
    .B(_0652_));
 sg13g2_or2_1 _4534_ (.X(_0669_),
    .B(_0668_),
    .A(net707));
 sg13g2_nand2b_1 _4535_ (.Y(_0670_),
    .B(_2393_),
    .A_N(_0653_));
 sg13g2_a21oi_1 _4536_ (.A1(net714),
    .A2(_0652_),
    .Y(_0671_),
    .B1(net722));
 sg13g2_o21ai_1 _4537_ (.B1(_0670_),
    .Y(_0672_),
    .A1(net708),
    .A2(_0656_));
 sg13g2_a22oi_1 _4538_ (.Y(_0673_),
    .B1(_0668_),
    .B2(net707),
    .A2(_0653_),
    .A1(net710));
 sg13g2_o21ai_1 _4539_ (.B1(_0673_),
    .Y(_0674_),
    .A1(_0667_),
    .A2(_0672_));
 sg13g2_a22oi_1 _4540_ (.Y(_0675_),
    .B1(_0674_),
    .B2(_0669_),
    .A2(_0671_),
    .A1(net705));
 sg13g2_o21ai_1 _4541_ (.B1(_2004_),
    .Y(_0676_),
    .A1(net705),
    .A2(_0671_));
 sg13g2_nor3_1 _4542_ (.A(net725),
    .B(_0675_),
    .C(_0676_),
    .Y(_0678_));
 sg13g2_nand3_1 _4543_ (.B(_0096_),
    .C(net813),
    .A(_0063_),
    .Y(_0679_));
 sg13g2_a22oi_1 _4544_ (.Y(_0680_),
    .B1(_0679_),
    .B2(_1347_),
    .A2(_2395_),
    .A1(net861));
 sg13g2_xnor2_1 _4545_ (.Y(_0681_),
    .A(_2390_),
    .B(net710));
 sg13g2_nand3b_1 _4546_ (.B(_1347_),
    .C(_0025_),
    .Y(_0682_),
    .A_N(net813));
 sg13g2_o21ai_1 _4547_ (.B1(_0682_),
    .Y(_0683_),
    .A1(net719),
    .A2(_0681_));
 sg13g2_xnor2_1 _4548_ (.Y(_0684_),
    .A(net707),
    .B(_0636_));
 sg13g2_a22oi_1 _4549_ (.Y(_0685_),
    .B1(_0684_),
    .B2(net711),
    .A2(_0681_),
    .A1(net719));
 sg13g2_o21ai_1 _4550_ (.B1(_0685_),
    .Y(_0686_),
    .A1(_0680_),
    .A2(_0683_));
 sg13g2_a21oi_1 _4551_ (.A1(net707),
    .A2(_0636_),
    .Y(_0687_),
    .B1(net704));
 sg13g2_nor2_1 _4552_ (.A(_0637_),
    .B(_0687_),
    .Y(_0689_));
 sg13g2_nor2_1 _4553_ (.A(net712),
    .B(_0684_),
    .Y(_0690_));
 sg13g2_a21oi_1 _4554_ (.A1(_2293_),
    .A2(_0689_),
    .Y(_0691_),
    .B1(_0690_));
 sg13g2_xnor2_1 _4555_ (.Y(_0692_),
    .A(_1993_),
    .B(_0637_));
 sg13g2_a22oi_1 _4556_ (.Y(_0693_),
    .B1(_0692_),
    .B2(net717),
    .A2(_0691_),
    .A1(_0686_));
 sg13g2_o21ai_1 _4557_ (.B1(_0693_),
    .Y(_0694_),
    .A1(_2293_),
    .A2(_0689_));
 sg13g2_xnor2_1 _4558_ (.Y(_0695_),
    .A(net724),
    .B(_0638_));
 sg13g2_nor2_1 _4559_ (.A(net717),
    .B(_0692_),
    .Y(_0696_));
 sg13g2_a21oi_1 _4560_ (.A1(net679),
    .A2(_0695_),
    .Y(_0697_),
    .B1(_0696_));
 sg13g2_o21ai_1 _4561_ (.B1(_2472_),
    .Y(_0698_),
    .A1(net679),
    .A2(_0695_));
 sg13g2_a21oi_1 _4562_ (.A1(_0694_),
    .A2(_0697_),
    .Y(_0700_),
    .B1(_0698_));
 sg13g2_a21oi_1 _4563_ (.A1(net679),
    .A2(_0651_),
    .Y(_0701_),
    .B1(_2370_));
 sg13g2_nor3_2 _4564_ (.A(_0678_),
    .B(_0700_),
    .C(_0701_),
    .Y(_0702_));
 sg13g2_nor3_2 _4565_ (.A(_0642_),
    .B(_0650_),
    .C(_0702_),
    .Y(_0703_));
 sg13g2_nor2b_2 _4566_ (.A(net853),
    .B_N(net857),
    .Y(_0704_));
 sg13g2_a21oi_1 _4567_ (.A1(net858),
    .A2(_1698_),
    .Y(_0705_),
    .B1(net853));
 sg13g2_nand2b_1 _4568_ (.Y(_0706_),
    .B(_0631_),
    .A_N(_0705_));
 sg13g2_nor2b_2 _4569_ (.A(net839),
    .B_N(net841),
    .Y(_0707_));
 sg13g2_a21oi_1 _4570_ (.A1(net841),
    .A2(_0617_),
    .Y(_0708_),
    .B1(net838));
 sg13g2_nand4_1 _4571_ (.B(_0616_),
    .C(_0704_),
    .A(net762),
    .Y(_0709_),
    .D(_0707_));
 sg13g2_and2_1 _4572_ (.A(net830),
    .B(_0709_),
    .X(_0711_));
 sg13g2_and3_1 _4573_ (.X(_0712_),
    .A(_0706_),
    .B(_0708_),
    .C(_0711_));
 sg13g2_nand3_1 _4574_ (.B(_0708_),
    .C(_0711_),
    .A(_0706_),
    .Y(_0713_));
 sg13g2_o21ai_1 _4575_ (.B1(net838),
    .Y(_0714_),
    .A1(net841),
    .A2(_0617_));
 sg13g2_o21ai_1 _4576_ (.B1(net768),
    .Y(_0715_),
    .A1(_0129_),
    .A2(_0616_));
 sg13g2_nand2_1 _4577_ (.Y(_0716_),
    .A(net865),
    .B(net828));
 sg13g2_nor2_1 _4578_ (.A(net860),
    .B(net857),
    .Y(_0717_));
 sg13g2_nand2_1 _4579_ (.Y(_0718_),
    .A(net854),
    .B(net839));
 sg13g2_a21oi_2 _4580_ (.B1(_0718_),
    .Y(_0719_),
    .A2(_0717_),
    .A1(_0716_));
 sg13g2_nor3_1 _4581_ (.A(net833),
    .B(_0715_),
    .C(_0719_),
    .Y(_0720_));
 sg13g2_a21oi_2 _4582_ (.B1(net854),
    .Y(_0722_),
    .A2(net857),
    .A1(net860));
 sg13g2_o21ai_1 _4583_ (.B1(_0170_),
    .Y(_0723_),
    .A1(_1829_),
    .A2(_0722_));
 sg13g2_and2_1 _4584_ (.A(net833),
    .B(_0723_),
    .X(_0724_));
 sg13g2_nand2_1 _4585_ (.Y(_0725_),
    .A(net833),
    .B(_0723_));
 sg13g2_nor2_1 _4586_ (.A(net846),
    .B(_0151_),
    .Y(_0726_));
 sg13g2_o21ai_1 _4587_ (.B1(net853),
    .Y(_0727_),
    .A1(net856),
    .A2(_0414_));
 sg13g2_nand2b_1 _4588_ (.Y(_0728_),
    .B(_0726_),
    .A_N(_0727_));
 sg13g2_nand3b_1 _4589_ (.B(net845),
    .C(_0728_),
    .Y(_0729_),
    .A_N(net840));
 sg13g2_a21oi_2 _4590_ (.B1(net693),
    .Y(_0730_),
    .A2(_0729_),
    .A1(net839));
 sg13g2_nor2_2 _4591_ (.A(net740),
    .B(_0730_),
    .Y(_0731_));
 sg13g2_nor2_2 _4592_ (.A(net698),
    .B(_0731_),
    .Y(_0733_));
 sg13g2_nor2_2 _4593_ (.A(_1237_),
    .B(_0400_),
    .Y(_0734_));
 sg13g2_nand3_1 _4594_ (.B(_1226_),
    .C(net672),
    .A(_0973_),
    .Y(_0735_));
 sg13g2_nor2_2 _4595_ (.A(_0918_),
    .B(_1215_),
    .Y(_0736_));
 sg13g2_nand2_2 _4596_ (.Y(_0737_),
    .A(_0907_),
    .B(_1204_));
 sg13g2_nand2_2 _4597_ (.Y(_0738_),
    .A(net672),
    .B(_0736_));
 sg13g2_nand3_1 _4598_ (.B(_0401_),
    .C(net671),
    .A(net749),
    .Y(_0739_));
 sg13g2_a21o_1 _4599_ (.A2(_0739_),
    .A1(_0738_),
    .B1(net745),
    .X(_0740_));
 sg13g2_o21ai_1 _4600_ (.B1(_0740_),
    .Y(_0741_),
    .A1(_0733_),
    .A2(_0735_));
 sg13g2_a221oi_1 _4601_ (.B2(_0635_),
    .C1(_0741_),
    .B1(_0629_),
    .A1(_0627_),
    .Y(_0742_),
    .A2(_0628_));
 sg13g2_nand2b_1 _4602_ (.Y(_0744_),
    .B(_0742_),
    .A_N(_0703_));
 sg13g2_nor2_2 _4603_ (.A(net865),
    .B(net827),
    .Y(_0745_));
 sg13g2_nand2_2 _4604_ (.Y(_0746_),
    .A(_0096_),
    .B(_0107_));
 sg13g2_and2_1 _4605_ (.A(_0125_),
    .B(net758),
    .X(_0747_));
 sg13g2_nand2_1 _4606_ (.Y(_0748_),
    .A(_0125_),
    .B(net758));
 sg13g2_nand2_1 _4607_ (.Y(_0749_),
    .A(net859),
    .B(net769));
 sg13g2_a21oi_2 _4608_ (.B1(_0615_),
    .Y(_0750_),
    .A2(_0749_),
    .A1(_0618_));
 sg13g2_nand2_1 _4609_ (.Y(_0751_),
    .A(net829),
    .B(net769));
 sg13g2_nand3_1 _4610_ (.B(_2059_),
    .C(_0616_),
    .A(_0557_),
    .Y(_0752_));
 sg13g2_nor2_1 _4611_ (.A(_0751_),
    .B(_0752_),
    .Y(_0753_));
 sg13g2_nor2_2 _4612_ (.A(_0750_),
    .B(_0753_),
    .Y(_0755_));
 sg13g2_or2_2 _4613_ (.X(_0756_),
    .B(_0753_),
    .A(_0750_));
 sg13g2_nand2_1 _4614_ (.Y(_0757_),
    .A(_0425_),
    .B(_1709_));
 sg13g2_a21oi_1 _4615_ (.A1(_0469_),
    .A2(_0632_),
    .Y(_0758_),
    .B1(_0757_));
 sg13g2_o21ai_1 _4616_ (.B1(_0634_),
    .Y(_0759_),
    .A1(_0458_),
    .A2(_0758_));
 sg13g2_nor2b_2 _4617_ (.A(_0730_),
    .B_N(_0759_),
    .Y(_0760_));
 sg13g2_or2_1 _4618_ (.X(_0761_),
    .B(_0760_),
    .A(_0755_));
 sg13g2_nand2b_1 _4619_ (.Y(_0762_),
    .B(_0761_),
    .A_N(net740));
 sg13g2_nor2_1 _4620_ (.A(net729),
    .B(_0762_),
    .Y(_0763_));
 sg13g2_nand2_2 _4621_ (.Y(_0764_),
    .A(_1281_),
    .B(_0401_));
 sg13g2_nor3_1 _4622_ (.A(net699),
    .B(_0763_),
    .C(_0764_),
    .Y(_0766_));
 sg13g2_nor2_2 _4623_ (.A(_0819_),
    .B(_1116_),
    .Y(_0767_));
 sg13g2_or2_1 _4624_ (.X(_0768_),
    .B(_1116_),
    .A(_0819_));
 sg13g2_nor2_2 _4625_ (.A(_1061_),
    .B(_1237_),
    .Y(_0769_));
 sg13g2_nand2_2 _4626_ (.Y(_0770_),
    .A(_1050_),
    .B(_1226_));
 sg13g2_nor2_1 _4627_ (.A(_1116_),
    .B(_0770_),
    .Y(_0771_));
 sg13g2_nand2_2 _4628_ (.Y(_0772_),
    .A(_0767_),
    .B(_0769_));
 sg13g2_a21oi_1 _4629_ (.A1(net758),
    .A2(_0755_),
    .Y(_0773_),
    .B1(net741));
 sg13g2_nor2_1 _4630_ (.A(net735),
    .B(_0759_),
    .Y(_0774_));
 sg13g2_nand2_1 _4631_ (.Y(_0775_),
    .A(net693),
    .B(_0745_));
 sg13g2_nand2_1 _4632_ (.Y(_0776_),
    .A(net760),
    .B(_0729_));
 sg13g2_nand3_1 _4633_ (.B(_0775_),
    .C(net658),
    .A(_0756_),
    .Y(_0777_));
 sg13g2_o21ai_1 _4634_ (.B1(_0773_),
    .Y(_0778_),
    .A1(_0774_),
    .A2(_0777_));
 sg13g2_a21oi_1 _4635_ (.A1(net695),
    .A2(_0778_),
    .Y(_0779_),
    .B1(_0772_));
 sg13g2_nand2_2 _4636_ (.Y(_0780_),
    .A(_1248_),
    .B(_0402_));
 sg13g2_nand2_1 _4637_ (.Y(_0781_),
    .A(_0747_),
    .B(net658));
 sg13g2_nand2_1 _4638_ (.Y(_0782_),
    .A(net696),
    .B(net694));
 sg13g2_nand2_2 _4639_ (.Y(_0783_),
    .A(net699),
    .B(net735));
 sg13g2_a21oi_1 _4640_ (.A1(_0781_),
    .A2(_0782_),
    .Y(_0784_),
    .B1(_0780_));
 sg13g2_nand2_1 _4641_ (.Y(_0785_),
    .A(net830),
    .B(net768));
 sg13g2_nor2b_1 _4642_ (.A(net841),
    .B_N(net838),
    .Y(_0787_));
 sg13g2_and2_1 _4643_ (.A(_0612_),
    .B(_0787_),
    .X(_0788_));
 sg13g2_nand3_1 _4644_ (.B(_0414_),
    .C(_0788_),
    .A(_0403_),
    .Y(_0789_));
 sg13g2_a21oi_1 _4645_ (.A1(net838),
    .A2(_0546_),
    .Y(_0790_),
    .B1(_0785_));
 sg13g2_nand2_2 _4646_ (.Y(_0791_),
    .A(_0789_),
    .B(_0790_));
 sg13g2_nor2_1 _4647_ (.A(net831),
    .B(_0630_),
    .Y(_0792_));
 sg13g2_nand2_1 _4648_ (.Y(_0793_),
    .A(_0294_),
    .B(_0631_));
 sg13g2_nor3_1 _4649_ (.A(net829),
    .B(_1709_),
    .C(_1753_),
    .Y(_0794_));
 sg13g2_or2_2 _4650_ (.X(_0795_),
    .B(_0794_),
    .A(net757));
 sg13g2_nand2b_1 _4651_ (.Y(_0796_),
    .B(_0791_),
    .A_N(_0795_));
 sg13g2_nand2_2 _4652_ (.Y(_0798_),
    .A(_1050_),
    .B(_0509_));
 sg13g2_nor2_2 _4653_ (.A(net660),
    .B(_0798_),
    .Y(_0799_));
 sg13g2_nand3b_1 _4654_ (.B(_0796_),
    .C(_0799_),
    .Y(_0800_),
    .A_N(net741));
 sg13g2_nand2_1 _4655_ (.Y(_0801_),
    .A(_0612_),
    .B(_0707_));
 sg13g2_nand3_1 _4656_ (.B(_1720_),
    .C(_0707_),
    .A(_0612_),
    .Y(_0802_));
 sg13g2_inv_1 _4657_ (.Y(_0803_),
    .A(_0802_));
 sg13g2_o21ai_1 _4658_ (.B1(net829),
    .Y(_0804_),
    .A1(_0170_),
    .A2(_0803_));
 sg13g2_a21oi_2 _4659_ (.B1(_0804_),
    .Y(_0805_),
    .A2(_0803_),
    .A1(net779));
 sg13g2_a21o_1 _4660_ (.A2(_0803_),
    .A1(net779),
    .B1(_0804_),
    .X(_0806_));
 sg13g2_nand4_1 _4661_ (.B(net830),
    .C(_1720_),
    .A(net835),
    .Y(_0807_),
    .D(_0616_));
 sg13g2_and2_2 _4662_ (.A(_0785_),
    .B(_0807_),
    .X(_0809_));
 sg13g2_nand2_1 _4663_ (.Y(_0810_),
    .A(_0785_),
    .B(_0807_));
 sg13g2_nor2_1 _4664_ (.A(net837),
    .B(net779),
    .Y(_0811_));
 sg13g2_nor3_2 _4665_ (.A(net837),
    .B(net778),
    .C(_0153_),
    .Y(_0812_));
 sg13g2_nor2_1 _4666_ (.A(net726),
    .B(_0812_),
    .Y(_0813_));
 sg13g2_nand2b_1 _4667_ (.Y(_0814_),
    .B(_0809_),
    .A_N(_0812_));
 sg13g2_nor2_1 _4668_ (.A(_0805_),
    .B(_0813_),
    .Y(_0815_));
 sg13g2_nand2_1 _4669_ (.Y(_0816_),
    .A(net666),
    .B(_0814_));
 sg13g2_nor2_2 _4670_ (.A(_1006_),
    .B(_0510_),
    .Y(_0817_));
 sg13g2_nand2_1 _4671_ (.Y(_0818_),
    .A(_0995_),
    .B(_0509_));
 sg13g2_nand2_1 _4672_ (.Y(_0820_),
    .A(_0402_),
    .B(_0817_));
 sg13g2_o21ai_1 _4673_ (.B1(_0800_),
    .Y(_0821_),
    .A1(_0815_),
    .A2(_0820_));
 sg13g2_nand2_2 _4674_ (.Y(_0822_),
    .A(_0995_),
    .B(_1226_));
 sg13g2_nor2_2 _4675_ (.A(net670),
    .B(_0822_),
    .Y(_0823_));
 sg13g2_nand2_2 _4676_ (.Y(_0824_),
    .A(net695),
    .B(net740));
 sg13g2_and2_1 _4677_ (.A(net697),
    .B(_0759_),
    .X(_0825_));
 sg13g2_inv_1 _4678_ (.Y(_0826_),
    .A(_0825_));
 sg13g2_nand2_1 _4679_ (.Y(_0827_),
    .A(_0824_),
    .B(_0826_));
 sg13g2_nand2_1 _4680_ (.Y(_0828_),
    .A(net658),
    .B(_0827_));
 sg13g2_nor2_2 _4681_ (.A(_0755_),
    .B(_0759_),
    .Y(_0829_));
 sg13g2_nand2b_2 _4682_ (.Y(_0831_),
    .B(_0756_),
    .A_N(_0759_));
 sg13g2_nor2_2 _4683_ (.A(_0400_),
    .B(_0510_),
    .Y(_0832_));
 sg13g2_nand2_2 _4684_ (.Y(_0833_),
    .A(_0399_),
    .B(_0509_));
 sg13g2_nand2_2 _4685_ (.Y(_0834_),
    .A(_0231_),
    .B(_0832_));
 sg13g2_nor2_2 _4686_ (.A(net699),
    .B(net740),
    .Y(_0835_));
 sg13g2_nand2_1 _4687_ (.Y(_0836_),
    .A(net694),
    .B(_0835_));
 sg13g2_nor2_1 _4688_ (.A(_0834_),
    .B(_0836_),
    .Y(_0837_));
 sg13g2_nor3_1 _4689_ (.A(_0829_),
    .B(_0834_),
    .C(_0836_),
    .Y(_0838_));
 sg13g2_a21oi_2 _4690_ (.B1(net698),
    .Y(_0839_),
    .A2(_0729_),
    .A1(net760));
 sg13g2_nand2_2 _4691_ (.Y(_0840_),
    .A(net695),
    .B(net658));
 sg13g2_nor2_2 _4692_ (.A(_0829_),
    .B(_0840_),
    .Y(_0842_));
 sg13g2_nand2_1 _4693_ (.Y(_0843_),
    .A(_0831_),
    .B(_0839_));
 sg13g2_nor2_2 _4694_ (.A(net670),
    .B(_0833_),
    .Y(_0844_));
 sg13g2_nor2_1 _4695_ (.A(_0511_),
    .B(net670),
    .Y(_0845_));
 sg13g2_nand2_1 _4696_ (.Y(_0846_),
    .A(_0843_),
    .B(_0845_));
 sg13g2_o21ai_1 _4697_ (.B1(_0843_),
    .Y(_0847_),
    .A1(_0844_),
    .A2(_0845_));
 sg13g2_nor2_2 _4698_ (.A(_0235_),
    .B(net660),
    .Y(_0848_));
 sg13g2_nand3_1 _4699_ (.B(_1720_),
    .C(_0787_),
    .A(_0612_),
    .Y(_0849_));
 sg13g2_nor2_2 _4700_ (.A(_0129_),
    .B(_0153_),
    .Y(_0850_));
 sg13g2_a21oi_2 _4701_ (.B1(_0294_),
    .Y(_0851_),
    .A2(_0850_),
    .A1(_0849_));
 sg13g2_a21o_1 _4702_ (.A2(_0850_),
    .A1(_0849_),
    .B1(net772),
    .X(_0853_));
 sg13g2_nand2b_2 _4703_ (.Y(_0854_),
    .B(net778),
    .A_N(_0849_));
 sg13g2_and2_2 _4704_ (.A(_0851_),
    .B(_0854_),
    .X(_0855_));
 sg13g2_nand2_1 _4705_ (.Y(_0856_),
    .A(_0851_),
    .B(_0854_));
 sg13g2_nor2_2 _4706_ (.A(net831),
    .B(_0714_),
    .Y(_0857_));
 sg13g2_or2_2 _4707_ (.X(_0858_),
    .B(_0857_),
    .A(net747));
 sg13g2_nor2_1 _4708_ (.A(net742),
    .B(net737),
    .Y(_0859_));
 sg13g2_nand2_1 _4709_ (.Y(_0860_),
    .A(net746),
    .B(net731));
 sg13g2_nor3_1 _4710_ (.A(net690),
    .B(_0857_),
    .C(_0859_),
    .Y(_0861_));
 sg13g2_nand2b_1 _4711_ (.Y(_0862_),
    .B(_0848_),
    .A_N(_0861_));
 sg13g2_o21ai_1 _4712_ (.B1(net755),
    .Y(_0864_),
    .A1(_0714_),
    .A2(_0746_));
 sg13g2_a21oi_1 _4713_ (.A1(net742),
    .A2(_0864_),
    .Y(_0865_),
    .B1(_1105_));
 sg13g2_nand2_2 _4714_ (.Y(_0866_),
    .A(_0233_),
    .B(_0399_));
 sg13g2_nor2_2 _4715_ (.A(net661),
    .B(_0866_),
    .Y(_0867_));
 sg13g2_nor2_1 _4716_ (.A(net674),
    .B(_0822_),
    .Y(_0868_));
 sg13g2_nor2_1 _4717_ (.A(_0867_),
    .B(_0868_),
    .Y(_0869_));
 sg13g2_a21oi_1 _4718_ (.A1(net737),
    .A2(net756),
    .Y(_0870_),
    .B1(_0869_));
 sg13g2_o21ai_1 _4719_ (.B1(net687),
    .Y(_0871_),
    .A1(_0865_),
    .A2(_0870_));
 sg13g2_nand2_2 _4720_ (.Y(_0872_),
    .A(_0862_),
    .B(_0871_));
 sg13g2_nor2_2 _4721_ (.A(net661),
    .B(_0770_),
    .Y(_0873_));
 sg13g2_nand2_2 _4722_ (.Y(_0875_),
    .A(_0402_),
    .B(_0769_));
 sg13g2_nor3_1 _4723_ (.A(net768),
    .B(_0623_),
    .C(_1731_),
    .Y(_0876_));
 sg13g2_o21ai_1 _4724_ (.B1(net830),
    .Y(_0877_),
    .A1(_0601_),
    .A2(_0876_));
 sg13g2_and2_1 _4725_ (.A(net778),
    .B(_0876_),
    .X(_0878_));
 sg13g2_nor3_1 _4726_ (.A(net732),
    .B(_0877_),
    .C(_0878_),
    .Y(_0879_));
 sg13g2_nor2_1 _4727_ (.A(net727),
    .B(_0879_),
    .Y(_0880_));
 sg13g2_o21ai_1 _4728_ (.B1(_0634_),
    .Y(_0881_),
    .A1(net778),
    .A2(net732));
 sg13g2_o21ai_1 _4729_ (.B1(_0877_),
    .Y(_0882_),
    .A1(net755),
    .A2(_0881_));
 sg13g2_a21oi_2 _4730_ (.B1(_0875_),
    .Y(_0883_),
    .A2(_0882_),
    .A1(_0880_));
 sg13g2_nor2_1 _4731_ (.A(_1061_),
    .B(_0234_),
    .Y(_0884_));
 sg13g2_nand2_2 _4732_ (.Y(_0886_),
    .A(_1050_),
    .B(_0233_));
 sg13g2_nand2_1 _4733_ (.Y(_0887_),
    .A(_1270_),
    .B(_0884_));
 sg13g2_nor2_2 _4734_ (.A(_0841_),
    .B(_0887_),
    .Y(_0888_));
 sg13g2_nor2_2 _4735_ (.A(_1028_),
    .B(net670),
    .Y(_0889_));
 sg13g2_or2_1 _4736_ (.X(_0890_),
    .B(_0798_),
    .A(net664));
 sg13g2_inv_1 _4737_ (.Y(_0891_),
    .A(_0890_));
 sg13g2_nor2_2 _4738_ (.A(_0633_),
    .B(net726),
    .Y(_0892_));
 sg13g2_nand2_2 _4739_ (.Y(_0893_),
    .A(_0634_),
    .B(net728));
 sg13g2_nor2_2 _4740_ (.A(net765),
    .B(net739),
    .Y(_0894_));
 sg13g2_nor2_1 _4741_ (.A(net727),
    .B(_0894_),
    .Y(_0895_));
 sg13g2_inv_2 _4742_ (.Y(_0897_),
    .A(_0895_));
 sg13g2_nor2_2 _4743_ (.A(_1006_),
    .B(_0234_),
    .Y(_0898_));
 sg13g2_nand2_2 _4744_ (.Y(_0899_),
    .A(_0995_),
    .B(_0233_));
 sg13g2_nor2_2 _4745_ (.A(net661),
    .B(_0899_),
    .Y(_0900_));
 sg13g2_nor2_2 _4746_ (.A(net664),
    .B(_0866_),
    .Y(_0901_));
 sg13g2_nor2_2 _4747_ (.A(net669),
    .B(_0886_),
    .Y(_0902_));
 sg13g2_nand2_2 _4748_ (.Y(_0903_),
    .A(net671),
    .B(_0898_));
 sg13g2_nor2_2 _4749_ (.A(net765),
    .B(net733),
    .Y(_0904_));
 sg13g2_a21oi_1 _4750_ (.A1(net659),
    .A2(_0831_),
    .Y(_0905_),
    .B1(net730));
 sg13g2_nor3_2 _4751_ (.A(net699),
    .B(_0903_),
    .C(_0905_),
    .Y(_0906_));
 sg13g2_nand2_2 _4752_ (.Y(_0908_),
    .A(_0231_),
    .B(_0401_));
 sg13g2_nor2_2 _4753_ (.A(_1028_),
    .B(net668),
    .Y(_0909_));
 sg13g2_nor2_2 _4754_ (.A(_1083_),
    .B(net669),
    .Y(_0910_));
 sg13g2_nand2_2 _4755_ (.Y(_0911_),
    .A(_0513_),
    .B(_0634_));
 sg13g2_nor2_1 _4756_ (.A(_0908_),
    .B(_0911_),
    .Y(_0912_));
 sg13g2_nor2_2 _4757_ (.A(net668),
    .B(_0899_),
    .Y(_0913_));
 sg13g2_a21oi_1 _4758_ (.A1(_0853_),
    .A2(_0911_),
    .Y(_0914_),
    .B1(_0908_));
 sg13g2_a221oi_1 _4759_ (.B2(net692),
    .C1(_0910_),
    .B1(_0913_),
    .A1(net754),
    .Y(_0915_),
    .A2(_0909_));
 sg13g2_nand2b_1 _4760_ (.Y(_0916_),
    .B(_0915_),
    .A_N(_0914_));
 sg13g2_nor2_2 _4761_ (.A(net699),
    .B(_0755_),
    .Y(_0917_));
 sg13g2_nand2_2 _4762_ (.Y(_0919_),
    .A(net671),
    .B(_0817_));
 sg13g2_inv_1 _4763_ (.Y(_0920_),
    .A(_0919_));
 sg13g2_a21oi_1 _4764_ (.A1(net659),
    .A2(_0917_),
    .Y(_0921_),
    .B1(_0919_));
 sg13g2_a21oi_1 _4765_ (.A1(net808),
    .A2(_0413_),
    .Y(_0922_),
    .B1(net806));
 sg13g2_nor2b_1 _4766_ (.A(_0922_),
    .B_N(_1501_),
    .Y(_0923_));
 sg13g2_o21ai_1 _4767_ (.B1(_0310_),
    .Y(_0924_),
    .A1(_0677_),
    .A2(_0923_));
 sg13g2_nand2_1 _4768_ (.Y(_0925_),
    .A(_2858_),
    .B(_0527_));
 sg13g2_nor4_1 _4769_ (.A(_1622_),
    .B(_0409_),
    .C(_0442_),
    .D(_0925_),
    .Y(_0926_));
 sg13g2_a21o_2 _4770_ (.A2(_0926_),
    .A1(net763),
    .B1(_0924_),
    .X(_0927_));
 sg13g2_inv_1 _4771_ (.Y(_0928_),
    .A(_0927_));
 sg13g2_nor2_2 _4772_ (.A(net673),
    .B(_0770_),
    .Y(_0930_));
 sg13g2_nand2_1 _4773_ (.Y(_0931_),
    .A(net731),
    .B(_0805_));
 sg13g2_and2_2 _4774_ (.A(_0402_),
    .B(_0734_),
    .X(_0932_));
 sg13g2_nand3_1 _4775_ (.B(_0931_),
    .C(_0932_),
    .A(net764),
    .Y(_0933_));
 sg13g2_nand2_2 _4776_ (.Y(_0934_),
    .A(net666),
    .B(net726));
 sg13g2_nor2_2 _4777_ (.A(net673),
    .B(_0798_),
    .Y(_0935_));
 sg13g2_a21oi_1 _4778_ (.A1(net736),
    .A2(net659),
    .Y(_0936_),
    .B1(net693));
 sg13g2_nor2_2 _4779_ (.A(net662),
    .B(_0899_),
    .Y(_0937_));
 sg13g2_nand2_1 _4780_ (.Y(_0938_),
    .A(_1281_),
    .B(_0898_));
 sg13g2_nand2_2 _4781_ (.Y(_0939_),
    .A(net740),
    .B(net735));
 sg13g2_nand2_2 _4782_ (.Y(_0941_),
    .A(net696),
    .B(_0939_));
 sg13g2_nor3_1 _4783_ (.A(_0936_),
    .B(_0938_),
    .C(_0941_),
    .Y(_0942_));
 sg13g2_nand2b_1 _4784_ (.Y(_0943_),
    .B(net831),
    .A_N(net837));
 sg13g2_a21oi_2 _4785_ (.B1(_0943_),
    .Y(_0944_),
    .A2(_0375_),
    .A1(_0579_));
 sg13g2_a21o_2 _4786_ (.A2(_0375_),
    .A1(_0579_),
    .B1(_0943_),
    .X(_0945_));
 sg13g2_nand2_1 _4787_ (.Y(_0946_),
    .A(net733),
    .B(net751));
 sg13g2_nand2_1 _4788_ (.Y(_0947_),
    .A(_0579_),
    .B(_0811_));
 sg13g2_o21ai_1 _4789_ (.B1(net766),
    .Y(_0948_),
    .A1(_0377_),
    .A2(_0947_));
 sg13g2_nor2_2 _4790_ (.A(net746),
    .B(_0948_),
    .Y(_0949_));
 sg13g2_nand2b_1 _4791_ (.Y(_0950_),
    .B(_1818_),
    .A_N(_0948_));
 sg13g2_nand2_2 _4792_ (.Y(_0952_),
    .A(_1072_),
    .B(_1281_));
 sg13g2_and2_2 _4793_ (.A(net742),
    .B(_0948_),
    .X(_0953_));
 sg13g2_nand2_2 _4794_ (.Y(_0954_),
    .A(net742),
    .B(_0948_));
 sg13g2_nor2_2 _4795_ (.A(_1028_),
    .B(net664),
    .Y(_0955_));
 sg13g2_nand2_1 _4796_ (.Y(_0956_),
    .A(_0954_),
    .B(_0955_));
 sg13g2_o21ai_1 _4797_ (.B1(_0956_),
    .Y(_0957_),
    .A1(_0949_),
    .A2(_0952_));
 sg13g2_nand2_1 _4798_ (.Y(_0958_),
    .A(_0946_),
    .B(_0957_));
 sg13g2_nor2_2 _4799_ (.A(net660),
    .B(_0822_),
    .Y(_0959_));
 sg13g2_nand2_1 _4800_ (.Y(_0960_),
    .A(net695),
    .B(_0959_));
 sg13g2_nand2_1 _4801_ (.Y(_0961_),
    .A(net741),
    .B(net730));
 sg13g2_nor2_1 _4802_ (.A(_0730_),
    .B(_0960_),
    .Y(_0963_));
 sg13g2_nor2_2 _4803_ (.A(_0634_),
    .B(net727),
    .Y(_0964_));
 sg13g2_nand2_2 _4804_ (.Y(_0965_),
    .A(_0633_),
    .B(net728));
 sg13g2_a21oi_1 _4805_ (.A1(net765),
    .A2(net739),
    .Y(_0966_),
    .B1(_0965_));
 sg13g2_o21ai_1 _4806_ (.B1(_0964_),
    .Y(_0967_),
    .A1(_1149_),
    .A2(net731));
 sg13g2_a21oi_2 _4807_ (.B1(_0805_),
    .Y(_0968_),
    .A2(net726),
    .A1(net739));
 sg13g2_o21ai_1 _4808_ (.B1(net666),
    .Y(_0969_),
    .A1(net731),
    .A2(_0809_));
 sg13g2_nor2_1 _4809_ (.A(_0746_),
    .B(net667),
    .Y(_0970_));
 sg13g2_nor2_2 _4810_ (.A(_1083_),
    .B(net670),
    .Y(_0971_));
 sg13g2_o21ai_1 _4811_ (.B1(_0971_),
    .Y(_0972_),
    .A1(net758),
    .A2(net667));
 sg13g2_o21ai_1 _4812_ (.B1(_0971_),
    .Y(_0974_),
    .A1(_0966_),
    .A2(_0969_));
 sg13g2_nor2_1 _4813_ (.A(_0970_),
    .B(_0974_),
    .Y(_0975_));
 sg13g2_nor2_2 _4814_ (.A(net760),
    .B(_0805_),
    .Y(_0976_));
 sg13g2_nand2_1 _4815_ (.Y(_0977_),
    .A(net764),
    .B(net666));
 sg13g2_nor2_2 _4816_ (.A(net674),
    .B(_0866_),
    .Y(_0978_));
 sg13g2_nor2_2 _4817_ (.A(net668),
    .B(_0833_),
    .Y(_0979_));
 sg13g2_a22oi_1 _4818_ (.Y(_0980_),
    .B1(_0979_),
    .B2(_0839_),
    .A2(_0978_),
    .A1(_0976_));
 sg13g2_o21ai_1 _4819_ (.B1(_0813_),
    .Y(_0981_),
    .A1(_0633_),
    .A2(net733));
 sg13g2_nand2_1 _4820_ (.Y(_0982_),
    .A(net667),
    .B(_0981_));
 sg13g2_nor2_1 _4821_ (.A(_1116_),
    .B(_1259_),
    .Y(_0983_));
 sg13g2_nor2_1 _4822_ (.A(_1259_),
    .B(net669),
    .Y(_0985_));
 sg13g2_nand2_1 _4823_ (.Y(_0986_),
    .A(_1248_),
    .B(_0767_));
 sg13g2_nor2_2 _4824_ (.A(net662),
    .B(_0833_),
    .Y(_0987_));
 sg13g2_nand2_1 _4825_ (.Y(_0988_),
    .A(net733),
    .B(net691));
 sg13g2_and3_1 _4826_ (.X(_0989_),
    .A(_1720_),
    .B(_0707_),
    .C(_0726_));
 sg13g2_o21ai_1 _4827_ (.B1(net830),
    .Y(_0990_),
    .A1(_0708_),
    .A2(_0989_));
 sg13g2_a21o_2 _4828_ (.A2(_0989_),
    .A1(net778),
    .B1(_0990_),
    .X(_0991_));
 sg13g2_nand2_2 _4829_ (.Y(_0992_),
    .A(net734),
    .B(net756));
 sg13g2_nand3_1 _4830_ (.B(net732),
    .C(net755),
    .A(_0715_),
    .Y(_0993_));
 sg13g2_nand3_1 _4831_ (.B(_0991_),
    .C(_0993_),
    .A(_0988_),
    .Y(_0994_));
 sg13g2_nand2_1 _4832_ (.Y(_0996_),
    .A(_0734_),
    .B(_0767_));
 sg13g2_nor2b_1 _4833_ (.A(_0996_),
    .B_N(_0946_),
    .Y(_0997_));
 sg13g2_nand2_1 _4834_ (.Y(_0998_),
    .A(net733),
    .B(_0949_));
 sg13g2_nor2_2 _4835_ (.A(_0235_),
    .B(net670),
    .Y(_0999_));
 sg13g2_o21ai_1 _4836_ (.B1(_0999_),
    .Y(_1000_),
    .A1(_0904_),
    .A2(_0965_));
 sg13g2_nor2_1 _4837_ (.A(net670),
    .B(_0798_),
    .Y(_1001_));
 sg13g2_nand2_1 _4838_ (.Y(_1002_),
    .A(_0949_),
    .B(_1001_));
 sg13g2_o21ai_1 _4839_ (.B1(_1001_),
    .Y(_1003_),
    .A1(net751),
    .A2(_0949_));
 sg13g2_nor2_2 _4840_ (.A(net662),
    .B(_0235_),
    .Y(_1004_));
 sg13g2_a21o_2 _4841_ (.A2(_0546_),
    .A1(net772),
    .B1(net755),
    .X(_1005_));
 sg13g2_nor2_2 _4842_ (.A(net673),
    .B(_0886_),
    .Y(_1007_));
 sg13g2_nor4_1 _4843_ (.A(net674),
    .B(_0886_),
    .C(net751),
    .D(_1005_),
    .Y(_1008_));
 sg13g2_nand2_2 _4844_ (.Y(_1009_),
    .A(_0231_),
    .B(_0736_));
 sg13g2_nor2_2 _4845_ (.A(net742),
    .B(_1009_),
    .Y(_1010_));
 sg13g2_nand3_1 _4846_ (.B(_1226_),
    .C(_0767_),
    .A(_0995_),
    .Y(_1011_));
 sg13g2_nor2_1 _4847_ (.A(net664),
    .B(_0886_),
    .Y(_1012_));
 sg13g2_nor2_1 _4848_ (.A(_0235_),
    .B(net669),
    .Y(_1013_));
 sg13g2_nor2_1 _4849_ (.A(_1012_),
    .B(_1013_),
    .Y(_1014_));
 sg13g2_inv_1 _4850_ (.Y(_1015_),
    .A(_1014_));
 sg13g2_nor2_2 _4851_ (.A(net664),
    .B(_0818_),
    .Y(_1016_));
 sg13g2_nor2_2 _4852_ (.A(net674),
    .B(_0818_),
    .Y(_1018_));
 sg13g2_nand2_1 _4853_ (.Y(_1019_),
    .A(_0966_),
    .B(_1018_));
 sg13g2_nor2_2 _4854_ (.A(net664),
    .B(_0511_),
    .Y(_1020_));
 sg13g2_nor2_2 _4855_ (.A(_1083_),
    .B(net673),
    .Y(_1021_));
 sg13g2_nor2_2 _4856_ (.A(_0511_),
    .B(net668),
    .Y(_1022_));
 sg13g2_nand3_1 _4857_ (.B(_0631_),
    .C(_1022_),
    .A(net834),
    .Y(_1023_));
 sg13g2_nor3_2 _4858_ (.A(_1237_),
    .B(net674),
    .C(_0400_),
    .Y(_1024_));
 sg13g2_and2_1 _4859_ (.A(net764),
    .B(_1024_),
    .X(_1025_));
 sg13g2_nand3_1 _4860_ (.B(net739),
    .C(_0964_),
    .A(net764),
    .Y(_1026_));
 sg13g2_o21ai_1 _4861_ (.B1(_1026_),
    .Y(_1027_),
    .A1(net731),
    .A2(net728));
 sg13g2_nand2_1 _4862_ (.Y(_1029_),
    .A(net666),
    .B(_1027_));
 sg13g2_nor2_2 _4863_ (.A(_1259_),
    .B(net674),
    .Y(_1030_));
 sg13g2_nor2_2 _4864_ (.A(net664),
    .B(_0737_),
    .Y(_1031_));
 sg13g2_nand2_2 _4865_ (.Y(_1032_),
    .A(net745),
    .B(net735));
 sg13g2_nand2_1 _4866_ (.Y(_1033_),
    .A(_0945_),
    .B(_1032_));
 sg13g2_nand2_2 _4867_ (.Y(_1034_),
    .A(net738),
    .B(net751));
 sg13g2_nand2_1 _4868_ (.Y(_1035_),
    .A(_1033_),
    .B(_1034_));
 sg13g2_and2_2 _4869_ (.A(_1281_),
    .B(_0734_),
    .X(_1036_));
 sg13g2_o21ai_1 _4870_ (.B1(_1036_),
    .Y(_1037_),
    .A1(_0814_),
    .A2(_0904_));
 sg13g2_nand2_2 _4871_ (.Y(_1038_),
    .A(_1017_),
    .B(_0231_));
 sg13g2_or2_1 _4872_ (.X(_1040_),
    .B(_1038_),
    .A(_0917_));
 sg13g2_o21ai_1 _4873_ (.B1(net780),
    .Y(_1041_),
    .A1(net796),
    .A2(_0923_));
 sg13g2_nor2_1 _4874_ (.A(_1534_),
    .B(_0442_),
    .Y(_1042_));
 sg13g2_nor4_1 _4875_ (.A(net782),
    .B(_1534_),
    .C(_0442_),
    .D(_0925_),
    .Y(_1043_));
 sg13g2_or2_1 _4876_ (.X(_1044_),
    .B(_1043_),
    .A(_1041_));
 sg13g2_nand2b_1 _4877_ (.Y(_1045_),
    .B(_1044_),
    .A_N(_0310_));
 sg13g2_a21oi_1 _4878_ (.A1(net761),
    .A2(_0180_),
    .Y(_1046_),
    .B1(_0020_));
 sg13g2_nor3_1 _4879_ (.A(net814),
    .B(_0217_),
    .C(_2861_),
    .Y(_1047_));
 sg13g2_nor2_1 _4880_ (.A(_1046_),
    .B(_1047_),
    .Y(_1048_));
 sg13g2_nor2_1 _4881_ (.A(_1446_),
    .B(_0441_),
    .Y(_1049_));
 sg13g2_a21oi_1 _4882_ (.A1(_1048_),
    .A2(_1049_),
    .Y(_1051_),
    .B1(_1457_));
 sg13g2_or2_1 _4883_ (.X(_1052_),
    .B(_1051_),
    .A(net782));
 sg13g2_nor2_1 _4884_ (.A(_1314_),
    .B(_0125_),
    .Y(_1053_));
 sg13g2_nand4_1 _4885_ (.B(_1045_),
    .C(_1052_),
    .A(_0219_),
    .Y(_1054_),
    .D(_1053_));
 sg13g2_nor2_1 _4886_ (.A(_0743_),
    .B(_0441_),
    .Y(_1055_));
 sg13g2_nor2b_1 _4887_ (.A(_1046_),
    .B_N(_1055_),
    .Y(_1056_));
 sg13g2_o21ai_1 _4888_ (.B1(net794),
    .Y(_1057_),
    .A1(net797),
    .A2(net803));
 sg13g2_a21oi_1 _4889_ (.A1(_1047_),
    .A2(_1055_),
    .Y(_1058_),
    .B1(net782));
 sg13g2_o21ai_1 _4890_ (.B1(_1058_),
    .Y(_1059_),
    .A1(_1056_),
    .A2(_1057_));
 sg13g2_nor2_1 _4891_ (.A(net787),
    .B(_1059_),
    .Y(_1060_));
 sg13g2_or2_1 _4892_ (.X(_1062_),
    .B(_1052_),
    .A(net729));
 sg13g2_nand2_1 _4893_ (.Y(_1063_),
    .A(_1314_),
    .B(net758));
 sg13g2_nand4_1 _4894_ (.B(_0927_),
    .C(_1062_),
    .A(net693),
    .Y(_1064_),
    .D(_1063_));
 sg13g2_nor4_1 _4895_ (.A(net698),
    .B(_0829_),
    .C(_1060_),
    .D(_1064_),
    .Y(_1065_));
 sg13g2_nor2_2 _4896_ (.A(net670),
    .B(_0770_),
    .Y(_1066_));
 sg13g2_o21ai_1 _4897_ (.B1(_1066_),
    .Y(_1067_),
    .A1(net698),
    .A2(_0731_));
 sg13g2_nand2_1 _4898_ (.Y(_1068_),
    .A(_0824_),
    .B(_1066_));
 sg13g2_a21oi_1 _4899_ (.A1(_1054_),
    .A2(_1065_),
    .Y(_1069_),
    .B1(_1067_));
 sg13g2_a21oi_1 _4900_ (.A1(net760),
    .A2(_0729_),
    .Y(_1070_),
    .B1(net735));
 sg13g2_nand2_1 _4901_ (.Y(_1071_),
    .A(net729),
    .B(net658));
 sg13g2_nor2_1 _4902_ (.A(net735),
    .B(_0756_),
    .Y(_1073_));
 sg13g2_nand3_1 _4903_ (.B(_0835_),
    .C(_1071_),
    .A(_0761_),
    .Y(_1074_));
 sg13g2_nor2_2 _4904_ (.A(_0641_),
    .B(_0886_),
    .Y(_1075_));
 sg13g2_nand3_1 _4905_ (.B(_1074_),
    .C(_1075_),
    .A(_0783_),
    .Y(_1076_));
 sg13g2_nand2b_1 _4906_ (.Y(_1077_),
    .B(_0788_),
    .A_N(_0436_));
 sg13g2_a22oi_1 _4907_ (.Y(_1078_),
    .B1(_0850_),
    .B2(_1077_),
    .A2(_0788_),
    .A1(_0491_));
 sg13g2_a21oi_1 _4908_ (.A1(_1698_),
    .A2(_0704_),
    .Y(_1079_),
    .B1(_0173_));
 sg13g2_nand2_1 _4909_ (.Y(_1080_),
    .A(_1742_),
    .B(_0707_));
 sg13g2_o21ai_1 _4910_ (.B1(_0013_),
    .Y(_1081_),
    .A1(_1079_),
    .A2(_1080_));
 sg13g2_inv_1 _4911_ (.Y(_1082_),
    .A(_1081_));
 sg13g2_nand2_1 _4912_ (.Y(_1084_),
    .A(_0911_),
    .B(_1081_));
 sg13g2_nand3_1 _4913_ (.B(_0911_),
    .C(_1081_),
    .A(net755),
    .Y(_1085_));
 sg13g2_nor2_1 _4914_ (.A(_1078_),
    .B(_1085_),
    .Y(_1086_));
 sg13g2_nand3_1 _4915_ (.B(_2059_),
    .C(_0704_),
    .A(net828),
    .Y(_1087_));
 sg13g2_nand2_2 _4916_ (.Y(_1088_),
    .A(_0557_),
    .B(_0726_));
 sg13g2_nor2_2 _4917_ (.A(_0568_),
    .B(_0616_),
    .Y(_1089_));
 sg13g2_nand2_1 _4918_ (.Y(_1090_),
    .A(_0140_),
    .B(_0722_));
 sg13g2_nand2_1 _4919_ (.Y(_1091_),
    .A(_1089_),
    .B(_1090_));
 sg13g2_o21ai_1 _4920_ (.B1(_1091_),
    .Y(_1092_),
    .A1(_1087_),
    .A2(_1088_));
 sg13g2_nor2_1 _4921_ (.A(net834),
    .B(_1092_),
    .Y(_1093_));
 sg13g2_o21ai_1 _4922_ (.B1(net688),
    .Y(_1095_),
    .A1(_1086_),
    .A2(_1093_));
 sg13g2_o21ai_1 _4923_ (.B1(_0171_),
    .Y(_1096_),
    .A1(_0436_),
    .A2(_0801_));
 sg13g2_nand4_1 _4924_ (.B(_0469_),
    .C(_0612_),
    .A(_0403_),
    .Y(_1097_),
    .D(_0707_));
 sg13g2_nand3_1 _4925_ (.B(_1096_),
    .C(_1097_),
    .A(net828),
    .Y(_1098_));
 sg13g2_nand4_1 _4926_ (.B(_0817_),
    .C(_1095_),
    .A(_0767_),
    .Y(_1099_),
    .D(_1098_));
 sg13g2_nor2_2 _4927_ (.A(net668),
    .B(_0798_),
    .Y(_1100_));
 sg13g2_nor2b_1 _4928_ (.A(_0982_),
    .B_N(_1100_),
    .Y(_1101_));
 sg13g2_nor3_2 _4929_ (.A(net663),
    .B(_0770_),
    .C(net687),
    .Y(_1102_));
 sg13g2_nor2_1 _4930_ (.A(net662),
    .B(_0822_),
    .Y(_1103_));
 sg13g2_nor3_1 _4931_ (.A(net662),
    .B(net742),
    .C(_0822_),
    .Y(_1104_));
 sg13g2_nor3_1 _4932_ (.A(_1101_),
    .B(_1102_),
    .C(_1104_),
    .Y(_1106_));
 sg13g2_a21oi_1 _4933_ (.A1(net746),
    .A2(_1021_),
    .Y(_1107_),
    .B1(_1025_));
 sg13g2_nand2_1 _4934_ (.Y(_1108_),
    .A(_1011_),
    .B(_1023_));
 sg13g2_a221oi_1 _4935_ (.B2(_1035_),
    .C1(_1108_),
    .B1(_1031_),
    .A1(net746),
    .Y(_1109_),
    .A2(_0888_));
 sg13g2_nand4_1 _4936_ (.B(_1040_),
    .C(_1107_),
    .A(_1003_),
    .Y(_1110_),
    .D(_1109_));
 sg13g2_a21oi_1 _4937_ (.A1(_0897_),
    .A2(_0900_),
    .Y(_1111_),
    .B1(_1008_));
 sg13g2_a221oi_1 _4938_ (.B2(_0946_),
    .C1(_1010_),
    .B1(_1020_),
    .A1(_0997_),
    .Y(_1112_),
    .A2(_0998_));
 sg13g2_nand3_1 _4939_ (.B(_1111_),
    .C(_1112_),
    .A(_1014_),
    .Y(_1113_));
 sg13g2_nand3_1 _4940_ (.B(_0917_),
    .C(_1004_),
    .A(net694),
    .Y(_1114_));
 sg13g2_nand4_1 _4941_ (.B(_1019_),
    .C(_1037_),
    .A(_1000_),
    .Y(_1115_),
    .D(_1114_));
 sg13g2_nor4_1 _4942_ (.A(_0906_),
    .B(_1110_),
    .C(_1113_),
    .D(_1115_),
    .Y(_1117_));
 sg13g2_nor3_1 _4943_ (.A(_1101_),
    .B(_1102_),
    .C(_1104_),
    .Y(_1118_));
 sg13g2_nand4_1 _4944_ (.B(_0980_),
    .C(_1117_),
    .A(_0847_),
    .Y(_1119_),
    .D(_1118_));
 sg13g2_a22oi_1 _4945_ (.Y(_1120_),
    .B1(_0961_),
    .B2(_0963_),
    .A2(_0935_),
    .A1(_0934_));
 sg13g2_nor3_1 _4946_ (.A(_0889_),
    .B(_0891_),
    .C(_1016_),
    .Y(_1121_));
 sg13g2_o21ai_1 _4947_ (.B1(net765),
    .Y(_1122_),
    .A1(_0901_),
    .A2(_0902_));
 sg13g2_o21ai_1 _4948_ (.B1(_1122_),
    .Y(_1123_),
    .A1(_0633_),
    .A2(_1121_));
 sg13g2_a21o_1 _4949_ (.A2(_0828_),
    .A1(_0823_),
    .B1(_0784_),
    .X(_1124_));
 sg13g2_a221oi_1 _4950_ (.B2(net728),
    .C1(_1124_),
    .B1(_1123_),
    .A1(_0824_),
    .Y(_1125_),
    .A2(_0921_));
 sg13g2_a22oi_1 _4951_ (.Y(_1126_),
    .B1(_0982_),
    .B2(_0985_),
    .A2(_0930_),
    .A1(_0928_));
 sg13g2_nand3_1 _4952_ (.B(_0958_),
    .C(_1126_),
    .A(_0933_),
    .Y(_1128_));
 sg13g2_nor4_1 _4953_ (.A(_0838_),
    .B(_0872_),
    .C(_0916_),
    .D(_1128_),
    .Y(_1129_));
 sg13g2_nand4_1 _4954_ (.B(_1120_),
    .C(_1125_),
    .A(_1076_),
    .Y(_1130_),
    .D(_1129_));
 sg13g2_nor4_2 _4955_ (.A(_0883_),
    .B(_0975_),
    .C(_1119_),
    .Y(_1131_),
    .D(_1130_));
 sg13g2_nor2_1 _4956_ (.A(_0766_),
    .B(_0942_),
    .Y(_1132_));
 sg13g2_a221oi_1 _4957_ (.B2(_1030_),
    .C1(_0821_),
    .B1(_1029_),
    .A1(_0987_),
    .Y(_1133_),
    .A2(_0994_));
 sg13g2_nor2b_1 _4958_ (.A(_0779_),
    .B_N(_1099_),
    .Y(_1134_));
 sg13g2_nand4_1 _4959_ (.B(_1132_),
    .C(_1133_),
    .A(_1131_),
    .Y(_1135_),
    .D(_1134_));
 sg13g2_nor2_1 _4960_ (.A(net660),
    .B(_0886_),
    .Y(_1136_));
 sg13g2_nor4_1 _4961_ (.A(_0614_),
    .B(_0744_),
    .C(_1069_),
    .D(_1135_),
    .Y(_1137_));
 sg13g2_xnor2_1 _4962_ (.Y(_1139_),
    .A(net801),
    .B(_2865_));
 sg13g2_nor2_1 _4963_ (.A(_0140_),
    .B(_1139_),
    .Y(_1140_));
 sg13g2_nand2_1 _4964_ (.Y(_1141_),
    .A(_0160_),
    .B(_0412_));
 sg13g2_a22oi_1 _4965_ (.Y(_1142_),
    .B1(_0412_),
    .B2(net700),
    .A2(_0374_),
    .A1(_0191_));
 sg13g2_xor2_1 _4966_ (.B(_1139_),
    .A(net844),
    .X(_1143_));
 sg13g2_nand4_1 _4967_ (.B(_0295_),
    .C(_1141_),
    .A(_0192_),
    .Y(_1144_),
    .D(_1143_));
 sg13g2_o21ai_1 _4968_ (.B1(_1144_),
    .Y(_1145_),
    .A1(_1140_),
    .A2(_1142_));
 sg13g2_o21ai_1 _4969_ (.B1(_1145_),
    .Y(_1146_),
    .A1(_0160_),
    .A2(_0412_));
 sg13g2_nor2_1 _4970_ (.A(net810),
    .B(_0732_),
    .Y(_1147_));
 sg13g2_xnor2_1 _4971_ (.Y(_1148_),
    .A(_0015_),
    .B(_1147_));
 sg13g2_nor2_1 _4972_ (.A(_1140_),
    .B(_1143_),
    .Y(_1150_));
 sg13g2_a21oi_1 _4973_ (.A1(net703),
    .A2(_1148_),
    .Y(_1151_),
    .B1(_1150_));
 sg13g2_a21o_1 _4974_ (.A2(_2865_),
    .A1(_1424_),
    .B1(net773),
    .X(_1152_));
 sg13g2_nor3_1 _4975_ (.A(net810),
    .B(_0732_),
    .C(_1446_),
    .Y(_1153_));
 sg13g2_nand2b_1 _4976_ (.Y(_1154_),
    .B(_1152_),
    .A_N(_1153_));
 sg13g2_nor2_1 _4977_ (.A(net703),
    .B(_1148_),
    .Y(_1155_));
 sg13g2_a221oi_1 _4978_ (.B2(_0177_),
    .C1(_1155_),
    .B1(_1154_),
    .A1(_1146_),
    .Y(_1156_),
    .A2(_1151_));
 sg13g2_nand3_1 _4979_ (.B(net782),
    .C(net780),
    .A(net786),
    .Y(_1157_));
 sg13g2_o21ai_1 _4980_ (.B1(net763),
    .Y(_1158_),
    .A1(_0177_),
    .A2(_1153_));
 sg13g2_mux2_1 _4981_ (.A0(_1157_),
    .A1(_1158_),
    .S(_1152_),
    .X(_1159_));
 sg13g2_or2_2 _4982_ (.X(_1161_),
    .B(_1159_),
    .A(_1156_));
 sg13g2_nand2b_1 _4983_ (.Y(_1162_),
    .B(_1161_),
    .A_N(_0225_));
 sg13g2_nand2b_1 _4984_ (.Y(_1163_),
    .B(_0396_),
    .A_N(_0285_));
 sg13g2_nor2_1 _4985_ (.A(_0307_),
    .B(_1163_),
    .Y(_1164_));
 sg13g2_a21o_1 _4986_ (.A2(_1164_),
    .A1(net747),
    .B1(_1162_),
    .X(_1165_));
 sg13g2_nor2_2 _4987_ (.A(net673),
    .B(_0899_),
    .Y(_1166_));
 sg13g2_a22oi_1 _4988_ (.Y(_1167_),
    .B1(_1165_),
    .B2(_1166_),
    .A2(_0398_),
    .A1(_0230_));
 sg13g2_nand3_1 _4989_ (.B(_1137_),
    .C(_1167_),
    .A(_0508_),
    .Y(_1168_));
 sg13g2_nor2b_1 _4990_ (.A(_2593_),
    .B_N(_2653_),
    .Y(_1169_));
 sg13g2_nand2_1 _4991_ (.Y(_1170_),
    .A(_2652_),
    .B(_2820_));
 sg13g2_xnor2_1 _4992_ (.Y(_1172_),
    .A(_1169_),
    .B(_1170_));
 sg13g2_a22oi_1 _4993_ (.Y(_1173_),
    .B1(_1172_),
    .B2(_2838_),
    .A2(_2840_),
    .A1(_2839_));
 sg13g2_or3_1 _4994_ (.A(_2835_),
    .B(_2836_),
    .C(_1173_),
    .X(_1174_));
 sg13g2_a21oi_2 _4995_ (.B1(net784),
    .Y(_1175_),
    .A2(_0220_),
    .A1(_0732_));
 sg13g2_or4_2 _4996_ (.A(net783),
    .B(_0710_),
    .C(net723),
    .D(_0220_),
    .X(_1176_));
 sg13g2_nor4_2 _4997_ (.A(_2835_),
    .B(_2836_),
    .C(_1173_),
    .Y(_1177_),
    .D(_1176_));
 sg13g2_a21oi_2 _4998_ (.B1(_1039_),
    .Y(_1178_),
    .A2(_1177_),
    .A1(_2842_));
 sg13g2_a21oi_1 _4999_ (.A1(net769),
    .A2(_1698_),
    .Y(_1179_),
    .B1(_1088_));
 sg13g2_nor2b_1 _5000_ (.A(_1179_),
    .B_N(_1089_),
    .Y(_1180_));
 sg13g2_nand2_1 _5001_ (.Y(_1181_),
    .A(net769),
    .B(net762));
 sg13g2_o21ai_1 _5002_ (.B1(net830),
    .Y(_1183_),
    .A1(_1088_),
    .A2(_1181_));
 sg13g2_nor2_1 _5003_ (.A(_1180_),
    .B(_1183_),
    .Y(_1184_));
 sg13g2_nor2_1 _5004_ (.A(net760),
    .B(_1184_),
    .Y(_1185_));
 sg13g2_a21oi_1 _5005_ (.A1(net734),
    .A2(_1184_),
    .Y(_1186_),
    .B1(_1185_));
 sg13g2_nor2_1 _5006_ (.A(net731),
    .B(net667),
    .Y(_1187_));
 sg13g2_nand2_2 _5007_ (.Y(_1188_),
    .A(net737),
    .B(_0805_));
 sg13g2_o21ai_1 _5008_ (.B1(_1188_),
    .Y(_1189_),
    .A1(_0805_),
    .A2(_1186_));
 sg13g2_o21ai_1 _5009_ (.B1(_1178_),
    .Y(_1190_),
    .A1(_1177_),
    .A2(_1189_));
 sg13g2_o21ai_1 _5010_ (.B1(_2841_),
    .Y(_1191_),
    .A1(_2835_),
    .A2(_2836_));
 sg13g2_o21ai_1 _5011_ (.B1(net792),
    .Y(_1192_),
    .A1(net798),
    .A2(_0655_));
 sg13g2_a21oi_2 _5012_ (.B1(_2844_),
    .Y(_1194_),
    .A2(_1192_),
    .A1(_1314_));
 sg13g2_nand4_1 _5013_ (.B(_1175_),
    .C(_1191_),
    .A(_1174_),
    .Y(_1195_),
    .D(_1194_));
 sg13g2_nor2_2 _5014_ (.A(net661),
    .B(_0833_),
    .Y(_1196_));
 sg13g2_nand2_1 _5015_ (.Y(_1197_),
    .A(net687),
    .B(_0992_));
 sg13g2_nor2_2 _5016_ (.A(net660),
    .B(_0511_),
    .Y(_1198_));
 sg13g2_a22oi_1 _5017_ (.Y(_1199_),
    .B1(_1197_),
    .B2(_1198_),
    .A2(_1196_),
    .A1(_1195_));
 sg13g2_nor2_2 _5018_ (.A(net756),
    .B(net690),
    .Y(_1200_));
 sg13g2_nand2_2 _5019_ (.Y(_1201_),
    .A(net753),
    .B(net687));
 sg13g2_nor2_1 _5020_ (.A(_0737_),
    .B(net669),
    .Y(_1202_));
 sg13g2_nor3_1 _5021_ (.A(_0737_),
    .B(net669),
    .C(_1201_),
    .Y(_1203_));
 sg13g2_inv_2 _5022_ (.Y(_1205_),
    .A(_1203_));
 sg13g2_nand2_2 _5023_ (.Y(_1206_),
    .A(_0401_),
    .B(_0767_));
 sg13g2_nor2_1 _5024_ (.A(_0732_),
    .B(_0743_),
    .Y(_1207_));
 sg13g2_a21oi_1 _5025_ (.A1(_1402_),
    .A2(_1207_),
    .Y(_1208_),
    .B1(net773));
 sg13g2_o21ai_1 _5026_ (.B1(net688),
    .Y(_1209_),
    .A1(_0013_),
    .A2(_0590_));
 sg13g2_nor2_1 _5027_ (.A(_0305_),
    .B(_0579_),
    .Y(_1210_));
 sg13g2_o21ai_1 _5028_ (.B1(_1209_),
    .Y(_1211_),
    .A1(net688),
    .A2(_1210_));
 sg13g2_xnor2_1 _5029_ (.Y(_1212_),
    .A(net779),
    .B(_1211_));
 sg13g2_xnor2_1 _5030_ (.Y(_1213_),
    .A(net833),
    .B(_1211_));
 sg13g2_xnor2_1 _5031_ (.Y(_1214_),
    .A(_0151_),
    .B(net689));
 sg13g2_xnor2_1 _5032_ (.Y(_1216_),
    .A(_0154_),
    .B(net689));
 sg13g2_xnor2_1 _5033_ (.Y(_1217_),
    .A(net844),
    .B(net689));
 sg13g2_nand3_1 _5034_ (.B(_1216_),
    .C(_1217_),
    .A(_0174_),
    .Y(_1218_));
 sg13g2_xnor2_1 _5035_ (.Y(_1219_),
    .A(net855),
    .B(net689));
 sg13g2_xnor2_1 _5036_ (.Y(_1220_),
    .A(\flag.flag_abrosexual_inst.pix_y[1] ),
    .B(net689));
 sg13g2_xnor2_1 _5037_ (.Y(_1221_),
    .A(net858),
    .B(net689));
 sg13g2_xnor2_1 _5038_ (.Y(_1222_),
    .A(net862),
    .B(net689));
 sg13g2_nor4_1 _5039_ (.A(_1219_),
    .B(_1220_),
    .C(_1221_),
    .D(_1222_),
    .Y(_1223_));
 sg13g2_nor3_1 _5040_ (.A(_1214_),
    .B(_1218_),
    .C(_1223_),
    .Y(_1224_));
 sg13g2_or2_1 _5041_ (.X(_1225_),
    .B(_1224_),
    .A(_1212_));
 sg13g2_o21ai_1 _5042_ (.B1(_1225_),
    .Y(_1227_),
    .A1(net759),
    .A2(_1208_));
 sg13g2_nand2_1 _5043_ (.Y(_1228_),
    .A(net773),
    .B(_0418_));
 sg13g2_nor2_1 _5044_ (.A(_1534_),
    .B(_0441_),
    .Y(_1229_));
 sg13g2_nand4_1 _5045_ (.B(net814),
    .C(net817),
    .A(net824),
    .Y(_1230_),
    .D(net810));
 sg13g2_nand4_1 _5046_ (.B(net804),
    .C(_1523_),
    .A(_0206_),
    .Y(_1231_),
    .D(_1230_));
 sg13g2_o21ai_1 _5047_ (.B1(_0261_),
    .Y(_1232_),
    .A1(_0228_),
    .A2(net801));
 sg13g2_nor2_1 _5048_ (.A(_2861_),
    .B(_0553_),
    .Y(_1233_));
 sg13g2_a221oi_1 _5049_ (.B2(_1229_),
    .C1(net759),
    .B1(_1233_),
    .A1(_1231_),
    .Y(_1234_),
    .A2(_1232_));
 sg13g2_and2_1 _5050_ (.A(_0206_),
    .B(_1230_),
    .X(_1235_));
 sg13g2_nor2_2 _5051_ (.A(_0206_),
    .B(_1230_),
    .Y(_1236_));
 sg13g2_nor2_1 _5052_ (.A(_1235_),
    .B(_1236_),
    .Y(_1238_));
 sg13g2_xnor2_1 _5053_ (.Y(_1239_),
    .A(net808),
    .B(_2872_));
 sg13g2_mux2_2 _5054_ (.A0(_1239_),
    .A1(_1238_),
    .S(_1234_),
    .X(_1240_));
 sg13g2_nand2b_1 _5055_ (.Y(_1241_),
    .B(net811),
    .A_N(net807));
 sg13g2_o21ai_1 _5056_ (.B1(net806),
    .Y(_1242_),
    .A1(_2854_),
    .A2(_1241_));
 sg13g2_xnor2_1 _5057_ (.Y(_1243_),
    .A(net776),
    .B(_1242_));
 sg13g2_xnor2_1 _5058_ (.Y(_1244_),
    .A(net802),
    .B(_1235_));
 sg13g2_mux2_2 _5059_ (.A0(_1243_),
    .A1(_1244_),
    .S(_1234_),
    .X(_1245_));
 sg13g2_nand2_2 _5060_ (.Y(_1246_),
    .A(_1240_),
    .B(_1245_));
 sg13g2_inv_1 _5061_ (.Y(_1247_),
    .A(_1246_));
 sg13g2_and2_1 _5062_ (.A(_0016_),
    .B(_0621_),
    .X(_1249_));
 sg13g2_xnor2_1 _5063_ (.Y(_1250_),
    .A(_0140_),
    .B(_1249_));
 sg13g2_xor2_1 _5064_ (.B(_0377_),
    .A(net845),
    .X(_1251_));
 sg13g2_mux2_1 _5065_ (.A0(_1251_),
    .A1(_1250_),
    .S(_0627_),
    .X(_1252_));
 sg13g2_xnor2_1 _5066_ (.Y(_1253_),
    .A(net844),
    .B(_0376_));
 sg13g2_nor2_1 _5067_ (.A(net752),
    .B(_1253_),
    .Y(_1254_));
 sg13g2_nor2_1 _5068_ (.A(_0016_),
    .B(_0621_),
    .Y(_1255_));
 sg13g2_xnor2_1 _5069_ (.Y(_1256_),
    .A(net847),
    .B(_1255_));
 sg13g2_a22oi_1 _5070_ (.Y(_1257_),
    .B1(_1256_),
    .B2(net752),
    .A2(_1254_),
    .A1(net691));
 sg13g2_o21ai_1 _5071_ (.B1(_1257_),
    .Y(_1258_),
    .A1(net691),
    .A2(_1252_));
 sg13g2_o21ai_1 _5072_ (.B1(_0378_),
    .Y(_1260_),
    .A1(_0622_),
    .A2(_0626_));
 sg13g2_or4_1 _5073_ (.A(_0622_),
    .B(_0626_),
    .C(_1249_),
    .D(_1255_),
    .X(_1261_));
 sg13g2_nand3_1 _5074_ (.B(_1260_),
    .C(_1261_),
    .A(_0856_),
    .Y(_1262_));
 sg13g2_nand2_1 _5075_ (.Y(_1263_),
    .A(_0620_),
    .B(net752));
 sg13g2_xnor2_1 _5076_ (.Y(_1264_),
    .A(_0378_),
    .B(_1263_));
 sg13g2_nand2_2 _5077_ (.Y(_1265_),
    .A(net691),
    .B(_1264_));
 sg13g2_and2_1 _5078_ (.A(_1262_),
    .B(_1265_),
    .X(_1266_));
 sg13g2_nand2_2 _5079_ (.Y(_1267_),
    .A(_1262_),
    .B(_1265_));
 sg13g2_nand2_2 _5080_ (.Y(_1268_),
    .A(_1258_),
    .B(_1266_));
 sg13g2_nor2_2 _5081_ (.A(_1246_),
    .B(_1268_),
    .Y(_1269_));
 sg13g2_nand2_1 _5082_ (.Y(_1271_),
    .A(_1245_),
    .B(_1258_));
 sg13g2_or2_1 _5083_ (.X(_1272_),
    .B(_1258_),
    .A(net685));
 sg13g2_a21oi_1 _5084_ (.A1(_1271_),
    .A2(_1272_),
    .Y(_1273_),
    .B1(_1269_));
 sg13g2_mux2_2 _5085_ (.A0(_2875_),
    .A1(_2877_),
    .S(_1234_),
    .X(_1274_));
 sg13g2_nand2_2 _5086_ (.Y(_1275_),
    .A(net685),
    .B(net684));
 sg13g2_nand2b_1 _5087_ (.Y(_1276_),
    .B(_1240_),
    .A_N(net684));
 sg13g2_nand2_1 _5088_ (.Y(_1277_),
    .A(_1275_),
    .B(_1276_));
 sg13g2_nand2_1 _5089_ (.Y(_1278_),
    .A(_1266_),
    .B(_1277_));
 sg13g2_nand3b_1 _5090_ (.B(net684),
    .C(net686),
    .Y(_1279_),
    .A_N(net685));
 sg13g2_nor2_1 _5091_ (.A(_1246_),
    .B(net683),
    .Y(_1280_));
 sg13g2_xor2_1 _5092_ (.B(_1280_),
    .A(_1268_),
    .X(_1282_));
 sg13g2_a21oi_1 _5093_ (.A1(_1278_),
    .A2(_1279_),
    .Y(_1283_),
    .B1(_1282_));
 sg13g2_a21oi_1 _5094_ (.A1(_1247_),
    .A2(net683),
    .Y(_1284_),
    .B1(_1269_));
 sg13g2_xnor2_1 _5095_ (.Y(_1285_),
    .A(_1283_),
    .B(_1284_));
 sg13g2_nand2b_1 _5096_ (.Y(_1286_),
    .B(_1285_),
    .A_N(_1273_));
 sg13g2_a21oi_1 _5097_ (.A1(_1271_),
    .A2(_1286_),
    .Y(_1287_),
    .B1(_1269_));
 sg13g2_xnor2_1 _5098_ (.Y(_1288_),
    .A(_1273_),
    .B(_1285_));
 sg13g2_nand3_1 _5099_ (.B(_1279_),
    .C(_1282_),
    .A(_1278_),
    .Y(_1289_));
 sg13g2_nand2b_1 _5100_ (.Y(_1290_),
    .B(_1289_),
    .A_N(_1283_));
 sg13g2_a221oi_1 _5101_ (.B2(_0854_),
    .C1(_0622_),
    .B1(_0851_),
    .A1(_0619_),
    .Y(_1291_),
    .A2(_0625_));
 sg13g2_nor2_1 _5102_ (.A(net752),
    .B(_1291_),
    .Y(_1293_));
 sg13g2_or3_1 _5103_ (.A(net852),
    .B(net752),
    .C(_1291_),
    .X(_1294_));
 sg13g2_o21ai_1 _5104_ (.B1(_1294_),
    .Y(_1295_),
    .A1(_0658_),
    .A2(_1293_));
 sg13g2_mux2_2 _5105_ (.A0(_0658_),
    .A1(net852),
    .S(_1293_),
    .X(_1296_));
 sg13g2_nand2_1 _5106_ (.Y(_1297_),
    .A(_1266_),
    .B(_1295_));
 sg13g2_mux2_2 _5107_ (.A0(_2928_),
    .A1(_2926_),
    .S(_1234_),
    .X(_1298_));
 sg13g2_inv_2 _5108_ (.Y(_1299_),
    .A(_1298_));
 sg13g2_o21ai_1 _5109_ (.B1(_1299_),
    .Y(_1300_),
    .A1(net686),
    .A2(net685));
 sg13g2_nor2_1 _5110_ (.A(_1247_),
    .B(_1300_),
    .Y(_1301_));
 sg13g2_inv_1 _5111_ (.Y(_1302_),
    .A(_1301_));
 sg13g2_nand2_1 _5112_ (.Y(_1304_),
    .A(net685),
    .B(_1299_));
 sg13g2_nand3_1 _5113_ (.B(net685),
    .C(_1299_),
    .A(net686),
    .Y(_1305_));
 sg13g2_o21ai_1 _5114_ (.B1(_1305_),
    .Y(_1306_),
    .A1(_1297_),
    .A2(_1302_));
 sg13g2_xnor2_1 _5115_ (.Y(_1307_),
    .A(_1267_),
    .B(_1277_));
 sg13g2_nand2_2 _5116_ (.Y(_1308_),
    .A(_1258_),
    .B(_1295_));
 sg13g2_nand3b_1 _5117_ (.B(_0019_),
    .C(_0945_),
    .Y(_1309_),
    .A_N(_1291_));
 sg13g2_o21ai_1 _5118_ (.B1(_2321_),
    .Y(_1310_),
    .A1(net752),
    .A2(_1291_));
 sg13g2_nand2_2 _5119_ (.Y(_1311_),
    .A(_1309_),
    .B(_1310_));
 sg13g2_nor2_1 _5120_ (.A(_1267_),
    .B(_1311_),
    .Y(_1312_));
 sg13g2_nand4_1 _5121_ (.B(_1265_),
    .C(_1309_),
    .A(_1262_),
    .Y(_1313_),
    .D(_1310_));
 sg13g2_xnor2_1 _5122_ (.Y(_1315_),
    .A(_1306_),
    .B(_1307_));
 sg13g2_nor3_1 _5123_ (.A(_1308_),
    .B(_1312_),
    .C(_1315_),
    .Y(_1316_));
 sg13g2_a21oi_1 _5124_ (.A1(_1306_),
    .A2(_1307_),
    .Y(_1317_),
    .B1(_1316_));
 sg13g2_or2_1 _5125_ (.X(_1318_),
    .B(_1317_),
    .A(_1290_));
 sg13g2_nor2_1 _5126_ (.A(_1275_),
    .B(_1308_),
    .Y(_1319_));
 sg13g2_nor2_2 _5127_ (.A(_1296_),
    .B(_1311_),
    .Y(_1320_));
 sg13g2_inv_1 _5128_ (.Y(_1321_),
    .A(_1320_));
 sg13g2_nor2_1 _5129_ (.A(_1268_),
    .B(_1320_),
    .Y(_1322_));
 sg13g2_xnor2_1 _5130_ (.Y(_1323_),
    .A(_1247_),
    .B(_1322_));
 sg13g2_nor2b_1 _5131_ (.A(_1323_),
    .B_N(_1319_),
    .Y(_1324_));
 sg13g2_xor2_1 _5132_ (.B(_1323_),
    .A(_1319_),
    .X(_1326_));
 sg13g2_xnor2_1 _5133_ (.Y(_1327_),
    .A(_1290_),
    .B(_1317_));
 sg13g2_o21ai_1 _5134_ (.B1(_1318_),
    .Y(_1328_),
    .A1(_1326_),
    .A2(_1327_));
 sg13g2_nor2_1 _5135_ (.A(_1308_),
    .B(_1313_),
    .Y(_1329_));
 sg13g2_a21oi_1 _5136_ (.A1(_1246_),
    .A2(_1329_),
    .Y(_1330_),
    .B1(_1324_));
 sg13g2_xor2_1 _5137_ (.B(_1328_),
    .A(_1288_),
    .X(_1331_));
 sg13g2_nor2b_1 _5138_ (.A(_1330_),
    .B_N(_1331_),
    .Y(_1332_));
 sg13g2_a21o_1 _5139_ (.A2(_1328_),
    .A1(_1288_),
    .B1(_1332_),
    .X(_1333_));
 sg13g2_xnor2_1 _5140_ (.Y(_1334_),
    .A(_1287_),
    .B(_1333_));
 sg13g2_mux2_2 _5141_ (.A0(net818),
    .A1(_1939_),
    .S(_1234_),
    .X(_1335_));
 sg13g2_mux2_2 _5142_ (.A0(_0195_),
    .A1(_1950_),
    .S(_1234_),
    .X(_1337_));
 sg13g2_nand2_2 _5143_ (.Y(_1338_),
    .A(net685),
    .B(_1337_));
 sg13g2_nor2_1 _5144_ (.A(_1313_),
    .B(_1338_),
    .Y(_1339_));
 sg13g2_xor2_1 _5145_ (.B(_1338_),
    .A(_1313_),
    .X(_1340_));
 sg13g2_o21ai_1 _5146_ (.B1(net683),
    .Y(_1341_),
    .A1(_1299_),
    .A2(_1340_));
 sg13g2_xnor2_1 _5147_ (.Y(_1342_),
    .A(_1297_),
    .B(_1301_));
 sg13g2_inv_1 _5148_ (.Y(_1343_),
    .A(_1342_));
 sg13g2_o21ai_1 _5149_ (.B1(_2069_),
    .Y(_1344_),
    .A1(net752),
    .A2(_1291_));
 sg13g2_nand3b_1 _5150_ (.B(_0022_),
    .C(_0945_),
    .Y(_1345_),
    .A_N(_1291_));
 sg13g2_nand2_2 _5151_ (.Y(_1346_),
    .A(_1344_),
    .B(_1345_));
 sg13g2_and2_2 _5152_ (.A(_1344_),
    .B(_1345_),
    .X(_1348_));
 sg13g2_nand2_2 _5153_ (.Y(_1349_),
    .A(_1258_),
    .B(_1348_));
 sg13g2_xnor2_1 _5154_ (.Y(_1350_),
    .A(_1295_),
    .B(_1313_));
 sg13g2_nand2b_1 _5155_ (.Y(_1351_),
    .B(_1350_),
    .A_N(_1349_));
 sg13g2_o21ai_1 _5156_ (.B1(_1351_),
    .Y(_1352_),
    .A1(_1296_),
    .A2(_1313_));
 sg13g2_nand2b_1 _5157_ (.Y(_1353_),
    .B(_1258_),
    .A_N(_1311_));
 sg13g2_a21oi_1 _5158_ (.A1(_1297_),
    .A2(_1353_),
    .Y(_1354_),
    .B1(_1329_));
 sg13g2_and2_1 _5159_ (.A(_1339_),
    .B(_1354_),
    .X(_1355_));
 sg13g2_xor2_1 _5160_ (.B(_1354_),
    .A(_1339_),
    .X(_1356_));
 sg13g2_xnor2_1 _5161_ (.Y(_1357_),
    .A(_1352_),
    .B(_1356_));
 sg13g2_xnor2_1 _5162_ (.Y(_1359_),
    .A(_1341_),
    .B(_1342_));
 sg13g2_nand2b_1 _5163_ (.Y(_1360_),
    .B(_1359_),
    .A_N(_1357_));
 sg13g2_o21ai_1 _5164_ (.B1(_1360_),
    .Y(_1361_),
    .A1(_1341_),
    .A2(_1343_));
 sg13g2_o21ai_1 _5165_ (.B1(_1315_),
    .Y(_1362_),
    .A1(_1308_),
    .A2(_1312_));
 sg13g2_nor2b_1 _5166_ (.A(_1316_),
    .B_N(_1362_),
    .Y(_1363_));
 sg13g2_and2_1 _5167_ (.A(_1361_),
    .B(_1363_),
    .X(_1364_));
 sg13g2_or2_1 _5168_ (.X(_1365_),
    .B(_1353_),
    .A(_1304_));
 sg13g2_a21oi_1 _5169_ (.A1(_1352_),
    .A2(_1356_),
    .Y(_1366_),
    .B1(_1355_));
 sg13g2_xor2_1 _5170_ (.B(_1308_),
    .A(_1275_),
    .X(_1367_));
 sg13g2_nand2b_1 _5171_ (.Y(_1368_),
    .B(_1367_),
    .A_N(_1366_));
 sg13g2_xor2_1 _5172_ (.B(_1367_),
    .A(_1366_),
    .X(_1370_));
 sg13g2_xor2_1 _5173_ (.B(_1370_),
    .A(_1365_),
    .X(_1371_));
 sg13g2_xor2_1 _5174_ (.B(_1363_),
    .A(_1361_),
    .X(_1372_));
 sg13g2_a21oi_1 _5175_ (.A1(_1371_),
    .A2(_1372_),
    .Y(_1373_),
    .B1(_1364_));
 sg13g2_xor2_1 _5176_ (.B(_1327_),
    .A(_1326_),
    .X(_1374_));
 sg13g2_nor2b_1 _5177_ (.A(_1373_),
    .B_N(_1374_),
    .Y(_1375_));
 sg13g2_o21ai_1 _5178_ (.B1(_1368_),
    .Y(_1376_),
    .A1(_1365_),
    .A2(_1370_));
 sg13g2_xnor2_1 _5179_ (.Y(_1377_),
    .A(_1373_),
    .B(_1374_));
 sg13g2_a21oi_1 _5180_ (.A1(_1376_),
    .A2(_1377_),
    .Y(_1378_),
    .B1(_1375_));
 sg13g2_xnor2_1 _5181_ (.Y(_1379_),
    .A(_1330_),
    .B(_1331_));
 sg13g2_nor2b_1 _5182_ (.A(_1378_),
    .B_N(_1379_),
    .Y(_1381_));
 sg13g2_and2_1 _5183_ (.A(net686),
    .B(_1337_),
    .X(_1382_));
 sg13g2_nand2_1 _5184_ (.Y(_1383_),
    .A(net827),
    .B(net686));
 sg13g2_and4_1 _5185_ (.A(net826),
    .B(net686),
    .C(net683),
    .D(_1337_),
    .X(_1384_));
 sg13g2_nand4_1 _5186_ (.B(net686),
    .C(net683),
    .A(net826),
    .Y(_1385_),
    .D(_1337_));
 sg13g2_a22oi_1 _5187_ (.Y(_1386_),
    .B1(net683),
    .B2(_1337_),
    .A2(net686),
    .A1(net826));
 sg13g2_nor2_1 _5188_ (.A(_1384_),
    .B(_1386_),
    .Y(_1387_));
 sg13g2_or3_1 _5189_ (.A(_1298_),
    .B(_1384_),
    .C(_1386_),
    .X(_1388_));
 sg13g2_o21ai_1 _5190_ (.B1(_1385_),
    .Y(_1389_),
    .A1(_1298_),
    .A2(_1386_));
 sg13g2_nand2_1 _5191_ (.Y(_1390_),
    .A(_1382_),
    .B(_1389_));
 sg13g2_xnor2_1 _5192_ (.Y(_1392_),
    .A(_1382_),
    .B(_1389_));
 sg13g2_nor2_2 _5193_ (.A(_1267_),
    .B(_1346_),
    .Y(_1393_));
 sg13g2_nand4_1 _5194_ (.B(_1265_),
    .C(_1344_),
    .A(_1262_),
    .Y(_1394_),
    .D(_1345_));
 sg13g2_nand2_2 _5195_ (.Y(_1395_),
    .A(net826),
    .B(net685));
 sg13g2_or2_1 _5196_ (.X(_1396_),
    .B(_1383_),
    .A(_1338_));
 sg13g2_xor2_1 _5197_ (.B(_1395_),
    .A(_1382_),
    .X(_1397_));
 sg13g2_xnor2_1 _5198_ (.Y(_1398_),
    .A(_1394_),
    .B(_1397_));
 sg13g2_o21ai_1 _5199_ (.B1(_1390_),
    .Y(_1399_),
    .A1(_1392_),
    .A2(_1398_));
 sg13g2_inv_1 _5200_ (.Y(_1400_),
    .A(_1399_));
 sg13g2_nand2_1 _5201_ (.Y(_1401_),
    .A(net684),
    .B(_1298_));
 sg13g2_xor2_1 _5202_ (.B(_1401_),
    .A(_1340_),
    .X(_1403_));
 sg13g2_nor2_1 _5203_ (.A(_1400_),
    .B(_1403_),
    .Y(_1404_));
 sg13g2_xnor2_1 _5204_ (.Y(_1405_),
    .A(_1399_),
    .B(_1403_));
 sg13g2_o21ai_1 _5205_ (.B1(_1396_),
    .Y(_1406_),
    .A1(_1394_),
    .A2(_1397_));
 sg13g2_xnor2_1 _5206_ (.Y(_1407_),
    .A(_1349_),
    .B(_1350_));
 sg13g2_nand2_1 _5207_ (.Y(_1408_),
    .A(_1406_),
    .B(_1407_));
 sg13g2_xnor2_1 _5208_ (.Y(_1409_),
    .A(_1406_),
    .B(_1407_));
 sg13g2_xnor2_1 _5209_ (.Y(_1410_),
    .A(_1320_),
    .B(_1409_));
 sg13g2_a21oi_1 _5210_ (.A1(_1405_),
    .A2(_1410_),
    .Y(_1411_),
    .B1(_1404_));
 sg13g2_xnor2_1 _5211_ (.Y(_1412_),
    .A(_1357_),
    .B(_1359_));
 sg13g2_nor2b_1 _5212_ (.A(_1411_),
    .B_N(_1412_),
    .Y(_1414_));
 sg13g2_o21ai_1 _5213_ (.B1(_1408_),
    .Y(_1415_),
    .A1(_1321_),
    .A2(_1409_));
 sg13g2_xor2_1 _5214_ (.B(_1353_),
    .A(_1304_),
    .X(_1416_));
 sg13g2_xnor2_1 _5215_ (.Y(_1417_),
    .A(_1415_),
    .B(_1416_));
 sg13g2_nor3_1 _5216_ (.A(_1338_),
    .B(_1349_),
    .C(_1417_),
    .Y(_1418_));
 sg13g2_o21ai_1 _5217_ (.B1(_1417_),
    .Y(_1419_),
    .A1(_1338_),
    .A2(_1349_));
 sg13g2_nor2b_1 _5218_ (.A(_1418_),
    .B_N(_1419_),
    .Y(_1420_));
 sg13g2_xnor2_1 _5219_ (.Y(_1421_),
    .A(_1411_),
    .B(_1412_));
 sg13g2_a21oi_1 _5220_ (.A1(_1420_),
    .A2(_1421_),
    .Y(_1422_),
    .B1(_1414_));
 sg13g2_xnor2_1 _5221_ (.Y(_1423_),
    .A(_1371_),
    .B(_1372_));
 sg13g2_nor2_1 _5222_ (.A(_1422_),
    .B(_1423_),
    .Y(_1425_));
 sg13g2_a21o_1 _5223_ (.A2(_1416_),
    .A1(_1415_),
    .B1(_1418_),
    .X(_1426_));
 sg13g2_xor2_1 _5224_ (.B(_1423_),
    .A(_1422_),
    .X(_1427_));
 sg13g2_a21oi_1 _5225_ (.A1(_1426_),
    .A2(_1427_),
    .Y(_1428_),
    .B1(_1425_));
 sg13g2_xnor2_1 _5226_ (.Y(_1429_),
    .A(_1376_),
    .B(_1377_));
 sg13g2_or2_1 _5227_ (.X(_1430_),
    .B(_1429_),
    .A(_1428_));
 sg13g2_nor3_2 _5228_ (.A(net821),
    .B(_1298_),
    .C(_1335_),
    .Y(_1431_));
 sg13g2_and2_2 _5229_ (.A(net683),
    .B(_1431_),
    .X(_1432_));
 sg13g2_inv_1 _5230_ (.Y(_1433_),
    .A(_1432_));
 sg13g2_nor2b_1 _5231_ (.A(_1383_),
    .B_N(_1432_),
    .Y(_1434_));
 sg13g2_nand2b_1 _5232_ (.Y(_1436_),
    .B(_1432_),
    .A_N(_1383_));
 sg13g2_o21ai_1 _5233_ (.B1(_1298_),
    .Y(_1437_),
    .A1(_1384_),
    .A2(_1386_));
 sg13g2_a21oi_1 _5234_ (.A1(_1388_),
    .A2(_1437_),
    .Y(_1438_),
    .B1(_1432_));
 sg13g2_nand3_1 _5235_ (.B(_1262_),
    .C(_1265_),
    .A(net864),
    .Y(_1439_));
 sg13g2_xor2_1 _5236_ (.B(_1439_),
    .A(_1387_),
    .X(_1440_));
 sg13g2_or3_1 _5237_ (.A(_1434_),
    .B(_1438_),
    .C(_1440_),
    .X(_1441_));
 sg13g2_o21ai_1 _5238_ (.B1(_1436_),
    .Y(_1442_),
    .A1(_1438_),
    .A2(_1440_));
 sg13g2_xor2_1 _5239_ (.B(_1398_),
    .A(_1392_),
    .X(_1443_));
 sg13g2_xnor2_1 _5240_ (.Y(_1444_),
    .A(_1442_),
    .B(_1443_));
 sg13g2_nand2_1 _5241_ (.Y(_1445_),
    .A(_1295_),
    .B(_1348_));
 sg13g2_o21ai_1 _5242_ (.B1(_1385_),
    .Y(_1447_),
    .A1(_1386_),
    .A2(_1439_));
 sg13g2_xnor2_1 _5243_ (.Y(_1448_),
    .A(_1393_),
    .B(_1447_));
 sg13g2_nor2_1 _5244_ (.A(_1445_),
    .B(_1448_),
    .Y(_1449_));
 sg13g2_xnor2_1 _5245_ (.Y(_1450_),
    .A(_1445_),
    .B(_1448_));
 sg13g2_nor2_1 _5246_ (.A(_1444_),
    .B(_1450_),
    .Y(_1451_));
 sg13g2_a21oi_1 _5247_ (.A1(_1442_),
    .A2(_1443_),
    .Y(_1452_),
    .B1(_1451_));
 sg13g2_xnor2_1 _5248_ (.Y(_1453_),
    .A(_1405_),
    .B(_1410_));
 sg13g2_or2_1 _5249_ (.X(_1454_),
    .B(_1453_),
    .A(_1452_));
 sg13g2_xnor2_1 _5250_ (.Y(_1455_),
    .A(_1452_),
    .B(_1453_));
 sg13g2_nand2_1 _5251_ (.Y(_1456_),
    .A(net864),
    .B(_1258_));
 sg13g2_inv_1 _5252_ (.Y(_1458_),
    .A(_1456_));
 sg13g2_a21oi_2 _5253_ (.B1(_1449_),
    .Y(_1459_),
    .A2(_1447_),
    .A1(_1393_));
 sg13g2_xnor2_1 _5254_ (.Y(_1460_),
    .A(_1338_),
    .B(_1349_));
 sg13g2_nor2_1 _5255_ (.A(_1459_),
    .B(_1460_),
    .Y(_1461_));
 sg13g2_xor2_1 _5256_ (.B(_1460_),
    .A(_1459_),
    .X(_1462_));
 sg13g2_xnor2_1 _5257_ (.Y(_1463_),
    .A(_1458_),
    .B(_1462_));
 sg13g2_o21ai_1 _5258_ (.B1(_1454_),
    .Y(_1464_),
    .A1(_1455_),
    .A2(_1463_));
 sg13g2_xnor2_1 _5259_ (.Y(_1465_),
    .A(_1420_),
    .B(_1421_));
 sg13g2_nor2b_1 _5260_ (.A(_1465_),
    .B_N(_1464_),
    .Y(_1466_));
 sg13g2_a21oi_1 _5261_ (.A1(_1458_),
    .A2(_1462_),
    .Y(_1467_),
    .B1(_1461_));
 sg13g2_xor2_1 _5262_ (.B(_1465_),
    .A(_1464_),
    .X(_1469_));
 sg13g2_nor2_1 _5263_ (.A(_1467_),
    .B(_1469_),
    .Y(_1470_));
 sg13g2_nor2_1 _5264_ (.A(_1466_),
    .B(_1470_),
    .Y(_1471_));
 sg13g2_xnor2_1 _5265_ (.Y(_1472_),
    .A(_1426_),
    .B(_1427_));
 sg13g2_nor2_1 _5266_ (.A(_1471_),
    .B(_1472_),
    .Y(_1473_));
 sg13g2_a22oi_1 _5267_ (.Y(_1474_),
    .B1(_1299_),
    .B2(_1337_),
    .A2(net683),
    .A1(_0349_));
 sg13g2_nor2_1 _5268_ (.A(_1432_),
    .B(_1474_),
    .Y(_1475_));
 sg13g2_o21ai_1 _5269_ (.B1(_1440_),
    .Y(_1476_),
    .A1(_1434_),
    .A2(_1438_));
 sg13g2_nand3_1 _5270_ (.B(_1475_),
    .C(_1476_),
    .A(_1441_),
    .Y(_1477_));
 sg13g2_a21oi_1 _5271_ (.A1(_1441_),
    .A2(_1476_),
    .Y(_1478_),
    .B1(_1475_));
 sg13g2_a21o_1 _5272_ (.A2(_1476_),
    .A1(_1441_),
    .B1(_1475_),
    .X(_1480_));
 sg13g2_nor2_1 _5273_ (.A(_1311_),
    .B(_1348_),
    .Y(_1481_));
 sg13g2_xnor2_1 _5274_ (.Y(_1482_),
    .A(_1432_),
    .B(_1481_));
 sg13g2_inv_1 _5275_ (.Y(_1483_),
    .A(_1482_));
 sg13g2_and3_1 _5276_ (.X(_1484_),
    .A(_1477_),
    .B(_1480_),
    .C(_1483_));
 sg13g2_o21ai_1 _5277_ (.B1(_1477_),
    .Y(_1485_),
    .A1(_1478_),
    .A2(_1482_));
 sg13g2_xor2_1 _5278_ (.B(_1450_),
    .A(_1444_),
    .X(_1486_));
 sg13g2_nand2_1 _5279_ (.Y(_1487_),
    .A(_1485_),
    .B(_1486_));
 sg13g2_a21oi_2 _5280_ (.B1(_1311_),
    .Y(_1488_),
    .A2(_1433_),
    .A1(_1346_));
 sg13g2_inv_1 _5281_ (.Y(_1489_),
    .A(_1488_));
 sg13g2_nor2_1 _5282_ (.A(_1395_),
    .B(_1489_),
    .Y(_1491_));
 sg13g2_xor2_1 _5283_ (.B(_1488_),
    .A(_1395_),
    .X(_1492_));
 sg13g2_xnor2_1 _5284_ (.Y(_1493_),
    .A(_1485_),
    .B(_1486_));
 sg13g2_o21ai_1 _5285_ (.B1(_1487_),
    .Y(_1494_),
    .A1(_1492_),
    .A2(_1493_));
 sg13g2_xor2_1 _5286_ (.B(_1463_),
    .A(_1455_),
    .X(_1495_));
 sg13g2_xnor2_1 _5287_ (.Y(_1496_),
    .A(_1494_),
    .B(_1495_));
 sg13g2_nor3_1 _5288_ (.A(_1395_),
    .B(_1489_),
    .C(_1496_),
    .Y(_1497_));
 sg13g2_a21oi_1 _5289_ (.A1(_1494_),
    .A2(_1495_),
    .Y(_1498_),
    .B1(_1497_));
 sg13g2_xor2_1 _5290_ (.B(_1469_),
    .A(_1467_),
    .X(_1499_));
 sg13g2_nand2b_1 _5291_ (.Y(_1500_),
    .B(_1499_),
    .A_N(_1498_));
 sg13g2_xor2_1 _5292_ (.B(_1499_),
    .A(_1498_),
    .X(_1502_));
 sg13g2_nor3_1 _5293_ (.A(net821),
    .B(_1298_),
    .C(_1337_),
    .Y(_1503_));
 sg13g2_nand3_1 _5294_ (.B(_1309_),
    .C(_1310_),
    .A(_0063_),
    .Y(_1504_));
 sg13g2_nor2_2 _5295_ (.A(_1346_),
    .B(_1504_),
    .Y(_1505_));
 sg13g2_inv_1 _5296_ (.Y(_1506_),
    .A(_1505_));
 sg13g2_nor2_1 _5297_ (.A(_0025_),
    .B(_1296_),
    .Y(_1507_));
 sg13g2_nand2_1 _5298_ (.Y(_1508_),
    .A(_1431_),
    .B(_1507_));
 sg13g2_xnor2_1 _5299_ (.Y(_1509_),
    .A(_1431_),
    .B(_1507_));
 sg13g2_xnor2_1 _5300_ (.Y(_1510_),
    .A(_1505_),
    .B(_1509_));
 sg13g2_nand2_1 _5301_ (.Y(_1511_),
    .A(_1503_),
    .B(_1510_));
 sg13g2_a21oi_1 _5302_ (.A1(_1477_),
    .A2(_1480_),
    .Y(_1513_),
    .B1(_1483_));
 sg13g2_nor3_1 _5303_ (.A(_1484_),
    .B(_1511_),
    .C(_1513_),
    .Y(_1514_));
 sg13g2_or3_1 _5304_ (.A(_1484_),
    .B(_1511_),
    .C(_1513_),
    .X(_1515_));
 sg13g2_o21ai_1 _5305_ (.B1(_1508_),
    .Y(_1516_),
    .A1(_1506_),
    .A2(_1509_));
 sg13g2_nand2b_1 _5306_ (.Y(_1517_),
    .B(_1516_),
    .A_N(_1439_));
 sg13g2_xnor2_1 _5307_ (.Y(_1518_),
    .A(_1439_),
    .B(_1516_));
 sg13g2_o21ai_1 _5308_ (.B1(_1511_),
    .Y(_1519_),
    .A1(_1484_),
    .A2(_1513_));
 sg13g2_and3_1 _5309_ (.X(_1520_),
    .A(_1515_),
    .B(_1518_),
    .C(_1519_));
 sg13g2_a21oi_1 _5310_ (.A1(_1518_),
    .A2(_1519_),
    .Y(_1521_),
    .B1(_1514_));
 sg13g2_xnor2_1 _5311_ (.Y(_1522_),
    .A(_1492_),
    .B(_1493_));
 sg13g2_xor2_1 _5312_ (.B(_1522_),
    .A(_1521_),
    .X(_1524_));
 sg13g2_nand2b_1 _5313_ (.Y(_1525_),
    .B(_1524_),
    .A_N(_1517_));
 sg13g2_o21ai_1 _5314_ (.B1(_1525_),
    .Y(_1526_),
    .A1(_1521_),
    .A2(_1522_));
 sg13g2_xor2_1 _5315_ (.B(_1496_),
    .A(_1491_),
    .X(_1527_));
 sg13g2_nor2b_1 _5316_ (.A(_1527_),
    .B_N(_1526_),
    .Y(_1528_));
 sg13g2_nand2b_1 _5317_ (.Y(_1529_),
    .B(_1526_),
    .A_N(_1527_));
 sg13g2_xnor2_1 _5318_ (.Y(_1530_),
    .A(_1348_),
    .B(_1504_));
 sg13g2_nand2_1 _5319_ (.Y(_1531_),
    .A(net826),
    .B(_1530_));
 sg13g2_o21ai_1 _5320_ (.B1(_1337_),
    .Y(_1532_),
    .A1(net826),
    .A2(_1530_));
 sg13g2_nor2b_1 _5321_ (.A(_1532_),
    .B_N(_1531_),
    .Y(_1533_));
 sg13g2_nor2_1 _5322_ (.A(_1335_),
    .B(_1531_),
    .Y(_1535_));
 sg13g2_nand2_1 _5323_ (.Y(_1536_),
    .A(net863),
    .B(_1295_));
 sg13g2_nor3_2 _5324_ (.A(_1335_),
    .B(_1531_),
    .C(_1536_),
    .Y(_1537_));
 sg13g2_xnor2_1 _5325_ (.Y(_1538_),
    .A(_1535_),
    .B(_1536_));
 sg13g2_nor2_1 _5326_ (.A(_1503_),
    .B(_1533_),
    .Y(_1539_));
 sg13g2_xnor2_1 _5327_ (.Y(_1540_),
    .A(_1510_),
    .B(_1539_));
 sg13g2_a22oi_1 _5328_ (.Y(_1541_),
    .B1(_1538_),
    .B2(_1540_),
    .A2(_1533_),
    .A1(_1510_));
 sg13g2_a21oi_1 _5329_ (.A1(_1515_),
    .A2(_1519_),
    .Y(_1542_),
    .B1(_1518_));
 sg13g2_nor3_1 _5330_ (.A(_1520_),
    .B(_1541_),
    .C(_1542_),
    .Y(_1543_));
 sg13g2_or3_1 _5331_ (.A(_1520_),
    .B(_1541_),
    .C(_1542_),
    .X(_1544_));
 sg13g2_o21ai_1 _5332_ (.B1(_1541_),
    .Y(_1546_),
    .A1(_1520_),
    .A2(_1542_));
 sg13g2_and3_1 _5333_ (.X(_1547_),
    .A(_1537_),
    .B(_1544_),
    .C(_1546_));
 sg13g2_a21oi_1 _5334_ (.A1(_1537_),
    .A2(_1546_),
    .Y(_1548_),
    .B1(_1543_));
 sg13g2_xnor2_1 _5335_ (.Y(_1549_),
    .A(_1517_),
    .B(_1524_));
 sg13g2_nand2b_1 _5336_ (.Y(_1550_),
    .B(_1549_),
    .A_N(_1548_));
 sg13g2_xor2_1 _5337_ (.B(_1549_),
    .A(_1548_),
    .X(_1551_));
 sg13g2_a21oi_1 _5338_ (.A1(_1544_),
    .A2(_1546_),
    .Y(_1552_),
    .B1(_1537_));
 sg13g2_nor2_1 _5339_ (.A(_1538_),
    .B(_1540_),
    .Y(_1553_));
 sg13g2_nand2_1 _5340_ (.Y(_1554_),
    .A(net863),
    .B(_1348_));
 sg13g2_a221oi_1 _5341_ (.B2(_1504_),
    .C1(_1533_),
    .B1(_1554_),
    .A1(_1335_),
    .Y(_1555_),
    .A2(_1505_));
 sg13g2_a21oi_1 _5342_ (.A1(net863),
    .A2(_1505_),
    .Y(_1557_),
    .B1(_1555_));
 sg13g2_a21o_1 _5343_ (.A2(_1540_),
    .A1(_1538_),
    .B1(_1557_),
    .X(_1558_));
 sg13g2_or4_1 _5344_ (.A(_1547_),
    .B(_1552_),
    .C(_1553_),
    .D(_1558_),
    .X(_1559_));
 sg13g2_o21ai_1 _5345_ (.B1(_1550_),
    .Y(_1560_),
    .A1(_1551_),
    .A2(_1559_));
 sg13g2_nand2b_1 _5346_ (.Y(_1561_),
    .B(_1527_),
    .A_N(_1526_));
 sg13g2_a21oi_1 _5347_ (.A1(_1560_),
    .A2(_1561_),
    .Y(_1562_),
    .B1(_1528_));
 sg13g2_o21ai_1 _5348_ (.B1(_1500_),
    .Y(_1563_),
    .A1(_1502_),
    .A2(_1562_));
 sg13g2_xor2_1 _5349_ (.B(_1472_),
    .A(_1471_),
    .X(_1564_));
 sg13g2_a21oi_1 _5350_ (.A1(_1563_),
    .A2(_1564_),
    .Y(_1565_),
    .B1(_1473_));
 sg13g2_xnor2_1 _5351_ (.Y(_1566_),
    .A(_1428_),
    .B(_1429_));
 sg13g2_o21ai_1 _5352_ (.B1(_1430_),
    .Y(_1568_),
    .A1(_1565_),
    .A2(_1566_));
 sg13g2_xnor2_1 _5353_ (.Y(_1569_),
    .A(_1378_),
    .B(_1379_));
 sg13g2_a21oi_1 _5354_ (.A1(_1568_),
    .A2(_1569_),
    .Y(_1570_),
    .B1(_1381_));
 sg13g2_a21oi_1 _5355_ (.A1(_1287_),
    .A2(_1333_),
    .Y(_1571_),
    .B1(_1269_));
 sg13g2_o21ai_1 _5356_ (.B1(_1571_),
    .Y(_1572_),
    .A1(_1334_),
    .A2(_1570_));
 sg13g2_xnor2_1 _5357_ (.Y(_1573_),
    .A(_1568_),
    .B(_1569_));
 sg13g2_xor2_1 _5358_ (.B(_1566_),
    .A(_1565_),
    .X(_1574_));
 sg13g2_xnor2_1 _5359_ (.Y(_1575_),
    .A(_1502_),
    .B(_1562_));
 sg13g2_a21oi_1 _5360_ (.A1(_1529_),
    .A2(_1561_),
    .Y(_1576_),
    .B1(_1560_));
 sg13g2_xnor2_1 _5361_ (.Y(_1577_),
    .A(_1551_),
    .B(_1559_));
 sg13g2_o21ai_1 _5362_ (.B1(_1575_),
    .Y(_1579_),
    .A1(_1576_),
    .A2(_1577_));
 sg13g2_xor2_1 _5363_ (.B(_1564_),
    .A(_1563_),
    .X(_1580_));
 sg13g2_a21oi_2 _5364_ (.B1(_1574_),
    .Y(_1581_),
    .A2(_1580_),
    .A1(_1579_));
 sg13g2_a22oi_1 _5365_ (.Y(_1582_),
    .B1(_1573_),
    .B2(_1581_),
    .A2(_1570_),
    .A1(_1334_));
 sg13g2_o21ai_1 _5366_ (.B1(_1227_),
    .Y(_1583_),
    .A1(_1572_),
    .A2(_1582_));
 sg13g2_o21ai_1 _5367_ (.B1(net801),
    .Y(_1584_),
    .A1(_0442_),
    .A2(_0553_));
 sg13g2_nor2_2 _5368_ (.A(net800),
    .B(_1584_),
    .Y(_1585_));
 sg13g2_nor2_2 _5369_ (.A(_0219_),
    .B(_1585_),
    .Y(_1586_));
 sg13g2_o21ai_1 _5370_ (.B1(net775),
    .Y(_1587_),
    .A1(net773),
    .A2(_1585_));
 sg13g2_nor2b_1 _5371_ (.A(_1586_),
    .B_N(_1587_),
    .Y(_1588_));
 sg13g2_nor2_1 _5372_ (.A(net806),
    .B(_0553_),
    .Y(_1590_));
 sg13g2_xnor2_1 _5373_ (.Y(_1591_),
    .A(net776),
    .B(_1590_));
 sg13g2_or2_1 _5374_ (.X(_1592_),
    .B(_1591_),
    .A(_1217_));
 sg13g2_xnor2_1 _5375_ (.Y(_1593_),
    .A(net796),
    .B(_1584_));
 sg13g2_o21ai_1 _5376_ (.B1(_1592_),
    .Y(_1594_),
    .A1(_1216_),
    .A2(_1593_));
 sg13g2_xnor2_1 _5377_ (.Y(_1595_),
    .A(_0316_),
    .B(_0553_));
 sg13g2_nor2_1 _5378_ (.A(_1214_),
    .B(_1595_),
    .Y(_1596_));
 sg13g2_nor2_1 _5379_ (.A(_0181_),
    .B(_1219_),
    .Y(_1597_));
 sg13g2_a21oi_1 _5380_ (.A1(_1214_),
    .A2(_1595_),
    .Y(_1598_),
    .B1(_1597_));
 sg13g2_a22oi_1 _5381_ (.Y(_1599_),
    .B1(_1221_),
    .B2(net816),
    .A2(_1219_),
    .A1(_0181_));
 sg13g2_xnor2_1 _5382_ (.Y(_1601_),
    .A(net771),
    .B(_1222_));
 sg13g2_nor2_1 _5383_ (.A(_0023_),
    .B(_1220_),
    .Y(_1602_));
 sg13g2_or2_1 _5384_ (.X(_1603_),
    .B(_1220_),
    .A(_0023_));
 sg13g2_nand2_1 _5385_ (.Y(_1604_),
    .A(_0023_),
    .B(_1220_));
 sg13g2_nand3_1 _5386_ (.B(_1603_),
    .C(_1604_),
    .A(_1601_),
    .Y(_1605_));
 sg13g2_xnor2_1 _5387_ (.Y(_1606_),
    .A(_0272_),
    .B(_1586_));
 sg13g2_nor2_1 _5388_ (.A(_1605_),
    .B(_1606_),
    .Y(_1607_));
 sg13g2_nor2_1 _5389_ (.A(_0107_),
    .B(_1222_),
    .Y(_1608_));
 sg13g2_a21oi_1 _5390_ (.A1(_1604_),
    .A2(_1608_),
    .Y(_1609_),
    .B1(_1602_));
 sg13g2_o21ai_1 _5391_ (.B1(_1609_),
    .Y(_1610_),
    .A1(net816),
    .A2(_1221_));
 sg13g2_o21ai_1 _5392_ (.B1(_1599_),
    .Y(_1612_),
    .A1(_1607_),
    .A2(_1610_));
 sg13g2_a221oi_1 _5393_ (.B2(_1612_),
    .C1(_1596_),
    .B1(_1598_),
    .A1(_1217_),
    .Y(_1613_),
    .A2(_1591_));
 sg13g2_xnor2_1 _5394_ (.Y(_1614_),
    .A(net773),
    .B(_1585_));
 sg13g2_a22oi_1 _5395_ (.Y(_1615_),
    .B1(_1614_),
    .B2(_0174_),
    .A2(_1593_),
    .A1(_1216_));
 sg13g2_o21ai_1 _5396_ (.B1(_1615_),
    .Y(_1616_),
    .A1(_1594_),
    .A2(_1613_));
 sg13g2_nor2_1 _5397_ (.A(_0174_),
    .B(_1614_),
    .Y(_1617_));
 sg13g2_a21oi_1 _5398_ (.A1(_1213_),
    .A2(_1588_),
    .Y(_1618_),
    .B1(_1617_));
 sg13g2_nand2_1 _5399_ (.Y(_1619_),
    .A(_1616_),
    .B(_1618_));
 sg13g2_o21ai_1 _5400_ (.B1(_1619_),
    .Y(_1620_),
    .A1(_1213_),
    .A2(_1588_));
 sg13g2_nor2_1 _5401_ (.A(_0666_),
    .B(_0553_),
    .Y(_1621_));
 sg13g2_nor3_1 _5402_ (.A(net786),
    .B(_1446_),
    .C(_1621_),
    .Y(_1623_));
 sg13g2_a21oi_1 _5403_ (.A1(_0378_),
    .A2(_1223_),
    .Y(_1624_),
    .B1(_1218_));
 sg13g2_nor2_1 _5404_ (.A(_1212_),
    .B(_1624_),
    .Y(_1625_));
 sg13g2_nor4_1 _5405_ (.A(net784),
    .B(_1586_),
    .C(_1623_),
    .D(_1625_),
    .Y(_1626_));
 sg13g2_nand3_1 _5406_ (.B(_1620_),
    .C(_1626_),
    .A(_1583_),
    .Y(_1627_));
 sg13g2_xnor2_1 _5407_ (.Y(_1628_),
    .A(net785),
    .B(_1213_));
 sg13g2_nand2_1 _5408_ (.Y(_1629_),
    .A(net781),
    .B(_1628_));
 sg13g2_xnor2_1 _5409_ (.Y(_1630_),
    .A(net773),
    .B(_0172_));
 sg13g2_o21ai_1 _5410_ (.B1(_1630_),
    .Y(_1631_),
    .A1(net796),
    .A2(_1216_));
 sg13g2_a21oi_1 _5411_ (.A1(net796),
    .A2(_1216_),
    .Y(_1632_),
    .B1(_1631_));
 sg13g2_and2_1 _5412_ (.A(net777),
    .B(_1217_),
    .X(_1634_));
 sg13g2_and2_1 _5413_ (.A(net813),
    .B(_1221_),
    .X(_1635_));
 sg13g2_nor2_1 _5414_ (.A(_1609_),
    .B(_1635_),
    .Y(_1636_));
 sg13g2_xnor2_1 _5415_ (.Y(_1637_),
    .A(net809),
    .B(_1219_));
 sg13g2_nor2_1 _5416_ (.A(net813),
    .B(_1221_),
    .Y(_1638_));
 sg13g2_nor3_1 _5417_ (.A(_1636_),
    .B(_1637_),
    .C(_1638_),
    .Y(_1639_));
 sg13g2_nor2_1 _5418_ (.A(_0316_),
    .B(_1214_),
    .Y(_1640_));
 sg13g2_a21oi_1 _5419_ (.A1(_0217_),
    .A2(_1219_),
    .Y(_1641_),
    .B1(_1640_));
 sg13g2_nor2b_1 _5420_ (.A(_1639_),
    .B_N(_1641_),
    .Y(_1642_));
 sg13g2_and2_1 _5421_ (.A(_0316_),
    .B(_1214_),
    .X(_1643_));
 sg13g2_xnor2_1 _5422_ (.Y(_1645_),
    .A(net802),
    .B(_1217_));
 sg13g2_nor3_1 _5423_ (.A(_1642_),
    .B(_1643_),
    .C(_1645_),
    .Y(_1646_));
 sg13g2_o21ai_1 _5424_ (.B1(_1632_),
    .Y(_1647_),
    .A1(_1634_),
    .A2(_1646_));
 sg13g2_a21oi_1 _5425_ (.A1(net790),
    .A2(_0172_),
    .Y(_1648_),
    .B1(net800));
 sg13g2_a22oi_1 _5426_ (.Y(_1649_),
    .B1(_1216_),
    .B2(_1648_),
    .A2(_0174_),
    .A1(net773));
 sg13g2_a21oi_1 _5427_ (.A1(_1647_),
    .A2(_1649_),
    .Y(_1650_),
    .B1(_1629_));
 sg13g2_a21oi_1 _5428_ (.A1(net763),
    .A2(_1212_),
    .Y(_1651_),
    .B1(_1650_));
 sg13g2_or4_1 _5429_ (.A(_1635_),
    .B(_1638_),
    .C(_1640_),
    .D(_1643_),
    .X(_1652_));
 sg13g2_nor3_1 _5430_ (.A(_1637_),
    .B(_1645_),
    .C(_1652_),
    .Y(_1653_));
 sg13g2_nor2b_1 _5431_ (.A(_1605_),
    .B_N(_1632_),
    .Y(_1654_));
 sg13g2_nand4_1 _5432_ (.B(_1628_),
    .C(_1653_),
    .A(net781),
    .Y(_1656_),
    .D(_1654_));
 sg13g2_nor2b_2 _5433_ (.A(_1651_),
    .B_N(_1656_),
    .Y(_1657_));
 sg13g2_nor2_1 _5434_ (.A(_1200_),
    .B(_1657_),
    .Y(_1658_));
 sg13g2_a21o_1 _5435_ (.A2(_1658_),
    .A1(_1627_),
    .B1(_1206_),
    .X(_1659_));
 sg13g2_a221oi_1 _5436_ (.B2(_1198_),
    .C1(_1168_),
    .B1(_1197_),
    .A1(_1195_),
    .Y(_1660_),
    .A2(_1196_));
 sg13g2_and4_1 _5437_ (.A(_1190_),
    .B(_1205_),
    .C(_1659_),
    .D(_1660_),
    .X(_1661_));
 sg13g2_a21oi_2 _5438_ (.B1(_1193_),
    .Y(uo_out[4]),
    .A2(_1661_),
    .A1(_2853_));
 sg13g2_nand2_1 _5439_ (.Y(_1662_),
    .A(_0616_),
    .B(_0630_));
 sg13g2_nand3_1 _5440_ (.B(_0616_),
    .C(_0630_),
    .A(_1709_),
    .Y(_1663_));
 sg13g2_nand2_1 _5441_ (.Y(_1664_),
    .A(net835),
    .B(_1663_));
 sg13g2_o21ai_1 _5442_ (.B1(_0806_),
    .Y(_1666_),
    .A1(_1184_),
    .A2(_1664_));
 sg13g2_nand2b_1 _5443_ (.Y(_1667_),
    .B(_1666_),
    .A_N(_1177_));
 sg13g2_or4_1 _5444_ (.A(net739),
    .B(_1177_),
    .C(_1180_),
    .D(_1183_),
    .X(_1668_));
 sg13g2_nand3_1 _5445_ (.B(_1667_),
    .C(_1668_),
    .A(_1178_),
    .Y(_1669_));
 sg13g2_a21oi_1 _5446_ (.A1(_0396_),
    .A2(_0858_),
    .Y(_1670_),
    .B1(_0285_));
 sg13g2_nor2_1 _5447_ (.A(_0307_),
    .B(_1670_),
    .Y(_1671_));
 sg13g2_o21ai_1 _5448_ (.B1(_1166_),
    .Y(_1672_),
    .A1(_1162_),
    .A2(_1671_));
 sg13g2_nand2b_1 _5449_ (.Y(_1673_),
    .B(_0635_),
    .A_N(_0627_));
 sg13g2_or2_1 _5450_ (.X(_1674_),
    .B(_0629_),
    .A(_0628_));
 sg13g2_nor2_1 _5451_ (.A(net749),
    .B(_0642_),
    .Y(_1675_));
 sg13g2_nor2_2 _5452_ (.A(net751),
    .B(_0953_),
    .Y(_1677_));
 sg13g2_nor2b_1 _5453_ (.A(_0738_),
    .B_N(net657),
    .Y(_1678_));
 sg13g2_a21oi_1 _5454_ (.A1(net742),
    .A2(_1675_),
    .Y(_1679_),
    .B1(_1678_));
 sg13g2_nand2b_1 _5455_ (.Y(_1680_),
    .B(_1679_),
    .A_N(_0703_));
 sg13g2_a21oi_1 _5456_ (.A1(_1673_),
    .A2(_1674_),
    .Y(_1681_),
    .B1(_1680_));
 sg13g2_o21ai_1 _5457_ (.B1(net688),
    .Y(_1682_),
    .A1(_1078_),
    .A2(_1085_));
 sg13g2_a21o_1 _5458_ (.A2(_1087_),
    .A1(_0722_),
    .B1(_1753_),
    .X(_1683_));
 sg13g2_nand3_1 _5459_ (.B(_0630_),
    .C(_1683_),
    .A(net779),
    .Y(_1684_));
 sg13g2_nand3_1 _5460_ (.B(_0817_),
    .C(_1684_),
    .A(_0767_),
    .Y(_1685_));
 sg13g2_a21oi_1 _5461_ (.A1(_1098_),
    .A2(_1682_),
    .Y(_1686_),
    .B1(_1685_));
 sg13g2_nand2_1 _5462_ (.Y(_1688_),
    .A(_0957_),
    .B(_1034_));
 sg13g2_and2_1 _5463_ (.A(net759),
    .B(_1059_),
    .X(_1689_));
 sg13g2_nand2_1 _5464_ (.Y(_1690_),
    .A(net759),
    .B(_1059_));
 sg13g2_nand2_2 _5465_ (.Y(_1691_),
    .A(_0924_),
    .B(_1689_));
 sg13g2_inv_1 _5466_ (.Y(_1692_),
    .A(_1691_));
 sg13g2_a21oi_1 _5467_ (.A1(net658),
    .A2(_0917_),
    .Y(_1693_),
    .B1(_1038_));
 sg13g2_nand2_1 _5468_ (.Y(_1694_),
    .A(_0512_),
    .B(net657));
 sg13g2_nand2b_2 _5469_ (.Y(_1695_),
    .B(_0976_),
    .A_N(_0820_));
 sg13g2_nand2_1 _5470_ (.Y(_1696_),
    .A(_1694_),
    .B(_1695_));
 sg13g2_nand2_1 _5471_ (.Y(_1697_),
    .A(_0735_),
    .B(_0834_));
 sg13g2_nand2_1 _5472_ (.Y(_1699_),
    .A(net693),
    .B(_0795_));
 sg13g2_nand2_1 _5473_ (.Y(_1700_),
    .A(_0791_),
    .B(_1699_));
 sg13g2_o21ai_1 _5474_ (.B1(_0799_),
    .Y(_1701_),
    .A1(net740),
    .A2(_1700_));
 sg13g2_a22oi_1 _5475_ (.Y(_1702_),
    .B1(_1697_),
    .B2(_0839_),
    .A2(net657),
    .A1(_0512_));
 sg13g2_and2_1 _5476_ (.A(_1695_),
    .B(_1701_),
    .X(_1703_));
 sg13g2_o21ai_1 _5477_ (.B1(_0773_),
    .Y(_1704_),
    .A1(net729),
    .A2(_0759_));
 sg13g2_a21oi_1 _5478_ (.A1(_0759_),
    .A2(_0775_),
    .Y(_1705_),
    .B1(_1704_));
 sg13g2_a21oi_1 _5479_ (.A1(net695),
    .A2(_1705_),
    .Y(_1706_),
    .B1(_0772_));
 sg13g2_nand2_2 _5480_ (.Y(_1707_),
    .A(_0764_),
    .B(_0903_));
 sg13g2_nor4_1 _5481_ (.A(net662),
    .B(_0235_),
    .C(net699),
    .D(_0831_),
    .Y(_1708_));
 sg13g2_nand2_1 _5482_ (.Y(_1710_),
    .A(net769),
    .B(_1742_));
 sg13g2_nand3_1 _5483_ (.B(_0630_),
    .C(_1710_),
    .A(net830),
    .Y(_1711_));
 sg13g2_nand2_1 _5484_ (.Y(_1712_),
    .A(_1007_),
    .B(_1711_));
 sg13g2_nand3_1 _5485_ (.B(_0736_),
    .C(_1005_),
    .A(_0231_),
    .Y(_1713_));
 sg13g2_nor2b_1 _5486_ (.A(_1709_),
    .B_N(_0788_),
    .Y(_1714_));
 sg13g2_nand2_1 _5487_ (.Y(_1715_),
    .A(net768),
    .B(_1764_));
 sg13g2_o21ai_1 _5488_ (.B1(_0948_),
    .Y(_1716_),
    .A1(_1714_),
    .A2(_1715_));
 sg13g2_a22oi_1 _5489_ (.Y(_1717_),
    .B1(_1716_),
    .B2(_1005_),
    .A2(_1713_),
    .A1(_1712_));
 sg13g2_nor2_2 _5490_ (.A(net668),
    .B(_0866_),
    .Y(_1718_));
 sg13g2_nand2_2 _5491_ (.Y(_1719_),
    .A(_0402_),
    .B(_0736_));
 sg13g2_nand2_1 _5492_ (.Y(_1721_),
    .A(net753),
    .B(_0867_));
 sg13g2_nand3_1 _5493_ (.B(_0631_),
    .C(_0868_),
    .A(net834),
    .Y(_1722_));
 sg13g2_nand2b_1 _5494_ (.Y(_1723_),
    .B(_1303_),
    .A_N(_1336_));
 sg13g2_nand2_2 _5495_ (.Y(_1724_),
    .A(_0996_),
    .B(_1011_));
 sg13g2_o21ai_1 _5496_ (.B1(_0967_),
    .Y(_1725_),
    .A1(_0971_),
    .A2(_1018_));
 sg13g2_nor3_1 _5497_ (.A(_0823_),
    .B(_0845_),
    .C(_1066_),
    .Y(_1726_));
 sg13g2_nor2_1 _5498_ (.A(_0840_),
    .B(_1726_),
    .Y(_1727_));
 sg13g2_nand3_1 _5499_ (.B(_0399_),
    .C(net671),
    .A(_0233_),
    .Y(_1728_));
 sg13g2_nor2_1 _5500_ (.A(_0900_),
    .B(_1024_),
    .Y(_1729_));
 sg13g2_a21oi_1 _5501_ (.A1(_1728_),
    .A2(_1729_),
    .Y(_1730_),
    .B1(_0964_));
 sg13g2_nor2_1 _5502_ (.A(_0892_),
    .B(_0986_),
    .Y(_1732_));
 sg13g2_nand2_1 _5503_ (.Y(_1733_),
    .A(net666),
    .B(_0935_));
 sg13g2_o21ai_1 _5504_ (.B1(_0873_),
    .Y(_1734_),
    .A1(net690),
    .A2(_0880_));
 sg13g2_and2_1 _5505_ (.A(net666),
    .B(_0902_),
    .X(_1735_));
 sg13g2_and2_1 _5506_ (.A(_1020_),
    .B(_1034_),
    .X(_1736_));
 sg13g2_nand2_1 _5507_ (.Y(_1737_),
    .A(_0888_),
    .B(_0954_));
 sg13g2_o21ai_1 _5508_ (.B1(_0858_),
    .Y(_1738_),
    .A1(_0848_),
    .A2(_1021_));
 sg13g2_nand2_1 _5509_ (.Y(_1739_),
    .A(net764),
    .B(net733));
 sg13g2_nor2_1 _5510_ (.A(net764),
    .B(net726),
    .Y(_1740_));
 sg13g2_nand2_1 _5511_ (.Y(_1741_),
    .A(net728),
    .B(_0904_));
 sg13g2_and2_2 _5512_ (.A(net696),
    .B(_0762_),
    .X(_1743_));
 sg13g2_and2_1 _5513_ (.A(_0844_),
    .B(_1743_),
    .X(_1744_));
 sg13g2_nand2_1 _5514_ (.Y(_1745_),
    .A(_0987_),
    .B(_0988_));
 sg13g2_nor3_1 _5515_ (.A(net662),
    .B(_0833_),
    .C(_0994_),
    .Y(_1746_));
 sg13g2_or3_1 _5516_ (.A(net699),
    .B(_0760_),
    .C(_0919_),
    .X(_1747_));
 sg13g2_a221oi_1 _5517_ (.B2(_0930_),
    .C1(_1727_),
    .B1(_1691_),
    .A1(_0816_),
    .Y(_1748_),
    .A2(_1100_));
 sg13g2_o21ai_1 _5518_ (.B1(_0976_),
    .Y(_1749_),
    .A1(_0889_),
    .A2(_0902_));
 sg13g2_nand4_1 _5519_ (.B(_1734_),
    .C(_1748_),
    .A(_1688_),
    .Y(_1750_),
    .D(_1749_));
 sg13g2_nor2_1 _5520_ (.A(_1686_),
    .B(_1750_),
    .Y(_1751_));
 sg13g2_a221oi_1 _5521_ (.B2(net694),
    .C1(_1732_),
    .B1(_1075_),
    .A1(_0892_),
    .Y(_1752_),
    .A2(_1016_));
 sg13g2_a21oi_1 _5522_ (.A1(_0633_),
    .A2(_1739_),
    .Y(_1754_),
    .B1(net726));
 sg13g2_a22oi_1 _5523_ (.Y(_1755_),
    .B1(_1754_),
    .B2(_0891_),
    .A2(_0901_),
    .A1(_0892_));
 sg13g2_a22oi_1 _5524_ (.Y(_1756_),
    .B1(_1103_),
    .B2(_0954_),
    .A2(_1036_),
    .A1(_0897_));
 sg13g2_nand4_1 _5525_ (.B(_1752_),
    .C(_1755_),
    .A(_0980_),
    .Y(_1757_),
    .D(_1756_));
 sg13g2_a221oi_1 _5526_ (.B2(_0950_),
    .C1(_1102_),
    .B1(_1736_),
    .A1(_0954_),
    .Y(_1758_),
    .A2(_1136_));
 sg13g2_nand2_1 _5527_ (.Y(_1759_),
    .A(_0780_),
    .B(_1719_));
 sg13g2_nor3_1 _5528_ (.A(_0914_),
    .B(_1718_),
    .C(_1759_),
    .Y(_1760_));
 sg13g2_nand4_1 _5529_ (.B(_1738_),
    .C(_1758_),
    .A(_0915_),
    .Y(_1761_),
    .D(_1760_));
 sg13g2_a221oi_1 _5530_ (.B2(_1034_),
    .C1(_1724_),
    .B1(_1031_),
    .A1(net753),
    .Y(_1762_),
    .A2(_0867_));
 sg13g2_o21ai_1 _5531_ (.B1(_1723_),
    .Y(_1763_),
    .A1(_1105_),
    .A2(net746));
 sg13g2_a221oi_1 _5532_ (.B2(net753),
    .C1(_1763_),
    .B1(_1198_),
    .A1(net766),
    .Y(_1765_),
    .A2(_1030_));
 sg13g2_nand2b_1 _5533_ (.Y(_1766_),
    .B(_1722_),
    .A_N(_1010_));
 sg13g2_nor4_1 _5534_ (.A(_0932_),
    .B(_1015_),
    .C(_1196_),
    .D(_1766_),
    .Y(_1767_));
 sg13g2_nand4_1 _5535_ (.B(_1762_),
    .C(_1765_),
    .A(_1003_),
    .Y(_1768_),
    .D(_1767_));
 sg13g2_a22oi_1 _5536_ (.Y(_1769_),
    .B1(_0959_),
    .B2(net658),
    .A2(_0935_),
    .A1(net667));
 sg13g2_a21oi_1 _5537_ (.A1(_0999_),
    .A2(_1741_),
    .Y(_1770_),
    .B1(_1717_));
 sg13g2_o21ai_1 _5538_ (.B1(_1725_),
    .Y(_1771_),
    .A1(_0825_),
    .A2(_0938_));
 sg13g2_a221oi_1 _5539_ (.B2(_0835_),
    .C1(_1771_),
    .B1(_1707_),
    .A1(_1022_),
    .Y(_1772_),
    .A2(_1201_));
 sg13g2_nor4_1 _5540_ (.A(net754),
    .B(_0908_),
    .C(_1078_),
    .D(_1082_),
    .Y(_1773_));
 sg13g2_nor4_1 _5541_ (.A(_1708_),
    .B(_1730_),
    .C(_1746_),
    .D(_1773_),
    .Y(_1774_));
 sg13g2_nand4_1 _5542_ (.B(_1770_),
    .C(_1772_),
    .A(_1769_),
    .Y(_1776_),
    .D(_1774_));
 sg13g2_nor4_2 _5543_ (.A(_1757_),
    .B(_1761_),
    .C(_1768_),
    .Y(_1777_),
    .D(_1776_));
 sg13g2_nand3_1 _5544_ (.B(_1703_),
    .C(_1747_),
    .A(_1702_),
    .Y(_1778_));
 sg13g2_nor4_2 _5545_ (.A(_1693_),
    .B(_1706_),
    .C(_1744_),
    .Y(_1779_),
    .D(_1778_));
 sg13g2_nand4_1 _5546_ (.B(_1751_),
    .C(_1777_),
    .A(_1681_),
    .Y(_1780_),
    .D(_1779_));
 sg13g2_nand3_1 _5547_ (.B(_0396_),
    .C(_0858_),
    .A(_0335_),
    .Y(_1781_));
 sg13g2_nand2b_1 _5548_ (.Y(_1782_),
    .B(_0396_),
    .A_N(_0365_));
 sg13g2_nand3_1 _5549_ (.B(_1781_),
    .C(_1782_),
    .A(_0309_),
    .Y(_1783_));
 sg13g2_a221oi_1 _5550_ (.B2(_0236_),
    .C1(_1780_),
    .B1(_1783_),
    .A1(_0405_),
    .Y(_1784_),
    .A2(_0507_));
 sg13g2_and4_1 _5551_ (.A(_1205_),
    .B(_1659_),
    .C(_1672_),
    .D(_1784_),
    .X(_1785_));
 sg13g2_a21oi_2 _5552_ (.B1(_1193_),
    .Y(uo_out[0]),
    .A2(_1785_),
    .A1(_1669_));
 sg13g2_nand2_1 _5553_ (.Y(_1787_),
    .A(_1479_),
    .B(net737));
 sg13g2_a21oi_1 _5554_ (.A1(_2837_),
    .A2(_2850_),
    .Y(_1788_),
    .B1(_1479_));
 sg13g2_nand2_1 _5555_ (.Y(_1789_),
    .A(_1325_),
    .B(_2849_));
 sg13g2_a22oi_1 _5556_ (.Y(_1790_),
    .B1(_1788_),
    .B2(_1789_),
    .A2(net737),
    .A1(_1479_));
 sg13g2_nor3_2 _5557_ (.A(net792),
    .B(net759),
    .C(net736),
    .Y(_1791_));
 sg13g2_nor3_1 _5558_ (.A(_1259_),
    .B(net665),
    .C(_1791_),
    .Y(_1792_));
 sg13g2_o21ai_1 _5559_ (.B1(_1792_),
    .Y(_1793_),
    .A1(_1336_),
    .A2(_1790_));
 sg13g2_o21ai_1 _5560_ (.B1(_1178_),
    .Y(_1794_),
    .A1(net760),
    .A2(_1667_));
 sg13g2_nor2b_1 _5561_ (.A(_1206_),
    .B_N(_1657_),
    .Y(_1795_));
 sg13g2_nor2_1 _5562_ (.A(net743),
    .B(net689),
    .Y(_1797_));
 sg13g2_a21oi_1 _5563_ (.A1(_0396_),
    .A2(_1797_),
    .Y(_1798_),
    .B1(_0285_));
 sg13g2_o21ai_1 _5564_ (.B1(_1161_),
    .Y(_1799_),
    .A1(_0308_),
    .A2(_1798_));
 sg13g2_nand2_1 _5565_ (.Y(_1800_),
    .A(_1166_),
    .B(_1799_));
 sg13g2_nor2_1 _5566_ (.A(_0496_),
    .B(_0506_),
    .Y(_1801_));
 sg13g2_nor2_1 _5567_ (.A(_0501_),
    .B(_0503_),
    .Y(_1802_));
 sg13g2_nand2_1 _5568_ (.Y(_1803_),
    .A(_0500_),
    .B(_1802_));
 sg13g2_a21oi_1 _5569_ (.A1(_1801_),
    .A2(_1803_),
    .Y(_1804_),
    .B1(_0494_));
 sg13g2_o21ai_1 _5570_ (.B1(_0497_),
    .Y(_1805_),
    .A1(_0499_),
    .A2(_1802_));
 sg13g2_nand2_1 _5571_ (.Y(_1806_),
    .A(_0489_),
    .B(_1801_));
 sg13g2_nor2_1 _5572_ (.A(_0493_),
    .B(_1806_),
    .Y(_1808_));
 sg13g2_a21oi_2 _5573_ (.B1(_1804_),
    .Y(_1809_),
    .A2(_1808_),
    .A1(_1805_));
 sg13g2_nand2_1 _5574_ (.Y(_1810_),
    .A(_0405_),
    .B(_1809_));
 sg13g2_a21oi_1 _5575_ (.A1(_1380_),
    .A2(_1457_),
    .Y(_1811_),
    .B1(net759));
 sg13g2_a22oi_1 _5576_ (.Y(_1812_),
    .B1(_0553_),
    .B2(_1049_),
    .A2(_0410_),
    .A1(_1457_));
 sg13g2_a221oi_1 _5577_ (.B2(_1042_),
    .C1(_2863_),
    .B1(_0556_),
    .A1(net774),
    .Y(_1813_),
    .A2(_0272_));
 sg13g2_nand3_1 _5578_ (.B(_2858_),
    .C(_1042_),
    .A(_1347_),
    .Y(_1814_));
 sg13g2_nand2b_1 _5579_ (.Y(_1815_),
    .B(_1814_),
    .A_N(_1813_));
 sg13g2_o21ai_1 _5580_ (.B1(_1229_),
    .Y(_1816_),
    .A1(_0217_),
    .A2(_1380_));
 sg13g2_nand3_1 _5581_ (.B(_1232_),
    .C(_1816_),
    .A(net759),
    .Y(_1817_));
 sg13g2_nand3_1 _5582_ (.B(_0180_),
    .C(_1229_),
    .A(_1347_),
    .Y(_1819_));
 sg13g2_nand3_1 _5583_ (.B(_1817_),
    .C(_1819_),
    .A(_1815_),
    .Y(_1820_));
 sg13g2_o21ai_1 _5584_ (.B1(_1820_),
    .Y(_1821_),
    .A1(_1811_),
    .A2(_1812_));
 sg13g2_nand2_1 _5585_ (.Y(_1822_),
    .A(_0469_),
    .B(_1709_));
 sg13g2_nand4_1 _5586_ (.B(_0612_),
    .C(_1709_),
    .A(_0469_),
    .Y(_1823_),
    .D(_0630_));
 sg13g2_nand4_1 _5587_ (.B(_0612_),
    .C(_1709_),
    .A(_0425_),
    .Y(_1824_),
    .D(_0630_));
 sg13g2_a21oi_1 _5588_ (.A1(_0633_),
    .A2(_1824_),
    .Y(_1825_),
    .B1(_0627_));
 sg13g2_nand4_1 _5589_ (.B(_1821_),
    .C(_1823_),
    .A(_0424_),
    .Y(_1826_),
    .D(_1825_));
 sg13g2_o21ai_1 _5590_ (.B1(net763),
    .Y(_1827_),
    .A1(_0688_),
    .A2(_1048_));
 sg13g2_nor3_1 _5591_ (.A(net772),
    .B(_1088_),
    .C(_1822_),
    .Y(_1828_));
 sg13g2_o21ai_1 _5592_ (.B1(_1089_),
    .Y(_1830_),
    .A1(_0757_),
    .A2(_1088_));
 sg13g2_nand3_1 _5593_ (.B(_2860_),
    .C(_1207_),
    .A(_2858_),
    .Y(_1831_));
 sg13g2_nand4_1 _5594_ (.B(_0272_),
    .C(_1830_),
    .A(net779),
    .Y(_1832_),
    .D(_1831_));
 sg13g2_a21oi_1 _5595_ (.A1(_2856_),
    .A2(_1207_),
    .Y(_1833_),
    .B1(_0219_));
 sg13g2_nor4_2 _5596_ (.A(net863),
    .B(_0118_),
    .C(_1764_),
    .Y(_1834_),
    .D(_0751_));
 sg13g2_or2_2 _5597_ (.X(_1835_),
    .B(_1710_),
    .A(_0425_));
 sg13g2_o21ai_1 _5598_ (.B1(net768),
    .Y(_1836_),
    .A1(_0129_),
    .A2(_1835_));
 sg13g2_o21ai_1 _5599_ (.B1(_1827_),
    .Y(_1837_),
    .A1(_1834_),
    .A2(_1836_));
 sg13g2_or4_1 _5600_ (.A(_1828_),
    .B(_1832_),
    .C(_1833_),
    .D(_1837_),
    .X(_1838_));
 sg13g2_a21oi_2 _5601_ (.B1(_1205_),
    .Y(_1839_),
    .A2(_1838_),
    .A1(_1826_));
 sg13g2_a22oi_1 _5602_ (.Y(_1841_),
    .B1(_0901_),
    .B2(_0931_),
    .A2(_0889_),
    .A1(net666));
 sg13g2_nor2_1 _5603_ (.A(_0964_),
    .B(_1841_),
    .Y(_1842_));
 sg13g2_a21oi_1 _5604_ (.A1(_0761_),
    .A2(_0939_),
    .Y(_1843_),
    .B1(_0960_));
 sg13g2_nor2_1 _5605_ (.A(net730),
    .B(_0829_),
    .Y(_1844_));
 sg13g2_a221oi_1 _5606_ (.B2(_0724_),
    .C1(net740),
    .B1(_1070_),
    .A1(net735),
    .Y(_1845_),
    .A2(_0829_));
 sg13g2_nor4_1 _5607_ (.A(net668),
    .B(_0833_),
    .C(_0941_),
    .D(_1845_),
    .Y(_1846_));
 sg13g2_nor3_1 _5608_ (.A(_1842_),
    .B(_1843_),
    .C(_1846_),
    .Y(_1847_));
 sg13g2_o21ai_1 _5609_ (.B1(_0911_),
    .Y(_1848_),
    .A1(net754),
    .A2(_1081_));
 sg13g2_nand2_2 _5610_ (.Y(_1849_),
    .A(net737),
    .B(net754));
 sg13g2_nor2_2 _5611_ (.A(net692),
    .B(_1849_),
    .Y(_1850_));
 sg13g2_a21oi_1 _5612_ (.A1(net688),
    .A2(_1848_),
    .Y(_1852_),
    .B1(_1850_));
 sg13g2_a21o_1 _5613_ (.A2(_1852_),
    .A1(_1098_),
    .B1(_1685_),
    .X(_1853_));
 sg13g2_o21ai_1 _5614_ (.B1(_0827_),
    .Y(_1854_),
    .A1(_0731_),
    .A2(net730));
 sg13g2_nand2b_1 _5615_ (.Y(_1855_),
    .B(_1854_),
    .A_N(_0780_));
 sg13g2_nand2_2 _5616_ (.Y(_1856_),
    .A(_0809_),
    .B(_0812_));
 sg13g2_inv_1 _5617_ (.Y(_1857_),
    .A(_1856_));
 sg13g2_nand2_1 _5618_ (.Y(_1858_),
    .A(_0968_),
    .B(_1024_));
 sg13g2_nand2_1 _5619_ (.Y(_1859_),
    .A(_1733_),
    .B(_1858_));
 sg13g2_a21oi_1 _5620_ (.A1(_0714_),
    .A2(net755),
    .Y(_1860_),
    .B1(net690));
 sg13g2_nand2b_1 _5621_ (.Y(_1861_),
    .B(_0873_),
    .A_N(_1860_));
 sg13g2_a21oi_1 _5622_ (.A1(_0715_),
    .A2(net732),
    .Y(_1863_),
    .B1(net753));
 sg13g2_o21ai_1 _5623_ (.B1(_1861_),
    .Y(_1864_),
    .A1(_1745_),
    .A2(_1863_));
 sg13g2_a22oi_1 _5624_ (.Y(_1865_),
    .B1(_1864_),
    .B2(_0991_),
    .A2(_1859_),
    .A1(_1856_));
 sg13g2_nand4_1 _5625_ (.B(_1853_),
    .C(_1855_),
    .A(_1847_),
    .Y(_1866_),
    .D(_1865_));
 sg13g2_o21ai_1 _5626_ (.B1(_0020_),
    .Y(_1867_),
    .A1(_1347_),
    .A2(_2859_));
 sg13g2_nand2_1 _5627_ (.Y(_1868_),
    .A(_1042_),
    .B(_1867_));
 sg13g2_nand4_1 _5628_ (.B(_0014_),
    .C(_1228_),
    .A(net774),
    .Y(_1869_),
    .D(_1868_));
 sg13g2_nor2b_1 _5629_ (.A(_0125_),
    .B_N(_1869_),
    .Y(_1870_));
 sg13g2_a21oi_1 _5630_ (.A1(net783),
    .A2(_1870_),
    .Y(_1871_),
    .B1(_0745_));
 sg13g2_o21ai_1 _5631_ (.B1(net806),
    .Y(_1872_),
    .A1(_1369_),
    .A2(_1241_));
 sg13g2_nand2_1 _5632_ (.Y(_1874_),
    .A(net796),
    .B(_1138_));
 sg13g2_a21oi_1 _5633_ (.A1(_0407_),
    .A2(_1872_),
    .Y(_1875_),
    .B1(_1874_));
 sg13g2_nor4_1 _5634_ (.A(net780),
    .B(_1690_),
    .C(_1871_),
    .D(_1875_),
    .Y(_1876_));
 sg13g2_nor3_1 _5635_ (.A(net787),
    .B(_0125_),
    .C(_1059_),
    .Y(_1877_));
 sg13g2_nor3_1 _5636_ (.A(_1336_),
    .B(_1876_),
    .C(_1877_),
    .Y(_1878_));
 sg13g2_nor3_1 _5637_ (.A(net787),
    .B(net792),
    .C(_1044_),
    .Y(_1879_));
 sg13g2_nor3_1 _5638_ (.A(_1791_),
    .B(_1878_),
    .C(_1879_),
    .Y(_1880_));
 sg13g2_a21oi_1 _5639_ (.A1(net758),
    .A2(_1879_),
    .Y(_1881_),
    .B1(_0724_));
 sg13g2_o21ai_1 _5640_ (.B1(_1881_),
    .Y(_1882_),
    .A1(net787),
    .A2(_1052_));
 sg13g2_o21ai_1 _5641_ (.B1(_0842_),
    .Y(_1883_),
    .A1(_1880_),
    .A2(_1882_));
 sg13g2_nand2b_1 _5642_ (.Y(_1885_),
    .B(_1883_),
    .A_N(_1068_));
 sg13g2_nand3_1 _5643_ (.B(_0761_),
    .C(_0939_),
    .A(net695),
    .Y(_1886_));
 sg13g2_a22oi_1 _5644_ (.Y(_1887_),
    .B1(_1684_),
    .B2(_0912_),
    .A2(_1021_),
    .A1(net745));
 sg13g2_a221oi_1 _5645_ (.B2(_0729_),
    .C1(_0772_),
    .B1(_0894_),
    .A1(net698),
    .Y(_1888_),
    .A2(net729));
 sg13g2_nand2b_1 _5646_ (.Y(_1889_),
    .B(_1888_),
    .A_N(_1705_));
 sg13g2_o21ai_1 _5647_ (.B1(_1889_),
    .Y(_1890_),
    .A1(net692),
    .A2(_1887_));
 sg13g2_nand2b_1 _5648_ (.Y(_1891_),
    .B(_0756_),
    .A_N(_0730_));
 sg13g2_and2_1 _5649_ (.A(net695),
    .B(_1891_),
    .X(_1892_));
 sg13g2_inv_1 _5650_ (.Y(_1893_),
    .A(_1892_));
 sg13g2_nand2_1 _5651_ (.Y(_1894_),
    .A(_1849_),
    .B(_1860_));
 sg13g2_nor2_1 _5652_ (.A(net730),
    .B(_0991_),
    .Y(_1896_));
 sg13g2_a21oi_1 _5653_ (.A1(_0991_),
    .A2(_1894_),
    .Y(_1897_),
    .B1(_1896_));
 sg13g2_a221oi_1 _5654_ (.B2(_0848_),
    .C1(_1890_),
    .B1(_1897_),
    .A1(_0823_),
    .Y(_1898_),
    .A2(_1893_));
 sg13g2_o21ai_1 _5655_ (.B1(_1898_),
    .Y(_1899_),
    .A1(_0903_),
    .A2(_1743_));
 sg13g2_a21oi_1 _5656_ (.A1(_0937_),
    .A2(_1886_),
    .Y(_1900_),
    .B1(_1899_));
 sg13g2_nand2_1 _5657_ (.Y(_1901_),
    .A(net738),
    .B(net690));
 sg13g2_nand3_1 _5658_ (.B(_1201_),
    .C(_1901_),
    .A(_1022_),
    .Y(_1902_));
 sg13g2_nand2_1 _5659_ (.Y(_1903_),
    .A(net738),
    .B(_0953_));
 sg13g2_a21oi_1 _5660_ (.A1(net738),
    .A2(_0953_),
    .Y(_1904_),
    .B1(net751));
 sg13g2_nand3_1 _5661_ (.B(_0998_),
    .C(_1904_),
    .A(_0955_),
    .Y(_1905_));
 sg13g2_a21oi_1 _5662_ (.A1(net738),
    .A2(_0949_),
    .Y(_1907_),
    .B1(_0952_));
 sg13g2_nand3_1 _5663_ (.B(_0945_),
    .C(_1907_),
    .A(_0860_),
    .Y(_1908_));
 sg13g2_a21oi_1 _5664_ (.A1(_1259_),
    .A2(_0866_),
    .Y(_1909_),
    .B1(net673));
 sg13g2_nand2_1 _5665_ (.Y(_1910_),
    .A(net738),
    .B(_1016_));
 sg13g2_nand3_1 _5666_ (.B(_1728_),
    .C(_1910_),
    .A(_0820_),
    .Y(_1911_));
 sg13g2_o21ai_1 _5667_ (.B1(_0892_),
    .Y(_1912_),
    .A1(_1909_),
    .A2(_1911_));
 sg13g2_nand4_1 _5668_ (.B(_1905_),
    .C(_1908_),
    .A(_1902_),
    .Y(_1913_),
    .D(_1912_));
 sg13g2_o21ai_1 _5669_ (.B1(net672),
    .Y(_1914_),
    .A1(_0734_),
    .A2(_0832_));
 sg13g2_a221oi_1 _5670_ (.B2(_0884_),
    .C1(_0910_),
    .B1(net671),
    .A1(_1281_),
    .Y(_1915_),
    .A2(_0401_));
 sg13g2_a21oi_2 _5671_ (.B1(_0842_),
    .Y(_1916_),
    .A2(_1915_),
    .A1(_1914_));
 sg13g2_a21oi_1 _5672_ (.A1(_0964_),
    .A2(_1739_),
    .Y(_1918_),
    .B1(_0890_));
 sg13g2_nand2_1 _5673_ (.Y(_1919_),
    .A(_0968_),
    .B(_1918_));
 sg13g2_a22oi_1 _5674_ (.Y(_1920_),
    .B1(_0855_),
    .B2(net729),
    .A2(net757),
    .A1(_0125_));
 sg13g2_o21ai_1 _5675_ (.B1(_1919_),
    .Y(_1921_),
    .A1(_1719_),
    .A2(_1920_));
 sg13g2_nor4_1 _5676_ (.A(_0837_),
    .B(_1913_),
    .C(_1916_),
    .D(_1921_),
    .Y(_1922_));
 sg13g2_nand3_1 _5677_ (.B(_0745_),
    .C(net757),
    .A(_0715_),
    .Y(_1923_));
 sg13g2_nand3_1 _5678_ (.B(_1032_),
    .C(_1923_),
    .A(net688),
    .Y(_1924_));
 sg13g2_nand2_1 _5679_ (.Y(_1925_),
    .A(_0991_),
    .B(_1924_));
 sg13g2_nand2_1 _5680_ (.Y(_1926_),
    .A(_0826_),
    .B(_1004_));
 sg13g2_a21oi_1 _5681_ (.A1(_0783_),
    .A2(_0941_),
    .Y(_1927_),
    .B1(_1926_));
 sg13g2_a221oi_1 _5682_ (.B2(_1094_),
    .C1(_1927_),
    .B1(_1925_),
    .A1(_0909_),
    .Y(_1929_),
    .A2(_1850_));
 sg13g2_a22oi_1 _5683_ (.Y(_1930_),
    .B1(_0967_),
    .B2(_0999_),
    .A2(_0900_),
    .A1(_0897_));
 sg13g2_o21ai_1 _5684_ (.B1(_0974_),
    .Y(_1931_),
    .A1(_1187_),
    .A2(_1930_));
 sg13g2_nor2_1 _5685_ (.A(net693),
    .B(_1070_),
    .Y(_1932_));
 sg13g2_nor4_2 _5686_ (.A(_0235_),
    .B(net668),
    .C(_0941_),
    .Y(_1933_),
    .D(_1932_));
 sg13g2_nand2_1 _5687_ (.Y(_1934_),
    .A(_0831_),
    .B(_1933_));
 sg13g2_nand3_1 _5688_ (.B(_1204_),
    .C(net671),
    .A(net750),
    .Y(_1935_));
 sg13g2_o21ai_1 _5689_ (.B1(_1934_),
    .Y(_1936_),
    .A1(_0733_),
    .A2(_1935_));
 sg13g2_nand3_1 _5690_ (.B(_1003_),
    .C(_1011_),
    .A(_0800_),
    .Y(_1937_));
 sg13g2_and2_1 _5691_ (.A(_0867_),
    .B(_0988_),
    .X(_1938_));
 sg13g2_nand2_1 _5692_ (.Y(_1940_),
    .A(_1741_),
    .B(_1856_));
 sg13g2_a221oi_1 _5693_ (.B2(_1036_),
    .C1(_1937_),
    .B1(_1940_),
    .A1(_0992_),
    .Y(_1941_),
    .A2(_1938_));
 sg13g2_a22oi_1 _5694_ (.Y(_1942_),
    .B1(_1031_),
    .B2(_0953_),
    .A2(_1012_),
    .A1(net753));
 sg13g2_nand3b_1 _5695_ (.B(net762),
    .C(_0704_),
    .Y(_1943_),
    .A_N(net842));
 sg13g2_a21oi_1 _5696_ (.A1(_0705_),
    .A2(_1943_),
    .Y(_1944_),
    .B1(_1764_));
 sg13g2_or2_1 _5697_ (.X(_1945_),
    .B(_1944_),
    .A(_0785_));
 sg13g2_nor3_2 _5698_ (.A(net741),
    .B(_0756_),
    .C(_1038_),
    .Y(_1946_));
 sg13g2_a21oi_1 _5699_ (.A1(_1010_),
    .A2(_1945_),
    .Y(_1947_),
    .B1(_1946_));
 sg13g2_o21ai_1 _5700_ (.B1(_1737_),
    .Y(_1948_),
    .A1(_0738_),
    .A2(_0950_));
 sg13g2_a221oi_1 _5701_ (.B2(_0902_),
    .C1(_1948_),
    .B1(_1857_),
    .A1(_0932_),
    .Y(_1949_),
    .A2(_0965_));
 sg13g2_nand4_1 _5702_ (.B(_1942_),
    .C(_1947_),
    .A(_1941_),
    .Y(_1951_),
    .D(_1949_));
 sg13g2_o21ai_1 _5703_ (.B1(_0945_),
    .Y(_1952_),
    .A1(net746),
    .A2(_1005_));
 sg13g2_nand3_1 _5704_ (.B(_1711_),
    .C(_1952_),
    .A(_1007_),
    .Y(_1953_));
 sg13g2_nand2b_1 _5705_ (.Y(_1954_),
    .B(_1198_),
    .A_N(_1197_));
 sg13g2_nand2_1 _5706_ (.Y(_1955_),
    .A(net732),
    .B(net753));
 sg13g2_nand4_1 _5707_ (.B(net753),
    .C(net687),
    .A(net732),
    .Y(_1956_),
    .D(_0913_));
 sg13g2_a21o_1 _5708_ (.A2(_0953_),
    .A1(net733),
    .B1(_0996_),
    .X(_1957_));
 sg13g2_nand3_1 _5709_ (.B(_0892_),
    .C(_0985_),
    .A(net731),
    .Y(_1958_));
 sg13g2_nand2_1 _5710_ (.Y(_1959_),
    .A(_1957_),
    .B(_1958_));
 sg13g2_a221oi_1 _5711_ (.B2(_1677_),
    .C1(_1959_),
    .B1(_1020_),
    .A1(_0840_),
    .Y(_1960_),
    .A2(_0920_));
 sg13g2_nand4_1 _5712_ (.B(_1954_),
    .C(_1956_),
    .A(_1953_),
    .Y(_1962_),
    .D(_1960_));
 sg13g2_nor4_1 _5713_ (.A(_1931_),
    .B(_1936_),
    .C(_1951_),
    .D(_1962_),
    .Y(_1963_));
 sg13g2_nand4_1 _5714_ (.B(_1922_),
    .C(_1929_),
    .A(_1106_),
    .Y(_1964_),
    .D(_1963_));
 sg13g2_nand3b_1 _5715_ (.B(_1885_),
    .C(_1900_),
    .Y(_1965_),
    .A_N(_1964_));
 sg13g2_nand4_1 _5716_ (.B(net694),
    .C(_0832_),
    .A(_0231_),
    .Y(_1966_),
    .D(_0835_));
 sg13g2_or4_1 _5717_ (.A(_0703_),
    .B(_1839_),
    .C(_1866_),
    .D(_1965_),
    .X(_1967_));
 sg13g2_a221oi_1 _5718_ (.B2(_0614_),
    .C1(_1967_),
    .B1(net657),
    .A1(_0627_),
    .Y(_1968_),
    .A2(_1674_));
 sg13g2_nand3_1 _5719_ (.B(_1810_),
    .C(_1968_),
    .A(_1800_),
    .Y(_1969_));
 sg13g2_nand3_1 _5720_ (.B(_0396_),
    .C(_1797_),
    .A(_0335_),
    .Y(_1970_));
 sg13g2_a21oi_1 _5721_ (.A1(_1782_),
    .A2(_1970_),
    .Y(_1971_),
    .B1(_0285_));
 sg13g2_nor2_1 _5722_ (.A(_0308_),
    .B(_1971_),
    .Y(_1973_));
 sg13g2_nor2_1 _5723_ (.A(_0237_),
    .B(_1973_),
    .Y(_1974_));
 sg13g2_a221oi_1 _5724_ (.B2(_0230_),
    .C1(_1969_),
    .B1(_1974_),
    .A1(_1627_),
    .Y(_1975_),
    .A2(_1795_));
 sg13g2_nand3_1 _5725_ (.B(_1195_),
    .C(_1196_),
    .A(net737),
    .Y(_1976_));
 sg13g2_and3_1 _5726_ (.X(_1977_),
    .A(_1794_),
    .B(_1975_),
    .C(_1976_));
 sg13g2_a21oi_2 _5727_ (.B1(_1193_),
    .Y(uo_out[5]),
    .A2(_1977_),
    .A1(_1793_));
 sg13g2_nand2b_1 _5728_ (.Y(_1978_),
    .B(_2849_),
    .A_N(_1479_));
 sg13g2_a21oi_1 _5729_ (.A1(_1787_),
    .A2(_1978_),
    .Y(_1979_),
    .B1(_1336_));
 sg13g2_o21ai_1 _5730_ (.B1(_1303_),
    .Y(_1980_),
    .A1(_1791_),
    .A2(_1979_));
 sg13g2_o21ai_1 _5731_ (.B1(_1178_),
    .Y(_1981_),
    .A1(_1177_),
    .A2(_1185_));
 sg13g2_nor2_1 _5732_ (.A(net691),
    .B(_1657_),
    .Y(_1983_));
 sg13g2_a21o_1 _5733_ (.A2(_1983_),
    .A1(_1627_),
    .B1(_1206_),
    .X(_1984_));
 sg13g2_and2_2 _5734_ (.A(net754),
    .B(_0991_),
    .X(_1985_));
 sg13g2_inv_1 _5735_ (.Y(_1986_),
    .A(_1985_));
 sg13g2_nand2_1 _5736_ (.Y(_1987_),
    .A(_0366_),
    .B(_1985_));
 sg13g2_nand3_1 _5737_ (.B(_0396_),
    .C(_1987_),
    .A(_0309_),
    .Y(_1988_));
 sg13g2_nand3_1 _5738_ (.B(_0236_),
    .C(_1988_),
    .A(_0230_),
    .Y(_1989_));
 sg13g2_nand2b_1 _5739_ (.Y(_1990_),
    .B(_0405_),
    .A_N(_1809_));
 sg13g2_nor2_1 _5740_ (.A(_0307_),
    .B(_1162_),
    .Y(_1991_));
 sg13g2_o21ai_1 _5741_ (.B1(_1991_),
    .Y(_1992_),
    .A1(_1163_),
    .A2(_1986_));
 sg13g2_a22oi_1 _5742_ (.Y(_1994_),
    .B1(_1078_),
    .B2(_1081_),
    .A2(_0634_),
    .A1(_0513_));
 sg13g2_a21o_1 _5743_ (.A2(_1994_),
    .A1(net757),
    .B1(_1685_),
    .X(_1995_));
 sg13g2_nand2_1 _5744_ (.Y(_1996_),
    .A(_1085_),
    .B(_1098_));
 sg13g2_a21oi_1 _5745_ (.A1(_1684_),
    .A2(_1996_),
    .Y(_1997_),
    .B1(_0908_));
 sg13g2_and2_1 _5746_ (.A(_0934_),
    .B(_1036_),
    .X(_1998_));
 sg13g2_o21ai_1 _5747_ (.B1(_1998_),
    .Y(_1999_),
    .A1(_0805_),
    .A2(_0894_));
 sg13g2_nand2_1 _5748_ (.Y(_2000_),
    .A(_0934_),
    .B(_1188_));
 sg13g2_nand2_1 _5749_ (.Y(_2001_),
    .A(_0900_),
    .B(_2000_));
 sg13g2_nand2_1 _5750_ (.Y(_2002_),
    .A(_1999_),
    .B(_2001_));
 sg13g2_o21ai_1 _5751_ (.B1(_0839_),
    .Y(_2003_),
    .A1(_1075_),
    .A2(_1707_));
 sg13g2_nor3_1 _5752_ (.A(_1028_),
    .B(net663),
    .C(net746),
    .Y(_2005_));
 sg13g2_nor2_2 _5753_ (.A(_1013_),
    .B(_1100_),
    .Y(_2006_));
 sg13g2_nor2_2 _5754_ (.A(_1009_),
    .B(_1711_),
    .Y(_2007_));
 sg13g2_nor3_1 _5755_ (.A(_0918_),
    .B(_0940_),
    .C(net664),
    .Y(_2008_));
 sg13g2_o21ai_1 _5756_ (.B1(net657),
    .Y(_2009_),
    .A1(_1020_),
    .A2(_2008_));
 sg13g2_or4_1 _5757_ (.A(net698),
    .B(net729),
    .C(_0755_),
    .D(_0759_),
    .X(_2010_));
 sg13g2_nand3_1 _5758_ (.B(_0999_),
    .C(_1026_),
    .A(_0931_),
    .Y(_2011_));
 sg13g2_nor2b_1 _5759_ (.A(_1719_),
    .B_N(_1920_),
    .Y(_2012_));
 sg13g2_nand3_1 _5760_ (.B(_0783_),
    .C(_1004_),
    .A(net693),
    .Y(_2013_));
 sg13g2_a22oi_1 _5761_ (.Y(_2014_),
    .B1(_0987_),
    .B2(_0993_),
    .A2(_0848_),
    .A1(net739));
 sg13g2_nor3_1 _5762_ (.A(net663),
    .B(_0770_),
    .C(net756),
    .Y(_2016_));
 sg13g2_o21ai_1 _5763_ (.B1(_0939_),
    .Y(_2017_),
    .A1(_0937_),
    .A2(_0959_));
 sg13g2_a21oi_1 _5764_ (.A1(_1038_),
    .A2(_2017_),
    .Y(_2018_),
    .B1(_0782_));
 sg13g2_nand2_2 _5765_ (.Y(_2019_),
    .A(_0954_),
    .B(_1001_));
 sg13g2_o21ai_1 _5766_ (.B1(net764),
    .Y(_2020_),
    .A1(_0889_),
    .A2(_0935_));
 sg13g2_nand2_1 _5767_ (.Y(_2021_),
    .A(_0948_),
    .B(_1005_));
 sg13g2_nand2_1 _5768_ (.Y(_2022_),
    .A(_1007_),
    .B(_1945_));
 sg13g2_o21ai_1 _5769_ (.B1(_2022_),
    .Y(_2023_),
    .A1(net751),
    .A2(_1009_));
 sg13g2_a22oi_1 _5770_ (.Y(_2024_),
    .B1(_2021_),
    .B2(_2023_),
    .A2(_0971_),
    .A1(_0968_));
 sg13g2_nand3b_1 _5771_ (.B(_0968_),
    .C(_0932_),
    .Y(_2025_),
    .A_N(_1740_));
 sg13g2_nand2_2 _5772_ (.Y(_2027_),
    .A(_0868_),
    .B(_1201_));
 sg13g2_o21ai_1 _5773_ (.B1(_0867_),
    .Y(_2028_),
    .A1(net733),
    .A2(_1200_));
 sg13g2_nand2_1 _5774_ (.Y(_2029_),
    .A(_0816_),
    .B(_1718_));
 sg13g2_nand3_1 _5775_ (.B(_0901_),
    .C(_1188_),
    .A(net764),
    .Y(_2030_));
 sg13g2_a21o_2 _5776_ (.A2(_0840_),
    .A1(net735),
    .B1(_0772_),
    .X(_2031_));
 sg13g2_a21oi_1 _5777_ (.A1(net736),
    .A2(_0755_),
    .Y(_2032_),
    .B1(_0780_));
 sg13g2_nand2_1 _5778_ (.Y(_2033_),
    .A(net697),
    .B(_2032_));
 sg13g2_a21oi_2 _5779_ (.B1(_1727_),
    .Y(_2034_),
    .A2(_0844_),
    .A1(_0839_));
 sg13g2_a21oi_1 _5780_ (.A1(_1021_),
    .A2(_1985_),
    .Y(_2035_),
    .B1(_1997_));
 sg13g2_nand4_1 _5781_ (.B(_1703_),
    .C(_2024_),
    .A(_1702_),
    .Y(_2036_),
    .D(_2035_));
 sg13g2_nor4_1 _5782_ (.A(_1022_),
    .B(_1025_),
    .C(_1675_),
    .D(_1724_),
    .Y(_2038_));
 sg13g2_a22oi_1 _5783_ (.Y(_2039_),
    .B1(_2010_),
    .B2(_0979_),
    .A2(_1692_),
    .A1(_0930_));
 sg13g2_nand3_1 _5784_ (.B(_2011_),
    .C(_2029_),
    .A(_2003_),
    .Y(_2040_));
 sg13g2_nor3_1 _5785_ (.A(_2012_),
    .B(_2018_),
    .C(_2040_),
    .Y(_2041_));
 sg13g2_nand3_1 _5786_ (.B(_2039_),
    .C(_2041_),
    .A(_2030_),
    .Y(_2042_));
 sg13g2_nor4_2 _5787_ (.A(_1909_),
    .B(_2005_),
    .C(_2007_),
    .Y(_2043_),
    .D(_2016_));
 sg13g2_nor2_1 _5788_ (.A(_1678_),
    .B(_1735_),
    .Y(_2044_));
 sg13g2_nand4_1 _5789_ (.B(_2014_),
    .C(_2043_),
    .A(_2006_),
    .Y(_2045_),
    .D(_2044_));
 sg13g2_nand2_1 _5790_ (.Y(_2046_),
    .A(_0813_),
    .B(_1739_));
 sg13g2_nand3_1 _5791_ (.B(_1016_),
    .C(_2046_),
    .A(net667),
    .Y(_2047_));
 sg13g2_o21ai_1 _5792_ (.B1(net687),
    .Y(_2049_),
    .A1(_0909_),
    .A2(_0913_));
 sg13g2_nand2_1 _5793_ (.Y(_2050_),
    .A(_2020_),
    .B(_2049_));
 sg13g2_nand4_1 _5794_ (.B(_0887_),
    .C(_0890_),
    .A(_0875_),
    .Y(_2051_),
    .D(_0986_));
 sg13g2_nor4_1 _5795_ (.A(_0910_),
    .B(_1104_),
    .C(_2050_),
    .D(_2051_),
    .Y(_2052_));
 sg13g2_nand3_1 _5796_ (.B(_2047_),
    .C(_2052_),
    .A(_2025_),
    .Y(_2053_));
 sg13g2_nor3_1 _5797_ (.A(_2042_),
    .B(_2045_),
    .C(_2053_),
    .Y(_2054_));
 sg13g2_o21ai_1 _5798_ (.B1(_0991_),
    .Y(_2055_),
    .A1(_1094_),
    .A2(_0848_));
 sg13g2_o21ai_1 _5799_ (.B1(_1995_),
    .Y(_2056_),
    .A1(_1932_),
    .A2(_2033_));
 sg13g2_o21ai_1 _5800_ (.B1(_2031_),
    .Y(_2057_),
    .A1(_0828_),
    .A2(_0919_));
 sg13g2_nand3_1 _5801_ (.B(_2028_),
    .C(_2034_),
    .A(_2027_),
    .Y(_2058_));
 sg13g2_nor4_1 _5802_ (.A(_2002_),
    .B(_2056_),
    .C(_2057_),
    .D(_2058_),
    .Y(_2060_));
 sg13g2_nand4_1 _5803_ (.B(_2013_),
    .C(_2055_),
    .A(_2009_),
    .Y(_2061_),
    .D(_2060_));
 sg13g2_nor2_1 _5804_ (.A(_1839_),
    .B(_2061_),
    .Y(_2062_));
 sg13g2_nand4_1 _5805_ (.B(_2038_),
    .C(_2054_),
    .A(_2019_),
    .Y(_2063_),
    .D(_2062_));
 sg13g2_nor4_1 _5806_ (.A(_0628_),
    .B(_0703_),
    .C(_2036_),
    .D(_2063_),
    .Y(_2064_));
 sg13g2_a22oi_1 _5807_ (.Y(_2065_),
    .B1(_1992_),
    .B2(_1166_),
    .A2(_1673_),
    .A1(_0629_));
 sg13g2_and4_1 _5808_ (.A(_1989_),
    .B(_1990_),
    .C(_2064_),
    .D(_2065_),
    .X(_2066_));
 sg13g2_and4_1 _5809_ (.A(_1199_),
    .B(_1981_),
    .C(_1984_),
    .D(_2066_),
    .X(_2067_));
 sg13g2_a21oi_2 _5810_ (.B1(_1193_),
    .Y(uo_out[1]),
    .A2(_2067_),
    .A1(_1980_));
 sg13g2_nor2_1 _5811_ (.A(_1201_),
    .B(_1657_),
    .Y(_2068_));
 sg13g2_nor2_1 _5812_ (.A(_1206_),
    .B(_2068_),
    .Y(_2070_));
 sg13g2_o21ai_1 _5813_ (.B1(_1991_),
    .Y(_2071_),
    .A1(net754),
    .A2(_1163_));
 sg13g2_and2_1 _5814_ (.A(_1166_),
    .B(_2071_),
    .X(_2072_));
 sg13g2_a21oi_2 _5815_ (.B1(_1093_),
    .Y(_2073_),
    .A2(_0911_),
    .A1(net754));
 sg13g2_nand2_1 _5816_ (.Y(_2074_),
    .A(_1098_),
    .B(_2073_));
 sg13g2_a21oi_1 _5817_ (.A1(_1684_),
    .A2(_2074_),
    .Y(_2075_),
    .B1(_0908_));
 sg13g2_nand3_1 _5818_ (.B(_1005_),
    .C(_1007_),
    .A(_0948_),
    .Y(_2076_));
 sg13g2_nand2_1 _5819_ (.Y(_2077_),
    .A(_1713_),
    .B(_2076_));
 sg13g2_nor4_2 _5820_ (.A(_2007_),
    .B(_2072_),
    .C(_2075_),
    .Y(_2078_),
    .D(_2077_));
 sg13g2_nand2_1 _5821_ (.Y(_2079_),
    .A(_0496_),
    .B(_0500_));
 sg13g2_nor3_1 _5822_ (.A(_0503_),
    .B(_0506_),
    .C(_2079_),
    .Y(_2081_));
 sg13g2_a21o_1 _5823_ (.A2(_2079_),
    .A1(_0506_),
    .B1(_2081_),
    .X(_2082_));
 sg13g2_inv_1 _5824_ (.Y(_2083_),
    .A(_2082_));
 sg13g2_o21ai_1 _5825_ (.B1(_0405_),
    .Y(_2084_),
    .A1(_0494_),
    .A2(_2083_));
 sg13g2_nand3_1 _5826_ (.B(_0900_),
    .C(_0965_),
    .A(net667),
    .Y(_2085_));
 sg13g2_nand3_1 _5827_ (.B(_0913_),
    .C(_1955_),
    .A(net687),
    .Y(_2086_));
 sg13g2_nand2_1 _5828_ (.Y(_2087_),
    .A(_1012_),
    .B(_1200_));
 sg13g2_nand3_1 _5829_ (.B(_1034_),
    .C(_1903_),
    .A(_1031_),
    .Y(_2088_));
 sg13g2_a22oi_1 _5830_ (.Y(_2089_),
    .B1(_1202_),
    .B2(net690),
    .A2(_1016_),
    .A1(_0893_));
 sg13g2_nor3_1 _5831_ (.A(net738),
    .B(_0952_),
    .C(net657),
    .Y(_2090_));
 sg13g2_o21ai_1 _5832_ (.B1(_0844_),
    .Y(_2092_),
    .A1(net698),
    .A2(_0731_));
 sg13g2_nor3_1 _5833_ (.A(net661),
    .B(_0511_),
    .C(_0992_),
    .Y(_2093_));
 sg13g2_nand3_1 _5834_ (.B(_0631_),
    .C(_0909_),
    .A(net834),
    .Y(_2094_));
 sg13g2_o21ai_1 _5835_ (.B1(_2094_),
    .Y(_2095_),
    .A1(net728),
    .A2(_1728_));
 sg13g2_nor2_1 _5836_ (.A(_2093_),
    .B(_2095_),
    .Y(_2096_));
 sg13g2_nor3_1 _5837_ (.A(_0511_),
    .B(net669),
    .C(net687),
    .Y(_2097_));
 sg13g2_a21oi_1 _5838_ (.A1(net831),
    .A2(net737),
    .Y(_2098_),
    .B1(net755));
 sg13g2_nand2_1 _5839_ (.Y(_2099_),
    .A(net728),
    .B(_2098_));
 sg13g2_a22oi_1 _5840_ (.Y(_2100_),
    .B1(_0955_),
    .B2(_0859_),
    .A2(_0892_),
    .A1(_0889_));
 sg13g2_nor2_1 _5841_ (.A(net726),
    .B(_0904_),
    .Y(_2101_));
 sg13g2_nor2_1 _5842_ (.A(net758),
    .B(net726),
    .Y(_2103_));
 sg13g2_o21ai_1 _5843_ (.B1(_0935_),
    .Y(_2104_),
    .A1(_0816_),
    .A2(_2103_));
 sg13g2_nand2_1 _5844_ (.Y(_2105_),
    .A(_0633_),
    .B(_0804_));
 sg13g2_a221oi_1 _5845_ (.B2(net657),
    .C1(_1102_),
    .B1(_1103_),
    .A1(net755),
    .Y(_2106_),
    .A2(_1021_));
 sg13g2_o21ai_1 _5846_ (.B1(_2106_),
    .Y(_2107_),
    .A1(_0826_),
    .A2(_1038_));
 sg13g2_o21ai_1 _5847_ (.B1(_0823_),
    .Y(_2108_),
    .A1(net698),
    .A2(_0760_));
 sg13g2_nor3_1 _5848_ (.A(net662),
    .B(_0866_),
    .C(_2000_),
    .Y(_2109_));
 sg13g2_o21ai_1 _5849_ (.B1(_0979_),
    .Y(_2110_),
    .A1(_0836_),
    .A2(_1844_));
 sg13g2_a21oi_1 _5850_ (.A1(_1084_),
    .A2(_2073_),
    .Y(_2111_),
    .B1(net692));
 sg13g2_nor2_1 _5851_ (.A(_1685_),
    .B(_2111_),
    .Y(_2112_));
 sg13g2_nand2_1 _5852_ (.Y(_2114_),
    .A(_0939_),
    .B(_1892_));
 sg13g2_nand3_1 _5853_ (.B(_1004_),
    .C(_2114_),
    .A(_0783_),
    .Y(_2115_));
 sg13g2_nor2_1 _5854_ (.A(_1070_),
    .B(_1891_),
    .Y(_2116_));
 sg13g2_nor3_1 _5855_ (.A(net740),
    .B(_0829_),
    .C(_2116_),
    .Y(_2117_));
 sg13g2_nor3_2 _5856_ (.A(_0780_),
    .B(_0941_),
    .C(_2117_),
    .Y(_2118_));
 sg13g2_o21ai_1 _5857_ (.B1(net695),
    .Y(_2119_),
    .A1(_0760_),
    .A2(_1073_));
 sg13g2_nand3_1 _5858_ (.B(_0959_),
    .C(_2119_),
    .A(_0824_),
    .Y(_2120_));
 sg13g2_nand2_1 _5859_ (.Y(_2121_),
    .A(_0969_),
    .B(_1018_));
 sg13g2_a22oi_1 _5860_ (.Y(_2122_),
    .B1(_1707_),
    .B2(net658),
    .A2(_1075_),
    .A1(net697));
 sg13g2_a21oi_1 _5861_ (.A1(net736),
    .A2(_0840_),
    .Y(_2123_),
    .B1(_2122_));
 sg13g2_nand2_1 _5862_ (.Y(_2125_),
    .A(_0977_),
    .B(_1100_));
 sg13g2_nand3_1 _5863_ (.B(_0991_),
    .C(_1032_),
    .A(_0848_),
    .Y(_2126_));
 sg13g2_nand2_2 _5864_ (.Y(_2127_),
    .A(_0917_),
    .B(_0937_));
 sg13g2_o21ai_1 _5865_ (.B1(_0987_),
    .Y(_2128_),
    .A1(net690),
    .A2(_0860_));
 sg13g2_nor2_1 _5866_ (.A(_1896_),
    .B(_2128_),
    .Y(_2129_));
 sg13g2_nor2_1 _5867_ (.A(_0932_),
    .B(_0999_),
    .Y(_2130_));
 sg13g2_a21oi_1 _5868_ (.A1(net731),
    .A2(_0812_),
    .Y(_2131_),
    .B1(_2130_));
 sg13g2_o21ai_1 _5869_ (.B1(net728),
    .Y(_2132_),
    .A1(_0902_),
    .A2(_2131_));
 sg13g2_a22oi_1 _5870_ (.Y(_2133_),
    .B1(_2099_),
    .B2(_0873_),
    .A2(_0983_),
    .A1(_0893_));
 sg13g2_a21oi_1 _5871_ (.A1(_1998_),
    .A2(_2105_),
    .Y(_2134_),
    .B1(_2123_));
 sg13g2_o21ai_1 _5872_ (.B1(_2092_),
    .Y(_2136_),
    .A1(_0919_),
    .A2(_1892_));
 sg13g2_nor3_1 _5873_ (.A(_2107_),
    .B(_2109_),
    .C(_2136_),
    .Y(_2137_));
 sg13g2_nand4_1 _5874_ (.B(_2108_),
    .C(_2134_),
    .A(_2104_),
    .Y(_2138_),
    .D(_2137_));
 sg13g2_o21ai_1 _5875_ (.B1(_2110_),
    .Y(_2139_),
    .A1(_0936_),
    .A2(_2127_));
 sg13g2_a22oi_1 _5876_ (.Y(_2140_),
    .B1(_1985_),
    .B2(_1094_),
    .A2(_0930_),
    .A1(_0927_));
 sg13g2_nand4_1 _5877_ (.B(_2121_),
    .C(_2132_),
    .A(_0846_),
    .Y(_2141_),
    .D(_2140_));
 sg13g2_nor3_1 _5878_ (.A(_2112_),
    .B(_2118_),
    .C(_2141_),
    .Y(_2142_));
 sg13g2_a221oi_1 _5879_ (.B2(_1024_),
    .C1(_2097_),
    .B1(_2101_),
    .A1(_0954_),
    .Y(_2143_),
    .A2(_1736_));
 sg13g2_a221oi_1 _5880_ (.B2(_0965_),
    .C1(_0997_),
    .B1(_0891_),
    .A1(_1072_),
    .Y(_2144_),
    .A2(_0767_));
 sg13g2_and4_1 _5881_ (.A(_1003_),
    .B(_1966_),
    .C(_2096_),
    .D(_2144_),
    .X(_2145_));
 sg13g2_and4_1 _5882_ (.A(_2100_),
    .B(_2133_),
    .C(_2143_),
    .D(_2145_),
    .X(_2147_));
 sg13g2_and4_1 _5883_ (.A(_2027_),
    .B(_2028_),
    .C(_2087_),
    .D(_2089_),
    .X(_2148_));
 sg13g2_nand4_1 _5884_ (.B(_2125_),
    .C(_2147_),
    .A(_0972_),
    .Y(_2149_),
    .D(_2148_));
 sg13g2_nor4_1 _5885_ (.A(net742),
    .B(net661),
    .C(_0886_),
    .D(net751),
    .Y(_2150_));
 sg13g2_nand2_1 _5886_ (.Y(_2151_),
    .A(_2031_),
    .B(_2085_));
 sg13g2_nor3_2 _5887_ (.A(_2090_),
    .B(_2150_),
    .C(_2151_),
    .Y(_2152_));
 sg13g2_nand4_1 _5888_ (.B(_2088_),
    .C(_2126_),
    .A(_2086_),
    .Y(_2153_),
    .D(_2152_));
 sg13g2_nor4_2 _5889_ (.A(_0821_),
    .B(_1933_),
    .C(_2149_),
    .Y(_2154_),
    .D(_2153_));
 sg13g2_o21ai_1 _5890_ (.B1(_0986_),
    .Y(_2155_),
    .A1(_0893_),
    .A2(_1011_));
 sg13g2_o21ai_1 _5891_ (.B1(net729),
    .Y(_2156_),
    .A1(_1998_),
    .A2(_2155_));
 sg13g2_nand3_1 _5892_ (.B(_2120_),
    .C(_2156_),
    .A(_2115_),
    .Y(_2158_));
 sg13g2_nor4_1 _5893_ (.A(_2129_),
    .B(_2138_),
    .C(_2139_),
    .D(_2158_),
    .Y(_2159_));
 sg13g2_nand3_1 _5894_ (.B(_2154_),
    .C(_2159_),
    .A(_2142_),
    .Y(_2160_));
 sg13g2_a22oi_1 _5895_ (.Y(_2161_),
    .B1(_1041_),
    .B2(_0551_),
    .A2(_0926_),
    .A1(_0424_));
 sg13g2_nor3_1 _5896_ (.A(net783),
    .B(_0125_),
    .C(_2161_),
    .Y(_2162_));
 sg13g2_a21oi_1 _5897_ (.A1(net736),
    .A2(_2161_),
    .Y(_2163_),
    .B1(_2162_));
 sg13g2_o21ai_1 _5898_ (.B1(_0479_),
    .Y(_2164_),
    .A1(_0745_),
    .A2(_1689_));
 sg13g2_a221oi_1 _5899_ (.B2(_0219_),
    .C1(_2164_),
    .B1(_1045_),
    .A1(net833),
    .Y(_2165_),
    .A2(_0723_));
 sg13g2_o21ai_1 _5900_ (.B1(_2165_),
    .Y(_2166_),
    .A1(_1690_),
    .A2(_2163_));
 sg13g2_a21oi_1 _5901_ (.A1(_0842_),
    .A2(_2166_),
    .Y(_2167_),
    .B1(_1068_));
 sg13g2_nor4_2 _5902_ (.A(_0614_),
    .B(_0744_),
    .C(_2160_),
    .Y(_2169_),
    .D(_2167_));
 sg13g2_nand3_1 _5903_ (.B(_2084_),
    .C(_2169_),
    .A(_2078_),
    .Y(_2170_));
 sg13g2_a21o_1 _5904_ (.A2(_2070_),
    .A1(_1627_),
    .B1(_2170_),
    .X(_2171_));
 sg13g2_a21oi_1 _5905_ (.A1(_0479_),
    .A2(_1788_),
    .Y(_2172_),
    .B1(_1723_));
 sg13g2_nor2b_1 _5906_ (.A(_1195_),
    .B_N(_1196_),
    .Y(_2173_));
 sg13g2_nand2_1 _5907_ (.Y(_2174_),
    .A(_0366_),
    .B(net757));
 sg13g2_a21o_1 _5908_ (.A2(_2174_),
    .A1(_1164_),
    .B1(_0225_),
    .X(_2175_));
 sg13g2_a21oi_2 _5909_ (.B1(_0237_),
    .Y(_2176_),
    .A2(_2175_),
    .A1(_0230_));
 sg13g2_nor3_1 _5910_ (.A(_0978_),
    .B(_2173_),
    .C(_2176_),
    .Y(_2177_));
 sg13g2_or3_1 _5911_ (.A(_0805_),
    .B(_1177_),
    .C(_1185_),
    .X(_2178_));
 sg13g2_nor4_1 _5912_ (.A(_0978_),
    .B(_2171_),
    .C(_2173_),
    .D(_2176_),
    .Y(_2180_));
 sg13g2_a22oi_1 _5913_ (.Y(_2181_),
    .B1(_2178_),
    .B2(_1178_),
    .A2(_2172_),
    .A1(_1790_));
 sg13g2_a21oi_2 _5914_ (.B1(_1193_),
    .Y(uo_out[6]),
    .A2(_2181_),
    .A1(_2180_));
 sg13g2_or2_1 _5915_ (.X(_2182_),
    .B(_1479_),
    .A(_1336_));
 sg13g2_o21ai_1 _5916_ (.B1(_1303_),
    .Y(_2183_),
    .A1(_2849_),
    .A2(_2182_));
 sg13g2_nand3_1 _5917_ (.B(_0495_),
    .C(_2082_),
    .A(_0405_),
    .Y(_2184_));
 sg13g2_nand2b_1 _5918_ (.Y(_2185_),
    .B(_2073_),
    .A_N(_1994_));
 sg13g2_a21oi_1 _5919_ (.A1(net688),
    .A2(_2185_),
    .Y(_2186_),
    .B1(_1685_));
 sg13g2_a22oi_1 _5920_ (.Y(_2187_),
    .B1(_1718_),
    .B2(_0977_),
    .A2(_1018_),
    .A1(_0968_));
 sg13g2_a22oi_1 _5921_ (.Y(_2188_),
    .B1(_1735_),
    .B2(_1856_),
    .A2(_0976_),
    .A1(_0901_));
 sg13g2_a21oi_1 _5922_ (.A1(net758),
    .A2(_1740_),
    .Y(_2190_),
    .B1(_1733_));
 sg13g2_a21oi_1 _5923_ (.A1(_0934_),
    .A2(_0999_),
    .Y(_2191_),
    .B1(_2190_));
 sg13g2_nor2_2 _5924_ (.A(_0952_),
    .B(_1904_),
    .Y(_2192_));
 sg13g2_nor2_1 _5925_ (.A(_0834_),
    .B(_0843_),
    .Y(_2193_));
 sg13g2_nor2_1 _5926_ (.A(_2192_),
    .B(_2193_),
    .Y(_2194_));
 sg13g2_nand4_1 _5927_ (.B(_2188_),
    .C(_2191_),
    .A(_2187_),
    .Y(_2195_),
    .D(_2194_));
 sg13g2_and2_1 _5928_ (.A(_2027_),
    .B(_2127_),
    .X(_2196_));
 sg13g2_nand2_1 _5929_ (.Y(_2197_),
    .A(_1745_),
    .B(_1957_));
 sg13g2_nor3_1 _5930_ (.A(_1732_),
    .B(_1918_),
    .C(_2197_),
    .Y(_2198_));
 sg13g2_nand4_1 _5931_ (.B(_2089_),
    .C(_2196_),
    .A(_2087_),
    .Y(_2199_),
    .D(_2198_));
 sg13g2_o21ai_1 _5932_ (.B1(_1707_),
    .Y(_2201_),
    .A1(net697),
    .A2(net736));
 sg13g2_o21ai_1 _5933_ (.B1(_1031_),
    .Y(_2202_),
    .A1(net738),
    .A2(_0954_));
 sg13g2_nor2_1 _5934_ (.A(_1201_),
    .B(_1719_),
    .Y(_2203_));
 sg13g2_a21oi_1 _5935_ (.A1(_0888_),
    .A2(net657),
    .Y(_2204_),
    .B1(_2203_));
 sg13g2_nand2_1 _5936_ (.Y(_2205_),
    .A(_0724_),
    .B(_0795_));
 sg13g2_and2_1 _5937_ (.A(_0939_),
    .B(_1004_),
    .X(_2206_));
 sg13g2_o21ai_1 _5938_ (.B1(net672),
    .Y(_2207_),
    .A1(_0734_),
    .A2(_0817_));
 sg13g2_nand2b_1 _5939_ (.Y(_2208_),
    .B(_0839_),
    .A_N(_2207_));
 sg13g2_o21ai_1 _5940_ (.B1(_2208_),
    .Y(_2209_),
    .A1(_0724_),
    .A2(_0960_));
 sg13g2_a221oi_1 _5941_ (.B2(_0839_),
    .C1(_2209_),
    .B1(_2206_),
    .A1(_0799_),
    .Y(_2210_),
    .A2(_2205_));
 sg13g2_nand4_1 _5942_ (.B(_2202_),
    .C(_2204_),
    .A(_2201_),
    .Y(_2212_),
    .D(_2210_));
 sg13g2_nor2_1 _5943_ (.A(_0815_),
    .B(_1011_),
    .Y(_2213_));
 sg13g2_a21oi_1 _5944_ (.A1(_0970_),
    .A2(_0971_),
    .Y(_2214_),
    .B1(_2213_));
 sg13g2_nand3_1 _5945_ (.B(_2034_),
    .C(_2214_),
    .A(_2025_),
    .Y(_2215_));
 sg13g2_nor3_1 _5946_ (.A(_0235_),
    .B(net660),
    .C(_0857_),
    .Y(_2216_));
 sg13g2_o21ai_1 _5947_ (.B1(_2006_),
    .Y(_2217_),
    .A1(net727),
    .A2(_1728_));
 sg13g2_nor4_1 _5948_ (.A(_0771_),
    .B(_0979_),
    .C(_1020_),
    .D(_1030_),
    .Y(_2218_));
 sg13g2_nand4_1 _5949_ (.B(_0875_),
    .C(_1721_),
    .A(_1105_),
    .Y(_2219_),
    .D(_2218_));
 sg13g2_nor3_1 _5950_ (.A(_2216_),
    .B(_2217_),
    .C(_2219_),
    .Y(_2220_));
 sg13g2_a22oi_1 _5951_ (.Y(_2221_),
    .B1(_1198_),
    .B2(net690),
    .A2(_1033_),
    .A1(_0955_));
 sg13g2_a22oi_1 _5952_ (.Y(_2223_),
    .B1(_1036_),
    .B2(_0893_),
    .A2(_1024_),
    .A1(_0895_));
 sg13g2_o21ai_1 _5953_ (.B1(_1075_),
    .Y(_2224_),
    .A1(net736),
    .A2(net659));
 sg13g2_nand2_1 _5954_ (.Y(_2225_),
    .A(_1002_),
    .B(_2224_));
 sg13g2_a221oi_1 _5955_ (.B2(_0900_),
    .C1(_2225_),
    .B1(_1856_),
    .A1(_0889_),
    .Y(_2226_),
    .A2(_0976_));
 sg13g2_nand4_1 _5956_ (.B(_2221_),
    .C(_2223_),
    .A(_2220_),
    .Y(_2227_),
    .D(_2226_));
 sg13g2_nor4_1 _5957_ (.A(_2199_),
    .B(_2212_),
    .C(_2215_),
    .D(_2227_),
    .Y(_2228_));
 sg13g2_nand3_1 _5958_ (.B(net671),
    .C(_1743_),
    .A(_1248_),
    .Y(_2229_));
 sg13g2_a22oi_1 _5959_ (.Y(_2230_),
    .B1(_2032_),
    .B2(net659),
    .A2(_0910_),
    .A1(net693));
 sg13g2_nor2b_1 _5960_ (.A(_2230_),
    .B_N(_0835_),
    .Y(_2231_));
 sg13g2_a21oi_1 _5961_ (.A1(_0909_),
    .A2(_1201_),
    .Y(_2232_),
    .B1(_0913_));
 sg13g2_nor2_1 _5962_ (.A(_1850_),
    .B(_2232_),
    .Y(_2234_));
 sg13g2_nor4_1 _5963_ (.A(_1696_),
    .B(_2107_),
    .C(_2231_),
    .D(_2234_),
    .Y(_2235_));
 sg13g2_nand3_1 _5964_ (.B(_2229_),
    .C(_2235_),
    .A(_2228_),
    .Y(_2236_));
 sg13g2_nand2_1 _5965_ (.Y(_2237_),
    .A(_1681_),
    .B(_2184_));
 sg13g2_nor4_1 _5966_ (.A(_2186_),
    .B(_2195_),
    .C(_2236_),
    .D(_2237_),
    .Y(_2238_));
 sg13g2_nand3_1 _5967_ (.B(_2183_),
    .C(_2238_),
    .A(_2078_),
    .Y(_2239_));
 sg13g2_a21oi_1 _5968_ (.A1(_1849_),
    .A2(_1983_),
    .Y(_2240_),
    .B1(_1206_));
 sg13g2_a221oi_1 _5969_ (.B2(_1627_),
    .C1(_2239_),
    .B1(_2240_),
    .A1(_1178_),
    .Y(_2241_),
    .A2(_1667_));
 sg13g2_a21oi_2 _5970_ (.B1(_1193_),
    .Y(uo_out[2]),
    .A2(_2241_),
    .A1(_2177_));
 sg13g2_or2_1 _5971_ (.X(_2242_),
    .B(\counter[0] ),
    .A(\counter[1] ));
 sg13g2_nand2b_2 _5972_ (.Y(_2244_),
    .B(_0074_),
    .A_N(_2242_));
 sg13g2_o21ai_1 _5973_ (.B1(\counter[4] ),
    .Y(_2245_),
    .A1(\counter[3] ),
    .A2(_2244_));
 sg13g2_o21ai_1 _5974_ (.B1(_0006_),
    .Y(_2246_),
    .A1(\counter[5] ),
    .A2(_2245_));
 sg13g2_nor2b_2 _5975_ (.A(_0005_),
    .B_N(_2246_),
    .Y(_2247_));
 sg13g2_o21ai_1 _5976_ (.B1(net5),
    .Y(_2248_),
    .A1(\counter[0] ),
    .A2(_2247_));
 sg13g2_a22oi_1 _5977_ (.Y(_2249_),
    .B1(_0283_),
    .B2(_0360_),
    .A2(net4),
    .A1(\counter[0] ));
 sg13g2_nor2_1 _5978_ (.A(\counter[0] ),
    .B(net770),
    .Y(_2250_));
 sg13g2_a21oi_1 _5979_ (.A1(_2248_),
    .A2(_2249_),
    .Y(_2251_),
    .B1(_0371_));
 sg13g2_nor3_1 _5980_ (.A(net6),
    .B(_2250_),
    .C(_2251_),
    .Y(_0026_));
 sg13g2_nand2_2 _5981_ (.Y(_2252_),
    .A(\counter[1] ),
    .B(\counter[0] ));
 sg13g2_nand2_1 _5982_ (.Y(_2254_),
    .A(_2242_),
    .B(_2252_));
 sg13g2_or3_1 _5983_ (.A(\counter[4] ),
    .B(\counter[3] ),
    .C(_2244_),
    .X(_2255_));
 sg13g2_or2_1 _5984_ (.X(_2256_),
    .B(_2255_),
    .A(\counter[5] ));
 sg13g2_o21ai_1 _5985_ (.B1(net4),
    .Y(_2257_),
    .A1(\counter[6] ),
    .A2(_2256_));
 sg13g2_nor2_2 _5986_ (.A(net5),
    .B(_2257_),
    .Y(_2258_));
 sg13g2_inv_1 _5987_ (.Y(_2259_),
    .A(_2258_));
 sg13g2_nor2b_2 _5988_ (.A(_2247_),
    .B_N(net5),
    .Y(_2260_));
 sg13g2_nand2b_1 _5989_ (.Y(_2261_),
    .B(net5),
    .A_N(_2247_));
 sg13g2_nand2b_1 _5990_ (.Y(_2262_),
    .B(_2260_),
    .A_N(_2254_));
 sg13g2_a221oi_1 _5991_ (.B2(_2258_),
    .C1(_0371_),
    .B1(_2254_),
    .A1(net8),
    .Y(_2263_),
    .A2(_0360_));
 sg13g2_a221oi_1 _5992_ (.B2(_2263_),
    .C1(net6),
    .B1(_2262_),
    .A1(_0085_),
    .Y(_0027_),
    .A2(_0371_));
 sg13g2_o21ai_1 _5993_ (.B1(_2260_),
    .Y(_2265_),
    .A1(_0008_),
    .A2(_2252_));
 sg13g2_a21o_1 _5994_ (.A2(_2252_),
    .A1(_0008_),
    .B1(_2265_),
    .X(_2266_));
 sg13g2_xor2_1 _5995_ (.B(_2242_),
    .A(_0008_),
    .X(_2267_));
 sg13g2_a221oi_1 _5996_ (.B2(_2267_),
    .C1(_0371_),
    .B1(_2258_),
    .A1(net9),
    .Y(_2268_),
    .A2(_0360_));
 sg13g2_a221oi_1 _5997_ (.B2(_2268_),
    .C1(net6),
    .B1(_2266_),
    .A1(_0074_),
    .Y(_0028_),
    .A2(_0371_));
 sg13g2_nand2_1 _5998_ (.Y(_2269_),
    .A(_2244_),
    .B(_2258_));
 sg13g2_nor2_1 _5999_ (.A(_2244_),
    .B(_2259_),
    .Y(_2270_));
 sg13g2_nor3_1 _6000_ (.A(_0008_),
    .B(_2252_),
    .C(_2261_),
    .Y(_2271_));
 sg13g2_o21ai_1 _6001_ (.B1(_0009_),
    .Y(_2272_),
    .A1(_2270_),
    .A2(_2271_));
 sg13g2_a21oi_1 _6002_ (.A1(_2265_),
    .A2(_2269_),
    .Y(_2274_),
    .B1(_0009_));
 sg13g2_a21oi_1 _6003_ (.A1(net10),
    .A2(_0360_),
    .Y(_2275_),
    .B1(_2274_));
 sg13g2_nand3_1 _6004_ (.B(_2272_),
    .C(_2275_),
    .A(net770),
    .Y(_2276_));
 sg13g2_o21ai_1 _6005_ (.B1(_2276_),
    .Y(_2277_),
    .A1(\counter[3] ),
    .A2(net770));
 sg13g2_nor2_1 _6006_ (.A(net6),
    .B(_2277_),
    .Y(_0029_));
 sg13g2_nand4_1 _6007_ (.B(\counter[2] ),
    .C(\counter[1] ),
    .A(\counter[3] ),
    .Y(_2278_),
    .D(\counter[0] ));
 sg13g2_inv_1 _6008_ (.Y(_2279_),
    .A(_2278_));
 sg13g2_o21ai_1 _6009_ (.B1(_2260_),
    .Y(_2280_),
    .A1(_0010_),
    .A2(_2278_));
 sg13g2_a21oi_1 _6010_ (.A1(_0010_),
    .A2(_2278_),
    .Y(_2281_),
    .B1(_2280_));
 sg13g2_nand3_1 _6011_ (.B(_2245_),
    .C(_2255_),
    .A(net4),
    .Y(_2282_));
 sg13g2_o21ai_1 _6012_ (.B1(_2282_),
    .Y(_2284_),
    .A1(net4),
    .A2(net11));
 sg13g2_o21ai_1 _6013_ (.B1(_0382_),
    .Y(_2285_),
    .A1(net5),
    .A2(_2284_));
 sg13g2_nor2_1 _6014_ (.A(_2281_),
    .B(_2285_),
    .Y(_2286_));
 sg13g2_nor2_1 _6015_ (.A(\counter[4] ),
    .B(net770),
    .Y(_2287_));
 sg13g2_nor3_1 _6016_ (.A(net6),
    .B(_2286_),
    .C(_2287_),
    .Y(_0030_));
 sg13g2_nand2_1 _6017_ (.Y(_2288_),
    .A(_2255_),
    .B(_2258_));
 sg13g2_nor2_1 _6018_ (.A(_2255_),
    .B(_2259_),
    .Y(_2289_));
 sg13g2_nor3_1 _6019_ (.A(_0010_),
    .B(_2261_),
    .C(_2278_),
    .Y(_2290_));
 sg13g2_o21ai_1 _6020_ (.B1(_0006_),
    .Y(_2291_),
    .A1(_2289_),
    .A2(_2290_));
 sg13g2_a21oi_1 _6021_ (.A1(_2280_),
    .A2(_2288_),
    .Y(_2292_),
    .B1(_0006_));
 sg13g2_a21oi_1 _6022_ (.A1(net12),
    .A2(_0360_),
    .Y(_2294_),
    .B1(_2292_));
 sg13g2_nand3_1 _6023_ (.B(_2291_),
    .C(_2294_),
    .A(net770),
    .Y(_2295_));
 sg13g2_o21ai_1 _6024_ (.B1(_2295_),
    .Y(_2296_),
    .A1(\counter[5] ),
    .A2(net770));
 sg13g2_nor2_1 _6025_ (.A(net6),
    .B(_2296_),
    .Y(_0031_));
 sg13g2_nand3_1 _6026_ (.B(\counter[4] ),
    .C(_2279_),
    .A(\counter[5] ),
    .Y(_2297_));
 sg13g2_xor2_1 _6027_ (.B(_2297_),
    .A(_0005_),
    .X(_2298_));
 sg13g2_a21o_1 _6028_ (.A2(_2256_),
    .A1(\counter[6] ),
    .B1(_2257_),
    .X(_2299_));
 sg13g2_o21ai_1 _6029_ (.B1(_2299_),
    .Y(_2300_),
    .A1(net4),
    .A2(net13));
 sg13g2_o21ai_1 _6030_ (.B1(net770),
    .Y(_2301_),
    .A1(net5),
    .A2(_2300_));
 sg13g2_a21oi_1 _6031_ (.A1(_2260_),
    .A2(_2298_),
    .Y(_2302_),
    .B1(_2301_));
 sg13g2_nor2_1 _6032_ (.A(\counter[6] ),
    .B(net770),
    .Y(_2304_));
 sg13g2_nor3_1 _6033_ (.A(net6),
    .B(_2302_),
    .C(_2304_),
    .Y(_0032_));
 sg13g2_nand3_1 _6034_ (.B(net782),
    .C(_2855_),
    .A(net789),
    .Y(_2305_));
 sg13g2_nor4_2 _6035_ (.A(net804),
    .B(_1446_),
    .C(_0411_),
    .Y(_2306_),
    .D(_2305_));
 sg13g2_nor2b_1 _6036_ (.A(_2306_),
    .B_N(net1),
    .Y(_2307_));
 sg13g2_nand2b_2 _6037_ (.Y(_2308_),
    .B(net1),
    .A_N(_2306_));
 sg13g2_nand2_1 _6038_ (.Y(_2309_),
    .A(net864),
    .B(net682));
 sg13g2_nand4_1 _6039_ (.B(\hvsync_gen.vpos[9] ),
    .C(net769),
    .A(net778),
    .Y(_2310_),
    .D(net762));
 sg13g2_o21ai_1 _6040_ (.B1(net1),
    .Y(_2311_),
    .A1(_1662_),
    .A2(_2310_));
 sg13g2_inv_1 _6041_ (.Y(_2312_),
    .A(_2311_));
 sg13g2_nand2_2 _6042_ (.Y(_2314_),
    .A(_2306_),
    .B(_2312_));
 sg13g2_o21ai_1 _6043_ (.B1(_2309_),
    .Y(_0033_),
    .A1(_0063_),
    .A2(_2314_));
 sg13g2_nand2_1 _6044_ (.Y(_2315_),
    .A(net859),
    .B(net682));
 sg13g2_o21ai_1 _6045_ (.B1(_2315_),
    .Y(_0034_),
    .A1(_2069_),
    .A2(_2314_));
 sg13g2_nand3_1 _6046_ (.B(_0414_),
    .C(_2308_),
    .A(net856),
    .Y(_2316_));
 sg13g2_nor2_2 _6047_ (.A(net682),
    .B(_2312_),
    .Y(_2317_));
 sg13g2_a21oi_1 _6048_ (.A1(_0414_),
    .A2(_2308_),
    .Y(_2318_),
    .B1(net856));
 sg13g2_nor2_1 _6049_ (.A(_2317_),
    .B(_2318_),
    .Y(_2319_));
 sg13g2_and2_1 _6050_ (.A(_2316_),
    .B(_2319_),
    .X(_0035_));
 sg13g2_nand2_1 _6051_ (.Y(_2320_),
    .A(net852),
    .B(net682));
 sg13g2_nor2_1 _6052_ (.A(net65),
    .B(_0425_),
    .Y(_2322_));
 sg13g2_xnor2_1 _6053_ (.Y(_2323_),
    .A(net852),
    .B(_2322_));
 sg13g2_o21ai_1 _6054_ (.B1(_2320_),
    .Y(_0036_),
    .A1(_2314_),
    .A2(_2323_));
 sg13g2_nor2_1 _6055_ (.A(_0376_),
    .B(_2316_),
    .Y(_2324_));
 sg13g2_a21oi_1 _6056_ (.A1(_0414_),
    .A2(_2308_),
    .Y(_2325_),
    .B1(net850));
 sg13g2_nor4_1 _6057_ (.A(_0535_),
    .B(_2317_),
    .C(_2324_),
    .D(_2325_),
    .Y(_0037_));
 sg13g2_nand2_1 _6058_ (.Y(_2326_),
    .A(net847),
    .B(net681));
 sg13g2_nand3b_1 _6059_ (.B(_0414_),
    .C(net769),
    .Y(_2327_),
    .A_N(_0016_));
 sg13g2_xnor2_1 _6060_ (.Y(_2328_),
    .A(_0140_),
    .B(_2327_));
 sg13g2_o21ai_1 _6061_ (.B1(_2326_),
    .Y(_0038_),
    .A1(_2314_),
    .A2(_2328_));
 sg13g2_nor2_1 _6062_ (.A(net841),
    .B(_2324_),
    .Y(_2330_));
 sg13g2_nor3_1 _6063_ (.A(_0590_),
    .B(_0376_),
    .C(_2316_),
    .Y(_2331_));
 sg13g2_nor4_1 _6064_ (.A(_0153_),
    .B(_2317_),
    .C(_2330_),
    .D(_2331_),
    .Y(_0039_));
 sg13g2_nand2_1 _6065_ (.Y(_2332_),
    .A(net837),
    .B(net681));
 sg13g2_nor2_1 _6066_ (.A(_0012_),
    .B(_1835_),
    .Y(_2333_));
 sg13g2_xnor2_1 _6067_ (.Y(_2334_),
    .A(net837),
    .B(_2333_));
 sg13g2_o21ai_1 _6068_ (.B1(_2332_),
    .Y(_0040_),
    .A1(_2314_),
    .A2(_2334_));
 sg13g2_or3_1 _6069_ (.A(net768),
    .B(_1835_),
    .C(net681),
    .X(_2335_));
 sg13g2_a221oi_1 _6070_ (.B2(net778),
    .C1(_2317_),
    .B1(_2335_),
    .A1(net760),
    .Y(_0041_),
    .A2(_2331_));
 sg13g2_nor3_1 _6071_ (.A(net830),
    .B(_0568_),
    .C(_1835_),
    .Y(_2336_));
 sg13g2_nor2_1 _6072_ (.A(net61),
    .B(_2336_),
    .Y(_2338_));
 sg13g2_a21oi_1 _6073_ (.A1(\hvsync_gen.vpos[9] ),
    .A2(_2336_),
    .Y(_2339_),
    .B1(_2314_));
 sg13g2_a21oi_1 _6074_ (.A1(net61),
    .A2(net681),
    .Y(_2340_),
    .B1(_2339_));
 sg13g2_nor2_1 _6075_ (.A(_2338_),
    .B(_2340_),
    .Y(_0042_));
 sg13g2_nor2_1 _6076_ (.A(_0349_),
    .B(_2308_),
    .Y(_0043_));
 sg13g2_nor2_1 _6077_ (.A(_1950_),
    .B(_2308_),
    .Y(_0044_));
 sg13g2_nor2_1 _6078_ (.A(_2925_),
    .B(_2308_),
    .Y(_0045_));
 sg13g2_nor2_1 _6079_ (.A(_2877_),
    .B(_2308_),
    .Y(_0046_));
 sg13g2_and2_1 _6080_ (.A(net1),
    .B(_1238_),
    .X(_0047_));
 sg13g2_o21ai_1 _6081_ (.B1(net681),
    .Y(_2341_),
    .A1(net761),
    .A2(_1591_));
 sg13g2_a21oi_1 _6082_ (.A1(net776),
    .A2(net761),
    .Y(_0048_),
    .B1(_2341_));
 sg13g2_nand2_2 _6083_ (.Y(_2343_),
    .A(net803),
    .B(_1236_));
 sg13g2_a21o_1 _6084_ (.A2(_1236_),
    .A1(_0418_),
    .B1(_2308_),
    .X(_2344_));
 sg13g2_a21oi_1 _6085_ (.A1(_0228_),
    .A2(_2343_),
    .Y(_0049_),
    .B1(_2344_));
 sg13g2_nor2_1 _6086_ (.A(net796),
    .B(_2343_),
    .Y(_2345_));
 sg13g2_o21ai_1 _6087_ (.B1(net681),
    .Y(_2346_),
    .A1(net794),
    .A2(_2345_));
 sg13g2_a21oi_1 _6088_ (.A1(net794),
    .A2(_2345_),
    .Y(_0050_),
    .B1(_2346_));
 sg13g2_nor2_1 _6089_ (.A(_0677_),
    .B(_2343_),
    .Y(_2347_));
 sg13g2_o21ai_1 _6090_ (.B1(net681),
    .Y(_2348_),
    .A1(net786),
    .A2(_2347_));
 sg13g2_a21oi_1 _6091_ (.A1(net786),
    .A2(_2347_),
    .Y(_0051_),
    .B1(_2348_));
 sg13g2_nor3_1 _6092_ (.A(net59),
    .B(_0677_),
    .C(_2343_),
    .Y(_2350_));
 sg13g2_o21ai_1 _6093_ (.B1(net681),
    .Y(_2351_),
    .A1(net782),
    .A2(_2350_));
 sg13g2_a21oi_1 _6094_ (.A1(net782),
    .A2(_2350_),
    .Y(_0052_),
    .B1(_2351_));
 sg13g2_dfrbp_1 _6095_ (.CLK(counter_clk),
    .RESET_B(net37),
    .D(_0026_),
    .Q_N(_3042_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _6096_ (.CLK(counter_clk),
    .RESET_B(net30),
    .D(_0027_),
    .Q_N(_3041_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _6097_ (.CLK(counter_clk),
    .RESET_B(net57),
    .D(_0028_),
    .Q_N(_0008_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _6098_ (.CLK(counter_clk),
    .RESET_B(net55),
    .D(_0029_),
    .Q_N(_0009_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _6099_ (.CLK(counter_clk),
    .RESET_B(net53),
    .D(_0030_),
    .Q_N(_0010_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _6100_ (.CLK(counter_clk),
    .RESET_B(net51),
    .D(_0031_),
    .Q_N(_0006_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _6101_ (.CLK(counter_clk),
    .RESET_B(net48),
    .D(_0032_),
    .Q_N(_0005_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _6102_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net49),
    .D(_0000_),
    .Q_N(_3040_),
    .Q(hsync));
 sg13g2_dfrbp_1 _6103_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net46),
    .D(_0033_),
    .Q_N(_0025_),
    .Q(\flag.flag_abrosexual_inst.pix_y[0] ));
 sg13g2_dfrbp_1 _6104_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net44),
    .D(_0034_),
    .Q_N(_0022_),
    .Q(\flag.flag_abrosexual_inst.pix_y[1] ));
 sg13g2_dfrbp_1 _6105_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net42),
    .D(_0035_),
    .Q_N(_0019_),
    .Q(\flag.flag_abrosexual_inst.pix_y[2] ));
 sg13g2_dfrbp_1 _6106_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net40),
    .D(_0036_),
    .Q_N(_0002_),
    .Q(\flag.flag_abrosexual_inst.pix_y[3] ));
 sg13g2_dfrbp_1 _6107_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net38),
    .D(_0037_),
    .Q_N(_0016_),
    .Q(\flag.flag_abrosexual_inst.pix_y[4] ));
 sg13g2_dfrbp_1 _6108_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net35),
    .D(_0038_),
    .Q_N(_0003_),
    .Q(\flag.flag_abrosexual_inst.pix_y[5] ));
 sg13g2_dfrbp_1 _6109_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net33),
    .D(_0039_),
    .Q_N(_0012_),
    .Q(\flag.flag_abrosexual_inst.pix_y[6] ));
 sg13g2_dfrbp_1 _6110_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net31),
    .D(_0040_),
    .Q_N(_0013_),
    .Q(\flag.flag_abrosexual_inst.pix_y[7] ));
 sg13g2_dfrbp_1 _6111_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net56),
    .D(_0041_),
    .Q_N(_0011_),
    .Q(\flag.flag_abrosexual_inst.pix_y[8] ));
 sg13g2_dfrbp_1 _6112_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net50),
    .D(net62),
    .Q_N(_3043_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _6113_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net52),
    .D(_0001_),
    .Q_N(_3039_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 _6114_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net47),
    .D(_0043_),
    .Q_N(_0024_),
    .Q(\flag.flag_abrosexual_inst.pix_x[0] ));
 sg13g2_dfrbp_1 _6115_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net45),
    .D(_0044_),
    .Q_N(_0023_),
    .Q(\flag.flag_abrosexual_inst.pix_x[1] ));
 sg13g2_dfrbp_1 _6116_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net43),
    .D(_0045_),
    .Q_N(_0021_),
    .Q(\flag.flag_abrosexual_inst.pix_x[2] ));
 sg13g2_dfrbp_1 _6117_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net41),
    .D(_0046_),
    .Q_N(_0020_),
    .Q(\flag.flag_abrosexual_inst.pix_x[3] ));
 sg13g2_dfrbp_1 _6118_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net39),
    .D(_0047_),
    .Q_N(_0018_),
    .Q(\flag.flag_abrosexual_inst.pix_x[4] ));
 sg13g2_dfrbp_1 _6119_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net36),
    .D(_0048_),
    .Q_N(_0017_),
    .Q(\flag.flag_abrosexual_inst.pix_x[5] ));
 sg13g2_dfrbp_1 _6120_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net34),
    .D(_0049_),
    .Q_N(_0015_),
    .Q(\flag.flag_abrosexual_inst.pix_x[6] ));
 sg13g2_dfrbp_1 _6121_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net32),
    .D(_0050_),
    .Q_N(_0014_),
    .Q(\flag.flag_abrosexual_inst.pix_x[7] ));
 sg13g2_dfrbp_1 _6122_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net58),
    .D(_0051_),
    .Q_N(_0007_),
    .Q(\flag.flag_abrosexual_inst.pix_x[8] ));
 sg13g2_dfrbp_1 _6123_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net54),
    .D(_0052_),
    .Q_N(_0004_),
    .Q(\flag.flag_abrosexual_inst.pix_x[9] ));
 sg13g2_tiehi _6110__31 (.L_HI(net31));
 sg13g2_tiehi _6121__32 (.L_HI(net32));
 sg13g2_tiehi _6109__33 (.L_HI(net33));
 sg13g2_tiehi _6120__34 (.L_HI(net34));
 sg13g2_tiehi _6108__35 (.L_HI(net35));
 sg13g2_tiehi _6119__36 (.L_HI(net36));
 sg13g2_tiehi _6095__37 (.L_HI(net37));
 sg13g2_tiehi _6107__38 (.L_HI(net38));
 sg13g2_tiehi _6118__39 (.L_HI(net39));
 sg13g2_tiehi _6106__40 (.L_HI(net40));
 sg13g2_tiehi _6117__41 (.L_HI(net41));
 sg13g2_tiehi _6105__42 (.L_HI(net42));
 sg13g2_tiehi _6116__43 (.L_HI(net43));
 sg13g2_tiehi _6104__44 (.L_HI(net44));
 sg13g2_tiehi _6115__45 (.L_HI(net45));
 sg13g2_tiehi _6103__46 (.L_HI(net46));
 sg13g2_tiehi _6114__47 (.L_HI(net47));
 sg13g2_tiehi _6101__48 (.L_HI(net48));
 sg13g2_tiehi _6102__49 (.L_HI(net49));
 sg13g2_tiehi _6112__50 (.L_HI(net50));
 sg13g2_tiehi _6100__51 (.L_HI(net51));
 sg13g2_tiehi _6113__52 (.L_HI(net52));
 sg13g2_tiehi _6099__53 (.L_HI(net53));
 sg13g2_tiehi _6123__54 (.L_HI(net54));
 sg13g2_tiehi _6098__55 (.L_HI(net55));
 sg13g2_tiehi _6111__56 (.L_HI(net56));
 sg13g2_tiehi _6097__57 (.L_HI(net57));
 sg13g2_tiehi _6122__58 (.L_HI(net58));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_15 (.L_LO(net15));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_16 (.L_LO(net16));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_17 (.L_LO(net17));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_18 (.L_LO(net18));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_19 (.L_LO(net19));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_20 (.L_LO(net20));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_21 (.L_LO(net21));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_22 (.L_LO(net22));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_23 (.L_LO(net23));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_24 (.L_LO(net24));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_25 (.L_LO(net25));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_26 (.L_LO(net26));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_27 (.L_LO(net27));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_28 (.L_LO(net28));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_29 (.L_LO(net29));
 sg13g2_tiehi _6096__30 (.L_HI(net30));
 sg13g2_buf_1 _6169_ (.A(\hvsync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _6170_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout657 (.X(net657),
    .A(_1677_));
 sg13g2_buf_4 fanout658 (.X(net658),
    .A(_0776_));
 sg13g2_buf_2 fanout659 (.A(_0776_),
    .X(net659));
 sg13g2_buf_4 fanout660 (.X(net660),
    .A(_0404_));
 sg13g2_buf_2 fanout661 (.A(_0404_),
    .X(net661));
 sg13g2_buf_4 fanout662 (.X(net662),
    .A(net663));
 sg13g2_buf_2 fanout663 (.A(net665),
    .X(net663));
 sg13g2_buf_4 fanout664 (.X(net664),
    .A(net665));
 sg13g2_buf_2 fanout665 (.A(_1292_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(net667),
    .X(net666));
 sg13g2_buf_4 fanout667 (.X(net667),
    .A(_0806_));
 sg13g2_buf_4 fanout668 (.X(net668),
    .A(_0768_));
 sg13g2_buf_2 fanout669 (.A(_0768_),
    .X(net669));
 sg13g2_buf_4 fanout670 (.X(net670),
    .A(_0641_));
 sg13g2_buf_4 fanout671 (.X(net671),
    .A(_0640_));
 sg13g2_buf_2 fanout672 (.A(_0640_),
    .X(net672));
 sg13g2_buf_4 fanout673 (.X(net673),
    .A(_0232_));
 sg13g2_buf_4 fanout674 (.X(net674),
    .A(_0232_));
 sg13g2_buf_4 fanout675 (.X(net675),
    .A(_0176_));
 sg13g2_buf_4 fanout676 (.X(net676),
    .A(_2879_));
 sg13g2_buf_4 fanout677 (.X(net677),
    .A(_2542_));
 sg13g2_buf_4 fanout678 (.X(net678),
    .A(_2371_));
 sg13g2_buf_2 fanout679 (.A(net680),
    .X(net679));
 sg13g2_buf_4 fanout680 (.X(net680),
    .A(_2355_));
 sg13g2_buf_4 fanout681 (.X(net681),
    .A(_2307_));
 sg13g2_buf_1 fanout682 (.A(_2307_),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(_1274_),
    .X(net683));
 sg13g2_buf_1 fanout684 (.A(_1274_),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(_1245_),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(_1240_),
    .X(net686));
 sg13g2_buf_4 fanout687 (.X(net687),
    .A(net688));
 sg13g2_buf_4 fanout688 (.X(net688),
    .A(_0856_));
 sg13g2_buf_4 fanout689 (.X(net689),
    .A(_0855_));
 sg13g2_buf_4 fanout690 (.X(net690),
    .A(net691));
 sg13g2_buf_4 fanout691 (.X(net691),
    .A(net692));
 sg13g2_buf_2 fanout692 (.A(_0855_),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(net694),
    .X(net693));
 sg13g2_buf_4 fanout694 (.X(net694),
    .A(_0725_));
 sg13g2_buf_2 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_1 fanout696 (.A(net697),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(_0713_),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(net699),
    .X(net698));
 sg13g2_buf_4 fanout699 (.X(net699),
    .A(_0712_));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(_0160_));
 sg13g2_buf_4 fanout701 (.X(net701),
    .A(net703));
 sg13g2_buf_1 fanout702 (.A(net703),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(_0155_),
    .X(net703));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(_2415_));
 sg13g2_buf_1 fanout705 (.A(_2415_),
    .X(net705));
 sg13g2_buf_4 fanout706 (.X(net706),
    .A(_2405_));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(_2405_));
 sg13g2_buf_4 fanout708 (.X(net708),
    .A(_2396_));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(_2392_));
 sg13g2_buf_2 fanout710 (.A(_2392_),
    .X(net710));
 sg13g2_buf_4 fanout711 (.X(net711),
    .A(_2329_));
 sg13g2_buf_2 fanout712 (.A(_2329_),
    .X(net712));
 sg13g2_buf_4 fanout713 (.X(net713),
    .A(_2283_));
 sg13g2_buf_2 fanout714 (.A(net715),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(net716),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(_2243_),
    .X(net716));
 sg13g2_buf_4 fanout717 (.X(net717),
    .A(net718));
 sg13g2_buf_4 fanout718 (.X(net718),
    .A(_2211_));
 sg13g2_buf_4 fanout719 (.X(net719),
    .A(_2102_));
 sg13g2_buf_4 fanout720 (.X(net720),
    .A(_2091_));
 sg13g2_buf_2 fanout721 (.A(net723),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(net723),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_1884_),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(net725),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(_1665_),
    .X(net725));
 sg13g2_buf_4 fanout726 (.X(net726),
    .A(net727));
 sg13g2_buf_2 fanout727 (.A(_0810_),
    .X(net727));
 sg13g2_buf_4 fanout728 (.X(net728),
    .A(_0809_));
 sg13g2_buf_2 fanout729 (.A(_0748_),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(_0748_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(net734),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(net734),
    .X(net732));
 sg13g2_buf_4 fanout733 (.X(net733),
    .A(net734));
 sg13g2_buf_4 fanout734 (.X(net734),
    .A(_0748_));
 sg13g2_buf_4 fanout735 (.X(net735),
    .A(net736));
 sg13g2_buf_4 fanout736 (.X(net736),
    .A(_0747_));
 sg13g2_buf_4 fanout737 (.X(net737),
    .A(net739));
 sg13g2_buf_2 fanout738 (.A(net739),
    .X(net738));
 sg13g2_buf_4 fanout739 (.X(net739),
    .A(_0747_));
 sg13g2_buf_4 fanout740 (.X(net740),
    .A(net741));
 sg13g2_buf_2 fanout741 (.A(_0720_),
    .X(net741));
 sg13g2_buf_4 fanout742 (.X(net742),
    .A(net743));
 sg13g2_buf_4 fanout743 (.X(net743),
    .A(_1818_));
 sg13g2_buf_4 fanout744 (.X(net744),
    .A(net745));
 sg13g2_buf_4 fanout745 (.X(net745),
    .A(net746));
 sg13g2_buf_4 fanout746 (.X(net746),
    .A(net747));
 sg13g2_buf_4 fanout747 (.X(net747),
    .A(_1807_));
 sg13g2_buf_4 fanout748 (.X(net748),
    .A(net749));
 sg13g2_buf_2 fanout749 (.A(_1611_),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(_0896_),
    .X(net750));
 sg13g2_buf_4 fanout751 (.X(net751),
    .A(_0944_));
 sg13g2_buf_2 fanout752 (.A(_0944_),
    .X(net752));
 sg13g2_buf_4 fanout753 (.X(net753),
    .A(net754));
 sg13g2_buf_4 fanout754 (.X(net754),
    .A(_0793_));
 sg13g2_buf_4 fanout755 (.X(net755),
    .A(net757));
 sg13g2_buf_1 fanout756 (.A(net757),
    .X(net756));
 sg13g2_buf_4 fanout757 (.X(net757),
    .A(_0792_));
 sg13g2_buf_4 fanout758 (.X(net758),
    .A(_0746_));
 sg13g2_buf_2 fanout759 (.A(_1325_),
    .X(net759));
 sg13g2_buf_4 fanout760 (.X(net760),
    .A(_1149_));
 sg13g2_buf_4 fanout761 (.X(net761),
    .A(_1928_));
 sg13g2_buf_2 fanout762 (.A(_1687_),
    .X(net762));
 sg13g2_buf_4 fanout763 (.X(net763),
    .A(_1314_));
 sg13g2_buf_2 fanout764 (.A(net766),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(net766),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(_1160_),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(_0721_),
    .X(net767));
 sg13g2_buf_4 fanout768 (.X(net768),
    .A(_0568_));
 sg13g2_buf_4 fanout769 (.X(net769),
    .A(_0524_));
 sg13g2_buf_2 fanout770 (.A(_0382_),
    .X(net770));
 sg13g2_buf_4 fanout771 (.X(net771),
    .A(_0349_));
 sg13g2_buf_4 fanout772 (.X(net772),
    .A(_0294_));
 sg13g2_buf_4 fanout773 (.X(net773),
    .A(_0261_));
 sg13g2_buf_4 fanout774 (.X(net774),
    .A(net775));
 sg13g2_buf_4 fanout775 (.X(net775),
    .A(_0250_));
 sg13g2_buf_4 fanout776 (.X(net776),
    .A(net777));
 sg13g2_buf_4 fanout777 (.X(net777),
    .A(_0239_));
 sg13g2_buf_4 fanout778 (.X(net778),
    .A(net779));
 sg13g2_buf_4 fanout779 (.X(net779),
    .A(_0162_));
 sg13g2_buf_4 fanout780 (.X(net780),
    .A(net781));
 sg13g2_buf_2 fanout781 (.A(_0004_),
    .X(net781));
 sg13g2_buf_4 fanout782 (.X(net782),
    .A(net784));
 sg13g2_buf_4 fanout783 (.X(net783),
    .A(net784));
 sg13g2_buf_2 fanout784 (.A(\flag.flag_abrosexual_inst.pix_x[9] ),
    .X(net784));
 sg13g2_buf_4 fanout785 (.X(net785),
    .A(_0007_));
 sg13g2_buf_4 fanout786 (.X(net786),
    .A(net789));
 sg13g2_buf_4 fanout787 (.X(net787),
    .A(net789));
 sg13g2_buf_2 fanout788 (.A(net789),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(\flag.flag_abrosexual_inst.pix_x[8] ),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(net795),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(net795),
    .X(net791));
 sg13g2_buf_4 fanout792 (.X(net792),
    .A(net795));
 sg13g2_buf_2 fanout793 (.A(net795),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(net795),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(\flag.flag_abrosexual_inst.pix_x[7] ),
    .X(net795));
 sg13g2_buf_4 fanout796 (.X(net796),
    .A(net64));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(net799));
 sg13g2_buf_2 fanout798 (.A(net799),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(net800),
    .X(net799));
 sg13g2_buf_4 fanout800 (.X(net800),
    .A(\flag.flag_abrosexual_inst.pix_x[6] ));
 sg13g2_buf_4 fanout801 (.X(net801),
    .A(net802));
 sg13g2_buf_4 fanout802 (.X(net802),
    .A(_0017_));
 sg13g2_buf_4 fanout803 (.X(net803),
    .A(net804));
 sg13g2_buf_4 fanout804 (.X(net804),
    .A(\flag.flag_abrosexual_inst.pix_x[5] ));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(_0018_));
 sg13g2_buf_4 fanout806 (.X(net806),
    .A(_0018_));
 sg13g2_buf_4 fanout807 (.X(net807),
    .A(\flag.flag_abrosexual_inst.pix_x[4] ));
 sg13g2_buf_2 fanout808 (.A(\flag.flag_abrosexual_inst.pix_x[4] ),
    .X(net808));
 sg13g2_buf_4 fanout809 (.X(net809),
    .A(_0020_));
 sg13g2_buf_2 fanout810 (.A(net811),
    .X(net810));
 sg13g2_buf_4 fanout811 (.X(net811),
    .A(net812));
 sg13g2_buf_4 fanout812 (.X(net812),
    .A(\flag.flag_abrosexual_inst.pix_x[3] ));
 sg13g2_buf_4 fanout813 (.X(net813),
    .A(_0021_));
 sg13g2_buf_2 fanout814 (.A(net815),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(net816),
    .X(net815));
 sg13g2_buf_4 fanout816 (.X(net816),
    .A(\flag.flag_abrosexual_inst.pix_x[2] ));
 sg13g2_buf_2 fanout817 (.A(net819),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(net819),
    .X(net818));
 sg13g2_buf_4 fanout819 (.X(net819),
    .A(\flag.flag_abrosexual_inst.pix_x[1] ));
 sg13g2_buf_4 fanout820 (.X(net820),
    .A(net821));
 sg13g2_buf_4 fanout821 (.X(net821),
    .A(net60));
 sg13g2_buf_2 fanout822 (.A(net825),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(net825),
    .X(net823));
 sg13g2_buf_4 fanout824 (.X(net824),
    .A(net825));
 sg13g2_buf_2 fanout825 (.A(\flag.flag_abrosexual_inst.pix_x[0] ),
    .X(net825));
 sg13g2_buf_4 fanout826 (.X(net826),
    .A(net827));
 sg13g2_buf_2 fanout827 (.A(\flag.flag_abrosexual_inst.pix_x[0] ),
    .X(net827));
 sg13g2_buf_4 fanout828 (.X(net828),
    .A(net829));
 sg13g2_buf_2 fanout829 (.A(net832),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(net832),
    .X(net830));
 sg13g2_buf_1 fanout831 (.A(net832),
    .X(net831));
 sg13g2_buf_4 fanout832 (.X(net832),
    .A(_0011_));
 sg13g2_buf_4 fanout833 (.X(net833),
    .A(net836));
 sg13g2_buf_4 fanout834 (.X(net834),
    .A(net836));
 sg13g2_buf_2 fanout835 (.A(net836),
    .X(net835));
 sg13g2_buf_4 fanout836 (.X(net836),
    .A(\flag.flag_abrosexual_inst.pix_y[8] ));
 sg13g2_buf_2 fanout837 (.A(net838),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(net839),
    .X(net838));
 sg13g2_buf_4 fanout839 (.X(net839),
    .A(\flag.flag_abrosexual_inst.pix_y[7] ));
 sg13g2_buf_2 fanout840 (.A(net843),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(net843),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(net843),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(\flag.flag_abrosexual_inst.pix_y[6] ),
    .X(net843));
 sg13g2_buf_8 fanout844 (.A(_0003_),
    .X(net844));
 sg13g2_buf_4 fanout845 (.X(net845),
    .A(_0003_));
 sg13g2_buf_2 fanout846 (.A(net848),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(net848),
    .X(net847));
 sg13g2_buf_4 fanout848 (.X(net848),
    .A(net849));
 sg13g2_buf_8 fanout849 (.A(\flag.flag_abrosexual_inst.pix_y[5] ),
    .X(net849));
 sg13g2_buf_4 fanout850 (.X(net850),
    .A(net851));
 sg13g2_buf_4 fanout851 (.X(net851),
    .A(\flag.flag_abrosexual_inst.pix_y[4] ));
 sg13g2_buf_2 fanout852 (.A(net853),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(net854),
    .X(net853));
 sg13g2_buf_4 fanout854 (.X(net854),
    .A(net855));
 sg13g2_buf_4 fanout855 (.X(net855),
    .A(\flag.flag_abrosexual_inst.pix_y[3] ));
 sg13g2_buf_2 fanout856 (.A(net857),
    .X(net856));
 sg13g2_buf_4 fanout857 (.X(net857),
    .A(net858));
 sg13g2_buf_4 fanout858 (.X(net858),
    .A(\flag.flag_abrosexual_inst.pix_y[2] ));
 sg13g2_buf_2 fanout859 (.A(net860),
    .X(net859));
 sg13g2_buf_4 fanout860 (.X(net860),
    .A(\flag.flag_abrosexual_inst.pix_y[1] ));
 sg13g2_buf_2 fanout861 (.A(net866),
    .X(net861));
 sg13g2_buf_4 fanout862 (.X(net862),
    .A(net866));
 sg13g2_buf_4 fanout863 (.X(net863),
    .A(net865));
 sg13g2_buf_2 fanout864 (.A(net865),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(net866),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(\flag.flag_abrosexual_inst.pix_y[0] ),
    .X(net866));
 sg13g2_buf_4 fanout867 (.X(net867),
    .A(net2));
 sg13g2_buf_4 input1 (.X(net1),
    .A(rst_n));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[5]));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[6]));
 sg13g2_buf_2 input6 (.A(ui_in[7]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[0]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[1]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[4]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[5]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[6]),
    .X(net13));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_14 (.L_LO(net14));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0007_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0024_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold3 (.A(\hvsync_gen.vpos[9] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0042_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold5 (.A(\flag.flag_abrosexual_inst.pix_y[4] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0015_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0019_),
    .X(net65));
 sg13g2_antennanp ANTENNA_1 (.A(_0000_));
 sg13g2_antennanp ANTENNA_2 (.A(_0000_));
 sg13g2_antennanp ANTENNA_3 (.A(_0000_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_4 FILLER_0_214 ();
 sg13g2_fill_1 FILLER_0_228 ();
 sg13g2_decap_8 FILLER_0_233 ();
 sg13g2_decap_8 FILLER_0_240 ();
 sg13g2_decap_8 FILLER_0_247 ();
 sg13g2_decap_8 FILLER_0_254 ();
 sg13g2_decap_8 FILLER_0_261 ();
 sg13g2_decap_8 FILLER_0_268 ();
 sg13g2_decap_8 FILLER_0_275 ();
 sg13g2_decap_8 FILLER_0_282 ();
 sg13g2_decap_8 FILLER_0_289 ();
 sg13g2_decap_8 FILLER_0_296 ();
 sg13g2_fill_2 FILLER_0_303 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_fill_2 FILLER_0_329 ();
 sg13g2_decap_4 FILLER_0_346 ();
 sg13g2_fill_1 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_356 ();
 sg13g2_decap_8 FILLER_0_368 ();
 sg13g2_decap_8 FILLER_0_375 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_389 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_4 FILLER_0_403 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_fill_2 FILLER_1_196 ();
 sg13g2_fill_2 FILLER_1_222 ();
 sg13g2_fill_1 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_249 ();
 sg13g2_decap_8 FILLER_1_256 ();
 sg13g2_decap_8 FILLER_1_263 ();
 sg13g2_decap_8 FILLER_1_270 ();
 sg13g2_decap_8 FILLER_1_277 ();
 sg13g2_decap_8 FILLER_1_284 ();
 sg13g2_decap_8 FILLER_1_291 ();
 sg13g2_fill_1 FILLER_1_298 ();
 sg13g2_decap_8 FILLER_1_375 ();
 sg13g2_decap_8 FILLER_1_382 ();
 sg13g2_decap_8 FILLER_1_389 ();
 sg13g2_decap_8 FILLER_1_396 ();
 sg13g2_decap_4 FILLER_1_403 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_fill_2 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_fill_1 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_195 ();
 sg13g2_fill_2 FILLER_2_202 ();
 sg13g2_fill_1 FILLER_2_204 ();
 sg13g2_decap_4 FILLER_2_214 ();
 sg13g2_fill_1 FILLER_2_218 ();
 sg13g2_fill_1 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_234 ();
 sg13g2_fill_2 FILLER_2_241 ();
 sg13g2_fill_1 FILLER_2_254 ();
 sg13g2_decap_8 FILLER_2_258 ();
 sg13g2_decap_8 FILLER_2_265 ();
 sg13g2_decap_8 FILLER_2_272 ();
 sg13g2_decap_8 FILLER_2_279 ();
 sg13g2_decap_8 FILLER_2_286 ();
 sg13g2_decap_8 FILLER_2_293 ();
 sg13g2_decap_4 FILLER_2_300 ();
 sg13g2_fill_2 FILLER_2_308 ();
 sg13g2_fill_1 FILLER_2_310 ();
 sg13g2_decap_8 FILLER_2_316 ();
 sg13g2_decap_8 FILLER_2_323 ();
 sg13g2_fill_1 FILLER_2_330 ();
 sg13g2_fill_2 FILLER_2_334 ();
 sg13g2_fill_2 FILLER_2_349 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_4 FILLER_3_168 ();
 sg13g2_fill_1 FILLER_3_172 ();
 sg13g2_fill_1 FILLER_3_204 ();
 sg13g2_decap_8 FILLER_3_265 ();
 sg13g2_decap_8 FILLER_3_272 ();
 sg13g2_decap_8 FILLER_3_279 ();
 sg13g2_fill_2 FILLER_3_286 ();
 sg13g2_fill_1 FILLER_3_288 ();
 sg13g2_decap_4 FILLER_3_295 ();
 sg13g2_fill_2 FILLER_3_338 ();
 sg13g2_fill_1 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_346 ();
 sg13g2_decap_4 FILLER_3_353 ();
 sg13g2_fill_2 FILLER_3_357 ();
 sg13g2_decap_4 FILLER_3_368 ();
 sg13g2_fill_1 FILLER_3_372 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_fill_2 FILLER_4_175 ();
 sg13g2_fill_1 FILLER_4_177 ();
 sg13g2_decap_8 FILLER_4_187 ();
 sg13g2_decap_4 FILLER_4_194 ();
 sg13g2_decap_8 FILLER_4_211 ();
 sg13g2_fill_2 FILLER_4_218 ();
 sg13g2_fill_1 FILLER_4_220 ();
 sg13g2_decap_8 FILLER_4_225 ();
 sg13g2_fill_1 FILLER_4_232 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_4 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_258 ();
 sg13g2_decap_8 FILLER_4_265 ();
 sg13g2_decap_8 FILLER_4_272 ();
 sg13g2_decap_8 FILLER_4_279 ();
 sg13g2_fill_2 FILLER_4_286 ();
 sg13g2_fill_1 FILLER_4_288 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_fill_1 FILLER_4_301 ();
 sg13g2_fill_2 FILLER_4_369 ();
 sg13g2_fill_1 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_fill_2 FILLER_5_181 ();
 sg13g2_fill_1 FILLER_5_183 ();
 sg13g2_fill_1 FILLER_5_202 ();
 sg13g2_fill_2 FILLER_5_208 ();
 sg13g2_fill_1 FILLER_5_210 ();
 sg13g2_fill_1 FILLER_5_216 ();
 sg13g2_decap_8 FILLER_5_274 ();
 sg13g2_decap_4 FILLER_5_281 ();
 sg13g2_fill_2 FILLER_5_285 ();
 sg13g2_fill_1 FILLER_5_295 ();
 sg13g2_fill_1 FILLER_5_314 ();
 sg13g2_decap_8 FILLER_5_320 ();
 sg13g2_decap_4 FILLER_5_337 ();
 sg13g2_fill_2 FILLER_5_341 ();
 sg13g2_fill_2 FILLER_5_347 ();
 sg13g2_fill_1 FILLER_5_349 ();
 sg13g2_decap_4 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_375 ();
 sg13g2_decap_8 FILLER_5_382 ();
 sg13g2_decap_8 FILLER_5_389 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_decap_4 FILLER_5_403 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_4 FILLER_6_161 ();
 sg13g2_fill_2 FILLER_6_165 ();
 sg13g2_fill_2 FILLER_6_183 ();
 sg13g2_fill_1 FILLER_6_185 ();
 sg13g2_fill_1 FILLER_6_222 ();
 sg13g2_decap_4 FILLER_6_229 ();
 sg13g2_fill_1 FILLER_6_233 ();
 sg13g2_decap_4 FILLER_6_246 ();
 sg13g2_decap_8 FILLER_6_254 ();
 sg13g2_fill_1 FILLER_6_271 ();
 sg13g2_decap_4 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_289 ();
 sg13g2_fill_2 FILLER_6_296 ();
 sg13g2_fill_1 FILLER_6_298 ();
 sg13g2_fill_2 FILLER_6_304 ();
 sg13g2_fill_1 FILLER_6_306 ();
 sg13g2_decap_4 FILLER_6_320 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_fill_1 FILLER_6_374 ();
 sg13g2_decap_8 FILLER_6_388 ();
 sg13g2_decap_8 FILLER_6_395 ();
 sg13g2_decap_8 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_4 FILLER_7_168 ();
 sg13g2_fill_2 FILLER_7_172 ();
 sg13g2_decap_8 FILLER_7_179 ();
 sg13g2_decap_8 FILLER_7_186 ();
 sg13g2_decap_4 FILLER_7_193 ();
 sg13g2_fill_1 FILLER_7_197 ();
 sg13g2_decap_8 FILLER_7_214 ();
 sg13g2_fill_2 FILLER_7_221 ();
 sg13g2_fill_1 FILLER_7_223 ();
 sg13g2_decap_4 FILLER_7_230 ();
 sg13g2_fill_2 FILLER_7_234 ();
 sg13g2_decap_8 FILLER_7_239 ();
 sg13g2_fill_2 FILLER_7_246 ();
 sg13g2_fill_1 FILLER_7_248 ();
 sg13g2_fill_2 FILLER_7_268 ();
 sg13g2_fill_1 FILLER_7_283 ();
 sg13g2_decap_4 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_354 ();
 sg13g2_fill_1 FILLER_7_361 ();
 sg13g2_fill_2 FILLER_7_372 ();
 sg13g2_fill_1 FILLER_7_374 ();
 sg13g2_decap_8 FILLER_7_387 ();
 sg13g2_decap_8 FILLER_7_394 ();
 sg13g2_decap_8 FILLER_7_401 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_4 FILLER_8_168 ();
 sg13g2_fill_2 FILLER_8_172 ();
 sg13g2_decap_8 FILLER_8_194 ();
 sg13g2_fill_1 FILLER_8_213 ();
 sg13g2_fill_1 FILLER_8_272 ();
 sg13g2_fill_1 FILLER_8_282 ();
 sg13g2_decap_8 FILLER_8_299 ();
 sg13g2_fill_1 FILLER_8_306 ();
 sg13g2_decap_8 FILLER_8_318 ();
 sg13g2_decap_4 FILLER_8_325 ();
 sg13g2_fill_1 FILLER_8_329 ();
 sg13g2_decap_4 FILLER_8_339 ();
 sg13g2_fill_1 FILLER_8_343 ();
 sg13g2_fill_1 FILLER_8_352 ();
 sg13g2_decap_4 FILLER_8_366 ();
 sg13g2_decap_4 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_decap_4 FILLER_8_404 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_fill_2 FILLER_9_161 ();
 sg13g2_fill_1 FILLER_9_163 ();
 sg13g2_fill_2 FILLER_9_180 ();
 sg13g2_fill_1 FILLER_9_182 ();
 sg13g2_fill_2 FILLER_9_195 ();
 sg13g2_fill_2 FILLER_9_209 ();
 sg13g2_decap_8 FILLER_9_222 ();
 sg13g2_decap_8 FILLER_9_235 ();
 sg13g2_decap_4 FILLER_9_242 ();
 sg13g2_fill_1 FILLER_9_246 ();
 sg13g2_fill_2 FILLER_9_256 ();
 sg13g2_fill_1 FILLER_9_258 ();
 sg13g2_fill_2 FILLER_9_267 ();
 sg13g2_decap_4 FILLER_9_291 ();
 sg13g2_fill_1 FILLER_9_295 ();
 sg13g2_decap_4 FILLER_9_304 ();
 sg13g2_fill_1 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_4 FILLER_10_161 ();
 sg13g2_fill_1 FILLER_10_165 ();
 sg13g2_fill_2 FILLER_10_169 ();
 sg13g2_fill_2 FILLER_10_181 ();
 sg13g2_fill_1 FILLER_10_193 ();
 sg13g2_fill_1 FILLER_10_200 ();
 sg13g2_fill_1 FILLER_10_206 ();
 sg13g2_fill_2 FILLER_10_211 ();
 sg13g2_fill_1 FILLER_10_213 ();
 sg13g2_decap_4 FILLER_10_226 ();
 sg13g2_fill_2 FILLER_10_275 ();
 sg13g2_fill_2 FILLER_10_289 ();
 sg13g2_fill_2 FILLER_10_304 ();
 sg13g2_fill_1 FILLER_10_306 ();
 sg13g2_fill_2 FILLER_10_315 ();
 sg13g2_fill_1 FILLER_10_322 ();
 sg13g2_decap_4 FILLER_10_332 ();
 sg13g2_fill_1 FILLER_10_336 ();
 sg13g2_fill_2 FILLER_10_353 ();
 sg13g2_fill_1 FILLER_10_355 ();
 sg13g2_fill_2 FILLER_10_360 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_fill_2 FILLER_11_161 ();
 sg13g2_fill_1 FILLER_11_184 ();
 sg13g2_decap_4 FILLER_11_246 ();
 sg13g2_decap_4 FILLER_11_263 ();
 sg13g2_fill_2 FILLER_11_267 ();
 sg13g2_decap_8 FILLER_11_277 ();
 sg13g2_fill_1 FILLER_11_284 ();
 sg13g2_fill_1 FILLER_11_299 ();
 sg13g2_fill_2 FILLER_11_312 ();
 sg13g2_fill_1 FILLER_11_314 ();
 sg13g2_decap_8 FILLER_11_338 ();
 sg13g2_decap_4 FILLER_11_345 ();
 sg13g2_fill_2 FILLER_11_349 ();
 sg13g2_decap_4 FILLER_11_359 ();
 sg13g2_fill_1 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_fill_2 FILLER_12_161 ();
 sg13g2_fill_1 FILLER_12_163 ();
 sg13g2_fill_2 FILLER_12_169 ();
 sg13g2_fill_2 FILLER_12_180 ();
 sg13g2_decap_8 FILLER_12_190 ();
 sg13g2_fill_2 FILLER_12_197 ();
 sg13g2_decap_4 FILLER_12_204 ();
 sg13g2_fill_2 FILLER_12_208 ();
 sg13g2_fill_2 FILLER_12_214 ();
 sg13g2_fill_1 FILLER_12_216 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_fill_2 FILLER_12_238 ();
 sg13g2_fill_1 FILLER_12_255 ();
 sg13g2_fill_1 FILLER_12_276 ();
 sg13g2_fill_1 FILLER_12_296 ();
 sg13g2_fill_1 FILLER_12_322 ();
 sg13g2_fill_2 FILLER_12_329 ();
 sg13g2_fill_1 FILLER_12_331 ();
 sg13g2_fill_1 FILLER_12_340 ();
 sg13g2_fill_1 FILLER_12_359 ();
 sg13g2_fill_2 FILLER_12_369 ();
 sg13g2_fill_1 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_380 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_fill_1 FILLER_13_161 ();
 sg13g2_fill_2 FILLER_13_170 ();
 sg13g2_fill_2 FILLER_13_180 ();
 sg13g2_decap_4 FILLER_13_192 ();
 sg13g2_fill_2 FILLER_13_196 ();
 sg13g2_fill_2 FILLER_13_203 ();
 sg13g2_fill_1 FILLER_13_216 ();
 sg13g2_fill_1 FILLER_13_223 ();
 sg13g2_decap_8 FILLER_13_277 ();
 sg13g2_fill_2 FILLER_13_284 ();
 sg13g2_fill_1 FILLER_13_286 ();
 sg13g2_fill_1 FILLER_13_295 ();
 sg13g2_fill_2 FILLER_13_304 ();
 sg13g2_fill_1 FILLER_13_306 ();
 sg13g2_fill_2 FILLER_13_324 ();
 sg13g2_fill_1 FILLER_13_336 ();
 sg13g2_fill_2 FILLER_13_351 ();
 sg13g2_fill_1 FILLER_13_363 ();
 sg13g2_decap_4 FILLER_13_369 ();
 sg13g2_fill_1 FILLER_13_373 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_decap_8 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_fill_2 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_216 ();
 sg13g2_fill_2 FILLER_14_223 ();
 sg13g2_decap_8 FILLER_14_237 ();
 sg13g2_decap_8 FILLER_14_244 ();
 sg13g2_decap_4 FILLER_14_251 ();
 sg13g2_decap_4 FILLER_14_272 ();
 sg13g2_fill_2 FILLER_14_276 ();
 sg13g2_fill_1 FILLER_14_318 ();
 sg13g2_fill_2 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_4 FILLER_15_154 ();
 sg13g2_fill_2 FILLER_15_158 ();
 sg13g2_fill_2 FILLER_15_173 ();
 sg13g2_fill_1 FILLER_15_175 ();
 sg13g2_decap_4 FILLER_15_193 ();
 sg13g2_fill_2 FILLER_15_197 ();
 sg13g2_fill_2 FILLER_15_203 ();
 sg13g2_fill_1 FILLER_15_222 ();
 sg13g2_fill_1 FILLER_15_231 ();
 sg13g2_fill_2 FILLER_15_244 ();
 sg13g2_fill_1 FILLER_15_246 ();
 sg13g2_decap_4 FILLER_15_268 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_fill_2 FILLER_15_287 ();
 sg13g2_fill_2 FILLER_15_297 ();
 sg13g2_fill_2 FILLER_15_308 ();
 sg13g2_fill_1 FILLER_15_310 ();
 sg13g2_fill_1 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_324 ();
 sg13g2_decap_8 FILLER_15_331 ();
 sg13g2_fill_1 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_4 FILLER_16_154 ();
 sg13g2_fill_1 FILLER_16_158 ();
 sg13g2_decap_8 FILLER_16_166 ();
 sg13g2_fill_1 FILLER_16_173 ();
 sg13g2_decap_8 FILLER_16_179 ();
 sg13g2_decap_8 FILLER_16_186 ();
 sg13g2_decap_4 FILLER_16_193 ();
 sg13g2_fill_1 FILLER_16_197 ();
 sg13g2_decap_4 FILLER_16_208 ();
 sg13g2_fill_1 FILLER_16_212 ();
 sg13g2_fill_1 FILLER_16_221 ();
 sg13g2_fill_2 FILLER_16_254 ();
 sg13g2_fill_2 FILLER_16_260 ();
 sg13g2_fill_1 FILLER_16_262 ();
 sg13g2_decap_8 FILLER_16_271 ();
 sg13g2_decap_4 FILLER_16_310 ();
 sg13g2_fill_2 FILLER_16_314 ();
 sg13g2_decap_4 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_fill_2 FILLER_17_147 ();
 sg13g2_fill_1 FILLER_17_149 ();
 sg13g2_fill_2 FILLER_17_163 ();
 sg13g2_decap_4 FILLER_17_176 ();
 sg13g2_fill_1 FILLER_17_206 ();
 sg13g2_fill_2 FILLER_17_219 ();
 sg13g2_fill_1 FILLER_17_221 ();
 sg13g2_decap_4 FILLER_17_228 ();
 sg13g2_decap_4 FILLER_17_238 ();
 sg13g2_fill_1 FILLER_17_242 ();
 sg13g2_fill_2 FILLER_17_251 ();
 sg13g2_fill_1 FILLER_17_253 ();
 sg13g2_fill_1 FILLER_17_262 ();
 sg13g2_fill_1 FILLER_17_297 ();
 sg13g2_decap_8 FILLER_17_330 ();
 sg13g2_fill_1 FILLER_17_337 ();
 sg13g2_fill_2 FILLER_17_343 ();
 sg13g2_fill_1 FILLER_17_345 ();
 sg13g2_decap_8 FILLER_17_351 ();
 sg13g2_decap_4 FILLER_17_358 ();
 sg13g2_fill_2 FILLER_17_362 ();
 sg13g2_fill_1 FILLER_17_372 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_4 FILLER_18_166 ();
 sg13g2_decap_4 FILLER_18_190 ();
 sg13g2_fill_1 FILLER_18_194 ();
 sg13g2_decap_4 FILLER_18_199 ();
 sg13g2_fill_1 FILLER_18_203 ();
 sg13g2_decap_4 FILLER_18_243 ();
 sg13g2_fill_2 FILLER_18_253 ();
 sg13g2_fill_1 FILLER_18_255 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_fill_1 FILLER_18_284 ();
 sg13g2_decap_8 FILLER_18_304 ();
 sg13g2_decap_4 FILLER_18_311 ();
 sg13g2_fill_1 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_320 ();
 sg13g2_fill_1 FILLER_18_327 ();
 sg13g2_fill_2 FILLER_18_352 ();
 sg13g2_fill_1 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_18_389 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_fill_2 FILLER_19_147 ();
 sg13g2_fill_2 FILLER_19_158 ();
 sg13g2_fill_1 FILLER_19_160 ();
 sg13g2_decap_8 FILLER_19_166 ();
 sg13g2_decap_4 FILLER_19_178 ();
 sg13g2_fill_2 FILLER_19_182 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_207 ();
 sg13g2_decap_8 FILLER_19_214 ();
 sg13g2_decap_8 FILLER_19_239 ();
 sg13g2_fill_2 FILLER_19_267 ();
 sg13g2_fill_1 FILLER_19_269 ();
 sg13g2_decap_8 FILLER_19_286 ();
 sg13g2_decap_8 FILLER_19_293 ();
 sg13g2_fill_1 FILLER_19_300 ();
 sg13g2_fill_2 FILLER_19_314 ();
 sg13g2_fill_2 FILLER_19_321 ();
 sg13g2_fill_2 FILLER_19_334 ();
 sg13g2_fill_1 FILLER_19_336 ();
 sg13g2_fill_2 FILLER_19_342 ();
 sg13g2_fill_1 FILLER_19_344 ();
 sg13g2_decap_4 FILLER_19_371 ();
 sg13g2_fill_2 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_4 FILLER_20_140 ();
 sg13g2_fill_1 FILLER_20_144 ();
 sg13g2_decap_4 FILLER_20_150 ();
 sg13g2_fill_2 FILLER_20_154 ();
 sg13g2_fill_2 FILLER_20_168 ();
 sg13g2_fill_2 FILLER_20_201 ();
 sg13g2_fill_1 FILLER_20_203 ();
 sg13g2_fill_1 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_243 ();
 sg13g2_fill_2 FILLER_20_250 ();
 sg13g2_fill_1 FILLER_20_289 ();
 sg13g2_fill_1 FILLER_20_307 ();
 sg13g2_decap_4 FILLER_20_313 ();
 sg13g2_fill_2 FILLER_20_331 ();
 sg13g2_fill_1 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_348 ();
 sg13g2_decap_8 FILLER_20_355 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_381 ();
 sg13g2_decap_8 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_4 FILLER_21_133 ();
 sg13g2_fill_2 FILLER_21_137 ();
 sg13g2_decap_8 FILLER_21_184 ();
 sg13g2_fill_2 FILLER_21_191 ();
 sg13g2_decap_4 FILLER_21_214 ();
 sg13g2_fill_1 FILLER_21_218 ();
 sg13g2_fill_2 FILLER_21_224 ();
 sg13g2_fill_1 FILLER_21_226 ();
 sg13g2_fill_1 FILLER_21_232 ();
 sg13g2_fill_1 FILLER_21_264 ();
 sg13g2_decap_4 FILLER_21_275 ();
 sg13g2_fill_1 FILLER_21_300 ();
 sg13g2_fill_1 FILLER_21_340 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_4 FILLER_22_154 ();
 sg13g2_fill_2 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_208 ();
 sg13g2_fill_1 FILLER_22_214 ();
 sg13g2_fill_2 FILLER_22_226 ();
 sg13g2_decap_4 FILLER_22_238 ();
 sg13g2_fill_2 FILLER_22_242 ();
 sg13g2_fill_2 FILLER_22_250 ();
 sg13g2_fill_1 FILLER_22_252 ();
 sg13g2_fill_1 FILLER_22_269 ();
 sg13g2_fill_2 FILLER_22_278 ();
 sg13g2_fill_2 FILLER_22_294 ();
 sg13g2_decap_4 FILLER_22_304 ();
 sg13g2_fill_1 FILLER_22_313 ();
 sg13g2_fill_1 FILLER_22_320 ();
 sg13g2_fill_2 FILLER_22_325 ();
 sg13g2_decap_4 FILLER_22_342 ();
 sg13g2_fill_2 FILLER_22_346 ();
 sg13g2_decap_8 FILLER_22_354 ();
 sg13g2_fill_1 FILLER_22_361 ();
 sg13g2_decap_4 FILLER_22_371 ();
 sg13g2_decap_4 FILLER_22_387 ();
 sg13g2_fill_2 FILLER_22_391 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_fill_2 FILLER_23_147 ();
 sg13g2_fill_1 FILLER_23_149 ();
 sg13g2_fill_2 FILLER_23_168 ();
 sg13g2_fill_2 FILLER_23_175 ();
 sg13g2_fill_1 FILLER_23_177 ();
 sg13g2_fill_1 FILLER_23_182 ();
 sg13g2_fill_1 FILLER_23_213 ();
 sg13g2_fill_1 FILLER_23_223 ();
 sg13g2_fill_1 FILLER_23_238 ();
 sg13g2_fill_2 FILLER_23_256 ();
 sg13g2_fill_1 FILLER_23_258 ();
 sg13g2_fill_1 FILLER_23_272 ();
 sg13g2_fill_2 FILLER_23_284 ();
 sg13g2_fill_1 FILLER_23_286 ();
 sg13g2_fill_2 FILLER_23_295 ();
 sg13g2_fill_1 FILLER_23_297 ();
 sg13g2_fill_2 FILLER_23_309 ();
 sg13g2_fill_1 FILLER_23_311 ();
 sg13g2_fill_2 FILLER_23_335 ();
 sg13g2_fill_1 FILLER_23_353 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_147 ();
 sg13g2_fill_2 FILLER_24_174 ();
 sg13g2_fill_1 FILLER_24_176 ();
 sg13g2_fill_2 FILLER_24_191 ();
 sg13g2_fill_1 FILLER_24_193 ();
 sg13g2_fill_2 FILLER_24_216 ();
 sg13g2_decap_8 FILLER_24_228 ();
 sg13g2_fill_1 FILLER_24_235 ();
 sg13g2_decap_8 FILLER_24_242 ();
 sg13g2_fill_2 FILLER_24_249 ();
 sg13g2_fill_1 FILLER_24_251 ();
 sg13g2_decap_8 FILLER_24_262 ();
 sg13g2_decap_4 FILLER_24_278 ();
 sg13g2_fill_2 FILLER_24_282 ();
 sg13g2_fill_2 FILLER_24_290 ();
 sg13g2_fill_1 FILLER_24_292 ();
 sg13g2_decap_8 FILLER_24_297 ();
 sg13g2_decap_4 FILLER_24_304 ();
 sg13g2_fill_1 FILLER_24_308 ();
 sg13g2_fill_1 FILLER_24_317 ();
 sg13g2_decap_8 FILLER_24_326 ();
 sg13g2_decap_4 FILLER_24_333 ();
 sg13g2_fill_2 FILLER_24_357 ();
 sg13g2_decap_4 FILLER_24_368 ();
 sg13g2_fill_2 FILLER_24_372 ();
 sg13g2_decap_4 FILLER_24_380 ();
 sg13g2_fill_2 FILLER_24_388 ();
 sg13g2_fill_2 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_fill_2 FILLER_25_147 ();
 sg13g2_decap_4 FILLER_25_154 ();
 sg13g2_fill_1 FILLER_25_158 ();
 sg13g2_fill_2 FILLER_25_185 ();
 sg13g2_fill_1 FILLER_25_187 ();
 sg13g2_decap_4 FILLER_25_202 ();
 sg13g2_fill_2 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_215 ();
 sg13g2_fill_2 FILLER_25_243 ();
 sg13g2_fill_1 FILLER_25_245 ();
 sg13g2_fill_2 FILLER_25_253 ();
 sg13g2_fill_1 FILLER_25_255 ();
 sg13g2_fill_2 FILLER_25_261 ();
 sg13g2_fill_1 FILLER_25_274 ();
 sg13g2_fill_1 FILLER_25_292 ();
 sg13g2_decap_4 FILLER_25_319 ();
 sg13g2_decap_8 FILLER_25_335 ();
 sg13g2_decap_4 FILLER_25_345 ();
 sg13g2_fill_1 FILLER_25_349 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_4 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_120 ();
 sg13g2_decap_8 FILLER_26_127 ();
 sg13g2_decap_8 FILLER_26_134 ();
 sg13g2_fill_2 FILLER_26_147 ();
 sg13g2_fill_2 FILLER_26_175 ();
 sg13g2_fill_1 FILLER_26_177 ();
 sg13g2_fill_1 FILLER_26_192 ();
 sg13g2_fill_2 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_207 ();
 sg13g2_fill_2 FILLER_26_218 ();
 sg13g2_fill_1 FILLER_26_220 ();
 sg13g2_fill_2 FILLER_26_233 ();
 sg13g2_fill_2 FILLER_26_240 ();
 sg13g2_fill_1 FILLER_26_242 ();
 sg13g2_fill_1 FILLER_26_248 ();
 sg13g2_fill_2 FILLER_26_255 ();
 sg13g2_fill_1 FILLER_26_280 ();
 sg13g2_decap_4 FILLER_26_285 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_fill_1 FILLER_26_303 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_4 FILLER_26_322 ();
 sg13g2_fill_1 FILLER_26_326 ();
 sg13g2_fill_2 FILLER_26_333 ();
 sg13g2_fill_1 FILLER_26_335 ();
 sg13g2_decap_4 FILLER_26_350 ();
 sg13g2_fill_1 FILLER_26_354 ();
 sg13g2_fill_2 FILLER_26_363 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_376 ();
 sg13g2_decap_4 FILLER_26_383 ();
 sg13g2_fill_2 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_4 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_93 ();
 sg13g2_decap_4 FILLER_27_100 ();
 sg13g2_decap_8 FILLER_27_130 ();
 sg13g2_fill_1 FILLER_27_141 ();
 sg13g2_fill_2 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_149 ();
 sg13g2_fill_1 FILLER_27_160 ();
 sg13g2_fill_2 FILLER_27_172 ();
 sg13g2_fill_1 FILLER_27_174 ();
 sg13g2_fill_2 FILLER_27_188 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_fill_2 FILLER_27_203 ();
 sg13g2_fill_1 FILLER_27_210 ();
 sg13g2_fill_1 FILLER_27_216 ();
 sg13g2_fill_1 FILLER_27_225 ();
 sg13g2_fill_2 FILLER_27_230 ();
 sg13g2_fill_2 FILLER_27_247 ();
 sg13g2_fill_1 FILLER_27_254 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_fill_1 FILLER_27_262 ();
 sg13g2_fill_1 FILLER_27_285 ();
 sg13g2_fill_2 FILLER_27_294 ();
 sg13g2_fill_1 FILLER_27_332 ();
 sg13g2_fill_2 FILLER_27_358 ();
 sg13g2_fill_1 FILLER_27_360 ();
 sg13g2_decap_4 FILLER_27_382 ();
 sg13g2_fill_1 FILLER_27_386 ();
 sg13g2_fill_1 FILLER_27_392 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_fill_2 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_77 ();
 sg13g2_fill_2 FILLER_28_96 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_decap_4 FILLER_28_108 ();
 sg13g2_decap_4 FILLER_28_121 ();
 sg13g2_fill_2 FILLER_28_140 ();
 sg13g2_fill_2 FILLER_28_161 ();
 sg13g2_fill_1 FILLER_28_163 ();
 sg13g2_fill_1 FILLER_28_178 ();
 sg13g2_fill_1 FILLER_28_212 ();
 sg13g2_fill_2 FILLER_28_218 ();
 sg13g2_fill_1 FILLER_28_220 ();
 sg13g2_fill_1 FILLER_28_232 ();
 sg13g2_fill_1 FILLER_28_248 ();
 sg13g2_decap_4 FILLER_28_264 ();
 sg13g2_fill_2 FILLER_28_268 ();
 sg13g2_decap_4 FILLER_28_274 ();
 sg13g2_fill_1 FILLER_28_278 ();
 sg13g2_fill_2 FILLER_28_305 ();
 sg13g2_fill_2 FILLER_28_326 ();
 sg13g2_fill_1 FILLER_28_344 ();
 sg13g2_decap_4 FILLER_28_366 ();
 sg13g2_fill_2 FILLER_28_375 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_fill_1 FILLER_29_56 ();
 sg13g2_fill_2 FILLER_29_63 ();
 sg13g2_fill_1 FILLER_29_70 ();
 sg13g2_fill_2 FILLER_29_80 ();
 sg13g2_fill_2 FILLER_29_89 ();
 sg13g2_fill_2 FILLER_29_102 ();
 sg13g2_fill_1 FILLER_29_104 ();
 sg13g2_fill_2 FILLER_29_115 ();
 sg13g2_fill_1 FILLER_29_127 ();
 sg13g2_fill_1 FILLER_29_139 ();
 sg13g2_decap_8 FILLER_29_144 ();
 sg13g2_decap_8 FILLER_29_151 ();
 sg13g2_decap_4 FILLER_29_167 ();
 sg13g2_decap_8 FILLER_29_185 ();
 sg13g2_decap_8 FILLER_29_208 ();
 sg13g2_fill_1 FILLER_29_219 ();
 sg13g2_fill_1 FILLER_29_228 ();
 sg13g2_fill_1 FILLER_29_238 ();
 sg13g2_fill_2 FILLER_29_244 ();
 sg13g2_fill_1 FILLER_29_246 ();
 sg13g2_fill_2 FILLER_29_255 ();
 sg13g2_fill_1 FILLER_29_270 ();
 sg13g2_decap_4 FILLER_29_276 ();
 sg13g2_fill_2 FILLER_29_288 ();
 sg13g2_decap_4 FILLER_29_316 ();
 sg13g2_fill_1 FILLER_29_365 ();
 sg13g2_fill_1 FILLER_29_374 ();
 sg13g2_decap_4 FILLER_29_383 ();
 sg13g2_fill_1 FILLER_29_387 ();
 sg13g2_fill_2 FILLER_29_397 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_4 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_67 ();
 sg13g2_decap_8 FILLER_30_83 ();
 sg13g2_fill_2 FILLER_30_90 ();
 sg13g2_fill_1 FILLER_30_92 ();
 sg13g2_fill_2 FILLER_30_102 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_fill_1 FILLER_30_110 ();
 sg13g2_fill_2 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_172 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_fill_2 FILLER_30_220 ();
 sg13g2_fill_1 FILLER_30_227 ();
 sg13g2_decap_8 FILLER_30_247 ();
 sg13g2_fill_2 FILLER_30_254 ();
 sg13g2_fill_1 FILLER_30_256 ();
 sg13g2_decap_8 FILLER_30_286 ();
 sg13g2_fill_1 FILLER_30_293 ();
 sg13g2_decap_4 FILLER_30_301 ();
 sg13g2_fill_2 FILLER_30_305 ();
 sg13g2_fill_2 FILLER_30_311 ();
 sg13g2_fill_1 FILLER_30_313 ();
 sg13g2_fill_2 FILLER_30_322 ();
 sg13g2_fill_1 FILLER_30_324 ();
 sg13g2_fill_1 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_334 ();
 sg13g2_decap_8 FILLER_30_341 ();
 sg13g2_fill_1 FILLER_30_348 ();
 sg13g2_decap_4 FILLER_30_357 ();
 sg13g2_fill_2 FILLER_30_361 ();
 sg13g2_decap_8 FILLER_30_368 ();
 sg13g2_fill_2 FILLER_30_375 ();
 sg13g2_fill_1 FILLER_30_377 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_4 FILLER_31_42 ();
 sg13g2_fill_2 FILLER_31_46 ();
 sg13g2_fill_2 FILLER_31_57 ();
 sg13g2_fill_1 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_87 ();
 sg13g2_fill_2 FILLER_31_93 ();
 sg13g2_fill_1 FILLER_31_108 ();
 sg13g2_decap_8 FILLER_31_115 ();
 sg13g2_decap_4 FILLER_31_122 ();
 sg13g2_fill_2 FILLER_31_126 ();
 sg13g2_decap_4 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_147 ();
 sg13g2_fill_2 FILLER_31_153 ();
 sg13g2_fill_1 FILLER_31_155 ();
 sg13g2_decap_8 FILLER_31_162 ();
 sg13g2_decap_4 FILLER_31_169 ();
 sg13g2_fill_2 FILLER_31_178 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_4 FILLER_31_212 ();
 sg13g2_fill_1 FILLER_31_216 ();
 sg13g2_fill_2 FILLER_31_237 ();
 sg13g2_fill_2 FILLER_31_261 ();
 sg13g2_decap_8 FILLER_31_268 ();
 sg13g2_fill_2 FILLER_31_275 ();
 sg13g2_fill_1 FILLER_31_277 ();
 sg13g2_fill_2 FILLER_31_294 ();
 sg13g2_fill_1 FILLER_31_322 ();
 sg13g2_fill_1 FILLER_31_346 ();
 sg13g2_fill_1 FILLER_31_352 ();
 sg13g2_fill_2 FILLER_31_362 ();
 sg13g2_fill_1 FILLER_31_398 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_fill_2 FILLER_32_49 ();
 sg13g2_fill_1 FILLER_32_51 ();
 sg13g2_fill_2 FILLER_32_60 ();
 sg13g2_fill_1 FILLER_32_62 ();
 sg13g2_fill_2 FILLER_32_68 ();
 sg13g2_fill_1 FILLER_32_70 ();
 sg13g2_fill_2 FILLER_32_81 ();
 sg13g2_fill_2 FILLER_32_87 ();
 sg13g2_fill_2 FILLER_32_99 ();
 sg13g2_fill_1 FILLER_32_105 ();
 sg13g2_fill_2 FILLER_32_114 ();
 sg13g2_fill_1 FILLER_32_126 ();
 sg13g2_decap_4 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_158 ();
 sg13g2_fill_2 FILLER_32_169 ();
 sg13g2_fill_2 FILLER_32_182 ();
 sg13g2_fill_1 FILLER_32_184 ();
 sg13g2_fill_2 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_209 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_fill_1 FILLER_32_224 ();
 sg13g2_decap_4 FILLER_32_241 ();
 sg13g2_fill_2 FILLER_32_288 ();
 sg13g2_decap_4 FILLER_32_301 ();
 sg13g2_fill_1 FILLER_32_305 ();
 sg13g2_fill_1 FILLER_32_312 ();
 sg13g2_decap_4 FILLER_32_321 ();
 sg13g2_decap_4 FILLER_32_334 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_fill_2 FILLER_32_345 ();
 sg13g2_fill_2 FILLER_32_377 ();
 sg13g2_fill_2 FILLER_32_393 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_fill_2 FILLER_33_49 ();
 sg13g2_fill_2 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_58 ();
 sg13g2_fill_1 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_93 ();
 sg13g2_fill_2 FILLER_33_113 ();
 sg13g2_fill_1 FILLER_33_115 ();
 sg13g2_fill_2 FILLER_33_137 ();
 sg13g2_fill_1 FILLER_33_139 ();
 sg13g2_fill_1 FILLER_33_154 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_fill_2 FILLER_33_176 ();
 sg13g2_fill_1 FILLER_33_178 ();
 sg13g2_fill_1 FILLER_33_192 ();
 sg13g2_decap_4 FILLER_33_197 ();
 sg13g2_fill_1 FILLER_33_201 ();
 sg13g2_fill_1 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_232 ();
 sg13g2_decap_4 FILLER_33_257 ();
 sg13g2_fill_2 FILLER_33_261 ();
 sg13g2_decap_8 FILLER_33_267 ();
 sg13g2_decap_8 FILLER_33_274 ();
 sg13g2_decap_4 FILLER_33_309 ();
 sg13g2_fill_1 FILLER_33_313 ();
 sg13g2_fill_2 FILLER_33_320 ();
 sg13g2_fill_1 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_335 ();
 sg13g2_fill_2 FILLER_33_342 ();
 sg13g2_fill_1 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_349 ();
 sg13g2_decap_4 FILLER_33_361 ();
 sg13g2_fill_1 FILLER_33_365 ();
 sg13g2_fill_2 FILLER_33_383 ();
 sg13g2_decap_4 FILLER_33_393 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_fill_2 FILLER_34_49 ();
 sg13g2_fill_1 FILLER_34_51 ();
 sg13g2_fill_2 FILLER_34_65 ();
 sg13g2_fill_1 FILLER_34_67 ();
 sg13g2_fill_1 FILLER_34_82 ();
 sg13g2_decap_4 FILLER_34_88 ();
 sg13g2_fill_2 FILLER_34_92 ();
 sg13g2_fill_2 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_116 ();
 sg13g2_decap_8 FILLER_34_123 ();
 sg13g2_fill_2 FILLER_34_130 ();
 sg13g2_fill_1 FILLER_34_149 ();
 sg13g2_fill_2 FILLER_34_155 ();
 sg13g2_fill_2 FILLER_34_187 ();
 sg13g2_fill_2 FILLER_34_194 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_fill_1 FILLER_34_205 ();
 sg13g2_decap_8 FILLER_34_211 ();
 sg13g2_decap_4 FILLER_34_218 ();
 sg13g2_fill_2 FILLER_34_222 ();
 sg13g2_decap_8 FILLER_34_235 ();
 sg13g2_decap_8 FILLER_34_242 ();
 sg13g2_decap_4 FILLER_34_249 ();
 sg13g2_fill_1 FILLER_34_253 ();
 sg13g2_fill_1 FILLER_34_293 ();
 sg13g2_decap_4 FILLER_34_299 ();
 sg13g2_decap_8 FILLER_34_319 ();
 sg13g2_fill_2 FILLER_34_326 ();
 sg13g2_decap_8 FILLER_34_374 ();
 sg13g2_decap_8 FILLER_34_381 ();
 sg13g2_fill_1 FILLER_34_388 ();
 sg13g2_fill_2 FILLER_34_397 ();
 sg13g2_fill_1 FILLER_34_399 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_4 FILLER_35_42 ();
 sg13g2_fill_1 FILLER_35_46 ();
 sg13g2_fill_1 FILLER_35_61 ();
 sg13g2_fill_1 FILLER_35_69 ();
 sg13g2_fill_2 FILLER_35_92 ();
 sg13g2_fill_1 FILLER_35_94 ();
 sg13g2_fill_1 FILLER_35_136 ();
 sg13g2_fill_2 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_163 ();
 sg13g2_decap_8 FILLER_35_173 ();
 sg13g2_fill_1 FILLER_35_184 ();
 sg13g2_fill_2 FILLER_35_195 ();
 sg13g2_fill_2 FILLER_35_213 ();
 sg13g2_decap_4 FILLER_35_223 ();
 sg13g2_fill_1 FILLER_35_238 ();
 sg13g2_fill_2 FILLER_35_279 ();
 sg13g2_fill_2 FILLER_35_299 ();
 sg13g2_fill_2 FILLER_35_309 ();
 sg13g2_decap_8 FILLER_35_341 ();
 sg13g2_fill_1 FILLER_35_348 ();
 sg13g2_fill_1 FILLER_35_366 ();
 sg13g2_fill_2 FILLER_35_375 ();
 sg13g2_fill_1 FILLER_35_377 ();
 sg13g2_fill_1 FILLER_35_390 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_fill_2 FILLER_36_56 ();
 sg13g2_decap_4 FILLER_36_63 ();
 sg13g2_fill_2 FILLER_36_67 ();
 sg13g2_fill_1 FILLER_36_74 ();
 sg13g2_decap_8 FILLER_36_80 ();
 sg13g2_decap_4 FILLER_36_87 ();
 sg13g2_fill_2 FILLER_36_91 ();
 sg13g2_fill_1 FILLER_36_108 ();
 sg13g2_decap_4 FILLER_36_117 ();
 sg13g2_fill_2 FILLER_36_121 ();
 sg13g2_fill_1 FILLER_36_128 ();
 sg13g2_decap_4 FILLER_36_134 ();
 sg13g2_fill_1 FILLER_36_138 ();
 sg13g2_fill_2 FILLER_36_151 ();
 sg13g2_fill_1 FILLER_36_153 ();
 sg13g2_fill_2 FILLER_36_159 ();
 sg13g2_fill_1 FILLER_36_161 ();
 sg13g2_fill_2 FILLER_36_187 ();
 sg13g2_fill_1 FILLER_36_189 ();
 sg13g2_fill_1 FILLER_36_198 ();
 sg13g2_decap_8 FILLER_36_204 ();
 sg13g2_decap_4 FILLER_36_211 ();
 sg13g2_fill_1 FILLER_36_215 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_fill_1 FILLER_36_227 ();
 sg13g2_fill_2 FILLER_36_238 ();
 sg13g2_fill_2 FILLER_36_257 ();
 sg13g2_fill_1 FILLER_36_259 ();
 sg13g2_fill_2 FILLER_36_270 ();
 sg13g2_fill_2 FILLER_36_290 ();
 sg13g2_fill_1 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_307 ();
 sg13g2_decap_8 FILLER_36_314 ();
 sg13g2_decap_4 FILLER_36_321 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_fill_1 FILLER_36_346 ();
 sg13g2_fill_2 FILLER_36_352 ();
 sg13g2_fill_1 FILLER_36_354 ();
 sg13g2_fill_2 FILLER_36_367 ();
 sg13g2_fill_1 FILLER_36_369 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_fill_2 FILLER_37_42 ();
 sg13g2_fill_1 FILLER_37_44 ();
 sg13g2_decap_4 FILLER_37_61 ();
 sg13g2_fill_2 FILLER_37_85 ();
 sg13g2_fill_1 FILLER_37_87 ();
 sg13g2_fill_2 FILLER_37_93 ();
 sg13g2_fill_1 FILLER_37_95 ();
 sg13g2_fill_2 FILLER_37_111 ();
 sg13g2_fill_1 FILLER_37_113 ();
 sg13g2_fill_1 FILLER_37_119 ();
 sg13g2_fill_2 FILLER_37_126 ();
 sg13g2_fill_1 FILLER_37_133 ();
 sg13g2_fill_2 FILLER_37_140 ();
 sg13g2_fill_2 FILLER_37_152 ();
 sg13g2_fill_1 FILLER_37_170 ();
 sg13g2_fill_2 FILLER_37_195 ();
 sg13g2_fill_1 FILLER_37_197 ();
 sg13g2_fill_1 FILLER_37_222 ();
 sg13g2_fill_2 FILLER_37_233 ();
 sg13g2_fill_1 FILLER_37_274 ();
 sg13g2_decap_4 FILLER_37_303 ();
 sg13g2_fill_1 FILLER_37_307 ();
 sg13g2_fill_2 FILLER_37_337 ();
 sg13g2_fill_1 FILLER_37_339 ();
 sg13g2_fill_2 FILLER_37_344 ();
 sg13g2_fill_1 FILLER_37_346 ();
 sg13g2_decap_4 FILLER_37_375 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_59 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_fill_1 FILLER_38_80 ();
 sg13g2_fill_2 FILLER_38_101 ();
 sg13g2_fill_1 FILLER_38_103 ();
 sg13g2_fill_1 FILLER_38_110 ();
 sg13g2_decap_4 FILLER_38_115 ();
 sg13g2_fill_2 FILLER_38_125 ();
 sg13g2_fill_1 FILLER_38_127 ();
 sg13g2_fill_1 FILLER_38_142 ();
 sg13g2_fill_1 FILLER_38_161 ();
 sg13g2_fill_2 FILLER_38_170 ();
 sg13g2_decap_8 FILLER_38_178 ();
 sg13g2_decap_4 FILLER_38_185 ();
 sg13g2_fill_1 FILLER_38_189 ();
 sg13g2_fill_2 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_205 ();
 sg13g2_fill_2 FILLER_38_212 ();
 sg13g2_fill_1 FILLER_38_214 ();
 sg13g2_decap_4 FILLER_38_219 ();
 sg13g2_fill_2 FILLER_38_232 ();
 sg13g2_fill_1 FILLER_38_234 ();
 sg13g2_decap_4 FILLER_38_249 ();
 sg13g2_fill_2 FILLER_38_258 ();
 sg13g2_fill_2 FILLER_38_269 ();
 sg13g2_decap_8 FILLER_38_276 ();
 sg13g2_fill_2 FILLER_38_283 ();
 sg13g2_decap_4 FILLER_38_290 ();
 sg13g2_fill_1 FILLER_38_294 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_decap_4 FILLER_38_342 ();
 sg13g2_fill_2 FILLER_38_346 ();
 sg13g2_fill_1 FILLER_38_354 ();
 sg13g2_decap_8 FILLER_38_360 ();
 sg13g2_decap_4 FILLER_38_367 ();
 sg13g2_fill_1 FILLER_38_371 ();
 sg13g2_fill_1 FILLER_38_380 ();
 sg13g2_fill_2 FILLER_38_393 ();
 sg13g2_fill_1 FILLER_38_395 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_fill_2 FILLER_39_49 ();
 sg13g2_fill_2 FILLER_39_90 ();
 sg13g2_fill_1 FILLER_39_121 ();
 sg13g2_fill_2 FILLER_39_130 ();
 sg13g2_fill_2 FILLER_39_155 ();
 sg13g2_fill_1 FILLER_39_157 ();
 sg13g2_decap_8 FILLER_39_162 ();
 sg13g2_decap_4 FILLER_39_177 ();
 sg13g2_fill_2 FILLER_39_190 ();
 sg13g2_fill_2 FILLER_39_195 ();
 sg13g2_fill_1 FILLER_39_203 ();
 sg13g2_fill_2 FILLER_39_238 ();
 sg13g2_fill_1 FILLER_39_240 ();
 sg13g2_fill_2 FILLER_39_274 ();
 sg13g2_fill_1 FILLER_39_276 ();
 sg13g2_decap_8 FILLER_39_296 ();
 sg13g2_decap_4 FILLER_39_303 ();
 sg13g2_fill_2 FILLER_39_307 ();
 sg13g2_fill_2 FILLER_39_316 ();
 sg13g2_fill_1 FILLER_39_331 ();
 sg13g2_decap_4 FILLER_39_352 ();
 sg13g2_fill_1 FILLER_39_356 ();
 sg13g2_decap_4 FILLER_39_365 ();
 sg13g2_fill_2 FILLER_39_377 ();
 sg13g2_fill_1 FILLER_39_379 ();
 sg13g2_fill_2 FILLER_39_388 ();
 sg13g2_fill_1 FILLER_39_397 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_4 FILLER_40_35 ();
 sg13g2_fill_1 FILLER_40_39 ();
 sg13g2_decap_8 FILLER_40_48 ();
 sg13g2_decap_8 FILLER_40_75 ();
 sg13g2_fill_2 FILLER_40_94 ();
 sg13g2_fill_2 FILLER_40_102 ();
 sg13g2_fill_2 FILLER_40_109 ();
 sg13g2_fill_1 FILLER_40_111 ();
 sg13g2_decap_8 FILLER_40_118 ();
 sg13g2_decap_8 FILLER_40_125 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_fill_2 FILLER_40_147 ();
 sg13g2_fill_1 FILLER_40_154 ();
 sg13g2_decap_4 FILLER_40_172 ();
 sg13g2_fill_1 FILLER_40_201 ();
 sg13g2_decap_8 FILLER_40_207 ();
 sg13g2_fill_2 FILLER_40_214 ();
 sg13g2_fill_1 FILLER_40_216 ();
 sg13g2_fill_1 FILLER_40_235 ();
 sg13g2_fill_1 FILLER_40_241 ();
 sg13g2_fill_2 FILLER_40_246 ();
 sg13g2_fill_1 FILLER_40_248 ();
 sg13g2_fill_2 FILLER_40_254 ();
 sg13g2_fill_1 FILLER_40_256 ();
 sg13g2_decap_4 FILLER_40_262 ();
 sg13g2_fill_2 FILLER_40_266 ();
 sg13g2_fill_1 FILLER_40_272 ();
 sg13g2_fill_2 FILLER_40_300 ();
 sg13g2_fill_1 FILLER_40_302 ();
 sg13g2_fill_2 FILLER_40_329 ();
 sg13g2_fill_2 FILLER_40_363 ();
 sg13g2_fill_1 FILLER_40_365 ();
 sg13g2_decap_4 FILLER_40_378 ();
 sg13g2_fill_1 FILLER_40_382 ();
 sg13g2_fill_2 FILLER_40_395 ();
 sg13g2_fill_1 FILLER_40_397 ();
 sg13g2_fill_2 FILLER_40_406 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_4 FILLER_41_35 ();
 sg13g2_fill_1 FILLER_41_58 ();
 sg13g2_fill_2 FILLER_41_64 ();
 sg13g2_fill_1 FILLER_41_79 ();
 sg13g2_decap_4 FILLER_41_85 ();
 sg13g2_fill_2 FILLER_41_89 ();
 sg13g2_fill_2 FILLER_41_102 ();
 sg13g2_fill_1 FILLER_41_104 ();
 sg13g2_fill_1 FILLER_41_111 ();
 sg13g2_decap_4 FILLER_41_138 ();
 sg13g2_decap_8 FILLER_41_156 ();
 sg13g2_decap_4 FILLER_41_167 ();
 sg13g2_fill_1 FILLER_41_171 ();
 sg13g2_decap_4 FILLER_41_182 ();
 sg13g2_fill_2 FILLER_41_219 ();
 sg13g2_fill_1 FILLER_41_221 ();
 sg13g2_fill_1 FILLER_41_230 ();
 sg13g2_fill_2 FILLER_41_241 ();
 sg13g2_fill_1 FILLER_41_243 ();
 sg13g2_decap_8 FILLER_41_300 ();
 sg13g2_decap_8 FILLER_41_307 ();
 sg13g2_decap_4 FILLER_41_314 ();
 sg13g2_fill_2 FILLER_41_326 ();
 sg13g2_fill_1 FILLER_41_328 ();
 sg13g2_fill_2 FILLER_41_337 ();
 sg13g2_fill_1 FILLER_41_339 ();
 sg13g2_decap_4 FILLER_41_348 ();
 sg13g2_fill_2 FILLER_41_357 ();
 sg13g2_fill_2 FILLER_41_388 ();
 sg13g2_fill_1 FILLER_41_390 ();
 sg13g2_fill_2 FILLER_41_399 ();
 sg13g2_fill_2 FILLER_41_406 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_4 FILLER_42_35 ();
 sg13g2_fill_2 FILLER_42_58 ();
 sg13g2_fill_1 FILLER_42_64 ();
 sg13g2_decap_4 FILLER_42_70 ();
 sg13g2_fill_2 FILLER_42_109 ();
 sg13g2_fill_1 FILLER_42_111 ();
 sg13g2_decap_4 FILLER_42_122 ();
 sg13g2_fill_2 FILLER_42_132 ();
 sg13g2_fill_1 FILLER_42_134 ();
 sg13g2_fill_1 FILLER_42_143 ();
 sg13g2_fill_2 FILLER_42_149 ();
 sg13g2_decap_8 FILLER_42_169 ();
 sg13g2_decap_4 FILLER_42_176 ();
 sg13g2_fill_2 FILLER_42_189 ();
 sg13g2_fill_1 FILLER_42_191 ();
 sg13g2_fill_2 FILLER_42_200 ();
 sg13g2_fill_1 FILLER_42_202 ();
 sg13g2_fill_1 FILLER_42_211 ();
 sg13g2_fill_2 FILLER_42_223 ();
 sg13g2_decap_8 FILLER_42_230 ();
 sg13g2_decap_8 FILLER_42_237 ();
 sg13g2_fill_1 FILLER_42_244 ();
 sg13g2_decap_8 FILLER_42_253 ();
 sg13g2_decap_8 FILLER_42_265 ();
 sg13g2_fill_2 FILLER_42_272 ();
 sg13g2_fill_1 FILLER_42_274 ();
 sg13g2_decap_8 FILLER_42_285 ();
 sg13g2_fill_1 FILLER_42_292 ();
 sg13g2_decap_4 FILLER_42_298 ();
 sg13g2_decap_4 FILLER_42_329 ();
 sg13g2_fill_2 FILLER_42_333 ();
 sg13g2_fill_2 FILLER_42_343 ();
 sg13g2_fill_1 FILLER_42_362 ();
 sg13g2_fill_2 FILLER_42_367 ();
 sg13g2_decap_4 FILLER_42_382 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_4 FILLER_43_28 ();
 sg13g2_fill_2 FILLER_43_32 ();
 sg13g2_decap_8 FILLER_43_43 ();
 sg13g2_fill_1 FILLER_43_50 ();
 sg13g2_decap_4 FILLER_43_77 ();
 sg13g2_fill_2 FILLER_43_109 ();
 sg13g2_fill_2 FILLER_43_117 ();
 sg13g2_fill_1 FILLER_43_128 ();
 sg13g2_fill_2 FILLER_43_134 ();
 sg13g2_fill_1 FILLER_43_136 ();
 sg13g2_fill_2 FILLER_43_147 ();
 sg13g2_fill_1 FILLER_43_149 ();
 sg13g2_fill_2 FILLER_43_172 ();
 sg13g2_fill_1 FILLER_43_174 ();
 sg13g2_fill_2 FILLER_43_192 ();
 sg13g2_fill_1 FILLER_43_194 ();
 sg13g2_decap_8 FILLER_43_201 ();
 sg13g2_fill_2 FILLER_43_212 ();
 sg13g2_fill_2 FILLER_43_222 ();
 sg13g2_fill_1 FILLER_43_229 ();
 sg13g2_fill_2 FILLER_43_244 ();
 sg13g2_fill_1 FILLER_43_246 ();
 sg13g2_fill_1 FILLER_43_263 ();
 sg13g2_fill_2 FILLER_43_282 ();
 sg13g2_fill_2 FILLER_43_291 ();
 sg13g2_fill_1 FILLER_43_293 ();
 sg13g2_fill_1 FILLER_43_303 ();
 sg13g2_fill_2 FILLER_43_327 ();
 sg13g2_fill_1 FILLER_43_329 ();
 sg13g2_fill_2 FILLER_43_338 ();
 sg13g2_fill_1 FILLER_43_362 ();
 sg13g2_fill_2 FILLER_43_368 ();
 sg13g2_fill_1 FILLER_43_370 ();
 sg13g2_fill_2 FILLER_43_376 ();
 sg13g2_fill_1 FILLER_43_383 ();
 sg13g2_decap_4 FILLER_43_405 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_4 FILLER_44_28 ();
 sg13g2_fill_1 FILLER_44_32 ();
 sg13g2_fill_2 FILLER_44_38 ();
 sg13g2_fill_1 FILLER_44_40 ();
 sg13g2_fill_2 FILLER_44_46 ();
 sg13g2_decap_8 FILLER_44_53 ();
 sg13g2_fill_2 FILLER_44_60 ();
 sg13g2_fill_2 FILLER_44_73 ();
 sg13g2_fill_1 FILLER_44_87 ();
 sg13g2_decap_4 FILLER_44_92 ();
 sg13g2_fill_1 FILLER_44_96 ();
 sg13g2_fill_2 FILLER_44_102 ();
 sg13g2_fill_1 FILLER_44_110 ();
 sg13g2_fill_2 FILLER_44_124 ();
 sg13g2_fill_1 FILLER_44_126 ();
 sg13g2_fill_2 FILLER_44_131 ();
 sg13g2_fill_1 FILLER_44_133 ();
 sg13g2_fill_2 FILLER_44_145 ();
 sg13g2_fill_1 FILLER_44_147 ();
 sg13g2_fill_1 FILLER_44_172 ();
 sg13g2_fill_1 FILLER_44_194 ();
 sg13g2_fill_2 FILLER_44_200 ();
 sg13g2_fill_1 FILLER_44_208 ();
 sg13g2_fill_2 FILLER_44_214 ();
 sg13g2_fill_2 FILLER_44_221 ();
 sg13g2_fill_1 FILLER_44_223 ();
 sg13g2_fill_1 FILLER_44_228 ();
 sg13g2_decap_4 FILLER_44_240 ();
 sg13g2_decap_4 FILLER_44_252 ();
 sg13g2_fill_2 FILLER_44_256 ();
 sg13g2_decap_4 FILLER_44_274 ();
 sg13g2_decap_8 FILLER_44_297 ();
 sg13g2_fill_2 FILLER_44_316 ();
 sg13g2_fill_1 FILLER_44_318 ();
 sg13g2_fill_1 FILLER_44_328 ();
 sg13g2_decap_4 FILLER_44_348 ();
 sg13g2_fill_1 FILLER_44_352 ();
 sg13g2_fill_1 FILLER_44_388 ();
 sg13g2_fill_2 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_fill_2 FILLER_45_28 ();
 sg13g2_decap_4 FILLER_45_55 ();
 sg13g2_decap_4 FILLER_45_67 ();
 sg13g2_decap_4 FILLER_45_96 ();
 sg13g2_fill_1 FILLER_45_100 ();
 sg13g2_fill_1 FILLER_45_119 ();
 sg13g2_fill_2 FILLER_45_131 ();
 sg13g2_fill_1 FILLER_45_154 ();
 sg13g2_fill_1 FILLER_45_159 ();
 sg13g2_decap_8 FILLER_45_164 ();
 sg13g2_fill_2 FILLER_45_171 ();
 sg13g2_fill_1 FILLER_45_173 ();
 sg13g2_fill_2 FILLER_45_189 ();
 sg13g2_fill_2 FILLER_45_203 ();
 sg13g2_fill_2 FILLER_45_213 ();
 sg13g2_fill_1 FILLER_45_215 ();
 sg13g2_fill_2 FILLER_45_224 ();
 sg13g2_fill_2 FILLER_45_232 ();
 sg13g2_fill_1 FILLER_45_234 ();
 sg13g2_fill_1 FILLER_45_244 ();
 sg13g2_fill_1 FILLER_45_253 ();
 sg13g2_decap_4 FILLER_45_264 ();
 sg13g2_fill_1 FILLER_45_268 ();
 sg13g2_fill_2 FILLER_45_281 ();
 sg13g2_fill_1 FILLER_45_300 ();
 sg13g2_fill_1 FILLER_45_325 ();
 sg13g2_decap_8 FILLER_45_332 ();
 sg13g2_fill_2 FILLER_45_339 ();
 sg13g2_fill_2 FILLER_45_347 ();
 sg13g2_decap_4 FILLER_45_354 ();
 sg13g2_fill_1 FILLER_45_358 ();
 sg13g2_decap_4 FILLER_45_365 ();
 sg13g2_fill_2 FILLER_45_369 ();
 sg13g2_fill_1 FILLER_45_376 ();
 sg13g2_fill_2 FILLER_45_397 ();
 sg13g2_fill_2 FILLER_45_407 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_fill_1 FILLER_46_39 ();
 sg13g2_decap_8 FILLER_46_45 ();
 sg13g2_decap_8 FILLER_46_52 ();
 sg13g2_fill_2 FILLER_46_59 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_fill_2 FILLER_46_97 ();
 sg13g2_fill_1 FILLER_46_99 ();
 sg13g2_decap_8 FILLER_46_117 ();
 sg13g2_fill_2 FILLER_46_124 ();
 sg13g2_fill_2 FILLER_46_135 ();
 sg13g2_decap_8 FILLER_46_146 ();
 sg13g2_fill_2 FILLER_46_153 ();
 sg13g2_fill_2 FILLER_46_165 ();
 sg13g2_fill_1 FILLER_46_183 ();
 sg13g2_fill_1 FILLER_46_195 ();
 sg13g2_decap_4 FILLER_46_201 ();
 sg13g2_fill_2 FILLER_46_205 ();
 sg13g2_fill_2 FILLER_46_285 ();
 sg13g2_decap_8 FILLER_46_292 ();
 sg13g2_decap_8 FILLER_46_299 ();
 sg13g2_decap_4 FILLER_46_306 ();
 sg13g2_decap_4 FILLER_46_315 ();
 sg13g2_fill_1 FILLER_46_319 ();
 sg13g2_fill_2 FILLER_46_324 ();
 sg13g2_fill_1 FILLER_46_326 ();
 sg13g2_fill_2 FILLER_46_359 ();
 sg13g2_fill_1 FILLER_46_369 ();
 sg13g2_fill_2 FILLER_46_394 ();
 sg13g2_fill_1 FILLER_46_396 ();
 sg13g2_decap_4 FILLER_46_405 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_4 FILLER_47_21 ();
 sg13g2_fill_2 FILLER_47_25 ();
 sg13g2_fill_1 FILLER_47_52 ();
 sg13g2_decap_8 FILLER_47_58 ();
 sg13g2_fill_2 FILLER_47_65 ();
 sg13g2_fill_1 FILLER_47_67 ();
 sg13g2_fill_1 FILLER_47_82 ();
 sg13g2_decap_4 FILLER_47_110 ();
 sg13g2_fill_1 FILLER_47_114 ();
 sg13g2_fill_2 FILLER_47_126 ();
 sg13g2_fill_1 FILLER_47_128 ();
 sg13g2_fill_2 FILLER_47_135 ();
 sg13g2_fill_1 FILLER_47_137 ();
 sg13g2_fill_1 FILLER_47_157 ();
 sg13g2_fill_2 FILLER_47_171 ();
 sg13g2_fill_1 FILLER_47_177 ();
 sg13g2_fill_1 FILLER_47_182 ();
 sg13g2_fill_2 FILLER_47_195 ();
 sg13g2_fill_1 FILLER_47_197 ();
 sg13g2_decap_4 FILLER_47_207 ();
 sg13g2_fill_1 FILLER_47_211 ();
 sg13g2_decap_4 FILLER_47_217 ();
 sg13g2_decap_4 FILLER_47_229 ();
 sg13g2_fill_1 FILLER_47_254 ();
 sg13g2_fill_1 FILLER_47_260 ();
 sg13g2_fill_2 FILLER_47_269 ();
 sg13g2_fill_1 FILLER_47_271 ();
 sg13g2_fill_1 FILLER_47_335 ();
 sg13g2_decap_8 FILLER_47_341 ();
 sg13g2_fill_2 FILLER_47_352 ();
 sg13g2_fill_1 FILLER_47_354 ();
 sg13g2_decap_4 FILLER_47_365 ();
 sg13g2_fill_1 FILLER_47_369 ();
 sg13g2_decap_4 FILLER_47_375 ();
 sg13g2_fill_1 FILLER_47_383 ();
 sg13g2_fill_2 FILLER_47_389 ();
 sg13g2_fill_1 FILLER_47_391 ();
 sg13g2_fill_2 FILLER_47_407 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_fill_1 FILLER_48_28 ();
 sg13g2_fill_2 FILLER_48_34 ();
 sg13g2_fill_1 FILLER_48_36 ();
 sg13g2_fill_2 FILLER_48_60 ();
 sg13g2_decap_8 FILLER_48_71 ();
 sg13g2_fill_2 FILLER_48_78 ();
 sg13g2_fill_2 FILLER_48_92 ();
 sg13g2_fill_1 FILLER_48_116 ();
 sg13g2_decap_4 FILLER_48_125 ();
 sg13g2_fill_1 FILLER_48_144 ();
 sg13g2_fill_2 FILLER_48_178 ();
 sg13g2_fill_1 FILLER_48_187 ();
 sg13g2_fill_2 FILLER_48_203 ();
 sg13g2_fill_1 FILLER_48_218 ();
 sg13g2_decap_8 FILLER_48_274 ();
 sg13g2_decap_8 FILLER_48_281 ();
 sg13g2_decap_8 FILLER_48_288 ();
 sg13g2_decap_8 FILLER_48_295 ();
 sg13g2_fill_2 FILLER_48_302 ();
 sg13g2_fill_2 FILLER_48_324 ();
 sg13g2_fill_1 FILLER_48_326 ();
 sg13g2_fill_1 FILLER_48_332 ();
 sg13g2_fill_2 FILLER_48_353 ();
 sg13g2_fill_1 FILLER_48_363 ();
 sg13g2_decap_4 FILLER_48_376 ();
 sg13g2_fill_1 FILLER_48_389 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_4 FILLER_49_28 ();
 sg13g2_decap_4 FILLER_49_36 ();
 sg13g2_fill_2 FILLER_49_44 ();
 sg13g2_fill_1 FILLER_49_46 ();
 sg13g2_fill_2 FILLER_49_52 ();
 sg13g2_fill_2 FILLER_49_66 ();
 sg13g2_decap_4 FILLER_49_84 ();
 sg13g2_fill_2 FILLER_49_88 ();
 sg13g2_decap_8 FILLER_49_96 ();
 sg13g2_decap_4 FILLER_49_113 ();
 sg13g2_fill_1 FILLER_49_129 ();
 sg13g2_fill_2 FILLER_49_139 ();
 sg13g2_decap_4 FILLER_49_147 ();
 sg13g2_decap_4 FILLER_49_155 ();
 sg13g2_fill_1 FILLER_49_159 ();
 sg13g2_decap_4 FILLER_49_166 ();
 sg13g2_decap_8 FILLER_49_173 ();
 sg13g2_fill_2 FILLER_49_192 ();
 sg13g2_fill_1 FILLER_49_199 ();
 sg13g2_fill_2 FILLER_49_204 ();
 sg13g2_fill_1 FILLER_49_206 ();
 sg13g2_fill_2 FILLER_49_211 ();
 sg13g2_decap_8 FILLER_49_217 ();
 sg13g2_fill_2 FILLER_49_224 ();
 sg13g2_fill_1 FILLER_49_226 ();
 sg13g2_decap_8 FILLER_49_233 ();
 sg13g2_decap_8 FILLER_49_240 ();
 sg13g2_fill_2 FILLER_49_247 ();
 sg13g2_fill_1 FILLER_49_249 ();
 sg13g2_decap_8 FILLER_49_254 ();
 sg13g2_fill_1 FILLER_49_261 ();
 sg13g2_fill_2 FILLER_49_267 ();
 sg13g2_decap_8 FILLER_49_297 ();
 sg13g2_fill_1 FILLER_49_304 ();
 sg13g2_decap_8 FILLER_49_345 ();
 sg13g2_fill_1 FILLER_49_360 ();
 sg13g2_fill_1 FILLER_49_378 ();
 sg13g2_fill_2 FILLER_49_387 ();
 sg13g2_fill_1 FILLER_49_389 ();
 sg13g2_decap_4 FILLER_49_405 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_fill_1 FILLER_50_21 ();
 sg13g2_fill_1 FILLER_50_37 ();
 sg13g2_fill_2 FILLER_50_44 ();
 sg13g2_decap_4 FILLER_50_57 ();
 sg13g2_fill_1 FILLER_50_61 ();
 sg13g2_decap_4 FILLER_50_73 ();
 sg13g2_fill_2 FILLER_50_89 ();
 sg13g2_fill_1 FILLER_50_91 ();
 sg13g2_fill_1 FILLER_50_115 ();
 sg13g2_decap_8 FILLER_50_122 ();
 sg13g2_decap_4 FILLER_50_129 ();
 sg13g2_fill_1 FILLER_50_133 ();
 sg13g2_fill_1 FILLER_50_138 ();
 sg13g2_fill_1 FILLER_50_145 ();
 sg13g2_fill_2 FILLER_50_158 ();
 sg13g2_decap_4 FILLER_50_165 ();
 sg13g2_fill_1 FILLER_50_169 ();
 sg13g2_fill_1 FILLER_50_184 ();
 sg13g2_fill_1 FILLER_50_214 ();
 sg13g2_fill_2 FILLER_50_226 ();
 sg13g2_decap_8 FILLER_50_233 ();
 sg13g2_fill_1 FILLER_50_240 ();
 sg13g2_decap_4 FILLER_50_280 ();
 sg13g2_decap_4 FILLER_50_292 ();
 sg13g2_fill_2 FILLER_50_324 ();
 sg13g2_fill_1 FILLER_50_326 ();
 sg13g2_fill_1 FILLER_50_355 ();
 sg13g2_fill_2 FILLER_50_373 ();
 sg13g2_decap_4 FILLER_50_380 ();
 sg13g2_fill_1 FILLER_50_384 ();
 sg13g2_fill_2 FILLER_50_398 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_4 FILLER_51_21 ();
 sg13g2_fill_1 FILLER_51_25 ();
 sg13g2_fill_2 FILLER_51_45 ();
 sg13g2_fill_2 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_88 ();
 sg13g2_decap_4 FILLER_51_95 ();
 sg13g2_fill_2 FILLER_51_111 ();
 sg13g2_fill_1 FILLER_51_113 ();
 sg13g2_fill_1 FILLER_51_124 ();
 sg13g2_fill_1 FILLER_51_135 ();
 sg13g2_fill_2 FILLER_51_154 ();
 sg13g2_decap_8 FILLER_51_162 ();
 sg13g2_fill_2 FILLER_51_220 ();
 sg13g2_decap_4 FILLER_51_227 ();
 sg13g2_fill_2 FILLER_51_243 ();
 sg13g2_fill_1 FILLER_51_245 ();
 sg13g2_fill_2 FILLER_51_250 ();
 sg13g2_fill_1 FILLER_51_252 ();
 sg13g2_decap_4 FILLER_51_266 ();
 sg13g2_fill_1 FILLER_51_270 ();
 sg13g2_decap_8 FILLER_51_281 ();
 sg13g2_fill_2 FILLER_51_298 ();
 sg13g2_decap_4 FILLER_51_324 ();
 sg13g2_fill_1 FILLER_51_340 ();
 sg13g2_fill_1 FILLER_51_345 ();
 sg13g2_decap_8 FILLER_51_354 ();
 sg13g2_fill_1 FILLER_51_375 ();
 sg13g2_fill_2 FILLER_51_390 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_fill_1 FILLER_52_28 ();
 sg13g2_fill_2 FILLER_52_36 ();
 sg13g2_fill_1 FILLER_52_38 ();
 sg13g2_fill_2 FILLER_52_43 ();
 sg13g2_decap_4 FILLER_52_65 ();
 sg13g2_fill_2 FILLER_52_74 ();
 sg13g2_fill_1 FILLER_52_76 ();
 sg13g2_fill_1 FILLER_52_92 ();
 sg13g2_fill_2 FILLER_52_103 ();
 sg13g2_decap_4 FILLER_52_121 ();
 sg13g2_fill_2 FILLER_52_130 ();
 sg13g2_fill_1 FILLER_52_132 ();
 sg13g2_decap_8 FILLER_52_138 ();
 sg13g2_decap_4 FILLER_52_145 ();
 sg13g2_fill_1 FILLER_52_149 ();
 sg13g2_fill_2 FILLER_52_158 ();
 sg13g2_fill_2 FILLER_52_178 ();
 sg13g2_fill_1 FILLER_52_180 ();
 sg13g2_fill_2 FILLER_52_190 ();
 sg13g2_fill_2 FILLER_52_214 ();
 sg13g2_fill_2 FILLER_52_234 ();
 sg13g2_fill_1 FILLER_52_236 ();
 sg13g2_fill_1 FILLER_52_249 ();
 sg13g2_decap_4 FILLER_52_256 ();
 sg13g2_fill_2 FILLER_52_260 ();
 sg13g2_fill_1 FILLER_52_270 ();
 sg13g2_fill_2 FILLER_52_279 ();
 sg13g2_fill_1 FILLER_52_281 ();
 sg13g2_fill_1 FILLER_52_290 ();
 sg13g2_fill_1 FILLER_52_296 ();
 sg13g2_decap_8 FILLER_52_319 ();
 sg13g2_fill_2 FILLER_52_326 ();
 sg13g2_fill_2 FILLER_52_336 ();
 sg13g2_fill_1 FILLER_52_338 ();
 sg13g2_fill_1 FILLER_52_354 ();
 sg13g2_fill_2 FILLER_52_368 ();
 sg13g2_fill_1 FILLER_52_370 ();
 sg13g2_decap_4 FILLER_52_380 ();
 sg13g2_fill_1 FILLER_52_384 ();
 sg13g2_fill_1 FILLER_52_401 ();
 sg13g2_fill_2 FILLER_52_407 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_fill_2 FILLER_53_28 ();
 sg13g2_fill_1 FILLER_53_34 ();
 sg13g2_fill_1 FILLER_53_45 ();
 sg13g2_fill_2 FILLER_53_51 ();
 sg13g2_fill_1 FILLER_53_53 ();
 sg13g2_fill_1 FILLER_53_64 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_fill_2 FILLER_53_91 ();
 sg13g2_fill_2 FILLER_53_104 ();
 sg13g2_decap_4 FILLER_53_122 ();
 sg13g2_fill_1 FILLER_53_156 ();
 sg13g2_fill_1 FILLER_53_162 ();
 sg13g2_fill_2 FILLER_53_171 ();
 sg13g2_fill_2 FILLER_53_187 ();
 sg13g2_fill_1 FILLER_53_189 ();
 sg13g2_decap_4 FILLER_53_205 ();
 sg13g2_fill_2 FILLER_53_209 ();
 sg13g2_decap_4 FILLER_53_218 ();
 sg13g2_fill_1 FILLER_53_222 ();
 sg13g2_fill_1 FILLER_53_237 ();
 sg13g2_fill_1 FILLER_53_247 ();
 sg13g2_fill_2 FILLER_53_284 ();
 sg13g2_fill_1 FILLER_53_286 ();
 sg13g2_fill_1 FILLER_53_292 ();
 sg13g2_decap_4 FILLER_53_298 ();
 sg13g2_fill_2 FILLER_53_326 ();
 sg13g2_fill_1 FILLER_53_328 ();
 sg13g2_fill_1 FILLER_53_333 ();
 sg13g2_decap_8 FILLER_53_339 ();
 sg13g2_fill_2 FILLER_53_346 ();
 sg13g2_fill_2 FILLER_53_400 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_4 FILLER_54_21 ();
 sg13g2_fill_2 FILLER_54_25 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_fill_2 FILLER_54_47 ();
 sg13g2_fill_2 FILLER_54_54 ();
 sg13g2_fill_1 FILLER_54_56 ();
 sg13g2_decap_4 FILLER_54_63 ();
 sg13g2_fill_1 FILLER_54_67 ();
 sg13g2_decap_4 FILLER_54_72 ();
 sg13g2_fill_2 FILLER_54_76 ();
 sg13g2_fill_2 FILLER_54_89 ();
 sg13g2_fill_1 FILLER_54_91 ();
 sg13g2_fill_2 FILLER_54_98 ();
 sg13g2_fill_1 FILLER_54_100 ();
 sg13g2_decap_4 FILLER_54_107 ();
 sg13g2_fill_1 FILLER_54_111 ();
 sg13g2_fill_2 FILLER_54_117 ();
 sg13g2_decap_4 FILLER_54_142 ();
 sg13g2_fill_2 FILLER_54_157 ();
 sg13g2_fill_2 FILLER_54_167 ();
 sg13g2_fill_2 FILLER_54_178 ();
 sg13g2_fill_2 FILLER_54_193 ();
 sg13g2_decap_8 FILLER_54_207 ();
 sg13g2_fill_2 FILLER_54_214 ();
 sg13g2_fill_1 FILLER_54_216 ();
 sg13g2_fill_2 FILLER_54_223 ();
 sg13g2_fill_1 FILLER_54_225 ();
 sg13g2_decap_8 FILLER_54_231 ();
 sg13g2_fill_1 FILLER_54_238 ();
 sg13g2_decap_4 FILLER_54_244 ();
 sg13g2_fill_1 FILLER_54_248 ();
 sg13g2_decap_4 FILLER_54_257 ();
 sg13g2_fill_1 FILLER_54_261 ();
 sg13g2_fill_1 FILLER_54_279 ();
 sg13g2_fill_2 FILLER_54_306 ();
 sg13g2_fill_2 FILLER_54_318 ();
 sg13g2_decap_4 FILLER_54_347 ();
 sg13g2_decap_8 FILLER_54_360 ();
 sg13g2_decap_8 FILLER_54_367 ();
 sg13g2_decap_8 FILLER_54_374 ();
 sg13g2_decap_8 FILLER_54_385 ();
 sg13g2_fill_2 FILLER_54_392 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_4 FILLER_55_28 ();
 sg13g2_fill_2 FILLER_55_32 ();
 sg13g2_fill_2 FILLER_55_39 ();
 sg13g2_fill_1 FILLER_55_41 ();
 sg13g2_fill_1 FILLER_55_46 ();
 sg13g2_decap_4 FILLER_55_51 ();
 sg13g2_fill_1 FILLER_55_55 ();
 sg13g2_fill_1 FILLER_55_62 ();
 sg13g2_fill_1 FILLER_55_72 ();
 sg13g2_fill_1 FILLER_55_78 ();
 sg13g2_fill_1 FILLER_55_83 ();
 sg13g2_decap_4 FILLER_55_131 ();
 sg13g2_fill_1 FILLER_55_135 ();
 sg13g2_fill_1 FILLER_55_141 ();
 sg13g2_fill_2 FILLER_55_150 ();
 sg13g2_fill_1 FILLER_55_152 ();
 sg13g2_decap_4 FILLER_55_175 ();
 sg13g2_decap_8 FILLER_55_195 ();
 sg13g2_decap_4 FILLER_55_207 ();
 sg13g2_fill_1 FILLER_55_211 ();
 sg13g2_fill_1 FILLER_55_243 ();
 sg13g2_decap_4 FILLER_55_252 ();
 sg13g2_decap_8 FILLER_55_265 ();
 sg13g2_fill_1 FILLER_55_272 ();
 sg13g2_fill_2 FILLER_55_277 ();
 sg13g2_fill_1 FILLER_55_279 ();
 sg13g2_decap_4 FILLER_55_299 ();
 sg13g2_fill_1 FILLER_55_303 ();
 sg13g2_decap_4 FILLER_55_309 ();
 sg13g2_decap_4 FILLER_55_319 ();
 sg13g2_fill_2 FILLER_55_328 ();
 sg13g2_fill_2 FILLER_55_334 ();
 sg13g2_fill_1 FILLER_55_343 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_fill_2 FILLER_56_21 ();
 sg13g2_fill_2 FILLER_56_37 ();
 sg13g2_fill_1 FILLER_56_39 ();
 sg13g2_decap_4 FILLER_56_56 ();
 sg13g2_fill_2 FILLER_56_60 ();
 sg13g2_decap_4 FILLER_56_70 ();
 sg13g2_fill_2 FILLER_56_85 ();
 sg13g2_fill_2 FILLER_56_92 ();
 sg13g2_fill_1 FILLER_56_94 ();
 sg13g2_decap_8 FILLER_56_101 ();
 sg13g2_decap_4 FILLER_56_112 ();
 sg13g2_decap_4 FILLER_56_120 ();
 sg13g2_fill_2 FILLER_56_143 ();
 sg13g2_fill_1 FILLER_56_145 ();
 sg13g2_fill_2 FILLER_56_160 ();
 sg13g2_fill_1 FILLER_56_162 ();
 sg13g2_decap_4 FILLER_56_168 ();
 sg13g2_fill_1 FILLER_56_182 ();
 sg13g2_fill_2 FILLER_56_199 ();
 sg13g2_fill_2 FILLER_56_211 ();
 sg13g2_fill_1 FILLER_56_213 ();
 sg13g2_fill_2 FILLER_56_224 ();
 sg13g2_fill_1 FILLER_56_226 ();
 sg13g2_decap_8 FILLER_56_245 ();
 sg13g2_decap_4 FILLER_56_262 ();
 sg13g2_fill_1 FILLER_56_266 ();
 sg13g2_fill_2 FILLER_56_283 ();
 sg13g2_fill_1 FILLER_56_285 ();
 sg13g2_decap_4 FILLER_56_295 ();
 sg13g2_fill_1 FILLER_56_303 ();
 sg13g2_fill_2 FILLER_56_318 ();
 sg13g2_fill_1 FILLER_56_320 ();
 sg13g2_fill_1 FILLER_56_335 ();
 sg13g2_decap_4 FILLER_56_341 ();
 sg13g2_fill_2 FILLER_56_345 ();
 sg13g2_fill_2 FILLER_56_352 ();
 sg13g2_fill_1 FILLER_56_354 ();
 sg13g2_fill_2 FILLER_56_368 ();
 sg13g2_fill_1 FILLER_56_370 ();
 sg13g2_decap_4 FILLER_56_391 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_4 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_36 ();
 sg13g2_fill_2 FILLER_57_47 ();
 sg13g2_fill_1 FILLER_57_58 ();
 sg13g2_fill_1 FILLER_57_68 ();
 sg13g2_fill_2 FILLER_57_102 ();
 sg13g2_fill_1 FILLER_57_104 ();
 sg13g2_fill_1 FILLER_57_155 ();
 sg13g2_decap_8 FILLER_57_161 ();
 sg13g2_decap_8 FILLER_57_168 ();
 sg13g2_fill_2 FILLER_57_188 ();
 sg13g2_decap_4 FILLER_57_195 ();
 sg13g2_fill_1 FILLER_57_199 ();
 sg13g2_fill_1 FILLER_57_205 ();
 sg13g2_fill_2 FILLER_57_221 ();
 sg13g2_fill_1 FILLER_57_223 ();
 sg13g2_fill_2 FILLER_57_229 ();
 sg13g2_fill_2 FILLER_57_244 ();
 sg13g2_decap_4 FILLER_57_251 ();
 sg13g2_decap_4 FILLER_57_273 ();
 sg13g2_fill_2 FILLER_57_277 ();
 sg13g2_fill_2 FILLER_57_285 ();
 sg13g2_fill_1 FILLER_57_287 ();
 sg13g2_fill_1 FILLER_57_339 ();
 sg13g2_fill_2 FILLER_57_352 ();
 sg13g2_decap_4 FILLER_57_364 ();
 sg13g2_fill_2 FILLER_57_368 ();
 sg13g2_decap_8 FILLER_57_375 ();
 sg13g2_fill_1 FILLER_57_382 ();
 sg13g2_fill_1 FILLER_57_401 ();
 sg13g2_fill_2 FILLER_57_406 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_4 FILLER_58_21 ();
 sg13g2_fill_1 FILLER_58_25 ();
 sg13g2_decap_4 FILLER_58_65 ();
 sg13g2_fill_1 FILLER_58_69 ();
 sg13g2_decap_4 FILLER_58_75 ();
 sg13g2_fill_2 FILLER_58_79 ();
 sg13g2_fill_2 FILLER_58_86 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_fill_1 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_109 ();
 sg13g2_decap_8 FILLER_58_121 ();
 sg13g2_fill_1 FILLER_58_128 ();
 sg13g2_decap_4 FILLER_58_138 ();
 sg13g2_fill_2 FILLER_58_142 ();
 sg13g2_fill_1 FILLER_58_148 ();
 sg13g2_decap_8 FILLER_58_181 ();
 sg13g2_decap_4 FILLER_58_194 ();
 sg13g2_fill_1 FILLER_58_198 ();
 sg13g2_decap_8 FILLER_58_208 ();
 sg13g2_fill_2 FILLER_58_221 ();
 sg13g2_fill_1 FILLER_58_228 ();
 sg13g2_decap_4 FILLER_58_237 ();
 sg13g2_decap_8 FILLER_58_257 ();
 sg13g2_fill_2 FILLER_58_264 ();
 sg13g2_decap_8 FILLER_58_296 ();
 sg13g2_decap_4 FILLER_58_303 ();
 sg13g2_fill_1 FILLER_58_307 ();
 sg13g2_fill_1 FILLER_58_326 ();
 sg13g2_decap_8 FILLER_58_332 ();
 sg13g2_fill_2 FILLER_58_339 ();
 sg13g2_decap_4 FILLER_58_346 ();
 sg13g2_decap_4 FILLER_58_382 ();
 sg13g2_fill_2 FILLER_58_406 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_fill_2 FILLER_59_28 ();
 sg13g2_fill_1 FILLER_59_30 ();
 sg13g2_fill_1 FILLER_59_46 ();
 sg13g2_fill_1 FILLER_59_56 ();
 sg13g2_fill_2 FILLER_59_61 ();
 sg13g2_fill_1 FILLER_59_67 ();
 sg13g2_fill_2 FILLER_59_77 ();
 sg13g2_fill_2 FILLER_59_105 ();
 sg13g2_fill_1 FILLER_59_107 ();
 sg13g2_fill_2 FILLER_59_114 ();
 sg13g2_fill_1 FILLER_59_116 ();
 sg13g2_fill_2 FILLER_59_138 ();
 sg13g2_fill_1 FILLER_59_140 ();
 sg13g2_fill_2 FILLER_59_146 ();
 sg13g2_fill_1 FILLER_59_148 ();
 sg13g2_decap_8 FILLER_59_155 ();
 sg13g2_fill_1 FILLER_59_162 ();
 sg13g2_fill_2 FILLER_59_171 ();
 sg13g2_fill_2 FILLER_59_184 ();
 sg13g2_fill_1 FILLER_59_192 ();
 sg13g2_fill_1 FILLER_59_202 ();
 sg13g2_fill_2 FILLER_59_219 ();
 sg13g2_decap_4 FILLER_59_229 ();
 sg13g2_decap_4 FILLER_59_237 ();
 sg13g2_fill_1 FILLER_59_241 ();
 sg13g2_fill_1 FILLER_59_246 ();
 sg13g2_decap_4 FILLER_59_251 ();
 sg13g2_fill_2 FILLER_59_276 ();
 sg13g2_fill_1 FILLER_59_278 ();
 sg13g2_decap_4 FILLER_59_313 ();
 sg13g2_fill_2 FILLER_59_324 ();
 sg13g2_fill_1 FILLER_59_342 ();
 sg13g2_decap_4 FILLER_59_357 ();
 sg13g2_fill_1 FILLER_59_361 ();
 sg13g2_fill_2 FILLER_59_375 ();
 sg13g2_decap_4 FILLER_59_393 ();
 sg13g2_fill_1 FILLER_59_397 ();
 sg13g2_fill_2 FILLER_59_406 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_4 FILLER_60_28 ();
 sg13g2_fill_2 FILLER_60_32 ();
 sg13g2_fill_2 FILLER_60_50 ();
 sg13g2_fill_1 FILLER_60_52 ();
 sg13g2_fill_1 FILLER_60_69 ();
 sg13g2_fill_2 FILLER_60_80 ();
 sg13g2_fill_1 FILLER_60_82 ();
 sg13g2_fill_2 FILLER_60_108 ();
 sg13g2_fill_2 FILLER_60_114 ();
 sg13g2_fill_1 FILLER_60_116 ();
 sg13g2_fill_1 FILLER_60_123 ();
 sg13g2_fill_2 FILLER_60_142 ();
 sg13g2_fill_2 FILLER_60_162 ();
 sg13g2_decap_4 FILLER_60_183 ();
 sg13g2_decap_8 FILLER_60_192 ();
 sg13g2_decap_4 FILLER_60_199 ();
 sg13g2_fill_1 FILLER_60_237 ();
 sg13g2_fill_2 FILLER_60_263 ();
 sg13g2_decap_8 FILLER_60_269 ();
 sg13g2_decap_4 FILLER_60_285 ();
 sg13g2_fill_2 FILLER_60_289 ();
 sg13g2_fill_1 FILLER_60_299 ();
 sg13g2_decap_8 FILLER_60_308 ();
 sg13g2_fill_1 FILLER_60_315 ();
 sg13g2_fill_2 FILLER_60_336 ();
 sg13g2_fill_1 FILLER_60_338 ();
 sg13g2_fill_1 FILLER_60_347 ();
 sg13g2_decap_4 FILLER_60_372 ();
 sg13g2_fill_2 FILLER_60_386 ();
 sg13g2_fill_1 FILLER_60_388 ();
 sg13g2_fill_2 FILLER_60_398 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_4 FILLER_61_28 ();
 sg13g2_fill_1 FILLER_61_38 ();
 sg13g2_decap_4 FILLER_61_43 ();
 sg13g2_decap_8 FILLER_61_52 ();
 sg13g2_decap_4 FILLER_61_59 ();
 sg13g2_fill_2 FILLER_61_63 ();
 sg13g2_fill_1 FILLER_61_78 ();
 sg13g2_fill_1 FILLER_61_84 ();
 sg13g2_fill_2 FILLER_61_93 ();
 sg13g2_fill_1 FILLER_61_95 ();
 sg13g2_fill_1 FILLER_61_105 ();
 sg13g2_decap_4 FILLER_61_111 ();
 sg13g2_fill_2 FILLER_61_115 ();
 sg13g2_fill_2 FILLER_61_125 ();
 sg13g2_fill_1 FILLER_61_127 ();
 sg13g2_decap_4 FILLER_61_134 ();
 sg13g2_fill_2 FILLER_61_148 ();
 sg13g2_fill_1 FILLER_61_164 ();
 sg13g2_fill_1 FILLER_61_186 ();
 sg13g2_fill_2 FILLER_61_196 ();
 sg13g2_fill_1 FILLER_61_198 ();
 sg13g2_decap_4 FILLER_61_211 ();
 sg13g2_fill_2 FILLER_61_227 ();
 sg13g2_fill_1 FILLER_61_229 ();
 sg13g2_decap_8 FILLER_61_236 ();
 sg13g2_fill_1 FILLER_61_247 ();
 sg13g2_decap_4 FILLER_61_252 ();
 sg13g2_fill_1 FILLER_61_269 ();
 sg13g2_fill_1 FILLER_61_302 ();
 sg13g2_decap_8 FILLER_61_314 ();
 sg13g2_fill_2 FILLER_61_338 ();
 sg13g2_decap_4 FILLER_61_344 ();
 sg13g2_fill_2 FILLER_61_348 ();
 sg13g2_decap_8 FILLER_61_359 ();
 sg13g2_fill_2 FILLER_61_379 ();
 sg13g2_fill_1 FILLER_61_389 ();
 sg13g2_fill_2 FILLER_61_406 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_fill_2 FILLER_62_41 ();
 sg13g2_fill_1 FILLER_62_75 ();
 sg13g2_fill_1 FILLER_62_100 ();
 sg13g2_fill_2 FILLER_62_119 ();
 sg13g2_fill_1 FILLER_62_130 ();
 sg13g2_fill_2 FILLER_62_141 ();
 sg13g2_fill_1 FILLER_62_143 ();
 sg13g2_fill_1 FILLER_62_163 ();
 sg13g2_fill_1 FILLER_62_175 ();
 sg13g2_fill_2 FILLER_62_184 ();
 sg13g2_fill_2 FILLER_62_195 ();
 sg13g2_fill_1 FILLER_62_197 ();
 sg13g2_fill_1 FILLER_62_206 ();
 sg13g2_decap_4 FILLER_62_217 ();
 sg13g2_decap_4 FILLER_62_225 ();
 sg13g2_fill_2 FILLER_62_269 ();
 sg13g2_decap_4 FILLER_62_287 ();
 sg13g2_fill_2 FILLER_62_302 ();
 sg13g2_fill_1 FILLER_62_326 ();
 sg13g2_decap_4 FILLER_62_334 ();
 sg13g2_fill_2 FILLER_62_338 ();
 sg13g2_decap_8 FILLER_62_353 ();
 sg13g2_decap_8 FILLER_62_367 ();
 sg13g2_fill_1 FILLER_62_388 ();
 sg13g2_fill_2 FILLER_62_406 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_4 FILLER_63_28 ();
 sg13g2_decap_4 FILLER_63_46 ();
 sg13g2_fill_2 FILLER_63_54 ();
 sg13g2_decap_4 FILLER_63_62 ();
 sg13g2_fill_1 FILLER_63_66 ();
 sg13g2_decap_4 FILLER_63_81 ();
 sg13g2_decap_8 FILLER_63_89 ();
 sg13g2_fill_1 FILLER_63_100 ();
 sg13g2_decap_4 FILLER_63_132 ();
 sg13g2_fill_1 FILLER_63_152 ();
 sg13g2_fill_2 FILLER_63_161 ();
 sg13g2_fill_1 FILLER_63_163 ();
 sg13g2_fill_1 FILLER_63_171 ();
 sg13g2_decap_4 FILLER_63_196 ();
 sg13g2_fill_2 FILLER_63_236 ();
 sg13g2_fill_1 FILLER_63_238 ();
 sg13g2_fill_2 FILLER_63_296 ();
 sg13g2_fill_1 FILLER_63_298 ();
 sg13g2_decap_4 FILLER_63_305 ();
 sg13g2_fill_1 FILLER_63_309 ();
 sg13g2_fill_2 FILLER_63_326 ();
 sg13g2_fill_1 FILLER_63_328 ();
 sg13g2_fill_2 FILLER_63_342 ();
 sg13g2_fill_1 FILLER_63_344 ();
 sg13g2_fill_1 FILLER_63_374 ();
 sg13g2_fill_1 FILLER_63_399 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_fill_1 FILLER_64_42 ();
 sg13g2_fill_2 FILLER_64_57 ();
 sg13g2_fill_1 FILLER_64_92 ();
 sg13g2_fill_2 FILLER_64_99 ();
 sg13g2_fill_1 FILLER_64_101 ();
 sg13g2_decap_8 FILLER_64_106 ();
 sg13g2_fill_2 FILLER_64_113 ();
 sg13g2_decap_4 FILLER_64_121 ();
 sg13g2_fill_2 FILLER_64_141 ();
 sg13g2_fill_1 FILLER_64_143 ();
 sg13g2_decap_8 FILLER_64_149 ();
 sg13g2_decap_4 FILLER_64_156 ();
 sg13g2_fill_1 FILLER_64_160 ();
 sg13g2_fill_1 FILLER_64_166 ();
 sg13g2_decap_8 FILLER_64_176 ();
 sg13g2_fill_1 FILLER_64_183 ();
 sg13g2_fill_2 FILLER_64_192 ();
 sg13g2_decap_4 FILLER_64_205 ();
 sg13g2_decap_8 FILLER_64_214 ();
 sg13g2_decap_8 FILLER_64_221 ();
 sg13g2_fill_1 FILLER_64_253 ();
 sg13g2_decap_8 FILLER_64_272 ();
 sg13g2_fill_2 FILLER_64_279 ();
 sg13g2_fill_1 FILLER_64_300 ();
 sg13g2_fill_2 FILLER_64_318 ();
 sg13g2_fill_1 FILLER_64_320 ();
 sg13g2_fill_2 FILLER_64_329 ();
 sg13g2_fill_1 FILLER_64_331 ();
 sg13g2_fill_2 FILLER_64_345 ();
 sg13g2_fill_2 FILLER_64_355 ();
 sg13g2_fill_1 FILLER_64_357 ();
 sg13g2_decap_4 FILLER_64_368 ();
 sg13g2_fill_1 FILLER_64_372 ();
 sg13g2_decap_8 FILLER_64_384 ();
 sg13g2_fill_1 FILLER_64_391 ();
 sg13g2_fill_1 FILLER_64_401 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_fill_1 FILLER_65_35 ();
 sg13g2_fill_2 FILLER_65_52 ();
 sg13g2_decap_4 FILLER_65_58 ();
 sg13g2_fill_2 FILLER_65_62 ();
 sg13g2_fill_1 FILLER_65_80 ();
 sg13g2_fill_1 FILLER_65_92 ();
 sg13g2_fill_1 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_118 ();
 sg13g2_fill_1 FILLER_65_125 ();
 sg13g2_decap_4 FILLER_65_136 ();
 sg13g2_fill_1 FILLER_65_140 ();
 sg13g2_fill_2 FILLER_65_164 ();
 sg13g2_fill_1 FILLER_65_166 ();
 sg13g2_fill_2 FILLER_65_173 ();
 sg13g2_decap_4 FILLER_65_185 ();
 sg13g2_decap_4 FILLER_65_206 ();
 sg13g2_fill_1 FILLER_65_242 ();
 sg13g2_fill_2 FILLER_65_305 ();
 sg13g2_fill_1 FILLER_65_307 ();
 sg13g2_fill_2 FILLER_65_320 ();
 sg13g2_fill_2 FILLER_65_330 ();
 sg13g2_fill_1 FILLER_65_332 ();
 sg13g2_decap_4 FILLER_65_341 ();
 sg13g2_fill_1 FILLER_65_345 ();
 sg13g2_fill_1 FILLER_65_384 ();
 sg13g2_fill_2 FILLER_65_406 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_fill_2 FILLER_66_42 ();
 sg13g2_fill_1 FILLER_66_55 ();
 sg13g2_fill_2 FILLER_66_68 ();
 sg13g2_decap_4 FILLER_66_96 ();
 sg13g2_fill_2 FILLER_66_100 ();
 sg13g2_decap_4 FILLER_66_108 ();
 sg13g2_fill_2 FILLER_66_112 ();
 sg13g2_fill_1 FILLER_66_134 ();
 sg13g2_fill_2 FILLER_66_150 ();
 sg13g2_fill_1 FILLER_66_152 ();
 sg13g2_fill_1 FILLER_66_180 ();
 sg13g2_decap_8 FILLER_66_221 ();
 sg13g2_fill_1 FILLER_66_228 ();
 sg13g2_fill_2 FILLER_66_238 ();
 sg13g2_fill_1 FILLER_66_240 ();
 sg13g2_fill_2 FILLER_66_245 ();
 sg13g2_fill_1 FILLER_66_247 ();
 sg13g2_fill_2 FILLER_66_258 ();
 sg13g2_fill_1 FILLER_66_266 ();
 sg13g2_decap_8 FILLER_66_271 ();
 sg13g2_decap_4 FILLER_66_278 ();
 sg13g2_fill_1 FILLER_66_282 ();
 sg13g2_decap_4 FILLER_66_289 ();
 sg13g2_fill_2 FILLER_66_307 ();
 sg13g2_fill_2 FILLER_66_318 ();
 sg13g2_fill_1 FILLER_66_320 ();
 sg13g2_fill_1 FILLER_66_364 ();
 sg13g2_decap_4 FILLER_66_369 ();
 sg13g2_fill_2 FILLER_66_373 ();
 sg13g2_decap_4 FILLER_66_394 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_fill_2 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_55 ();
 sg13g2_decap_8 FILLER_67_78 ();
 sg13g2_fill_2 FILLER_67_85 ();
 sg13g2_fill_1 FILLER_67_98 ();
 sg13g2_decap_4 FILLER_67_104 ();
 sg13g2_fill_2 FILLER_67_108 ();
 sg13g2_fill_1 FILLER_67_116 ();
 sg13g2_fill_2 FILLER_67_130 ();
 sg13g2_fill_1 FILLER_67_132 ();
 sg13g2_decap_8 FILLER_67_146 ();
 sg13g2_decap_4 FILLER_67_153 ();
 sg13g2_fill_1 FILLER_67_157 ();
 sg13g2_fill_1 FILLER_67_168 ();
 sg13g2_fill_2 FILLER_67_177 ();
 sg13g2_fill_2 FILLER_67_183 ();
 sg13g2_fill_1 FILLER_67_190 ();
 sg13g2_decap_4 FILLER_67_196 ();
 sg13g2_decap_8 FILLER_67_242 ();
 sg13g2_fill_2 FILLER_67_249 ();
 sg13g2_fill_1 FILLER_67_251 ();
 sg13g2_decap_8 FILLER_67_257 ();
 sg13g2_fill_2 FILLER_67_274 ();
 sg13g2_fill_2 FILLER_67_304 ();
 sg13g2_fill_1 FILLER_67_306 ();
 sg13g2_decap_4 FILLER_67_313 ();
 sg13g2_fill_2 FILLER_67_317 ();
 sg13g2_decap_8 FILLER_67_328 ();
 sg13g2_decap_4 FILLER_67_350 ();
 sg13g2_fill_2 FILLER_67_367 ();
 sg13g2_decap_4 FILLER_67_377 ();
 sg13g2_fill_1 FILLER_67_391 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_4 FILLER_68_42 ();
 sg13g2_fill_1 FILLER_68_60 ();
 sg13g2_fill_2 FILLER_68_66 ();
 sg13g2_fill_1 FILLER_68_72 ();
 sg13g2_fill_2 FILLER_68_79 ();
 sg13g2_fill_1 FILLER_68_97 ();
 sg13g2_fill_2 FILLER_68_114 ();
 sg13g2_fill_1 FILLER_68_116 ();
 sg13g2_decap_4 FILLER_68_123 ();
 sg13g2_fill_2 FILLER_68_132 ();
 sg13g2_fill_2 FILLER_68_139 ();
 sg13g2_decap_8 FILLER_68_161 ();
 sg13g2_fill_2 FILLER_68_168 ();
 sg13g2_fill_1 FILLER_68_174 ();
 sg13g2_fill_2 FILLER_68_178 ();
 sg13g2_fill_1 FILLER_68_180 ();
 sg13g2_fill_1 FILLER_68_208 ();
 sg13g2_fill_2 FILLER_68_217 ();
 sg13g2_fill_1 FILLER_68_219 ();
 sg13g2_fill_2 FILLER_68_257 ();
 sg13g2_fill_1 FILLER_68_259 ();
 sg13g2_decap_8 FILLER_68_275 ();
 sg13g2_decap_8 FILLER_68_282 ();
 sg13g2_decap_4 FILLER_68_289 ();
 sg13g2_fill_1 FILLER_68_293 ();
 sg13g2_fill_2 FILLER_68_325 ();
 sg13g2_fill_1 FILLER_68_335 ();
 sg13g2_decap_8 FILLER_68_341 ();
 sg13g2_decap_8 FILLER_68_348 ();
 sg13g2_decap_4 FILLER_68_355 ();
 sg13g2_fill_2 FILLER_68_364 ();
 sg13g2_fill_2 FILLER_68_371 ();
 sg13g2_fill_1 FILLER_68_373 ();
 sg13g2_decap_4 FILLER_68_379 ();
 sg13g2_fill_2 FILLER_68_398 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_4 FILLER_69_42 ();
 sg13g2_fill_1 FILLER_69_46 ();
 sg13g2_fill_1 FILLER_69_82 ();
 sg13g2_decap_4 FILLER_69_99 ();
 sg13g2_fill_1 FILLER_69_108 ();
 sg13g2_fill_2 FILLER_69_132 ();
 sg13g2_decap_8 FILLER_69_148 ();
 sg13g2_decap_4 FILLER_69_155 ();
 sg13g2_decap_4 FILLER_69_185 ();
 sg13g2_fill_1 FILLER_69_189 ();
 sg13g2_fill_2 FILLER_69_198 ();
 sg13g2_fill_1 FILLER_69_224 ();
 sg13g2_fill_1 FILLER_69_263 ();
 sg13g2_fill_2 FILLER_69_305 ();
 sg13g2_decap_4 FILLER_69_316 ();
 sg13g2_fill_1 FILLER_69_320 ();
 sg13g2_fill_1 FILLER_69_364 ();
 sg13g2_decap_8 FILLER_69_384 ();
 sg13g2_fill_2 FILLER_69_391 ();
 sg13g2_fill_1 FILLER_69_393 ();
 sg13g2_fill_2 FILLER_69_406 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_4 FILLER_70_56 ();
 sg13g2_fill_1 FILLER_70_60 ();
 sg13g2_fill_1 FILLER_70_67 ();
 sg13g2_fill_2 FILLER_70_77 ();
 sg13g2_fill_1 FILLER_70_79 ();
 sg13g2_fill_2 FILLER_70_104 ();
 sg13g2_fill_2 FILLER_70_124 ();
 sg13g2_fill_1 FILLER_70_126 ();
 sg13g2_fill_2 FILLER_70_142 ();
 sg13g2_fill_1 FILLER_70_144 ();
 sg13g2_decap_4 FILLER_70_175 ();
 sg13g2_decap_8 FILLER_70_224 ();
 sg13g2_decap_4 FILLER_70_231 ();
 sg13g2_fill_1 FILLER_70_235 ();
 sg13g2_fill_2 FILLER_70_252 ();
 sg13g2_fill_1 FILLER_70_273 ();
 sg13g2_decap_4 FILLER_70_280 ();
 sg13g2_fill_2 FILLER_70_292 ();
 sg13g2_fill_2 FILLER_70_308 ();
 sg13g2_fill_1 FILLER_70_321 ();
 sg13g2_fill_2 FILLER_70_335 ();
 sg13g2_fill_2 FILLER_70_349 ();
 sg13g2_fill_1 FILLER_70_363 ();
 sg13g2_decap_4 FILLER_70_369 ();
 sg13g2_fill_2 FILLER_70_373 ();
 sg13g2_decap_4 FILLER_70_395 ();
 sg13g2_fill_2 FILLER_70_399 ();
 sg13g2_decap_4 FILLER_70_405 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_fill_1 FILLER_71_62 ();
 sg13g2_fill_2 FILLER_71_69 ();
 sg13g2_fill_2 FILLER_71_77 ();
 sg13g2_fill_1 FILLER_71_79 ();
 sg13g2_decap_8 FILLER_71_96 ();
 sg13g2_decap_8 FILLER_71_103 ();
 sg13g2_decap_8 FILLER_71_110 ();
 sg13g2_decap_4 FILLER_71_117 ();
 sg13g2_fill_1 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_142 ();
 sg13g2_fill_1 FILLER_71_163 ();
 sg13g2_fill_2 FILLER_71_189 ();
 sg13g2_fill_1 FILLER_71_191 ();
 sg13g2_fill_2 FILLER_71_205 ();
 sg13g2_fill_1 FILLER_71_207 ();
 sg13g2_fill_2 FILLER_71_242 ();
 sg13g2_fill_1 FILLER_71_244 ();
 sg13g2_decap_4 FILLER_71_268 ();
 sg13g2_fill_1 FILLER_71_282 ();
 sg13g2_fill_2 FILLER_71_287 ();
 sg13g2_fill_1 FILLER_71_289 ();
 sg13g2_fill_1 FILLER_71_295 ();
 sg13g2_fill_2 FILLER_71_300 ();
 sg13g2_fill_1 FILLER_71_302 ();
 sg13g2_decap_4 FILLER_71_307 ();
 sg13g2_fill_1 FILLER_71_311 ();
 sg13g2_fill_2 FILLER_71_317 ();
 sg13g2_decap_4 FILLER_71_329 ();
 sg13g2_fill_1 FILLER_71_333 ();
 sg13g2_decap_8 FILLER_71_338 ();
 sg13g2_fill_2 FILLER_71_345 ();
 sg13g2_fill_1 FILLER_71_359 ();
 sg13g2_decap_8 FILLER_71_373 ();
 sg13g2_fill_1 FILLER_71_380 ();
 sg13g2_decap_8 FILLER_71_386 ();
 sg13g2_decap_8 FILLER_71_393 ();
 sg13g2_decap_8 FILLER_71_400 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_4 FILLER_72_49 ();
 sg13g2_fill_1 FILLER_72_53 ();
 sg13g2_decap_4 FILLER_72_62 ();
 sg13g2_fill_1 FILLER_72_66 ();
 sg13g2_fill_2 FILLER_72_73 ();
 sg13g2_fill_1 FILLER_72_75 ();
 sg13g2_fill_1 FILLER_72_108 ();
 sg13g2_fill_1 FILLER_72_121 ();
 sg13g2_decap_4 FILLER_72_139 ();
 sg13g2_fill_1 FILLER_72_157 ();
 sg13g2_fill_2 FILLER_72_194 ();
 sg13g2_decap_8 FILLER_72_222 ();
 sg13g2_fill_1 FILLER_72_229 ();
 sg13g2_fill_2 FILLER_72_238 ();
 sg13g2_fill_1 FILLER_72_240 ();
 sg13g2_fill_2 FILLER_72_263 ();
 sg13g2_fill_1 FILLER_72_265 ();
 sg13g2_fill_2 FILLER_72_282 ();
 sg13g2_fill_1 FILLER_72_293 ();
 sg13g2_fill_1 FILLER_72_306 ();
 sg13g2_decap_4 FILLER_72_317 ();
 sg13g2_fill_2 FILLER_72_321 ();
 sg13g2_fill_2 FILLER_72_328 ();
 sg13g2_decap_4 FILLER_72_362 ();
 sg13g2_fill_1 FILLER_72_366 ();
 sg13g2_fill_1 FILLER_72_380 ();
 sg13g2_decap_8 FILLER_72_394 ();
 sg13g2_decap_8 FILLER_72_401 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_4 FILLER_73_56 ();
 sg13g2_fill_1 FILLER_73_60 ();
 sg13g2_decap_8 FILLER_73_67 ();
 sg13g2_decap_8 FILLER_73_74 ();
 sg13g2_decap_4 FILLER_73_81 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_4 FILLER_73_98 ();
 sg13g2_fill_2 FILLER_73_102 ();
 sg13g2_decap_8 FILLER_73_115 ();
 sg13g2_fill_2 FILLER_73_122 ();
 sg13g2_fill_1 FILLER_73_124 ();
 sg13g2_fill_2 FILLER_73_134 ();
 sg13g2_fill_1 FILLER_73_136 ();
 sg13g2_decap_8 FILLER_73_167 ();
 sg13g2_fill_2 FILLER_73_203 ();
 sg13g2_decap_4 FILLER_73_209 ();
 sg13g2_fill_1 FILLER_73_213 ();
 sg13g2_fill_2 FILLER_73_248 ();
 sg13g2_fill_1 FILLER_73_255 ();
 sg13g2_decap_4 FILLER_73_274 ();
 sg13g2_fill_2 FILLER_73_278 ();
 sg13g2_fill_2 FILLER_73_293 ();
 sg13g2_fill_1 FILLER_73_295 ();
 sg13g2_fill_1 FILLER_73_304 ();
 sg13g2_decap_4 FILLER_73_379 ();
 sg13g2_decap_8 FILLER_73_396 ();
 sg13g2_decap_4 FILLER_73_403 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_4 FILLER_74_63 ();
 sg13g2_fill_1 FILLER_74_67 ();
 sg13g2_fill_2 FILLER_74_82 ();
 sg13g2_fill_1 FILLER_74_91 ();
 sg13g2_decap_4 FILLER_74_98 ();
 sg13g2_fill_1 FILLER_74_114 ();
 sg13g2_fill_1 FILLER_74_127 ();
 sg13g2_decap_4 FILLER_74_139 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_fill_2 FILLER_74_161 ();
 sg13g2_fill_1 FILLER_74_176 ();
 sg13g2_decap_4 FILLER_74_182 ();
 sg13g2_fill_2 FILLER_74_186 ();
 sg13g2_decap_8 FILLER_74_193 ();
 sg13g2_decap_8 FILLER_74_200 ();
 sg13g2_decap_8 FILLER_74_211 ();
 sg13g2_decap_8 FILLER_74_218 ();
 sg13g2_decap_8 FILLER_74_229 ();
 sg13g2_fill_2 FILLER_74_236 ();
 sg13g2_fill_1 FILLER_74_238 ();
 sg13g2_fill_1 FILLER_74_244 ();
 sg13g2_decap_8 FILLER_74_258 ();
 sg13g2_fill_2 FILLER_74_265 ();
 sg13g2_fill_2 FILLER_74_289 ();
 sg13g2_fill_2 FILLER_74_296 ();
 sg13g2_fill_1 FILLER_74_298 ();
 sg13g2_decap_8 FILLER_74_309 ();
 sg13g2_decap_8 FILLER_74_316 ();
 sg13g2_fill_1 FILLER_74_323 ();
 sg13g2_fill_2 FILLER_74_332 ();
 sg13g2_fill_1 FILLER_74_334 ();
 sg13g2_decap_8 FILLER_74_348 ();
 sg13g2_decap_8 FILLER_74_367 ();
 sg13g2_decap_4 FILLER_74_374 ();
 sg13g2_fill_2 FILLER_74_378 ();
 sg13g2_decap_8 FILLER_74_385 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_decap_8 FILLER_74_399 ();
 sg13g2_fill_2 FILLER_74_406 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_4 FILLER_75_84 ();
 sg13g2_fill_1 FILLER_75_88 ();
 sg13g2_fill_2 FILLER_75_96 ();
 sg13g2_fill_1 FILLER_75_98 ();
 sg13g2_fill_2 FILLER_75_120 ();
 sg13g2_fill_1 FILLER_75_122 ();
 sg13g2_fill_2 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_166 ();
 sg13g2_decap_4 FILLER_75_173 ();
 sg13g2_fill_2 FILLER_75_184 ();
 sg13g2_fill_1 FILLER_75_186 ();
 sg13g2_fill_1 FILLER_75_200 ();
 sg13g2_fill_1 FILLER_75_208 ();
 sg13g2_decap_4 FILLER_75_215 ();
 sg13g2_fill_2 FILLER_75_219 ();
 sg13g2_fill_1 FILLER_75_247 ();
 sg13g2_decap_4 FILLER_75_253 ();
 sg13g2_fill_2 FILLER_75_270 ();
 sg13g2_fill_1 FILLER_75_272 ();
 sg13g2_fill_2 FILLER_75_276 ();
 sg13g2_decap_4 FILLER_75_316 ();
 sg13g2_decap_8 FILLER_75_335 ();
 sg13g2_decap_8 FILLER_75_391 ();
 sg13g2_decap_8 FILLER_75_398 ();
 sg13g2_decap_4 FILLER_75_405 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_4 FILLER_76_100 ();
 sg13g2_fill_2 FILLER_76_110 ();
 sg13g2_decap_4 FILLER_76_158 ();
 sg13g2_fill_2 FILLER_76_181 ();
 sg13g2_fill_1 FILLER_76_255 ();
 sg13g2_fill_1 FILLER_76_261 ();
 sg13g2_decap_4 FILLER_76_289 ();
 sg13g2_fill_1 FILLER_76_293 ();
 sg13g2_decap_4 FILLER_76_324 ();
 sg13g2_fill_1 FILLER_76_339 ();
 sg13g2_decap_4 FILLER_76_345 ();
 sg13g2_fill_1 FILLER_76_349 ();
 sg13g2_fill_1 FILLER_76_368 ();
 sg13g2_fill_2 FILLER_76_379 ();
 sg13g2_decap_8 FILLER_76_386 ();
 sg13g2_decap_8 FILLER_76_393 ();
 sg13g2_decap_8 FILLER_76_400 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_fill_2 FILLER_77_84 ();
 sg13g2_fill_1 FILLER_77_86 ();
 sg13g2_fill_2 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_136 ();
 sg13g2_fill_2 FILLER_77_143 ();
 sg13g2_fill_1 FILLER_77_157 ();
 sg13g2_decap_4 FILLER_77_164 ();
 sg13g2_fill_2 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_195 ();
 sg13g2_fill_2 FILLER_77_202 ();
 sg13g2_fill_2 FILLER_77_207 ();
 sg13g2_fill_1 FILLER_77_209 ();
 sg13g2_decap_4 FILLER_77_213 ();
 sg13g2_fill_1 FILLER_77_217 ();
 sg13g2_decap_8 FILLER_77_222 ();
 sg13g2_decap_8 FILLER_77_229 ();
 sg13g2_fill_2 FILLER_77_236 ();
 sg13g2_decap_8 FILLER_77_244 ();
 sg13g2_fill_2 FILLER_77_251 ();
 sg13g2_fill_1 FILLER_77_253 ();
 sg13g2_fill_2 FILLER_77_267 ();
 sg13g2_fill_1 FILLER_77_269 ();
 sg13g2_decap_4 FILLER_77_286 ();
 sg13g2_fill_2 FILLER_77_312 ();
 sg13g2_decap_4 FILLER_77_322 ();
 sg13g2_decap_8 FILLER_77_351 ();
 sg13g2_fill_2 FILLER_77_358 ();
 sg13g2_decap_8 FILLER_77_389 ();
 sg13g2_decap_8 FILLER_77_396 ();
 sg13g2_decap_4 FILLER_77_403 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_fill_2 FILLER_78_91 ();
 sg13g2_fill_2 FILLER_78_103 ();
 sg13g2_fill_2 FILLER_78_121 ();
 sg13g2_fill_2 FILLER_78_149 ();
 sg13g2_decap_4 FILLER_78_169 ();
 sg13g2_fill_1 FILLER_78_197 ();
 sg13g2_decap_4 FILLER_78_243 ();
 sg13g2_decap_8 FILLER_78_272 ();
 sg13g2_fill_1 FILLER_78_279 ();
 sg13g2_decap_4 FILLER_78_290 ();
 sg13g2_fill_1 FILLER_78_294 ();
 sg13g2_fill_2 FILLER_78_308 ();
 sg13g2_fill_1 FILLER_78_310 ();
 sg13g2_decap_8 FILLER_78_344 ();
 sg13g2_fill_2 FILLER_78_364 ();
 sg13g2_fill_1 FILLER_78_366 ();
 sg13g2_decap_8 FILLER_78_376 ();
 sg13g2_decap_8 FILLER_78_383 ();
 sg13g2_decap_8 FILLER_78_390 ();
 sg13g2_decap_8 FILLER_78_397 ();
 sg13g2_decap_4 FILLER_78_404 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_4 FILLER_79_91 ();
 sg13g2_fill_2 FILLER_79_95 ();
 sg13g2_fill_1 FILLER_79_109 ();
 sg13g2_decap_8 FILLER_79_121 ();
 sg13g2_fill_2 FILLER_79_157 ();
 sg13g2_fill_2 FILLER_79_185 ();
 sg13g2_fill_1 FILLER_79_187 ();
 sg13g2_decap_8 FILLER_79_204 ();
 sg13g2_decap_8 FILLER_79_211 ();
 sg13g2_fill_1 FILLER_79_218 ();
 sg13g2_decap_8 FILLER_79_227 ();
 sg13g2_decap_4 FILLER_79_234 ();
 sg13g2_fill_1 FILLER_79_238 ();
 sg13g2_decap_4 FILLER_79_244 ();
 sg13g2_fill_2 FILLER_79_261 ();
 sg13g2_decap_8 FILLER_79_393 ();
 sg13g2_decap_8 FILLER_79_400 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_fill_1 FILLER_80_100 ();
 sg13g2_fill_2 FILLER_80_109 ();
 sg13g2_fill_1 FILLER_80_111 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_fill_2 FILLER_80_158 ();
 sg13g2_fill_1 FILLER_80_183 ();
 sg13g2_fill_1 FILLER_80_193 ();
 sg13g2_fill_1 FILLER_80_199 ();
 sg13g2_fill_2 FILLER_80_280 ();
 sg13g2_fill_1 FILLER_80_282 ();
 sg13g2_fill_2 FILLER_80_296 ();
 sg13g2_fill_2 FILLER_80_318 ();
 sg13g2_fill_2 FILLER_80_345 ();
 sg13g2_fill_1 FILLER_80_347 ();
 sg13g2_decap_4 FILLER_80_358 ();
 sg13g2_fill_2 FILLER_80_366 ();
 sg13g2_fill_2 FILLER_80_373 ();
 sg13g2_fill_1 FILLER_80_375 ();
 sg13g2_decap_8 FILLER_80_384 ();
 sg13g2_decap_8 FILLER_80_391 ();
 sg13g2_decap_8 FILLER_80_398 ();
 sg13g2_decap_4 FILLER_80_405 ();
 assign uio_oe[0] = net14;
 assign uio_oe[1] = net15;
 assign uio_oe[2] = net16;
 assign uio_oe[3] = net17;
 assign uio_oe[4] = net18;
 assign uio_oe[5] = net19;
 assign uio_oe[6] = net20;
 assign uio_oe[7] = net21;
 assign uio_out[0] = net22;
 assign uio_out[1] = net23;
 assign uio_out[2] = net24;
 assign uio_out[3] = net25;
 assign uio_out[4] = net26;
 assign uio_out[5] = net27;
 assign uio_out[6] = net28;
 assign uio_out[7] = net29;
endmodule

module tt_um_bilal_trng (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \TRNG.NOISE_SAMPLER.Sample_Out ;
 wire \TRNG.NOISE_SOURCE.Loop1.NOT2_OUT_TO_NAND1_IN2 ;
 wire \TRNG.NOISE_SOURCE.Loop2.NOT2_OUT_TO_NAND1_IN2 ;
 wire \TRNG.NOISE_SOURCE.Loop3.NOT2_OUT_TO_NAND1_IN2 ;
 wire \TRNG.NOISE_SOURCE.Loop4.NOT2_OUT_TO_NAND1_IN2 ;
 wire \TRNG.NOISE_SOURCE.Loop5.NOT2_OUT_TO_NAND1_IN2 ;
 wire \TRNG.NOISE_SOURCE.Noise_Source_Out ;
 wire \TRNG.Padded_Out[100] ;
 wire \TRNG.Padded_Out[101] ;
 wire \TRNG.Padded_Out[102] ;
 wire \TRNG.Padded_Out[103] ;
 wire \TRNG.Padded_Out[104] ;
 wire \TRNG.Padded_Out[105] ;
 wire \TRNG.Padded_Out[106] ;
 wire \TRNG.Padded_Out[107] ;
 wire \TRNG.Padded_Out[108] ;
 wire \TRNG.Padded_Out[109] ;
 wire \TRNG.Padded_Out[110] ;
 wire \TRNG.Padded_Out[111] ;
 wire \TRNG.Padded_Out[112] ;
 wire \TRNG.Padded_Out[113] ;
 wire \TRNG.Padded_Out[114] ;
 wire \TRNG.Padded_Out[115] ;
 wire \TRNG.Padded_Out[116] ;
 wire \TRNG.Padded_Out[117] ;
 wire \TRNG.Padded_Out[118] ;
 wire \TRNG.Padded_Out[119] ;
 wire \TRNG.Padded_Out[120] ;
 wire \TRNG.Padded_Out[121] ;
 wire \TRNG.Padded_Out[122] ;
 wire \TRNG.Padded_Out[123] ;
 wire \TRNG.Padded_Out[124] ;
 wire \TRNG.Padded_Out[125] ;
 wire \TRNG.Padded_Out[126] ;
 wire \TRNG.Padded_Out[127] ;
 wire \TRNG.Padded_Out[128] ;
 wire \TRNG.Padded_Out[129] ;
 wire \TRNG.Padded_Out[130] ;
 wire \TRNG.Padded_Out[131] ;
 wire \TRNG.Padded_Out[132] ;
 wire \TRNG.Padded_Out[133] ;
 wire \TRNG.Padded_Out[134] ;
 wire \TRNG.Padded_Out[135] ;
 wire \TRNG.Padded_Out[136] ;
 wire \TRNG.Padded_Out[137] ;
 wire \TRNG.Padded_Out[138] ;
 wire \TRNG.Padded_Out[139] ;
 wire \TRNG.Padded_Out[140] ;
 wire \TRNG.Padded_Out[141] ;
 wire \TRNG.Padded_Out[142] ;
 wire \TRNG.Padded_Out[143] ;
 wire \TRNG.Padded_Out[144] ;
 wire \TRNG.Padded_Out[145] ;
 wire \TRNG.Padded_Out[146] ;
 wire \TRNG.Padded_Out[147] ;
 wire \TRNG.Padded_Out[148] ;
 wire \TRNG.Padded_Out[149] ;
 wire \TRNG.Padded_Out[150] ;
 wire \TRNG.Padded_Out[151] ;
 wire \TRNG.Padded_Out[152] ;
 wire \TRNG.Padded_Out[153] ;
 wire \TRNG.Padded_Out[154] ;
 wire \TRNG.Padded_Out[155] ;
 wire \TRNG.Padded_Out[156] ;
 wire \TRNG.Padded_Out[157] ;
 wire \TRNG.Padded_Out[158] ;
 wire \TRNG.Padded_Out[159] ;
 wire \TRNG.Padded_Out[160] ;
 wire \TRNG.Padded_Out[161] ;
 wire \TRNG.Padded_Out[162] ;
 wire \TRNG.Padded_Out[163] ;
 wire \TRNG.Padded_Out[164] ;
 wire \TRNG.Padded_Out[165] ;
 wire \TRNG.Padded_Out[166] ;
 wire \TRNG.Padded_Out[167] ;
 wire \TRNG.Padded_Out[168] ;
 wire \TRNG.Padded_Out[169] ;
 wire \TRNG.Padded_Out[170] ;
 wire \TRNG.Padded_Out[171] ;
 wire \TRNG.Padded_Out[172] ;
 wire \TRNG.Padded_Out[173] ;
 wire \TRNG.Padded_Out[174] ;
 wire \TRNG.Padded_Out[175] ;
 wire \TRNG.Padded_Out[176] ;
 wire \TRNG.Padded_Out[177] ;
 wire \TRNG.Padded_Out[178] ;
 wire \TRNG.Padded_Out[179] ;
 wire \TRNG.Padded_Out[180] ;
 wire \TRNG.Padded_Out[181] ;
 wire \TRNG.Padded_Out[182] ;
 wire \TRNG.Padded_Out[183] ;
 wire \TRNG.Padded_Out[184] ;
 wire \TRNG.Padded_Out[185] ;
 wire \TRNG.Padded_Out[186] ;
 wire \TRNG.Padded_Out[187] ;
 wire \TRNG.Padded_Out[188] ;
 wire \TRNG.Padded_Out[189] ;
 wire \TRNG.Padded_Out[190] ;
 wire \TRNG.Padded_Out[191] ;
 wire \TRNG.Padded_Out[192] ;
 wire \TRNG.Padded_Out[193] ;
 wire \TRNG.Padded_Out[194] ;
 wire \TRNG.Padded_Out[195] ;
 wire \TRNG.Padded_Out[196] ;
 wire \TRNG.Padded_Out[197] ;
 wire \TRNG.Padded_Out[198] ;
 wire \TRNG.Padded_Out[199] ;
 wire \TRNG.Padded_Out[200] ;
 wire \TRNG.Padded_Out[201] ;
 wire \TRNG.Padded_Out[202] ;
 wire \TRNG.Padded_Out[203] ;
 wire \TRNG.Padded_Out[204] ;
 wire \TRNG.Padded_Out[205] ;
 wire \TRNG.Padded_Out[206] ;
 wire \TRNG.Padded_Out[207] ;
 wire \TRNG.Padded_Out[208] ;
 wire \TRNG.Padded_Out[209] ;
 wire \TRNG.Padded_Out[210] ;
 wire \TRNG.Padded_Out[211] ;
 wire \TRNG.Padded_Out[212] ;
 wire \TRNG.Padded_Out[213] ;
 wire \TRNG.Padded_Out[214] ;
 wire \TRNG.Padded_Out[215] ;
 wire \TRNG.Padded_Out[216] ;
 wire \TRNG.Padded_Out[217] ;
 wire \TRNG.Padded_Out[218] ;
 wire \TRNG.Padded_Out[219] ;
 wire \TRNG.Padded_Out[220] ;
 wire \TRNG.Padded_Out[221] ;
 wire \TRNG.Padded_Out[222] ;
 wire \TRNG.Padded_Out[223] ;
 wire \TRNG.Padded_Out[224] ;
 wire \TRNG.Padded_Out[225] ;
 wire \TRNG.Padded_Out[226] ;
 wire \TRNG.Padded_Out[227] ;
 wire \TRNG.Padded_Out[228] ;
 wire \TRNG.Padded_Out[229] ;
 wire \TRNG.Padded_Out[230] ;
 wire \TRNG.Padded_Out[231] ;
 wire \TRNG.Padded_Out[232] ;
 wire \TRNG.Padded_Out[233] ;
 wire \TRNG.Padded_Out[234] ;
 wire \TRNG.Padded_Out[235] ;
 wire \TRNG.Padded_Out[236] ;
 wire \TRNG.Padded_Out[237] ;
 wire \TRNG.Padded_Out[238] ;
 wire \TRNG.Padded_Out[239] ;
 wire \TRNG.Padded_Out[240] ;
 wire \TRNG.Padded_Out[241] ;
 wire \TRNG.Padded_Out[242] ;
 wire \TRNG.Padded_Out[243] ;
 wire \TRNG.Padded_Out[244] ;
 wire \TRNG.Padded_Out[245] ;
 wire \TRNG.Padded_Out[246] ;
 wire \TRNG.Padded_Out[247] ;
 wire \TRNG.Padded_Out[248] ;
 wire \TRNG.Padded_Out[249] ;
 wire \TRNG.Padded_Out[250] ;
 wire \TRNG.Padded_Out[251] ;
 wire \TRNG.Padded_Out[252] ;
 wire \TRNG.Padded_Out[253] ;
 wire \TRNG.Padded_Out[254] ;
 wire \TRNG.Padded_Out[255] ;
 wire \TRNG.Padded_Out[256] ;
 wire \TRNG.Padded_Out[257] ;
 wire \TRNG.Padded_Out[258] ;
 wire \TRNG.Padded_Out[259] ;
 wire \TRNG.Padded_Out[260] ;
 wire \TRNG.Padded_Out[261] ;
 wire \TRNG.Padded_Out[262] ;
 wire \TRNG.Padded_Out[263] ;
 wire \TRNG.Padded_Out[264] ;
 wire \TRNG.Padded_Out[265] ;
 wire \TRNG.Padded_Out[266] ;
 wire \TRNG.Padded_Out[267] ;
 wire \TRNG.Padded_Out[268] ;
 wire \TRNG.Padded_Out[269] ;
 wire \TRNG.Padded_Out[270] ;
 wire \TRNG.Padded_Out[271] ;
 wire \TRNG.Padded_Out[272] ;
 wire \TRNG.Padded_Out[273] ;
 wire \TRNG.Padded_Out[274] ;
 wire \TRNG.Padded_Out[275] ;
 wire \TRNG.Padded_Out[276] ;
 wire \TRNG.Padded_Out[277] ;
 wire \TRNG.Padded_Out[278] ;
 wire \TRNG.Padded_Out[279] ;
 wire \TRNG.Padded_Out[280] ;
 wire \TRNG.Padded_Out[281] ;
 wire \TRNG.Padded_Out[282] ;
 wire \TRNG.Padded_Out[283] ;
 wire \TRNG.Padded_Out[284] ;
 wire \TRNG.Padded_Out[285] ;
 wire \TRNG.Padded_Out[286] ;
 wire \TRNG.Padded_Out[287] ;
 wire \TRNG.Padded_Out[288] ;
 wire \TRNG.Padded_Out[289] ;
 wire \TRNG.Padded_Out[290] ;
 wire \TRNG.Padded_Out[291] ;
 wire \TRNG.Padded_Out[292] ;
 wire \TRNG.Padded_Out[293] ;
 wire \TRNG.Padded_Out[294] ;
 wire \TRNG.Padded_Out[295] ;
 wire \TRNG.Padded_Out[296] ;
 wire \TRNG.Padded_Out[297] ;
 wire \TRNG.Padded_Out[298] ;
 wire \TRNG.Padded_Out[299] ;
 wire \TRNG.Padded_Out[300] ;
 wire \TRNG.Padded_Out[301] ;
 wire \TRNG.Padded_Out[302] ;
 wire \TRNG.Padded_Out[303] ;
 wire \TRNG.Padded_Out[304] ;
 wire \TRNG.Padded_Out[305] ;
 wire \TRNG.Padded_Out[306] ;
 wire \TRNG.Padded_Out[307] ;
 wire \TRNG.Padded_Out[308] ;
 wire \TRNG.Padded_Out[309] ;
 wire \TRNG.Padded_Out[310] ;
 wire \TRNG.Padded_Out[311] ;
 wire \TRNG.Padded_Out[312] ;
 wire \TRNG.Padded_Out[313] ;
 wire \TRNG.Padded_Out[314] ;
 wire \TRNG.Padded_Out[315] ;
 wire \TRNG.Padded_Out[316] ;
 wire \TRNG.Padded_Out[317] ;
 wire \TRNG.Padded_Out[318] ;
 wire \TRNG.Padded_Out[319] ;
 wire \TRNG.Padded_Out[320] ;
 wire \TRNG.Padded_Out[321] ;
 wire \TRNG.Padded_Out[322] ;
 wire \TRNG.Padded_Out[323] ;
 wire \TRNG.Padded_Out[324] ;
 wire \TRNG.Padded_Out[325] ;
 wire \TRNG.Padded_Out[326] ;
 wire \TRNG.Padded_Out[327] ;
 wire \TRNG.Padded_Out[328] ;
 wire \TRNG.Padded_Out[329] ;
 wire \TRNG.Padded_Out[330] ;
 wire \TRNG.Padded_Out[331] ;
 wire \TRNG.Padded_Out[332] ;
 wire \TRNG.Padded_Out[333] ;
 wire \TRNG.Padded_Out[334] ;
 wire \TRNG.Padded_Out[335] ;
 wire \TRNG.Padded_Out[336] ;
 wire \TRNG.Padded_Out[337] ;
 wire \TRNG.Padded_Out[338] ;
 wire \TRNG.Padded_Out[339] ;
 wire \TRNG.Padded_Out[340] ;
 wire \TRNG.Padded_Out[341] ;
 wire \TRNG.Padded_Out[342] ;
 wire \TRNG.Padded_Out[343] ;
 wire \TRNG.Padded_Out[344] ;
 wire \TRNG.Padded_Out[345] ;
 wire \TRNG.Padded_Out[346] ;
 wire \TRNG.Padded_Out[347] ;
 wire \TRNG.Padded_Out[348] ;
 wire \TRNG.Padded_Out[349] ;
 wire \TRNG.Padded_Out[350] ;
 wire \TRNG.Padded_Out[351] ;
 wire \TRNG.Padded_Out[352] ;
 wire \TRNG.Padded_Out[353] ;
 wire \TRNG.Padded_Out[354] ;
 wire \TRNG.Padded_Out[355] ;
 wire \TRNG.Padded_Out[356] ;
 wire \TRNG.Padded_Out[357] ;
 wire \TRNG.Padded_Out[358] ;
 wire \TRNG.Padded_Out[359] ;
 wire \TRNG.Padded_Out[360] ;
 wire \TRNG.Padded_Out[361] ;
 wire \TRNG.Padded_Out[362] ;
 wire \TRNG.Padded_Out[363] ;
 wire \TRNG.Padded_Out[364] ;
 wire \TRNG.Padded_Out[365] ;
 wire \TRNG.Padded_Out[366] ;
 wire \TRNG.Padded_Out[367] ;
 wire \TRNG.Padded_Out[368] ;
 wire \TRNG.Padded_Out[369] ;
 wire \TRNG.Padded_Out[370] ;
 wire \TRNG.Padded_Out[371] ;
 wire \TRNG.Padded_Out[372] ;
 wire \TRNG.Padded_Out[373] ;
 wire \TRNG.Padded_Out[374] ;
 wire \TRNG.Padded_Out[375] ;
 wire \TRNG.Padded_Out[376] ;
 wire \TRNG.Padded_Out[377] ;
 wire \TRNG.Padded_Out[378] ;
 wire \TRNG.Padded_Out[379] ;
 wire \TRNG.Padded_Out[380] ;
 wire \TRNG.Padded_Out[381] ;
 wire \TRNG.Padded_Out[382] ;
 wire \TRNG.Padded_Out[383] ;
 wire \TRNG.Padded_Out[384] ;
 wire \TRNG.Padded_Out[385] ;
 wire \TRNG.Padded_Out[386] ;
 wire \TRNG.Padded_Out[387] ;
 wire \TRNG.Padded_Out[388] ;
 wire \TRNG.Padded_Out[389] ;
 wire \TRNG.Padded_Out[390] ;
 wire \TRNG.Padded_Out[391] ;
 wire \TRNG.Padded_Out[392] ;
 wire \TRNG.Padded_Out[393] ;
 wire \TRNG.Padded_Out[394] ;
 wire \TRNG.Padded_Out[395] ;
 wire \TRNG.Padded_Out[396] ;
 wire \TRNG.Padded_Out[397] ;
 wire \TRNG.Padded_Out[398] ;
 wire \TRNG.Padded_Out[399] ;
 wire \TRNG.Padded_Out[400] ;
 wire \TRNG.Padded_Out[401] ;
 wire \TRNG.Padded_Out[402] ;
 wire \TRNG.Padded_Out[403] ;
 wire \TRNG.Padded_Out[404] ;
 wire \TRNG.Padded_Out[405] ;
 wire \TRNG.Padded_Out[406] ;
 wire \TRNG.Padded_Out[407] ;
 wire \TRNG.Padded_Out[408] ;
 wire \TRNG.Padded_Out[409] ;
 wire \TRNG.Padded_Out[410] ;
 wire \TRNG.Padded_Out[411] ;
 wire \TRNG.Padded_Out[412] ;
 wire \TRNG.Padded_Out[413] ;
 wire \TRNG.Padded_Out[414] ;
 wire \TRNG.Padded_Out[415] ;
 wire \TRNG.Padded_Out[416] ;
 wire \TRNG.Padded_Out[417] ;
 wire \TRNG.Padded_Out[418] ;
 wire \TRNG.Padded_Out[419] ;
 wire \TRNG.Padded_Out[420] ;
 wire \TRNG.Padded_Out[421] ;
 wire \TRNG.Padded_Out[422] ;
 wire \TRNG.Padded_Out[423] ;
 wire \TRNG.Padded_Out[424] ;
 wire \TRNG.Padded_Out[425] ;
 wire \TRNG.Padded_Out[426] ;
 wire \TRNG.Padded_Out[427] ;
 wire \TRNG.Padded_Out[428] ;
 wire \TRNG.Padded_Out[429] ;
 wire \TRNG.Padded_Out[430] ;
 wire \TRNG.Padded_Out[431] ;
 wire \TRNG.Padded_Out[432] ;
 wire \TRNG.Padded_Out[433] ;
 wire \TRNG.Padded_Out[434] ;
 wire \TRNG.Padded_Out[435] ;
 wire \TRNG.Padded_Out[436] ;
 wire \TRNG.Padded_Out[437] ;
 wire \TRNG.Padded_Out[438] ;
 wire \TRNG.Padded_Out[439] ;
 wire \TRNG.Padded_Out[440] ;
 wire \TRNG.Padded_Out[441] ;
 wire \TRNG.Padded_Out[442] ;
 wire \TRNG.Padded_Out[443] ;
 wire \TRNG.Padded_Out[444] ;
 wire \TRNG.Padded_Out[445] ;
 wire \TRNG.Padded_Out[446] ;
 wire \TRNG.Padded_Out[447] ;
 wire \TRNG.Padded_Out[448] ;
 wire \TRNG.Padded_Out[449] ;
 wire \TRNG.Padded_Out[450] ;
 wire \TRNG.Padded_Out[451] ;
 wire \TRNG.Padded_Out[452] ;
 wire \TRNG.Padded_Out[453] ;
 wire \TRNG.Padded_Out[454] ;
 wire \TRNG.Padded_Out[455] ;
 wire \TRNG.Padded_Out[456] ;
 wire \TRNG.Padded_Out[457] ;
 wire \TRNG.Padded_Out[458] ;
 wire \TRNG.Padded_Out[459] ;
 wire \TRNG.Padded_Out[460] ;
 wire \TRNG.Padded_Out[461] ;
 wire \TRNG.Padded_Out[462] ;
 wire \TRNG.Padded_Out[463] ;
 wire \TRNG.Padded_Out[464] ;
 wire \TRNG.Padded_Out[465] ;
 wire \TRNG.Padded_Out[466] ;
 wire \TRNG.Padded_Out[467] ;
 wire \TRNG.Padded_Out[468] ;
 wire \TRNG.Padded_Out[469] ;
 wire \TRNG.Padded_Out[470] ;
 wire \TRNG.Padded_Out[471] ;
 wire \TRNG.Padded_Out[472] ;
 wire \TRNG.Padded_Out[473] ;
 wire \TRNG.Padded_Out[474] ;
 wire \TRNG.Padded_Out[475] ;
 wire \TRNG.Padded_Out[476] ;
 wire \TRNG.Padded_Out[477] ;
 wire \TRNG.Padded_Out[478] ;
 wire \TRNG.Padded_Out[479] ;
 wire \TRNG.Padded_Out[480] ;
 wire \TRNG.Padded_Out[481] ;
 wire \TRNG.Padded_Out[482] ;
 wire \TRNG.Padded_Out[483] ;
 wire \TRNG.Padded_Out[484] ;
 wire \TRNG.Padded_Out[485] ;
 wire \TRNG.Padded_Out[486] ;
 wire \TRNG.Padded_Out[487] ;
 wire \TRNG.Padded_Out[488] ;
 wire \TRNG.Padded_Out[489] ;
 wire \TRNG.Padded_Out[490] ;
 wire \TRNG.Padded_Out[491] ;
 wire \TRNG.Padded_Out[492] ;
 wire \TRNG.Padded_Out[493] ;
 wire \TRNG.Padded_Out[494] ;
 wire \TRNG.Padded_Out[495] ;
 wire \TRNG.Padded_Out[496] ;
 wire \TRNG.Padded_Out[497] ;
 wire \TRNG.Padded_Out[498] ;
 wire \TRNG.Padded_Out[499] ;
 wire \TRNG.Padded_Out[500] ;
 wire \TRNG.Padded_Out[501] ;
 wire \TRNG.Padded_Out[502] ;
 wire \TRNG.Padded_Out[503] ;
 wire \TRNG.Padded_Out[504] ;
 wire \TRNG.Padded_Out[505] ;
 wire \TRNG.Padded_Out[506] ;
 wire \TRNG.Padded_Out[507] ;
 wire \TRNG.Padded_Out[508] ;
 wire \TRNG.Padded_Out[509] ;
 wire \TRNG.Padded_Out[510] ;
 wire \TRNG.Padded_Out[511] ;
 wire \TRNG.Padded_Out[64] ;
 wire \TRNG.Padded_Out[65] ;
 wire \TRNG.Padded_Out[66] ;
 wire \TRNG.Padded_Out[67] ;
 wire \TRNG.Padded_Out[68] ;
 wire \TRNG.Padded_Out[69] ;
 wire \TRNG.Padded_Out[70] ;
 wire \TRNG.Padded_Out[71] ;
 wire \TRNG.Padded_Out[72] ;
 wire \TRNG.Padded_Out[73] ;
 wire \TRNG.Padded_Out[74] ;
 wire \TRNG.Padded_Out[75] ;
 wire \TRNG.Padded_Out[76] ;
 wire \TRNG.Padded_Out[77] ;
 wire \TRNG.Padded_Out[78] ;
 wire \TRNG.Padded_Out[79] ;
 wire \TRNG.Padded_Out[80] ;
 wire \TRNG.Padded_Out[81] ;
 wire \TRNG.Padded_Out[82] ;
 wire \TRNG.Padded_Out[83] ;
 wire \TRNG.Padded_Out[84] ;
 wire \TRNG.Padded_Out[85] ;
 wire \TRNG.Padded_Out[86] ;
 wire \TRNG.Padded_Out[87] ;
 wire \TRNG.Padded_Out[88] ;
 wire \TRNG.Padded_Out[89] ;
 wire \TRNG.Padded_Out[90] ;
 wire \TRNG.Padded_Out[91] ;
 wire \TRNG.Padded_Out[92] ;
 wire \TRNG.Padded_Out[93] ;
 wire \TRNG.Padded_Out[94] ;
 wire \TRNG.Padded_Out[95] ;
 wire \TRNG.Padded_Out[96] ;
 wire \TRNG.Padded_Out[97] ;
 wire \TRNG.Padded_Out[98] ;
 wire \TRNG.Padded_Out[99] ;
 wire \TRNG.Repetition_Count_Test.count[0] ;
 wire \TRNG.Repetition_Count_Test.count[1] ;
 wire \TRNG.Repetition_Count_Test.count[2] ;
 wire \TRNG.Repetition_Count_Test.count[3] ;
 wire \TRNG.Repetition_Count_Test.count[4] ;
 wire \TRNG.Repetition_Count_Test.count[5] ;
 wire \TRNG.Repetition_Count_Test.failure ;
 wire \TRNG.Repetition_Count_Test.prev_bit ;
 wire \TRNG.UART_Tx ;
 wire \TRNG.Word_Out[0] ;
 wire \TRNG.Word_Out[100] ;
 wire \TRNG.Word_Out[101] ;
 wire \TRNG.Word_Out[102] ;
 wire \TRNG.Word_Out[103] ;
 wire \TRNG.Word_Out[104] ;
 wire \TRNG.Word_Out[105] ;
 wire \TRNG.Word_Out[106] ;
 wire \TRNG.Word_Out[107] ;
 wire \TRNG.Word_Out[108] ;
 wire \TRNG.Word_Out[109] ;
 wire \TRNG.Word_Out[10] ;
 wire \TRNG.Word_Out[110] ;
 wire \TRNG.Word_Out[111] ;
 wire \TRNG.Word_Out[112] ;
 wire \TRNG.Word_Out[113] ;
 wire \TRNG.Word_Out[114] ;
 wire \TRNG.Word_Out[115] ;
 wire \TRNG.Word_Out[116] ;
 wire \TRNG.Word_Out[117] ;
 wire \TRNG.Word_Out[118] ;
 wire \TRNG.Word_Out[119] ;
 wire \TRNG.Word_Out[11] ;
 wire \TRNG.Word_Out[120] ;
 wire \TRNG.Word_Out[121] ;
 wire \TRNG.Word_Out[122] ;
 wire \TRNG.Word_Out[123] ;
 wire \TRNG.Word_Out[124] ;
 wire \TRNG.Word_Out[125] ;
 wire \TRNG.Word_Out[126] ;
 wire \TRNG.Word_Out[127] ;
 wire \TRNG.Word_Out[128] ;
 wire \TRNG.Word_Out[129] ;
 wire \TRNG.Word_Out[12] ;
 wire \TRNG.Word_Out[130] ;
 wire \TRNG.Word_Out[131] ;
 wire \TRNG.Word_Out[132] ;
 wire \TRNG.Word_Out[133] ;
 wire \TRNG.Word_Out[134] ;
 wire \TRNG.Word_Out[135] ;
 wire \TRNG.Word_Out[136] ;
 wire \TRNG.Word_Out[137] ;
 wire \TRNG.Word_Out[138] ;
 wire \TRNG.Word_Out[139] ;
 wire \TRNG.Word_Out[13] ;
 wire \TRNG.Word_Out[140] ;
 wire \TRNG.Word_Out[141] ;
 wire \TRNG.Word_Out[142] ;
 wire \TRNG.Word_Out[143] ;
 wire \TRNG.Word_Out[144] ;
 wire \TRNG.Word_Out[145] ;
 wire \TRNG.Word_Out[146] ;
 wire \TRNG.Word_Out[147] ;
 wire \TRNG.Word_Out[148] ;
 wire \TRNG.Word_Out[149] ;
 wire \TRNG.Word_Out[14] ;
 wire \TRNG.Word_Out[150] ;
 wire \TRNG.Word_Out[151] ;
 wire \TRNG.Word_Out[152] ;
 wire \TRNG.Word_Out[153] ;
 wire \TRNG.Word_Out[154] ;
 wire \TRNG.Word_Out[155] ;
 wire \TRNG.Word_Out[156] ;
 wire \TRNG.Word_Out[157] ;
 wire \TRNG.Word_Out[158] ;
 wire \TRNG.Word_Out[159] ;
 wire \TRNG.Word_Out[15] ;
 wire \TRNG.Word_Out[160] ;
 wire \TRNG.Word_Out[161] ;
 wire \TRNG.Word_Out[162] ;
 wire \TRNG.Word_Out[163] ;
 wire \TRNG.Word_Out[164] ;
 wire \TRNG.Word_Out[165] ;
 wire \TRNG.Word_Out[166] ;
 wire \TRNG.Word_Out[167] ;
 wire \TRNG.Word_Out[168] ;
 wire \TRNG.Word_Out[169] ;
 wire \TRNG.Word_Out[16] ;
 wire \TRNG.Word_Out[170] ;
 wire \TRNG.Word_Out[171] ;
 wire \TRNG.Word_Out[172] ;
 wire \TRNG.Word_Out[173] ;
 wire \TRNG.Word_Out[174] ;
 wire \TRNG.Word_Out[175] ;
 wire \TRNG.Word_Out[176] ;
 wire \TRNG.Word_Out[177] ;
 wire \TRNG.Word_Out[178] ;
 wire \TRNG.Word_Out[179] ;
 wire \TRNG.Word_Out[17] ;
 wire \TRNG.Word_Out[180] ;
 wire \TRNG.Word_Out[181] ;
 wire \TRNG.Word_Out[182] ;
 wire \TRNG.Word_Out[183] ;
 wire \TRNG.Word_Out[184] ;
 wire \TRNG.Word_Out[185] ;
 wire \TRNG.Word_Out[186] ;
 wire \TRNG.Word_Out[187] ;
 wire \TRNG.Word_Out[188] ;
 wire \TRNG.Word_Out[189] ;
 wire \TRNG.Word_Out[18] ;
 wire \TRNG.Word_Out[190] ;
 wire \TRNG.Word_Out[191] ;
 wire \TRNG.Word_Out[192] ;
 wire \TRNG.Word_Out[193] ;
 wire \TRNG.Word_Out[194] ;
 wire \TRNG.Word_Out[195] ;
 wire \TRNG.Word_Out[196] ;
 wire \TRNG.Word_Out[197] ;
 wire \TRNG.Word_Out[198] ;
 wire \TRNG.Word_Out[199] ;
 wire \TRNG.Word_Out[19] ;
 wire \TRNG.Word_Out[1] ;
 wire \TRNG.Word_Out[200] ;
 wire \TRNG.Word_Out[201] ;
 wire \TRNG.Word_Out[202] ;
 wire \TRNG.Word_Out[203] ;
 wire \TRNG.Word_Out[204] ;
 wire \TRNG.Word_Out[205] ;
 wire \TRNG.Word_Out[206] ;
 wire \TRNG.Word_Out[207] ;
 wire \TRNG.Word_Out[208] ;
 wire \TRNG.Word_Out[209] ;
 wire \TRNG.Word_Out[20] ;
 wire \TRNG.Word_Out[210] ;
 wire \TRNG.Word_Out[211] ;
 wire \TRNG.Word_Out[212] ;
 wire \TRNG.Word_Out[213] ;
 wire \TRNG.Word_Out[214] ;
 wire \TRNG.Word_Out[215] ;
 wire \TRNG.Word_Out[216] ;
 wire \TRNG.Word_Out[217] ;
 wire \TRNG.Word_Out[218] ;
 wire \TRNG.Word_Out[219] ;
 wire \TRNG.Word_Out[21] ;
 wire \TRNG.Word_Out[220] ;
 wire \TRNG.Word_Out[221] ;
 wire \TRNG.Word_Out[222] ;
 wire \TRNG.Word_Out[223] ;
 wire \TRNG.Word_Out[224] ;
 wire \TRNG.Word_Out[225] ;
 wire \TRNG.Word_Out[226] ;
 wire \TRNG.Word_Out[227] ;
 wire \TRNG.Word_Out[228] ;
 wire \TRNG.Word_Out[229] ;
 wire \TRNG.Word_Out[22] ;
 wire \TRNG.Word_Out[230] ;
 wire \TRNG.Word_Out[231] ;
 wire \TRNG.Word_Out[232] ;
 wire \TRNG.Word_Out[233] ;
 wire \TRNG.Word_Out[234] ;
 wire \TRNG.Word_Out[235] ;
 wire \TRNG.Word_Out[236] ;
 wire \TRNG.Word_Out[237] ;
 wire \TRNG.Word_Out[238] ;
 wire \TRNG.Word_Out[239] ;
 wire \TRNG.Word_Out[23] ;
 wire \TRNG.Word_Out[240] ;
 wire \TRNG.Word_Out[241] ;
 wire \TRNG.Word_Out[242] ;
 wire \TRNG.Word_Out[243] ;
 wire \TRNG.Word_Out[244] ;
 wire \TRNG.Word_Out[245] ;
 wire \TRNG.Word_Out[246] ;
 wire \TRNG.Word_Out[247] ;
 wire \TRNG.Word_Out[248] ;
 wire \TRNG.Word_Out[249] ;
 wire \TRNG.Word_Out[24] ;
 wire \TRNG.Word_Out[250] ;
 wire \TRNG.Word_Out[251] ;
 wire \TRNG.Word_Out[252] ;
 wire \TRNG.Word_Out[253] ;
 wire \TRNG.Word_Out[254] ;
 wire \TRNG.Word_Out[255] ;
 wire \TRNG.Word_Out[256] ;
 wire \TRNG.Word_Out[257] ;
 wire \TRNG.Word_Out[258] ;
 wire \TRNG.Word_Out[259] ;
 wire \TRNG.Word_Out[25] ;
 wire \TRNG.Word_Out[260] ;
 wire \TRNG.Word_Out[261] ;
 wire \TRNG.Word_Out[262] ;
 wire \TRNG.Word_Out[263] ;
 wire \TRNG.Word_Out[264] ;
 wire \TRNG.Word_Out[265] ;
 wire \TRNG.Word_Out[266] ;
 wire \TRNG.Word_Out[267] ;
 wire \TRNG.Word_Out[268] ;
 wire \TRNG.Word_Out[269] ;
 wire \TRNG.Word_Out[26] ;
 wire \TRNG.Word_Out[270] ;
 wire \TRNG.Word_Out[271] ;
 wire \TRNG.Word_Out[272] ;
 wire \TRNG.Word_Out[273] ;
 wire \TRNG.Word_Out[274] ;
 wire \TRNG.Word_Out[275] ;
 wire \TRNG.Word_Out[276] ;
 wire \TRNG.Word_Out[277] ;
 wire \TRNG.Word_Out[278] ;
 wire \TRNG.Word_Out[279] ;
 wire \TRNG.Word_Out[27] ;
 wire \TRNG.Word_Out[280] ;
 wire \TRNG.Word_Out[281] ;
 wire \TRNG.Word_Out[282] ;
 wire \TRNG.Word_Out[283] ;
 wire \TRNG.Word_Out[284] ;
 wire \TRNG.Word_Out[285] ;
 wire \TRNG.Word_Out[286] ;
 wire \TRNG.Word_Out[287] ;
 wire \TRNG.Word_Out[288] ;
 wire \TRNG.Word_Out[289] ;
 wire \TRNG.Word_Out[28] ;
 wire \TRNG.Word_Out[290] ;
 wire \TRNG.Word_Out[291] ;
 wire \TRNG.Word_Out[292] ;
 wire \TRNG.Word_Out[293] ;
 wire \TRNG.Word_Out[294] ;
 wire \TRNG.Word_Out[295] ;
 wire \TRNG.Word_Out[296] ;
 wire \TRNG.Word_Out[297] ;
 wire \TRNG.Word_Out[298] ;
 wire \TRNG.Word_Out[299] ;
 wire \TRNG.Word_Out[29] ;
 wire \TRNG.Word_Out[2] ;
 wire \TRNG.Word_Out[300] ;
 wire \TRNG.Word_Out[301] ;
 wire \TRNG.Word_Out[302] ;
 wire \TRNG.Word_Out[303] ;
 wire \TRNG.Word_Out[304] ;
 wire \TRNG.Word_Out[305] ;
 wire \TRNG.Word_Out[306] ;
 wire \TRNG.Word_Out[307] ;
 wire \TRNG.Word_Out[308] ;
 wire \TRNG.Word_Out[309] ;
 wire \TRNG.Word_Out[30] ;
 wire \TRNG.Word_Out[310] ;
 wire \TRNG.Word_Out[311] ;
 wire \TRNG.Word_Out[312] ;
 wire \TRNG.Word_Out[313] ;
 wire \TRNG.Word_Out[314] ;
 wire \TRNG.Word_Out[315] ;
 wire \TRNG.Word_Out[316] ;
 wire \TRNG.Word_Out[317] ;
 wire \TRNG.Word_Out[318] ;
 wire \TRNG.Word_Out[319] ;
 wire \TRNG.Word_Out[31] ;
 wire \TRNG.Word_Out[320] ;
 wire \TRNG.Word_Out[321] ;
 wire \TRNG.Word_Out[322] ;
 wire \TRNG.Word_Out[323] ;
 wire \TRNG.Word_Out[324] ;
 wire \TRNG.Word_Out[325] ;
 wire \TRNG.Word_Out[326] ;
 wire \TRNG.Word_Out[327] ;
 wire \TRNG.Word_Out[328] ;
 wire \TRNG.Word_Out[329] ;
 wire \TRNG.Word_Out[32] ;
 wire \TRNG.Word_Out[330] ;
 wire \TRNG.Word_Out[331] ;
 wire \TRNG.Word_Out[332] ;
 wire \TRNG.Word_Out[333] ;
 wire \TRNG.Word_Out[334] ;
 wire \TRNG.Word_Out[335] ;
 wire \TRNG.Word_Out[336] ;
 wire \TRNG.Word_Out[337] ;
 wire \TRNG.Word_Out[338] ;
 wire \TRNG.Word_Out[339] ;
 wire \TRNG.Word_Out[33] ;
 wire \TRNG.Word_Out[340] ;
 wire \TRNG.Word_Out[341] ;
 wire \TRNG.Word_Out[342] ;
 wire \TRNG.Word_Out[343] ;
 wire \TRNG.Word_Out[344] ;
 wire \TRNG.Word_Out[345] ;
 wire \TRNG.Word_Out[346] ;
 wire \TRNG.Word_Out[347] ;
 wire \TRNG.Word_Out[348] ;
 wire \TRNG.Word_Out[349] ;
 wire \TRNG.Word_Out[34] ;
 wire \TRNG.Word_Out[350] ;
 wire \TRNG.Word_Out[351] ;
 wire \TRNG.Word_Out[352] ;
 wire \TRNG.Word_Out[353] ;
 wire \TRNG.Word_Out[354] ;
 wire \TRNG.Word_Out[355] ;
 wire \TRNG.Word_Out[356] ;
 wire \TRNG.Word_Out[357] ;
 wire \TRNG.Word_Out[358] ;
 wire \TRNG.Word_Out[359] ;
 wire \TRNG.Word_Out[35] ;
 wire \TRNG.Word_Out[360] ;
 wire \TRNG.Word_Out[361] ;
 wire \TRNG.Word_Out[362] ;
 wire \TRNG.Word_Out[363] ;
 wire \TRNG.Word_Out[364] ;
 wire \TRNG.Word_Out[365] ;
 wire \TRNG.Word_Out[366] ;
 wire \TRNG.Word_Out[367] ;
 wire \TRNG.Word_Out[368] ;
 wire \TRNG.Word_Out[369] ;
 wire \TRNG.Word_Out[36] ;
 wire \TRNG.Word_Out[370] ;
 wire \TRNG.Word_Out[371] ;
 wire \TRNG.Word_Out[372] ;
 wire \TRNG.Word_Out[373] ;
 wire \TRNG.Word_Out[374] ;
 wire \TRNG.Word_Out[375] ;
 wire \TRNG.Word_Out[376] ;
 wire \TRNG.Word_Out[377] ;
 wire \TRNG.Word_Out[378] ;
 wire \TRNG.Word_Out[379] ;
 wire \TRNG.Word_Out[37] ;
 wire \TRNG.Word_Out[380] ;
 wire \TRNG.Word_Out[381] ;
 wire \TRNG.Word_Out[382] ;
 wire \TRNG.Word_Out[383] ;
 wire \TRNG.Word_Out[384] ;
 wire \TRNG.Word_Out[385] ;
 wire \TRNG.Word_Out[386] ;
 wire \TRNG.Word_Out[387] ;
 wire \TRNG.Word_Out[388] ;
 wire \TRNG.Word_Out[389] ;
 wire \TRNG.Word_Out[38] ;
 wire \TRNG.Word_Out[390] ;
 wire \TRNG.Word_Out[391] ;
 wire \TRNG.Word_Out[392] ;
 wire \TRNG.Word_Out[393] ;
 wire \TRNG.Word_Out[394] ;
 wire \TRNG.Word_Out[395] ;
 wire \TRNG.Word_Out[396] ;
 wire \TRNG.Word_Out[397] ;
 wire \TRNG.Word_Out[398] ;
 wire \TRNG.Word_Out[399] ;
 wire \TRNG.Word_Out[39] ;
 wire \TRNG.Word_Out[3] ;
 wire \TRNG.Word_Out[400] ;
 wire \TRNG.Word_Out[401] ;
 wire \TRNG.Word_Out[402] ;
 wire \TRNG.Word_Out[403] ;
 wire \TRNG.Word_Out[404] ;
 wire \TRNG.Word_Out[405] ;
 wire \TRNG.Word_Out[406] ;
 wire \TRNG.Word_Out[407] ;
 wire \TRNG.Word_Out[408] ;
 wire \TRNG.Word_Out[409] ;
 wire \TRNG.Word_Out[40] ;
 wire \TRNG.Word_Out[410] ;
 wire \TRNG.Word_Out[411] ;
 wire \TRNG.Word_Out[412] ;
 wire \TRNG.Word_Out[413] ;
 wire \TRNG.Word_Out[414] ;
 wire \TRNG.Word_Out[415] ;
 wire \TRNG.Word_Out[416] ;
 wire \TRNG.Word_Out[417] ;
 wire \TRNG.Word_Out[418] ;
 wire \TRNG.Word_Out[419] ;
 wire \TRNG.Word_Out[41] ;
 wire \TRNG.Word_Out[420] ;
 wire \TRNG.Word_Out[421] ;
 wire \TRNG.Word_Out[422] ;
 wire \TRNG.Word_Out[423] ;
 wire \TRNG.Word_Out[424] ;
 wire \TRNG.Word_Out[425] ;
 wire \TRNG.Word_Out[426] ;
 wire \TRNG.Word_Out[427] ;
 wire \TRNG.Word_Out[428] ;
 wire \TRNG.Word_Out[429] ;
 wire \TRNG.Word_Out[42] ;
 wire \TRNG.Word_Out[430] ;
 wire \TRNG.Word_Out[431] ;
 wire \TRNG.Word_Out[432] ;
 wire \TRNG.Word_Out[433] ;
 wire \TRNG.Word_Out[434] ;
 wire \TRNG.Word_Out[435] ;
 wire \TRNG.Word_Out[436] ;
 wire \TRNG.Word_Out[437] ;
 wire \TRNG.Word_Out[438] ;
 wire \TRNG.Word_Out[439] ;
 wire \TRNG.Word_Out[43] ;
 wire \TRNG.Word_Out[440] ;
 wire \TRNG.Word_Out[441] ;
 wire \TRNG.Word_Out[442] ;
 wire \TRNG.Word_Out[443] ;
 wire \TRNG.Word_Out[444] ;
 wire \TRNG.Word_Out[445] ;
 wire \TRNG.Word_Out[446] ;
 wire \TRNG.Word_Out[44] ;
 wire \TRNG.Word_Out[45] ;
 wire \TRNG.Word_Out[46] ;
 wire \TRNG.Word_Out[47] ;
 wire \TRNG.Word_Out[48] ;
 wire \TRNG.Word_Out[49] ;
 wire \TRNG.Word_Out[4] ;
 wire \TRNG.Word_Out[50] ;
 wire \TRNG.Word_Out[51] ;
 wire \TRNG.Word_Out[52] ;
 wire \TRNG.Word_Out[53] ;
 wire \TRNG.Word_Out[54] ;
 wire \TRNG.Word_Out[55] ;
 wire \TRNG.Word_Out[56] ;
 wire \TRNG.Word_Out[57] ;
 wire \TRNG.Word_Out[58] ;
 wire \TRNG.Word_Out[59] ;
 wire \TRNG.Word_Out[5] ;
 wire \TRNG.Word_Out[60] ;
 wire \TRNG.Word_Out[61] ;
 wire \TRNG.Word_Out[62] ;
 wire \TRNG.Word_Out[63] ;
 wire \TRNG.Word_Out[64] ;
 wire \TRNG.Word_Out[65] ;
 wire \TRNG.Word_Out[66] ;
 wire \TRNG.Word_Out[67] ;
 wire \TRNG.Word_Out[68] ;
 wire \TRNG.Word_Out[69] ;
 wire \TRNG.Word_Out[6] ;
 wire \TRNG.Word_Out[70] ;
 wire \TRNG.Word_Out[71] ;
 wire \TRNG.Word_Out[72] ;
 wire \TRNG.Word_Out[73] ;
 wire \TRNG.Word_Out[74] ;
 wire \TRNG.Word_Out[75] ;
 wire \TRNG.Word_Out[76] ;
 wire \TRNG.Word_Out[77] ;
 wire \TRNG.Word_Out[78] ;
 wire \TRNG.Word_Out[79] ;
 wire \TRNG.Word_Out[7] ;
 wire \TRNG.Word_Out[80] ;
 wire \TRNG.Word_Out[81] ;
 wire \TRNG.Word_Out[82] ;
 wire \TRNG.Word_Out[83] ;
 wire \TRNG.Word_Out[84] ;
 wire \TRNG.Word_Out[85] ;
 wire \TRNG.Word_Out[86] ;
 wire \TRNG.Word_Out[87] ;
 wire \TRNG.Word_Out[88] ;
 wire \TRNG.Word_Out[89] ;
 wire \TRNG.Word_Out[8] ;
 wire \TRNG.Word_Out[90] ;
 wire \TRNG.Word_Out[91] ;
 wire \TRNG.Word_Out[92] ;
 wire \TRNG.Word_Out[93] ;
 wire \TRNG.Word_Out[94] ;
 wire \TRNG.Word_Out[95] ;
 wire \TRNG.Word_Out[96] ;
 wire \TRNG.Word_Out[97] ;
 wire \TRNG.Word_Out[98] ;
 wire \TRNG.Word_Out[99] ;
 wire \TRNG.Word_Out[9] ;
 wire \TRNG.Word_Valid ;
 wire \TRNG.bit_counter[0] ;
 wire \TRNG.bit_counter[1] ;
 wire \TRNG.bit_counter[2] ;
 wire \TRNG.bit_counter[3] ;
 wire \TRNG.bit_counter[4] ;
 wire \TRNG.bit_counter[5] ;
 wire \TRNG.bit_counter[6] ;
 wire \TRNG.bit_counter[7] ;
 wire \TRNG.bit_counter[8] ;
 wire \TRNG.chunk_index[0] ;
 wire \TRNG.chunk_index[1] ;
 wire \TRNG.chunk_index[2] ;
 wire \TRNG.chunk_index[3] ;
 wire \TRNG.chunk_index[4] ;
 wire \TRNG.chunk_reg[0] ;
 wire \TRNG.chunk_reg[1] ;
 wire \TRNG.chunk_reg[2] ;
 wire \TRNG.chunk_reg[3] ;
 wire \TRNG.chunk_reg[4] ;
 wire \TRNG.chunk_reg[5] ;
 wire \TRNG.chunk_reg[6] ;
 wire \TRNG.chunk_reg[7] ;
 wire \TRNG.ctrl_mode_sync[0] ;
 wire \TRNG.ctrl_mode_sync[1] ;
 wire \TRNG.discard ;
 wire \TRNG.hash[0] ;
 wire \TRNG.hash[100] ;
 wire \TRNG.hash[101] ;
 wire \TRNG.hash[102] ;
 wire \TRNG.hash[103] ;
 wire \TRNG.hash[104] ;
 wire \TRNG.hash[105] ;
 wire \TRNG.hash[106] ;
 wire \TRNG.hash[107] ;
 wire \TRNG.hash[108] ;
 wire \TRNG.hash[109] ;
 wire \TRNG.hash[10] ;
 wire \TRNG.hash[110] ;
 wire \TRNG.hash[111] ;
 wire \TRNG.hash[112] ;
 wire \TRNG.hash[113] ;
 wire \TRNG.hash[114] ;
 wire \TRNG.hash[115] ;
 wire \TRNG.hash[116] ;
 wire \TRNG.hash[117] ;
 wire \TRNG.hash[118] ;
 wire \TRNG.hash[119] ;
 wire \TRNG.hash[11] ;
 wire \TRNG.hash[120] ;
 wire \TRNG.hash[121] ;
 wire \TRNG.hash[122] ;
 wire \TRNG.hash[123] ;
 wire \TRNG.hash[124] ;
 wire \TRNG.hash[125] ;
 wire \TRNG.hash[126] ;
 wire \TRNG.hash[127] ;
 wire \TRNG.hash[128] ;
 wire \TRNG.hash[129] ;
 wire \TRNG.hash[12] ;
 wire \TRNG.hash[130] ;
 wire \TRNG.hash[131] ;
 wire \TRNG.hash[132] ;
 wire \TRNG.hash[133] ;
 wire \TRNG.hash[134] ;
 wire \TRNG.hash[135] ;
 wire \TRNG.hash[136] ;
 wire \TRNG.hash[137] ;
 wire \TRNG.hash[138] ;
 wire \TRNG.hash[139] ;
 wire \TRNG.hash[13] ;
 wire \TRNG.hash[140] ;
 wire \TRNG.hash[141] ;
 wire \TRNG.hash[142] ;
 wire \TRNG.hash[143] ;
 wire \TRNG.hash[144] ;
 wire \TRNG.hash[145] ;
 wire \TRNG.hash[146] ;
 wire \TRNG.hash[147] ;
 wire \TRNG.hash[148] ;
 wire \TRNG.hash[149] ;
 wire \TRNG.hash[14] ;
 wire \TRNG.hash[150] ;
 wire \TRNG.hash[151] ;
 wire \TRNG.hash[152] ;
 wire \TRNG.hash[153] ;
 wire \TRNG.hash[154] ;
 wire \TRNG.hash[155] ;
 wire \TRNG.hash[156] ;
 wire \TRNG.hash[157] ;
 wire \TRNG.hash[158] ;
 wire \TRNG.hash[159] ;
 wire \TRNG.hash[15] ;
 wire \TRNG.hash[160] ;
 wire \TRNG.hash[161] ;
 wire \TRNG.hash[162] ;
 wire \TRNG.hash[163] ;
 wire \TRNG.hash[164] ;
 wire \TRNG.hash[165] ;
 wire \TRNG.hash[166] ;
 wire \TRNG.hash[167] ;
 wire \TRNG.hash[168] ;
 wire \TRNG.hash[169] ;
 wire \TRNG.hash[16] ;
 wire \TRNG.hash[170] ;
 wire \TRNG.hash[171] ;
 wire \TRNG.hash[172] ;
 wire \TRNG.hash[173] ;
 wire \TRNG.hash[174] ;
 wire \TRNG.hash[175] ;
 wire \TRNG.hash[176] ;
 wire \TRNG.hash[177] ;
 wire \TRNG.hash[178] ;
 wire \TRNG.hash[179] ;
 wire \TRNG.hash[17] ;
 wire \TRNG.hash[180] ;
 wire \TRNG.hash[181] ;
 wire \TRNG.hash[182] ;
 wire \TRNG.hash[183] ;
 wire \TRNG.hash[184] ;
 wire \TRNG.hash[185] ;
 wire \TRNG.hash[186] ;
 wire \TRNG.hash[187] ;
 wire \TRNG.hash[188] ;
 wire \TRNG.hash[189] ;
 wire \TRNG.hash[18] ;
 wire \TRNG.hash[190] ;
 wire \TRNG.hash[191] ;
 wire \TRNG.hash[192] ;
 wire \TRNG.hash[193] ;
 wire \TRNG.hash[194] ;
 wire \TRNG.hash[195] ;
 wire \TRNG.hash[196] ;
 wire \TRNG.hash[197] ;
 wire \TRNG.hash[198] ;
 wire \TRNG.hash[199] ;
 wire \TRNG.hash[19] ;
 wire \TRNG.hash[1] ;
 wire \TRNG.hash[200] ;
 wire \TRNG.hash[201] ;
 wire \TRNG.hash[202] ;
 wire \TRNG.hash[203] ;
 wire \TRNG.hash[204] ;
 wire \TRNG.hash[205] ;
 wire \TRNG.hash[206] ;
 wire \TRNG.hash[207] ;
 wire \TRNG.hash[208] ;
 wire \TRNG.hash[209] ;
 wire \TRNG.hash[20] ;
 wire \TRNG.hash[210] ;
 wire \TRNG.hash[211] ;
 wire \TRNG.hash[212] ;
 wire \TRNG.hash[213] ;
 wire \TRNG.hash[214] ;
 wire \TRNG.hash[215] ;
 wire \TRNG.hash[216] ;
 wire \TRNG.hash[217] ;
 wire \TRNG.hash[218] ;
 wire \TRNG.hash[219] ;
 wire \TRNG.hash[21] ;
 wire \TRNG.hash[220] ;
 wire \TRNG.hash[221] ;
 wire \TRNG.hash[222] ;
 wire \TRNG.hash[223] ;
 wire \TRNG.hash[224] ;
 wire \TRNG.hash[225] ;
 wire \TRNG.hash[226] ;
 wire \TRNG.hash[227] ;
 wire \TRNG.hash[228] ;
 wire \TRNG.hash[229] ;
 wire \TRNG.hash[22] ;
 wire \TRNG.hash[230] ;
 wire \TRNG.hash[231] ;
 wire \TRNG.hash[232] ;
 wire \TRNG.hash[233] ;
 wire \TRNG.hash[234] ;
 wire \TRNG.hash[235] ;
 wire \TRNG.hash[236] ;
 wire \TRNG.hash[237] ;
 wire \TRNG.hash[238] ;
 wire \TRNG.hash[239] ;
 wire \TRNG.hash[23] ;
 wire \TRNG.hash[240] ;
 wire \TRNG.hash[241] ;
 wire \TRNG.hash[242] ;
 wire \TRNG.hash[243] ;
 wire \TRNG.hash[244] ;
 wire \TRNG.hash[245] ;
 wire \TRNG.hash[246] ;
 wire \TRNG.hash[247] ;
 wire \TRNG.hash[248] ;
 wire \TRNG.hash[249] ;
 wire \TRNG.hash[24] ;
 wire \TRNG.hash[250] ;
 wire \TRNG.hash[251] ;
 wire \TRNG.hash[252] ;
 wire \TRNG.hash[253] ;
 wire \TRNG.hash[254] ;
 wire \TRNG.hash[255] ;
 wire \TRNG.hash[25] ;
 wire \TRNG.hash[26] ;
 wire \TRNG.hash[27] ;
 wire \TRNG.hash[28] ;
 wire \TRNG.hash[29] ;
 wire \TRNG.hash[2] ;
 wire \TRNG.hash[30] ;
 wire \TRNG.hash[31] ;
 wire \TRNG.hash[32] ;
 wire \TRNG.hash[33] ;
 wire \TRNG.hash[34] ;
 wire \TRNG.hash[35] ;
 wire \TRNG.hash[36] ;
 wire \TRNG.hash[37] ;
 wire \TRNG.hash[38] ;
 wire \TRNG.hash[39] ;
 wire \TRNG.hash[3] ;
 wire \TRNG.hash[40] ;
 wire \TRNG.hash[41] ;
 wire \TRNG.hash[42] ;
 wire \TRNG.hash[43] ;
 wire \TRNG.hash[44] ;
 wire \TRNG.hash[45] ;
 wire \TRNG.hash[46] ;
 wire \TRNG.hash[47] ;
 wire \TRNG.hash[48] ;
 wire \TRNG.hash[49] ;
 wire \TRNG.hash[4] ;
 wire \TRNG.hash[50] ;
 wire \TRNG.hash[51] ;
 wire \TRNG.hash[52] ;
 wire \TRNG.hash[53] ;
 wire \TRNG.hash[54] ;
 wire \TRNG.hash[55] ;
 wire \TRNG.hash[56] ;
 wire \TRNG.hash[57] ;
 wire \TRNG.hash[58] ;
 wire \TRNG.hash[59] ;
 wire \TRNG.hash[5] ;
 wire \TRNG.hash[60] ;
 wire \TRNG.hash[61] ;
 wire \TRNG.hash[62] ;
 wire \TRNG.hash[63] ;
 wire \TRNG.hash[64] ;
 wire \TRNG.hash[65] ;
 wire \TRNG.hash[66] ;
 wire \TRNG.hash[67] ;
 wire \TRNG.hash[68] ;
 wire \TRNG.hash[69] ;
 wire \TRNG.hash[6] ;
 wire \TRNG.hash[70] ;
 wire \TRNG.hash[71] ;
 wire \TRNG.hash[72] ;
 wire \TRNG.hash[73] ;
 wire \TRNG.hash[74] ;
 wire \TRNG.hash[75] ;
 wire \TRNG.hash[76] ;
 wire \TRNG.hash[77] ;
 wire \TRNG.hash[78] ;
 wire \TRNG.hash[79] ;
 wire \TRNG.hash[7] ;
 wire \TRNG.hash[80] ;
 wire \TRNG.hash[81] ;
 wire \TRNG.hash[82] ;
 wire \TRNG.hash[83] ;
 wire \TRNG.hash[84] ;
 wire \TRNG.hash[85] ;
 wire \TRNG.hash[86] ;
 wire \TRNG.hash[87] ;
 wire \TRNG.hash[88] ;
 wire \TRNG.hash[89] ;
 wire \TRNG.hash[8] ;
 wire \TRNG.hash[90] ;
 wire \TRNG.hash[91] ;
 wire \TRNG.hash[92] ;
 wire \TRNG.hash[93] ;
 wire \TRNG.hash[94] ;
 wire \TRNG.hash[95] ;
 wire \TRNG.hash[96] ;
 wire \TRNG.hash[97] ;
 wire \TRNG.hash[98] ;
 wire \TRNG.hash[99] ;
 wire \TRNG.hash[9] ;
 wire \TRNG.hash_rdy ;
 wire \TRNG.prev_ctrl_mode ;
 wire \TRNG.raw_bit_counter[0] ;
 wire \TRNG.raw_bit_counter[1] ;
 wire \TRNG.raw_bit_counter[2] ;
 wire \TRNG.raw_byte[0] ;
 wire \TRNG.raw_byte[1] ;
 wire \TRNG.raw_byte[2] ;
 wire \TRNG.raw_byte[3] ;
 wire \TRNG.raw_byte[4] ;
 wire \TRNG.raw_byte[5] ;
 wire \TRNG.raw_byte[6] ;
 wire \TRNG.raw_byte[7] ;
 wire \TRNG.sha256.K[0] ;
 wire \TRNG.sha256.K[10] ;
 wire \TRNG.sha256.K[11] ;
 wire \TRNG.sha256.K[12] ;
 wire \TRNG.sha256.K[13] ;
 wire \TRNG.sha256.K[14] ;
 wire \TRNG.sha256.K[15] ;
 wire \TRNG.sha256.K[16] ;
 wire \TRNG.sha256.K[17] ;
 wire \TRNG.sha256.K[18] ;
 wire \TRNG.sha256.K[19] ;
 wire \TRNG.sha256.K[1] ;
 wire \TRNG.sha256.K[20] ;
 wire \TRNG.sha256.K[21] ;
 wire \TRNG.sha256.K[22] ;
 wire \TRNG.sha256.K[23] ;
 wire \TRNG.sha256.K[24] ;
 wire \TRNG.sha256.K[25] ;
 wire \TRNG.sha256.K[26] ;
 wire \TRNG.sha256.K[27] ;
 wire \TRNG.sha256.K[28] ;
 wire \TRNG.sha256.K[29] ;
 wire \TRNG.sha256.K[2] ;
 wire \TRNG.sha256.K[30] ;
 wire \TRNG.sha256.K[31] ;
 wire \TRNG.sha256.K[3] ;
 wire \TRNG.sha256.K[4] ;
 wire \TRNG.sha256.K[5] ;
 wire \TRNG.sha256.K[6] ;
 wire \TRNG.sha256.K[7] ;
 wire \TRNG.sha256.K[8] ;
 wire \TRNG.sha256.K[9] ;
 wire \TRNG.sha256.W[0] ;
 wire \TRNG.sha256.W[10] ;
 wire \TRNG.sha256.W[11] ;
 wire \TRNG.sha256.W[12] ;
 wire \TRNG.sha256.W[13] ;
 wire \TRNG.sha256.W[14] ;
 wire \TRNG.sha256.W[15] ;
 wire \TRNG.sha256.W[16] ;
 wire \TRNG.sha256.W[17] ;
 wire \TRNG.sha256.W[18] ;
 wire \TRNG.sha256.W[19] ;
 wire \TRNG.sha256.W[1] ;
 wire \TRNG.sha256.W[20] ;
 wire \TRNG.sha256.W[21] ;
 wire \TRNG.sha256.W[22] ;
 wire \TRNG.sha256.W[23] ;
 wire \TRNG.sha256.W[24] ;
 wire \TRNG.sha256.W[25] ;
 wire \TRNG.sha256.W[26] ;
 wire \TRNG.sha256.W[27] ;
 wire \TRNG.sha256.W[28] ;
 wire \TRNG.sha256.W[29] ;
 wire \TRNG.sha256.W[2] ;
 wire \TRNG.sha256.W[30] ;
 wire \TRNG.sha256.W[31] ;
 wire \TRNG.sha256.W[3] ;
 wire \TRNG.sha256.W[4] ;
 wire \TRNG.sha256.W[5] ;
 wire \TRNG.sha256.W[6] ;
 wire \TRNG.sha256.W[7] ;
 wire \TRNG.sha256.W[8] ;
 wire \TRNG.sha256.W[9] ;
 wire \TRNG.sha256.compress.count[0] ;
 wire \TRNG.sha256.compress.count[1] ;
 wire \TRNG.sha256.compress.count[2] ;
 wire \TRNG.sha256.compress.count[3] ;
 wire \TRNG.sha256.compress.count[4] ;
 wire \TRNG.sha256.compress.done ;
 wire \TRNG.sha256.compress.hash_gen.temp[0] ;
 wire \TRNG.sha256.compress.hash_gen.temp[1] ;
 wire \TRNG.sha256.compress.hash_gen.temp[2] ;
 wire \TRNG.sha256.compress.hash_gen.temp[3] ;
 wire \TRNG.sha256.compress.hash_gen.temp[4] ;
 wire \TRNG.sha256.compress.hash_gen.w_rdy ;
 wire \TRNG.sha256.connect[0] ;
 wire \TRNG.sha256.connect[1] ;
 wire \TRNG.sha256.connect[2] ;
 wire \TRNG.sha256.connect[3] ;
 wire \TRNG.sha256.connect[4] ;
 wire \TRNG.sha256.connect[5] ;
 wire \TRNG.sha256.control.iteration[6] ;
 wire \TRNG.sha256.control.iteration[7] ;
 wire \TRNG.sha256.control.iteration[8] ;
 wire \TRNG.sha256.expand.address1[0] ;
 wire \TRNG.sha256.expand.address1[1] ;
 wire \TRNG.sha256.expand.address1[2] ;
 wire \TRNG.sha256.expand.address1[3] ;
 wire \TRNG.sha256.expand.address2[0] ;
 wire \TRNG.sha256.expand.address2[1] ;
 wire \TRNG.sha256.expand.address2[2] ;
 wire \TRNG.sha256.expand.address2[3] ;
 wire \TRNG.sha256.expand.data1_to_ram[0] ;
 wire \TRNG.sha256.expand.data1_to_ram[10] ;
 wire \TRNG.sha256.expand.data1_to_ram[11] ;
 wire \TRNG.sha256.expand.data1_to_ram[12] ;
 wire \TRNG.sha256.expand.data1_to_ram[13] ;
 wire \TRNG.sha256.expand.data1_to_ram[14] ;
 wire \TRNG.sha256.expand.data1_to_ram[15] ;
 wire \TRNG.sha256.expand.data1_to_ram[16] ;
 wire \TRNG.sha256.expand.data1_to_ram[17] ;
 wire \TRNG.sha256.expand.data1_to_ram[18] ;
 wire \TRNG.sha256.expand.data1_to_ram[19] ;
 wire \TRNG.sha256.expand.data1_to_ram[1] ;
 wire \TRNG.sha256.expand.data1_to_ram[20] ;
 wire \TRNG.sha256.expand.data1_to_ram[21] ;
 wire \TRNG.sha256.expand.data1_to_ram[22] ;
 wire \TRNG.sha256.expand.data1_to_ram[23] ;
 wire \TRNG.sha256.expand.data1_to_ram[24] ;
 wire \TRNG.sha256.expand.data1_to_ram[25] ;
 wire \TRNG.sha256.expand.data1_to_ram[26] ;
 wire \TRNG.sha256.expand.data1_to_ram[27] ;
 wire \TRNG.sha256.expand.data1_to_ram[28] ;
 wire \TRNG.sha256.expand.data1_to_ram[29] ;
 wire \TRNG.sha256.expand.data1_to_ram[2] ;
 wire \TRNG.sha256.expand.data1_to_ram[30] ;
 wire \TRNG.sha256.expand.data1_to_ram[31] ;
 wire \TRNG.sha256.expand.data1_to_ram[3] ;
 wire \TRNG.sha256.expand.data1_to_ram[4] ;
 wire \TRNG.sha256.expand.data1_to_ram[5] ;
 wire \TRNG.sha256.expand.data1_to_ram[6] ;
 wire \TRNG.sha256.expand.data1_to_ram[7] ;
 wire \TRNG.sha256.expand.data1_to_ram[8] ;
 wire \TRNG.sha256.expand.data1_to_ram[9] ;
 wire \TRNG.sha256.expand.dout1[0] ;
 wire \TRNG.sha256.expand.dout1[10] ;
 wire \TRNG.sha256.expand.dout1[11] ;
 wire \TRNG.sha256.expand.dout1[12] ;
 wire \TRNG.sha256.expand.dout1[13] ;
 wire \TRNG.sha256.expand.dout1[14] ;
 wire \TRNG.sha256.expand.dout1[15] ;
 wire \TRNG.sha256.expand.dout1[16] ;
 wire \TRNG.sha256.expand.dout1[17] ;
 wire \TRNG.sha256.expand.dout1[18] ;
 wire \TRNG.sha256.expand.dout1[19] ;
 wire \TRNG.sha256.expand.dout1[1] ;
 wire \TRNG.sha256.expand.dout1[20] ;
 wire \TRNG.sha256.expand.dout1[21] ;
 wire \TRNG.sha256.expand.dout1[22] ;
 wire \TRNG.sha256.expand.dout1[23] ;
 wire \TRNG.sha256.expand.dout1[24] ;
 wire \TRNG.sha256.expand.dout1[25] ;
 wire \TRNG.sha256.expand.dout1[26] ;
 wire \TRNG.sha256.expand.dout1[27] ;
 wire \TRNG.sha256.expand.dout1[28] ;
 wire \TRNG.sha256.expand.dout1[29] ;
 wire \TRNG.sha256.expand.dout1[2] ;
 wire \TRNG.sha256.expand.dout1[30] ;
 wire \TRNG.sha256.expand.dout1[31] ;
 wire \TRNG.sha256.expand.dout1[3] ;
 wire \TRNG.sha256.expand.dout1[4] ;
 wire \TRNG.sha256.expand.dout1[5] ;
 wire \TRNG.sha256.expand.dout1[6] ;
 wire \TRNG.sha256.expand.dout1[7] ;
 wire \TRNG.sha256.expand.dout1[8] ;
 wire \TRNG.sha256.expand.dout1[9] ;
 wire \TRNG.sha256.expand.dout2[0] ;
 wire \TRNG.sha256.expand.dout2[10] ;
 wire \TRNG.sha256.expand.dout2[11] ;
 wire \TRNG.sha256.expand.dout2[12] ;
 wire \TRNG.sha256.expand.dout2[13] ;
 wire \TRNG.sha256.expand.dout2[14] ;
 wire \TRNG.sha256.expand.dout2[15] ;
 wire \TRNG.sha256.expand.dout2[16] ;
 wire \TRNG.sha256.expand.dout2[17] ;
 wire \TRNG.sha256.expand.dout2[18] ;
 wire \TRNG.sha256.expand.dout2[19] ;
 wire \TRNG.sha256.expand.dout2[1] ;
 wire \TRNG.sha256.expand.dout2[20] ;
 wire \TRNG.sha256.expand.dout2[21] ;
 wire \TRNG.sha256.expand.dout2[22] ;
 wire \TRNG.sha256.expand.dout2[23] ;
 wire \TRNG.sha256.expand.dout2[24] ;
 wire \TRNG.sha256.expand.dout2[25] ;
 wire \TRNG.sha256.expand.dout2[26] ;
 wire \TRNG.sha256.expand.dout2[27] ;
 wire \TRNG.sha256.expand.dout2[28] ;
 wire \TRNG.sha256.expand.dout2[29] ;
 wire \TRNG.sha256.expand.dout2[2] ;
 wire \TRNG.sha256.expand.dout2[30] ;
 wire \TRNG.sha256.expand.dout2[31] ;
 wire \TRNG.sha256.expand.dout2[3] ;
 wire \TRNG.sha256.expand.dout2[4] ;
 wire \TRNG.sha256.expand.dout2[5] ;
 wire \TRNG.sha256.expand.dout2[6] ;
 wire \TRNG.sha256.expand.dout2[7] ;
 wire \TRNG.sha256.expand.dout2[8] ;
 wire \TRNG.sha256.expand.dout2[9] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[0] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[10] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[11] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[12] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[13] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[14] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[15] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[16] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[17] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[18] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[19] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[1] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[20] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[21] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[22] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[23] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[24] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[25] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[26] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[27] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[28] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[29] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[2] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[30] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[31] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[3] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[4] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[5] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[6] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[7] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[8] ;
 wire \TRNG.sha256.expand.exp_ctrl.final_sum[9] ;
 wire \TRNG.sha256.expand.exp_ctrl.j[0] ;
 wire \TRNG.sha256.expand.exp_ctrl.j[1] ;
 wire \TRNG.sha256.expand.exp_ctrl.j[2] ;
 wire \TRNG.sha256.expand.exp_ctrl.j[3] ;
 wire \TRNG.sha256.expand.exp_ctrl.j_15[0] ;
 wire \TRNG.sha256.expand.exp_ctrl.j_15[1] ;
 wire \TRNG.sha256.expand.exp_ctrl.j_15[2] ;
 wire \TRNG.sha256.expand.exp_ctrl.j_15[3] ;
 wire \TRNG.sha256.expand.exp_ctrl.j_2[0] ;
 wire \TRNG.sha256.expand.exp_ctrl.j_2[1] ;
 wire \TRNG.sha256.expand.exp_ctrl.j_2[2] ;
 wire \TRNG.sha256.expand.exp_ctrl.j_2[3] ;
 wire \TRNG.sha256.expand.exp_ctrl.j_7[0] ;
 wire \TRNG.sha256.expand.exp_ctrl.j_7[1] ;
 wire \TRNG.sha256.expand.exp_ctrl.j_7[2] ;
 wire \TRNG.sha256.expand.exp_ctrl.j_7[3] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[0] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[10] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[11] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[12] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[13] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[14] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[15] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[16] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[17] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[18] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[19] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[1] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[20] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[21] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[22] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[23] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[24] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[25] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[26] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[27] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[28] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[29] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[2] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[30] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[31] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[3] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[4] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[5] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[6] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[7] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[8] ;
 wire \TRNG.sha256.expand.exp_ctrl.sum[9] ;
 wire \TRNG.sha256.expand.exp_ctrl.write_en1 ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][0] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][10] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][11] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][12] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][13] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][14] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][15] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][16] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][17] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][18] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][19] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][1] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][20] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][21] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][22] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][23] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][24] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][25] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][26] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][27] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][28] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][29] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][2] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][30] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][31] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][3] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][4] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][5] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][6] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][7] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][8] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[0][9] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][0] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][10] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][11] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][12] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][13] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][14] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][15] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][16] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][17] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][18] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][19] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][1] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][20] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][21] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][22] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][23] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][24] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][25] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][26] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][27] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][28] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][29] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][2] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][30] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][31] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][3] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][4] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][5] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][6] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][7] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][8] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[10][9] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][0] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][10] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][11] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][12] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][13] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][14] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][15] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][16] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][17] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][18] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][19] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][1] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][20] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][21] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][22] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][23] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][24] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][25] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][26] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][27] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][28] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][29] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][2] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][30] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][31] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][3] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][4] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][5] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][6] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][7] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][8] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[11][9] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][0] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][10] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][11] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][12] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][13] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][14] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][15] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][16] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][17] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][18] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][19] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][1] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][20] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][21] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][22] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][23] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][24] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][25] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][26] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][27] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][28] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][29] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][2] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][30] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][31] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][3] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][4] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][5] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][6] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][7] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][8] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[12][9] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][0] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][10] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][11] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][12] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][13] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][14] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][15] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][16] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][17] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][18] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][19] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][1] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][20] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][21] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][22] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][23] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][24] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][25] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][26] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][27] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][28] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][29] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][2] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][30] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][31] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][3] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][4] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][5] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][6] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][7] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][8] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[13][9] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][0] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][10] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][11] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][12] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][13] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][14] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][15] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][16] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][17] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][18] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][19] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][1] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][20] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][21] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][22] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][23] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][24] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][25] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][26] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][27] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][28] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][29] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][2] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][30] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][31] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][3] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][4] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][5] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][6] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][7] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][8] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[14][9] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][0] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][10] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][11] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][12] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][13] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][14] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][15] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][16] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][17] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][18] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][19] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][1] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][20] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][21] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][22] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][23] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][24] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][25] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][26] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][27] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][28] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][29] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][2] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][30] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][31] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][3] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][4] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][5] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][6] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][7] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][8] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[15][9] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][0] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][10] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][11] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][12] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][13] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][14] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][15] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][16] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][17] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][18] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][19] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][1] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][20] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][21] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][22] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][23] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][24] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][25] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][26] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][27] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][28] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][29] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][2] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][30] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][31] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][3] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][4] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][5] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][6] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][7] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][8] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[1][9] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][0] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][10] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][11] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][12] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][13] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][14] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][15] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][16] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][17] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][18] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][19] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][1] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][20] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][21] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][22] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][23] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][24] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][25] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][26] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][27] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][28] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][29] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][2] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][30] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][31] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][3] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][4] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][5] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][6] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][7] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][8] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[2][9] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][0] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][10] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][11] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][12] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][13] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][14] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][15] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][16] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][17] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][18] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][19] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][1] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][20] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][21] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][22] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][23] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][24] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][25] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][26] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][27] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][28] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][29] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][2] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][30] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][31] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][3] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][4] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][5] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][6] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][7] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][8] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[3][9] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][0] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][10] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][11] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][12] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][13] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][14] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][15] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][16] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][17] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][18] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][19] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][1] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][20] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][21] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][22] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][23] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][24] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][25] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][26] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][27] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][28] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][29] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][2] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][30] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][31] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][3] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][4] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][5] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][6] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][7] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][8] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[4][9] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][0] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][10] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][11] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][12] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][13] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][14] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][15] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][16] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][17] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][18] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][19] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][1] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][20] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][21] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][22] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][23] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][24] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][25] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][26] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][27] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][28] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][29] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][2] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][30] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][31] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][3] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][4] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][5] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][6] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][7] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][8] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[5][9] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][0] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][10] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][11] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][12] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][13] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][14] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][15] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][16] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][17] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][18] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][19] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][1] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][20] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][21] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][22] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][23] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][24] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][25] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][26] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][27] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][28] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][29] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][2] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][30] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][31] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][3] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][4] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][5] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][6] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][7] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][8] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[6][9] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][0] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][10] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][11] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][12] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][13] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][14] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][15] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][16] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][17] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][18] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][19] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][1] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][20] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][21] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][22] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][23] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][24] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][25] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][26] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][27] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][28] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][29] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][2] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][30] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][31] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][3] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][4] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][5] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][6] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][7] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][8] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[7][9] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][0] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][10] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][11] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][12] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][13] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][14] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][15] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][16] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][17] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][18] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][19] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][1] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][20] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][21] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][22] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][23] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][24] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][25] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][26] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][27] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][28] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][29] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][2] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][30] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][31] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][3] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][4] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][5] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][6] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][7] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][8] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[8][9] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][0] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][10] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][11] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][12] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][13] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][14] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][15] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][16] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][17] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][18] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][19] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][1] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][20] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][21] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][22] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][23] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][24] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][25] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][26] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][27] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][28] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][29] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][2] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][30] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][31] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][3] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][4] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][5] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][6] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][7] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][8] ;
 wire \TRNG.sha256.expand.msg_schdl.RAM[9][9] ;
 wire \TRNG.sha256.expand.sm0.sum_0[0] ;
 wire \TRNG.sha256.expand.sm0.sum_0[10] ;
 wire \TRNG.sha256.expand.sm0.sum_0[11] ;
 wire \TRNG.sha256.expand.sm0.sum_0[12] ;
 wire \TRNG.sha256.expand.sm0.sum_0[13] ;
 wire \TRNG.sha256.expand.sm0.sum_0[14] ;
 wire \TRNG.sha256.expand.sm0.sum_0[15] ;
 wire \TRNG.sha256.expand.sm0.sum_0[16] ;
 wire \TRNG.sha256.expand.sm0.sum_0[17] ;
 wire \TRNG.sha256.expand.sm0.sum_0[18] ;
 wire \TRNG.sha256.expand.sm0.sum_0[19] ;
 wire \TRNG.sha256.expand.sm0.sum_0[1] ;
 wire \TRNG.sha256.expand.sm0.sum_0[20] ;
 wire \TRNG.sha256.expand.sm0.sum_0[21] ;
 wire \TRNG.sha256.expand.sm0.sum_0[22] ;
 wire \TRNG.sha256.expand.sm0.sum_0[23] ;
 wire \TRNG.sha256.expand.sm0.sum_0[24] ;
 wire \TRNG.sha256.expand.sm0.sum_0[25] ;
 wire \TRNG.sha256.expand.sm0.sum_0[26] ;
 wire \TRNG.sha256.expand.sm0.sum_0[27] ;
 wire \TRNG.sha256.expand.sm0.sum_0[28] ;
 wire \TRNG.sha256.expand.sm0.sum_0[29] ;
 wire \TRNG.sha256.expand.sm0.sum_0[2] ;
 wire \TRNG.sha256.expand.sm0.sum_0[30] ;
 wire \TRNG.sha256.expand.sm0.sum_0[31] ;
 wire \TRNG.sha256.expand.sm0.sum_0[3] ;
 wire \TRNG.sha256.expand.sm0.sum_0[4] ;
 wire \TRNG.sha256.expand.sm0.sum_0[5] ;
 wire \TRNG.sha256.expand.sm0.sum_0[6] ;
 wire \TRNG.sha256.expand.sm0.sum_0[7] ;
 wire \TRNG.sha256.expand.sm0.sum_0[8] ;
 wire \TRNG.sha256.expand.sm0.sum_0[9] ;
 wire \TRNG.state[0] ;
 wire \TRNG.state[1] ;
 wire \TRNG.state[2] ;
 wire \TRNG.uart_start ;
 wire \TRNG.uart_tx_inst.currentState[0] ;
 wire \TRNG.uart_tx_inst.currentState[1] ;
 wire \TRNG.uart_tx_inst.currentState[2] ;
 wire \TRNG.uart_tx_inst.currentState[3] ;
 wire \TRNG.uart_tx_inst.currentState[4] ;
 wire \TRNG.uart_tx_inst.ticks_counter[0] ;
 wire \TRNG.uart_tx_inst.ticks_counter[1] ;
 wire \TRNG.uart_tx_inst.ticks_counter[2] ;
 wire \TRNG.uart_tx_inst.ticks_counter[3] ;
 wire \TRNG.uart_tx_inst.ticks_counter[4] ;
 wire \TRNG.uart_tx_inst.ticks_counter[5] ;
 wire \TRNG.uart_tx_inst.ticks_counter[6] ;
 wire \TRNG.uart_tx_inst.ticks_counter[7] ;
 wire \TRNG.uart_tx_inst.ticks_counter[8] ;
 wire \TRNG.uart_tx_inst.tx_bit_counter[0] ;
 wire \TRNG.uart_tx_inst.tx_bit_counter[1] ;
 wire \TRNG.uart_tx_inst.tx_bit_counter[2] ;
 wire \TRNG.uart_tx_inst.tx_bit_counter[3] ;
 wire \TRNG.uart_tx_inst.tx_reg[0] ;
 wire \TRNG.uart_tx_inst.tx_reg[1] ;
 wire \TRNG.uart_tx_inst.tx_reg[2] ;
 wire \TRNG.uart_tx_inst.tx_reg[3] ;
 wire \TRNG.uart_tx_inst.tx_reg[4] ;
 wire \TRNG.uart_tx_inst.tx_reg[5] ;
 wire \TRNG.uart_tx_inst.tx_reg[6] ;
 wire \TRNG.uart_tx_inst.tx_reg[7] ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire clknet_leaf_0_clk;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net4570;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4625;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net4630;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4644;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net4997;
 wire net4998;
 wire net4999;
 wire net5000;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net5010;
 wire net5011;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5023;
 wire net5024;
 wire net5025;
 wire net5026;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5035;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5227;
 wire net5228;
 wire net5229;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net5260;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5278;
 wire net5279;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5346;
 wire net5347;
 wire net5348;
 wire net5349;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net5360;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net5386;
 wire net5387;
 wire net5388;
 wire net5389;
 wire net5390;
 wire net5391;
 wire net5392;
 wire net5393;
 wire net5394;
 wire net5395;
 wire net5396;
 wire net5397;
 wire net5398;
 wire net5399;
 wire net5400;
 wire net5401;
 wire net5402;
 wire net5403;
 wire net5404;
 wire net5405;
 wire net5406;
 wire net5407;
 wire net5408;
 wire net5409;
 wire net5410;
 wire net5411;
 wire net5412;
 wire net5413;
 wire net5414;
 wire net5415;
 wire net5416;
 wire net5417;
 wire net5418;
 wire net5419;
 wire net5420;
 wire net5421;
 wire net5422;
 wire net5423;
 wire net5424;
 wire net5425;
 wire net5426;
 wire net5427;
 wire net5428;
 wire net5429;
 wire net5430;
 wire net5431;
 wire net5432;
 wire net5433;
 wire net5434;
 wire net5435;
 wire net5436;
 wire net5437;
 wire net5438;
 wire net5439;
 wire net5440;
 wire net5441;
 wire net5442;
 wire net5443;
 wire net5444;
 wire net5445;
 wire net5446;
 wire net5447;
 wire net5448;
 wire net5449;
 wire net5450;
 wire net5451;
 wire net5452;
 wire net5453;
 wire net5454;
 wire net5455;
 wire net5456;
 wire net5457;
 wire net5458;
 wire net5459;
 wire net5460;
 wire net5461;
 wire net5462;
 wire net5463;
 wire net5464;
 wire net5465;
 wire net5466;
 wire net5467;
 wire net5468;
 wire net5469;
 wire net5470;
 wire net5471;
 wire net5472;
 wire net5473;
 wire net5474;
 wire net5475;
 wire net5476;
 wire net5477;
 wire net5478;
 wire net5479;
 wire net5480;
 wire net5481;
 wire net5482;
 wire net5483;
 wire net5484;
 wire net5485;
 wire net5486;
 wire net5487;
 wire net5488;
 wire net5489;
 wire net5490;
 wire net5491;
 wire net5492;
 wire net5493;
 wire net5494;
 wire net5495;
 wire net5496;
 wire net5497;
 wire net5498;
 wire net5499;
 wire net5500;
 wire net5501;
 wire net5502;
 wire net5503;
 wire net5504;
 wire net5505;
 wire net5506;
 wire net5507;
 wire net5508;
 wire net5509;
 wire net5510;
 wire net5511;
 wire net5512;
 wire net5513;
 wire net5514;
 wire net5515;
 wire net5516;
 wire net5517;
 wire net5518;
 wire net5519;
 wire net5520;
 wire net5521;
 wire net5522;
 wire net5523;
 wire net5524;
 wire net5525;
 wire net5526;
 wire net5527;
 wire net5528;
 wire net5529;
 wire net5530;
 wire net5531;
 wire net5532;
 wire net5533;
 wire net5534;
 wire net5535;
 wire net5536;
 wire net5537;
 wire net5538;
 wire net5539;
 wire net5540;
 wire net5541;
 wire net5542;
 wire net5543;
 wire net5544;
 wire net5545;
 wire net5546;
 wire net5547;
 wire net5548;
 wire net5549;
 wire net5550;
 wire net5551;
 wire net5552;
 wire net5553;
 wire net5554;
 wire net5555;
 wire net5556;
 wire net5557;
 wire net5558;
 wire net5559;
 wire net5560;
 wire net5561;
 wire net5562;
 wire net5563;
 wire net5564;
 wire net5565;
 wire net5566;
 wire net5567;
 wire net5568;
 wire net5569;
 wire net5570;
 wire net5571;
 wire net5572;
 wire net5573;
 wire net5574;
 wire net5575;
 wire net5576;
 wire net5577;
 wire net5578;
 wire net5579;
 wire net5580;
 wire net5581;
 wire net5582;
 wire net5583;
 wire net5584;
 wire net5585;
 wire net5586;
 wire net5587;
 wire net5588;
 wire net5589;
 wire net5590;
 wire net5591;
 wire net5592;
 wire net5593;
 wire net5594;
 wire net5595;
 wire net5596;
 wire net5597;
 wire net5598;
 wire net5599;
 wire net5600;
 wire net5601;
 wire net5602;
 wire net5603;
 wire net5604;
 wire net5605;
 wire net5606;
 wire net5607;
 wire net5608;
 wire net5609;
 wire net5610;
 wire net5611;
 wire net5612;
 wire net5613;
 wire net5614;
 wire net5615;
 wire net5616;
 wire net5617;
 wire net5618;
 wire net5619;
 wire net5620;
 wire net5621;
 wire net5622;
 wire net5623;
 wire net5624;
 wire net5625;
 wire net5626;
 wire net5627;
 wire net5628;
 wire net5629;
 wire net5630;
 wire net5631;
 wire net5632;
 wire net5633;
 wire net5634;
 wire net5635;
 wire net5636;
 wire net5637;
 wire net5638;
 wire net5639;
 wire net5640;
 wire net5641;
 wire net5642;
 wire net5643;
 wire net5644;
 wire net5645;
 wire net5646;
 wire net5647;
 wire net5648;
 wire net5649;
 wire net5650;
 wire net5651;
 wire net5652;
 wire net5653;
 wire net5654;
 wire net5655;
 wire net5656;
 wire net5657;
 wire net5658;
 wire net5659;
 wire net5660;
 wire net5661;
 wire net5662;
 wire net5663;
 wire net5664;
 wire net5665;
 wire net5666;
 wire net5667;
 wire net5668;
 wire net5669;
 wire net5670;
 wire net5671;
 wire net5672;
 wire net5673;
 wire net5674;
 wire net5675;
 wire net5676;
 wire net5677;
 wire net5678;
 wire net5679;
 wire net5680;
 wire net5681;
 wire net5682;
 wire net5683;
 wire net5684;
 wire net5685;
 wire net5686;
 wire net5687;
 wire net5688;
 wire net5689;
 wire net5690;
 wire net5691;
 wire net5692;
 wire net5693;
 wire net5694;
 wire net5695;
 wire net5696;
 wire net5697;
 wire net5698;
 wire net5699;
 wire net5700;
 wire net5701;
 wire net5702;
 wire net5703;
 wire net5704;
 wire net5705;
 wire net5706;
 wire net5707;
 wire net5708;
 wire net5709;
 wire net5710;
 wire net5711;
 wire net5712;
 wire net5713;
 wire net5714;
 wire net5715;
 wire net5716;
 wire net5717;
 wire net5718;
 wire net5719;
 wire net5720;
 wire net5721;
 wire net5722;
 wire net5723;
 wire net5724;
 wire net5725;
 wire net5726;
 wire net5727;
 wire net5728;
 wire net5729;
 wire net5730;
 wire net5731;
 wire net5732;
 wire net5733;
 wire net5734;
 wire net5735;
 wire net5736;
 wire net5737;
 wire net5738;
 wire net5739;
 wire net5740;
 wire net5741;
 wire net5742;
 wire net5743;
 wire net5744;
 wire net5745;
 wire net5746;
 wire net5747;
 wire net5748;
 wire net5749;
 wire net5750;
 wire net5751;
 wire net5752;
 wire net5753;
 wire net5754;
 wire net5755;
 wire net5756;
 wire net5757;
 wire net5758;
 wire net5759;
 wire net5760;
 wire net5761;
 wire net5762;
 wire net5763;
 wire net5764;
 wire net5765;
 wire net5766;
 wire net5767;
 wire net5768;
 wire net5769;
 wire net5770;
 wire net5771;
 wire net5772;
 wire net5773;
 wire net5774;
 wire net5775;
 wire net5776;
 wire net5777;
 wire net5778;
 wire net5779;
 wire net5780;
 wire net5781;
 wire net5782;
 wire net5783;
 wire net5784;
 wire net5785;
 wire net5786;
 wire net5787;
 wire net5788;
 wire net5789;
 wire net5790;
 wire net5791;
 wire net5792;
 wire net5793;
 wire net5794;
 wire net5795;
 wire net5796;
 wire net5797;
 wire net5798;
 wire net5799;
 wire net5800;
 wire net5801;
 wire net5802;
 wire net5803;
 wire net5804;
 wire net5805;
 wire net5806;
 wire net5807;
 wire net5808;
 wire net5809;
 wire net5810;
 wire net5811;
 wire net5812;
 wire net5813;
 wire net5814;
 wire net5815;
 wire net5816;
 wire net5817;
 wire net5818;
 wire net5819;
 wire net5820;
 wire net5821;
 wire net5822;
 wire net5823;
 wire net5824;
 wire net5825;
 wire net5826;
 wire net5827;
 wire net5828;
 wire net5829;
 wire net5830;
 wire net5831;
 wire net5832;
 wire net5833;
 wire net5834;
 wire net5835;
 wire net5836;
 wire net5837;
 wire net5838;
 wire net5839;
 wire net5840;
 wire net5841;
 wire net5842;
 wire net5843;
 wire net5844;
 wire net5845;
 wire net5846;
 wire net5847;
 wire net5848;
 wire net5849;
 wire net5850;
 wire net5851;
 wire net5852;
 wire net5853;
 wire net5854;
 wire net5855;
 wire net5856;
 wire net5857;
 wire net5858;
 wire net5859;
 wire net5860;
 wire net5861;
 wire net5862;
 wire net5863;
 wire net5864;
 wire net5865;
 wire net5866;
 wire net5867;
 wire net5868;
 wire net5869;
 wire net5870;
 wire net5871;
 wire net5872;
 wire net5873;
 wire net5874;
 wire net5875;
 wire net5876;
 wire net5877;
 wire net5878;
 wire net5879;
 wire net5880;
 wire net5881;
 wire net5882;
 wire net5883;
 wire net5884;
 wire net5885;
 wire net5886;
 wire net5887;
 wire net5888;
 wire net5889;
 wire net5890;
 wire net5891;
 wire net5892;
 wire net5893;
 wire net5894;
 wire net5895;
 wire net5896;
 wire net5897;
 wire net5898;
 wire net5899;
 wire net5900;
 wire net5901;
 wire net5902;
 wire net5903;
 wire net5904;
 wire net5905;
 wire net5906;
 wire net5907;
 wire net5908;
 wire net5909;
 wire net5910;
 wire net5911;
 wire net5912;
 wire net5913;
 wire net5914;
 wire net5915;
 wire net5916;
 wire net5917;
 wire net5918;
 wire net5919;
 wire net5920;
 wire net5921;
 wire net5922;
 wire net5923;
 wire net5924;
 wire net5925;
 wire net5926;
 wire net5927;
 wire net5928;
 wire net5929;
 wire net5930;
 wire net5931;
 wire net5932;
 wire net5933;
 wire net5934;
 wire net5935;
 wire net5936;
 wire net5937;
 wire net5938;
 wire net5939;
 wire net5940;
 wire net5941;
 wire net5942;
 wire net5943;
 wire net5944;
 wire net5945;
 wire net5946;
 wire net5947;
 wire net5948;
 wire net5949;
 wire net5950;
 wire net5951;
 wire net5952;
 wire net5953;
 wire net5954;
 wire net5955;
 wire net5956;
 wire net5957;
 wire net5958;
 wire net5959;
 wire net5960;
 wire net5961;
 wire net5962;
 wire net5963;
 wire net5964;
 wire net5965;
 wire net5966;
 wire net5967;
 wire net5968;
 wire net5969;
 wire net5970;
 wire net5971;
 wire net5972;
 wire net5973;
 wire net5974;
 wire net5975;
 wire net5976;
 wire net5977;
 wire net5978;
 wire net5979;
 wire net5980;
 wire net5981;
 wire net5982;
 wire net5983;
 wire net5984;
 wire net5985;
 wire net5986;
 wire net5987;
 wire net5988;
 wire net5989;
 wire net5990;
 wire net5991;
 wire net5992;
 wire net5993;
 wire net5994;
 wire net5995;
 wire net5996;
 wire net5997;
 wire net5998;
 wire net5999;
 wire net6000;
 wire net6001;
 wire net6002;
 wire net6003;
 wire net6004;
 wire net6005;
 wire net6006;
 wire net6007;
 wire net6008;
 wire net6009;
 wire net6010;
 wire net6011;
 wire net6012;
 wire net6013;
 wire net6014;
 wire net6015;
 wire net6016;
 wire net6017;
 wire net6018;
 wire net6019;
 wire net6020;
 wire net6021;
 wire net6022;
 wire net6023;
 wire net6024;
 wire net6025;
 wire net6026;
 wire net6027;
 wire net6028;
 wire net6029;
 wire net6030;
 wire net6031;
 wire net6032;
 wire net6033;
 wire net6034;
 wire net6035;
 wire net6036;
 wire net6037;
 wire net6038;
 wire net6039;
 wire net6040;
 wire net6041;
 wire net6042;
 wire net6043;
 wire net6044;
 wire net6045;
 wire net6046;
 wire net6047;
 wire net6048;
 wire net6049;
 wire net6050;
 wire net6051;
 wire net6052;
 wire net6053;
 wire net6054;
 wire net6055;
 wire net6056;
 wire net6057;
 wire net6058;
 wire net6059;
 wire net6060;
 wire net6061;
 wire net6062;
 wire net6063;
 wire net6064;
 wire net6065;
 wire net6066;
 wire net1;
 wire net2;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0_0_clk;
 wire clknet_6_1_0_clk;
 wire clknet_6_2_0_clk;
 wire clknet_6_3_0_clk;
 wire clknet_6_4_0_clk;
 wire clknet_6_5_0_clk;
 wire clknet_6_6_0_clk;
 wire clknet_6_7_0_clk;
 wire clknet_6_8_0_clk;
 wire clknet_6_9_0_clk;
 wire clknet_6_10_0_clk;
 wire clknet_6_11_0_clk;
 wire clknet_6_12_0_clk;
 wire clknet_6_13_0_clk;
 wire clknet_6_14_0_clk;
 wire clknet_6_15_0_clk;
 wire clknet_6_16_0_clk;
 wire clknet_6_17_0_clk;
 wire clknet_6_18_0_clk;
 wire clknet_6_19_0_clk;
 wire clknet_6_20_0_clk;
 wire clknet_6_21_0_clk;
 wire clknet_6_22_0_clk;
 wire clknet_6_23_0_clk;
 wire clknet_6_24_0_clk;
 wire clknet_6_25_0_clk;
 wire clknet_6_26_0_clk;
 wire clknet_6_27_0_clk;
 wire clknet_6_28_0_clk;
 wire clknet_6_29_0_clk;
 wire clknet_6_30_0_clk;
 wire clknet_6_31_0_clk;
 wire clknet_6_32_0_clk;
 wire clknet_6_33_0_clk;
 wire clknet_6_34_0_clk;
 wire clknet_6_35_0_clk;
 wire clknet_6_36_0_clk;
 wire clknet_6_37_0_clk;
 wire clknet_6_38_0_clk;
 wire clknet_6_39_0_clk;
 wire clknet_6_40_0_clk;
 wire clknet_6_41_0_clk;
 wire clknet_6_42_0_clk;
 wire clknet_6_43_0_clk;
 wire clknet_6_44_0_clk;
 wire clknet_6_45_0_clk;
 wire clknet_6_46_0_clk;
 wire clknet_6_47_0_clk;
 wire clknet_6_48_0_clk;
 wire clknet_6_49_0_clk;
 wire clknet_6_50_0_clk;
 wire clknet_6_51_0_clk;
 wire clknet_6_52_0_clk;
 wire clknet_6_53_0_clk;
 wire clknet_6_54_0_clk;
 wire clknet_6_55_0_clk;
 wire clknet_6_56_0_clk;
 wire clknet_6_57_0_clk;
 wire clknet_6_58_0_clk;
 wire clknet_6_59_0_clk;
 wire clknet_6_60_0_clk;
 wire clknet_6_61_0_clk;
 wire clknet_6_62_0_clk;
 wire clknet_6_63_0_clk;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;

 sg13g2_inv_1 _12194_ (.Y(_04220_),
    .A(\TRNG.hash[71] ));
 sg13g2_inv_1 _12195_ (.Y(_04221_),
    .A(\TRNG.hash[126] ));
 sg13g2_inv_1 _12196_ (.Y(_04222_),
    .A(\TRNG.hash[105] ));
 sg13g2_inv_1 _12197_ (.Y(_04223_),
    .A(net3784));
 sg13g2_inv_1 _12198_ (.Y(_04224_),
    .A(\TRNG.hash[213] ));
 sg13g2_inv_1 _12199_ (.Y(_04225_),
    .A(net3513));
 sg13g2_inv_1 _12200_ (.Y(_04226_),
    .A(\TRNG.hash[240] ));
 sg13g2_inv_1 _12201_ (.Y(_04227_),
    .A(net2873));
 sg13g2_inv_8 _12202_ (.Y(_04228_),
    .A(net5572));
 sg13g2_inv_1 _12203_ (.Y(_04229_),
    .A(net3655));
 sg13g2_inv_2 _12204_ (.Y(_04230_),
    .A(net3534));
 sg13g2_inv_2 _12205_ (.Y(_04231_),
    .A(net3675));
 sg13g2_inv_1 _12206_ (.Y(_04232_),
    .A(net3842));
 sg13g2_inv_1 _12207_ (.Y(_04233_),
    .A(net3465));
 sg13g2_inv_1 _12208_ (.Y(_04234_),
    .A(net3852));
 sg13g2_inv_1 _12209_ (.Y(_04235_),
    .A(net5576));
 sg13g2_inv_1 _12210_ (.Y(_04236_),
    .A(net5581));
 sg13g2_inv_1 _12211_ (.Y(_04237_),
    .A(net5600));
 sg13g2_inv_1 _12212_ (.Y(_04238_),
    .A(net5610));
 sg13g2_inv_2 _12213_ (.Y(_04239_),
    .A(net5614));
 sg13g2_inv_1 _12214_ (.Y(_04240_),
    .A(net2478));
 sg13g2_inv_1 _12215_ (.Y(_04241_),
    .A(net2512));
 sg13g2_inv_1 _12216_ (.Y(_04242_),
    .A(net1931));
 sg13g2_inv_1 _12217_ (.Y(_04243_),
    .A(net2271));
 sg13g2_inv_1 _12218_ (.Y(_04244_),
    .A(net2134));
 sg13g2_inv_1 _12219_ (.Y(_04245_),
    .A(net2458));
 sg13g2_inv_1 _12220_ (.Y(_04246_),
    .A(net2623));
 sg13g2_inv_1 _12221_ (.Y(_04247_),
    .A(net2305));
 sg13g2_inv_1 _12222_ (.Y(_04248_),
    .A(net2344));
 sg13g2_inv_1 _12223_ (.Y(_04249_),
    .A(net1853));
 sg13g2_inv_1 _12224_ (.Y(_04250_),
    .A(net2661));
 sg13g2_inv_1 _12225_ (.Y(_04251_),
    .A(net1886));
 sg13g2_inv_1 _12226_ (.Y(_04252_),
    .A(net2394));
 sg13g2_inv_1 _12227_ (.Y(_04253_),
    .A(net2269));
 sg13g2_inv_1 _12228_ (.Y(_04254_),
    .A(net2634));
 sg13g2_inv_1 _12229_ (.Y(_04255_),
    .A(net2392));
 sg13g2_inv_1 _12230_ (.Y(_04256_),
    .A(net2476));
 sg13g2_inv_1 _12231_ (.Y(_04257_),
    .A(net2467));
 sg13g2_inv_1 _12232_ (.Y(_04258_),
    .A(net2229));
 sg13g2_inv_1 _12233_ (.Y(_04259_),
    .A(net2342));
 sg13g2_inv_1 _12234_ (.Y(_04260_),
    .A(net2536));
 sg13g2_inv_1 _12235_ (.Y(_04261_),
    .A(net2443));
 sg13g2_inv_1 _12236_ (.Y(_04262_),
    .A(net2209));
 sg13g2_inv_1 _12237_ (.Y(_04263_),
    .A(net2415));
 sg13g2_inv_1 _12238_ (.Y(_04264_),
    .A(net2226));
 sg13g2_inv_1 _12239_ (.Y(_04265_),
    .A(net2299));
 sg13g2_inv_1 _12240_ (.Y(_04266_),
    .A(net2038));
 sg13g2_inv_1 _12241_ (.Y(_04267_),
    .A(net2307));
 sg13g2_inv_1 _12242_ (.Y(_04268_),
    .A(net2403));
 sg13g2_inv_1 _12243_ (.Y(_04269_),
    .A(net2265));
 sg13g2_inv_1 _12244_ (.Y(_04270_),
    .A(net2352));
 sg13g2_inv_1 _12245_ (.Y(_04271_),
    .A(net2541));
 sg13g2_inv_1 _12246_ (.Y(_04272_),
    .A(\TRNG.sha256.expand.exp_ctrl.j_15[0] ));
 sg13g2_inv_1 _12247_ (.Y(_04273_),
    .A(\TRNG.sha256.expand.exp_ctrl.j_7[0] ));
 sg13g2_inv_1 _12248_ (.Y(_04274_),
    .A(net1180));
 sg13g2_inv_1 _12249_ (.Y(_04275_),
    .A(net1136));
 sg13g2_inv_2 _12250_ (.Y(_04276_),
    .A(net3232));
 sg13g2_inv_1 _12251_ (.Y(_04277_),
    .A(\TRNG.sha256.expand.address1[3] ));
 sg13g2_inv_1 _12252_ (.Y(_04278_),
    .A(\TRNG.sha256.expand.address1[2] ));
 sg13g2_inv_2 _12253_ (.Y(_04279_),
    .A(net5857));
 sg13g2_inv_1 _12254_ (.Y(_04280_),
    .A(\TRNG.hash[250] ));
 sg13g2_inv_1 _12255_ (.Y(_04281_),
    .A(\TRNG.hash[246] ));
 sg13g2_inv_1 _12256_ (.Y(_04282_),
    .A(net5881));
 sg13g2_inv_1 _12257_ (.Y(_04283_),
    .A(\TRNG.hash[235] ));
 sg13g2_inv_1 _12258_ (.Y(_04284_),
    .A(\TRNG.hash[231] ));
 sg13g2_inv_1 _12259_ (.Y(_04285_),
    .A(\TRNG.hash[222] ));
 sg13g2_inv_1 _12260_ (.Y(_04286_),
    .A(\TRNG.hash[218] ));
 sg13g2_inv_1 _12261_ (.Y(_04287_),
    .A(\TRNG.hash[212] ));
 sg13g2_inv_1 _12262_ (.Y(_04288_),
    .A(\TRNG.hash[190] ));
 sg13g2_inv_1 _12263_ (.Y(_04289_),
    .A(net3579));
 sg13g2_inv_1 _12264_ (.Y(_04290_),
    .A(\TRNG.hash[176] ));
 sg13g2_inv_1 _12265_ (.Y(_04291_),
    .A(\TRNG.hash[171] ));
 sg13g2_inv_1 _12266_ (.Y(_04292_),
    .A(\TRNG.hash[167] ));
 sg13g2_inv_1 _12267_ (.Y(_04293_),
    .A(\TRNG.hash[118] ));
 sg13g2_inv_1 _12268_ (.Y(_04294_),
    .A(\TRNG.hash[93] ));
 sg13g2_inv_1 _12269_ (.Y(_04295_),
    .A(net3558));
 sg13g2_inv_1 _12270_ (.Y(_04296_),
    .A(\TRNG.hash[42] ));
 sg13g2_inv_1 _12271_ (.Y(_04297_),
    .A(\TRNG.hash[16] ));
 sg13g2_inv_1 _12272_ (.Y(_04298_),
    .A(\TRNG.hash[156] ));
 sg13g2_inv_1 _12273_ (.Y(_04299_),
    .A(\TRNG.hash[137] ));
 sg13g2_inv_1 _12274_ (.Y(_04300_),
    .A(\TRNG.hash[135] ));
 sg13g2_inv_1 _12275_ (.Y(_04301_),
    .A(\TRNG.uart_tx_inst.ticks_counter[0] ));
 sg13g2_inv_1 _12276_ (.Y(_04302_),
    .A(\TRNG.uart_tx_inst.ticks_counter[1] ));
 sg13g2_inv_1 _12277_ (.Y(_04303_),
    .A(net3727));
 sg13g2_inv_8 _12278_ (.Y(_04304_),
    .A(net5539));
 sg13g2_inv_1 _12279_ (.Y(_04305_),
    .A(\TRNG.state[0] ));
 sg13g2_inv_1 _12280_ (.Y(_04306_),
    .A(net2936));
 sg13g2_inv_1 _12281_ (.Y(_04307_),
    .A(\TRNG.bit_counter[3] ));
 sg13g2_inv_1 _12282_ (.Y(_04308_),
    .A(net2557));
 sg13g2_inv_1 _12283_ (.Y(_04309_),
    .A(net3780));
 sg13g2_inv_1 _12284_ (.Y(_04310_),
    .A(net2354));
 sg13g2_inv_1 _12285_ (.Y(_04311_),
    .A(net2213));
 sg13g2_inv_1 _12286_ (.Y(_04312_),
    .A(net1980));
 sg13g2_inv_1 _12287_ (.Y(_04313_),
    .A(net2809));
 sg13g2_inv_1 _12288_ (.Y(_04314_),
    .A(\TRNG.Padded_Out[485] ));
 sg13g2_inv_1 _12289_ (.Y(_04315_),
    .A(net1508));
 sg13g2_inv_1 _12290_ (.Y(_04316_),
    .A(net1272));
 sg13g2_inv_1 _12291_ (.Y(_04317_),
    .A(net1663));
 sg13g2_inv_1 _12292_ (.Y(_04318_),
    .A(net2582));
 sg13g2_inv_1 _12293_ (.Y(_04319_),
    .A(net2480));
 sg13g2_inv_1 _12294_ (.Y(_04320_),
    .A(\TRNG.Padded_Out[491] ));
 sg13g2_inv_1 _12295_ (.Y(_04321_),
    .A(net2441));
 sg13g2_inv_1 _12296_ (.Y(_04322_),
    .A(net2293));
 sg13g2_inv_1 _12297_ (.Y(_04323_),
    .A(net2472));
 sg13g2_inv_1 _12298_ (.Y(_04324_),
    .A(net2666));
 sg13g2_inv_1 _12299_ (.Y(_04325_),
    .A(\TRNG.Padded_Out[496] ));
 sg13g2_inv_1 _12300_ (.Y(_04326_),
    .A(net2733));
 sg13g2_inv_1 _12301_ (.Y(_04327_),
    .A(\TRNG.Padded_Out[498] ));
 sg13g2_inv_1 _12302_ (.Y(_04328_),
    .A(net2685));
 sg13g2_inv_1 _12303_ (.Y(_04329_),
    .A(\TRNG.Padded_Out[500] ));
 sg13g2_inv_1 _12304_ (.Y(_04330_),
    .A(net2997));
 sg13g2_inv_1 _12305_ (.Y(_04331_),
    .A(net2700));
 sg13g2_inv_1 _12306_ (.Y(_04332_),
    .A(net2464));
 sg13g2_inv_1 _12307_ (.Y(_04333_),
    .A(net2575));
 sg13g2_inv_1 _12308_ (.Y(_04334_),
    .A(net2378));
 sg13g2_inv_1 _12309_ (.Y(_04335_),
    .A(net2580));
 sg13g2_inv_1 _12310_ (.Y(_04336_),
    .A(net1356));
 sg13g2_inv_1 _12311_ (.Y(_04337_),
    .A(net2364));
 sg13g2_inv_1 _12312_ (.Y(_04338_),
    .A(net2357));
 sg13g2_inv_1 _12313_ (.Y(_04339_),
    .A(net1608));
 sg13g2_inv_1 _12314_ (.Y(_04340_),
    .A(net3309));
 sg13g2_inv_4 _12315_ (.A(net5508),
    .Y(_04341_));
 sg13g2_inv_2 _12316_ (.Y(_04342_),
    .A(net5512));
 sg13g2_inv_1 _12317_ (.Y(_04343_),
    .A(net3544));
 sg13g2_inv_1 _12318_ (.Y(_04344_),
    .A(net3101));
 sg13g2_inv_1 _12319_ (.Y(_04345_),
    .A(net3105));
 sg13g2_inv_1 _12320_ (.Y(_04346_),
    .A(net3147));
 sg13g2_inv_1 _12321_ (.Y(_04347_),
    .A(net3071));
 sg13g2_inv_1 _12322_ (.Y(_04348_),
    .A(net3175));
 sg13g2_inv_1 _12323_ (.Y(_04349_),
    .A(net2950));
 sg13g2_inv_1 _12324_ (.Y(_04350_),
    .A(net2853));
 sg13g2_inv_1 _12325_ (.Y(_04351_),
    .A(net3005));
 sg13g2_inv_1 _12326_ (.Y(_04352_),
    .A(net2758));
 sg13g2_inv_1 _12327_ (.Y(_04353_),
    .A(net3007));
 sg13g2_inv_1 _12328_ (.Y(_04354_),
    .A(net2912));
 sg13g2_inv_1 _12329_ (.Y(_04355_),
    .A(net3032));
 sg13g2_inv_1 _12330_ (.Y(_04356_),
    .A(net3047));
 sg13g2_inv_1 _12331_ (.Y(_04357_),
    .A(net2735));
 sg13g2_inv_1 _12332_ (.Y(_04358_),
    .A(net3192));
 sg13g2_inv_1 _12333_ (.Y(_04359_),
    .A(net2898));
 sg13g2_inv_1 _12334_ (.Y(_04360_),
    .A(net2956));
 sg13g2_inv_1 _12335_ (.Y(_04361_),
    .A(net3140));
 sg13g2_inv_1 _12336_ (.Y(_04362_),
    .A(net2932));
 sg13g2_inv_1 _12337_ (.Y(_04363_),
    .A(net3096));
 sg13g2_inv_1 _12338_ (.Y(_04364_),
    .A(net3191));
 sg13g2_inv_1 _12339_ (.Y(_04365_),
    .A(net2864));
 sg13g2_inv_1 _12340_ (.Y(_04366_),
    .A(net3070));
 sg13g2_inv_1 _12341_ (.Y(_04367_),
    .A(net2934));
 sg13g2_inv_1 _12342_ (.Y(_04368_),
    .A(net3181));
 sg13g2_inv_1 _12343_ (.Y(_04369_),
    .A(net3208));
 sg13g2_inv_1 _12344_ (.Y(_04370_),
    .A(net3179));
 sg13g2_inv_1 _12345_ (.Y(_04371_),
    .A(net3023));
 sg13g2_inv_1 _12346_ (.Y(_04372_),
    .A(net3130));
 sg13g2_inv_1 _12347_ (.Y(_04373_),
    .A(net3164));
 sg13g2_inv_1 _12348_ (.Y(_04374_),
    .A(_00132_));
 sg13g2_inv_1 _12349_ (.Y(_04375_),
    .A(_00134_));
 sg13g2_inv_1 _12350_ (.Y(_04376_),
    .A(net3505));
 sg13g2_inv_1 _12351_ (.Y(_04377_),
    .A(net3654));
 sg13g2_inv_1 _12352_ (.Y(_04378_),
    .A(_00192_));
 sg13g2_inv_1 _12353_ (.Y(_04379_),
    .A(net3439));
 sg13g2_inv_1 _12354_ (.Y(_04380_),
    .A(_00230_));
 sg13g2_inv_1 _12355_ (.Y(_04381_),
    .A(net1864));
 sg13g2_inv_1 _12356_ (.Y(_04382_),
    .A(\TRNG.Word_Out[1] ));
 sg13g2_inv_2 _12357_ (.Y(_04383_),
    .A(net2611));
 sg13g2_inv_1 _12358_ (.Y(_04384_),
    .A(\TRNG.Word_Out[3] ));
 sg13g2_inv_1 _12359_ (.Y(_04385_),
    .A(net1937));
 sg13g2_inv_1 _12360_ (.Y(_04386_),
    .A(\TRNG.Word_Out[5] ));
 sg13g2_inv_1 _12361_ (.Y(_04387_),
    .A(net1820));
 sg13g2_inv_1 _12362_ (.Y(_04388_),
    .A(net1193));
 sg13g2_inv_1 _12363_ (.Y(_04389_),
    .A(\TRNG.Word_Out[8] ));
 sg13g2_inv_1 _12364_ (.Y(_04390_),
    .A(net1718));
 sg13g2_inv_1 _12365_ (.Y(_04391_),
    .A(\TRNG.Word_Out[10] ));
 sg13g2_inv_1 _12366_ (.Y(_04392_),
    .A(\TRNG.Word_Out[11] ));
 sg13g2_inv_1 _12367_ (.Y(_04393_),
    .A(\TRNG.Word_Out[12] ));
 sg13g2_inv_1 _12368_ (.Y(_04394_),
    .A(net1229));
 sg13g2_inv_1 _12369_ (.Y(_04395_),
    .A(\TRNG.Word_Out[14] ));
 sg13g2_inv_1 _12370_ (.Y(_04396_),
    .A(net1362));
 sg13g2_inv_1 _12371_ (.Y(_04397_),
    .A(\TRNG.Word_Out[16] ));
 sg13g2_inv_1 _12372_ (.Y(_04398_),
    .A(net1978));
 sg13g2_inv_1 _12373_ (.Y(_04399_),
    .A(\TRNG.Word_Out[18] ));
 sg13g2_inv_1 _12374_ (.Y(_04400_),
    .A(\TRNG.Word_Out[19] ));
 sg13g2_inv_1 _12375_ (.Y(_04401_),
    .A(net2757));
 sg13g2_inv_1 _12376_ (.Y(_04402_),
    .A(net2548));
 sg13g2_inv_1 _12377_ (.Y(_04403_),
    .A(net2129));
 sg13g2_inv_1 _12378_ (.Y(_04404_),
    .A(\TRNG.Word_Out[23] ));
 sg13g2_inv_1 _12379_ (.Y(_04405_),
    .A(net1150));
 sg13g2_inv_1 _12380_ (.Y(_04406_),
    .A(\TRNG.Word_Out[25] ));
 sg13g2_inv_1 _12381_ (.Y(_04407_),
    .A(net2280));
 sg13g2_inv_1 _12382_ (.Y(_04408_),
    .A(\TRNG.Word_Out[27] ));
 sg13g2_inv_1 _12383_ (.Y(_04409_),
    .A(\TRNG.Word_Out[28] ));
 sg13g2_inv_1 _12384_ (.Y(_04410_),
    .A(net1231));
 sg13g2_inv_1 _12385_ (.Y(_04411_),
    .A(net1191));
 sg13g2_inv_1 _12386_ (.Y(_04412_),
    .A(\TRNG.Word_Out[31] ));
 sg13g2_inv_1 _12387_ (.Y(_04413_),
    .A(\TRNG.Word_Out[32] ));
 sg13g2_inv_1 _12388_ (.Y(_04414_),
    .A(\TRNG.Word_Out[33] ));
 sg13g2_inv_1 _12389_ (.Y(_04415_),
    .A(\TRNG.Word_Out[34] ));
 sg13g2_inv_1 _12390_ (.Y(_04416_),
    .A(net2113));
 sg13g2_inv_1 _12391_ (.Y(_04417_),
    .A(net1223));
 sg13g2_inv_1 _12392_ (.Y(_04418_),
    .A(net2549));
 sg13g2_inv_1 _12393_ (.Y(_04419_),
    .A(net1239));
 sg13g2_inv_1 _12394_ (.Y(_04420_),
    .A(\TRNG.Word_Out[39] ));
 sg13g2_inv_1 _12395_ (.Y(_04421_),
    .A(net1653));
 sg13g2_inv_1 _12396_ (.Y(_04422_),
    .A(\TRNG.Word_Out[41] ));
 sg13g2_inv_1 _12397_ (.Y(_04423_),
    .A(net2850));
 sg13g2_inv_1 _12398_ (.Y(_04424_),
    .A(net2586));
 sg13g2_inv_1 _12399_ (.Y(_04425_),
    .A(net2268));
 sg13g2_inv_1 _12400_ (.Y(_04426_),
    .A(net2112));
 sg13g2_inv_1 _12401_ (.Y(_04427_),
    .A(net1821));
 sg13g2_inv_1 _12402_ (.Y(_04428_),
    .A(\TRNG.Word_Out[47] ));
 sg13g2_inv_1 _12403_ (.Y(_04429_),
    .A(\TRNG.Word_Out[48] ));
 sg13g2_inv_1 _12404_ (.Y(_04430_),
    .A(net2351));
 sg13g2_inv_1 _12405_ (.Y(_04431_),
    .A(net2108));
 sg13g2_inv_1 _12406_ (.Y(_04432_),
    .A(\TRNG.Word_Out[51] ));
 sg13g2_inv_1 _12407_ (.Y(_04433_),
    .A(net2244));
 sg13g2_inv_1 _12408_ (.Y(_04434_),
    .A(net1941));
 sg13g2_inv_1 _12409_ (.Y(_04435_),
    .A(\TRNG.Word_Out[54] ));
 sg13g2_inv_1 _12410_ (.Y(_04436_),
    .A(net1722));
 sg13g2_inv_1 _12411_ (.Y(_04437_),
    .A(\TRNG.Word_Out[56] ));
 sg13g2_inv_1 _12412_ (.Y(_04438_),
    .A(\TRNG.Word_Out[57] ));
 sg13g2_inv_1 _12413_ (.Y(_04439_),
    .A(net2578));
 sg13g2_inv_1 _12414_ (.Y(_04440_),
    .A(\TRNG.Word_Out[59] ));
 sg13g2_inv_1 _12415_ (.Y(_04441_),
    .A(net1215));
 sg13g2_inv_1 _12416_ (.Y(_04442_),
    .A(\TRNG.Word_Out[61] ));
 sg13g2_inv_1 _12417_ (.Y(_04443_),
    .A(net2106));
 sg13g2_inv_1 _12418_ (.Y(_04444_),
    .A(net1170));
 sg13g2_inv_1 _12419_ (.Y(_04445_),
    .A(\TRNG.Word_Out[64] ));
 sg13g2_inv_1 _12420_ (.Y(_04446_),
    .A(\TRNG.Word_Out[65] ));
 sg13g2_inv_1 _12421_ (.Y(_04447_),
    .A(net1857));
 sg13g2_inv_1 _12422_ (.Y(_04448_),
    .A(net2123));
 sg13g2_inv_1 _12423_ (.Y(_04449_),
    .A(\TRNG.Word_Out[68] ));
 sg13g2_inv_1 _12424_ (.Y(_04450_),
    .A(net2189));
 sg13g2_inv_1 _12425_ (.Y(_04451_),
    .A(net1206));
 sg13g2_inv_1 _12426_ (.Y(_04452_),
    .A(net1577));
 sg13g2_inv_1 _12427_ (.Y(_04453_),
    .A(net1724));
 sg13g2_inv_1 _12428_ (.Y(_04454_),
    .A(\TRNG.Word_Out[73] ));
 sg13g2_inv_1 _12429_ (.Y(_04455_),
    .A(net2153));
 sg13g2_inv_1 _12430_ (.Y(_04456_),
    .A(\TRNG.Word_Out[75] ));
 sg13g2_inv_1 _12431_ (.Y(_04457_),
    .A(net3193));
 sg13g2_inv_1 _12432_ (.Y(_04458_),
    .A(net2474));
 sg13g2_inv_1 _12433_ (.Y(_04459_),
    .A(net1200));
 sg13g2_inv_1 _12434_ (.Y(_04460_),
    .A(\TRNG.Word_Out[79] ));
 sg13g2_inv_1 _12435_ (.Y(_04461_),
    .A(\TRNG.Word_Out[80] ));
 sg13g2_inv_1 _12436_ (.Y(_04462_),
    .A(\TRNG.Word_Out[81] ));
 sg13g2_inv_1 _12437_ (.Y(_04463_),
    .A(\TRNG.Word_Out[82] ));
 sg13g2_inv_1 _12438_ (.Y(_04464_),
    .A(\TRNG.Word_Out[83] ));
 sg13g2_inv_1 _12439_ (.Y(_04465_),
    .A(net2284));
 sg13g2_inv_1 _12440_ (.Y(_04466_),
    .A(\TRNG.Word_Out[85] ));
 sg13g2_inv_1 _12441_ (.Y(_04467_),
    .A(net2211));
 sg13g2_inv_1 _12442_ (.Y(_04468_),
    .A(net1341));
 sg13g2_inv_1 _12443_ (.Y(_04469_),
    .A(net1241));
 sg13g2_inv_1 _12444_ (.Y(_04470_),
    .A(\TRNG.Word_Out[89] ));
 sg13g2_inv_1 _12445_ (.Y(_04471_),
    .A(net2202));
 sg13g2_inv_1 _12446_ (.Y(_04472_),
    .A(\TRNG.Word_Out[91] ));
 sg13g2_inv_1 _12447_ (.Y(_04473_),
    .A(\TRNG.Word_Out[92] ));
 sg13g2_inv_1 _12448_ (.Y(_04474_),
    .A(net1176));
 sg13g2_inv_1 _12449_ (.Y(_04475_),
    .A(\TRNG.Word_Out[94] ));
 sg13g2_inv_1 _12450_ (.Y(_04476_),
    .A(net2058));
 sg13g2_inv_1 _12451_ (.Y(_04477_),
    .A(\TRNG.Word_Out[96] ));
 sg13g2_inv_1 _12452_ (.Y(_04478_),
    .A(net2075));
 sg13g2_inv_1 _12453_ (.Y(_04479_),
    .A(net1816));
 sg13g2_inv_1 _12454_ (.Y(_04480_),
    .A(\TRNG.Word_Out[99] ));
 sg13g2_inv_1 _12455_ (.Y(_04481_),
    .A(net1879));
 sg13g2_inv_1 _12456_ (.Y(_04482_),
    .A(\TRNG.Word_Out[101] ));
 sg13g2_inv_1 _12457_ (.Y(_04483_),
    .A(net1736));
 sg13g2_inv_1 _12458_ (.Y(_04484_),
    .A(net1182));
 sg13g2_inv_1 _12459_ (.Y(_04485_),
    .A(\TRNG.Word_Out[104] ));
 sg13g2_inv_1 _12460_ (.Y(_04486_),
    .A(\TRNG.Word_Out[105] ));
 sg13g2_inv_1 _12461_ (.Y(_04487_),
    .A(\TRNG.Word_Out[106] ));
 sg13g2_inv_1 _12462_ (.Y(_04488_),
    .A(net1832));
 sg13g2_inv_1 _12463_ (.Y(_04489_),
    .A(\TRNG.Word_Out[108] ));
 sg13g2_inv_1 _12464_ (.Y(_04490_),
    .A(\TRNG.Word_Out[109] ));
 sg13g2_inv_1 _12465_ (.Y(_04491_),
    .A(net1964));
 sg13g2_inv_1 _12466_ (.Y(_04492_),
    .A(net1506));
 sg13g2_inv_1 _12467_ (.Y(_04493_),
    .A(net1225));
 sg13g2_inv_1 _12468_ (.Y(_04494_),
    .A(net1461));
 sg13g2_inv_1 _12469_ (.Y(_04495_),
    .A(\TRNG.Word_Out[114] ));
 sg13g2_inv_1 _12470_ (.Y(_04496_),
    .A(net2267));
 sg13g2_inv_1 _12471_ (.Y(_04497_),
    .A(net2240));
 sg13g2_inv_1 _12472_ (.Y(_04498_),
    .A(\TRNG.Word_Out[117] ));
 sg13g2_inv_1 _12473_ (.Y(_04499_),
    .A(net2014));
 sg13g2_inv_1 _12474_ (.Y(_04500_),
    .A(\TRNG.Word_Out[119] ));
 sg13g2_inv_1 _12475_ (.Y(_04501_),
    .A(net1549));
 sg13g2_inv_1 _12476_ (.Y(_04502_),
    .A(net1681));
 sg13g2_inv_1 _12477_ (.Y(_04503_),
    .A(net2070));
 sg13g2_inv_1 _12478_ (.Y(_04504_),
    .A(net2287));
 sg13g2_inv_1 _12479_ (.Y(_04505_),
    .A(net2242));
 sg13g2_inv_1 _12480_ (.Y(_04506_),
    .A(net1217));
 sg13g2_inv_1 _12481_ (.Y(_04507_),
    .A(\TRNG.Word_Out[126] ));
 sg13g2_inv_1 _12482_ (.Y(_04508_),
    .A(net1152));
 sg13g2_inv_1 _12483_ (.Y(_04509_),
    .A(net1927));
 sg13g2_inv_1 _12484_ (.Y(_04510_),
    .A(\TRNG.Word_Out[129] ));
 sg13g2_inv_1 _12485_ (.Y(_04511_),
    .A(net2786));
 sg13g2_inv_1 _12486_ (.Y(_04512_),
    .A(net1367));
 sg13g2_inv_1 _12487_ (.Y(_04513_),
    .A(\TRNG.Word_Out[132] ));
 sg13g2_inv_1 _12488_ (.Y(_04514_),
    .A(net1160));
 sg13g2_inv_1 _12489_ (.Y(_04515_),
    .A(\TRNG.Word_Out[134] ));
 sg13g2_inv_1 _12490_ (.Y(_04516_),
    .A(net1221));
 sg13g2_inv_1 _12491_ (.Y(_04517_),
    .A(\TRNG.Word_Out[136] ));
 sg13g2_inv_1 _12492_ (.Y(_04518_),
    .A(net2118));
 sg13g2_inv_1 _12493_ (.Y(_04519_),
    .A(net1144));
 sg13g2_inv_1 _12494_ (.Y(_04520_),
    .A(\TRNG.Word_Out[139] ));
 sg13g2_inv_1 _12495_ (.Y(_04521_),
    .A(\TRNG.Word_Out[140] ));
 sg13g2_inv_1 _12496_ (.Y(_04522_),
    .A(net1162));
 sg13g2_inv_1 _12497_ (.Y(_04523_),
    .A(\TRNG.Word_Out[142] ));
 sg13g2_inv_1 _12498_ (.Y(_04524_),
    .A(\TRNG.Word_Out[143] ));
 sg13g2_inv_1 _12499_ (.Y(_04525_),
    .A(\TRNG.Word_Out[144] ));
 sg13g2_inv_1 _12500_ (.Y(_04526_),
    .A(\TRNG.Word_Out[145] ));
 sg13g2_inv_1 _12501_ (.Y(_04527_),
    .A(\TRNG.Word_Out[146] ));
 sg13g2_inv_1 _12502_ (.Y(_04528_),
    .A(net2396));
 sg13g2_inv_1 _12503_ (.Y(_04529_),
    .A(\TRNG.Word_Out[148] ));
 sg13g2_inv_1 _12504_ (.Y(_04530_),
    .A(net1541));
 sg13g2_inv_1 _12505_ (.Y(_04531_),
    .A(net1866));
 sg13g2_inv_1 _12506_ (.Y(_04532_),
    .A(net1921));
 sg13g2_inv_1 _12507_ (.Y(_04533_),
    .A(\TRNG.Word_Out[152] ));
 sg13g2_inv_1 _12508_ (.Y(_04534_),
    .A(\TRNG.Word_Out[153] ));
 sg13g2_inv_1 _12509_ (.Y(_04535_),
    .A(net1189));
 sg13g2_inv_1 _12510_ (.Y(_04536_),
    .A(\TRNG.Word_Out[155] ));
 sg13g2_inv_1 _12511_ (.Y(_04537_),
    .A(net2454));
 sg13g2_inv_1 _12512_ (.Y(_04538_),
    .A(net1236));
 sg13g2_inv_1 _12513_ (.Y(_04539_),
    .A(net1960));
 sg13g2_inv_1 _12514_ (.Y(_04540_),
    .A(\TRNG.Word_Out[159] ));
 sg13g2_inv_1 _12515_ (.Y(_04541_),
    .A(\TRNG.Word_Out[160] ));
 sg13g2_inv_1 _12516_ (.Y(_04542_),
    .A(net2410));
 sg13g2_inv_1 _12517_ (.Y(_04543_),
    .A(\TRNG.Word_Out[162] ));
 sg13g2_inv_1 _12518_ (.Y(_04544_),
    .A(net1823));
 sg13g2_inv_1 _12519_ (.Y(_04545_),
    .A(net1579));
 sg13g2_inv_1 _12520_ (.Y(_04546_),
    .A(\TRNG.Word_Out[165] ));
 sg13g2_inv_1 _12521_ (.Y(_04547_),
    .A(net1493));
 sg13g2_inv_1 _12522_ (.Y(_04548_),
    .A(\TRNG.Word_Out[167] ));
 sg13g2_inv_1 _12523_ (.Y(_04549_),
    .A(\TRNG.Word_Out[168] ));
 sg13g2_inv_1 _12524_ (.Y(_04550_),
    .A(net1569));
 sg13g2_inv_1 _12525_ (.Y(_04551_),
    .A(\TRNG.Word_Out[170] ));
 sg13g2_inv_1 _12526_ (.Y(_04552_),
    .A(\TRNG.Word_Out[171] ));
 sg13g2_inv_1 _12527_ (.Y(_04553_),
    .A(net2233));
 sg13g2_inv_1 _12528_ (.Y(_04554_),
    .A(\TRNG.Word_Out[173] ));
 sg13g2_inv_1 _12529_ (.Y(_04555_),
    .A(net1156));
 sg13g2_inv_1 _12530_ (.Y(_04556_),
    .A(\TRNG.Word_Out[175] ));
 sg13g2_inv_1 _12531_ (.Y(_04557_),
    .A(\TRNG.Word_Out[176] ));
 sg13g2_inv_1 _12532_ (.Y(_04558_),
    .A(net2103));
 sg13g2_inv_1 _12533_ (.Y(_04559_),
    .A(\TRNG.Word_Out[178] ));
 sg13g2_inv_1 _12534_ (.Y(_04560_),
    .A(net2465));
 sg13g2_inv_1 _12535_ (.Y(_04561_),
    .A(\TRNG.Word_Out[180] ));
 sg13g2_inv_1 _12536_ (.Y(_04562_),
    .A(net2054));
 sg13g2_inv_1 _12537_ (.Y(_04563_),
    .A(\TRNG.Word_Out[182] ));
 sg13g2_inv_1 _12538_ (.Y(_04564_),
    .A(net2219));
 sg13g2_inv_1 _12539_ (.Y(_04565_),
    .A(\TRNG.Word_Out[184] ));
 sg13g2_inv_1 _12540_ (.Y(_04566_),
    .A(net1954));
 sg13g2_inv_1 _12541_ (.Y(_04567_),
    .A(\TRNG.Word_Out[186] ));
 sg13g2_inv_1 _12542_ (.Y(_04568_),
    .A(\TRNG.Word_Out[187] ));
 sg13g2_inv_1 _12543_ (.Y(_04569_),
    .A(\TRNG.Word_Out[188] ));
 sg13g2_inv_1 _12544_ (.Y(_04570_),
    .A(net1202));
 sg13g2_inv_1 _12545_ (.Y(_04571_),
    .A(\TRNG.Word_Out[190] ));
 sg13g2_inv_1 _12546_ (.Y(_04572_),
    .A(\TRNG.Word_Out[191] ));
 sg13g2_inv_1 _12547_ (.Y(_04573_),
    .A(net1133));
 sg13g2_inv_1 _12548_ (.Y(_04574_),
    .A(\TRNG.Word_Out[193] ));
 sg13g2_inv_1 _12549_ (.Y(_04575_),
    .A(net2875));
 sg13g2_inv_1 _12550_ (.Y(_04576_),
    .A(net1962));
 sg13g2_inv_1 _12551_ (.Y(_04577_),
    .A(\TRNG.Word_Out[196] ));
 sg13g2_inv_1 _12552_ (.Y(_04578_),
    .A(net1573));
 sg13g2_inv_1 _12553_ (.Y(_04579_),
    .A(\TRNG.Word_Out[198] ));
 sg13g2_inv_1 _12554_ (.Y(_04580_),
    .A(\TRNG.Word_Out[199] ));
 sg13g2_inv_1 _12555_ (.Y(_04581_),
    .A(net1280));
 sg13g2_inv_1 _12556_ (.Y(_04582_),
    .A(\TRNG.Word_Out[201] ));
 sg13g2_inv_1 _12557_ (.Y(_04583_),
    .A(\TRNG.Word_Out[202] ));
 sg13g2_inv_1 _12558_ (.Y(_04584_),
    .A(net3044));
 sg13g2_inv_1 _12559_ (.Y(_04585_),
    .A(net2648));
 sg13g2_inv_1 _12560_ (.Y(_04586_),
    .A(net2105));
 sg13g2_inv_1 _12561_ (.Y(_04587_),
    .A(net2005));
 sg13g2_inv_1 _12562_ (.Y(_04588_),
    .A(\TRNG.Word_Out[207] ));
 sg13g2_inv_1 _12563_ (.Y(_04589_),
    .A(net1891));
 sg13g2_inv_1 _12564_ (.Y(_04590_),
    .A(\TRNG.Word_Out[209] ));
 sg13g2_inv_1 _12565_ (.Y(_04591_),
    .A(\TRNG.Word_Out[210] ));
 sg13g2_inv_1 _12566_ (.Y(_04592_),
    .A(\TRNG.Word_Out[211] ));
 sg13g2_inv_1 _12567_ (.Y(_04593_),
    .A(net2564));
 sg13g2_inv_1 _12568_ (.Y(_04594_),
    .A(net2446));
 sg13g2_inv_1 _12569_ (.Y(_04595_),
    .A(\TRNG.Word_Out[214] ));
 sg13g2_inv_1 _12570_ (.Y(_04596_),
    .A(net1904));
 sg13g2_inv_1 _12571_ (.Y(_04597_),
    .A(net2225));
 sg13g2_inv_1 _12572_ (.Y(_04598_),
    .A(net2017));
 sg13g2_inv_1 _12573_ (.Y(_04599_),
    .A(net1994));
 sg13g2_inv_1 _12574_ (.Y(_04600_),
    .A(\TRNG.Word_Out[219] ));
 sg13g2_inv_1 _12575_ (.Y(_04601_),
    .A(net2366));
 sg13g2_inv_1 _12576_ (.Y(_04602_),
    .A(\TRNG.Word_Out[221] ));
 sg13g2_inv_1 _12577_ (.Y(_04603_),
    .A(net1947));
 sg13g2_inv_1 _12578_ (.Y(_04604_),
    .A(\TRNG.Word_Out[223] ));
 sg13g2_inv_1 _12579_ (.Y(_04605_),
    .A(net1158));
 sg13g2_inv_1 _12580_ (.Y(_04606_),
    .A(\TRNG.Word_Out[225] ));
 sg13g2_inv_1 _12581_ (.Y(_04607_),
    .A(net3229));
 sg13g2_inv_1 _12582_ (.Y(_04608_),
    .A(net1956));
 sg13g2_inv_1 _12583_ (.Y(_04609_),
    .A(net1208));
 sg13g2_inv_1 _12584_ (.Y(_04610_),
    .A(\TRNG.Word_Out[229] ));
 sg13g2_inv_1 _12585_ (.Y(_04611_),
    .A(net2283));
 sg13g2_inv_1 _12586_ (.Y(_04612_),
    .A(net1836));
 sg13g2_inv_1 _12587_ (.Y(_04613_),
    .A(net2204));
 sg13g2_inv_1 _12588_ (.Y(_04614_),
    .A(\TRNG.Word_Out[233] ));
 sg13g2_inv_1 _12589_ (.Y(_04615_),
    .A(net2274));
 sg13g2_inv_1 _12590_ (.Y(_04616_),
    .A(\TRNG.Word_Out[235] ));
 sg13g2_inv_1 _12591_ (.Y(_04617_),
    .A(\TRNG.Word_Out[236] ));
 sg13g2_inv_1 _12592_ (.Y(_04618_),
    .A(net2243));
 sg13g2_inv_1 _12593_ (.Y(_04619_),
    .A(net2094));
 sg13g2_inv_1 _12594_ (.Y(_04620_),
    .A(\TRNG.Word_Out[239] ));
 sg13g2_inv_1 _12595_ (.Y(_04621_),
    .A(net1428));
 sg13g2_inv_1 _12596_ (.Y(_04622_),
    .A(net2339));
 sg13g2_inv_1 _12597_ (.Y(_04623_),
    .A(\TRNG.Word_Out[242] ));
 sg13g2_inv_1 _12598_ (.Y(_04624_),
    .A(net3127));
 sg13g2_inv_1 _12599_ (.Y(_04625_),
    .A(net2488));
 sg13g2_inv_1 _12600_ (.Y(_04626_),
    .A(net2425));
 sg13g2_inv_1 _12601_ (.Y(_04627_),
    .A(\TRNG.Word_Out[246] ));
 sg13g2_inv_1 _12602_ (.Y(_04628_),
    .A(net1560));
 sg13g2_inv_1 _12603_ (.Y(_04629_),
    .A(\TRNG.Word_Out[248] ));
 sg13g2_inv_1 _12604_ (.Y(_04630_),
    .A(net1348));
 sg13g2_inv_1 _12605_ (.Y(_04631_),
    .A(\TRNG.Word_Out[250] ));
 sg13g2_inv_1 _12606_ (.Y(_04632_),
    .A(net2431));
 sg13g2_inv_1 _12607_ (.Y(_04633_),
    .A(\TRNG.Word_Out[252] ));
 sg13g2_inv_1 _12608_ (.Y(_04634_),
    .A(net2254));
 sg13g2_inv_1 _12609_ (.Y(_04635_),
    .A(net1195));
 sg13g2_inv_1 _12610_ (.Y(_04636_),
    .A(\TRNG.Word_Out[255] ));
 sg13g2_inv_1 _12611_ (.Y(_04637_),
    .A(net2206));
 sg13g2_inv_1 _12612_ (.Y(_04638_),
    .A(\TRNG.Word_Out[257] ));
 sg13g2_inv_1 _12613_ (.Y(_04639_),
    .A(net1851));
 sg13g2_inv_1 _12614_ (.Y(_04640_),
    .A(\TRNG.Word_Out[259] ));
 sg13g2_inv_1 _12615_ (.Y(_04641_),
    .A(net1759));
 sg13g2_inv_1 _12616_ (.Y(_04642_),
    .A(\TRNG.Word_Out[261] ));
 sg13g2_inv_1 _12617_ (.Y(_04643_),
    .A(net1788));
 sg13g2_inv_1 _12618_ (.Y(_04644_),
    .A(net1371));
 sg13g2_inv_1 _12619_ (.Y(_04645_),
    .A(net2188));
 sg13g2_inv_1 _12620_ (.Y(_04646_),
    .A(net1253));
 sg13g2_inv_1 _12621_ (.Y(_04647_),
    .A(\TRNG.Word_Out[266] ));
 sg13g2_inv_1 _12622_ (.Y(_04648_),
    .A(\TRNG.Word_Out[267] ));
 sg13g2_inv_1 _12623_ (.Y(_04649_),
    .A(\TRNG.Word_Out[268] ));
 sg13g2_inv_1 _12624_ (.Y(_04650_),
    .A(\TRNG.Word_Out[269] ));
 sg13g2_inv_1 _12625_ (.Y(_04651_),
    .A(net1998));
 sg13g2_inv_1 _12626_ (.Y(_04652_),
    .A(\TRNG.Word_Out[271] ));
 sg13g2_inv_1 _12627_ (.Y(_04653_),
    .A(net2081));
 sg13g2_inv_1 _12628_ (.Y(_04654_),
    .A(\TRNG.Word_Out[273] ));
 sg13g2_inv_1 _12629_ (.Y(_04655_),
    .A(net2436));
 sg13g2_inv_1 _12630_ (.Y(_04656_),
    .A(\TRNG.Word_Out[275] ));
 sg13g2_inv_1 _12631_ (.Y(_04657_),
    .A(\TRNG.Word_Out[276] ));
 sg13g2_inv_1 _12632_ (.Y(_04658_),
    .A(net2865));
 sg13g2_inv_1 _12633_ (.Y(_04659_),
    .A(net2380));
 sg13g2_inv_1 _12634_ (.Y(_04660_),
    .A(\TRNG.Word_Out[279] ));
 sg13g2_inv_1 _12635_ (.Y(_04661_),
    .A(net1138));
 sg13g2_inv_1 _12636_ (.Y(_04662_),
    .A(\TRNG.Word_Out[281] ));
 sg13g2_inv_1 _12637_ (.Y(_04663_),
    .A(net2669));
 sg13g2_inv_1 _12638_ (.Y(_04664_),
    .A(net1935));
 sg13g2_inv_1 _12639_ (.Y(_04665_),
    .A(\TRNG.Word_Out[284] ));
 sg13g2_inv_1 _12640_ (.Y(_04666_),
    .A(net1410));
 sg13g2_inv_1 _12641_ (.Y(_04667_),
    .A(\TRNG.Word_Out[286] ));
 sg13g2_inv_1 _12642_ (.Y(_04668_),
    .A(\TRNG.Word_Out[287] ));
 sg13g2_inv_1 _12643_ (.Y(_04669_),
    .A(net2286));
 sg13g2_inv_1 _12644_ (.Y(_04670_),
    .A(net1751));
 sg13g2_inv_1 _12645_ (.Y(_04671_),
    .A(\TRNG.Word_Out[290] ));
 sg13g2_inv_1 _12646_ (.Y(_04672_),
    .A(net1212));
 sg13g2_inv_1 _12647_ (.Y(_04673_),
    .A(\TRNG.Word_Out[292] ));
 sg13g2_inv_1 _12648_ (.Y(_04674_),
    .A(\TRNG.Word_Out[293] ));
 sg13g2_inv_1 _12649_ (.Y(_04675_),
    .A(net1245));
 sg13g2_inv_1 _12650_ (.Y(_04676_),
    .A(net1911));
 sg13g2_inv_1 _12651_ (.Y(_04677_),
    .A(\TRNG.Word_Out[296] ));
 sg13g2_inv_1 _12652_ (.Y(_04678_),
    .A(net2121));
 sg13g2_inv_1 _12653_ (.Y(_04679_),
    .A(\TRNG.Word_Out[298] ));
 sg13g2_inv_1 _12654_ (.Y(_04680_),
    .A(\TRNG.Word_Out[299] ));
 sg13g2_inv_1 _12655_ (.Y(_04681_),
    .A(\TRNG.Word_Out[300] ));
 sg13g2_inv_1 _12656_ (.Y(_04682_),
    .A(net2730));
 sg13g2_inv_1 _12657_ (.Y(_04683_),
    .A(net2237));
 sg13g2_inv_1 _12658_ (.Y(_04684_),
    .A(net1298));
 sg13g2_inv_1 _12659_ (.Y(_04685_),
    .A(\TRNG.Word_Out[304] ));
 sg13g2_inv_1 _12660_ (.Y(_04686_),
    .A(net2349));
 sg13g2_inv_1 _12661_ (.Y(_04687_),
    .A(\TRNG.Word_Out[306] ));
 sg13g2_inv_1 _12662_ (.Y(_04688_),
    .A(net2916));
 sg13g2_inv_1 _12663_ (.Y(_04689_),
    .A(net2683));
 sg13g2_inv_1 _12664_ (.Y(_04690_),
    .A(net2034));
 sg13g2_inv_1 _12665_ (.Y(_04691_),
    .A(\TRNG.Word_Out[310] ));
 sg13g2_inv_1 _12666_ (.Y(_04692_),
    .A(\TRNG.Word_Out[311] ));
 sg13g2_inv_1 _12667_ (.Y(_04693_),
    .A(net1198));
 sg13g2_inv_1 _12668_ (.Y(_04694_),
    .A(net1286));
 sg13g2_inv_1 _12669_ (.Y(_04695_),
    .A(net2255));
 sg13g2_inv_1 _12670_ (.Y(_04696_),
    .A(net2356));
 sg13g2_inv_1 _12671_ (.Y(_04697_),
    .A(net2627));
 sg13g2_inv_1 _12672_ (.Y(_04698_),
    .A(net1959));
 sg13g2_inv_1 _12673_ (.Y(_04699_),
    .A(net1290));
 sg13g2_inv_1 _12674_ (.Y(_04700_),
    .A(\TRNG.Word_Out[319] ));
 sg13g2_inv_1 _12675_ (.Y(_04701_),
    .A(\TRNG.Word_Out[320] ));
 sg13g2_inv_1 _12676_ (.Y(_04702_),
    .A(net1140));
 sg13g2_inv_1 _12677_ (.Y(_04703_),
    .A(net1166));
 sg13g2_inv_1 _12678_ (.Y(_04704_),
    .A(net1197));
 sg13g2_inv_1 _12679_ (.Y(_04705_),
    .A(net1172));
 sg13g2_inv_1 _12680_ (.Y(_04706_),
    .A(\TRNG.Word_Out[325] ));
 sg13g2_inv_1 _12681_ (.Y(_04707_),
    .A(net1602));
 sg13g2_inv_1 _12682_ (.Y(_04708_),
    .A(net1393));
 sg13g2_inv_1 _12683_ (.Y(_04709_),
    .A(\TRNG.Word_Out[328] ));
 sg13g2_inv_1 _12684_ (.Y(_04710_),
    .A(\TRNG.Word_Out[329] ));
 sg13g2_inv_1 _12685_ (.Y(_04711_),
    .A(net3098));
 sg13g2_inv_1 _12686_ (.Y(_04712_),
    .A(net2556));
 sg13g2_inv_1 _12687_ (.Y(_04713_),
    .A(net1680));
 sg13g2_inv_1 _12688_ (.Y(_04714_),
    .A(net1154));
 sg13g2_inv_1 _12689_ (.Y(_04715_),
    .A(\TRNG.Word_Out[334] ));
 sg13g2_inv_1 _12690_ (.Y(_04716_),
    .A(\TRNG.Word_Out[335] ));
 sg13g2_inv_1 _12691_ (.Y(_04717_),
    .A(net2199));
 sg13g2_inv_1 _12692_ (.Y(_04718_),
    .A(\TRNG.Word_Out[337] ));
 sg13g2_inv_1 _12693_ (.Y(_04719_),
    .A(net2629));
 sg13g2_inv_1 _12694_ (.Y(_04720_),
    .A(\TRNG.Word_Out[339] ));
 sg13g2_inv_1 _12695_ (.Y(_04721_),
    .A(net2770));
 sg13g2_inv_1 _12696_ (.Y(_04722_),
    .A(net2597));
 sg13g2_inv_1 _12697_ (.Y(_04723_),
    .A(net2184));
 sg13g2_inv_1 _12698_ (.Y(_04724_),
    .A(\TRNG.Word_Out[343] ));
 sg13g2_inv_1 _12699_ (.Y(_04725_),
    .A(net2292));
 sg13g2_inv_1 _12700_ (.Y(_04726_),
    .A(net1164));
 sg13g2_inv_1 _12701_ (.Y(_04727_),
    .A(\TRNG.Word_Out[346] ));
 sg13g2_inv_1 _12702_ (.Y(_04728_),
    .A(net2461));
 sg13g2_inv_1 _12703_ (.Y(_04729_),
    .A(net1185));
 sg13g2_inv_1 _12704_ (.Y(_04730_),
    .A(net1381));
 sg13g2_inv_1 _12705_ (.Y(_04731_),
    .A(\TRNG.Word_Out[350] ));
 sg13g2_inv_1 _12706_ (.Y(_04732_),
    .A(\TRNG.Word_Out[351] ));
 sg13g2_inv_1 _12707_ (.Y(_04733_),
    .A(net2087));
 sg13g2_inv_1 _12708_ (.Y(_04734_),
    .A(net2071));
 sg13g2_inv_1 _12709_ (.Y(_04735_),
    .A(\TRNG.Word_Out[354] ));
 sg13g2_inv_1 _12710_ (.Y(_04736_),
    .A(net1187));
 sg13g2_inv_1 _12711_ (.Y(_04737_),
    .A(\TRNG.Word_Out[356] ));
 sg13g2_inv_1 _12712_ (.Y(_04738_),
    .A(net1599));
 sg13g2_inv_1 _12713_ (.Y(_04739_),
    .A(\TRNG.Word_Out[358] ));
 sg13g2_inv_1 _12714_ (.Y(_04740_),
    .A(net1219));
 sg13g2_inv_1 _12715_ (.Y(_04741_),
    .A(\TRNG.Word_Out[360] ));
 sg13g2_inv_1 _12716_ (.Y(_04742_),
    .A(net2588));
 sg13g2_inv_1 _12717_ (.Y(_04743_),
    .A(\TRNG.Word_Out[362] ));
 sg13g2_inv_1 _12718_ (.Y(_04744_),
    .A(net1982));
 sg13g2_inv_1 _12719_ (.Y(_04745_),
    .A(\TRNG.Word_Out[364] ));
 sg13g2_inv_1 _12720_ (.Y(_04746_),
    .A(net2139));
 sg13g2_inv_1 _12721_ (.Y(_04747_),
    .A(\TRNG.Word_Out[366] ));
 sg13g2_inv_1 _12722_ (.Y(_04748_),
    .A(\TRNG.Word_Out[367] ));
 sg13g2_inv_1 _12723_ (.Y(_04749_),
    .A(net2128));
 sg13g2_inv_1 _12724_ (.Y(_04750_),
    .A(net1985));
 sg13g2_inv_1 _12725_ (.Y(_04751_),
    .A(\TRNG.Word_Out[370] ));
 sg13g2_inv_1 _12726_ (.Y(_04752_),
    .A(net2584));
 sg13g2_inv_1 _12727_ (.Y(_04753_),
    .A(\TRNG.Word_Out[372] ));
 sg13g2_inv_1 _12728_ (.Y(_04754_),
    .A(net2414));
 sg13g2_inv_1 _12729_ (.Y(_04755_),
    .A(net2228));
 sg13g2_inv_1 _12730_ (.Y(_04756_),
    .A(net2078));
 sg13g2_inv_1 _12731_ (.Y(_04757_),
    .A(net1178));
 sg13g2_inv_1 _12732_ (.Y(_04758_),
    .A(\TRNG.Word_Out[377] ));
 sg13g2_inv_1 _12733_ (.Y(_04759_),
    .A(net2455));
 sg13g2_inv_1 _12734_ (.Y(_04760_),
    .A(\TRNG.Word_Out[379] ));
 sg13g2_inv_1 _12735_ (.Y(_04761_),
    .A(net2497));
 sg13g2_inv_1 _12736_ (.Y(_04762_),
    .A(net1204));
 sg13g2_inv_1 _12737_ (.Y(_04763_),
    .A(\TRNG.Word_Out[382] ));
 sg13g2_inv_1 _12738_ (.Y(_04764_),
    .A(net2689));
 sg13g2_inv_1 _12739_ (.Y(_04765_),
    .A(net1818));
 sg13g2_inv_1 _12740_ (.Y(_04766_),
    .A(\TRNG.Word_Out[385] ));
 sg13g2_inv_1 _12741_ (.Y(_04767_),
    .A(\TRNG.Word_Out[386] ));
 sg13g2_inv_1 _12742_ (.Y(_04768_),
    .A(net1607));
 sg13g2_inv_1 _12743_ (.Y(_04769_),
    .A(net1425));
 sg13g2_inv_1 _12744_ (.Y(_04770_),
    .A(net1174));
 sg13g2_inv_1 _12745_ (.Y(_04771_),
    .A(net1661));
 sg13g2_inv_1 _12746_ (.Y(_04772_),
    .A(\TRNG.Word_Out[391] ));
 sg13g2_inv_1 _12747_ (.Y(_04773_),
    .A(\TRNG.Word_Out[392] ));
 sg13g2_inv_1 _12748_ (.Y(_04774_),
    .A(net1232));
 sg13g2_inv_1 _12749_ (.Y(_04775_),
    .A(\TRNG.Word_Out[394] ));
 sg13g2_inv_1 _12750_ (.Y(_04776_),
    .A(net1387));
 sg13g2_inv_1 _12751_ (.Y(_04777_),
    .A(\TRNG.Word_Out[396] ));
 sg13g2_inv_1 _12752_ (.Y(_04778_),
    .A(net1227));
 sg13g2_inv_1 _12753_ (.Y(_04779_),
    .A(\TRNG.Word_Out[398] ));
 sg13g2_inv_1 _12754_ (.Y(_04780_),
    .A(\TRNG.Word_Out[399] ));
 sg13g2_inv_1 _12755_ (.Y(_04781_),
    .A(net1471));
 sg13g2_inv_1 _12756_ (.Y(_04782_),
    .A(\TRNG.Word_Out[401] ));
 sg13g2_inv_1 _12757_ (.Y(_04783_),
    .A(\TRNG.Word_Out[402] ));
 sg13g2_inv_1 _12758_ (.Y(_04784_),
    .A(\TRNG.Word_Out[403] ));
 sg13g2_inv_1 _12759_ (.Y(_04785_),
    .A(net2881));
 sg13g2_inv_1 _12760_ (.Y(_04786_),
    .A(net1874));
 sg13g2_inv_1 _12761_ (.Y(_04787_),
    .A(\TRNG.Word_Out[406] ));
 sg13g2_inv_1 _12762_ (.Y(_04788_),
    .A(\TRNG.Word_Out[407] ));
 sg13g2_inv_1 _12763_ (.Y(_04789_),
    .A(net2490));
 sg13g2_inv_1 _12764_ (.Y(_04790_),
    .A(net1168));
 sg13g2_inv_1 _12765_ (.Y(_04791_),
    .A(\TRNG.Word_Out[410] ));
 sg13g2_inv_1 _12766_ (.Y(_04792_),
    .A(net2943));
 sg13g2_inv_1 _12767_ (.Y(_04793_),
    .A(net2641));
 sg13g2_inv_1 _12768_ (.Y(_04794_),
    .A(net1398));
 sg13g2_inv_1 _12769_ (.Y(_04795_),
    .A(\TRNG.Word_Out[414] ));
 sg13g2_inv_1 _12770_ (.Y(_04796_),
    .A(net2030));
 sg13g2_inv_1 _12771_ (.Y(_04797_),
    .A(\TRNG.Word_Out[416] ));
 sg13g2_inv_1 _12772_ (.Y(_04798_),
    .A(net2161));
 sg13g2_inv_1 _12773_ (.Y(_04799_),
    .A(\TRNG.Word_Out[418] ));
 sg13g2_inv_1 _12774_ (.Y(_04800_),
    .A(net2755));
 sg13g2_inv_1 _12775_ (.Y(_04801_),
    .A(net1633));
 sg13g2_inv_1 _12776_ (.Y(_04802_),
    .A(\TRNG.Word_Out[421] ));
 sg13g2_inv_1 _12777_ (.Y(_04803_),
    .A(net2245));
 sg13g2_inv_1 _12778_ (.Y(_04804_),
    .A(net2024));
 sg13g2_inv_1 _12779_ (.Y(_04805_),
    .A(net2231));
 sg13g2_inv_1 _12780_ (.Y(_04806_),
    .A(\TRNG.Word_Out[425] ));
 sg13g2_inv_1 _12781_ (.Y(_04807_),
    .A(net1469));
 sg13g2_inv_1 _12782_ (.Y(_04808_),
    .A(net2273));
 sg13g2_inv_1 _12783_ (.Y(_04809_),
    .A(net1650));
 sg13g2_inv_1 _12784_ (.Y(_04810_),
    .A(net2279));
 sg13g2_inv_1 _12785_ (.Y(_04811_),
    .A(net1795));
 sg13g2_inv_1 _12786_ (.Y(_04812_),
    .A(net2132));
 sg13g2_inv_1 _12787_ (.Y(_04813_),
    .A(\TRNG.Word_Out[432] ));
 sg13g2_inv_1 _12788_ (.Y(_04814_),
    .A(net2298));
 sg13g2_inv_1 _12789_ (.Y(_04815_),
    .A(net1913));
 sg13g2_inv_1 _12790_ (.Y(_04816_),
    .A(net1804));
 sg13g2_inv_1 _12791_ (.Y(_04817_),
    .A(net2346));
 sg13g2_inv_1 _12792_ (.Y(_04818_),
    .A(net2143));
 sg13g2_inv_1 _12793_ (.Y(_04819_),
    .A(net2026));
 sg13g2_inv_1 _12794_ (.Y(_04820_),
    .A(\TRNG.Word_Out[439] ));
 sg13g2_inv_1 _12795_ (.Y(_04821_),
    .A(net2514));
 sg13g2_inv_1 _12796_ (.Y(_04822_),
    .A(net2116));
 sg13g2_inv_1 _12797_ (.Y(_04823_),
    .A(\TRNG.Word_Out[442] ));
 sg13g2_inv_1 _12798_ (.Y(_04824_),
    .A(net2163));
 sg13g2_inv_1 _12799_ (.Y(_04825_),
    .A(net2316));
 sg13g2_inv_1 _12800_ (.Y(_04826_),
    .A(net2217));
 sg13g2_inv_1 _12801_ (.Y(_04827_),
    .A(net1130));
 sg13g2_inv_1 _12802_ (.Y(_04828_),
    .A(\TRNG.Word_Out[446] ));
 sg13g2_nor3_1 _12803_ (.A(net2679),
    .B(\TRNG.uart_tx_inst.currentState[1] ),
    .C(\TRNG.uart_tx_inst.currentState[0] ),
    .Y(_04829_));
 sg13g2_nand3b_1 _12804_ (.B(_04829_),
    .C(\TRNG.uart_tx_inst.currentState[2] ),
    .Y(_04830_),
    .A_N(\TRNG.uart_tx_inst.currentState[3] ));
 sg13g2_inv_1 _12805_ (.Y(_04831_),
    .A(_04830_));
 sg13g2_nor2_1 _12806_ (.A(\TRNG.uart_tx_inst.currentState[2] ),
    .B(\TRNG.uart_tx_inst.currentState[3] ),
    .Y(_04832_));
 sg13g2_nor3_1 _12807_ (.A(\TRNG.uart_tx_inst.currentState[0] ),
    .B(\TRNG.uart_tx_inst.currentState[2] ),
    .C(\TRNG.uart_tx_inst.currentState[3] ),
    .Y(_04833_));
 sg13g2_nand3_1 _12808_ (.B(net3291),
    .C(_04833_),
    .A(\TRNG.uart_tx_inst.currentState[1] ),
    .Y(_04834_));
 sg13g2_nand2_1 _12809_ (.Y(_04835_),
    .A(_04830_),
    .B(_04834_));
 sg13g2_nor2_1 _12810_ (.A(\TRNG.uart_tx_inst.tx_bit_counter[3] ),
    .B(\TRNG.uart_tx_inst.tx_reg[0] ),
    .Y(_04836_));
 sg13g2_o21ai_1 _12811_ (.B1(_04835_),
    .Y(\TRNG.UART_Tx ),
    .A1(_04830_),
    .A2(_04836_));
 sg13g2_nand2_1 _12812_ (.Y(_04837_),
    .A(\TRNG.state[1] ),
    .B(net3378));
 sg13g2_nand3_1 _12813_ (.B(\TRNG.state[0] ),
    .C(net3886),
    .A(\TRNG.state[1] ),
    .Y(_04838_));
 sg13g2_nor2b_1 _12814_ (.A(\TRNG.state[1] ),
    .B_N(_00119_),
    .Y(_04839_));
 sg13g2_and2_2 _12815_ (.A(_04305_),
    .B(_04839_),
    .X(_04840_));
 sg13g2_inv_1 _12816_ (.Y(_04841_),
    .A(_04840_));
 sg13g2_nand2b_1 _12817_ (.Y(_04842_),
    .B(_04840_),
    .A_N(net5517));
 sg13g2_o21ai_1 _12818_ (.B1(_04842_),
    .Y(_04843_),
    .A1(_04305_),
    .A2(\TRNG.state[2] ));
 sg13g2_and2_1 _12819_ (.A(_04838_),
    .B(_04843_),
    .X(_04844_));
 sg13g2_and2_2 _12820_ (.A(\TRNG.state[0] ),
    .B(_04839_),
    .X(_04845_));
 sg13g2_nand2_2 _12821_ (.Y(_04846_),
    .A(\TRNG.state[0] ),
    .B(_04839_));
 sg13g2_nand3b_1 _12822_ (.B(\TRNG.discard ),
    .C(net5237),
    .Y(_04847_),
    .A_N(\TRNG.Repetition_Count_Test.failure ));
 sg13g2_xnor2_1 _12823_ (.Y(_04848_),
    .A(net5517),
    .B(\TRNG.prev_ctrl_mode ));
 sg13g2_inv_2 _12824_ (.Y(_04849_),
    .A(net5457));
 sg13g2_a21oi_2 _12825_ (.B1(_04849_),
    .Y(_04850_),
    .A2(_04847_),
    .A1(_04844_));
 sg13g2_nor2_2 _12826_ (.A(\TRNG.Repetition_Count_Test.failure ),
    .B(net2936),
    .Y(_04851_));
 sg13g2_or2_2 _12827_ (.X(_04852_),
    .B(\TRNG.discard ),
    .A(\TRNG.Repetition_Count_Test.failure ));
 sg13g2_nor2_1 _12828_ (.A(_04846_),
    .B(_04852_),
    .Y(_04853_));
 sg13g2_nor3_2 _12829_ (.A(\TRNG.state[2] ),
    .B(_04846_),
    .C(_04852_),
    .Y(_04854_));
 sg13g2_a22oi_1 _12830_ (.Y(_04855_),
    .B1(_04854_),
    .B2(net1131),
    .A2(_04850_),
    .A1(\TRNG.bit_counter[0] ));
 sg13g2_inv_1 _12831_ (.Y(_02148_),
    .A(net1132));
 sg13g2_a21oi_1 _12832_ (.A1(\TRNG.bit_counter[0] ),
    .A2(_04854_),
    .Y(_04856_),
    .B1(net2331));
 sg13g2_nand2_1 _12833_ (.Y(_04857_),
    .A(net2331),
    .B(\TRNG.bit_counter[0] ));
 sg13g2_a21oi_1 _12834_ (.A1(net5100),
    .A2(_04857_),
    .Y(_04858_),
    .B1(_04850_));
 sg13g2_nor2_1 _12835_ (.A(net2332),
    .B(_04858_),
    .Y(_02149_));
 sg13g2_nand3_1 _12836_ (.B(\TRNG.bit_counter[0] ),
    .C(net3009),
    .A(net2331),
    .Y(_04859_));
 sg13g2_xnor2_1 _12837_ (.Y(_04860_),
    .A(net3009),
    .B(_04857_));
 sg13g2_a22oi_1 _12838_ (.Y(_04861_),
    .B1(net5100),
    .B2(_04860_),
    .A2(_04850_),
    .A1(net3009));
 sg13g2_inv_1 _12839_ (.Y(_02150_),
    .A(net3010));
 sg13g2_nor2_1 _12840_ (.A(_04307_),
    .B(_04859_),
    .Y(_04862_));
 sg13g2_xnor2_1 _12841_ (.Y(_04863_),
    .A(net3073),
    .B(_04859_));
 sg13g2_a22oi_1 _12842_ (.Y(_04864_),
    .B1(net5100),
    .B2(_04863_),
    .A2(_04850_),
    .A1(net3073));
 sg13g2_inv_1 _12843_ (.Y(_02151_),
    .A(net3074));
 sg13g2_nand2_1 _12844_ (.Y(_04865_),
    .A(net2329),
    .B(_04850_));
 sg13g2_and2_1 _12845_ (.A(net2329),
    .B(_04862_),
    .X(_04866_));
 sg13g2_o21ai_1 _12846_ (.B1(net5100),
    .Y(_04867_),
    .A1(net2329),
    .A2(_04862_));
 sg13g2_o21ai_1 _12847_ (.B1(_04865_),
    .Y(_02152_),
    .A1(_04866_),
    .A2(_04867_));
 sg13g2_nand2_1 _12848_ (.Y(_04868_),
    .A(net2361),
    .B(_04850_));
 sg13g2_and2_1 _12849_ (.A(net2361),
    .B(_04866_),
    .X(_04869_));
 sg13g2_o21ai_1 _12850_ (.B1(net5100),
    .Y(_04870_),
    .A1(net2361),
    .A2(_04866_));
 sg13g2_o21ai_1 _12851_ (.B1(_04868_),
    .Y(_02153_),
    .A1(_04869_),
    .A2(_04870_));
 sg13g2_nand2_1 _12852_ (.Y(_04871_),
    .A(net2754),
    .B(_04850_));
 sg13g2_and2_1 _12853_ (.A(net2754),
    .B(_04869_),
    .X(_04872_));
 sg13g2_o21ai_1 _12854_ (.B1(net5100),
    .Y(_04873_),
    .A1(net2754),
    .A2(_04869_));
 sg13g2_o21ai_1 _12855_ (.B1(_04871_),
    .Y(_02154_),
    .A1(_04872_),
    .A2(_04873_));
 sg13g2_xnor2_1 _12856_ (.Y(_04874_),
    .A(_04308_),
    .B(_04872_));
 sg13g2_a22oi_1 _12857_ (.Y(_04875_),
    .B1(net5100),
    .B2(_04874_),
    .A2(_04850_),
    .A1(net2557));
 sg13g2_inv_1 _12858_ (.Y(_02155_),
    .A(_04875_));
 sg13g2_nand3_1 _12859_ (.B(net2557),
    .C(_04872_),
    .A(_04306_),
    .Y(_04876_));
 sg13g2_nor4_1 _12860_ (.A(\TRNG.state[2] ),
    .B(\TRNG.Repetition_Count_Test.failure ),
    .C(_04846_),
    .D(_04849_),
    .Y(_04877_));
 sg13g2_xnor2_1 _12861_ (.Y(_04878_),
    .A(net2652),
    .B(_04876_));
 sg13g2_o21ai_1 _12862_ (.B1(_04878_),
    .Y(_04879_),
    .A1(net5100),
    .A2(_04877_));
 sg13g2_nand2_1 _12863_ (.Y(_04880_),
    .A(net2652),
    .B(net5457));
 sg13g2_o21ai_1 _12864_ (.B1(_04879_),
    .Y(_02156_),
    .A1(_04844_),
    .A2(_04880_));
 sg13g2_nand2_1 _12865_ (.Y(_04881_),
    .A(net3525),
    .B(_04848_));
 sg13g2_nor2b_2 _12866_ (.A(\TRNG.state[1] ),
    .B_N(\TRNG.state[2] ),
    .Y(_04882_));
 sg13g2_nand2_1 _12867_ (.Y(_04883_),
    .A(\TRNG.state[0] ),
    .B(_04882_));
 sg13g2_nand3b_1 _12868_ (.B(net3391),
    .C(_04829_),
    .Y(_04884_),
    .A_N(\TRNG.uart_tx_inst.currentState[2] ));
 sg13g2_nand3_1 _12869_ (.B(_04834_),
    .C(_04884_),
    .A(_04830_),
    .Y(_04885_));
 sg13g2_nand2_1 _12870_ (.Y(_04886_),
    .A(net2679),
    .B(_04833_));
 sg13g2_o21ai_1 _12871_ (.B1(net2670),
    .Y(_04887_),
    .A1(\TRNG.uart_tx_inst.currentState[1] ),
    .A2(_04886_));
 sg13g2_or2_1 _12872_ (.X(_04888_),
    .B(_04887_),
    .A(_04885_));
 sg13g2_inv_1 _12873_ (.Y(_04889_),
    .A(_04888_));
 sg13g2_nor2_1 _12874_ (.A(_04883_),
    .B(_04889_),
    .Y(_04890_));
 sg13g2_nand2_2 _12875_ (.Y(_04891_),
    .A(net1146),
    .B(_04840_));
 sg13g2_o21ai_1 _12876_ (.B1(_04891_),
    .Y(_04892_),
    .A1(_04840_),
    .A2(_04882_));
 sg13g2_nor2_1 _12877_ (.A(_04890_),
    .B(_04892_),
    .Y(_04893_));
 sg13g2_o21ai_1 _12878_ (.B1(_04306_),
    .Y(_04894_),
    .A1(_04840_),
    .A2(_04882_));
 sg13g2_nand2_1 _12879_ (.Y(_04895_),
    .A(_04881_),
    .B(_04894_));
 sg13g2_and2_1 _12880_ (.A(_04305_),
    .B(_04882_),
    .X(_04896_));
 sg13g2_nor2b_1 _12881_ (.A(net3449),
    .B_N(net5219),
    .Y(_04897_));
 sg13g2_nand2_1 _12882_ (.Y(_04898_),
    .A(_04306_),
    .B(net3525));
 sg13g2_nand3_1 _12883_ (.B(_04897_),
    .C(_04898_),
    .A(_04895_),
    .Y(_04899_));
 sg13g2_o21ai_1 _12884_ (.B1(_04899_),
    .Y(_02145_),
    .A1(_04881_),
    .A2(_04893_));
 sg13g2_nand2_1 _12885_ (.Y(_04900_),
    .A(net3400),
    .B(_04848_));
 sg13g2_nand3_1 _12886_ (.B(net3400),
    .C(net5457),
    .A(net2936),
    .Y(_04901_));
 sg13g2_nand2_1 _12887_ (.Y(_04902_),
    .A(\TRNG.raw_bit_counter[0] ),
    .B(\TRNG.raw_bit_counter[1] ));
 sg13g2_xnor2_1 _12888_ (.Y(_04903_),
    .A(\TRNG.raw_bit_counter[0] ),
    .B(net3400));
 sg13g2_o21ai_1 _12889_ (.B1(_04901_),
    .Y(_04904_),
    .A1(_04894_),
    .A2(_04903_));
 sg13g2_nand2_1 _12890_ (.Y(_04905_),
    .A(_04897_),
    .B(_04904_));
 sg13g2_o21ai_1 _12891_ (.B1(_04905_),
    .Y(_02146_),
    .A1(_04893_),
    .A2(net3401));
 sg13g2_nand2_1 _12892_ (.Y(_04906_),
    .A(net3314),
    .B(net5457));
 sg13g2_nand3_1 _12893_ (.B(net3314),
    .C(net5457),
    .A(net2936),
    .Y(_04907_));
 sg13g2_xor2_1 _12894_ (.B(_04902_),
    .A(net3314),
    .X(_04908_));
 sg13g2_o21ai_1 _12895_ (.B1(_04907_),
    .Y(_04909_),
    .A1(_04894_),
    .A2(_04908_));
 sg13g2_nand2_1 _12896_ (.Y(_04910_),
    .A(_04897_),
    .B(_04909_));
 sg13g2_o21ai_1 _12897_ (.B1(_04910_),
    .Y(_02147_),
    .A1(_04893_),
    .A2(_04906_));
 sg13g2_a21oi_1 _12898_ (.A1(net3041),
    .A2(net5458),
    .Y(_04911_),
    .B1(net2937));
 sg13g2_o21ai_1 _12899_ (.B1(net5218),
    .Y(_04912_),
    .A1(net2880),
    .A2(net5456));
 sg13g2_or2_1 _12900_ (.X(_04913_),
    .B(net5218),
    .A(_04840_));
 sg13g2_a21oi_2 _12901_ (.B1(_04849_),
    .Y(_04914_),
    .A2(_04913_),
    .A1(_04891_));
 sg13g2_nand2_1 _12902_ (.Y(_04915_),
    .A(net3041),
    .B(_04914_));
 sg13g2_o21ai_1 _12903_ (.B1(_04915_),
    .Y(_02160_),
    .A1(_04911_),
    .A2(_04912_));
 sg13g2_and2_2 _12904_ (.A(_04851_),
    .B(_04913_),
    .X(_04916_));
 sg13g2_a21oi_1 _12905_ (.A1(net3132),
    .A2(net5458),
    .Y(_04917_),
    .B1(_04916_));
 sg13g2_o21ai_1 _12906_ (.B1(net5219),
    .Y(_04918_),
    .A1(net3041),
    .A2(net5456));
 sg13g2_nand2_1 _12907_ (.Y(_04919_),
    .A(net3132),
    .B(_04914_));
 sg13g2_o21ai_1 _12908_ (.B1(_04919_),
    .Y(_02161_),
    .A1(_04917_),
    .A2(_04918_));
 sg13g2_a21oi_1 _12909_ (.A1(net2869),
    .A2(net5458),
    .Y(_04920_),
    .B1(_04916_));
 sg13g2_o21ai_1 _12910_ (.B1(net5218),
    .Y(_04921_),
    .A1(\TRNG.raw_byte[1] ),
    .A2(net5456));
 sg13g2_nand2_1 _12911_ (.Y(_04922_),
    .A(net2869),
    .B(_04914_));
 sg13g2_o21ai_1 _12912_ (.B1(_04922_),
    .Y(_02162_),
    .A1(_04920_),
    .A2(_04921_));
 sg13g2_a21oi_1 _12913_ (.A1(net2795),
    .A2(net5458),
    .Y(_04923_),
    .B1(_04916_));
 sg13g2_o21ai_1 _12914_ (.B1(net5218),
    .Y(_04924_),
    .A1(net2869),
    .A2(net5456));
 sg13g2_nand2_1 _12915_ (.Y(_04925_),
    .A(net2795),
    .B(_04914_));
 sg13g2_o21ai_1 _12916_ (.B1(_04925_),
    .Y(_02163_),
    .A1(_04923_),
    .A2(_04924_));
 sg13g2_a21oi_1 _12917_ (.A1(net2520),
    .A2(net5458),
    .Y(_04926_),
    .B1(_04916_));
 sg13g2_o21ai_1 _12918_ (.B1(net5218),
    .Y(_04927_),
    .A1(net2795),
    .A2(net5456));
 sg13g2_nand2_1 _12919_ (.Y(_04928_),
    .A(net2520),
    .B(_04914_));
 sg13g2_o21ai_1 _12920_ (.B1(_04928_),
    .Y(_02164_),
    .A1(_04926_),
    .A2(_04927_));
 sg13g2_a21oi_1 _12921_ (.A1(net2725),
    .A2(net5458),
    .Y(_04929_),
    .B1(_04916_));
 sg13g2_o21ai_1 _12922_ (.B1(net5218),
    .Y(_04930_),
    .A1(net2520),
    .A2(net5456));
 sg13g2_nand2_1 _12923_ (.Y(_04931_),
    .A(net2725),
    .B(_04914_));
 sg13g2_o21ai_1 _12924_ (.B1(_04931_),
    .Y(_02165_),
    .A1(_04929_),
    .A2(_04930_));
 sg13g2_a21oi_1 _12925_ (.A1(net3123),
    .A2(net5458),
    .Y(_04932_),
    .B1(_04916_));
 sg13g2_o21ai_1 _12926_ (.B1(net5218),
    .Y(_04933_),
    .A1(net2725),
    .A2(net5456));
 sg13g2_nand2_1 _12927_ (.Y(_04934_),
    .A(net3123),
    .B(_04914_));
 sg13g2_o21ai_1 _12928_ (.B1(_04934_),
    .Y(_02166_),
    .A1(_04932_),
    .A2(_04933_));
 sg13g2_a21oi_1 _12929_ (.A1(net2528),
    .A2(net5458),
    .Y(_04935_),
    .B1(_04916_));
 sg13g2_o21ai_1 _12930_ (.B1(net5218),
    .Y(_04936_),
    .A1(\TRNG.raw_byte[6] ),
    .A2(net5456));
 sg13g2_nand2_1 _12931_ (.Y(_04937_),
    .A(net2528),
    .B(_04914_));
 sg13g2_o21ai_1 _12932_ (.B1(_04937_),
    .Y(_02167_),
    .A1(_04935_),
    .A2(_04936_));
 sg13g2_and4_1 _12933_ (.A(\TRNG.raw_bit_counter[0] ),
    .B(\TRNG.raw_bit_counter[1] ),
    .C(\TRNG.raw_bit_counter[2] ),
    .D(net5219),
    .X(_04938_));
 sg13g2_a22oi_1 _12934_ (.Y(_04939_),
    .B1(_04851_),
    .B2(_04938_),
    .A2(net5457),
    .A1(\TRNG.state[0] ));
 sg13g2_nor4_1 _12935_ (.A(\TRNG.bit_counter[6] ),
    .B(_04308_),
    .C(_00120_),
    .D(_04852_),
    .Y(_04940_));
 sg13g2_and2_1 _12936_ (.A(_04869_),
    .B(_04940_),
    .X(_04941_));
 sg13g2_nor2_1 _12937_ (.A(_04846_),
    .B(_04941_),
    .Y(_04942_));
 sg13g2_nor3_1 _12938_ (.A(_04890_),
    .B(_04938_),
    .C(_04942_),
    .Y(_04943_));
 sg13g2_nor2_1 _12939_ (.A(_04939_),
    .B(_04943_),
    .Y(_04944_));
 sg13g2_nand4_1 _12940_ (.B(\TRNG.state[1] ),
    .C(_04305_),
    .A(net2873),
    .Y(_04945_),
    .D(net3378));
 sg13g2_inv_1 _12941_ (.Y(_04946_),
    .A(_04945_));
 sg13g2_nand2b_1 _12942_ (.Y(_04947_),
    .B(net5457),
    .A_N(_04837_));
 sg13g2_o21ai_1 _12943_ (.B1(_04842_),
    .Y(_04948_),
    .A1(_04838_),
    .A2(_04849_));
 sg13g2_or3_1 _12944_ (.A(_04944_),
    .B(_04946_),
    .C(_04948_),
    .X(_02157_));
 sg13g2_nand2_2 _12945_ (.Y(_04949_),
    .A(net5237),
    .B(_04941_));
 sg13g2_nand3_1 _12946_ (.B(_04947_),
    .C(net4606),
    .A(net3379),
    .Y(_02158_));
 sg13g2_a21oi_1 _12947_ (.A1(\TRNG.hash_rdy ),
    .A2(_04305_),
    .Y(_04950_),
    .B1(_04837_));
 sg13g2_a22oi_1 _12948_ (.Y(_04951_),
    .B1(_04851_),
    .B2(_04938_),
    .A2(net5457),
    .A1(\TRNG.state[2] ));
 sg13g2_o21ai_1 _12949_ (.B1(_04951_),
    .Y(_04952_),
    .A1(_04883_),
    .A2(_04888_));
 sg13g2_o21ai_1 _12950_ (.B1(_04952_),
    .Y(_04953_),
    .A1(_04882_),
    .A2(_04950_));
 sg13g2_o21ai_1 _12951_ (.B1(_04953_),
    .Y(_02159_),
    .A1(net1146),
    .A2(_04841_));
 sg13g2_nand2_1 _12952_ (.Y(_04954_),
    .A(_04277_),
    .B(\TRNG.sha256.expand.address1[2] ));
 sg13g2_nor2b_1 _12953_ (.A(\TRNG.sha256.expand.address1[1] ),
    .B_N(\TRNG.sha256.expand.address1[0] ),
    .Y(_04955_));
 sg13g2_nor2b_1 _12954_ (.A(\TRNG.sha256.expand.address1[0] ),
    .B_N(\TRNG.sha256.expand.address1[1] ),
    .Y(_04956_));
 sg13g2_a22oi_1 _12955_ (.Y(_04957_),
    .B1(net5412),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][0] ),
    .A2(net5434),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][0] ));
 sg13g2_nor2_2 _12956_ (.A(\TRNG.sha256.expand.address1[1] ),
    .B(\TRNG.sha256.expand.address1[0] ),
    .Y(_04958_));
 sg13g2_and2_1 _12957_ (.A(\TRNG.sha256.expand.address1[1] ),
    .B(\TRNG.sha256.expand.address1[0] ),
    .X(_04959_));
 sg13g2_a22oi_1 _12958_ (.Y(_04960_),
    .B1(net5365),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][0] ),
    .A2(net5388),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][0] ));
 sg13g2_a21oi_1 _12959_ (.A1(_04957_),
    .A2(_04960_),
    .Y(_04961_),
    .B1(net5214));
 sg13g2_nand2_1 _12960_ (.Y(_04962_),
    .A(\TRNG.sha256.expand.address1[3] ),
    .B(_04278_));
 sg13g2_a22oi_1 _12961_ (.Y(_04963_),
    .B1(net5412),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][0] ),
    .A2(net5434),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][0] ));
 sg13g2_a22oi_1 _12962_ (.Y(_04964_),
    .B1(net5365),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][0] ),
    .A2(net5388),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][0] ));
 sg13g2_a21oi_1 _12963_ (.A1(_04963_),
    .A2(_04964_),
    .Y(_04965_),
    .B1(net5208));
 sg13g2_nand2_1 _12964_ (.Y(_04966_),
    .A(_04277_),
    .B(_04278_));
 sg13g2_a22oi_1 _12965_ (.Y(_04967_),
    .B1(net5412),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][0] ),
    .A2(net5434),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][0] ));
 sg13g2_a22oi_1 _12966_ (.Y(_04968_),
    .B1(net5365),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][0] ),
    .A2(net5388),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][0] ));
 sg13g2_a21oi_1 _12967_ (.A1(_04967_),
    .A2(_04968_),
    .Y(_04969_),
    .B1(net5203));
 sg13g2_nand2_1 _12968_ (.Y(_04970_),
    .A(\TRNG.sha256.expand.address1[3] ),
    .B(\TRNG.sha256.expand.address1[2] ));
 sg13g2_a22oi_1 _12969_ (.Y(_04971_),
    .B1(net5412),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][0] ),
    .A2(net5434),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][0] ));
 sg13g2_a22oi_1 _12970_ (.Y(_04972_),
    .B1(net5365),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][0] ),
    .A2(net5388),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][0] ));
 sg13g2_a21oi_1 _12971_ (.A1(_04971_),
    .A2(_04972_),
    .Y(_04973_),
    .B1(net5361));
 sg13g2_or4_2 _12972_ (.A(_04961_),
    .B(_04965_),
    .C(_04969_),
    .D(_04973_),
    .X(_00064_));
 sg13g2_a22oi_1 _12973_ (.Y(_04974_),
    .B1(net5414),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][1] ),
    .A2(net5436),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][1] ));
 sg13g2_a22oi_1 _12974_ (.Y(_04975_),
    .B1(net5367),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][1] ),
    .A2(net5390),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][1] ));
 sg13g2_a21oi_1 _12975_ (.A1(_04974_),
    .A2(_04975_),
    .Y(_04976_),
    .B1(net5214));
 sg13g2_a22oi_1 _12976_ (.Y(_04977_),
    .B1(net5414),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][1] ),
    .A2(net5436),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][1] ));
 sg13g2_a22oi_1 _12977_ (.Y(_04978_),
    .B1(net5367),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][1] ),
    .A2(net5390),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][1] ));
 sg13g2_a21oi_1 _12978_ (.A1(_04977_),
    .A2(_04978_),
    .Y(_04979_),
    .B1(net5361));
 sg13g2_a22oi_1 _12979_ (.Y(_04980_),
    .B1(net5414),
    .B2(net2723),
    .A2(net5436),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][1] ));
 sg13g2_a22oi_1 _12980_ (.Y(_04981_),
    .B1(net5367),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][1] ),
    .A2(net5390),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][1] ));
 sg13g2_a21oi_1 _12981_ (.A1(_04980_),
    .A2(_04981_),
    .Y(_04982_),
    .B1(net5203));
 sg13g2_a22oi_1 _12982_ (.Y(_04983_),
    .B1(net5414),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][1] ),
    .A2(net5436),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][1] ));
 sg13g2_a22oi_1 _12983_ (.Y(_04984_),
    .B1(net5367),
    .B2(net3915),
    .A2(net5390),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][1] ));
 sg13g2_a21oi_1 _12984_ (.A1(_04983_),
    .A2(_04984_),
    .Y(_04985_),
    .B1(net5208));
 sg13g2_or4_1 _12985_ (.A(_04976_),
    .B(_04979_),
    .C(_04982_),
    .D(net3916),
    .X(_00075_));
 sg13g2_a22oi_1 _12986_ (.Y(_04986_),
    .B1(net5418),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][2] ),
    .A2(net5440),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][2] ));
 sg13g2_a22oi_1 _12987_ (.Y(_04987_),
    .B1(net5371),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][2] ),
    .A2(net5395),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][2] ));
 sg13g2_a21oi_1 _12988_ (.A1(_04986_),
    .A2(_04987_),
    .Y(_04988_),
    .B1(net5202));
 sg13g2_a22oi_1 _12989_ (.Y(_04989_),
    .B1(net5418),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][2] ),
    .A2(net5440),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][2] ));
 sg13g2_a22oi_1 _12990_ (.Y(_04990_),
    .B1(net5371),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][2] ),
    .A2(net5395),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][2] ));
 sg13g2_a21oi_1 _12991_ (.A1(_04989_),
    .A2(_04990_),
    .Y(_04991_),
    .B1(net5360));
 sg13g2_a22oi_1 _12992_ (.Y(_04992_),
    .B1(net5418),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][2] ),
    .A2(net5440),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][2] ));
 sg13g2_a22oi_1 _12993_ (.Y(_04993_),
    .B1(net5371),
    .B2(net3936),
    .A2(net5395),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][2] ));
 sg13g2_a21oi_1 _12994_ (.A1(_04992_),
    .A2(_04993_),
    .Y(_04994_),
    .B1(net5213));
 sg13g2_a22oi_1 _12995_ (.Y(_04995_),
    .B1(net5418),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][2] ),
    .A2(net5440),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][2] ));
 sg13g2_a22oi_1 _12996_ (.Y(_04996_),
    .B1(net5371),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][2] ),
    .A2(net5395),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][2] ));
 sg13g2_a21oi_1 _12997_ (.A1(_04995_),
    .A2(_04996_),
    .Y(_04997_),
    .B1(net5207));
 sg13g2_or4_2 _12998_ (.A(_04988_),
    .B(_04991_),
    .C(_04994_),
    .D(_04997_),
    .X(_00086_));
 sg13g2_a22oi_1 _12999_ (.Y(_04998_),
    .B1(net5425),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][3] ),
    .A2(net5447),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][3] ));
 sg13g2_a22oi_1 _13000_ (.Y(_04999_),
    .B1(net5378),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][3] ),
    .A2(net5403),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][3] ));
 sg13g2_a21oi_1 _13001_ (.A1(_04998_),
    .A2(_04999_),
    .Y(_05000_),
    .B1(net5205));
 sg13g2_a22oi_1 _13002_ (.Y(_05001_),
    .B1(net5423),
    .B2(net3920),
    .A2(net5445),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][3] ));
 sg13g2_a22oi_1 _13003_ (.Y(_05002_),
    .B1(net5376),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][3] ),
    .A2(net5400),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][3] ));
 sg13g2_a21oi_1 _13004_ (.A1(_05001_),
    .A2(_05002_),
    .Y(_05003_),
    .B1(net5363));
 sg13g2_a22oi_1 _13005_ (.Y(_05004_),
    .B1(net5425),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][3] ),
    .A2(net5447),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][3] ));
 sg13g2_a22oi_1 _13006_ (.Y(_05005_),
    .B1(net5378),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][3] ),
    .A2(net5403),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][3] ));
 sg13g2_a21oi_1 _13007_ (.A1(_05004_),
    .A2(_05005_),
    .Y(_05006_),
    .B1(net5215));
 sg13g2_a22oi_1 _13008_ (.Y(_05007_),
    .B1(net5425),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][3] ),
    .A2(net5447),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][3] ));
 sg13g2_a22oi_1 _13009_ (.Y(_05008_),
    .B1(net5378),
    .B2(net2974),
    .A2(net5403),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][3] ));
 sg13g2_a21oi_1 _13010_ (.A1(_05007_),
    .A2(_05008_),
    .Y(_05009_),
    .B1(net5209));
 sg13g2_or4_1 _13011_ (.A(_05000_),
    .B(_05003_),
    .C(_05006_),
    .D(_05009_),
    .X(_00089_));
 sg13g2_a22oi_1 _13012_ (.Y(_05010_),
    .B1(net5421),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][4] ),
    .A2(net5443),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][4] ));
 sg13g2_a22oi_1 _13013_ (.Y(_05011_),
    .B1(net5374),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][4] ),
    .A2(net5394),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][4] ));
 sg13g2_a21oi_1 _13014_ (.A1(_05010_),
    .A2(_05011_),
    .Y(_05012_),
    .B1(net5202));
 sg13g2_a22oi_1 _13015_ (.Y(_05013_),
    .B1(net5417),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][4] ),
    .A2(net5439),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][4] ));
 sg13g2_a22oi_1 _13016_ (.Y(_05014_),
    .B1(net5370),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][4] ),
    .A2(net5393),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][4] ));
 sg13g2_a21oi_1 _13017_ (.A1(_05013_),
    .A2(_05014_),
    .Y(_05015_),
    .B1(net5207));
 sg13g2_a22oi_1 _13018_ (.Y(_05016_),
    .B1(net5417),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][4] ),
    .A2(net5439),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][4] ));
 sg13g2_a22oi_1 _13019_ (.Y(_05017_),
    .B1(net5370),
    .B2(net3932),
    .A2(net5394),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][4] ));
 sg13g2_a21oi_1 _13020_ (.A1(_05016_),
    .A2(_05017_),
    .Y(_05018_),
    .B1(net5213));
 sg13g2_a22oi_1 _13021_ (.Y(_05019_),
    .B1(net5417),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][4] ),
    .A2(net5439),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][4] ));
 sg13g2_a22oi_1 _13022_ (.Y(_05020_),
    .B1(net5370),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][4] ),
    .A2(net5393),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][4] ));
 sg13g2_a21oi_1 _13023_ (.A1(_05019_),
    .A2(_05020_),
    .Y(_05021_),
    .B1(net5360));
 sg13g2_or4_2 _13024_ (.A(_05012_),
    .B(_05015_),
    .C(_05018_),
    .D(_05021_),
    .X(_00090_));
 sg13g2_a22oi_1 _13025_ (.Y(_05022_),
    .B1(net5419),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][5] ),
    .A2(net5441),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][5] ));
 sg13g2_a22oi_1 _13026_ (.Y(_05023_),
    .B1(net5372),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][5] ),
    .A2(net5396),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][5] ));
 sg13g2_a21oi_1 _13027_ (.A1(_05022_),
    .A2(_05023_),
    .Y(_05024_),
    .B1(net5202));
 sg13g2_a22oi_1 _13028_ (.Y(_05025_),
    .B1(net5419),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][5] ),
    .A2(net5441),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][5] ));
 sg13g2_a22oi_1 _13029_ (.Y(_05026_),
    .B1(net5372),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][5] ),
    .A2(net5396),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][5] ));
 sg13g2_a21oi_1 _13030_ (.A1(_05025_),
    .A2(_05026_),
    .Y(_05027_),
    .B1(net5207));
 sg13g2_a22oi_1 _13031_ (.Y(_05028_),
    .B1(net5420),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][5] ),
    .A2(net5442),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][5] ));
 sg13g2_a22oi_1 _13032_ (.Y(_05029_),
    .B1(net5373),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][5] ),
    .A2(net5397),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][5] ));
 sg13g2_a21oi_1 _13033_ (.A1(_05028_),
    .A2(_05029_),
    .Y(_05030_),
    .B1(net5213));
 sg13g2_a22oi_1 _13034_ (.Y(_05031_),
    .B1(net5417),
    .B2(net3909),
    .A2(net5439),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][5] ));
 sg13g2_a22oi_1 _13035_ (.Y(_05032_),
    .B1(net5370),
    .B2(net3071),
    .A2(net5396),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][5] ));
 sg13g2_a21oi_1 _13036_ (.A1(_05031_),
    .A2(_05032_),
    .Y(_05033_),
    .B1(net5360));
 sg13g2_or4_1 _13037_ (.A(_05024_),
    .B(_05027_),
    .C(_05030_),
    .D(_05033_),
    .X(_00091_));
 sg13g2_a22oi_1 _13038_ (.Y(_05034_),
    .B1(net5421),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][6] ),
    .A2(net5443),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][6] ));
 sg13g2_a22oi_1 _13039_ (.Y(_05035_),
    .B1(net5374),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][6] ),
    .A2(net5393),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][6] ));
 sg13g2_a21oi_1 _13040_ (.A1(_05034_),
    .A2(_05035_),
    .Y(_05036_),
    .B1(net5213));
 sg13g2_a22oi_1 _13041_ (.Y(_05037_),
    .B1(net5417),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][6] ),
    .A2(net5439),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][6] ));
 sg13g2_a22oi_1 _13042_ (.Y(_05038_),
    .B1(net5370),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][6] ),
    .A2(net5394),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][6] ));
 sg13g2_a21oi_1 _13043_ (.A1(_05037_),
    .A2(_05038_),
    .Y(_05039_),
    .B1(net5207));
 sg13g2_a22oi_1 _13044_ (.Y(_05040_),
    .B1(net5417),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][6] ),
    .A2(net5439),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][6] ));
 sg13g2_a22oi_1 _13045_ (.Y(_05041_),
    .B1(net5370),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][6] ),
    .A2(net5393),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][6] ));
 sg13g2_a21oi_1 _13046_ (.A1(_05040_),
    .A2(_05041_),
    .Y(_05042_),
    .B1(net5202));
 sg13g2_a22oi_1 _13047_ (.Y(_05043_),
    .B1(net5417),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][6] ),
    .A2(net5439),
    .A1(net3902));
 sg13g2_a22oi_1 _13048_ (.Y(_05044_),
    .B1(net5370),
    .B2(net3175),
    .A2(net5394),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][6] ));
 sg13g2_a21oi_1 _13049_ (.A1(net3903),
    .A2(_05044_),
    .Y(_05045_),
    .B1(net5360));
 sg13g2_or4_1 _13050_ (.A(_05036_),
    .B(_05039_),
    .C(_05042_),
    .D(net3904),
    .X(_00092_));
 sg13g2_a22oi_1 _13051_ (.Y(_05046_),
    .B1(net5427),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][7] ),
    .A2(net5449),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][7] ));
 sg13g2_a22oi_1 _13052_ (.Y(_05047_),
    .B1(net5380),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][7] ),
    .A2(net5406),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][7] ));
 sg13g2_a21oi_1 _13053_ (.A1(_05046_),
    .A2(_05047_),
    .Y(_05048_),
    .B1(net5206));
 sg13g2_a22oi_1 _13054_ (.Y(_05049_),
    .B1(net5427),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][7] ),
    .A2(net5449),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][7] ));
 sg13g2_a22oi_1 _13055_ (.Y(_05050_),
    .B1(net5380),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][7] ),
    .A2(net5406),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][7] ));
 sg13g2_a21oi_1 _13056_ (.A1(_05049_),
    .A2(_05050_),
    .Y(_05051_),
    .B1(net5210));
 sg13g2_a22oi_1 _13057_ (.Y(_05052_),
    .B1(net5427),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][7] ),
    .A2(net5449),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][7] ));
 sg13g2_a22oi_1 _13058_ (.Y(_05053_),
    .B1(net5380),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][7] ),
    .A2(net5405),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][7] ));
 sg13g2_a21oi_1 _13059_ (.A1(_05052_),
    .A2(_05053_),
    .Y(_05054_),
    .B1(net5216));
 sg13g2_a22oi_1 _13060_ (.Y(_05055_),
    .B1(net5427),
    .B2(net3907),
    .A2(net5449),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][7] ));
 sg13g2_a22oi_1 _13061_ (.Y(_05056_),
    .B1(net5381),
    .B2(net2950),
    .A2(net5406),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][7] ));
 sg13g2_a21oi_1 _13062_ (.A1(_05055_),
    .A2(_05056_),
    .Y(_05057_),
    .B1(net5362));
 sg13g2_or4_2 _13063_ (.A(_05048_),
    .B(_05051_),
    .C(_05054_),
    .D(_05057_),
    .X(_00093_));
 sg13g2_a22oi_1 _13064_ (.Y(_05058_),
    .B1(net5419),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][8] ),
    .A2(net5441),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][8] ));
 sg13g2_a22oi_1 _13065_ (.Y(_05059_),
    .B1(net5372),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][8] ),
    .A2(net5397),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][8] ));
 sg13g2_a21oi_1 _13066_ (.A1(_05058_),
    .A2(_05059_),
    .Y(_05060_),
    .B1(net5206));
 sg13g2_a22oi_1 _13067_ (.Y(_05061_),
    .B1(net5420),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][8] ),
    .A2(net5442),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][8] ));
 sg13g2_a22oi_1 _13068_ (.Y(_05062_),
    .B1(net5373),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][8] ),
    .A2(net5397),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][8] ));
 sg13g2_a21oi_1 _13069_ (.A1(_05061_),
    .A2(_05062_),
    .Y(_05063_),
    .B1(net5364));
 sg13g2_a22oi_1 _13070_ (.Y(_05064_),
    .B1(net5420),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][8] ),
    .A2(net5442),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][8] ));
 sg13g2_a22oi_1 _13071_ (.Y(_05065_),
    .B1(net5373),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][8] ),
    .A2(net5396),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][8] ));
 sg13g2_a21oi_1 _13072_ (.A1(_05064_),
    .A2(_05065_),
    .Y(_05066_),
    .B1(net5217));
 sg13g2_a22oi_1 _13073_ (.Y(_05067_),
    .B1(net5419),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][8] ),
    .A2(net5441),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][8] ));
 sg13g2_a22oi_1 _13074_ (.Y(_05068_),
    .B1(net5372),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][8] ),
    .A2(net5397),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][8] ));
 sg13g2_a21oi_1 _13075_ (.A1(_05067_),
    .A2(_05068_),
    .Y(_05069_),
    .B1(net5212));
 sg13g2_or4_1 _13076_ (.A(_05060_),
    .B(_05063_),
    .C(_05066_),
    .D(_05069_),
    .X(_00094_));
 sg13g2_a22oi_1 _13077_ (.Y(_05070_),
    .B1(net5430),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][9] ),
    .A2(net5452),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][9] ));
 sg13g2_a22oi_1 _13078_ (.Y(_05071_),
    .B1(net5383),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][9] ),
    .A2(net5408),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][9] ));
 sg13g2_a21oi_1 _13079_ (.A1(_05070_),
    .A2(_05071_),
    .Y(_05072_),
    .B1(net5217));
 sg13g2_a22oi_1 _13080_ (.Y(_05073_),
    .B1(net5429),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][9] ),
    .A2(net5451),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][9] ));
 sg13g2_a22oi_1 _13081_ (.Y(_05074_),
    .B1(net5382),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][9] ),
    .A2(net5407),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][9] ));
 sg13g2_a21oi_1 _13082_ (.A1(_05073_),
    .A2(_05074_),
    .Y(_05075_),
    .B1(net5362));
 sg13g2_a22oi_1 _13083_ (.Y(_05076_),
    .B1(net5427),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][9] ),
    .A2(net5449),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][9] ));
 sg13g2_a22oi_1 _13084_ (.Y(_05077_),
    .B1(net5383),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][9] ),
    .A2(net5408),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][9] ));
 sg13g2_a21oi_1 _13085_ (.A1(_05076_),
    .A2(_05077_),
    .Y(_05078_),
    .B1(net5205));
 sg13g2_a22oi_1 _13086_ (.Y(_05079_),
    .B1(net5428),
    .B2(net2866),
    .A2(net5450),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][9] ));
 sg13g2_a22oi_1 _13087_ (.Y(_05080_),
    .B1(net5382),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][9] ),
    .A2(net5407),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][9] ));
 sg13g2_a21oi_1 _13088_ (.A1(_05079_),
    .A2(_05080_),
    .Y(_05081_),
    .B1(net5210));
 sg13g2_or4_1 _13089_ (.A(_05072_),
    .B(_05075_),
    .C(_05078_),
    .D(_05081_),
    .X(_00095_));
 sg13g2_a22oi_1 _13090_ (.Y(_05082_),
    .B1(net5429),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][10] ),
    .A2(net5451),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][10] ));
 sg13g2_a22oi_1 _13091_ (.Y(_05083_),
    .B1(net5382),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][10] ),
    .A2(net5410),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][10] ));
 sg13g2_a21oi_1 _13092_ (.A1(_05082_),
    .A2(_05083_),
    .Y(_05084_),
    .B1(net5217));
 sg13g2_a22oi_1 _13093_ (.Y(_05085_),
    .B1(net5429),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][10] ),
    .A2(net5451),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][10] ));
 sg13g2_a22oi_1 _13094_ (.Y(_05086_),
    .B1(net5382),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][10] ),
    .A2(net5407),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][10] ));
 sg13g2_a21oi_1 _13095_ (.A1(_05085_),
    .A2(_05086_),
    .Y(_05087_),
    .B1(net5362));
 sg13g2_a22oi_1 _13096_ (.Y(_05088_),
    .B1(net5429),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][10] ),
    .A2(net5451),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][10] ));
 sg13g2_a22oi_1 _13097_ (.Y(_05089_),
    .B1(net5382),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][10] ),
    .A2(net5407),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][10] ));
 sg13g2_a21oi_1 _13098_ (.A1(_05088_),
    .A2(_05089_),
    .Y(_05090_),
    .B1(net5205));
 sg13g2_a22oi_1 _13099_ (.Y(_05091_),
    .B1(net5429),
    .B2(net3931),
    .A2(net5451),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][10] ));
 sg13g2_a22oi_1 _13100_ (.Y(_05092_),
    .B1(net5382),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][10] ),
    .A2(net5407),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][10] ));
 sg13g2_a21oi_1 _13101_ (.A1(_05091_),
    .A2(_05092_),
    .Y(_05093_),
    .B1(net5211));
 sg13g2_or4_1 _13102_ (.A(_05084_),
    .B(_05087_),
    .C(_05090_),
    .D(_05093_),
    .X(_00065_));
 sg13g2_a22oi_1 _13103_ (.Y(_05094_),
    .B1(net5415),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][11] ),
    .A2(net5437),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][11] ));
 sg13g2_a22oi_1 _13104_ (.Y(_05095_),
    .B1(net5368),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][11] ),
    .A2(net5391),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][11] ));
 sg13g2_a21oi_1 _13105_ (.A1(_05094_),
    .A2(_05095_),
    .Y(_05096_),
    .B1(net5214));
 sg13g2_a22oi_1 _13106_ (.Y(_05097_),
    .B1(net5415),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][11] ),
    .A2(net5437),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][11] ));
 sg13g2_a22oi_1 _13107_ (.Y(_05098_),
    .B1(net5368),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][11] ),
    .A2(net5391),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][11] ));
 sg13g2_a21oi_1 _13108_ (.A1(_05097_),
    .A2(_05098_),
    .Y(_05099_),
    .B1(net5208));
 sg13g2_a22oi_1 _13109_ (.Y(_05100_),
    .B1(net5415),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][11] ),
    .A2(net5437),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][11] ));
 sg13g2_a22oi_1 _13110_ (.Y(_05101_),
    .B1(net5368),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][11] ),
    .A2(net5391),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][11] ));
 sg13g2_a21oi_1 _13111_ (.A1(_05100_),
    .A2(_05101_),
    .Y(_05102_),
    .B1(net5203));
 sg13g2_a22oi_1 _13112_ (.Y(_05103_),
    .B1(net5415),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][11] ),
    .A2(net5437),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][11] ));
 sg13g2_a22oi_1 _13113_ (.Y(_05104_),
    .B1(net5368),
    .B2(net3935),
    .A2(net5391),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][11] ));
 sg13g2_a21oi_1 _13114_ (.A1(_05103_),
    .A2(_05104_),
    .Y(_05105_),
    .B1(net5361));
 sg13g2_or4_1 _13115_ (.A(_05096_),
    .B(_05099_),
    .C(_05102_),
    .D(_05105_),
    .X(_00066_));
 sg13g2_a22oi_1 _13116_ (.Y(_05106_),
    .B1(net5413),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][12] ),
    .A2(net5435),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][12] ));
 sg13g2_a22oi_1 _13117_ (.Y(_05107_),
    .B1(net5366),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][12] ),
    .A2(net5389),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][12] ));
 sg13g2_a21oi_1 _13118_ (.A1(_05106_),
    .A2(_05107_),
    .Y(_05108_),
    .B1(net5203));
 sg13g2_a22oi_1 _13119_ (.Y(_05109_),
    .B1(net5413),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][12] ),
    .A2(net5435),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][12] ));
 sg13g2_a22oi_1 _13120_ (.Y(_05110_),
    .B1(net5366),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][12] ),
    .A2(net5389),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][12] ));
 sg13g2_a21oi_1 _13121_ (.A1(_05109_),
    .A2(_05110_),
    .Y(_05111_),
    .B1(net5208));
 sg13g2_a22oi_1 _13122_ (.Y(_05112_),
    .B1(net5413),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][12] ),
    .A2(net5435),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][12] ));
 sg13g2_a22oi_1 _13123_ (.Y(_05113_),
    .B1(net5366),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][12] ),
    .A2(net5389),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][12] ));
 sg13g2_a21oi_1 _13124_ (.A1(_05112_),
    .A2(_05113_),
    .Y(_05114_),
    .B1(net5214));
 sg13g2_a22oi_1 _13125_ (.Y(_05115_),
    .B1(net5413),
    .B2(net3896),
    .A2(net5435),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][12] ));
 sg13g2_a22oi_1 _13126_ (.Y(_05116_),
    .B1(net5366),
    .B2(net2912),
    .A2(net5389),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][12] ));
 sg13g2_a21oi_1 _13127_ (.A1(_05115_),
    .A2(_05116_),
    .Y(_05117_),
    .B1(net5361));
 sg13g2_or4_2 _13128_ (.A(_05108_),
    .B(_05111_),
    .C(_05114_),
    .D(_05117_),
    .X(_00067_));
 sg13g2_a22oi_1 _13129_ (.Y(_05118_),
    .B1(net5412),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][13] ),
    .A2(net5434),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][13] ));
 sg13g2_a22oi_1 _13130_ (.Y(_05119_),
    .B1(net5365),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][13] ),
    .A2(net5388),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][13] ));
 sg13g2_a21oi_1 _13131_ (.A1(_05118_),
    .A2(_05119_),
    .Y(_05120_),
    .B1(net5214));
 sg13g2_a22oi_1 _13132_ (.Y(_05121_),
    .B1(net5412),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][13] ),
    .A2(net5434),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][13] ));
 sg13g2_a22oi_1 _13133_ (.Y(_05122_),
    .B1(net5365),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][13] ),
    .A2(net5388),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][13] ));
 sg13g2_a21oi_1 _13134_ (.A1(_05121_),
    .A2(_05122_),
    .Y(_05123_),
    .B1(net5361));
 sg13g2_a22oi_1 _13135_ (.Y(_05124_),
    .B1(net5412),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][13] ),
    .A2(net5434),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][13] ));
 sg13g2_a22oi_1 _13136_ (.Y(_05125_),
    .B1(net5365),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][13] ),
    .A2(net5388),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][13] ));
 sg13g2_a21oi_1 _13137_ (.A1(_05124_),
    .A2(_05125_),
    .Y(_05126_),
    .B1(net5203));
 sg13g2_a22oi_1 _13138_ (.Y(_05127_),
    .B1(net5412),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][13] ),
    .A2(net5434),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][13] ));
 sg13g2_a22oi_1 _13139_ (.Y(_05128_),
    .B1(net5365),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][13] ),
    .A2(net5388),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][13] ));
 sg13g2_a21oi_1 _13140_ (.A1(_05127_),
    .A2(_05128_),
    .Y(_05129_),
    .B1(net5208));
 sg13g2_or4_2 _13141_ (.A(_05120_),
    .B(_05123_),
    .C(_05126_),
    .D(_05129_),
    .X(_00068_));
 sg13g2_a22oi_1 _13142_ (.Y(_05130_),
    .B1(net5430),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][14] ),
    .A2(net5452),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][14] ));
 sg13g2_a22oi_1 _13143_ (.Y(_05131_),
    .B1(net5383),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][14] ),
    .A2(net5409),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][14] ));
 sg13g2_a21oi_1 _13144_ (.A1(_05130_),
    .A2(_05131_),
    .Y(_05132_),
    .B1(net5205));
 sg13g2_a22oi_1 _13145_ (.Y(_05133_),
    .B1(net5431),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][14] ),
    .A2(net5453),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][14] ));
 sg13g2_a22oi_1 _13146_ (.Y(_05134_),
    .B1(net5384),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][14] ),
    .A2(net5409),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][14] ));
 sg13g2_a21oi_1 _13147_ (.A1(_05133_),
    .A2(_05134_),
    .Y(_05135_),
    .B1(net5362));
 sg13g2_a22oi_1 _13148_ (.Y(_05136_),
    .B1(net5431),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][14] ),
    .A2(net5453),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][14] ));
 sg13g2_a22oi_1 _13149_ (.Y(_05137_),
    .B1(net5384),
    .B2(net3047),
    .A2(net5409),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][14] ));
 sg13g2_a21oi_1 _13150_ (.A1(_05136_),
    .A2(_05137_),
    .Y(_05138_),
    .B1(net5216));
 sg13g2_a22oi_1 _13151_ (.Y(_05139_),
    .B1(net5431),
    .B2(net3910),
    .A2(net5453),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][14] ));
 sg13g2_a22oi_1 _13152_ (.Y(_05140_),
    .B1(net5384),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][14] ),
    .A2(net5409),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][14] ));
 sg13g2_a21oi_1 _13153_ (.A1(net3911),
    .A2(_05140_),
    .Y(_05141_),
    .B1(net5210));
 sg13g2_or4_1 _13154_ (.A(_05132_),
    .B(_05135_),
    .C(_05138_),
    .D(_05141_),
    .X(_00069_));
 sg13g2_a22oi_1 _13155_ (.Y(_05142_),
    .B1(net5422),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][15] ),
    .A2(net5444),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][15] ));
 sg13g2_a22oi_1 _13156_ (.Y(_05143_),
    .B1(net5368),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][15] ),
    .A2(net5399),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][15] ));
 sg13g2_a21oi_1 _13157_ (.A1(_05142_),
    .A2(_05143_),
    .Y(_05144_),
    .B1(net5215));
 sg13g2_a22oi_1 _13158_ (.Y(_05145_),
    .B1(net5415),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][15] ),
    .A2(net5437),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][15] ));
 sg13g2_a22oi_1 _13159_ (.Y(_05146_),
    .B1(net5375),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][15] ),
    .A2(net5399),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][15] ));
 sg13g2_a21oi_1 _13160_ (.A1(_05145_),
    .A2(_05146_),
    .Y(_05147_),
    .B1(net5361));
 sg13g2_a22oi_1 _13161_ (.Y(_05148_),
    .B1(net5415),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][15] ),
    .A2(net5437),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][15] ));
 sg13g2_a22oi_1 _13162_ (.Y(_05149_),
    .B1(net5368),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][15] ),
    .A2(net5399),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][15] ));
 sg13g2_a21oi_1 _13163_ (.A1(_05148_),
    .A2(_05149_),
    .Y(_05150_),
    .B1(net5203));
 sg13g2_a22oi_1 _13164_ (.Y(_05151_),
    .B1(net5415),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][15] ),
    .A2(net5437),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][15] ));
 sg13g2_a22oi_1 _13165_ (.Y(_05152_),
    .B1(net5368),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][15] ),
    .A2(net5399),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][15] ));
 sg13g2_a21oi_1 _13166_ (.A1(_05151_),
    .A2(_05152_),
    .Y(_05153_),
    .B1(net5209));
 sg13g2_or4_1 _13167_ (.A(_05144_),
    .B(_05147_),
    .C(_05150_),
    .D(_05153_),
    .X(_00070_));
 sg13g2_a22oi_1 _13168_ (.Y(_05154_),
    .B1(net5430),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][16] ),
    .A2(net5452),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][16] ));
 sg13g2_a22oi_1 _13169_ (.Y(_05155_),
    .B1(net5384),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][16] ),
    .A2(net5408),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][16] ));
 sg13g2_a21oi_1 _13170_ (.A1(_05154_),
    .A2(_05155_),
    .Y(_05156_),
    .B1(net5205));
 sg13g2_a22oi_1 _13171_ (.Y(_05157_),
    .B1(net5430),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][16] ),
    .A2(net5452),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][16] ));
 sg13g2_a22oi_1 _13172_ (.Y(_05158_),
    .B1(net5383),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][16] ),
    .A2(net5408),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][16] ));
 sg13g2_a21oi_1 _13173_ (.A1(_05157_),
    .A2(_05158_),
    .Y(_05159_),
    .B1(net5362));
 sg13g2_a22oi_1 _13174_ (.Y(_05160_),
    .B1(net5430),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][16] ),
    .A2(net5452),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][16] ));
 sg13g2_a22oi_1 _13175_ (.Y(_05161_),
    .B1(net5383),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][16] ),
    .A2(net5408),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][16] ));
 sg13g2_a21oi_1 _13176_ (.A1(_05160_),
    .A2(_05161_),
    .Y(_05162_),
    .B1(net5216));
 sg13g2_a22oi_1 _13177_ (.Y(_05163_),
    .B1(net5430),
    .B2(net3933),
    .A2(net5452),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][16] ));
 sg13g2_a22oi_1 _13178_ (.Y(_05164_),
    .B1(net5383),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][16] ),
    .A2(net5408),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][16] ));
 sg13g2_a21oi_1 _13179_ (.A1(_05163_),
    .A2(_05164_),
    .Y(_05165_),
    .B1(net5210));
 sg13g2_or4_1 _13180_ (.A(_05156_),
    .B(_05159_),
    .C(_05162_),
    .D(_05165_),
    .X(_00071_));
 sg13g2_a22oi_1 _13181_ (.Y(_05166_),
    .B1(net5423),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][17] ),
    .A2(net5445),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][17] ));
 sg13g2_a22oi_1 _13182_ (.Y(_05167_),
    .B1(net5376),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][17] ),
    .A2(net5400),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][17] ));
 sg13g2_a21oi_1 _13183_ (.A1(_05166_),
    .A2(_05167_),
    .Y(_05168_),
    .B1(net5215));
 sg13g2_a22oi_1 _13184_ (.Y(_05169_),
    .B1(net5423),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][17] ),
    .A2(net5445),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][17] ));
 sg13g2_a22oi_1 _13185_ (.Y(_05170_),
    .B1(net5376),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][17] ),
    .A2(net5400),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][17] ));
 sg13g2_a21oi_1 _13186_ (.A1(_05169_),
    .A2(_05170_),
    .Y(_05171_),
    .B1(net5363));
 sg13g2_a22oi_1 _13187_ (.Y(_05172_),
    .B1(net5423),
    .B2(net3052),
    .A2(net5445),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][17] ));
 sg13g2_a22oi_1 _13188_ (.Y(_05173_),
    .B1(net5376),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][17] ),
    .A2(net5400),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][17] ));
 sg13g2_a21oi_1 _13189_ (.A1(_05172_),
    .A2(_05173_),
    .Y(_05174_),
    .B1(net5204));
 sg13g2_a22oi_1 _13190_ (.Y(_05175_),
    .B1(net5423),
    .B2(net3912),
    .A2(net5445),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][17] ));
 sg13g2_a22oi_1 _13191_ (.Y(_05176_),
    .B1(net5376),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][17] ),
    .A2(net5411),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][17] ));
 sg13g2_a21oi_1 _13192_ (.A1(_05175_),
    .A2(_05176_),
    .Y(_05177_),
    .B1(net5209));
 sg13g2_or4_1 _13193_ (.A(_05168_),
    .B(_05171_),
    .C(_05174_),
    .D(net3913),
    .X(_00072_));
 sg13g2_a22oi_1 _13194_ (.Y(_05178_),
    .B1(net5416),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][18] ),
    .A2(net5438),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][18] ));
 sg13g2_a22oi_1 _13195_ (.Y(_05179_),
    .B1(net5369),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][18] ),
    .A2(net5392),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][18] ));
 sg13g2_a21oi_1 _13196_ (.A1(_05178_),
    .A2(_05179_),
    .Y(_05180_),
    .B1(net5203));
 sg13g2_a22oi_1 _13197_ (.Y(_05181_),
    .B1(net5416),
    .B2(net3880),
    .A2(net5438),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][18] ));
 sg13g2_a22oi_1 _13198_ (.Y(_05182_),
    .B1(net5369),
    .B2(net2956),
    .A2(net5392),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][18] ));
 sg13g2_a21oi_1 _13199_ (.A1(_05181_),
    .A2(_05182_),
    .Y(_05183_),
    .B1(net5361));
 sg13g2_a22oi_1 _13200_ (.Y(_05184_),
    .B1(net5413),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][18] ),
    .A2(net5435),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][18] ));
 sg13g2_a22oi_1 _13201_ (.Y(_05185_),
    .B1(net5366),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][18] ),
    .A2(net5389),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][18] ));
 sg13g2_a21oi_1 _13202_ (.A1(_05184_),
    .A2(_05185_),
    .Y(_05186_),
    .B1(net5214));
 sg13g2_a22oi_1 _13203_ (.Y(_05187_),
    .B1(net5414),
    .B2(net2802),
    .A2(net5436),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][18] ));
 sg13g2_a22oi_1 _13204_ (.Y(_05188_),
    .B1(net5367),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][18] ),
    .A2(net5390),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][18] ));
 sg13g2_a21oi_1 _13205_ (.A1(_05187_),
    .A2(_05188_),
    .Y(_05189_),
    .B1(net5208));
 sg13g2_or4_1 _13206_ (.A(_05180_),
    .B(_05183_),
    .C(_05186_),
    .D(_05189_),
    .X(_00073_));
 sg13g2_a22oi_1 _13207_ (.Y(_05190_),
    .B1(net5416),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][19] ),
    .A2(net5438),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][19] ));
 sg13g2_a22oi_1 _13208_ (.Y(_05191_),
    .B1(net5369),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][19] ),
    .A2(net5391),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][19] ));
 sg13g2_a21oi_1 _13209_ (.A1(_05190_),
    .A2(_05191_),
    .Y(_05192_),
    .B1(net5203));
 sg13g2_a22oi_1 _13210_ (.Y(_05193_),
    .B1(net5416),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][19] ),
    .A2(net5438),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][19] ));
 sg13g2_a22oi_1 _13211_ (.Y(_05194_),
    .B1(net5369),
    .B2(net3140),
    .A2(net5391),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][19] ));
 sg13g2_a21oi_1 _13212_ (.A1(_05193_),
    .A2(_05194_),
    .Y(_05195_),
    .B1(net5361));
 sg13g2_a22oi_1 _13213_ (.Y(_05196_),
    .B1(net5415),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][19] ),
    .A2(net5438),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][19] ));
 sg13g2_a22oi_1 _13214_ (.Y(_05197_),
    .B1(net5369),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][19] ),
    .A2(net5391),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][19] ));
 sg13g2_a21oi_1 _13215_ (.A1(_05196_),
    .A2(_05197_),
    .Y(_05198_),
    .B1(net5214));
 sg13g2_a22oi_1 _13216_ (.Y(_05199_),
    .B1(net5416),
    .B2(net3922),
    .A2(net5437),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][19] ));
 sg13g2_a22oi_1 _13217_ (.Y(_05200_),
    .B1(net5368),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][19] ),
    .A2(net5391),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][19] ));
 sg13g2_a21oi_1 _13218_ (.A1(_05199_),
    .A2(_05200_),
    .Y(_05201_),
    .B1(net5208));
 sg13g2_or4_1 _13219_ (.A(_05192_),
    .B(_05195_),
    .C(_05198_),
    .D(_05201_),
    .X(_00074_));
 sg13g2_a22oi_1 _13220_ (.Y(_05202_),
    .B1(net5426),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][20] ),
    .A2(net5448),
    .A1(net3883));
 sg13g2_a22oi_1 _13221_ (.Y(_05203_),
    .B1(net5379),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][20] ),
    .A2(net5403),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][20] ));
 sg13g2_a21oi_1 _13222_ (.A1(net3884),
    .A2(_05203_),
    .Y(_05204_),
    .B1(net5204));
 sg13g2_a22oi_1 _13223_ (.Y(_05205_),
    .B1(net5425),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][20] ),
    .A2(net5447),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][20] ));
 sg13g2_a22oi_1 _13224_ (.Y(_05206_),
    .B1(net5378),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][20] ),
    .A2(net5404),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][20] ));
 sg13g2_a21oi_1 _13225_ (.A1(_05205_),
    .A2(_05206_),
    .Y(_05207_),
    .B1(net5209));
 sg13g2_a22oi_1 _13226_ (.Y(_05208_),
    .B1(net5426),
    .B2(net3879),
    .A2(net5448),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][20] ));
 sg13g2_a22oi_1 _13227_ (.Y(_05209_),
    .B1(net5378),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][20] ),
    .A2(net5403),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][20] ));
 sg13g2_a21oi_1 _13228_ (.A1(_05208_),
    .A2(_05209_),
    .Y(_05210_),
    .B1(net5215));
 sg13g2_a22oi_1 _13229_ (.Y(_05211_),
    .B1(net5425),
    .B2(net2620),
    .A2(net5447),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][20] ));
 sg13g2_a22oi_1 _13230_ (.Y(_05212_),
    .B1(net5378),
    .B2(net3025),
    .A2(net5403),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][20] ));
 sg13g2_a21oi_1 _13231_ (.A1(_05211_),
    .A2(_05212_),
    .Y(_05213_),
    .B1(net5363));
 sg13g2_or4_1 _13232_ (.A(net3885),
    .B(_05207_),
    .C(_05210_),
    .D(_05213_),
    .X(_00076_));
 sg13g2_a22oi_1 _13233_ (.Y(_05214_),
    .B1(net5423),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][21] ),
    .A2(net5445),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][21] ));
 sg13g2_a22oi_1 _13234_ (.Y(_05215_),
    .B1(net5376),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][21] ),
    .A2(net5400),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][21] ));
 sg13g2_a21oi_1 _13235_ (.A1(_05214_),
    .A2(_05215_),
    .Y(_05216_),
    .B1(net5204));
 sg13g2_a22oi_1 _13236_ (.Y(_05217_),
    .B1(net5422),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][21] ),
    .A2(net5444),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][21] ));
 sg13g2_a22oi_1 _13237_ (.Y(_05218_),
    .B1(net5375),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][21] ),
    .A2(net5400),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][21] ));
 sg13g2_a21oi_1 _13238_ (.A1(_05217_),
    .A2(_05218_),
    .Y(_05219_),
    .B1(net5363));
 sg13g2_a22oi_1 _13239_ (.Y(_05220_),
    .B1(net5422),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][21] ),
    .A2(net5444),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][21] ));
 sg13g2_a22oi_1 _13240_ (.Y(_05221_),
    .B1(net5375),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][21] ),
    .A2(net5401),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][21] ));
 sg13g2_a21oi_1 _13241_ (.A1(_05220_),
    .A2(_05221_),
    .Y(_05222_),
    .B1(net5216));
 sg13g2_a22oi_1 _13242_ (.Y(_05223_),
    .B1(net5422),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][21] ),
    .A2(net5444),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][21] ));
 sg13g2_a22oi_1 _13243_ (.Y(_05224_),
    .B1(net5375),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][21] ),
    .A2(net5400),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][21] ));
 sg13g2_a21oi_1 _13244_ (.A1(_05223_),
    .A2(_05224_),
    .Y(_05225_),
    .B1(net5209));
 sg13g2_or4_1 _13245_ (.A(_05216_),
    .B(_05219_),
    .C(_05222_),
    .D(_05225_),
    .X(_00077_));
 sg13g2_a22oi_1 _13246_ (.Y(_05226_),
    .B1(net5424),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][22] ),
    .A2(net5446),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][22] ));
 sg13g2_a22oi_1 _13247_ (.Y(_05227_),
    .B1(net5377),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][22] ),
    .A2(net5402),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][22] ));
 sg13g2_a21oi_1 _13248_ (.A1(_05226_),
    .A2(_05227_),
    .Y(_05228_),
    .B1(net5204));
 sg13g2_a22oi_1 _13249_ (.Y(_05229_),
    .B1(net5424),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][22] ),
    .A2(net5446),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][22] ));
 sg13g2_a22oi_1 _13250_ (.Y(_05230_),
    .B1(net5377),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][22] ),
    .A2(net5402),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][22] ));
 sg13g2_a21oi_1 _13251_ (.A1(_05229_),
    .A2(_05230_),
    .Y(_05231_),
    .B1(net5363));
 sg13g2_a22oi_1 _13252_ (.Y(_05232_),
    .B1(net5424),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][22] ),
    .A2(net5446),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][22] ));
 sg13g2_a22oi_1 _13253_ (.Y(_05233_),
    .B1(net5377),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][22] ),
    .A2(net5402),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][22] ));
 sg13g2_a21oi_1 _13254_ (.A1(_05232_),
    .A2(_05233_),
    .Y(_05234_),
    .B1(net5215));
 sg13g2_a22oi_1 _13255_ (.Y(_05235_),
    .B1(net5424),
    .B2(net3928),
    .A2(net5446),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][22] ));
 sg13g2_a22oi_1 _13256_ (.Y(_05236_),
    .B1(net5379),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][22] ),
    .A2(net5404),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][22] ));
 sg13g2_a21oi_1 _13257_ (.A1(_05235_),
    .A2(_05236_),
    .Y(_05237_),
    .B1(net5209));
 sg13g2_or4_1 _13258_ (.A(_05228_),
    .B(_05231_),
    .C(_05234_),
    .D(net3929),
    .X(_00078_));
 sg13g2_a22oi_1 _13259_ (.Y(_05238_),
    .B1(net5426),
    .B2(net2906),
    .A2(net5448),
    .A1(net3890));
 sg13g2_a22oi_1 _13260_ (.Y(_05239_),
    .B1(net5377),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][23] ),
    .A2(net5401),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][23] ));
 sg13g2_a21oi_1 _13261_ (.A1(_05238_),
    .A2(_05239_),
    .Y(_05240_),
    .B1(net5204));
 sg13g2_a22oi_1 _13262_ (.Y(_05241_),
    .B1(net5424),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][23] ),
    .A2(net5446),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][23] ));
 sg13g2_a22oi_1 _13263_ (.Y(_05242_),
    .B1(net5379),
    .B2(net2864),
    .A2(net5401),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][23] ));
 sg13g2_a21oi_1 _13264_ (.A1(_05241_),
    .A2(_05242_),
    .Y(_05243_),
    .B1(net5363));
 sg13g2_a22oi_1 _13265_ (.Y(_05244_),
    .B1(net5426),
    .B2(net2695),
    .A2(net5448),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][23] ));
 sg13g2_a22oi_1 _13266_ (.Y(_05245_),
    .B1(net5379),
    .B2(net3109),
    .A2(net5401),
    .A1(net3247));
 sg13g2_a21oi_1 _13267_ (.A1(_05244_),
    .A2(_05245_),
    .Y(_05246_),
    .B1(net5215));
 sg13g2_a22oi_1 _13268_ (.Y(_05247_),
    .B1(net5426),
    .B2(net2729),
    .A2(net5448),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][23] ));
 sg13g2_a22oi_1 _13269_ (.Y(_05248_),
    .B1(net5379),
    .B2(net2732),
    .A2(net5402),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][23] ));
 sg13g2_a21oi_1 _13270_ (.A1(_05247_),
    .A2(_05248_),
    .Y(_05249_),
    .B1(net5211));
 sg13g2_or4_1 _13271_ (.A(_05240_),
    .B(_05243_),
    .C(_05246_),
    .D(_05249_),
    .X(_00079_));
 sg13g2_a22oi_1 _13272_ (.Y(_05250_),
    .B1(net5424),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][24] ),
    .A2(net5446),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][24] ));
 sg13g2_a22oi_1 _13273_ (.Y(_05251_),
    .B1(net5377),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][24] ),
    .A2(net5401),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][24] ));
 sg13g2_a21oi_1 _13274_ (.A1(_05250_),
    .A2(_05251_),
    .Y(_05252_),
    .B1(net5204));
 sg13g2_a22oi_1 _13275_ (.Y(_05253_),
    .B1(net5424),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][24] ),
    .A2(net5446),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][24] ));
 sg13g2_a22oi_1 _13276_ (.Y(_05254_),
    .B1(net5377),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][24] ),
    .A2(net5401),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][24] ));
 sg13g2_a21oi_1 _13277_ (.A1(_05253_),
    .A2(_05254_),
    .Y(_05255_),
    .B1(net5363));
 sg13g2_a22oi_1 _13278_ (.Y(_05256_),
    .B1(net5424),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][24] ),
    .A2(net5446),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][24] ));
 sg13g2_a22oi_1 _13279_ (.Y(_05257_),
    .B1(net5377),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][24] ),
    .A2(net5401),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][24] ));
 sg13g2_a21oi_1 _13280_ (.A1(_05256_),
    .A2(_05257_),
    .Y(_05258_),
    .B1(net5216));
 sg13g2_a22oi_1 _13281_ (.Y(_05259_),
    .B1(net5425),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][24] ),
    .A2(net5447),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][24] ));
 sg13g2_a22oi_1 _13282_ (.Y(_05260_),
    .B1(net5377),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][24] ),
    .A2(net5401),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][24] ));
 sg13g2_a21oi_1 _13283_ (.A1(_05259_),
    .A2(_05260_),
    .Y(_05261_),
    .B1(net5209));
 sg13g2_or4_1 _13284_ (.A(_05252_),
    .B(_05255_),
    .C(_05258_),
    .D(_05261_),
    .X(_00080_));
 sg13g2_a22oi_1 _13285_ (.Y(_05262_),
    .B1(net5422),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][25] ),
    .A2(net5444),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][25] ));
 sg13g2_a22oi_1 _13286_ (.Y(_05263_),
    .B1(net5375),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][25] ),
    .A2(net5399),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][25] ));
 sg13g2_a21oi_1 _13287_ (.A1(_05262_),
    .A2(_05263_),
    .Y(_05264_),
    .B1(net5215));
 sg13g2_a22oi_1 _13288_ (.Y(_05265_),
    .B1(net5422),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][25] ),
    .A2(net5444),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][25] ));
 sg13g2_a22oi_1 _13289_ (.Y(_05266_),
    .B1(net5375),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][25] ),
    .A2(net5399),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][25] ));
 sg13g2_a21oi_1 _13290_ (.A1(_05265_),
    .A2(_05266_),
    .Y(_05267_),
    .B1(net5209));
 sg13g2_a22oi_1 _13291_ (.Y(_05268_),
    .B1(net5422),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][25] ),
    .A2(net5444),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][25] ));
 sg13g2_a22oi_1 _13292_ (.Y(_05269_),
    .B1(net5375),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][25] ),
    .A2(net5399),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][25] ));
 sg13g2_a21oi_1 _13293_ (.A1(_05268_),
    .A2(_05269_),
    .Y(_05270_),
    .B1(net5204));
 sg13g2_a22oi_1 _13294_ (.Y(_05271_),
    .B1(net5422),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][25] ),
    .A2(net5444),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][25] ));
 sg13g2_a22oi_1 _13295_ (.Y(_05272_),
    .B1(net5375),
    .B2(net3941),
    .A2(net5399),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][25] ));
 sg13g2_a21oi_1 _13296_ (.A1(_05271_),
    .A2(_05272_),
    .Y(_05273_),
    .B1(net5363));
 sg13g2_or4_2 _13297_ (.A(_05264_),
    .B(_05267_),
    .C(_05270_),
    .D(_05273_),
    .X(_00081_));
 sg13g2_a22oi_1 _13298_ (.Y(_05274_),
    .B1(net5425),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][26] ),
    .A2(net5447),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][26] ));
 sg13g2_a22oi_1 _13299_ (.Y(_05275_),
    .B1(net5378),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][26] ),
    .A2(net5403),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][26] ));
 sg13g2_a21oi_1 _13300_ (.A1(_05274_),
    .A2(_05275_),
    .Y(_05276_),
    .B1(net5215));
 sg13g2_a22oi_1 _13301_ (.Y(_05277_),
    .B1(net5431),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][26] ),
    .A2(net5453),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][26] ));
 sg13g2_a22oi_1 _13302_ (.Y(_05278_),
    .B1(net5385),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][26] ),
    .A2(net5407),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][26] ));
 sg13g2_a21oi_1 _13303_ (.A1(_05277_),
    .A2(_05278_),
    .Y(_05279_),
    .B1(net5210));
 sg13g2_a22oi_1 _13304_ (.Y(_05280_),
    .B1(net5425),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][26] ),
    .A2(net5447),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][26] ));
 sg13g2_a22oi_1 _13305_ (.Y(_05281_),
    .B1(net5378),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][26] ),
    .A2(net5403),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][26] ));
 sg13g2_a21oi_1 _13306_ (.A1(_05280_),
    .A2(_05281_),
    .Y(_05282_),
    .B1(net5204));
 sg13g2_a22oi_1 _13307_ (.Y(_05283_),
    .B1(net5429),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][26] ),
    .A2(net5451),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][26] ));
 sg13g2_a22oi_1 _13308_ (.Y(_05284_),
    .B1(net5385),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][26] ),
    .A2(net5410),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][26] ));
 sg13g2_a21oi_1 _13309_ (.A1(_05283_),
    .A2(_05284_),
    .Y(_05285_),
    .B1(net5364));
 sg13g2_or4_1 _13310_ (.A(_05276_),
    .B(_05279_),
    .C(_05282_),
    .D(_05285_),
    .X(_00082_));
 sg13g2_a22oi_1 _13311_ (.Y(_05286_),
    .B1(net5418),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][27] ),
    .A2(net5440),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][27] ));
 sg13g2_a22oi_1 _13312_ (.Y(_05287_),
    .B1(net5371),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][27] ),
    .A2(net5395),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][27] ));
 sg13g2_a21oi_1 _13313_ (.A1(_05286_),
    .A2(_05287_),
    .Y(_05288_),
    .B1(net5213));
 sg13g2_a22oi_1 _13314_ (.Y(_05289_),
    .B1(net5418),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][27] ),
    .A2(net5440),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][27] ));
 sg13g2_a22oi_1 _13315_ (.Y(_05290_),
    .B1(net5371),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][27] ),
    .A2(net5395),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][27] ));
 sg13g2_a21oi_1 _13316_ (.A1(_05289_),
    .A2(_05290_),
    .Y(_05291_),
    .B1(net5207));
 sg13g2_a22oi_1 _13317_ (.Y(_05292_),
    .B1(net5418),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][27] ),
    .A2(net5440),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][27] ));
 sg13g2_a22oi_1 _13318_ (.Y(_05293_),
    .B1(net5371),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][27] ),
    .A2(net5395),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][27] ));
 sg13g2_a21oi_1 _13319_ (.A1(_05292_),
    .A2(_05293_),
    .Y(_05294_),
    .B1(net5202));
 sg13g2_a22oi_1 _13320_ (.Y(_05295_),
    .B1(net5418),
    .B2(net3898),
    .A2(net5440),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][27] ));
 sg13g2_a22oi_1 _13321_ (.Y(_05296_),
    .B1(net5371),
    .B2(net3208),
    .A2(net5395),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][27] ));
 sg13g2_a21oi_1 _13322_ (.A1(_05295_),
    .A2(_05296_),
    .Y(_05297_),
    .B1(net5360));
 sg13g2_or4_1 _13323_ (.A(_05288_),
    .B(_05291_),
    .C(_05294_),
    .D(_05297_),
    .X(_00083_));
 sg13g2_a22oi_1 _13324_ (.Y(_05298_),
    .B1(net5428),
    .B2(net3893),
    .A2(net5450),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][28] ));
 sg13g2_a22oi_1 _13325_ (.Y(_05299_),
    .B1(net5381),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][28] ),
    .A2(net5406),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][28] ));
 sg13g2_a21oi_1 _13326_ (.A1(_05298_),
    .A2(_05299_),
    .Y(_05300_),
    .B1(net5206));
 sg13g2_a22oi_1 _13327_ (.Y(_05301_),
    .B1(net5428),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][28] ),
    .A2(net5450),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][28] ));
 sg13g2_a22oi_1 _13328_ (.Y(_05302_),
    .B1(net5380),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][28] ),
    .A2(net5405),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][28] ));
 sg13g2_a21oi_1 _13329_ (.A1(_05301_),
    .A2(_05302_),
    .Y(_05303_),
    .B1(net5210));
 sg13g2_a22oi_1 _13330_ (.Y(_05304_),
    .B1(net5428),
    .B2(net3045),
    .A2(net5450),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][28] ));
 sg13g2_a22oi_1 _13331_ (.Y(_05305_),
    .B1(net5380),
    .B2(net3179),
    .A2(net5405),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][28] ));
 sg13g2_a21oi_1 _13332_ (.A1(_05304_),
    .A2(_05305_),
    .Y(_05306_),
    .B1(net5216));
 sg13g2_a22oi_1 _13333_ (.Y(_05307_),
    .B1(net5427),
    .B2(net2609),
    .A2(net5449),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][28] ));
 sg13g2_a22oi_1 _13334_ (.Y(_05308_),
    .B1(net5381),
    .B2(net2967),
    .A2(net5405),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][28] ));
 sg13g2_a21oi_1 _13335_ (.A1(_05307_),
    .A2(_05308_),
    .Y(_05309_),
    .B1(net5362));
 sg13g2_or4_1 _13336_ (.A(net3894),
    .B(_05303_),
    .C(_05306_),
    .D(_05309_),
    .X(_00084_));
 sg13g2_a22oi_1 _13337_ (.Y(_05310_),
    .B1(net5429),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][29] ),
    .A2(net5451),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][29] ));
 sg13g2_a22oi_1 _13338_ (.Y(_05311_),
    .B1(net5382),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][29] ),
    .A2(net5407),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][29] ));
 sg13g2_a21oi_1 _13339_ (.A1(_05310_),
    .A2(_05311_),
    .Y(_05312_),
    .B1(net5217));
 sg13g2_a22oi_1 _13340_ (.Y(_05313_),
    .B1(net5429),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][29] ),
    .A2(net5451),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][29] ));
 sg13g2_a22oi_1 _13341_ (.Y(_05314_),
    .B1(net5382),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][29] ),
    .A2(net5407),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][29] ));
 sg13g2_a21oi_1 _13342_ (.A1(_05313_),
    .A2(_05314_),
    .Y(_05315_),
    .B1(net5362));
 sg13g2_a22oi_1 _13343_ (.Y(_05316_),
    .B1(net5428),
    .B2(net3925),
    .A2(net5450),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][29] ));
 sg13g2_a22oi_1 _13344_ (.Y(_05317_),
    .B1(net5380),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][29] ),
    .A2(net5405),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][29] ));
 sg13g2_a21oi_1 _13345_ (.A1(_05316_),
    .A2(_05317_),
    .Y(_05318_),
    .B1(net5205));
 sg13g2_a22oi_1 _13346_ (.Y(_05319_),
    .B1(net5428),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[10][29] ),
    .A2(net5450),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][29] ));
 sg13g2_a22oi_1 _13347_ (.Y(_05320_),
    .B1(net5380),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][29] ),
    .A2(net5405),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][29] ));
 sg13g2_a21oi_1 _13348_ (.A1(_05319_),
    .A2(_05320_),
    .Y(_05321_),
    .B1(net5210));
 sg13g2_or4_1 _13349_ (.A(_05312_),
    .B(_05315_),
    .C(net3926),
    .D(_05321_),
    .X(_00085_));
 sg13g2_a22oi_1 _13350_ (.Y(_05322_),
    .B1(net5419),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][30] ),
    .A2(net5441),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][30] ));
 sg13g2_a22oi_1 _13351_ (.Y(_05323_),
    .B1(net5372),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][30] ),
    .A2(net5396),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][30] ));
 sg13g2_a21oi_1 _13352_ (.A1(_05322_),
    .A2(_05323_),
    .Y(_05324_),
    .B1(net5206));
 sg13g2_a22oi_1 _13353_ (.Y(_05325_),
    .B1(net5419),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][30] ),
    .A2(net5441),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][30] ));
 sg13g2_a22oi_1 _13354_ (.Y(_05326_),
    .B1(net5372),
    .B2(net3130),
    .A2(net5396),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][30] ));
 sg13g2_a21oi_1 _13355_ (.A1(_05325_),
    .A2(_05326_),
    .Y(_05327_),
    .B1(net5364));
 sg13g2_a22oi_1 _13356_ (.Y(_05328_),
    .B1(net5419),
    .B2(net3899),
    .A2(net5441),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][30] ));
 sg13g2_a22oi_1 _13357_ (.Y(_05329_),
    .B1(net5372),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][30] ),
    .A2(net5396),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][30] ));
 sg13g2_a21oi_1 _13358_ (.A1(_05328_),
    .A2(_05329_),
    .Y(_05330_),
    .B1(net5217));
 sg13g2_a22oi_1 _13359_ (.Y(_05331_),
    .B1(net5419),
    .B2(net2839),
    .A2(net5441),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][30] ));
 sg13g2_a22oi_1 _13360_ (.Y(_05332_),
    .B1(net5372),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][30] ),
    .A2(net5396),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][30] ));
 sg13g2_a21oi_1 _13361_ (.A1(_05331_),
    .A2(_05332_),
    .Y(_05333_),
    .B1(net5212));
 sg13g2_or4_1 _13362_ (.A(_05324_),
    .B(_05327_),
    .C(net3900),
    .D(_05333_),
    .X(_00087_));
 sg13g2_a22oi_1 _13363_ (.Y(_05334_),
    .B1(net5430),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[6][31] ),
    .A2(net5452),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[5][31] ));
 sg13g2_a22oi_1 _13364_ (.Y(_05335_),
    .B1(net5383),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[7][31] ),
    .A2(net5408),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][31] ));
 sg13g2_a21oi_1 _13365_ (.A1(_05334_),
    .A2(_05335_),
    .Y(_05336_),
    .B1(net5216));
 sg13g2_a22oi_1 _13366_ (.Y(_05337_),
    .B1(net5427),
    .B2(net3938),
    .A2(net5449),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][31] ));
 sg13g2_a22oi_1 _13367_ (.Y(_05338_),
    .B1(net5381),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[11][31] ),
    .A2(net5405),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][31] ));
 sg13g2_a21oi_1 _13368_ (.A1(_05337_),
    .A2(_05338_),
    .Y(_05339_),
    .B1(net5210));
 sg13g2_a22oi_1 _13369_ (.Y(_05340_),
    .B1(net5427),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[2][31] ),
    .A2(net5449),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][31] ));
 sg13g2_a22oi_1 _13370_ (.Y(_05341_),
    .B1(net5380),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[3][31] ),
    .A2(net5405),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][31] ));
 sg13g2_a21oi_1 _13371_ (.A1(_05340_),
    .A2(_05341_),
    .Y(_05342_),
    .B1(net5205));
 sg13g2_a22oi_1 _13372_ (.Y(_05343_),
    .B1(net5430),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[14][31] ),
    .A2(net5452),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[13][31] ));
 sg13g2_a22oi_1 _13373_ (.Y(_05344_),
    .B1(net5383),
    .B2(\TRNG.sha256.expand.msg_schdl.RAM[15][31] ),
    .A2(net5408),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[12][31] ));
 sg13g2_a21oi_1 _13374_ (.A1(_05343_),
    .A2(_05344_),
    .Y(_05345_),
    .B1(net5362));
 sg13g2_or4_1 _13375_ (.A(_05336_),
    .B(_05339_),
    .C(_05342_),
    .D(_05345_),
    .X(_00088_));
 sg13g2_mux2_1 _13376_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[14][0] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[15][0] ),
    .S(net5761),
    .X(_05346_));
 sg13g2_nor2b_1 _13377_ (.A(net5761),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][0] ),
    .Y(_05347_));
 sg13g2_a21oi_1 _13378_ (.A1(net5761),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][0] ),
    .Y(_05348_),
    .B1(_05347_));
 sg13g2_o21ai_1 _13379_ (.B1(net5702),
    .Y(_05349_),
    .A1(net5726),
    .A2(_05348_));
 sg13g2_a21oi_1 _13380_ (.A1(net5726),
    .A2(_05346_),
    .Y(_05350_),
    .B1(_05349_));
 sg13g2_mux4_1 _13381_ (.S0(net5765),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][0] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][0] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][0] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][0] ),
    .S1(net5727),
    .X(_05351_));
 sg13g2_o21ai_1 _13382_ (.B1(net5691),
    .Y(_05352_),
    .A1(net5702),
    .A2(_05351_));
 sg13g2_mux4_1 _13383_ (.S0(net5761),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][0] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][0] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][0] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][0] ),
    .S1(net5726),
    .X(_05353_));
 sg13g2_mux2_1 _13384_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][0] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][0] ),
    .S(net5761),
    .X(_05354_));
 sg13g2_nor2b_1 _13385_ (.A(net5761),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][0] ),
    .Y(_05355_));
 sg13g2_a21oi_1 _13386_ (.A1(net5761),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][0] ),
    .Y(_05356_),
    .B1(_05355_));
 sg13g2_o21ai_1 _13387_ (.B1(net5702),
    .Y(_05357_),
    .A1(net5726),
    .A2(_05356_));
 sg13g2_a21oi_1 _13388_ (.A1(net5726),
    .A2(_05354_),
    .Y(_05358_),
    .B1(_05357_));
 sg13g2_nor2_1 _13389_ (.A(net5691),
    .B(_05358_),
    .Y(_05359_));
 sg13g2_o21ai_1 _13390_ (.B1(_05359_),
    .Y(_05360_),
    .A1(net5702),
    .A2(_05353_));
 sg13g2_o21ai_1 _13391_ (.B1(_05360_),
    .Y(_00032_),
    .A1(_05350_),
    .A2(_05352_));
 sg13g2_mux4_1 _13392_ (.S0(net5766),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][1] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][1] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][1] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][1] ),
    .S1(net5729),
    .X(_05361_));
 sg13g2_nor2_1 _13393_ (.A(net5704),
    .B(_05361_),
    .Y(_05362_));
 sg13g2_nor2b_1 _13394_ (.A(net5767),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][1] ),
    .Y(_05363_));
 sg13g2_a21oi_1 _13395_ (.A1(net5766),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][1] ),
    .Y(_05364_),
    .B1(_05363_));
 sg13g2_o21ai_1 _13396_ (.B1(net5733),
    .Y(_05365_),
    .A1(net5766),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][1] ));
 sg13g2_a21oi_1 _13397_ (.A1(net5766),
    .A2(_04344_),
    .Y(_05366_),
    .B1(_05365_));
 sg13g2_o21ai_1 _13398_ (.B1(net5704),
    .Y(_05367_),
    .A1(net5729),
    .A2(_05364_));
 sg13g2_o21ai_1 _13399_ (.B1(net5691),
    .Y(_05368_),
    .A1(_05366_),
    .A2(_05367_));
 sg13g2_mux4_1 _13400_ (.S0(net5766),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][1] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][1] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][1] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][1] ),
    .S1(net5729),
    .X(_05369_));
 sg13g2_mux2_1 _13401_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][1] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][1] ),
    .S(net5766),
    .X(_05370_));
 sg13g2_nor2b_1 _13402_ (.A(net5766),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][1] ),
    .Y(_05371_));
 sg13g2_a21oi_1 _13403_ (.A1(net5766),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][1] ),
    .Y(_05372_),
    .B1(_05371_));
 sg13g2_o21ai_1 _13404_ (.B1(net5704),
    .Y(_05373_),
    .A1(net5729),
    .A2(_05372_));
 sg13g2_a21oi_1 _13405_ (.A1(net5729),
    .A2(_05370_),
    .Y(_05374_),
    .B1(_05373_));
 sg13g2_nor2_1 _13406_ (.A(net5692),
    .B(_05374_),
    .Y(_05375_));
 sg13g2_o21ai_1 _13407_ (.B1(_05375_),
    .Y(_05376_),
    .A1(net5704),
    .A2(_05369_));
 sg13g2_o21ai_1 _13408_ (.B1(_05376_),
    .Y(_00043_),
    .A1(_05362_),
    .A2(_05368_));
 sg13g2_mux2_1 _13409_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[10][2] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[11][2] ),
    .S(net5774),
    .X(_05377_));
 sg13g2_nor2b_1 _13410_ (.A(net5774),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[8][2] ),
    .Y(_05378_));
 sg13g2_a21oi_1 _13411_ (.A1(net5775),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[9][2] ),
    .Y(_05379_),
    .B1(_05378_));
 sg13g2_a21oi_1 _13412_ (.A1(net5734),
    .A2(_05377_),
    .Y(_05380_),
    .B1(net5707));
 sg13g2_o21ai_1 _13413_ (.B1(_05380_),
    .Y(_05381_),
    .A1(net5735),
    .A2(_05379_));
 sg13g2_nor2b_1 _13414_ (.A(net5775),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][2] ),
    .Y(_05382_));
 sg13g2_a21oi_1 _13415_ (.A1(net5775),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][2] ),
    .Y(_05383_),
    .B1(_05382_));
 sg13g2_mux2_1 _13416_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[14][2] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[15][2] ),
    .S(net5775),
    .X(_05384_));
 sg13g2_o21ai_1 _13417_ (.B1(net5707),
    .Y(_05385_),
    .A1(net5735),
    .A2(_05383_));
 sg13g2_a21o_1 _13418_ (.A2(_05384_),
    .A1(net5734),
    .B1(_05385_),
    .X(_05386_));
 sg13g2_nand3_1 _13419_ (.B(_05381_),
    .C(_05386_),
    .A(net5693),
    .Y(_05387_));
 sg13g2_mux2_1 _13420_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[2][2] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[3][2] ),
    .S(net5775),
    .X(_05388_));
 sg13g2_nor2b_1 _13421_ (.A(net5775),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[0][2] ),
    .Y(_05389_));
 sg13g2_a21oi_1 _13422_ (.A1(net5775),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[1][2] ),
    .Y(_05390_),
    .B1(_05389_));
 sg13g2_a21oi_1 _13423_ (.A1(net5735),
    .A2(_05388_),
    .Y(_05391_),
    .B1(net5707));
 sg13g2_o21ai_1 _13424_ (.B1(_05391_),
    .Y(_05392_),
    .A1(net5735),
    .A2(_05390_));
 sg13g2_o21ai_1 _13425_ (.B1(net5735),
    .Y(_05393_),
    .A1(net5776),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[6][2] ));
 sg13g2_a21oi_1 _13426_ (.A1(net5776),
    .A2(_04345_),
    .Y(_05394_),
    .B1(_05393_));
 sg13g2_nor2b_1 _13427_ (.A(net5776),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][2] ),
    .Y(_05395_));
 sg13g2_a21oi_1 _13428_ (.A1(net5776),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][2] ),
    .Y(_05396_),
    .B1(_05395_));
 sg13g2_o21ai_1 _13429_ (.B1(net5707),
    .Y(_05397_),
    .A1(net5735),
    .A2(_05396_));
 sg13g2_o21ai_1 _13430_ (.B1(_05392_),
    .Y(_05398_),
    .A1(_05394_),
    .A2(_05397_));
 sg13g2_o21ai_1 _13431_ (.B1(_05387_),
    .Y(_00054_),
    .A1(net5693),
    .A2(_05398_));
 sg13g2_mux2_1 _13432_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[10][3] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[11][3] ),
    .S(net5799),
    .X(_05399_));
 sg13g2_nor2b_1 _13433_ (.A(net5799),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[8][3] ),
    .Y(_05400_));
 sg13g2_a21oi_1 _13434_ (.A1(net5799),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[9][3] ),
    .Y(_05401_),
    .B1(_05400_));
 sg13g2_a21oi_1 _13435_ (.A1(net5749),
    .A2(_05399_),
    .Y(_05402_),
    .B1(net5716));
 sg13g2_o21ai_1 _13436_ (.B1(_05402_),
    .Y(_05403_),
    .A1(net5749),
    .A2(_05401_));
 sg13g2_nor2b_1 _13437_ (.A(net5789),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][3] ),
    .Y(_05404_));
 sg13g2_a21oi_1 _13438_ (.A1(net5789),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][3] ),
    .Y(_05405_),
    .B1(_05404_));
 sg13g2_mux2_1 _13439_ (.A0(net2682),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[15][3] ),
    .S(net5789),
    .X(_05406_));
 sg13g2_o21ai_1 _13440_ (.B1(net5713),
    .Y(_05407_),
    .A1(net5744),
    .A2(_05405_));
 sg13g2_a21oi_1 _13441_ (.A1(net5744),
    .A2(_05406_),
    .Y(_05408_),
    .B1(_05407_));
 sg13g2_nand2_1 _13442_ (.Y(_05409_),
    .A(net5696),
    .B(_05403_));
 sg13g2_mux4_1 _13443_ (.S0(net5789),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][3] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][3] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][3] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][3] ),
    .S1(net5749),
    .X(_05410_));
 sg13g2_mux2_1 _13444_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][3] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][3] ),
    .S(net5799),
    .X(_05411_));
 sg13g2_nor2b_1 _13445_ (.A(net5799),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][3] ),
    .Y(_05412_));
 sg13g2_a21oi_1 _13446_ (.A1(net5799),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][3] ),
    .Y(_05413_),
    .B1(_05412_));
 sg13g2_o21ai_1 _13447_ (.B1(net5716),
    .Y(_05414_),
    .A1(net5749),
    .A2(_05413_));
 sg13g2_a21oi_1 _13448_ (.A1(net5749),
    .A2(_05411_),
    .Y(_05415_),
    .B1(_05414_));
 sg13g2_nor2_1 _13449_ (.A(net5696),
    .B(_05415_),
    .Y(_05416_));
 sg13g2_o21ai_1 _13450_ (.B1(_05416_),
    .Y(_05417_),
    .A1(net5716),
    .A2(_05410_));
 sg13g2_o21ai_1 _13451_ (.B1(_05417_),
    .Y(_00057_),
    .A1(_05408_),
    .A2(_05409_));
 sg13g2_mux4_1 _13452_ (.S0(net5779),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][4] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][4] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][4] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][4] ),
    .S1(net5737),
    .X(_05418_));
 sg13g2_nor2b_1 _13453_ (.A(net5779),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][4] ),
    .Y(_05419_));
 sg13g2_a21oi_1 _13454_ (.A1(net5779),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][4] ),
    .Y(_05420_),
    .B1(_05419_));
 sg13g2_mux2_1 _13455_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[14][4] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[15][4] ),
    .S(net5779),
    .X(_05421_));
 sg13g2_o21ai_1 _13456_ (.B1(net5706),
    .Y(_05422_),
    .A1(net5737),
    .A2(_05420_));
 sg13g2_a21oi_1 _13457_ (.A1(net5737),
    .A2(_05421_),
    .Y(_05423_),
    .B1(_05422_));
 sg13g2_nor2b_1 _13458_ (.A(_05423_),
    .B_N(net5693),
    .Y(_05424_));
 sg13g2_o21ai_1 _13459_ (.B1(_05424_),
    .Y(_05425_),
    .A1(net5706),
    .A2(_05418_));
 sg13g2_mux2_1 _13460_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[2][4] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[3][4] ),
    .S(net5777),
    .X(_05426_));
 sg13g2_nor2b_1 _13461_ (.A(net5777),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[0][4] ),
    .Y(_05427_));
 sg13g2_a21oi_1 _13462_ (.A1(net5777),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[1][4] ),
    .Y(_05428_),
    .B1(_05427_));
 sg13g2_a21oi_1 _13463_ (.A1(net5736),
    .A2(_05426_),
    .Y(_05429_),
    .B1(net5706));
 sg13g2_o21ai_1 _13464_ (.B1(_05429_),
    .Y(_05430_),
    .A1(net5736),
    .A2(_05428_));
 sg13g2_o21ai_1 _13465_ (.B1(net5736),
    .Y(_05431_),
    .A1(net5777),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[6][4] ));
 sg13g2_a21oi_1 _13466_ (.A1(net5777),
    .A2(_04346_),
    .Y(_05432_),
    .B1(_05431_));
 sg13g2_nor2b_1 _13467_ (.A(net5775),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][4] ),
    .Y(_05433_));
 sg13g2_a21oi_1 _13468_ (.A1(net5777),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][4] ),
    .Y(_05434_),
    .B1(_05433_));
 sg13g2_o21ai_1 _13469_ (.B1(net5710),
    .Y(_05435_),
    .A1(net5736),
    .A2(_05434_));
 sg13g2_o21ai_1 _13470_ (.B1(_05430_),
    .Y(_05436_),
    .A1(_05432_),
    .A2(_05435_));
 sg13g2_o21ai_1 _13471_ (.B1(_05425_),
    .Y(_00058_),
    .A1(net5693),
    .A2(_05436_));
 sg13g2_mux4_1 _13472_ (.S0(net5781),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][5] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][5] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][5] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][5] ),
    .S1(net5738),
    .X(_05437_));
 sg13g2_nor2_1 _13473_ (.A(net5708),
    .B(_05437_),
    .Y(_05438_));
 sg13g2_nor2b_1 _13474_ (.A(net5781),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][5] ),
    .Y(_05439_));
 sg13g2_a21oi_1 _13475_ (.A1(net5781),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][5] ),
    .Y(_05440_),
    .B1(_05439_));
 sg13g2_o21ai_1 _13476_ (.B1(net5738),
    .Y(_05441_),
    .A1(net5781),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][5] ));
 sg13g2_a21oi_1 _13477_ (.A1(net5781),
    .A2(_04347_),
    .Y(_05442_),
    .B1(_05441_));
 sg13g2_o21ai_1 _13478_ (.B1(net5708),
    .Y(_05443_),
    .A1(net5738),
    .A2(_05440_));
 sg13g2_o21ai_1 _13479_ (.B1(net5694),
    .Y(_05444_),
    .A1(_05442_),
    .A2(_05443_));
 sg13g2_mux4_1 _13480_ (.S0(net5781),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][5] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][5] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][5] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][5] ),
    .S1(net5738),
    .X(_05445_));
 sg13g2_mux2_1 _13481_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][5] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][5] ),
    .S(net5783),
    .X(_05446_));
 sg13g2_nor2b_1 _13482_ (.A(net5783),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][5] ),
    .Y(_05447_));
 sg13g2_a21oi_1 _13483_ (.A1(net5783),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][5] ),
    .Y(_05448_),
    .B1(_05447_));
 sg13g2_o21ai_1 _13484_ (.B1(net5709),
    .Y(_05449_),
    .A1(net5739),
    .A2(_05448_));
 sg13g2_a21oi_1 _13485_ (.A1(net5739),
    .A2(_05446_),
    .Y(_05450_),
    .B1(_05449_));
 sg13g2_nor2_1 _13486_ (.A(net5694),
    .B(_05450_),
    .Y(_05451_));
 sg13g2_o21ai_1 _13487_ (.B1(_05451_),
    .Y(_05452_),
    .A1(net5708),
    .A2(_05445_));
 sg13g2_o21ai_1 _13488_ (.B1(_05452_),
    .Y(_00059_),
    .A1(_05438_),
    .A2(_05444_));
 sg13g2_mux4_1 _13489_ (.S0(net5778),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][6] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][6] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][6] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][6] ),
    .S1(net5737),
    .X(_05453_));
 sg13g2_nor2_1 _13490_ (.A(net5706),
    .B(_05453_),
    .Y(_05454_));
 sg13g2_nor2b_1 _13491_ (.A(net5777),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][6] ),
    .Y(_05455_));
 sg13g2_a21oi_1 _13492_ (.A1(net5778),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][6] ),
    .Y(_05456_),
    .B1(_05455_));
 sg13g2_o21ai_1 _13493_ (.B1(net5736),
    .Y(_05457_),
    .A1(net5778),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][6] ));
 sg13g2_a21oi_1 _13494_ (.A1(net5777),
    .A2(_04348_),
    .Y(_05458_),
    .B1(_05457_));
 sg13g2_o21ai_1 _13495_ (.B1(net5706),
    .Y(_05459_),
    .A1(net5736),
    .A2(_05456_));
 sg13g2_o21ai_1 _13496_ (.B1(net5693),
    .Y(_05460_),
    .A1(_05458_),
    .A2(_05459_));
 sg13g2_mux4_1 _13497_ (.S0(net5779),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][6] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][6] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][6] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][6] ),
    .S1(net5737),
    .X(_05461_));
 sg13g2_mux2_1 _13498_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][6] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][6] ),
    .S(net5778),
    .X(_05462_));
 sg13g2_nor2b_1 _13499_ (.A(net5778),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][6] ),
    .Y(_05463_));
 sg13g2_a21oi_1 _13500_ (.A1(net5778),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][6] ),
    .Y(_05464_),
    .B1(_05463_));
 sg13g2_o21ai_1 _13501_ (.B1(net5706),
    .Y(_05465_),
    .A1(net5736),
    .A2(_05464_));
 sg13g2_a21oi_1 _13502_ (.A1(net5736),
    .A2(_05462_),
    .Y(_05466_),
    .B1(_05465_));
 sg13g2_nor2_1 _13503_ (.A(net5693),
    .B(_05466_),
    .Y(_05467_));
 sg13g2_o21ai_1 _13504_ (.B1(_05467_),
    .Y(_05468_),
    .A1(net5706),
    .A2(_05461_));
 sg13g2_o21ai_1 _13505_ (.B1(_05468_),
    .Y(_00060_),
    .A1(_05454_),
    .A2(_05460_));
 sg13g2_mux4_1 _13506_ (.S0(net5803),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][7] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][7] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][7] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][7] ),
    .S1(net5752),
    .X(_05469_));
 sg13g2_nor2_1 _13507_ (.A(net5724),
    .B(_05469_),
    .Y(_05470_));
 sg13g2_nor2b_1 _13508_ (.A(net5804),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][7] ),
    .Y(_05471_));
 sg13g2_a21oi_1 _13509_ (.A1(net5804),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][7] ),
    .Y(_05472_),
    .B1(_05471_));
 sg13g2_o21ai_1 _13510_ (.B1(net5753),
    .Y(_05473_),
    .A1(net5803),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][7] ));
 sg13g2_a21oi_1 _13511_ (.A1(net5802),
    .A2(_04349_),
    .Y(_05474_),
    .B1(_05473_));
 sg13g2_o21ai_1 _13512_ (.B1(net5724),
    .Y(_05475_),
    .A1(net5752),
    .A2(_05472_));
 sg13g2_o21ai_1 _13513_ (.B1(net5700),
    .Y(_05476_),
    .A1(_05474_),
    .A2(_05475_));
 sg13g2_mux4_1 _13514_ (.S0(net5803),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][7] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][7] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][7] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][7] ),
    .S1(net5752),
    .X(_05477_));
 sg13g2_mux2_1 _13515_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][7] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][7] ),
    .S(net5803),
    .X(_05478_));
 sg13g2_nor2b_1 _13516_ (.A(net5803),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][7] ),
    .Y(_05479_));
 sg13g2_a21oi_1 _13517_ (.A1(net5803),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][7] ),
    .Y(_05480_),
    .B1(_05479_));
 sg13g2_o21ai_1 _13518_ (.B1(net5718),
    .Y(_05481_),
    .A1(net5752),
    .A2(_05480_));
 sg13g2_a21oi_1 _13519_ (.A1(net5752),
    .A2(_05478_),
    .Y(_05482_),
    .B1(_05481_));
 sg13g2_nor2_1 _13520_ (.A(net5700),
    .B(_05482_),
    .Y(_05483_));
 sg13g2_o21ai_1 _13521_ (.B1(_05483_),
    .Y(_05484_),
    .A1(net5718),
    .A2(_05477_));
 sg13g2_o21ai_1 _13522_ (.B1(_05484_),
    .Y(_00061_),
    .A1(_05470_),
    .A2(_05476_));
 sg13g2_mux4_1 _13523_ (.S0(net5782),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][8] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][8] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][8] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][8] ),
    .S1(net5739),
    .X(_05485_));
 sg13g2_nor2b_1 _13524_ (.A(net5782),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][8] ),
    .Y(_05486_));
 sg13g2_a21oi_1 _13525_ (.A1(net5783),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][8] ),
    .Y(_05487_),
    .B1(_05486_));
 sg13g2_mux2_1 _13526_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[14][8] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[15][8] ),
    .S(net5782),
    .X(_05488_));
 sg13g2_o21ai_1 _13527_ (.B1(net5709),
    .Y(_05489_),
    .A1(net5740),
    .A2(_05487_));
 sg13g2_a21oi_1 _13528_ (.A1(net5739),
    .A2(_05488_),
    .Y(_05490_),
    .B1(_05489_));
 sg13g2_nor2b_1 _13529_ (.A(_05490_),
    .B_N(net5694),
    .Y(_05491_));
 sg13g2_o21ai_1 _13530_ (.B1(_05491_),
    .Y(_05492_),
    .A1(net5708),
    .A2(_05485_));
 sg13g2_mux2_1 _13531_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[2][8] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[3][8] ),
    .S(net5782),
    .X(_05493_));
 sg13g2_nor2b_1 _13532_ (.A(net5782),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[0][8] ),
    .Y(_05494_));
 sg13g2_a21oi_1 _13533_ (.A1(net5782),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[1][8] ),
    .Y(_05495_),
    .B1(_05494_));
 sg13g2_a21oi_1 _13534_ (.A1(net5739),
    .A2(_05493_),
    .Y(_05496_),
    .B1(net5709));
 sg13g2_o21ai_1 _13535_ (.B1(_05496_),
    .Y(_05497_),
    .A1(net5739),
    .A2(_05495_));
 sg13g2_o21ai_1 _13536_ (.B1(net5739),
    .Y(_05498_),
    .A1(net5782),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[6][8] ));
 sg13g2_a21oi_1 _13537_ (.A1(net5782),
    .A2(_04350_),
    .Y(_05499_),
    .B1(_05498_));
 sg13g2_nor2b_1 _13538_ (.A(net5783),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][8] ),
    .Y(_05500_));
 sg13g2_a21oi_1 _13539_ (.A1(net5783),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][8] ),
    .Y(_05501_),
    .B1(_05500_));
 sg13g2_o21ai_1 _13540_ (.B1(net5709),
    .Y(_05502_),
    .A1(net5739),
    .A2(_05501_));
 sg13g2_o21ai_1 _13541_ (.B1(_05497_),
    .Y(_05503_),
    .A1(_05499_),
    .A2(_05502_));
 sg13g2_o21ai_1 _13542_ (.B1(_05492_),
    .Y(_00062_),
    .A1(net5694),
    .A2(_05503_));
 sg13g2_mux4_1 _13543_ (.S0(net5801),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][9] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][9] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][9] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][9] ),
    .S1(net5755),
    .X(_05504_));
 sg13g2_nor2_1 _13544_ (.A(net5719),
    .B(_05504_),
    .Y(_05505_));
 sg13g2_nor2b_1 _13545_ (.A(net5808),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][9] ),
    .Y(_05506_));
 sg13g2_a21oi_1 _13546_ (.A1(net5808),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][9] ),
    .Y(_05507_),
    .B1(_05506_));
 sg13g2_o21ai_1 _13547_ (.B1(net5755),
    .Y(_05508_),
    .A1(net5808),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][9] ));
 sg13g2_a21oi_1 _13548_ (.A1(net5805),
    .A2(_04351_),
    .Y(_05509_),
    .B1(_05508_));
 sg13g2_o21ai_1 _13549_ (.B1(net5719),
    .Y(_05510_),
    .A1(net5755),
    .A2(_05507_));
 sg13g2_o21ai_1 _13550_ (.B1(net5698),
    .Y(_05511_),
    .A1(_05509_),
    .A2(_05510_));
 sg13g2_mux4_1 _13551_ (.S0(net5802),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][9] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][9] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][9] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][9] ),
    .S1(net5758),
    .X(_05512_));
 sg13g2_mux2_1 _13552_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][9] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][9] ),
    .S(net5810),
    .X(_05513_));
 sg13g2_nor2b_1 _13553_ (.A(net5810),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][9] ),
    .Y(_05514_));
 sg13g2_a21oi_1 _13554_ (.A1(net5810),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][9] ),
    .Y(_05515_),
    .B1(_05514_));
 sg13g2_o21ai_1 _13555_ (.B1(net5721),
    .Y(_05516_),
    .A1(net5758),
    .A2(_05515_));
 sg13g2_a21oi_1 _13556_ (.A1(net5758),
    .A2(_05513_),
    .Y(_05517_),
    .B1(_05516_));
 sg13g2_nor2_1 _13557_ (.A(net5698),
    .B(_05517_),
    .Y(_05518_));
 sg13g2_o21ai_1 _13558_ (.B1(_05518_),
    .Y(_05519_),
    .A1(net5721),
    .A2(_05512_));
 sg13g2_o21ai_1 _13559_ (.B1(_05519_),
    .Y(_00063_),
    .A1(_05505_),
    .A2(_05511_));
 sg13g2_mux4_1 _13560_ (.S0(net5807),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][10] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][10] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][10] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][10] ),
    .S1(net5759),
    .X(_05520_));
 sg13g2_nor2b_1 _13561_ (.A(net5807),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][10] ),
    .Y(_05521_));
 sg13g2_a21oi_1 _13562_ (.A1(net5807),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][10] ),
    .Y(_05522_),
    .B1(_05521_));
 sg13g2_mux2_1 _13563_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[14][10] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[15][10] ),
    .S(net5806),
    .X(_05523_));
 sg13g2_o21ai_1 _13564_ (.B1(net5720),
    .Y(_05524_),
    .A1(net5754),
    .A2(_05522_));
 sg13g2_a21oi_1 _13565_ (.A1(net5754),
    .A2(_05523_),
    .Y(_05525_),
    .B1(_05524_));
 sg13g2_nor2b_1 _13566_ (.A(_05525_),
    .B_N(net5698),
    .Y(_05526_));
 sg13g2_o21ai_1 _13567_ (.B1(_05526_),
    .Y(_05527_),
    .A1(net5719),
    .A2(_05520_));
 sg13g2_mux2_1 _13568_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[2][10] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[3][10] ),
    .S(net5806),
    .X(_05528_));
 sg13g2_nor2b_1 _13569_ (.A(net5806),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[0][10] ),
    .Y(_05529_));
 sg13g2_a21oi_1 _13570_ (.A1(net5806),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[1][10] ),
    .Y(_05530_),
    .B1(_05529_));
 sg13g2_a21oi_1 _13571_ (.A1(net5754),
    .A2(_05528_),
    .Y(_05531_),
    .B1(net5720));
 sg13g2_o21ai_1 _13572_ (.B1(_05531_),
    .Y(_05532_),
    .A1(net5754),
    .A2(_05530_));
 sg13g2_o21ai_1 _13573_ (.B1(net5759),
    .Y(_05533_),
    .A1(net5807),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[6][10] ));
 sg13g2_a21oi_1 _13574_ (.A1(net5807),
    .A2(_04352_),
    .Y(_05534_),
    .B1(_05533_));
 sg13g2_nor2b_1 _13575_ (.A(net5807),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][10] ),
    .Y(_05535_));
 sg13g2_a21oi_1 _13576_ (.A1(net5807),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][10] ),
    .Y(_05536_),
    .B1(_05535_));
 sg13g2_o21ai_1 _13577_ (.B1(net5719),
    .Y(_05537_),
    .A1(net5754),
    .A2(_05536_));
 sg13g2_o21ai_1 _13578_ (.B1(_05532_),
    .Y(_05538_),
    .A1(_05534_),
    .A2(_05537_));
 sg13g2_o21ai_1 _13579_ (.B1(_05527_),
    .Y(_00033_),
    .A1(net5698),
    .A2(_05538_));
 sg13g2_mux4_1 _13580_ (.S0(net5768),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][11] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][11] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][11] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][11] ),
    .S1(net5730),
    .X(_05539_));
 sg13g2_nor2_1 _13581_ (.A(net5705),
    .B(_05539_),
    .Y(_05540_));
 sg13g2_nor2b_1 _13582_ (.A(net5771),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][11] ),
    .Y(_05541_));
 sg13g2_a21oi_1 _13583_ (.A1(net5768),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][11] ),
    .Y(_05542_),
    .B1(_05541_));
 sg13g2_o21ai_1 _13584_ (.B1(net5730),
    .Y(_05543_),
    .A1(net5768),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][11] ));
 sg13g2_a21oi_1 _13585_ (.A1(net5768),
    .A2(_04353_),
    .Y(_05544_),
    .B1(_05543_));
 sg13g2_o21ai_1 _13586_ (.B1(net5705),
    .Y(_05545_),
    .A1(net5730),
    .A2(_05542_));
 sg13g2_o21ai_1 _13587_ (.B1(net5692),
    .Y(_05546_),
    .A1(_05544_),
    .A2(_05545_));
 sg13g2_mux4_1 _13588_ (.S0(net5768),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][11] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][11] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][11] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][11] ),
    .S1(net5730),
    .X(_05547_));
 sg13g2_mux2_1 _13589_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][11] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][11] ),
    .S(net5768),
    .X(_05548_));
 sg13g2_nor2b_1 _13590_ (.A(net5768),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][11] ),
    .Y(_05549_));
 sg13g2_a21oi_1 _13591_ (.A1(net5768),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][11] ),
    .Y(_05550_),
    .B1(_05549_));
 sg13g2_o21ai_1 _13592_ (.B1(net5705),
    .Y(_05551_),
    .A1(net5730),
    .A2(_05550_));
 sg13g2_a21oi_1 _13593_ (.A1(net5730),
    .A2(_05548_),
    .Y(_05552_),
    .B1(_05551_));
 sg13g2_nor2_1 _13594_ (.A(net5692),
    .B(_05552_),
    .Y(_05553_));
 sg13g2_o21ai_1 _13595_ (.B1(_05553_),
    .Y(_05554_),
    .A1(net5705),
    .A2(_05547_));
 sg13g2_o21ai_1 _13596_ (.B1(_05554_),
    .Y(_00034_),
    .A1(_05540_),
    .A2(_05546_));
 sg13g2_mux4_1 _13597_ (.S0(net5764),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][12] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][12] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][12] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][12] ),
    .S1(net5728),
    .X(_05555_));
 sg13g2_nor2_1 _13598_ (.A(net5703),
    .B(_05555_),
    .Y(_05556_));
 sg13g2_nor2b_1 _13599_ (.A(net5763),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][12] ),
    .Y(_05557_));
 sg13g2_a21oi_1 _13600_ (.A1(net5763),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][12] ),
    .Y(_05558_),
    .B1(_05557_));
 sg13g2_o21ai_1 _13601_ (.B1(net5728),
    .Y(_05559_),
    .A1(net5763),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][12] ));
 sg13g2_a21oi_1 _13602_ (.A1(net5763),
    .A2(_04354_),
    .Y(_05560_),
    .B1(_05559_));
 sg13g2_o21ai_1 _13603_ (.B1(net5703),
    .Y(_05561_),
    .A1(net5728),
    .A2(_05558_));
 sg13g2_o21ai_1 _13604_ (.B1(net5691),
    .Y(_05562_),
    .A1(_05560_),
    .A2(_05561_));
 sg13g2_mux4_1 _13605_ (.S0(net5763),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][12] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][12] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][12] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][12] ),
    .S1(net5728),
    .X(_05563_));
 sg13g2_mux2_1 _13606_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][12] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][12] ),
    .S(net5763),
    .X(_05564_));
 sg13g2_nor2b_1 _13607_ (.A(net5763),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][12] ),
    .Y(_05565_));
 sg13g2_a21oi_1 _13608_ (.A1(net5763),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][12] ),
    .Y(_05566_),
    .B1(_05565_));
 sg13g2_o21ai_1 _13609_ (.B1(net5703),
    .Y(_05567_),
    .A1(net5728),
    .A2(_05566_));
 sg13g2_a21oi_1 _13610_ (.A1(net5728),
    .A2(_05564_),
    .Y(_05568_),
    .B1(_05567_));
 sg13g2_nor2_1 _13611_ (.A(net5691),
    .B(_05568_),
    .Y(_05569_));
 sg13g2_o21ai_1 _13612_ (.B1(_05569_),
    .Y(_05570_),
    .A1(net5703),
    .A2(_05563_));
 sg13g2_o21ai_1 _13613_ (.B1(_05570_),
    .Y(_00035_),
    .A1(_05556_),
    .A2(_05562_));
 sg13g2_mux4_1 _13614_ (.S0(net5762),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][13] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][13] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][13] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][13] ),
    .S1(net5727),
    .X(_05571_));
 sg13g2_nor2_1 _13615_ (.A(net5702),
    .B(_05571_),
    .Y(_05572_));
 sg13g2_nor2b_1 _13616_ (.A(net5765),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][13] ),
    .Y(_05573_));
 sg13g2_a21oi_1 _13617_ (.A1(net5762),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][13] ),
    .Y(_05574_),
    .B1(_05573_));
 sg13g2_o21ai_1 _13618_ (.B1(net5727),
    .Y(_05575_),
    .A1(net5762),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][13] ));
 sg13g2_a21oi_1 _13619_ (.A1(net5762),
    .A2(_04355_),
    .Y(_05576_),
    .B1(_05575_));
 sg13g2_o21ai_1 _13620_ (.B1(net5702),
    .Y(_05577_),
    .A1(net5727),
    .A2(_05574_));
 sg13g2_o21ai_1 _13621_ (.B1(net5691),
    .Y(_05578_),
    .A1(_05576_),
    .A2(_05577_));
 sg13g2_mux4_1 _13622_ (.S0(net5761),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][13] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][13] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][13] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][13] ),
    .S1(net5726),
    .X(_05579_));
 sg13g2_mux2_1 _13623_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][13] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][13] ),
    .S(net5762),
    .X(_05580_));
 sg13g2_nor2b_1 _13624_ (.A(net5762),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][13] ),
    .Y(_05581_));
 sg13g2_a21oi_1 _13625_ (.A1(net5762),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][13] ),
    .Y(_05582_),
    .B1(_05581_));
 sg13g2_o21ai_1 _13626_ (.B1(net5702),
    .Y(_05583_),
    .A1(net5726),
    .A2(_05582_));
 sg13g2_a21oi_1 _13627_ (.A1(net5726),
    .A2(_05580_),
    .Y(_05584_),
    .B1(_05583_));
 sg13g2_nor2_1 _13628_ (.A(net5691),
    .B(_05584_),
    .Y(_05585_));
 sg13g2_o21ai_1 _13629_ (.B1(_05585_),
    .Y(_05586_),
    .A1(net5702),
    .A2(_05579_));
 sg13g2_o21ai_1 _13630_ (.B1(_05586_),
    .Y(_00036_),
    .A1(_05572_),
    .A2(_05578_));
 sg13g2_mux4_1 _13631_ (.S0(net5811),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][14] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][14] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][14] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][14] ),
    .S1(net5756),
    .X(_05587_));
 sg13g2_nor2b_1 _13632_ (.A(net5811),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][14] ),
    .Y(_05588_));
 sg13g2_a21oi_1 _13633_ (.A1(net5811),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][14] ),
    .Y(_05589_),
    .B1(_05588_));
 sg13g2_mux2_1 _13634_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[14][14] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[15][14] ),
    .S(net5811),
    .X(_05590_));
 sg13g2_o21ai_1 _13635_ (.B1(net5722),
    .Y(_05591_),
    .A1(net5756),
    .A2(_05589_));
 sg13g2_a21oi_1 _13636_ (.A1(net5756),
    .A2(_05590_),
    .Y(_05592_),
    .B1(_05591_));
 sg13g2_nor2b_1 _13637_ (.A(_05592_),
    .B_N(net5699),
    .Y(_05593_));
 sg13g2_o21ai_1 _13638_ (.B1(_05593_),
    .Y(_05594_),
    .A1(net5721),
    .A2(_05587_));
 sg13g2_mux2_1 _13639_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[2][14] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[3][14] ),
    .S(net5812),
    .X(_05595_));
 sg13g2_nor2b_1 _13640_ (.A(net5812),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[0][14] ),
    .Y(_05596_));
 sg13g2_a21oi_1 _13641_ (.A1(net5812),
    .A2(net3086),
    .Y(_05597_),
    .B1(_05596_));
 sg13g2_a21oi_1 _13642_ (.A1(net5756),
    .A2(_05595_),
    .Y(_05598_),
    .B1(net5722));
 sg13g2_o21ai_1 _13643_ (.B1(_05598_),
    .Y(_05599_),
    .A1(net5756),
    .A2(_05597_));
 sg13g2_o21ai_1 _13644_ (.B1(net5756),
    .Y(_05600_),
    .A1(net5811),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[6][14] ));
 sg13g2_a21oi_1 _13645_ (.A1(net5811),
    .A2(_04356_),
    .Y(_05601_),
    .B1(_05600_));
 sg13g2_nor2b_1 _13646_ (.A(net5811),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][14] ),
    .Y(_05602_));
 sg13g2_a21oi_1 _13647_ (.A1(net5811),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][14] ),
    .Y(_05603_),
    .B1(_05602_));
 sg13g2_o21ai_1 _13648_ (.B1(net5722),
    .Y(_05604_),
    .A1(net5756),
    .A2(_05603_));
 sg13g2_o21ai_1 _13649_ (.B1(_05599_),
    .Y(_05605_),
    .A1(_05601_),
    .A2(_05604_));
 sg13g2_o21ai_1 _13650_ (.B1(_05594_),
    .Y(_00037_),
    .A1(net5698),
    .A2(_05605_));
 sg13g2_mux4_1 _13651_ (.S0(net5769),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][15] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][15] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][15] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][15] ),
    .S1(net5743),
    .X(_05606_));
 sg13g2_nor2_1 _13652_ (.A(net5712),
    .B(_05606_),
    .Y(_05607_));
 sg13g2_nor2b_1 _13653_ (.A(net5786),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][15] ),
    .Y(_05608_));
 sg13g2_a21oi_1 _13654_ (.A1(net5786),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][15] ),
    .Y(_05609_),
    .B1(_05608_));
 sg13g2_o21ai_1 _13655_ (.B1(net5730),
    .Y(_05610_),
    .A1(net5769),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][15] ));
 sg13g2_a21oi_1 _13656_ (.A1(net5786),
    .A2(_04357_),
    .Y(_05611_),
    .B1(_05610_));
 sg13g2_o21ai_1 _13657_ (.B1(net5712),
    .Y(_05612_),
    .A1(net5742),
    .A2(_05609_));
 sg13g2_o21ai_1 _13658_ (.B1(net5697),
    .Y(_05613_),
    .A1(_05611_),
    .A2(_05612_));
 sg13g2_mux4_1 _13659_ (.S0(net5769),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][15] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][15] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][15] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][15] ),
    .S1(net5742),
    .X(_05614_));
 sg13g2_mux2_1 _13660_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][15] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][15] ),
    .S(net5785),
    .X(_05615_));
 sg13g2_nor2b_1 _13661_ (.A(net5785),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][15] ),
    .Y(_05616_));
 sg13g2_a21oi_1 _13662_ (.A1(net5785),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][15] ),
    .Y(_05617_),
    .B1(_05616_));
 sg13g2_o21ai_1 _13663_ (.B1(net5712),
    .Y(_05618_),
    .A1(net5742),
    .A2(_05617_));
 sg13g2_a21oi_1 _13664_ (.A1(net5742),
    .A2(_05615_),
    .Y(_05619_),
    .B1(_05618_));
 sg13g2_nor2_1 _13665_ (.A(net5697),
    .B(_05619_),
    .Y(_05620_));
 sg13g2_o21ai_1 _13666_ (.B1(_05620_),
    .Y(_05621_),
    .A1(net5712),
    .A2(_05614_));
 sg13g2_o21ai_1 _13667_ (.B1(_05621_),
    .Y(_00038_),
    .A1(_05607_),
    .A2(_05613_));
 sg13g2_mux4_1 _13668_ (.S0(net5809),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][16] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][16] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][16] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][16] ),
    .S1(net5756),
    .X(_05622_));
 sg13g2_nor2b_1 _13669_ (.A(net5809),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][16] ),
    .Y(_05623_));
 sg13g2_a21oi_1 _13670_ (.A1(net5810),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][16] ),
    .Y(_05624_),
    .B1(_05623_));
 sg13g2_mux2_1 _13671_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[14][16] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[15][16] ),
    .S(net5810),
    .X(_05625_));
 sg13g2_o21ai_1 _13672_ (.B1(net5721),
    .Y(_05626_),
    .A1(net5758),
    .A2(_05624_));
 sg13g2_a21oi_1 _13673_ (.A1(net5757),
    .A2(_05625_),
    .Y(_05627_),
    .B1(_05626_));
 sg13g2_nor2b_1 _13674_ (.A(_05627_),
    .B_N(net5699),
    .Y(_05628_));
 sg13g2_o21ai_1 _13675_ (.B1(_05628_),
    .Y(_05629_),
    .A1(net5721),
    .A2(_05622_));
 sg13g2_mux2_1 _13676_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[2][16] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[3][16] ),
    .S(net5813),
    .X(_05630_));
 sg13g2_nor2b_1 _13677_ (.A(net5812),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[0][16] ),
    .Y(_05631_));
 sg13g2_a21oi_1 _13678_ (.A1(net5812),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[1][16] ),
    .Y(_05632_),
    .B1(_05631_));
 sg13g2_a21oi_1 _13679_ (.A1(net5757),
    .A2(_05630_),
    .Y(_05633_),
    .B1(net5722));
 sg13g2_o21ai_1 _13680_ (.B1(_05633_),
    .Y(_05634_),
    .A1(net5757),
    .A2(_05632_));
 sg13g2_o21ai_1 _13681_ (.B1(net5757),
    .Y(_05635_),
    .A1(net5813),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[6][16] ));
 sg13g2_a21oi_1 _13682_ (.A1(net5813),
    .A2(_04358_),
    .Y(_05636_),
    .B1(_05635_));
 sg13g2_nor2b_1 _13683_ (.A(net5812),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][16] ),
    .Y(_05637_));
 sg13g2_a21oi_1 _13684_ (.A1(net5812),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][16] ),
    .Y(_05638_),
    .B1(_05637_));
 sg13g2_o21ai_1 _13685_ (.B1(net5721),
    .Y(_05639_),
    .A1(net5757),
    .A2(_05638_));
 sg13g2_o21ai_1 _13686_ (.B1(_05634_),
    .Y(_05640_),
    .A1(_05636_),
    .A2(_05639_));
 sg13g2_o21ai_1 _13687_ (.B1(_05629_),
    .Y(_00039_),
    .A1(net5699),
    .A2(_05640_));
 sg13g2_mux4_1 _13688_ (.S0(net5790),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][17] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][17] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][17] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][17] ),
    .S1(net5744),
    .X(_05641_));
 sg13g2_nor2_1 _13689_ (.A(net5725),
    .B(_05641_),
    .Y(_05642_));
 sg13g2_nor2b_1 _13690_ (.A(net5788),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][17] ),
    .Y(_05643_));
 sg13g2_a21oi_1 _13691_ (.A1(net5788),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][17] ),
    .Y(_05644_),
    .B1(_05643_));
 sg13g2_o21ai_1 _13692_ (.B1(net5751),
    .Y(_05645_),
    .A1(net5788),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][17] ));
 sg13g2_a21oi_1 _13693_ (.A1(net5788),
    .A2(_04359_),
    .Y(_05646_),
    .B1(_05645_));
 sg13g2_o21ai_1 _13694_ (.B1(net5713),
    .Y(_05647_),
    .A1(net5751),
    .A2(_05644_));
 sg13g2_o21ai_1 _13695_ (.B1(net5697),
    .Y(_05648_),
    .A1(_05646_),
    .A2(_05647_));
 sg13g2_mux4_1 _13696_ (.S0(net5788),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][17] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][17] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][17] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][17] ),
    .S1(net5744),
    .X(_05649_));
 sg13g2_mux2_1 _13697_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][17] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][17] ),
    .S(net5788),
    .X(_05650_));
 sg13g2_nor2b_1 _13698_ (.A(net5788),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][17] ),
    .Y(_05651_));
 sg13g2_a21oi_1 _13699_ (.A1(net5788),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][17] ),
    .Y(_05652_),
    .B1(_05651_));
 sg13g2_o21ai_1 _13700_ (.B1(net5713),
    .Y(_05653_),
    .A1(net5744),
    .A2(_05652_));
 sg13g2_a21oi_1 _13701_ (.A1(net5744),
    .A2(_05650_),
    .Y(_05654_),
    .B1(_05653_));
 sg13g2_nor2_1 _13702_ (.A(net5697),
    .B(_05654_),
    .Y(_05655_));
 sg13g2_o21ai_1 _13703_ (.B1(_05655_),
    .Y(_05656_),
    .A1(net5713),
    .A2(_05649_));
 sg13g2_o21ai_1 _13704_ (.B1(_05656_),
    .Y(_00040_),
    .A1(_05642_),
    .A2(_05648_));
 sg13g2_mux4_1 _13705_ (.S0(net5767),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][18] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][18] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][18] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][18] ),
    .S1(net5733),
    .X(_05657_));
 sg13g2_nor2_1 _13706_ (.A(net5704),
    .B(_05657_),
    .Y(_05658_));
 sg13g2_nor2b_1 _13707_ (.A(net5772),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][18] ),
    .Y(_05659_));
 sg13g2_a21oi_1 _13708_ (.A1(net5772),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][18] ),
    .Y(_05660_),
    .B1(_05659_));
 sg13g2_o21ai_1 _13709_ (.B1(net5732),
    .Y(_05661_),
    .A1(net5772),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][18] ));
 sg13g2_a21oi_1 _13710_ (.A1(net5772),
    .A2(_04360_),
    .Y(_05662_),
    .B1(_05661_));
 sg13g2_o21ai_1 _13711_ (.B1(net5704),
    .Y(_05663_),
    .A1(net5733),
    .A2(_05660_));
 sg13g2_o21ai_1 _13712_ (.B1(net5692),
    .Y(_05664_),
    .A1(_05662_),
    .A2(_05663_));
 sg13g2_mux4_1 _13713_ (.S0(net5772),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][18] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][18] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][18] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][18] ),
    .S1(net5732),
    .X(_05665_));
 sg13g2_mux2_1 _13714_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][18] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][18] ),
    .S(net5764),
    .X(_05666_));
 sg13g2_nor2b_1 _13715_ (.A(net5764),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][18] ),
    .Y(_05667_));
 sg13g2_a21oi_1 _13716_ (.A1(net5764),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][18] ),
    .Y(_05668_),
    .B1(_05667_));
 sg13g2_o21ai_1 _13717_ (.B1(net5703),
    .Y(_05669_),
    .A1(net5729),
    .A2(_05668_));
 sg13g2_a21oi_1 _13718_ (.A1(net5729),
    .A2(_05666_),
    .Y(_05670_),
    .B1(_05669_));
 sg13g2_nor2_1 _13719_ (.A(net5691),
    .B(_05670_),
    .Y(_05671_));
 sg13g2_o21ai_1 _13720_ (.B1(_05671_),
    .Y(_05672_),
    .A1(net5711),
    .A2(_05665_));
 sg13g2_o21ai_1 _13721_ (.B1(_05672_),
    .Y(_00041_),
    .A1(_05658_),
    .A2(_05664_));
 sg13g2_mux4_1 _13722_ (.S0(net5770),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][19] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][19] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][19] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][19] ),
    .S1(net5731),
    .X(_05673_));
 sg13g2_nor2_1 _13723_ (.A(net5705),
    .B(_05673_),
    .Y(_05674_));
 sg13g2_nor2b_1 _13724_ (.A(net5769),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][19] ),
    .Y(_05675_));
 sg13g2_a21oi_1 _13725_ (.A1(net5770),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][19] ),
    .Y(_05676_),
    .B1(_05675_));
 sg13g2_o21ai_1 _13726_ (.B1(net5731),
    .Y(_05677_),
    .A1(net5770),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][19] ));
 sg13g2_a21oi_1 _13727_ (.A1(net5770),
    .A2(_04361_),
    .Y(_05678_),
    .B1(_05677_));
 sg13g2_o21ai_1 _13728_ (.B1(net5705),
    .Y(_05679_),
    .A1(net5731),
    .A2(_05676_));
 sg13g2_o21ai_1 _13729_ (.B1(net5692),
    .Y(_05680_),
    .A1(_05678_),
    .A2(_05679_));
 sg13g2_mux4_1 _13730_ (.S0(net5769),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][19] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][19] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][19] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][19] ),
    .S1(net5730),
    .X(_05681_));
 sg13g2_mux2_1 _13731_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][19] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][19] ),
    .S(net5769),
    .X(_05682_));
 sg13g2_nor2b_1 _13732_ (.A(net5769),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][19] ),
    .Y(_05683_));
 sg13g2_a21oi_1 _13733_ (.A1(net5769),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][19] ),
    .Y(_05684_),
    .B1(_05683_));
 sg13g2_o21ai_1 _13734_ (.B1(net5705),
    .Y(_05685_),
    .A1(net5731),
    .A2(_05684_));
 sg13g2_a21oi_1 _13735_ (.A1(net5731),
    .A2(_05682_),
    .Y(_05686_),
    .B1(_05685_));
 sg13g2_nor2_1 _13736_ (.A(net5692),
    .B(_05686_),
    .Y(_05687_));
 sg13g2_o21ai_1 _13737_ (.B1(_05687_),
    .Y(_05688_),
    .A1(net5705),
    .A2(_05681_));
 sg13g2_o21ai_1 _13738_ (.B1(_05688_),
    .Y(_00042_),
    .A1(_05674_),
    .A2(_05680_));
 sg13g2_mux4_1 _13739_ (.S0(net5797),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][20] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][20] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][20] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][20] ),
    .S1(net5750),
    .X(_05689_));
 sg13g2_nor2b_1 _13740_ (.A(net5796),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][20] ),
    .Y(_05690_));
 sg13g2_a21oi_1 _13741_ (.A1(net5796),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][20] ),
    .Y(_05691_),
    .B1(_05690_));
 sg13g2_mux2_1 _13742_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[14][20] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[15][20] ),
    .S(net5796),
    .X(_05692_));
 sg13g2_o21ai_1 _13743_ (.B1(net5716),
    .Y(_05693_),
    .A1(net5749),
    .A2(_05691_));
 sg13g2_a21oi_1 _13744_ (.A1(net5749),
    .A2(_05692_),
    .Y(_05694_),
    .B1(_05693_));
 sg13g2_nor2b_1 _13745_ (.A(_05694_),
    .B_N(net5696),
    .Y(_05695_));
 sg13g2_o21ai_1 _13746_ (.B1(_05695_),
    .Y(_05696_),
    .A1(net5717),
    .A2(_05689_));
 sg13g2_mux2_1 _13747_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[2][20] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[3][20] ),
    .S(net5798),
    .X(_05697_));
 sg13g2_nor2b_1 _13748_ (.A(net5798),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[0][20] ),
    .Y(_05698_));
 sg13g2_a21oi_1 _13749_ (.A1(net5798),
    .A2(net2722),
    .Y(_05699_),
    .B1(_05698_));
 sg13g2_a21oi_1 _13750_ (.A1(net5748),
    .A2(_05697_),
    .Y(_05700_),
    .B1(net5716));
 sg13g2_o21ai_1 _13751_ (.B1(_05700_),
    .Y(_05701_),
    .A1(net5748),
    .A2(_05699_));
 sg13g2_o21ai_1 _13752_ (.B1(net5748),
    .Y(_05702_),
    .A1(net5798),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[6][20] ));
 sg13g2_a21oi_1 _13753_ (.A1(net5798),
    .A2(_04362_),
    .Y(_05703_),
    .B1(_05702_));
 sg13g2_nor2b_1 _13754_ (.A(net5798),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][20] ),
    .Y(_05704_));
 sg13g2_a21oi_1 _13755_ (.A1(net5798),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][20] ),
    .Y(_05705_),
    .B1(_05704_));
 sg13g2_o21ai_1 _13756_ (.B1(net5716),
    .Y(_05706_),
    .A1(net5748),
    .A2(_05705_));
 sg13g2_o21ai_1 _13757_ (.B1(_05701_),
    .Y(_05707_),
    .A1(_05703_),
    .A2(_05706_));
 sg13g2_o21ai_1 _13758_ (.B1(_05696_),
    .Y(_00044_),
    .A1(net5696),
    .A2(_05707_));
 sg13g2_mux4_1 _13759_ (.S0(net5787),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][21] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][21] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][21] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][21] ),
    .S1(net5743),
    .X(_05708_));
 sg13g2_nor2_1 _13760_ (.A(net5713),
    .B(_05708_),
    .Y(_05709_));
 sg13g2_nor2b_1 _13761_ (.A(net5787),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][21] ),
    .Y(_05710_));
 sg13g2_a21oi_1 _13762_ (.A1(net5787),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][21] ),
    .Y(_05711_),
    .B1(_05710_));
 sg13g2_o21ai_1 _13763_ (.B1(net5743),
    .Y(_05712_),
    .A1(net5787),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][21] ));
 sg13g2_a21oi_1 _13764_ (.A1(net5787),
    .A2(_04363_),
    .Y(_05713_),
    .B1(_05712_));
 sg13g2_o21ai_1 _13765_ (.B1(net5713),
    .Y(_05714_),
    .A1(net5743),
    .A2(_05711_));
 sg13g2_o21ai_1 _13766_ (.B1(net5697),
    .Y(_05715_),
    .A1(_05713_),
    .A2(_05714_));
 sg13g2_mux4_1 _13767_ (.S0(net5787),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][21] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][21] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][21] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][21] ),
    .S1(net5743),
    .X(_05716_));
 sg13g2_mux2_1 _13768_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][21] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][21] ),
    .S(net5791),
    .X(_05717_));
 sg13g2_nor2b_1 _13769_ (.A(net5790),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][21] ),
    .Y(_05718_));
 sg13g2_a21oi_1 _13770_ (.A1(net5791),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][21] ),
    .Y(_05719_),
    .B1(_05718_));
 sg13g2_o21ai_1 _13771_ (.B1(net5714),
    .Y(_05720_),
    .A1(net5743),
    .A2(_05719_));
 sg13g2_a21oi_1 _13772_ (.A1(net5747),
    .A2(_05717_),
    .Y(_05721_),
    .B1(_05720_));
 sg13g2_nor2_1 _13773_ (.A(net5695),
    .B(_05721_),
    .Y(_05722_));
 sg13g2_o21ai_1 _13774_ (.B1(_05722_),
    .Y(_05723_),
    .A1(net5712),
    .A2(_05716_));
 sg13g2_o21ai_1 _13775_ (.B1(_05723_),
    .Y(_00045_),
    .A1(_05709_),
    .A2(_05715_));
 sg13g2_mux4_1 _13776_ (.S0(net5798),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][22] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][22] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][22] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][22] ),
    .S1(net5745),
    .X(_05724_));
 sg13g2_nor2b_1 _13777_ (.A(net5793),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][22] ),
    .Y(_05725_));
 sg13g2_a21oi_1 _13778_ (.A1(net5794),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][22] ),
    .Y(_05726_),
    .B1(_05725_));
 sg13g2_mux2_1 _13779_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[14][22] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[15][22] ),
    .S(net5794),
    .X(_05727_));
 sg13g2_o21ai_1 _13780_ (.B1(net5714),
    .Y(_05728_),
    .A1(net5746),
    .A2(_05726_));
 sg13g2_a21oi_1 _13781_ (.A1(net5746),
    .A2(_05727_),
    .Y(_05729_),
    .B1(_05728_));
 sg13g2_nor2b_1 _13782_ (.A(_05729_),
    .B_N(net5695),
    .Y(_05730_));
 sg13g2_o21ai_1 _13783_ (.B1(_05730_),
    .Y(_05731_),
    .A1(net5715),
    .A2(_05724_));
 sg13g2_mux2_1 _13784_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[2][22] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[3][22] ),
    .S(net5793),
    .X(_05732_));
 sg13g2_nor2b_1 _13785_ (.A(net5793),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[0][22] ),
    .Y(_05733_));
 sg13g2_a21oi_1 _13786_ (.A1(net5793),
    .A2(net2904),
    .Y(_05734_),
    .B1(_05733_));
 sg13g2_a21oi_1 _13787_ (.A1(net5745),
    .A2(_05732_),
    .Y(_05735_),
    .B1(net5714));
 sg13g2_o21ai_1 _13788_ (.B1(_05735_),
    .Y(_05736_),
    .A1(net5746),
    .A2(_05734_));
 sg13g2_o21ai_1 _13789_ (.B1(net5746),
    .Y(_05737_),
    .A1(net5793),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[6][22] ));
 sg13g2_a21oi_1 _13790_ (.A1(net5793),
    .A2(_04364_),
    .Y(_05738_),
    .B1(_05737_));
 sg13g2_nor2b_1 _13791_ (.A(net5793),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][22] ),
    .Y(_05739_));
 sg13g2_a21oi_1 _13792_ (.A1(net5793),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][22] ),
    .Y(_05740_),
    .B1(_05739_));
 sg13g2_o21ai_1 _13793_ (.B1(net5714),
    .Y(_05741_),
    .A1(net5746),
    .A2(_05740_));
 sg13g2_o21ai_1 _13794_ (.B1(_05736_),
    .Y(_05742_),
    .A1(_05738_),
    .A2(_05741_));
 sg13g2_o21ai_1 _13795_ (.B1(_05731_),
    .Y(_00046_),
    .A1(net5695),
    .A2(_05742_));
 sg13g2_mux4_1 _13796_ (.S0(net5792),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][23] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][23] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][23] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][23] ),
    .S1(net5745),
    .X(_05743_));
 sg13g2_nor2_1 _13797_ (.A(net5715),
    .B(_05743_),
    .Y(_05744_));
 sg13g2_nor2b_1 _13798_ (.A(net5792),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][23] ),
    .Y(_05745_));
 sg13g2_a21oi_1 _13799_ (.A1(net5792),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][23] ),
    .Y(_05746_),
    .B1(_05745_));
 sg13g2_o21ai_1 _13800_ (.B1(net5745),
    .Y(_05747_),
    .A1(net5792),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][23] ));
 sg13g2_a21oi_1 _13801_ (.A1(net5792),
    .A2(_04365_),
    .Y(_05748_),
    .B1(_05747_));
 sg13g2_o21ai_1 _13802_ (.B1(net5715),
    .Y(_05749_),
    .A1(net5745),
    .A2(_05746_));
 sg13g2_o21ai_1 _13803_ (.B1(net5695),
    .Y(_05750_),
    .A1(_05748_),
    .A2(_05749_));
 sg13g2_mux4_1 _13804_ (.S0(net5792),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][23] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][23] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][23] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][23] ),
    .S1(net5745),
    .X(_05751_));
 sg13g2_mux2_1 _13805_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][23] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][23] ),
    .S(net5792),
    .X(_05752_));
 sg13g2_nor2b_1 _13806_ (.A(net5792),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][23] ),
    .Y(_05753_));
 sg13g2_a21oi_1 _13807_ (.A1(net5794),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][23] ),
    .Y(_05754_),
    .B1(_05753_));
 sg13g2_o21ai_1 _13808_ (.B1(net5715),
    .Y(_05755_),
    .A1(net5745),
    .A2(_05754_));
 sg13g2_a21oi_1 _13809_ (.A1(net5745),
    .A2(_05752_),
    .Y(_05756_),
    .B1(_05755_));
 sg13g2_nor2_1 _13810_ (.A(net5695),
    .B(_05756_),
    .Y(_05757_));
 sg13g2_o21ai_1 _13811_ (.B1(_05757_),
    .Y(_05758_),
    .A1(net5715),
    .A2(_05751_));
 sg13g2_o21ai_1 _13812_ (.B1(_05758_),
    .Y(_00047_),
    .A1(_05744_),
    .A2(_05750_));
 sg13g2_mux4_1 _13813_ (.S0(net5799),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][24] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][24] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][24] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][24] ),
    .S1(net5747),
    .X(_05759_));
 sg13g2_nor2_1 _13814_ (.A(net5714),
    .B(_05759_),
    .Y(_05760_));
 sg13g2_nor2b_1 _13815_ (.A(net5791),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][24] ),
    .Y(_05761_));
 sg13g2_a21oi_1 _13816_ (.A1(net5791),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][24] ),
    .Y(_05762_),
    .B1(_05761_));
 sg13g2_o21ai_1 _13817_ (.B1(net5747),
    .Y(_05763_),
    .A1(net5791),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][24] ));
 sg13g2_a21oi_1 _13818_ (.A1(net5791),
    .A2(_04366_),
    .Y(_05764_),
    .B1(_05763_));
 sg13g2_o21ai_1 _13819_ (.B1(net5714),
    .Y(_05765_),
    .A1(net5747),
    .A2(_05762_));
 sg13g2_o21ai_1 _13820_ (.B1(net5695),
    .Y(_05766_),
    .A1(_05764_),
    .A2(_05765_));
 sg13g2_mux4_1 _13821_ (.S0(net5791),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][24] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][24] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][24] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][24] ),
    .S1(net5747),
    .X(_05767_));
 sg13g2_mux2_1 _13822_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][24] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][24] ),
    .S(net5795),
    .X(_05768_));
 sg13g2_nor2b_1 _13823_ (.A(net5795),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][24] ),
    .Y(_05769_));
 sg13g2_a21oi_1 _13824_ (.A1(net5791),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][24] ),
    .Y(_05770_),
    .B1(_05769_));
 sg13g2_o21ai_1 _13825_ (.B1(net5714),
    .Y(_05771_),
    .A1(net5747),
    .A2(_05770_));
 sg13g2_a21oi_1 _13826_ (.A1(net5747),
    .A2(_05768_),
    .Y(_05772_),
    .B1(_05771_));
 sg13g2_nor2_1 _13827_ (.A(net5695),
    .B(_05772_),
    .Y(_05773_));
 sg13g2_o21ai_1 _13828_ (.B1(_05773_),
    .Y(_05774_),
    .A1(net5714),
    .A2(_05767_));
 sg13g2_o21ai_1 _13829_ (.B1(_05774_),
    .Y(_00048_),
    .A1(_05760_),
    .A2(_05766_));
 sg13g2_mux4_1 _13830_ (.S0(net5786),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][25] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][25] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][25] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][25] ),
    .S1(net5743),
    .X(_05775_));
 sg13g2_nor2_1 _13831_ (.A(net5712),
    .B(_05775_),
    .Y(_05776_));
 sg13g2_nor2b_1 _13832_ (.A(net5785),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][25] ),
    .Y(_05777_));
 sg13g2_a21oi_1 _13833_ (.A1(net5785),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][25] ),
    .Y(_05778_),
    .B1(_05777_));
 sg13g2_o21ai_1 _13834_ (.B1(net5742),
    .Y(_05779_),
    .A1(net5786),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][25] ));
 sg13g2_a21oi_1 _13835_ (.A1(net5786),
    .A2(_04367_),
    .Y(_05780_),
    .B1(_05779_));
 sg13g2_o21ai_1 _13836_ (.B1(net5712),
    .Y(_05781_),
    .A1(net5742),
    .A2(_05778_));
 sg13g2_o21ai_1 _13837_ (.B1(net5697),
    .Y(_05782_),
    .A1(_05780_),
    .A2(_05781_));
 sg13g2_mux4_1 _13838_ (.S0(net5785),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][25] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][25] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][25] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][25] ),
    .S1(net5742),
    .X(_05783_));
 sg13g2_mux2_1 _13839_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][25] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][25] ),
    .S(net5790),
    .X(_05784_));
 sg13g2_nor2b_1 _13840_ (.A(net5785),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][25] ),
    .Y(_05785_));
 sg13g2_a21oi_1 _13841_ (.A1(net5785),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][25] ),
    .Y(_05786_),
    .B1(_05785_));
 sg13g2_o21ai_1 _13842_ (.B1(net5713),
    .Y(_05787_),
    .A1(net5742),
    .A2(_05786_));
 sg13g2_a21oi_1 _13843_ (.A1(net5744),
    .A2(_05784_),
    .Y(_05788_),
    .B1(_05787_));
 sg13g2_nor2_1 _13844_ (.A(net5697),
    .B(_05788_),
    .Y(_05789_));
 sg13g2_o21ai_1 _13845_ (.B1(_05789_),
    .Y(_05790_),
    .A1(net5712),
    .A2(_05783_));
 sg13g2_o21ai_1 _13846_ (.B1(_05790_),
    .Y(_00049_),
    .A1(_05776_),
    .A2(_05782_));
 sg13g2_mux4_1 _13847_ (.S0(net5806),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][26] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][26] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][26] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][26] ),
    .S1(net5754),
    .X(_05791_));
 sg13g2_nor2b_1 _13848_ (.A(net5806),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][26] ),
    .Y(_05792_));
 sg13g2_a21oi_1 _13849_ (.A1(net5806),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][26] ),
    .Y(_05793_),
    .B1(_05792_));
 sg13g2_mux2_1 _13850_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[14][26] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[15][26] ),
    .S(net5806),
    .X(_05794_));
 sg13g2_o21ai_1 _13851_ (.B1(net5720),
    .Y(_05795_),
    .A1(net5754),
    .A2(_05793_));
 sg13g2_a21oi_1 _13852_ (.A1(net5754),
    .A2(_05794_),
    .Y(_05796_),
    .B1(_05795_));
 sg13g2_nor2b_1 _13853_ (.A(_05796_),
    .B_N(net5698),
    .Y(_05797_));
 sg13g2_o21ai_1 _13854_ (.B1(_05797_),
    .Y(_05798_),
    .A1(net5720),
    .A2(_05791_));
 sg13g2_mux2_1 _13855_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[2][26] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[3][26] ),
    .S(net5797),
    .X(_05799_));
 sg13g2_nor2b_1 _13856_ (.A(net5796),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[0][26] ),
    .Y(_05800_));
 sg13g2_a21oi_1 _13857_ (.A1(net5796),
    .A2(net2801),
    .Y(_05801_),
    .B1(_05800_));
 sg13g2_a21oi_1 _13858_ (.A1(net5748),
    .A2(_05799_),
    .Y(_05802_),
    .B1(net5716));
 sg13g2_o21ai_1 _13859_ (.B1(_05802_),
    .Y(_05803_),
    .A1(net5748),
    .A2(_05801_));
 sg13g2_o21ai_1 _13860_ (.B1(net5748),
    .Y(_05804_),
    .A1(net5797),
    .A2(net2827));
 sg13g2_a21oi_1 _13861_ (.A1(net5796),
    .A2(_04368_),
    .Y(_05805_),
    .B1(_05804_));
 sg13g2_nor2b_1 _13862_ (.A(net5796),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][26] ),
    .Y(_05806_));
 sg13g2_a21oi_1 _13863_ (.A1(net5796),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][26] ),
    .Y(_05807_),
    .B1(_05806_));
 sg13g2_o21ai_1 _13864_ (.B1(net5716),
    .Y(_05808_),
    .A1(net5748),
    .A2(_05807_));
 sg13g2_o21ai_1 _13865_ (.B1(_05803_),
    .Y(_05809_),
    .A1(_05805_),
    .A2(_05808_));
 sg13g2_o21ai_1 _13866_ (.B1(_05798_),
    .Y(_00050_),
    .A1(net5695),
    .A2(_05809_));
 sg13g2_mux4_1 _13867_ (.S0(net5773),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][27] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][27] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][27] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][27] ),
    .S1(net5734),
    .X(_05810_));
 sg13g2_nor2_1 _13868_ (.A(net5707),
    .B(_05810_),
    .Y(_05811_));
 sg13g2_nor2b_1 _13869_ (.A(net5773),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][27] ),
    .Y(_05812_));
 sg13g2_a21oi_1 _13870_ (.A1(net5773),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][27] ),
    .Y(_05813_),
    .B1(_05812_));
 sg13g2_o21ai_1 _13871_ (.B1(net5734),
    .Y(_05814_),
    .A1(net5773),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][27] ));
 sg13g2_a21oi_1 _13872_ (.A1(net5773),
    .A2(_04369_),
    .Y(_05815_),
    .B1(_05814_));
 sg13g2_o21ai_1 _13873_ (.B1(net5707),
    .Y(_05816_),
    .A1(net5734),
    .A2(_05813_));
 sg13g2_o21ai_1 _13874_ (.B1(net5693),
    .Y(_05817_),
    .A1(_05815_),
    .A2(_05816_));
 sg13g2_mux4_1 _13875_ (.S0(net5774),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][27] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][27] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][27] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][27] ),
    .S1(net5734),
    .X(_05818_));
 sg13g2_mux2_1 _13876_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][27] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][27] ),
    .S(net5773),
    .X(_05819_));
 sg13g2_nor2b_1 _13877_ (.A(net5773),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][27] ),
    .Y(_05820_));
 sg13g2_a21oi_1 _13878_ (.A1(net5773),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][27] ),
    .Y(_05821_),
    .B1(_05820_));
 sg13g2_o21ai_1 _13879_ (.B1(net5707),
    .Y(_05822_),
    .A1(net5734),
    .A2(_05821_));
 sg13g2_a21oi_1 _13880_ (.A1(net5734),
    .A2(_05819_),
    .Y(_05823_),
    .B1(_05822_));
 sg13g2_nor2_1 _13881_ (.A(net5693),
    .B(_05823_),
    .Y(_05824_));
 sg13g2_o21ai_1 _13882_ (.B1(_05824_),
    .Y(_05825_),
    .A1(net5707),
    .A2(_05818_));
 sg13g2_o21ai_1 _13883_ (.B1(_05825_),
    .Y(_00051_),
    .A1(_05811_),
    .A2(_05817_));
 sg13g2_mux4_1 _13884_ (.S0(net5804),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][28] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][28] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][28] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][28] ),
    .S1(net5753),
    .X(_05826_));
 sg13g2_nor2b_1 _13885_ (.A(net5803),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][28] ),
    .Y(_05827_));
 sg13g2_a21oi_1 _13886_ (.A1(net5802),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][28] ),
    .Y(_05828_),
    .B1(_05827_));
 sg13g2_mux2_1 _13887_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[14][28] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[15][28] ),
    .S(net5802),
    .X(_05829_));
 sg13g2_o21ai_1 _13888_ (.B1(net5718),
    .Y(_05830_),
    .A1(net5752),
    .A2(_05828_));
 sg13g2_a21oi_1 _13889_ (.A1(net5760),
    .A2(_05829_),
    .Y(_05831_),
    .B1(_05830_));
 sg13g2_nor2b_1 _13890_ (.A(_05831_),
    .B_N(net5700),
    .Y(_05832_));
 sg13g2_o21ai_1 _13891_ (.B1(_05832_),
    .Y(_05833_),
    .A1(net5718),
    .A2(_05826_));
 sg13g2_mux2_1 _13892_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[2][28] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[3][28] ),
    .S(net5802),
    .X(_05834_));
 sg13g2_nor2b_1 _13893_ (.A(net5804),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[0][28] ),
    .Y(_05835_));
 sg13g2_a21oi_1 _13894_ (.A1(net5801),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[1][28] ),
    .Y(_05836_),
    .B1(_05835_));
 sg13g2_a21oi_1 _13895_ (.A1(net5753),
    .A2(_05834_),
    .Y(_05837_),
    .B1(net5718));
 sg13g2_o21ai_1 _13896_ (.B1(_05837_),
    .Y(_05838_),
    .A1(net5753),
    .A2(_05836_));
 sg13g2_o21ai_1 _13897_ (.B1(net5753),
    .Y(_05839_),
    .A1(net5801),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[6][28] ));
 sg13g2_a21oi_1 _13898_ (.A1(net5801),
    .A2(_04370_),
    .Y(_05840_),
    .B1(_05839_));
 sg13g2_nor2b_1 _13899_ (.A(net5801),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][28] ),
    .Y(_05841_));
 sg13g2_a21oi_1 _13900_ (.A1(net5801),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][28] ),
    .Y(_05842_),
    .B1(_05841_));
 sg13g2_o21ai_1 _13901_ (.B1(net5718),
    .Y(_05843_),
    .A1(net5753),
    .A2(_05842_));
 sg13g2_o21ai_1 _13902_ (.B1(_05838_),
    .Y(_05844_),
    .A1(_05840_),
    .A2(_05843_));
 sg13g2_o21ai_1 _13903_ (.B1(_05833_),
    .Y(_00052_),
    .A1(net5700),
    .A2(_05844_));
 sg13g2_mux4_1 _13904_ (.S0(net5801),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][29] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][29] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][29] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][29] ),
    .S1(net5753),
    .X(_05845_));
 sg13g2_nor2_1 _13905_ (.A(net5719),
    .B(_05845_),
    .Y(_05846_));
 sg13g2_nor2b_1 _13906_ (.A(net5805),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][29] ),
    .Y(_05847_));
 sg13g2_a21oi_1 _13907_ (.A1(net5805),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][29] ),
    .Y(_05848_),
    .B1(_05847_));
 sg13g2_o21ai_1 _13908_ (.B1(net5755),
    .Y(_05849_),
    .A1(net5805),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][29] ));
 sg13g2_a21oi_1 _13909_ (.A1(net5805),
    .A2(_04371_),
    .Y(_05850_),
    .B1(_05849_));
 sg13g2_o21ai_1 _13910_ (.B1(net5719),
    .Y(_05851_),
    .A1(net5755),
    .A2(_05848_));
 sg13g2_o21ai_1 _13911_ (.B1(net5698),
    .Y(_05852_),
    .A1(_05850_),
    .A2(_05851_));
 sg13g2_mux4_1 _13912_ (.S0(net5801),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][29] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][29] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][29] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][29] ),
    .S1(net5755),
    .X(_05853_));
 sg13g2_mux2_1 _13913_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][29] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][29] ),
    .S(net5805),
    .X(_05854_));
 sg13g2_nor2b_1 _13914_ (.A(net5805),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][29] ),
    .Y(_05855_));
 sg13g2_a21oi_1 _13915_ (.A1(net5805),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][29] ),
    .Y(_05856_),
    .B1(_05855_));
 sg13g2_o21ai_1 _13916_ (.B1(net5719),
    .Y(_05857_),
    .A1(net5755),
    .A2(_05856_));
 sg13g2_a21oi_1 _13917_ (.A1(net5755),
    .A2(_05854_),
    .Y(_05858_),
    .B1(_05857_));
 sg13g2_nor2_1 _13918_ (.A(net5698),
    .B(_05858_),
    .Y(_05859_));
 sg13g2_o21ai_1 _13919_ (.B1(_05859_),
    .Y(_05860_),
    .A1(net5719),
    .A2(_05853_));
 sg13g2_o21ai_1 _13920_ (.B1(_05860_),
    .Y(_00053_),
    .A1(_05846_),
    .A2(_05852_));
 sg13g2_mux4_1 _13921_ (.S0(net5780),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][30] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][30] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][30] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][30] ),
    .S1(net5738),
    .X(_05861_));
 sg13g2_nor2_1 _13922_ (.A(net5708),
    .B(_05861_),
    .Y(_05862_));
 sg13g2_nor2b_1 _13923_ (.A(net5780),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][30] ),
    .Y(_05863_));
 sg13g2_a21oi_1 _13924_ (.A1(net5780),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][30] ),
    .Y(_05864_),
    .B1(_05863_));
 sg13g2_o21ai_1 _13925_ (.B1(net5740),
    .Y(_05865_),
    .A1(net5781),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][30] ));
 sg13g2_a21oi_1 _13926_ (.A1(net5780),
    .A2(_04372_),
    .Y(_05866_),
    .B1(_05865_));
 sg13g2_o21ai_1 _13927_ (.B1(net5708),
    .Y(_05867_),
    .A1(net5740),
    .A2(_05864_));
 sg13g2_o21ai_1 _13928_ (.B1(net5694),
    .Y(_05868_),
    .A1(_05866_),
    .A2(_05867_));
 sg13g2_mux4_1 _13929_ (.S0(net5780),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][30] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][30] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][30] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][30] ),
    .S1(net5738),
    .X(_05869_));
 sg13g2_mux2_1 _13930_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][30] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][30] ),
    .S(net5780),
    .X(_05870_));
 sg13g2_nor2b_1 _13931_ (.A(net5780),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][30] ),
    .Y(_05871_));
 sg13g2_a21oi_1 _13932_ (.A1(net5780),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][30] ),
    .Y(_05872_),
    .B1(_05871_));
 sg13g2_o21ai_1 _13933_ (.B1(net5708),
    .Y(_05873_),
    .A1(net5738),
    .A2(_05872_));
 sg13g2_a21oi_1 _13934_ (.A1(net5738),
    .A2(_05870_),
    .Y(_05874_),
    .B1(_05873_));
 sg13g2_nor2_1 _13935_ (.A(net5694),
    .B(_05874_),
    .Y(_05875_));
 sg13g2_o21ai_1 _13936_ (.B1(_05875_),
    .Y(_05876_),
    .A1(net5708),
    .A2(_05869_));
 sg13g2_o21ai_1 _13937_ (.B1(_05876_),
    .Y(_00055_),
    .A1(_05862_),
    .A2(_05868_));
 sg13g2_mux4_1 _13938_ (.S0(net5802),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[8][31] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[9][31] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[10][31] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[11][31] ),
    .S1(net5752),
    .X(_05877_));
 sg13g2_nor2_1 _13939_ (.A(net5718),
    .B(_05877_),
    .Y(_05878_));
 sg13g2_nor2b_1 _13940_ (.A(net5809),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[12][31] ),
    .Y(_05879_));
 sg13g2_a21oi_1 _13941_ (.A1(net5809),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[13][31] ),
    .Y(_05880_),
    .B1(_05879_));
 sg13g2_o21ai_1 _13942_ (.B1(net5758),
    .Y(_05881_),
    .A1(net5802),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[14][31] ));
 sg13g2_a21oi_1 _13943_ (.A1(net5809),
    .A2(_04373_),
    .Y(_05882_),
    .B1(_05881_));
 sg13g2_o21ai_1 _13944_ (.B1(net5721),
    .Y(_05883_),
    .A1(net5758),
    .A2(_05880_));
 sg13g2_o21ai_1 _13945_ (.B1(net5699),
    .Y(_05884_),
    .A1(_05882_),
    .A2(_05883_));
 sg13g2_mux4_1 _13946_ (.S0(net5802),
    .A0(\TRNG.sha256.expand.msg_schdl.RAM[0][31] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[1][31] ),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[2][31] ),
    .A3(\TRNG.sha256.expand.msg_schdl.RAM[3][31] ),
    .S1(net5752),
    .X(_05885_));
 sg13g2_mux2_1 _13947_ (.A0(\TRNG.sha256.expand.msg_schdl.RAM[6][31] ),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[7][31] ),
    .S(net5809),
    .X(_05886_));
 sg13g2_nor2b_1 _13948_ (.A(net5809),
    .B_N(\TRNG.sha256.expand.msg_schdl.RAM[4][31] ),
    .Y(_05887_));
 sg13g2_a21oi_1 _13949_ (.A1(net5809),
    .A2(\TRNG.sha256.expand.msg_schdl.RAM[5][31] ),
    .Y(_05888_),
    .B1(_05887_));
 sg13g2_o21ai_1 _13950_ (.B1(net5721),
    .Y(_05889_),
    .A1(net5758),
    .A2(_05888_));
 sg13g2_a21oi_1 _13951_ (.A1(net5758),
    .A2(_05886_),
    .Y(_05890_),
    .B1(_05889_));
 sg13g2_nor2_1 _13952_ (.A(net5699),
    .B(_05890_),
    .Y(_05891_));
 sg13g2_o21ai_1 _13953_ (.B1(_05891_),
    .Y(_05892_),
    .A1(net5718),
    .A2(_05885_));
 sg13g2_o21ai_1 _13954_ (.B1(_05892_),
    .Y(_00056_),
    .A1(_05878_),
    .A2(_05884_));
 sg13g2_nand2_1 _13955_ (.Y(_05893_),
    .A(\TRNG.uart_tx_inst.ticks_counter[7] ),
    .B(net3269));
 sg13g2_nor2_1 _13956_ (.A(net2400),
    .B(_05893_),
    .Y(_05894_));
 sg13g2_nor4_1 _13957_ (.A(\TRNG.uart_tx_inst.ticks_counter[0] ),
    .B(_04302_),
    .C(\TRNG.uart_tx_inst.ticks_counter[3] ),
    .D(net3354),
    .Y(_05895_));
 sg13g2_nand4_1 _13958_ (.B(\TRNG.uart_tx_inst.ticks_counter[4] ),
    .C(_05894_),
    .A(net3169),
    .Y(_05896_),
    .D(_05895_));
 sg13g2_inv_1 _13959_ (.Y(_05897_),
    .A(_05896_));
 sg13g2_nor2_1 _13960_ (.A(_04302_),
    .B(\TRNG.uart_tx_inst.ticks_counter[2] ),
    .Y(_05898_));
 sg13g2_nand4_1 _13961_ (.B(\TRNG.uart_tx_inst.ticks_counter[4] ),
    .C(_05894_),
    .A(\TRNG.uart_tx_inst.ticks_counter[5] ),
    .Y(_05899_),
    .D(_05898_));
 sg13g2_o21ai_1 _13962_ (.B1(_04831_),
    .Y(_05900_),
    .A1(\TRNG.uart_tx_inst.tx_bit_counter[0] ),
    .A2(_05896_));
 sg13g2_a21oi_1 _13963_ (.A1(\TRNG.uart_tx_inst.tx_bit_counter[0] ),
    .A2(_05896_),
    .Y(_05901_),
    .B1(_05900_));
 sg13g2_nand2_1 _13964_ (.Y(_05902_),
    .A(\TRNG.uart_tx_inst.currentState[0] ),
    .B(_04832_));
 sg13g2_nor3_2 _13965_ (.A(net2679),
    .B(\TRNG.uart_tx_inst.currentState[1] ),
    .C(_05902_),
    .Y(_05903_));
 sg13g2_nor2b_2 _13966_ (.A(net2670),
    .B_N(_05903_),
    .Y(_05904_));
 sg13g2_a21oi_1 _13967_ (.A1(net1564),
    .A2(_04830_),
    .Y(_05905_),
    .B1(_05904_));
 sg13g2_nor2b_1 _13968_ (.A(_05901_),
    .B_N(net1565),
    .Y(_00102_));
 sg13g2_nand2_1 _13969_ (.Y(_05906_),
    .A(_04831_),
    .B(_05897_));
 sg13g2_nor4_2 _13970_ (.A(\TRNG.uart_tx_inst.ticks_counter[0] ),
    .B(\TRNG.uart_tx_inst.ticks_counter[3] ),
    .C(_04830_),
    .Y(_05907_),
    .D(_05899_));
 sg13g2_a21oi_1 _13971_ (.A1(net2322),
    .A2(net4749),
    .Y(_05908_),
    .B1(_05904_));
 sg13g2_nand2_1 _13972_ (.Y(_05909_),
    .A(\TRNG.uart_tx_inst.tx_bit_counter[0] ),
    .B(\TRNG.uart_tx_inst.tx_bit_counter[1] ));
 sg13g2_xor2_1 _13973_ (.B(\TRNG.uart_tx_inst.tx_bit_counter[1] ),
    .A(\TRNG.uart_tx_inst.tx_bit_counter[0] ),
    .X(_05910_));
 sg13g2_o21ai_1 _13974_ (.B1(net2323),
    .Y(_05911_),
    .A1(net4749),
    .A2(_05910_));
 sg13g2_inv_1 _13975_ (.Y(_00103_),
    .A(net2324));
 sg13g2_o21ai_1 _13976_ (.B1(net2192),
    .Y(_05912_),
    .A1(net4749),
    .A2(_05909_));
 sg13g2_inv_1 _13977_ (.Y(_05913_),
    .A(net2193));
 sg13g2_nor3_1 _13978_ (.A(net2192),
    .B(net4749),
    .C(_05909_),
    .Y(_05914_));
 sg13g2_nor3_1 _13979_ (.A(_05904_),
    .B(_05913_),
    .C(_05914_),
    .Y(_00104_));
 sg13g2_xor2_1 _13980_ (.B(_05914_),
    .A(net1210),
    .X(_05915_));
 sg13g2_nor2_1 _13981_ (.A(_05904_),
    .B(_05915_),
    .Y(_00105_));
 sg13g2_and2_1 _13982_ (.A(\TRNG.uart_start ),
    .B(_05903_),
    .X(_05916_));
 sg13g2_nand2_1 _13983_ (.Y(_05917_),
    .A(net2999),
    .B(net2680));
 sg13g2_nor2b_1 _13984_ (.A(net5515),
    .B_N(\TRNG.chunk_reg[0] ),
    .Y(_05918_));
 sg13g2_a21oi_1 _13985_ (.A1(net5517),
    .A2(\TRNG.raw_byte[0] ),
    .Y(_05919_),
    .B1(_05918_));
 sg13g2_nand2_1 _13986_ (.Y(_05920_),
    .A(net2482),
    .B(_05907_));
 sg13g2_a21oi_1 _13987_ (.A1(\TRNG.uart_tx_inst.tx_reg[0] ),
    .A2(net4750),
    .Y(_05921_),
    .B1(net4979));
 sg13g2_a22oi_1 _13988_ (.Y(_00106_),
    .B1(net2483),
    .B2(_05921_),
    .A2(_05919_),
    .A1(net4979));
 sg13g2_nor2b_1 _13989_ (.A(net5516),
    .B_N(\TRNG.chunk_reg[1] ),
    .Y(_05922_));
 sg13g2_a21oi_1 _13990_ (.A1(net5516),
    .A2(\TRNG.raw_byte[1] ),
    .Y(_05923_),
    .B1(_05922_));
 sg13g2_nand2_1 _13991_ (.Y(_05924_),
    .A(net2358),
    .B(_05907_));
 sg13g2_a21oi_1 _13992_ (.A1(\TRNG.uart_tx_inst.tx_reg[1] ),
    .A2(net4750),
    .Y(_05925_),
    .B1(net4979));
 sg13g2_a22oi_1 _13993_ (.Y(_00107_),
    .B1(net2359),
    .B2(_05925_),
    .A2(_05923_),
    .A1(net4979));
 sg13g2_nor2b_1 _13994_ (.A(net5515),
    .B_N(\TRNG.chunk_reg[2] ),
    .Y(_05926_));
 sg13g2_a21oi_1 _13995_ (.A1(net5516),
    .A2(\TRNG.raw_byte[2] ),
    .Y(_05927_),
    .B1(_05926_));
 sg13g2_nand2_1 _13996_ (.Y(_05928_),
    .A(net2334),
    .B(_05907_));
 sg13g2_a21oi_1 _13997_ (.A1(\TRNG.uart_tx_inst.tx_reg[2] ),
    .A2(net4750),
    .Y(_05929_),
    .B1(net4979));
 sg13g2_a22oi_1 _13998_ (.Y(_00108_),
    .B1(net2335),
    .B2(_05929_),
    .A2(_05927_),
    .A1(net4978));
 sg13g2_nor2b_1 _13999_ (.A(net5515),
    .B_N(\TRNG.chunk_reg[3] ),
    .Y(_05930_));
 sg13g2_a21oi_1 _14000_ (.A1(net5515),
    .A2(\TRNG.raw_byte[3] ),
    .Y(_05931_),
    .B1(_05930_));
 sg13g2_nand2_1 _14001_ (.Y(_05932_),
    .A(net2325),
    .B(_05907_));
 sg13g2_a21oi_1 _14002_ (.A1(\TRNG.uart_tx_inst.tx_reg[3] ),
    .A2(net4750),
    .Y(_05933_),
    .B1(net4979));
 sg13g2_a22oi_1 _14003_ (.Y(_00109_),
    .B1(net2326),
    .B2(_05933_),
    .A2(_05931_),
    .A1(net4978));
 sg13g2_nor2b_1 _14004_ (.A(net5515),
    .B_N(\TRNG.chunk_reg[4] ),
    .Y(_05934_));
 sg13g2_a21oi_1 _14005_ (.A1(net5515),
    .A2(net2520),
    .Y(_05935_),
    .B1(_05934_));
 sg13g2_nand2_1 _14006_ (.Y(_05936_),
    .A(net2499),
    .B(_05907_));
 sg13g2_a21oi_1 _14007_ (.A1(net2325),
    .A2(net4749),
    .Y(_05937_),
    .B1(net4978));
 sg13g2_a22oi_1 _14008_ (.Y(_00110_),
    .B1(_05936_),
    .B2(_05937_),
    .A2(net2521),
    .A1(net4978));
 sg13g2_nor2b_1 _14009_ (.A(net5516),
    .B_N(\TRNG.chunk_reg[5] ),
    .Y(_05938_));
 sg13g2_a21oi_1 _14010_ (.A1(net5516),
    .A2(\TRNG.raw_byte[5] ),
    .Y(_05939_),
    .B1(_05938_));
 sg13g2_nand2_1 _14011_ (.Y(_05940_),
    .A(net2259),
    .B(_05907_));
 sg13g2_a21oi_1 _14012_ (.A1(net2499),
    .A2(net4749),
    .Y(_05941_),
    .B1(net4978));
 sg13g2_a22oi_1 _14013_ (.Y(_00111_),
    .B1(_05940_),
    .B2(_05941_),
    .A2(_05939_),
    .A1(net4978));
 sg13g2_nor2b_1 _14014_ (.A(net5515),
    .B_N(\TRNG.chunk_reg[6] ),
    .Y(_05942_));
 sg13g2_a21oi_1 _14015_ (.A1(net5515),
    .A2(\TRNG.raw_byte[6] ),
    .Y(_05943_),
    .B1(_05942_));
 sg13g2_nand2_1 _14016_ (.Y(_05944_),
    .A(net2214),
    .B(_05907_));
 sg13g2_a21oi_1 _14017_ (.A1(net2259),
    .A2(net4749),
    .Y(_05945_),
    .B1(net4978));
 sg13g2_a22oi_1 _14018_ (.Y(_00112_),
    .B1(_05944_),
    .B2(_05945_),
    .A2(_05943_),
    .A1(net4978));
 sg13g2_nand3_1 _14019_ (.B(net4749),
    .C(_05917_),
    .A(net2214),
    .Y(_05946_));
 sg13g2_nand2b_1 _14020_ (.Y(_05947_),
    .B(net5516),
    .A_N(\TRNG.raw_byte[7] ));
 sg13g2_o21ai_1 _14021_ (.B1(_05947_),
    .Y(_05948_),
    .A1(net5516),
    .A2(\TRNG.chunk_reg[7] ));
 sg13g2_o21ai_1 _14022_ (.B1(net2215),
    .Y(_00113_),
    .A1(_05917_),
    .A2(_05948_));
 sg13g2_nor2_2 _14023_ (.A(net5607),
    .B(net5614),
    .Y(_05949_));
 sg13g2_or2_2 _14024_ (.X(_05950_),
    .B(net5614),
    .A(net5607));
 sg13g2_nor2_2 _14025_ (.A(net5502),
    .B(_04239_),
    .Y(_05951_));
 sg13g2_nand2_2 _14026_ (.Y(_05952_),
    .A(net5600),
    .B(net5615));
 sg13g2_nor2_2 _14027_ (.A(net5500),
    .B(_05949_),
    .Y(_05953_));
 sg13g2_nand2_1 _14028_ (.Y(_05954_),
    .A(net5607),
    .B(net5614));
 sg13g2_nor2b_2 _14029_ (.A(net5610),
    .B_N(net5607),
    .Y(_05955_));
 sg13g2_nor2_2 _14030_ (.A(net5498),
    .B(net5613),
    .Y(_05956_));
 sg13g2_nand2_2 _14031_ (.Y(_05957_),
    .A(net5611),
    .B(_04239_));
 sg13g2_nand2_2 _14032_ (.Y(_05958_),
    .A(net5605),
    .B(_05957_));
 sg13g2_nor2_2 _14033_ (.A(net5612),
    .B(net5613),
    .Y(_05959_));
 sg13g2_nand2_2 _14034_ (.Y(_05960_),
    .A(net5498),
    .B(net5497));
 sg13g2_nand2_2 _14035_ (.Y(_05961_),
    .A(net5607),
    .B(net5497));
 sg13g2_nor2_2 _14036_ (.A(net5608),
    .B(net5498),
    .Y(_05962_));
 sg13g2_nand2b_2 _14037_ (.Y(_05963_),
    .B(net5610),
    .A_N(net5607));
 sg13g2_nand2_2 _14038_ (.Y(_05964_),
    .A(net5497),
    .B(_05963_));
 sg13g2_nor2_2 _14039_ (.A(_05955_),
    .B(_05962_),
    .Y(_05965_));
 sg13g2_nand2b_2 _14040_ (.Y(_05966_),
    .B(_05963_),
    .A_N(_05955_));
 sg13g2_a21oi_2 _14041_ (.B1(net5592),
    .Y(_05967_),
    .A2(_05965_),
    .A1(net5497));
 sg13g2_nor2_1 _14042_ (.A(net5580),
    .B(_05967_),
    .Y(_05968_));
 sg13g2_nor2_2 _14043_ (.A(net5503),
    .B(net5500),
    .Y(_05969_));
 sg13g2_nand2_2 _14044_ (.Y(_05970_),
    .A(net5584),
    .B(net5602));
 sg13g2_nor2_2 _14045_ (.A(net5503),
    .B(net5588),
    .Y(_05971_));
 sg13g2_nand2_2 _14046_ (.Y(_05972_),
    .A(net5584),
    .B(net5500));
 sg13g2_a221oi_1 _14047_ (.B2(_05960_),
    .C1(_05968_),
    .B1(_05971_),
    .A1(_05949_),
    .Y(_05973_),
    .A2(_05969_));
 sg13g2_a21oi_1 _14048_ (.A1(_05953_),
    .A2(_05958_),
    .Y(_05974_),
    .B1(_05973_));
 sg13g2_and2_2 _14049_ (.A(net5606),
    .B(_00131_),
    .X(_05975_));
 sg13g2_nand2_2 _14050_ (.Y(_05976_),
    .A(net5608),
    .B(_00131_));
 sg13g2_nor2_2 _14051_ (.A(net5604),
    .B(net5612),
    .Y(_05977_));
 sg13g2_or2_2 _14052_ (.X(_05978_),
    .B(net5612),
    .A(net5604));
 sg13g2_nor2_2 _14053_ (.A(net5609),
    .B(net5497),
    .Y(_05979_));
 sg13g2_nor2_2 _14054_ (.A(net5606),
    .B(_05956_),
    .Y(_05980_));
 sg13g2_o21ai_1 _14055_ (.B1(net5588),
    .Y(_05981_),
    .A1(_05975_),
    .A2(_05980_));
 sg13g2_and2_1 _14056_ (.A(net5503),
    .B(_05981_),
    .X(_05982_));
 sg13g2_nor2_2 _14057_ (.A(net5498),
    .B(net5497),
    .Y(_05983_));
 sg13g2_nand2_2 _14058_ (.Y(_05984_),
    .A(net5610),
    .B(net5614));
 sg13g2_nor2_1 _14059_ (.A(_05959_),
    .B(_05983_),
    .Y(_05985_));
 sg13g2_nand2_2 _14060_ (.Y(_05986_),
    .A(_05960_),
    .B(_05984_));
 sg13g2_nand2b_2 _14061_ (.Y(_05987_),
    .B(net5098),
    .A_N(net5606));
 sg13g2_nor2_2 _14062_ (.A(net5610),
    .B(net5497),
    .Y(_05988_));
 sg13g2_nand2_2 _14063_ (.Y(_05989_),
    .A(_04238_),
    .B(net5613));
 sg13g2_or2_1 _14064_ (.X(_05990_),
    .B(net5098),
    .A(net5606));
 sg13g2_nand2_1 _14065_ (.Y(_05991_),
    .A(_05961_),
    .B(_05987_));
 sg13g2_o21ai_1 _14066_ (.B1(_05982_),
    .Y(_05992_),
    .A1(net5588),
    .A2(_05991_));
 sg13g2_nor2_1 _14067_ (.A(net5589),
    .B(net5613),
    .Y(_05993_));
 sg13g2_nor2_2 _14068_ (.A(net5593),
    .B(net5498),
    .Y(_05994_));
 sg13g2_nor2_2 _14069_ (.A(net5593),
    .B(_05988_),
    .Y(_05995_));
 sg13g2_nand2_1 _14070_ (.Y(_05996_),
    .A(net5590),
    .B(_05963_));
 sg13g2_a22oi_1 _14071_ (.Y(_05997_),
    .B1(_05995_),
    .B2(_05950_),
    .A2(net5098),
    .A1(_05953_));
 sg13g2_a21oi_1 _14072_ (.A1(net5580),
    .A2(_05997_),
    .Y(_05998_),
    .B1(net5505));
 sg13g2_nand2_1 _14073_ (.Y(_05999_),
    .A(_05992_),
    .B(_05998_));
 sg13g2_o21ai_1 _14074_ (.B1(_05999_),
    .Y(_00000_),
    .A1(net5576),
    .A2(_05974_));
 sg13g2_and2_2 _14075_ (.A(net5608),
    .B(net5611),
    .X(_06000_));
 sg13g2_nand2_2 _14076_ (.Y(_06001_),
    .A(net5608),
    .B(net5611));
 sg13g2_nand2_2 _14077_ (.Y(_06002_),
    .A(net5608),
    .B(_05989_));
 sg13g2_nor2_2 _14078_ (.A(_05956_),
    .B(_06002_),
    .Y(_06003_));
 sg13g2_nand2_1 _14079_ (.Y(_06004_),
    .A(net5604),
    .B(_05986_));
 sg13g2_nand2_2 _14080_ (.Y(_06005_),
    .A(net5607),
    .B(_05984_));
 sg13g2_nand2_2 _14081_ (.Y(_06006_),
    .A(net5604),
    .B(net5098));
 sg13g2_inv_1 _14082_ (.Y(_06007_),
    .A(_06006_));
 sg13g2_nor3_2 _14083_ (.A(net5591),
    .B(_05949_),
    .C(_06003_),
    .Y(_06008_));
 sg13g2_inv_1 _14084_ (.Y(_06009_),
    .A(_06008_));
 sg13g2_nand2_1 _14085_ (.Y(_06010_),
    .A(_05978_),
    .B(_06008_));
 sg13g2_o21ai_1 _14086_ (.B1(_04236_),
    .Y(_06011_),
    .A1(net5606),
    .A2(_05952_));
 sg13g2_a21oi_1 _14087_ (.A1(_05978_),
    .A2(_06008_),
    .Y(_06012_),
    .B1(_06011_));
 sg13g2_nand2_1 _14088_ (.Y(_06013_),
    .A(net5583),
    .B(_05996_));
 sg13g2_nor2_2 _14089_ (.A(net5201),
    .B(_05979_),
    .Y(_06014_));
 sg13g2_o21ai_1 _14090_ (.B1(net5576),
    .Y(_06015_),
    .A1(_06013_),
    .A2(_06014_));
 sg13g2_nor2_2 _14091_ (.A(net5500),
    .B(net5606),
    .Y(_06016_));
 sg13g2_nand3b_1 _14092_ (.B(_05958_),
    .C(_05987_),
    .Y(_06017_),
    .A_N(_06016_));
 sg13g2_nand2_1 _14093_ (.Y(_06018_),
    .A(net5595),
    .B(net5099));
 sg13g2_nand2_1 _14094_ (.Y(_06019_),
    .A(net5098),
    .B(_06016_));
 sg13g2_nor2_1 _14095_ (.A(net5578),
    .B(net5504),
    .Y(_06020_));
 sg13g2_nand2_2 _14096_ (.Y(_06021_),
    .A(net5507),
    .B(net5584));
 sg13g2_nand2_1 _14097_ (.Y(_06022_),
    .A(net5584),
    .B(_06019_));
 sg13g2_nand3_1 _14098_ (.B(_06019_),
    .C(_06020_),
    .A(_06017_),
    .Y(_06023_));
 sg13g2_and2_1 _14099_ (.A(_05966_),
    .B(_05993_),
    .X(_06024_));
 sg13g2_nand2_2 _14100_ (.Y(_06025_),
    .A(net5590),
    .B(_05978_));
 sg13g2_nor2_1 _14101_ (.A(_06003_),
    .B(_06025_),
    .Y(_06026_));
 sg13g2_nor2_2 _14102_ (.A(net5578),
    .B(net5585),
    .Y(_06027_));
 sg13g2_nand2_1 _14103_ (.Y(_06028_),
    .A(net5506),
    .B(net5503));
 sg13g2_o21ai_1 _14104_ (.B1(_06027_),
    .Y(_06029_),
    .A1(_06024_),
    .A2(_06026_));
 sg13g2_o21ai_1 _14105_ (.B1(_06029_),
    .Y(_06030_),
    .A1(_06012_),
    .A2(_06015_));
 sg13g2_nand2b_2 _14106_ (.Y(_00011_),
    .B(_06023_),
    .A_N(_06030_));
 sg13g2_a21oi_1 _14107_ (.A1(_05963_),
    .A2(_05976_),
    .Y(_06031_),
    .B1(net5594));
 sg13g2_a21oi_1 _14108_ (.A1(net5501),
    .A2(_05979_),
    .Y(_06032_),
    .B1(_06031_));
 sg13g2_nand3_1 _14109_ (.B(_05952_),
    .C(_06032_),
    .A(net5585),
    .Y(_06033_));
 sg13g2_nand2_1 _14110_ (.Y(_06034_),
    .A(net5600),
    .B(_04239_));
 sg13g2_nand2_1 _14111_ (.Y(_06035_),
    .A(net5592),
    .B(_05956_));
 sg13g2_or2_1 _14112_ (.X(_06036_),
    .B(_06025_),
    .A(_05979_));
 sg13g2_nor2_1 _14113_ (.A(net5582),
    .B(_05994_),
    .Y(_06037_));
 sg13g2_a21oi_1 _14114_ (.A1(_06036_),
    .A2(_06037_),
    .Y(_06038_),
    .B1(net5578));
 sg13g2_nor2_1 _14115_ (.A(net5505),
    .B(net5580),
    .Y(_06039_));
 sg13g2_nand2_2 _14116_ (.Y(_06040_),
    .A(net5577),
    .B(net5504));
 sg13g2_nand2b_2 _14117_ (.Y(_06041_),
    .B(_00131_),
    .A_N(net5604));
 sg13g2_a21oi_1 _14118_ (.A1(_06002_),
    .A2(_06041_),
    .Y(_06042_),
    .B1(net5599));
 sg13g2_nor2_1 _14119_ (.A(net5501),
    .B(net5603),
    .Y(_06043_));
 sg13g2_nor2_1 _14120_ (.A(net5603),
    .B(_06018_),
    .Y(_06044_));
 sg13g2_o21ai_1 _14121_ (.B1(net5199),
    .Y(_06045_),
    .A1(_06042_),
    .A2(_06044_));
 sg13g2_nor2_1 _14122_ (.A(net5597),
    .B(net5201),
    .Y(_06046_));
 sg13g2_nor3_2 _14123_ (.A(net5595),
    .B(_05949_),
    .C(_05962_),
    .Y(_06047_));
 sg13g2_nand2_1 _14124_ (.Y(_06048_),
    .A(net5604),
    .B(_05956_));
 sg13g2_nor2_1 _14125_ (.A(net5506),
    .B(net5503),
    .Y(_06049_));
 sg13g2_nand2_2 _14126_ (.Y(_06050_),
    .A(net5579),
    .B(net5586));
 sg13g2_nand2_1 _14127_ (.Y(_06051_),
    .A(net5498),
    .B(net5603));
 sg13g2_a21oi_1 _14128_ (.A1(net5610),
    .A2(_00131_),
    .Y(_06052_),
    .B1(net5502));
 sg13g2_a221oi_1 _14129_ (.B2(_06052_),
    .C1(_06050_),
    .B1(_06051_),
    .A1(_05957_),
    .Y(_06053_),
    .A2(_06047_));
 sg13g2_a21oi_1 _14130_ (.A1(_06033_),
    .A2(_06038_),
    .Y(_06054_),
    .B1(_06053_));
 sg13g2_nand2_2 _14131_ (.Y(_00022_),
    .A(_06045_),
    .B(_06054_));
 sg13g2_nand2_2 _14132_ (.Y(_06055_),
    .A(net5606),
    .B(_05959_));
 sg13g2_and2_1 _14133_ (.A(_06041_),
    .B(_06055_),
    .X(_06056_));
 sg13g2_nand2_1 _14134_ (.Y(_06057_),
    .A(net5613),
    .B(_05955_));
 sg13g2_nand2_1 _14135_ (.Y(_06058_),
    .A(_06041_),
    .B(_06057_));
 sg13g2_a21oi_1 _14136_ (.A1(net5599),
    .A2(_06058_),
    .Y(_06059_),
    .B1(net5585));
 sg13g2_o21ai_1 _14137_ (.B1(_06059_),
    .Y(_06060_),
    .A1(net5598),
    .A2(_06056_));
 sg13g2_nor3_1 _14138_ (.A(net5598),
    .B(_05949_),
    .C(_05977_),
    .Y(_06061_));
 sg13g2_o21ai_1 _14139_ (.B1(_06060_),
    .Y(_06062_),
    .A1(_06022_),
    .A2(_06061_));
 sg13g2_nand2_1 _14140_ (.Y(_06063_),
    .A(net5498),
    .B(net5359));
 sg13g2_nand2_2 _14141_ (.Y(_06064_),
    .A(_05950_),
    .B(net5359));
 sg13g2_nor2_2 _14142_ (.A(net5610),
    .B(_06064_),
    .Y(_06065_));
 sg13g2_nand2_1 _14143_ (.Y(_06066_),
    .A(net5601),
    .B(_06065_));
 sg13g2_nand2_2 _14144_ (.Y(_06067_),
    .A(net5604),
    .B(_00132_));
 sg13g2_nor2b_1 _14145_ (.A(_05980_),
    .B_N(_06067_),
    .Y(_06068_));
 sg13g2_a22oi_1 _14146_ (.Y(_06069_),
    .B1(_06068_),
    .B2(net5586),
    .A2(_06066_),
    .A1(_05970_));
 sg13g2_nor2_1 _14147_ (.A(net5599),
    .B(_05986_),
    .Y(_06070_));
 sg13g2_nand2_1 _14148_ (.Y(_06071_),
    .A(net5501),
    .B(net5099));
 sg13g2_o21ai_1 _14149_ (.B1(net5579),
    .Y(_06072_),
    .A1(_06069_),
    .A2(_06070_));
 sg13g2_o21ai_1 _14150_ (.B1(_06072_),
    .Y(_00025_),
    .A1(net5579),
    .A2(_06062_));
 sg13g2_nand3_1 _14151_ (.B(_06014_),
    .C(_06067_),
    .A(net5499),
    .Y(_06073_));
 sg13g2_nand2_1 _14152_ (.Y(_06074_),
    .A(net5199),
    .B(_06073_));
 sg13g2_nand2_2 _14153_ (.Y(_06075_),
    .A(_05957_),
    .B(_06016_));
 sg13g2_o21ai_1 _14154_ (.B1(net5597),
    .Y(_06076_),
    .A1(_05980_),
    .A2(_06007_));
 sg13g2_inv_1 _14155_ (.Y(_06077_),
    .A(_06076_));
 sg13g2_nor2_1 _14156_ (.A(net5612),
    .B(_05950_),
    .Y(_06078_));
 sg13g2_o21ai_1 _14157_ (.B1(net5589),
    .Y(_06079_),
    .A1(_05975_),
    .A2(_06078_));
 sg13g2_nand2_1 _14158_ (.Y(_06080_),
    .A(net5501),
    .B(_06000_));
 sg13g2_nand3_1 _14159_ (.B(_06079_),
    .C(_06080_),
    .A(net5582),
    .Y(_06081_));
 sg13g2_nand2b_2 _14160_ (.Y(_06082_),
    .B(_00132_),
    .A_N(net5604));
 sg13g2_mux2_1 _14161_ (.A0(_06041_),
    .A1(_06082_),
    .S(net5499),
    .X(_06083_));
 sg13g2_a21oi_1 _14162_ (.A1(net5605),
    .A2(_05957_),
    .Y(_06084_),
    .B1(net5586));
 sg13g2_a21oi_1 _14163_ (.A1(_06083_),
    .A2(_06084_),
    .Y(_06085_),
    .B1(net5579));
 sg13g2_o21ai_1 _14164_ (.B1(_06035_),
    .Y(_06086_),
    .A1(net5098),
    .A2(_06016_));
 sg13g2_a22oi_1 _14165_ (.Y(_06087_),
    .B1(_06086_),
    .B2(_06049_),
    .A2(_06085_),
    .A1(_06081_));
 sg13g2_o21ai_1 _14166_ (.B1(_06087_),
    .Y(_00026_),
    .A1(_06074_),
    .A2(_06077_));
 sg13g2_a21oi_1 _14167_ (.A1(_06010_),
    .A2(_06036_),
    .Y(_06088_),
    .B1(_06028_));
 sg13g2_o21ai_1 _14168_ (.B1(net5359),
    .Y(_06089_),
    .A1(net5607),
    .A2(_05988_));
 sg13g2_nand2_1 _14169_ (.Y(_06090_),
    .A(net5593),
    .B(_06089_));
 sg13g2_a21oi_1 _14170_ (.A1(_06071_),
    .A2(_06090_),
    .Y(_06091_),
    .B1(_06040_));
 sg13g2_nand3_1 _14171_ (.B(_05978_),
    .C(_05986_),
    .A(net5499),
    .Y(_06092_));
 sg13g2_a21oi_1 _14172_ (.A1(_05996_),
    .A2(_06092_),
    .Y(_06093_),
    .B1(net5358));
 sg13g2_nor2_2 _14173_ (.A(net5608),
    .B(_05989_),
    .Y(_06094_));
 sg13g2_nand2_1 _14174_ (.Y(_06095_),
    .A(_04238_),
    .B(_05979_));
 sg13g2_nor3_1 _14175_ (.A(net5500),
    .B(_06003_),
    .C(_06094_),
    .Y(_06096_));
 sg13g2_nor2_2 _14176_ (.A(net5593),
    .B(_05955_),
    .Y(_06097_));
 sg13g2_nor3_1 _14177_ (.A(_06021_),
    .B(_06096_),
    .C(_06097_),
    .Y(_06098_));
 sg13g2_or4_1 _14178_ (.A(_06088_),
    .B(_06091_),
    .C(_06093_),
    .D(_06098_),
    .X(_00027_));
 sg13g2_nand2_1 _14179_ (.Y(_06099_),
    .A(net5499),
    .B(net5615));
 sg13g2_nor2_1 _14180_ (.A(net5588),
    .B(net5359),
    .Y(_06100_));
 sg13g2_o21ai_1 _14181_ (.B1(net5503),
    .Y(_06101_),
    .A1(_05956_),
    .A2(_06025_));
 sg13g2_nor3_1 _14182_ (.A(_06024_),
    .B(_06100_),
    .C(_06101_),
    .Y(_06102_));
 sg13g2_a21o_1 _14183_ (.A2(_05988_),
    .A1(_05971_),
    .B1(_06102_),
    .X(_06103_));
 sg13g2_nor2_1 _14184_ (.A(net5590),
    .B(_05979_),
    .Y(_06104_));
 sg13g2_inv_1 _14185_ (.Y(_06105_),
    .A(_06104_));
 sg13g2_nor2_1 _14186_ (.A(_05959_),
    .B(_06105_),
    .Y(_06106_));
 sg13g2_nor3_1 _14187_ (.A(net5505),
    .B(_06013_),
    .C(_06106_),
    .Y(_06107_));
 sg13g2_nand3_1 _14188_ (.B(_05990_),
    .C(_06005_),
    .A(net5588),
    .Y(_06108_));
 sg13g2_nor2_1 _14189_ (.A(_06024_),
    .B(_06040_),
    .Y(_06109_));
 sg13g2_a221oi_1 _14190_ (.B2(_06109_),
    .C1(_06107_),
    .B1(_06108_),
    .A1(net5505),
    .Y(_00028_),
    .A2(_06103_));
 sg13g2_nand3_1 _14191_ (.B(_05958_),
    .C(_05987_),
    .A(net5596),
    .Y(_06110_));
 sg13g2_nor2_2 _14192_ (.A(net5592),
    .B(_05950_),
    .Y(_06111_));
 sg13g2_nor2_2 _14193_ (.A(net5582),
    .B(_06111_),
    .Y(_06112_));
 sg13g2_nand2_1 _14194_ (.Y(_06113_),
    .A(_06110_),
    .B(_06112_));
 sg13g2_nand2_1 _14195_ (.Y(_06114_),
    .A(net5596),
    .B(_06014_));
 sg13g2_nand3_1 _14196_ (.B(_06092_),
    .C(_06114_),
    .A(net5584),
    .Y(_06115_));
 sg13g2_o21ai_1 _14197_ (.B1(_06115_),
    .Y(_06116_),
    .A1(_06100_),
    .A2(_06113_));
 sg13g2_nor2b_1 _14198_ (.A(_05970_),
    .B_N(net5359),
    .Y(_06117_));
 sg13g2_or2_1 _14199_ (.X(_06118_),
    .B(_00130_),
    .A(net5613));
 sg13g2_nor2_1 _14200_ (.A(net5612),
    .B(_06118_),
    .Y(_06119_));
 sg13g2_a22oi_1 _14201_ (.Y(_06120_),
    .B1(_06117_),
    .B2(_05966_),
    .A2(_06096_),
    .A1(net5504));
 sg13g2_o21ai_1 _14202_ (.B1(_06120_),
    .Y(_06121_),
    .A1(net5596),
    .A2(_06119_));
 sg13g2_nand2_1 _14203_ (.Y(_06122_),
    .A(net5507),
    .B(_06121_));
 sg13g2_o21ai_1 _14204_ (.B1(_06122_),
    .Y(_00029_),
    .A1(_04235_),
    .A2(_06116_));
 sg13g2_nand3_1 _14205_ (.B(net5611),
    .C(_05954_),
    .A(net5594),
    .Y(_06123_));
 sg13g2_a21oi_1 _14206_ (.A1(_06032_),
    .A2(_06123_),
    .Y(_06124_),
    .B1(net5585));
 sg13g2_nand2_1 _14207_ (.Y(_06125_),
    .A(_05976_),
    .B(_06095_));
 sg13g2_a21oi_1 _14208_ (.A1(_05976_),
    .A2(_06095_),
    .Y(_06126_),
    .B1(_05970_));
 sg13g2_nand2_1 _14209_ (.Y(_06127_),
    .A(net5605),
    .B(_05983_));
 sg13g2_a21oi_1 _14210_ (.A1(_06041_),
    .A2(_06127_),
    .Y(_06128_),
    .B1(_05972_));
 sg13g2_nor4_1 _14211_ (.A(net5507),
    .B(_06124_),
    .C(_06126_),
    .D(_06128_),
    .Y(_06129_));
 sg13g2_nor2_2 _14212_ (.A(net5594),
    .B(net5603),
    .Y(_06130_));
 sg13g2_a22oi_1 _14213_ (.Y(_06131_),
    .B1(_06130_),
    .B2(_05957_),
    .A2(_06094_),
    .A1(net5594));
 sg13g2_nor2_1 _14214_ (.A(_06021_),
    .B(_06131_),
    .Y(_06132_));
 sg13g2_nor2_2 _14215_ (.A(net5599),
    .B(_06065_),
    .Y(_06133_));
 sg13g2_o21ai_1 _14216_ (.B1(net5594),
    .Y(_06134_),
    .A1(net5613),
    .A2(_05966_));
 sg13g2_nand2_1 _14217_ (.Y(_06135_),
    .A(_06027_),
    .B(_06134_));
 sg13g2_a21oi_1 _14218_ (.A1(_06001_),
    .A2(_06133_),
    .Y(_06136_),
    .B1(_06135_));
 sg13g2_nor3_2 _14219_ (.A(_06129_),
    .B(_06132_),
    .C(_06136_),
    .Y(_00030_));
 sg13g2_nand2_1 _14220_ (.Y(_06137_),
    .A(net5497),
    .B(net5201));
 sg13g2_a21oi_1 _14221_ (.A1(_05952_),
    .A2(_05996_),
    .Y(_06138_),
    .B1(_05988_));
 sg13g2_o21ai_1 _14222_ (.B1(_06067_),
    .Y(_06139_),
    .A1(net5613),
    .A2(_05978_));
 sg13g2_o21ai_1 _14223_ (.B1(net5199),
    .Y(_06140_),
    .A1(net5590),
    .A2(_06139_));
 sg13g2_o21ai_1 _14224_ (.B1(net5590),
    .Y(_06141_),
    .A1(net5201),
    .A2(_05975_));
 sg13g2_nor2b_1 _14225_ (.A(_05979_),
    .B_N(_06141_),
    .Y(_06142_));
 sg13g2_nor3_1 _14226_ (.A(_05994_),
    .B(_06021_),
    .C(_06142_),
    .Y(_06143_));
 sg13g2_or2_2 _14227_ (.X(_06144_),
    .B(_00132_),
    .A(net5605));
 sg13g2_a21oi_1 _14228_ (.A1(_06048_),
    .A2(_06082_),
    .Y(_06145_),
    .B1(net5499));
 sg13g2_or2_1 _14229_ (.X(_06146_),
    .B(_06145_),
    .A(_05995_));
 sg13g2_o21ai_1 _14230_ (.B1(_05981_),
    .Y(_06147_),
    .A1(_05959_),
    .A2(_06105_));
 sg13g2_a221oi_1 _14231_ (.B2(net5198),
    .C1(_06143_),
    .B1(_06147_),
    .A1(_06027_),
    .Y(_06148_),
    .A2(_06146_));
 sg13g2_o21ai_1 _14232_ (.B1(_06148_),
    .Y(_00031_),
    .A1(_06138_),
    .A2(_06140_));
 sg13g2_nand3_1 _14233_ (.B(_06005_),
    .C(_06144_),
    .A(net5500),
    .Y(_06149_));
 sg13g2_a21oi_1 _14234_ (.A1(_06141_),
    .A2(_06149_),
    .Y(_06150_),
    .B1(net5580));
 sg13g2_a21oi_1 _14235_ (.A1(_05987_),
    .A2(_06067_),
    .Y(_06151_),
    .B1(_05972_));
 sg13g2_nor2_1 _14236_ (.A(_05970_),
    .B(_06014_),
    .Y(_06152_));
 sg13g2_nor3_1 _14237_ (.A(_06150_),
    .B(_06151_),
    .C(_06152_),
    .Y(_06153_));
 sg13g2_a21oi_2 _14238_ (.B1(net5596),
    .Y(_06154_),
    .A2(_06014_),
    .A1(_06004_));
 sg13g2_a21o_2 _14239_ (.A2(_05955_),
    .A1(net5592),
    .B1(net5504),
    .X(_06155_));
 sg13g2_a221oi_1 _14240_ (.B2(_05961_),
    .C1(net5580),
    .B1(_05994_),
    .A1(_05953_),
    .Y(_06156_),
    .A2(net5098));
 sg13g2_nor2_1 _14241_ (.A(net5505),
    .B(_06156_),
    .Y(_06157_));
 sg13g2_o21ai_1 _14242_ (.B1(_06157_),
    .Y(_06158_),
    .A1(_06154_),
    .A2(_06155_));
 sg13g2_o21ai_1 _14243_ (.B1(_06158_),
    .Y(_00001_),
    .A1(net5576),
    .A2(_06153_));
 sg13g2_nor2_1 _14244_ (.A(_04374_),
    .B(_06034_),
    .Y(_06159_));
 sg13g2_a21oi_2 _14245_ (.B1(_06159_),
    .Y(_06160_),
    .A2(_05951_),
    .A1(_00130_));
 sg13g2_a21oi_1 _14246_ (.A1(_05995_),
    .A2(_06118_),
    .Y(_06161_),
    .B1(net5586));
 sg13g2_o21ai_1 _14247_ (.B1(net5585),
    .Y(_06162_),
    .A1(net5099),
    .A2(_06025_));
 sg13g2_a21oi_1 _14248_ (.A1(_06160_),
    .A2(_06161_),
    .Y(_06163_),
    .B1(net5579));
 sg13g2_o21ai_1 _14249_ (.B1(_06163_),
    .Y(_06164_),
    .A1(_06042_),
    .A2(_06162_));
 sg13g2_nor2_1 _14250_ (.A(net5499),
    .B(_06056_),
    .Y(_06165_));
 sg13g2_o21ai_1 _14251_ (.B1(net5200),
    .Y(_06166_),
    .A1(_06133_),
    .A2(_06165_));
 sg13g2_nand3_1 _14252_ (.B(_05958_),
    .C(_06137_),
    .A(net5599),
    .Y(_06167_));
 sg13g2_nand3b_1 _14253_ (.B(_06167_),
    .C(net5198),
    .Y(_06168_),
    .A_N(_06111_));
 sg13g2_nand3_1 _14254_ (.B(_06166_),
    .C(_06168_),
    .A(_06164_),
    .Y(_00002_));
 sg13g2_a21oi_1 _14255_ (.A1(_05987_),
    .A2(_06055_),
    .Y(_06169_),
    .B1(net5589));
 sg13g2_nor4_1 _14256_ (.A(net5580),
    .B(_05949_),
    .C(_05956_),
    .D(_06169_),
    .Y(_06170_));
 sg13g2_and2_1 _14257_ (.A(_05969_),
    .B(_05987_),
    .X(_06171_));
 sg13g2_nand2_1 _14258_ (.Y(_06172_),
    .A(_05949_),
    .B(_05994_));
 sg13g2_a221oi_1 _14259_ (.B2(_06171_),
    .C1(_06170_),
    .B1(_06002_),
    .A1(_05949_),
    .Y(_06173_),
    .A2(_05994_));
 sg13g2_nand2_2 _14260_ (.Y(_06174_),
    .A(net5614),
    .B(net5201));
 sg13g2_nand3_1 _14261_ (.B(_06048_),
    .C(_06174_),
    .A(net5596),
    .Y(_06175_));
 sg13g2_o21ai_1 _14262_ (.B1(net5199),
    .Y(_06176_),
    .A1(net5597),
    .A2(_06119_));
 sg13g2_inv_1 _14263_ (.Y(_06177_),
    .A(_06176_));
 sg13g2_nor2_1 _14264_ (.A(_06046_),
    .B(net5358),
    .Y(_06178_));
 sg13g2_a22oi_1 _14265_ (.Y(_06179_),
    .B1(_06178_),
    .B2(_06076_),
    .A2(_06177_),
    .A1(_06175_));
 sg13g2_o21ai_1 _14266_ (.B1(_06179_),
    .Y(_00003_),
    .A1(net5576),
    .A2(_06173_));
 sg13g2_a21oi_2 _14267_ (.B1(net5588),
    .Y(_06180_),
    .A2(_06006_),
    .A1(_05990_));
 sg13g2_inv_1 _14268_ (.Y(_06181_),
    .A(_06180_));
 sg13g2_nand3_1 _14269_ (.B(_06002_),
    .C(_06082_),
    .A(net5590),
    .Y(_06182_));
 sg13g2_nand2_1 _14270_ (.Y(_06183_),
    .A(net5503),
    .B(_06182_));
 sg13g2_a22oi_1 _14271_ (.Y(_06184_),
    .B1(_05990_),
    .B2(_05969_),
    .A2(_05971_),
    .A1(_05964_));
 sg13g2_o21ai_1 _14272_ (.B1(_06184_),
    .Y(_06185_),
    .A1(_06180_),
    .A2(_06183_));
 sg13g2_nand3_1 _14273_ (.B(_05961_),
    .C(_05987_),
    .A(net5588),
    .Y(_06186_));
 sg13g2_nor2_1 _14274_ (.A(_05972_),
    .B(_05975_),
    .Y(_06187_));
 sg13g2_o21ai_1 _14275_ (.B1(net5505),
    .Y(_06188_),
    .A1(net5612),
    .A2(_05970_));
 sg13g2_a221oi_1 _14276_ (.B2(_05990_),
    .C1(_06188_),
    .B1(_06187_),
    .A1(_06112_),
    .Y(_06189_),
    .A2(_06186_));
 sg13g2_a21o_1 _14277_ (.A2(_06185_),
    .A1(net5576),
    .B1(_06189_),
    .X(_00004_));
 sg13g2_nor4_1 _14278_ (.A(net5584),
    .B(_05979_),
    .C(_06003_),
    .D(_06154_),
    .Y(_06190_));
 sg13g2_nand2_1 _14279_ (.Y(_06191_),
    .A(net5499),
    .B(_05977_));
 sg13g2_nand3_1 _14280_ (.B(_06167_),
    .C(_06191_),
    .A(net5585),
    .Y(_06192_));
 sg13g2_nand2_1 _14281_ (.Y(_06193_),
    .A(net5507),
    .B(_06192_));
 sg13g2_a21oi_1 _14282_ (.A1(_05976_),
    .A2(_06137_),
    .Y(_06194_),
    .B1(net5599));
 sg13g2_nand2b_1 _14283_ (.Y(_06195_),
    .B(_06160_),
    .A_N(_06194_));
 sg13g2_a21oi_1 _14284_ (.A1(_06001_),
    .A2(_06061_),
    .Y(_06196_),
    .B1(net5358));
 sg13g2_a22oi_1 _14285_ (.Y(_06197_),
    .B1(_06196_),
    .B2(_06110_),
    .A2(_06195_),
    .A1(net5199));
 sg13g2_o21ai_1 _14286_ (.B1(_06197_),
    .Y(_00005_),
    .A1(_06190_),
    .A2(_06193_));
 sg13g2_nand2_2 _14287_ (.Y(_06198_),
    .A(_06056_),
    .B(_06127_));
 sg13g2_a22oi_1 _14288_ (.Y(_06199_),
    .B1(_06198_),
    .B2(net5589),
    .A2(_06130_),
    .A1(_05956_));
 sg13g2_a21oi_1 _14289_ (.A1(net5592),
    .A2(_06064_),
    .Y(_06200_),
    .B1(_06031_));
 sg13g2_a22oi_1 _14290_ (.Y(_06201_),
    .B1(_06063_),
    .B2(_05971_),
    .A2(_05988_),
    .A1(_05969_));
 sg13g2_o21ai_1 _14291_ (.B1(_06201_),
    .Y(_06202_),
    .A1(net5581),
    .A2(_06200_));
 sg13g2_nand2_1 _14292_ (.Y(_06203_),
    .A(_06079_),
    .B(_06181_));
 sg13g2_a22oi_1 _14293_ (.Y(_06204_),
    .B1(_06203_),
    .B2(net5198),
    .A2(_06202_),
    .A1(net5506));
 sg13g2_o21ai_1 _14294_ (.B1(_06204_),
    .Y(_00006_),
    .A1(_06040_),
    .A2(_06199_));
 sg13g2_nand2_1 _14295_ (.Y(_06205_),
    .A(_06005_),
    .B(_06174_));
 sg13g2_nand3_1 _14296_ (.B(_06005_),
    .C(_06174_),
    .A(net5588),
    .Y(_06206_));
 sg13g2_a21oi_1 _14297_ (.A1(_06009_),
    .A2(_06206_),
    .Y(_06207_),
    .B1(net5580));
 sg13g2_a221oi_1 _14298_ (.B2(_06198_),
    .C1(_06207_),
    .B1(_05971_),
    .A1(_05964_),
    .Y(_06208_),
    .A2(_05969_));
 sg13g2_nand2_1 _14299_ (.Y(_06209_),
    .A(_06059_),
    .B(_06191_));
 sg13g2_a21oi_1 _14300_ (.A1(net5599),
    .A2(_06000_),
    .Y(_06210_),
    .B1(_06094_));
 sg13g2_nand3_1 _14301_ (.B(_06075_),
    .C(_06210_),
    .A(net5585),
    .Y(_06211_));
 sg13g2_nand3_1 _14302_ (.B(_06209_),
    .C(_06211_),
    .A(net3283),
    .Y(_06212_));
 sg13g2_o21ai_1 _14303_ (.B1(_06212_),
    .Y(_00007_),
    .A1(net5576),
    .A2(_06208_));
 sg13g2_nand3_1 _14304_ (.B(net5359),
    .C(_05986_),
    .A(net5598),
    .Y(_06213_));
 sg13g2_o21ai_1 _14305_ (.B1(_06213_),
    .Y(_06214_),
    .A1(_05966_),
    .A2(_06099_));
 sg13g2_a221oi_1 _14306_ (.B2(_05951_),
    .C1(_06040_),
    .B1(_05966_),
    .A1(net5501),
    .Y(_06215_),
    .A2(net5201));
 sg13g2_and3_1 _14307_ (.X(_06216_),
    .A(net5596),
    .B(_06006_),
    .C(_06041_));
 sg13g2_o21ai_1 _14308_ (.B1(_06020_),
    .Y(_06217_),
    .A1(net5590),
    .A2(_05977_));
 sg13g2_nand3_1 _14309_ (.B(_06048_),
    .C(_06144_),
    .A(net5598),
    .Y(_06218_));
 sg13g2_and2_1 _14310_ (.A(_05976_),
    .B(_06082_),
    .X(_06219_));
 sg13g2_o21ai_1 _14311_ (.B1(_06218_),
    .Y(_06220_),
    .A1(net5591),
    .A2(_06219_));
 sg13g2_a221oi_1 _14312_ (.B2(_06027_),
    .C1(_06215_),
    .B1(_06220_),
    .A1(net5198),
    .Y(_06221_),
    .A2(_06214_));
 sg13g2_o21ai_1 _14313_ (.B1(_06221_),
    .Y(_00008_),
    .A1(_06216_),
    .A2(_06217_));
 sg13g2_a21oi_1 _14314_ (.A1(_06002_),
    .A2(_06082_),
    .Y(_06222_),
    .B1(net5596));
 sg13g2_nand2_1 _14315_ (.Y(_06223_),
    .A(net5587),
    .B(_06160_));
 sg13g2_o21ai_1 _14316_ (.B1(_06113_),
    .Y(_06224_),
    .A1(_06222_),
    .A2(_06223_));
 sg13g2_a21oi_1 _14317_ (.A1(_06002_),
    .A2(_06104_),
    .Y(_06225_),
    .B1(_06028_));
 sg13g2_a21oi_1 _14318_ (.A1(_06099_),
    .A2(_06114_),
    .Y(_06226_),
    .B1(_06021_));
 sg13g2_a22oi_1 _14319_ (.Y(_06227_),
    .B1(_06226_),
    .B2(_06002_),
    .A2(_06225_),
    .A1(_06108_));
 sg13g2_o21ai_1 _14320_ (.B1(_06227_),
    .Y(_00009_),
    .A1(net5507),
    .A2(_06224_));
 sg13g2_nor2b_1 _14321_ (.A(_05955_),
    .B_N(_06171_),
    .Y(_06228_));
 sg13g2_a21oi_1 _14322_ (.A1(_05978_),
    .A2(net5098),
    .Y(_06229_),
    .B1(_05972_));
 sg13g2_a22oi_1 _14323_ (.Y(_06230_),
    .B1(_05995_),
    .B2(_05965_),
    .A2(_05978_),
    .A1(_05953_));
 sg13g2_nor2_1 _14324_ (.A(net5583),
    .B(_06230_),
    .Y(_06231_));
 sg13g2_nor3_1 _14325_ (.A(_06228_),
    .B(_06229_),
    .C(_06231_),
    .Y(_06232_));
 sg13g2_nand2_1 _14326_ (.Y(_06233_),
    .A(_00131_),
    .B(_05969_));
 sg13g2_o21ai_1 _14327_ (.B1(_06233_),
    .Y(_06234_),
    .A1(_05972_),
    .A2(_05980_));
 sg13g2_a21oi_1 _14328_ (.A1(net5597),
    .A2(_06119_),
    .Y(_06235_),
    .B1(_06074_));
 sg13g2_a21oi_1 _14329_ (.A1(net5579),
    .A2(_06234_),
    .Y(_06236_),
    .B1(_06235_));
 sg13g2_o21ai_1 _14330_ (.B1(_06236_),
    .Y(_00010_),
    .A1(net5579),
    .A2(_06232_));
 sg13g2_nand2_1 _14331_ (.Y(_06237_),
    .A(_06055_),
    .B(_06144_));
 sg13g2_nor2_1 _14332_ (.A(net5592),
    .B(_06237_),
    .Y(_06238_));
 sg13g2_o21ai_1 _14333_ (.B1(_06075_),
    .Y(_06239_),
    .A1(net5592),
    .A2(_06237_));
 sg13g2_a22oi_1 _14334_ (.Y(_06240_),
    .B1(_06239_),
    .B2(net5581),
    .A2(_06112_),
    .A1(_06075_));
 sg13g2_a21o_1 _14335_ (.A2(_06051_),
    .A1(_05984_),
    .B1(net5594),
    .X(_06241_));
 sg13g2_o21ai_1 _14336_ (.B1(_06241_),
    .Y(_06242_),
    .A1(net5501),
    .A2(_04374_));
 sg13g2_a21oi_1 _14337_ (.A1(_06064_),
    .A2(_06097_),
    .Y(_06243_),
    .B1(_06016_));
 sg13g2_a22oi_1 _14338_ (.Y(_06244_),
    .B1(_06243_),
    .B2(net5198),
    .A2(_06242_),
    .A1(net5200));
 sg13g2_o21ai_1 _14339_ (.B1(_06244_),
    .Y(_00012_),
    .A1(net5577),
    .A2(_06240_));
 sg13g2_o21ai_1 _14340_ (.B1(net5595),
    .Y(_06245_),
    .A1(_06000_),
    .A2(_06065_));
 sg13g2_nand3_1 _14341_ (.B(_06241_),
    .C(_06245_),
    .A(net5577),
    .Y(_06246_));
 sg13g2_nor2_1 _14342_ (.A(net5577),
    .B(_06047_),
    .Y(_06247_));
 sg13g2_a21oi_1 _14343_ (.A1(_06218_),
    .A2(_06247_),
    .Y(_06248_),
    .B1(net5504));
 sg13g2_nand2_1 _14344_ (.Y(_06249_),
    .A(_06246_),
    .B(_06248_));
 sg13g2_nand3_1 _14345_ (.B(net5200),
    .C(_06089_),
    .A(_06018_),
    .Y(_06250_));
 sg13g2_nor2_2 _14346_ (.A(_05965_),
    .B(_06034_),
    .Y(_06251_));
 sg13g2_o21ai_1 _14347_ (.B1(_06027_),
    .Y(_06252_),
    .A1(_06008_),
    .A2(_06251_));
 sg13g2_nand3_1 _14348_ (.B(_06250_),
    .C(_06252_),
    .A(_06249_),
    .Y(_00013_));
 sg13g2_a21oi_1 _14349_ (.A1(_06067_),
    .A2(_06137_),
    .Y(_06253_),
    .B1(net5599));
 sg13g2_nor3_1 _14350_ (.A(net5585),
    .B(_06044_),
    .C(_06253_),
    .Y(_06254_));
 sg13g2_nor2_1 _14351_ (.A(net5503),
    .B(_05975_),
    .Y(_06255_));
 sg13g2_a21oi_1 _14352_ (.A1(_06174_),
    .A2(_06255_),
    .Y(_06256_),
    .B1(_05971_));
 sg13g2_nor3_1 _14353_ (.A(_06024_),
    .B(_06100_),
    .C(_06256_),
    .Y(_06257_));
 sg13g2_nor3_1 _14354_ (.A(net5577),
    .B(_06254_),
    .C(_06257_),
    .Y(_06258_));
 sg13g2_nand2_1 _14355_ (.Y(_06259_),
    .A(_05960_),
    .B(_06130_));
 sg13g2_nand3_1 _14356_ (.B(net5610),
    .C(_05961_),
    .A(net5593),
    .Y(_06260_));
 sg13g2_a21oi_1 _14357_ (.A1(_06259_),
    .A2(_06260_),
    .Y(_06261_),
    .B1(_06040_));
 sg13g2_a221oi_1 _14358_ (.B2(_05950_),
    .C1(_06050_),
    .B1(_05995_),
    .A1(net5498),
    .Y(_06262_),
    .A2(net5359));
 sg13g2_or3_1 _14359_ (.A(_06258_),
    .B(_06261_),
    .C(_06262_),
    .X(_00014_));
 sg13g2_a21o_1 _14360_ (.A2(net5359),
    .A1(net5589),
    .B1(_06180_),
    .X(_06263_));
 sg13g2_a221oi_1 _14361_ (.B2(_06133_),
    .C1(net5581),
    .B1(_06001_),
    .A1(_05953_),
    .Y(_06264_),
    .A2(_05963_));
 sg13g2_a21oi_1 _14362_ (.A1(net5614),
    .A2(net5201),
    .Y(_06265_),
    .B1(net5593));
 sg13g2_a221oi_1 _14363_ (.B2(_06265_),
    .C1(net5504),
    .B1(_06057_),
    .A1(_05984_),
    .Y(_06266_),
    .A2(_06043_));
 sg13g2_nor3_1 _14364_ (.A(net5578),
    .B(_06264_),
    .C(_06266_),
    .Y(_06267_));
 sg13g2_o21ai_1 _14365_ (.B1(net5199),
    .Y(_06268_),
    .A1(net5500),
    .A2(_06139_));
 sg13g2_a21oi_1 _14366_ (.A1(net5198),
    .A2(_06263_),
    .Y(_06269_),
    .B1(_06267_));
 sg13g2_o21ai_1 _14367_ (.B1(_06269_),
    .Y(_00015_),
    .A1(_05967_),
    .A2(_06268_));
 sg13g2_o21ai_1 _14368_ (.B1(net5580),
    .Y(_06270_),
    .A1(_05952_),
    .A2(_05965_));
 sg13g2_nand2_1 _14369_ (.Y(_06271_),
    .A(net5612),
    .B(_05953_));
 sg13g2_a21oi_1 _14370_ (.A1(_05968_),
    .A2(_06271_),
    .Y(_06272_),
    .B1(net5576));
 sg13g2_o21ai_1 _14371_ (.B1(_06272_),
    .Y(_06273_),
    .A1(_06169_),
    .A2(_06270_));
 sg13g2_nor3_1 _14372_ (.A(_05956_),
    .B(_06025_),
    .C(_06064_),
    .Y(_06274_));
 sg13g2_or3_1 _14373_ (.A(_06031_),
    .B(_06111_),
    .C(_06274_),
    .X(_06275_));
 sg13g2_a22oi_1 _14374_ (.Y(_06276_),
    .B1(_06275_),
    .B2(net5200),
    .A2(net5198),
    .A1(_05993_));
 sg13g2_nand2_1 _14375_ (.Y(_00016_),
    .A(_06273_),
    .B(_06276_));
 sg13g2_a221oi_1 _14376_ (.B2(net5593),
    .C1(net5581),
    .B1(_06125_),
    .A1(_05965_),
    .Y(_06277_),
    .A2(_05995_));
 sg13g2_a21oi_1 _14377_ (.A1(_05964_),
    .A2(_06265_),
    .Y(_06278_),
    .B1(_06256_));
 sg13g2_nor3_1 _14378_ (.A(net5577),
    .B(_06277_),
    .C(_06278_),
    .Y(_06279_));
 sg13g2_nand4_1 _14379_ (.B(net5200),
    .C(_06172_),
    .A(_05961_),
    .Y(_06280_),
    .D(_06245_));
 sg13g2_a21oi_1 _14380_ (.A1(net5600),
    .A2(_06000_),
    .Y(_06281_),
    .B1(_06070_));
 sg13g2_o21ai_1 _14381_ (.B1(_06280_),
    .Y(_06282_),
    .A1(net5358),
    .A2(_06281_));
 sg13g2_or2_1 _14382_ (.X(_00017_),
    .B(_06282_),
    .A(_06279_));
 sg13g2_nand3_1 _14383_ (.B(_06006_),
    .C(_06174_),
    .A(net5597),
    .Y(_06283_));
 sg13g2_a21oi_1 _14384_ (.A1(_06061_),
    .A2(_06067_),
    .Y(_06284_),
    .B1(net5507));
 sg13g2_nand2_1 _14385_ (.Y(_06285_),
    .A(_06283_),
    .B(_06284_));
 sg13g2_a21oi_1 _14386_ (.A1(net5201),
    .A2(_06099_),
    .Y(_06286_),
    .B1(net5584));
 sg13g2_o21ai_1 _14387_ (.B1(_06285_),
    .Y(_06287_),
    .A1(net5199),
    .A2(_06286_));
 sg13g2_o21ai_1 _14388_ (.B1(net5502),
    .Y(_06288_),
    .A1(net5603),
    .A2(_05989_));
 sg13g2_a21oi_1 _14389_ (.A1(_05953_),
    .A2(_05978_),
    .Y(_06289_),
    .B1(_06021_));
 sg13g2_nand2_1 _14390_ (.Y(_06290_),
    .A(net5611),
    .B(net5603));
 sg13g2_a22oi_1 _14391_ (.Y(_06291_),
    .B1(_06290_),
    .B2(_05995_),
    .A2(_06065_),
    .A1(net5600));
 sg13g2_o21ai_1 _14392_ (.B1(_06287_),
    .Y(_06292_),
    .A1(net5358),
    .A2(_06291_));
 sg13g2_a21oi_1 _14393_ (.A1(_06288_),
    .A2(_06289_),
    .Y(_00018_),
    .B1(_06292_));
 sg13g2_nand2_1 _14394_ (.Y(_06293_),
    .A(_05984_),
    .B(_06097_));
 sg13g2_a21oi_1 _14395_ (.A1(_06134_),
    .A2(_06293_),
    .Y(_06294_),
    .B1(_06028_));
 sg13g2_a221oi_1 _14396_ (.B2(net5501),
    .C1(net5358),
    .B1(_05963_),
    .A1(_05953_),
    .Y(_06295_),
    .A2(_05958_));
 sg13g2_and3_1 _14397_ (.X(_06296_),
    .A(net5200),
    .B(_06095_),
    .C(_06172_));
 sg13g2_nor3_1 _14398_ (.A(net5589),
    .B(_05983_),
    .C(_06078_),
    .Y(_06297_));
 sg13g2_nand2_1 _14399_ (.Y(_06298_),
    .A(_06020_),
    .B(_06075_));
 sg13g2_nor2_1 _14400_ (.A(_06297_),
    .B(_06298_),
    .Y(_06299_));
 sg13g2_nor4_1 _14401_ (.A(_06294_),
    .B(_06295_),
    .C(_06296_),
    .D(_06299_),
    .Y(_00019_));
 sg13g2_o21ai_1 _14402_ (.B1(_05971_),
    .Y(_06300_),
    .A1(_05975_),
    .A2(_05980_));
 sg13g2_nor4_1 _14403_ (.A(net5583),
    .B(_05977_),
    .C(_05993_),
    .D(_06016_),
    .Y(_06301_));
 sg13g2_nor2_1 _14404_ (.A(_05970_),
    .B(_06219_),
    .Y(_06302_));
 sg13g2_nand2b_1 _14405_ (.Y(_06303_),
    .B(_05982_),
    .A_N(_06297_));
 sg13g2_nand3_1 _14406_ (.B(_06080_),
    .C(_06090_),
    .A(net5581),
    .Y(_06304_));
 sg13g2_nand2_1 _14407_ (.Y(_06305_),
    .A(_06303_),
    .B(_06304_));
 sg13g2_nor3_1 _14408_ (.A(net5506),
    .B(_06301_),
    .C(_06302_),
    .Y(_06306_));
 sg13g2_a22oi_1 _14409_ (.Y(_00020_),
    .B1(_06306_),
    .B2(_06300_),
    .A2(_06305_),
    .A1(net5505));
 sg13g2_nor2_1 _14410_ (.A(_06154_),
    .B(_06251_),
    .Y(_06307_));
 sg13g2_nor2_1 _14411_ (.A(net5584),
    .B(_06307_),
    .Y(_06308_));
 sg13g2_nor3_1 _14412_ (.A(_06152_),
    .B(_06229_),
    .C(_06308_),
    .Y(_06309_));
 sg13g2_nand3_1 _14413_ (.B(_06006_),
    .C(_06082_),
    .A(net5596),
    .Y(_06310_));
 sg13g2_a21oi_1 _14414_ (.A1(_06004_),
    .A2(_06046_),
    .Y(_06311_),
    .B1(net5358));
 sg13g2_a21o_1 _14415_ (.A2(_00132_),
    .A1(net5499),
    .B1(_06145_),
    .X(_06312_));
 sg13g2_a22oi_1 _14416_ (.Y(_06313_),
    .B1(_06312_),
    .B2(net5199),
    .A2(_06311_),
    .A1(_06310_));
 sg13g2_o21ai_1 _14417_ (.B1(_06313_),
    .Y(_00021_),
    .A1(net5578),
    .A2(_06309_));
 sg13g2_nand3_1 _14418_ (.B(_06005_),
    .C(_06144_),
    .A(net5592),
    .Y(_06314_));
 sg13g2_nand3_1 _14419_ (.B(_06259_),
    .C(_06314_),
    .A(net5581),
    .Y(_06315_));
 sg13g2_a21oi_1 _14420_ (.A1(_05965_),
    .A2(_06035_),
    .Y(_06316_),
    .B1(net5505));
 sg13g2_o21ai_1 _14421_ (.B1(_06315_),
    .Y(_06317_),
    .A1(net5198),
    .A2(_06316_));
 sg13g2_a21oi_1 _14422_ (.A1(net5501),
    .A2(_05988_),
    .Y(_06318_),
    .B1(net5581));
 sg13g2_o21ai_1 _14423_ (.B1(_06318_),
    .Y(_06319_),
    .A1(net5099),
    .A2(_06047_));
 sg13g2_o21ai_1 _14424_ (.B1(_06319_),
    .Y(_06320_),
    .A1(_06155_),
    .A2(_06238_));
 sg13g2_o21ai_1 _14425_ (.B1(_06317_),
    .Y(_00023_),
    .A1(net5577),
    .A2(_06320_));
 sg13g2_o21ai_1 _14426_ (.B1(_06001_),
    .Y(_06321_),
    .A1(net5594),
    .A2(_05977_));
 sg13g2_nand3_1 _14427_ (.B(_06014_),
    .C(_06055_),
    .A(net5590),
    .Y(_06322_));
 sg13g2_a221oi_1 _14428_ (.B2(_06037_),
    .C1(net5577),
    .B1(_06322_),
    .A1(net5582),
    .Y(_06323_),
    .A2(_06321_));
 sg13g2_o21ai_1 _14429_ (.B1(net5594),
    .Y(_06324_),
    .A1(net5603),
    .A2(_05984_));
 sg13g2_a21oi_1 _14430_ (.A1(_06080_),
    .A2(_06324_),
    .Y(_06325_),
    .B1(_06040_));
 sg13g2_nor2_1 _14431_ (.A(_06323_),
    .B(_06325_),
    .Y(_06326_));
 sg13g2_o21ai_1 _14432_ (.B1(_06326_),
    .Y(_00024_),
    .A1(_06025_),
    .A2(_06050_));
 sg13g2_xnor2_1 _14433_ (.Y(_06327_),
    .A(net3394),
    .B(\TRNG.NOISE_SAMPLER.Sample_Out ));
 sg13g2_xor2_1 _14434_ (.B(\TRNG.NOISE_SAMPLER.Sample_Out ),
    .A(net3937),
    .X(_06328_));
 sg13g2_nand2_1 _14435_ (.Y(_00096_),
    .A(net1257),
    .B(_06327_));
 sg13g2_and2_1 _14436_ (.A(net2312),
    .B(net1257),
    .X(_06329_));
 sg13g2_nor2_1 _14437_ (.A(net2312),
    .B(net1257),
    .Y(_06330_));
 sg13g2_nor3_1 _14438_ (.A(_06328_),
    .B(_06329_),
    .C(_06330_),
    .Y(_00097_));
 sg13g2_o21ai_1 _14439_ (.B1(_06327_),
    .Y(_06331_),
    .A1(net2368),
    .A2(_06329_));
 sg13g2_a21oi_1 _14440_ (.A1(net2368),
    .A2(_06329_),
    .Y(_00098_),
    .B1(_06331_));
 sg13g2_and3_1 _14441_ (.X(_06332_),
    .A(net1405),
    .B(net2368),
    .C(_06329_));
 sg13g2_a21oi_1 _14442_ (.A1(\TRNG.Repetition_Count_Test.count[2] ),
    .A2(_06329_),
    .Y(_06333_),
    .B1(net1405));
 sg13g2_nor3_1 _14443_ (.A(_06328_),
    .B(_06332_),
    .C(net1406),
    .Y(_00099_));
 sg13g2_and2_1 _14444_ (.A(net3370),
    .B(_06332_),
    .X(_06334_));
 sg13g2_o21ai_1 _14445_ (.B1(_06327_),
    .Y(_06335_),
    .A1(net3370),
    .A2(_06332_));
 sg13g2_nor2_1 _14446_ (.A(_06334_),
    .B(_06335_),
    .Y(_00100_));
 sg13g2_a21oi_1 _14447_ (.A1(net3149),
    .A2(_06334_),
    .Y(_06336_),
    .B1(_06328_));
 sg13g2_o21ai_1 _14448_ (.B1(_06336_),
    .Y(_06337_),
    .A1(net3149),
    .A2(_06334_));
 sg13g2_inv_1 _14449_ (.Y(_00101_),
    .A(_06337_));
 sg13g2_nand2_1 _14450_ (.Y(\TRNG.NOISE_SOURCE.Loop1.NOT2_OUT_TO_NAND1_IN2 ),
    .A(net5898),
    .B(\TRNG.NOISE_SOURCE.Loop1.NOT2_OUT_TO_NAND1_IN2 ));
 sg13g2_nand2_1 _14451_ (.Y(\TRNG.NOISE_SOURCE.Loop2.NOT2_OUT_TO_NAND1_IN2 ),
    .A(net5898),
    .B(\TRNG.NOISE_SOURCE.Loop2.NOT2_OUT_TO_NAND1_IN2 ));
 sg13g2_nand2_1 _14452_ (.Y(\TRNG.NOISE_SOURCE.Loop3.NOT2_OUT_TO_NAND1_IN2 ),
    .A(net5898),
    .B(\TRNG.NOISE_SOURCE.Loop3.NOT2_OUT_TO_NAND1_IN2 ));
 sg13g2_nand2_1 _14453_ (.Y(\TRNG.NOISE_SOURCE.Loop4.NOT2_OUT_TO_NAND1_IN2 ),
    .A(net5898),
    .B(\TRNG.NOISE_SOURCE.Loop4.NOT2_OUT_TO_NAND1_IN2 ));
 sg13g2_nand2_1 _14454_ (.Y(\TRNG.NOISE_SOURCE.Loop5.NOT2_OUT_TO_NAND1_IN2 ),
    .A(net5898),
    .B(\TRNG.NOISE_SOURCE.Loop5.NOT2_OUT_TO_NAND1_IN2 ));
 sg13g2_xnor2_1 _14455_ (.Y(_06338_),
    .A(\TRNG.sha256.expand.dout2[17] ),
    .B(\TRNG.sha256.expand.dout2[10] ));
 sg13g2_xnor2_1 _14456_ (.Y(_06339_),
    .A(\TRNG.sha256.expand.dout2[19] ),
    .B(_06338_));
 sg13g2_xnor2_1 _14457_ (.Y(_06340_),
    .A(\TRNG.sha256.expand.dout1[7] ),
    .B(\TRNG.sha256.expand.dout1[3] ));
 sg13g2_xnor2_1 _14458_ (.Y(_06341_),
    .A(\TRNG.sha256.expand.dout1[18] ),
    .B(_06340_));
 sg13g2_nand2_1 _14459_ (.Y(_06342_),
    .A(_06339_),
    .B(_06341_));
 sg13g2_xor2_1 _14460_ (.B(_06341_),
    .A(_06339_),
    .X(_00238_));
 sg13g2_xnor2_1 _14461_ (.Y(_06343_),
    .A(\TRNG.sha256.expand.dout2[18] ),
    .B(\TRNG.sha256.expand.dout2[11] ));
 sg13g2_xnor2_1 _14462_ (.Y(_06344_),
    .A(\TRNG.sha256.expand.dout2[20] ),
    .B(_06343_));
 sg13g2_xnor2_1 _14463_ (.Y(_06345_),
    .A(\TRNG.sha256.expand.dout1[8] ),
    .B(\TRNG.sha256.expand.dout1[4] ));
 sg13g2_xnor2_1 _14464_ (.Y(_06346_),
    .A(\TRNG.sha256.expand.dout1[19] ),
    .B(_06345_));
 sg13g2_nand2_1 _14465_ (.Y(_06347_),
    .A(_06344_),
    .B(_06346_));
 sg13g2_xnor2_1 _14466_ (.Y(_06348_),
    .A(_06344_),
    .B(_06346_));
 sg13g2_xor2_1 _14467_ (.B(_06348_),
    .A(_06342_),
    .X(_00249_));
 sg13g2_o21ai_1 _14468_ (.B1(_06347_),
    .Y(_06349_),
    .A1(_06342_),
    .A2(_06348_));
 sg13g2_xnor2_1 _14469_ (.Y(_06350_),
    .A(\TRNG.sha256.expand.dout2[21] ),
    .B(\TRNG.sha256.expand.dout2[12] ));
 sg13g2_xnor2_1 _14470_ (.Y(_06351_),
    .A(\TRNG.sha256.expand.dout2[19] ),
    .B(_06350_));
 sg13g2_xnor2_1 _14471_ (.Y(_06352_),
    .A(\TRNG.sha256.expand.dout1[9] ),
    .B(\TRNG.sha256.expand.dout1[5] ));
 sg13g2_xnor2_1 _14472_ (.Y(_06353_),
    .A(\TRNG.sha256.expand.dout1[20] ),
    .B(_06352_));
 sg13g2_and2_1 _14473_ (.A(_06351_),
    .B(_06353_),
    .X(_06354_));
 sg13g2_or2_1 _14474_ (.X(_06355_),
    .B(_06353_),
    .A(_06351_));
 sg13g2_nand2b_1 _14475_ (.Y(_06356_),
    .B(_06355_),
    .A_N(_06354_));
 sg13g2_xnor2_1 _14476_ (.Y(_00260_),
    .A(_06349_),
    .B(_06356_));
 sg13g2_a21o_1 _14477_ (.A2(_06355_),
    .A1(_06349_),
    .B1(_06354_),
    .X(_06357_));
 sg13g2_xnor2_1 _14478_ (.Y(_06358_),
    .A(\TRNG.sha256.expand.dout2[22] ),
    .B(\TRNG.sha256.expand.dout2[13] ));
 sg13g2_xnor2_1 _14479_ (.Y(_06359_),
    .A(\TRNG.sha256.expand.dout2[20] ),
    .B(_06358_));
 sg13g2_xnor2_1 _14480_ (.Y(_06360_),
    .A(\TRNG.sha256.expand.dout1[10] ),
    .B(\TRNG.sha256.expand.dout1[6] ));
 sg13g2_xnor2_1 _14481_ (.Y(_06361_),
    .A(\TRNG.sha256.expand.dout1[21] ),
    .B(_06360_));
 sg13g2_and2_1 _14482_ (.A(_06359_),
    .B(_06361_),
    .X(_06362_));
 sg13g2_xor2_1 _14483_ (.B(_06361_),
    .A(_06359_),
    .X(_06363_));
 sg13g2_xor2_1 _14484_ (.B(_06363_),
    .A(_06357_),
    .X(_00263_));
 sg13g2_a21oi_1 _14485_ (.A1(_06357_),
    .A2(_06363_),
    .Y(_06364_),
    .B1(_06362_));
 sg13g2_xnor2_1 _14486_ (.Y(_06365_),
    .A(\TRNG.sha256.expand.dout2[23] ),
    .B(\TRNG.sha256.expand.dout2[14] ));
 sg13g2_xnor2_1 _14487_ (.Y(_06366_),
    .A(\TRNG.sha256.expand.dout2[21] ),
    .B(_06365_));
 sg13g2_xnor2_1 _14488_ (.Y(_06367_),
    .A(\TRNG.sha256.expand.dout1[22] ),
    .B(\TRNG.sha256.expand.dout1[11] ));
 sg13g2_xnor2_1 _14489_ (.Y(_06368_),
    .A(\TRNG.sha256.expand.dout1[7] ),
    .B(_06367_));
 sg13g2_nand2_1 _14490_ (.Y(_06369_),
    .A(_06366_),
    .B(_06368_));
 sg13g2_xnor2_1 _14491_ (.Y(_06370_),
    .A(_06366_),
    .B(_06368_));
 sg13g2_xor2_1 _14492_ (.B(_06370_),
    .A(_06364_),
    .X(_00264_));
 sg13g2_o21ai_1 _14493_ (.B1(_06369_),
    .Y(_06371_),
    .A1(_06364_),
    .A2(_06370_));
 sg13g2_xnor2_1 _14494_ (.Y(_06372_),
    .A(\TRNG.sha256.expand.dout2[24] ),
    .B(\TRNG.sha256.expand.dout2[15] ));
 sg13g2_xnor2_1 _14495_ (.Y(_06373_),
    .A(\TRNG.sha256.expand.dout2[22] ),
    .B(_06372_));
 sg13g2_xnor2_1 _14496_ (.Y(_06374_),
    .A(\TRNG.sha256.expand.dout1[23] ),
    .B(\TRNG.sha256.expand.dout1[12] ));
 sg13g2_xnor2_1 _14497_ (.Y(_06375_),
    .A(\TRNG.sha256.expand.dout1[8] ),
    .B(_06374_));
 sg13g2_and2_1 _14498_ (.A(_06373_),
    .B(_06375_),
    .X(_06376_));
 sg13g2_xor2_1 _14499_ (.B(_06375_),
    .A(_06373_),
    .X(_06377_));
 sg13g2_xor2_1 _14500_ (.B(_06377_),
    .A(_06371_),
    .X(_00265_));
 sg13g2_a21oi_1 _14501_ (.A1(_06371_),
    .A2(_06377_),
    .Y(_06378_),
    .B1(_06376_));
 sg13g2_xnor2_1 _14502_ (.Y(_06379_),
    .A(\TRNG.sha256.expand.dout2[25] ),
    .B(\TRNG.sha256.expand.dout2[16] ));
 sg13g2_xnor2_1 _14503_ (.Y(_06380_),
    .A(\TRNG.sha256.expand.dout2[23] ),
    .B(_06379_));
 sg13g2_xnor2_1 _14504_ (.Y(_06381_),
    .A(\TRNG.sha256.expand.dout1[24] ),
    .B(\TRNG.sha256.expand.dout1[13] ));
 sg13g2_xnor2_1 _14505_ (.Y(_06382_),
    .A(\TRNG.sha256.expand.dout1[9] ),
    .B(_06381_));
 sg13g2_nand2_1 _14506_ (.Y(_06383_),
    .A(_06380_),
    .B(_06382_));
 sg13g2_xnor2_1 _14507_ (.Y(_06384_),
    .A(_06380_),
    .B(_06382_));
 sg13g2_xor2_1 _14508_ (.B(_06384_),
    .A(_06378_),
    .X(_00266_));
 sg13g2_o21ai_1 _14509_ (.B1(_06383_),
    .Y(_06385_),
    .A1(_06378_),
    .A2(_06384_));
 sg13g2_xnor2_1 _14510_ (.Y(_06386_),
    .A(\TRNG.sha256.expand.dout2[24] ),
    .B(\TRNG.sha256.expand.dout2[26] ));
 sg13g2_xnor2_1 _14511_ (.Y(_06387_),
    .A(\TRNG.sha256.expand.dout2[17] ),
    .B(_06386_));
 sg13g2_xnor2_1 _14512_ (.Y(_06388_),
    .A(\TRNG.sha256.expand.dout1[25] ),
    .B(\TRNG.sha256.expand.dout1[14] ));
 sg13g2_xnor2_1 _14513_ (.Y(_06389_),
    .A(\TRNG.sha256.expand.dout1[10] ),
    .B(_06388_));
 sg13g2_nand2_1 _14514_ (.Y(_06390_),
    .A(_06387_),
    .B(_06389_));
 sg13g2_inv_1 _14515_ (.Y(_06391_),
    .A(_06390_));
 sg13g2_xor2_1 _14516_ (.B(_06389_),
    .A(_06387_),
    .X(_06392_));
 sg13g2_xor2_1 _14517_ (.B(_06392_),
    .A(_06385_),
    .X(_00267_));
 sg13g2_xnor2_1 _14518_ (.Y(_06393_),
    .A(\TRNG.sha256.expand.dout2[25] ),
    .B(\TRNG.sha256.expand.dout2[27] ));
 sg13g2_xnor2_1 _14519_ (.Y(_06394_),
    .A(\TRNG.sha256.expand.dout2[18] ),
    .B(_06393_));
 sg13g2_xnor2_1 _14520_ (.Y(_06395_),
    .A(\TRNG.sha256.expand.dout1[26] ),
    .B(\TRNG.sha256.expand.dout1[15] ));
 sg13g2_xnor2_1 _14521_ (.Y(_06396_),
    .A(\TRNG.sha256.expand.dout1[11] ),
    .B(_06395_));
 sg13g2_nand2_1 _14522_ (.Y(_06397_),
    .A(_06394_),
    .B(_06396_));
 sg13g2_xnor2_1 _14523_ (.Y(_06398_),
    .A(_06394_),
    .B(_06396_));
 sg13g2_a21oi_2 _14524_ (.B1(_06391_),
    .Y(_06399_),
    .A2(_06392_),
    .A1(_06385_));
 sg13g2_xor2_1 _14525_ (.B(_06399_),
    .A(_06398_),
    .X(_00268_));
 sg13g2_xnor2_1 _14526_ (.Y(_06400_),
    .A(\TRNG.sha256.expand.dout2[26] ),
    .B(\TRNG.sha256.expand.dout2[28] ));
 sg13g2_xnor2_1 _14527_ (.Y(_06401_),
    .A(\TRNG.sha256.expand.dout2[19] ),
    .B(_06400_));
 sg13g2_xnor2_1 _14528_ (.Y(_06402_),
    .A(\TRNG.sha256.expand.dout1[27] ),
    .B(\TRNG.sha256.expand.dout1[16] ));
 sg13g2_xnor2_1 _14529_ (.Y(_06403_),
    .A(\TRNG.sha256.expand.dout1[12] ),
    .B(_06402_));
 sg13g2_nor2_1 _14530_ (.A(_06401_),
    .B(_06403_),
    .Y(_06404_));
 sg13g2_nand2_1 _14531_ (.Y(_06405_),
    .A(_06401_),
    .B(_06403_));
 sg13g2_nand2b_1 _14532_ (.Y(_06406_),
    .B(_06405_),
    .A_N(_06404_));
 sg13g2_o21ai_1 _14533_ (.B1(_06397_),
    .Y(_06407_),
    .A1(_06398_),
    .A2(_06399_));
 sg13g2_xnor2_1 _14534_ (.Y(_00269_),
    .A(_06406_),
    .B(_06407_));
 sg13g2_xnor2_1 _14535_ (.Y(_06408_),
    .A(\TRNG.sha256.expand.dout2[27] ),
    .B(\TRNG.sha256.expand.dout2[29] ));
 sg13g2_xnor2_1 _14536_ (.Y(_06409_),
    .A(\TRNG.sha256.expand.dout2[20] ),
    .B(_06408_));
 sg13g2_xnor2_1 _14537_ (.Y(_06410_),
    .A(\TRNG.sha256.expand.dout1[28] ),
    .B(\TRNG.sha256.expand.dout1[17] ));
 sg13g2_xnor2_1 _14538_ (.Y(_06411_),
    .A(\TRNG.sha256.expand.dout1[13] ),
    .B(_06410_));
 sg13g2_and2_1 _14539_ (.A(_06409_),
    .B(_06411_),
    .X(_06412_));
 sg13g2_xnor2_1 _14540_ (.Y(_06413_),
    .A(_06409_),
    .B(_06411_));
 sg13g2_inv_1 _14541_ (.Y(_06414_),
    .A(_06413_));
 sg13g2_and2_1 _14542_ (.A(_06397_),
    .B(_06405_),
    .X(_06415_));
 sg13g2_o21ai_1 _14543_ (.B1(_06415_),
    .Y(_06416_),
    .A1(_06398_),
    .A2(_06399_));
 sg13g2_nor2b_1 _14544_ (.A(_06404_),
    .B_N(_06416_),
    .Y(_06417_));
 sg13g2_nand3b_1 _14545_ (.B(_06414_),
    .C(_06416_),
    .Y(_06418_),
    .A_N(_06404_));
 sg13g2_xnor2_1 _14546_ (.Y(_00239_),
    .A(_06413_),
    .B(_06417_));
 sg13g2_nor2b_1 _14547_ (.A(_06412_),
    .B_N(_06418_),
    .Y(_06419_));
 sg13g2_xnor2_1 _14548_ (.Y(_06420_),
    .A(\TRNG.sha256.expand.dout2[28] ),
    .B(\TRNG.sha256.expand.dout2[30] ));
 sg13g2_xnor2_1 _14549_ (.Y(_06421_),
    .A(\TRNG.sha256.expand.dout2[21] ),
    .B(_06420_));
 sg13g2_inv_1 _14550_ (.Y(_06422_),
    .A(_06421_));
 sg13g2_xnor2_1 _14551_ (.Y(_06423_),
    .A(\TRNG.sha256.expand.dout1[14] ),
    .B(\TRNG.sha256.expand.dout1[29] ));
 sg13g2_xnor2_1 _14552_ (.Y(_06424_),
    .A(\TRNG.sha256.expand.dout1[18] ),
    .B(_06423_));
 sg13g2_inv_1 _14553_ (.Y(_06425_),
    .A(_06424_));
 sg13g2_nand2_1 _14554_ (.Y(_06426_),
    .A(_06422_),
    .B(_06425_));
 sg13g2_nand2_1 _14555_ (.Y(_06427_),
    .A(_06421_),
    .B(_06424_));
 sg13g2_nor2b_1 _14556_ (.A(_06412_),
    .B_N(_06427_),
    .Y(_06428_));
 sg13g2_nand2_1 _14557_ (.Y(_06429_),
    .A(_06418_),
    .B(_06428_));
 sg13g2_nand2_1 _14558_ (.Y(_06430_),
    .A(_06426_),
    .B(_06429_));
 sg13g2_nand2_1 _14559_ (.Y(_06431_),
    .A(_06426_),
    .B(_06427_));
 sg13g2_xor2_1 _14560_ (.B(_06431_),
    .A(_06419_),
    .X(_00240_));
 sg13g2_xnor2_1 _14561_ (.Y(_06432_),
    .A(\TRNG.sha256.expand.dout2[29] ),
    .B(\TRNG.sha256.expand.dout2[31] ));
 sg13g2_xnor2_1 _14562_ (.Y(_06433_),
    .A(\TRNG.sha256.expand.dout2[22] ),
    .B(_06432_));
 sg13g2_xnor2_1 _14563_ (.Y(_06434_),
    .A(\TRNG.sha256.expand.dout1[15] ),
    .B(\TRNG.sha256.expand.dout1[30] ));
 sg13g2_xnor2_1 _14564_ (.Y(_06435_),
    .A(\TRNG.sha256.expand.dout1[19] ),
    .B(_06434_));
 sg13g2_nand2_1 _14565_ (.Y(_06436_),
    .A(_06433_),
    .B(_06435_));
 sg13g2_xnor2_1 _14566_ (.Y(_06437_),
    .A(_06433_),
    .B(_06435_));
 sg13g2_xor2_1 _14567_ (.B(_06437_),
    .A(_06430_),
    .X(_00241_));
 sg13g2_o21ai_1 _14568_ (.B1(_06436_),
    .Y(_06438_),
    .A1(_06430_),
    .A2(_06437_));
 sg13g2_xnor2_1 _14569_ (.Y(_06439_),
    .A(\TRNG.sha256.expand.dout2[30] ),
    .B(\TRNG.sha256.expand.dout2[0] ));
 sg13g2_xnor2_1 _14570_ (.Y(_06440_),
    .A(\TRNG.sha256.expand.dout2[23] ),
    .B(_06439_));
 sg13g2_xnor2_1 _14571_ (.Y(_06441_),
    .A(\TRNG.sha256.expand.dout1[16] ),
    .B(\TRNG.sha256.expand.dout1[31] ));
 sg13g2_xnor2_1 _14572_ (.Y(_06442_),
    .A(\TRNG.sha256.expand.dout1[20] ),
    .B(_06441_));
 sg13g2_nand2_1 _14573_ (.Y(_06443_),
    .A(_06440_),
    .B(_06442_));
 sg13g2_nor2_1 _14574_ (.A(_06440_),
    .B(_06442_),
    .Y(_06444_));
 sg13g2_inv_1 _14575_ (.Y(_06445_),
    .A(_06444_));
 sg13g2_nand2_1 _14576_ (.Y(_06446_),
    .A(_06443_),
    .B(_06445_));
 sg13g2_xnor2_1 _14577_ (.Y(_00242_),
    .A(_06438_),
    .B(_06446_));
 sg13g2_xnor2_1 _14578_ (.Y(_06447_),
    .A(\TRNG.sha256.expand.dout2[31] ),
    .B(\TRNG.sha256.expand.dout2[1] ));
 sg13g2_xnor2_1 _14579_ (.Y(_06448_),
    .A(\TRNG.sha256.expand.dout2[24] ),
    .B(_06447_));
 sg13g2_xnor2_1 _14580_ (.Y(_06449_),
    .A(\TRNG.sha256.expand.dout1[17] ),
    .B(\TRNG.sha256.expand.dout1[0] ));
 sg13g2_xnor2_1 _14581_ (.Y(_06450_),
    .A(\TRNG.sha256.expand.dout1[21] ),
    .B(_06449_));
 sg13g2_nand2_1 _14582_ (.Y(_06451_),
    .A(_06448_),
    .B(_06450_));
 sg13g2_xnor2_1 _14583_ (.Y(_06452_),
    .A(_06448_),
    .B(_06450_));
 sg13g2_or2_1 _14584_ (.X(_06453_),
    .B(_06446_),
    .A(_06437_));
 sg13g2_a221oi_1 _14585_ (.B2(_06418_),
    .C1(_06453_),
    .B1(_06428_),
    .A1(_06422_),
    .Y(_06454_),
    .A2(_06425_));
 sg13g2_o21ai_1 _14586_ (.B1(_06443_),
    .Y(_06455_),
    .A1(_06436_),
    .A2(_06444_));
 sg13g2_nor2_1 _14587_ (.A(_06454_),
    .B(_06455_),
    .Y(_06456_));
 sg13g2_xor2_1 _14588_ (.B(_06456_),
    .A(_06452_),
    .X(_00243_));
 sg13g2_o21ai_1 _14589_ (.B1(_06451_),
    .Y(_06457_),
    .A1(_06452_),
    .A2(_06456_));
 sg13g2_xnor2_1 _14590_ (.Y(_06458_),
    .A(\TRNG.sha256.expand.dout2[0] ),
    .B(\TRNG.sha256.expand.dout2[2] ));
 sg13g2_xnor2_1 _14591_ (.Y(_06459_),
    .A(\TRNG.sha256.expand.dout2[25] ),
    .B(_06458_));
 sg13g2_xnor2_1 _14592_ (.Y(_06460_),
    .A(\TRNG.sha256.expand.dout1[22] ),
    .B(\TRNG.sha256.expand.dout1[1] ));
 sg13g2_xnor2_1 _14593_ (.Y(_06461_),
    .A(\TRNG.sha256.expand.dout1[18] ),
    .B(_06460_));
 sg13g2_nor2_1 _14594_ (.A(_06459_),
    .B(_06461_),
    .Y(_06462_));
 sg13g2_and2_1 _14595_ (.A(_06459_),
    .B(_06461_),
    .X(_06463_));
 sg13g2_or2_1 _14596_ (.X(_06464_),
    .B(_06463_),
    .A(_06462_));
 sg13g2_xnor2_1 _14597_ (.Y(_00244_),
    .A(_06457_),
    .B(_06464_));
 sg13g2_nor2_1 _14598_ (.A(_06452_),
    .B(_06464_),
    .Y(_06465_));
 sg13g2_o21ai_1 _14599_ (.B1(_06465_),
    .Y(_06466_),
    .A1(_06454_),
    .A2(_06455_));
 sg13g2_nor2_1 _14600_ (.A(_06451_),
    .B(_06462_),
    .Y(_06467_));
 sg13g2_nor2_1 _14601_ (.A(_06463_),
    .B(_06467_),
    .Y(_06468_));
 sg13g2_nand2_1 _14602_ (.Y(_06469_),
    .A(_06466_),
    .B(_06468_));
 sg13g2_inv_1 _14603_ (.Y(_06470_),
    .A(_06469_));
 sg13g2_xnor2_1 _14604_ (.Y(_06471_),
    .A(\TRNG.sha256.expand.dout2[1] ),
    .B(\TRNG.sha256.expand.dout2[3] ));
 sg13g2_xnor2_1 _14605_ (.Y(_06472_),
    .A(\TRNG.sha256.expand.dout2[26] ),
    .B(_06471_));
 sg13g2_xnor2_1 _14606_ (.Y(_06473_),
    .A(\TRNG.sha256.expand.dout1[23] ),
    .B(\TRNG.sha256.expand.dout1[2] ));
 sg13g2_xnor2_1 _14607_ (.Y(_06474_),
    .A(\TRNG.sha256.expand.dout1[19] ),
    .B(_06473_));
 sg13g2_nand2_1 _14608_ (.Y(_06475_),
    .A(_06472_),
    .B(_06474_));
 sg13g2_xnor2_1 _14609_ (.Y(_06476_),
    .A(_06472_),
    .B(_06474_));
 sg13g2_xnor2_1 _14610_ (.Y(_00245_),
    .A(_06469_),
    .B(_06476_));
 sg13g2_xnor2_1 _14611_ (.Y(_06477_),
    .A(\TRNG.sha256.expand.dout2[2] ),
    .B(\TRNG.sha256.expand.dout2[4] ));
 sg13g2_xnor2_1 _14612_ (.Y(_06478_),
    .A(\TRNG.sha256.expand.dout2[27] ),
    .B(_06477_));
 sg13g2_xnor2_1 _14613_ (.Y(_06479_),
    .A(\TRNG.sha256.expand.dout1[20] ),
    .B(\TRNG.sha256.expand.dout1[24] ));
 sg13g2_xnor2_1 _14614_ (.Y(_06480_),
    .A(\TRNG.sha256.expand.dout1[3] ),
    .B(_06479_));
 sg13g2_nand2_1 _14615_ (.Y(_06481_),
    .A(_06478_),
    .B(_06480_));
 sg13g2_nor2_1 _14616_ (.A(_06478_),
    .B(_06480_),
    .Y(_06482_));
 sg13g2_xnor2_1 _14617_ (.Y(_06483_),
    .A(_06478_),
    .B(_06480_));
 sg13g2_o21ai_1 _14618_ (.B1(_06475_),
    .Y(_06484_),
    .A1(_06470_),
    .A2(_06476_));
 sg13g2_xnor2_1 _14619_ (.Y(_00246_),
    .A(_06483_),
    .B(_06484_));
 sg13g2_or2_1 _14620_ (.X(_06485_),
    .B(_06483_),
    .A(_06476_));
 sg13g2_a21oi_1 _14621_ (.A1(_06466_),
    .A2(_06468_),
    .Y(_06486_),
    .B1(_06485_));
 sg13g2_o21ai_1 _14622_ (.B1(_06481_),
    .Y(_06487_),
    .A1(_06475_),
    .A2(_06482_));
 sg13g2_nor2_1 _14623_ (.A(_06486_),
    .B(_06487_),
    .Y(_06488_));
 sg13g2_xnor2_1 _14624_ (.Y(_06489_),
    .A(\TRNG.sha256.expand.dout2[3] ),
    .B(\TRNG.sha256.expand.dout2[5] ));
 sg13g2_xnor2_1 _14625_ (.Y(_06490_),
    .A(\TRNG.sha256.expand.dout2[28] ),
    .B(_06489_));
 sg13g2_xnor2_1 _14626_ (.Y(_06491_),
    .A(\TRNG.sha256.expand.dout1[21] ),
    .B(\TRNG.sha256.expand.dout1[25] ));
 sg13g2_xnor2_1 _14627_ (.Y(_06492_),
    .A(\TRNG.sha256.expand.dout1[4] ),
    .B(_06491_));
 sg13g2_nand2_1 _14628_ (.Y(_06493_),
    .A(_06490_),
    .B(_06492_));
 sg13g2_xnor2_1 _14629_ (.Y(_06494_),
    .A(_06490_),
    .B(_06492_));
 sg13g2_xor2_1 _14630_ (.B(_06494_),
    .A(_06488_),
    .X(_00247_));
 sg13g2_xnor2_1 _14631_ (.Y(_06495_),
    .A(\TRNG.sha256.expand.dout2[4] ),
    .B(\TRNG.sha256.expand.dout2[6] ));
 sg13g2_xnor2_1 _14632_ (.Y(_06496_),
    .A(\TRNG.sha256.expand.dout2[29] ),
    .B(_06495_));
 sg13g2_xnor2_1 _14633_ (.Y(_06497_),
    .A(\TRNG.sha256.expand.dout1[22] ),
    .B(\TRNG.sha256.expand.dout1[26] ));
 sg13g2_xnor2_1 _14634_ (.Y(_06498_),
    .A(\TRNG.sha256.expand.dout1[5] ),
    .B(_06497_));
 sg13g2_and2_1 _14635_ (.A(_06496_),
    .B(_06498_),
    .X(_06499_));
 sg13g2_nor2_1 _14636_ (.A(_06496_),
    .B(_06498_),
    .Y(_06500_));
 sg13g2_or2_1 _14637_ (.X(_06501_),
    .B(_06500_),
    .A(_06499_));
 sg13g2_o21ai_1 _14638_ (.B1(_06493_),
    .Y(_06502_),
    .A1(_06488_),
    .A2(_06494_));
 sg13g2_xnor2_1 _14639_ (.Y(_00248_),
    .A(_06501_),
    .B(_06502_));
 sg13g2_nor2_1 _14640_ (.A(_06494_),
    .B(_06501_),
    .Y(_06503_));
 sg13g2_o21ai_1 _14641_ (.B1(_06503_),
    .Y(_06504_),
    .A1(_06486_),
    .A2(_06487_));
 sg13g2_nor2_1 _14642_ (.A(_06493_),
    .B(_06500_),
    .Y(_06505_));
 sg13g2_nor2_1 _14643_ (.A(_06499_),
    .B(_06505_),
    .Y(_06506_));
 sg13g2_and2_1 _14644_ (.A(_06504_),
    .B(_06506_),
    .X(_06507_));
 sg13g2_xnor2_1 _14645_ (.Y(_06508_),
    .A(\TRNG.sha256.expand.dout2[5] ),
    .B(\TRNG.sha256.expand.dout2[7] ));
 sg13g2_xnor2_1 _14646_ (.Y(_06509_),
    .A(\TRNG.sha256.expand.dout2[30] ),
    .B(_06508_));
 sg13g2_xnor2_1 _14647_ (.Y(_06510_),
    .A(\TRNG.sha256.expand.dout1[23] ),
    .B(\TRNG.sha256.expand.dout1[27] ));
 sg13g2_xnor2_1 _14648_ (.Y(_06511_),
    .A(\TRNG.sha256.expand.dout1[6] ),
    .B(_06510_));
 sg13g2_nand2_1 _14649_ (.Y(_06512_),
    .A(_06509_),
    .B(_06511_));
 sg13g2_xnor2_1 _14650_ (.Y(_06513_),
    .A(_06509_),
    .B(_06511_));
 sg13g2_xor2_1 _14651_ (.B(_06513_),
    .A(_06507_),
    .X(_00250_));
 sg13g2_xnor2_1 _14652_ (.Y(_06514_),
    .A(\TRNG.sha256.expand.dout2[6] ),
    .B(\TRNG.sha256.expand.dout2[8] ));
 sg13g2_xnor2_1 _14653_ (.Y(_06515_),
    .A(\TRNG.sha256.expand.dout2[31] ),
    .B(_06514_));
 sg13g2_xnor2_1 _14654_ (.Y(_06516_),
    .A(\TRNG.sha256.expand.dout1[24] ),
    .B(\TRNG.sha256.expand.dout1[28] ));
 sg13g2_xnor2_1 _14655_ (.Y(_06517_),
    .A(\TRNG.sha256.expand.dout1[7] ),
    .B(_06516_));
 sg13g2_nand2_1 _14656_ (.Y(_06518_),
    .A(_06515_),
    .B(_06517_));
 sg13g2_xnor2_1 _14657_ (.Y(_06519_),
    .A(_06515_),
    .B(_06517_));
 sg13g2_o21ai_1 _14658_ (.B1(_06512_),
    .Y(_06520_),
    .A1(_06507_),
    .A2(_06513_));
 sg13g2_or2_1 _14659_ (.X(_06521_),
    .B(_06519_),
    .A(_06513_));
 sg13g2_a21oi_1 _14660_ (.A1(_06504_),
    .A2(_06506_),
    .Y(_06522_),
    .B1(_06521_));
 sg13g2_xnor2_1 _14661_ (.Y(_00251_),
    .A(_06519_),
    .B(_06520_));
 sg13g2_xnor2_1 _14662_ (.Y(_06523_),
    .A(\TRNG.sha256.expand.dout1[25] ),
    .B(\TRNG.sha256.expand.dout1[29] ));
 sg13g2_xnor2_1 _14663_ (.Y(_06524_),
    .A(\TRNG.sha256.expand.dout1[8] ),
    .B(_06523_));
 sg13g2_xor2_1 _14664_ (.B(\TRNG.sha256.expand.dout2[9] ),
    .A(\TRNG.sha256.expand.dout2[7] ),
    .X(_06525_));
 sg13g2_and2_1 _14665_ (.A(_06524_),
    .B(_06525_),
    .X(_06526_));
 sg13g2_xnor2_1 _14666_ (.Y(_06527_),
    .A(_06524_),
    .B(_06525_));
 sg13g2_o21ai_1 _14667_ (.B1(_06518_),
    .Y(_06528_),
    .A1(_06512_),
    .A2(_06519_));
 sg13g2_nor2_1 _14668_ (.A(_06522_),
    .B(_06528_),
    .Y(_06529_));
 sg13g2_nor2_1 _14669_ (.A(_06527_),
    .B(_06529_),
    .Y(_06530_));
 sg13g2_xor2_1 _14670_ (.B(_06529_),
    .A(_06527_),
    .X(_00252_));
 sg13g2_nor2_1 _14671_ (.A(_06526_),
    .B(_06530_),
    .Y(_06531_));
 sg13g2_xnor2_1 _14672_ (.Y(_06532_),
    .A(\TRNG.sha256.expand.dout1[26] ),
    .B(\TRNG.sha256.expand.dout1[30] ));
 sg13g2_xnor2_1 _14673_ (.Y(_06533_),
    .A(\TRNG.sha256.expand.dout1[9] ),
    .B(_06532_));
 sg13g2_xor2_1 _14674_ (.B(\TRNG.sha256.expand.dout2[8] ),
    .A(\TRNG.sha256.expand.dout2[10] ),
    .X(_06534_));
 sg13g2_and2_1 _14675_ (.A(_06533_),
    .B(_06534_),
    .X(_06535_));
 sg13g2_xor2_1 _14676_ (.B(_06534_),
    .A(_06533_),
    .X(_06536_));
 sg13g2_xnor2_1 _14677_ (.Y(_00253_),
    .A(_06531_),
    .B(_06536_));
 sg13g2_xnor2_1 _14678_ (.Y(_06537_),
    .A(\TRNG.sha256.expand.dout1[27] ),
    .B(\TRNG.sha256.expand.dout1[31] ));
 sg13g2_xnor2_1 _14679_ (.Y(_06538_),
    .A(\TRNG.sha256.expand.dout1[10] ),
    .B(_06537_));
 sg13g2_xor2_1 _14680_ (.B(\TRNG.sha256.expand.dout2[9] ),
    .A(\TRNG.sha256.expand.dout2[11] ),
    .X(_06539_));
 sg13g2_nand2_1 _14681_ (.Y(_06540_),
    .A(_06538_),
    .B(_06539_));
 sg13g2_xnor2_1 _14682_ (.Y(_06541_),
    .A(_06538_),
    .B(_06539_));
 sg13g2_nor2b_1 _14683_ (.A(_06527_),
    .B_N(_06536_),
    .Y(_06542_));
 sg13g2_o21ai_1 _14684_ (.B1(_06542_),
    .Y(_06543_),
    .A1(_06522_),
    .A2(_06528_));
 sg13g2_a21oi_1 _14685_ (.A1(_06526_),
    .A2(_06536_),
    .Y(_06544_),
    .B1(_06535_));
 sg13g2_a21o_1 _14686_ (.A2(_06544_),
    .A1(_06543_),
    .B1(_06541_),
    .X(_06545_));
 sg13g2_nand3_1 _14687_ (.B(_06543_),
    .C(_06544_),
    .A(_06541_),
    .Y(_06546_));
 sg13g2_and2_1 _14688_ (.A(_06545_),
    .B(_06546_),
    .X(_00254_));
 sg13g2_xnor2_1 _14689_ (.Y(_06547_),
    .A(\TRNG.sha256.expand.dout1[28] ),
    .B(\TRNG.sha256.expand.dout1[0] ));
 sg13g2_xnor2_1 _14690_ (.Y(_06548_),
    .A(\TRNG.sha256.expand.dout1[11] ),
    .B(_06547_));
 sg13g2_inv_1 _14691_ (.Y(_06549_),
    .A(_06548_));
 sg13g2_xnor2_1 _14692_ (.Y(_06550_),
    .A(\TRNG.sha256.expand.dout2[10] ),
    .B(\TRNG.sha256.expand.dout2[12] ));
 sg13g2_inv_1 _14693_ (.Y(_06551_),
    .A(_06550_));
 sg13g2_xnor2_1 _14694_ (.Y(_06552_),
    .A(_06548_),
    .B(_06551_));
 sg13g2_nand2_1 _14695_ (.Y(_06553_),
    .A(_06540_),
    .B(_06545_));
 sg13g2_xnor2_1 _14696_ (.Y(_00255_),
    .A(_06552_),
    .B(_06553_));
 sg13g2_a22oi_1 _14697_ (.Y(_06554_),
    .B1(_06548_),
    .B2(_06551_),
    .A2(_06539_),
    .A1(_06538_));
 sg13g2_a22oi_1 _14698_ (.Y(_06555_),
    .B1(_06554_),
    .B2(_06545_),
    .A2(_06550_),
    .A1(_06549_));
 sg13g2_xnor2_1 _14699_ (.Y(_06556_),
    .A(\TRNG.sha256.expand.dout1[29] ),
    .B(\TRNG.sha256.expand.dout1[1] ));
 sg13g2_xnor2_1 _14700_ (.Y(_06557_),
    .A(\TRNG.sha256.expand.dout1[12] ),
    .B(_06556_));
 sg13g2_xor2_1 _14701_ (.B(\TRNG.sha256.expand.dout2[13] ),
    .A(\TRNG.sha256.expand.dout2[11] ),
    .X(_06558_));
 sg13g2_and2_1 _14702_ (.A(_06557_),
    .B(_06558_),
    .X(_06559_));
 sg13g2_xor2_1 _14703_ (.B(_06558_),
    .A(_06557_),
    .X(_06560_));
 sg13g2_and2_1 _14704_ (.A(_06555_),
    .B(_06560_),
    .X(_06561_));
 sg13g2_xor2_1 _14705_ (.B(_06560_),
    .A(_06555_),
    .X(_00256_));
 sg13g2_xnor2_1 _14706_ (.Y(_06562_),
    .A(\TRNG.sha256.expand.dout1[30] ),
    .B(\TRNG.sha256.expand.dout1[2] ));
 sg13g2_xnor2_1 _14707_ (.Y(_06563_),
    .A(\TRNG.sha256.expand.dout1[13] ),
    .B(_06562_));
 sg13g2_xor2_1 _14708_ (.B(\TRNG.sha256.expand.dout2[14] ),
    .A(\TRNG.sha256.expand.dout2[12] ),
    .X(_06564_));
 sg13g2_nand2_1 _14709_ (.Y(_06565_),
    .A(_06563_),
    .B(_06564_));
 sg13g2_xor2_1 _14710_ (.B(_06564_),
    .A(_06563_),
    .X(_06566_));
 sg13g2_o21ai_1 _14711_ (.B1(_06566_),
    .Y(_06567_),
    .A1(_06559_),
    .A2(_06561_));
 sg13g2_or3_1 _14712_ (.A(_06559_),
    .B(_06561_),
    .C(_06566_),
    .X(_06568_));
 sg13g2_and2_1 _14713_ (.A(_06567_),
    .B(_06568_),
    .X(_00257_));
 sg13g2_nand2_1 _14714_ (.Y(_06569_),
    .A(_06565_),
    .B(_06567_));
 sg13g2_xnor2_1 _14715_ (.Y(_06570_),
    .A(\TRNG.sha256.expand.dout1[14] ),
    .B(\TRNG.sha256.expand.dout1[31] ));
 sg13g2_xnor2_1 _14716_ (.Y(_06571_),
    .A(\TRNG.sha256.expand.dout1[3] ),
    .B(_06570_));
 sg13g2_xor2_1 _14717_ (.B(\TRNG.sha256.expand.dout2[15] ),
    .A(\TRNG.sha256.expand.dout2[13] ),
    .X(_06572_));
 sg13g2_and2_1 _14718_ (.A(_06571_),
    .B(_06572_),
    .X(_06573_));
 sg13g2_xor2_1 _14719_ (.B(_06572_),
    .A(_06571_),
    .X(_06574_));
 sg13g2_xor2_1 _14720_ (.B(_06574_),
    .A(_06569_),
    .X(_00258_));
 sg13g2_xor2_1 _14721_ (.B(\TRNG.sha256.expand.dout2[16] ),
    .A(\TRNG.sha256.expand.dout2[14] ),
    .X(_06575_));
 sg13g2_xor2_1 _14722_ (.B(\TRNG.sha256.expand.dout1[15] ),
    .A(\TRNG.sha256.expand.dout1[4] ),
    .X(_06576_));
 sg13g2_nand2_1 _14723_ (.Y(_06577_),
    .A(_06575_),
    .B(_06576_));
 sg13g2_xnor2_1 _14724_ (.Y(_06578_),
    .A(_06575_),
    .B(_06576_));
 sg13g2_a21oi_1 _14725_ (.A1(_06569_),
    .A2(_06574_),
    .Y(_06579_),
    .B1(_06573_));
 sg13g2_xor2_1 _14726_ (.B(_06579_),
    .A(_06578_),
    .X(_00259_));
 sg13g2_xor2_1 _14727_ (.B(\TRNG.sha256.expand.dout2[15] ),
    .A(\TRNG.sha256.expand.dout2[17] ),
    .X(_06580_));
 sg13g2_xor2_1 _14728_ (.B(\TRNG.sha256.expand.dout1[16] ),
    .A(\TRNG.sha256.expand.dout1[5] ),
    .X(_06581_));
 sg13g2_and2_1 _14729_ (.A(_06580_),
    .B(_06581_),
    .X(_06582_));
 sg13g2_xnor2_1 _14730_ (.Y(_06583_),
    .A(_06580_),
    .B(_06581_));
 sg13g2_inv_1 _14731_ (.Y(_06584_),
    .A(_06583_));
 sg13g2_o21ai_1 _14732_ (.B1(_06577_),
    .Y(_06585_),
    .A1(_06578_),
    .A2(_06579_));
 sg13g2_xnor2_1 _14733_ (.Y(_00261_),
    .A(_06583_),
    .B(_06585_));
 sg13g2_a21oi_1 _14734_ (.A1(_06584_),
    .A2(_06585_),
    .Y(_06586_),
    .B1(_06582_));
 sg13g2_xnor2_1 _14735_ (.Y(_06587_),
    .A(\TRNG.sha256.expand.dout2[18] ),
    .B(\TRNG.sha256.expand.dout1[6] ));
 sg13g2_xor2_1 _14736_ (.B(\TRNG.sha256.expand.dout1[17] ),
    .A(\TRNG.sha256.expand.dout2[16] ),
    .X(_06588_));
 sg13g2_xnor2_1 _14737_ (.Y(_06589_),
    .A(_06587_),
    .B(_06588_));
 sg13g2_xnor2_1 _14738_ (.Y(_00262_),
    .A(_06586_),
    .B(_06589_));
 sg13g2_nand2_1 _14739_ (.Y(_06590_),
    .A(\TRNG.sha256.expand.dout1[0] ),
    .B(net3790));
 sg13g2_xor2_1 _14740_ (.B(\TRNG.sha256.expand.sm0.sum_0[0] ),
    .A(\TRNG.sha256.expand.dout1[0] ),
    .X(_06591_));
 sg13g2_nand2_1 _14741_ (.Y(_06592_),
    .A(\TRNG.sha256.expand.dout2[0] ),
    .B(_06591_));
 sg13g2_xor2_1 _14742_ (.B(_06591_),
    .A(net3484),
    .X(_00276_));
 sg13g2_and2_1 _14743_ (.A(\TRNG.sha256.expand.dout1[1] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[1] ),
    .X(_06593_));
 sg13g2_xor2_1 _14744_ (.B(\TRNG.sha256.expand.sm0.sum_0[1] ),
    .A(\TRNG.sha256.expand.dout1[1] ),
    .X(_06594_));
 sg13g2_xnor2_1 _14745_ (.Y(_06595_),
    .A(\TRNG.sha256.expand.dout2[1] ),
    .B(_06594_));
 sg13g2_a21oi_2 _14746_ (.B1(_06595_),
    .Y(_06596_),
    .A2(_06592_),
    .A1(_06590_));
 sg13g2_nand3_1 _14747_ (.B(_06592_),
    .C(_06595_),
    .A(_06590_),
    .Y(_06597_));
 sg13g2_nor2b_1 _14748_ (.A(_06596_),
    .B_N(net3791),
    .Y(_00277_));
 sg13g2_a21oi_1 _14749_ (.A1(\TRNG.sha256.expand.dout2[1] ),
    .A2(_06594_),
    .Y(_06598_),
    .B1(_06593_));
 sg13g2_and2_1 _14750_ (.A(\TRNG.sha256.expand.dout1[2] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[2] ),
    .X(_06599_));
 sg13g2_xor2_1 _14751_ (.B(\TRNG.sha256.expand.sm0.sum_0[2] ),
    .A(\TRNG.sha256.expand.dout1[2] ),
    .X(_06600_));
 sg13g2_xnor2_1 _14752_ (.Y(_06601_),
    .A(\TRNG.sha256.expand.dout2[2] ),
    .B(_06600_));
 sg13g2_nor2_1 _14753_ (.A(_06598_),
    .B(_06601_),
    .Y(_06602_));
 sg13g2_xor2_1 _14754_ (.B(_06601_),
    .A(_06598_),
    .X(_06603_));
 sg13g2_xor2_1 _14755_ (.B(_06603_),
    .A(_06596_),
    .X(_00298_));
 sg13g2_a21oi_2 _14756_ (.B1(_06602_),
    .Y(_06604_),
    .A2(_06603_),
    .A1(_06596_));
 sg13g2_a21oi_1 _14757_ (.A1(\TRNG.sha256.expand.dout2[2] ),
    .A2(_06600_),
    .Y(_06605_),
    .B1(_06599_));
 sg13g2_and2_1 _14758_ (.A(\TRNG.sha256.expand.dout1[3] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[3] ),
    .X(_06606_));
 sg13g2_xor2_1 _14759_ (.B(\TRNG.sha256.expand.sm0.sum_0[3] ),
    .A(\TRNG.sha256.expand.dout1[3] ),
    .X(_06607_));
 sg13g2_xnor2_1 _14760_ (.Y(_06608_),
    .A(\TRNG.sha256.expand.dout2[3] ),
    .B(_06607_));
 sg13g2_or2_1 _14761_ (.X(_06609_),
    .B(_06608_),
    .A(_06605_));
 sg13g2_xnor2_1 _14762_ (.Y(_06610_),
    .A(_06605_),
    .B(_06608_));
 sg13g2_xor2_1 _14763_ (.B(_06610_),
    .A(_06604_),
    .X(_00301_));
 sg13g2_o21ai_1 _14764_ (.B1(_06609_),
    .Y(_06611_),
    .A1(_06604_),
    .A2(_06610_));
 sg13g2_a21oi_2 _14765_ (.B1(_06606_),
    .Y(_06612_),
    .A2(_06607_),
    .A1(\TRNG.sha256.expand.dout2[3] ));
 sg13g2_nand2_1 _14766_ (.Y(_06613_),
    .A(\TRNG.sha256.expand.dout1[4] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[4] ));
 sg13g2_xor2_1 _14767_ (.B(\TRNG.sha256.expand.sm0.sum_0[4] ),
    .A(\TRNG.sha256.expand.dout1[4] ),
    .X(_06614_));
 sg13g2_nand2_1 _14768_ (.Y(_06615_),
    .A(\TRNG.sha256.expand.dout2[4] ),
    .B(_06614_));
 sg13g2_xnor2_1 _14769_ (.Y(_06616_),
    .A(\TRNG.sha256.expand.dout2[4] ),
    .B(_06614_));
 sg13g2_nor2_1 _14770_ (.A(_06612_),
    .B(_06616_),
    .Y(_06617_));
 sg13g2_xor2_1 _14771_ (.B(_06616_),
    .A(_06612_),
    .X(_06618_));
 sg13g2_xor2_1 _14772_ (.B(_06618_),
    .A(_06611_),
    .X(_00302_));
 sg13g2_a21oi_1 _14773_ (.A1(_06611_),
    .A2(_06618_),
    .Y(_06619_),
    .B1(_06617_));
 sg13g2_nand2_1 _14774_ (.Y(_06620_),
    .A(_06613_),
    .B(_06615_));
 sg13g2_and2_1 _14775_ (.A(\TRNG.sha256.expand.dout1[5] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[5] ),
    .X(_06621_));
 sg13g2_xor2_1 _14776_ (.B(\TRNG.sha256.expand.sm0.sum_0[5] ),
    .A(\TRNG.sha256.expand.dout1[5] ),
    .X(_06622_));
 sg13g2_xnor2_1 _14777_ (.Y(_06623_),
    .A(\TRNG.sha256.expand.dout2[5] ),
    .B(_06622_));
 sg13g2_inv_1 _14778_ (.Y(_06624_),
    .A(_06623_));
 sg13g2_nand3_1 _14779_ (.B(_06615_),
    .C(_06623_),
    .A(_06613_),
    .Y(_06625_));
 sg13g2_inv_1 _14780_ (.Y(_06626_),
    .A(_06625_));
 sg13g2_xnor2_1 _14781_ (.Y(_06627_),
    .A(_06620_),
    .B(_06623_));
 sg13g2_xnor2_1 _14782_ (.Y(_00303_),
    .A(_06619_),
    .B(_06627_));
 sg13g2_a21oi_1 _14783_ (.A1(\TRNG.sha256.expand.dout2[5] ),
    .A2(_06622_),
    .Y(_06628_),
    .B1(_06621_));
 sg13g2_and2_1 _14784_ (.A(\TRNG.sha256.expand.dout1[6] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[6] ),
    .X(_06629_));
 sg13g2_xor2_1 _14785_ (.B(\TRNG.sha256.expand.sm0.sum_0[6] ),
    .A(\TRNG.sha256.expand.dout1[6] ),
    .X(_06630_));
 sg13g2_xnor2_1 _14786_ (.Y(_06631_),
    .A(\TRNG.sha256.expand.dout2[6] ),
    .B(_06630_));
 sg13g2_or2_1 _14787_ (.X(_06632_),
    .B(_06631_),
    .A(_06628_));
 sg13g2_xnor2_1 _14788_ (.Y(_06633_),
    .A(_06628_),
    .B(_06631_));
 sg13g2_a221oi_1 _14789_ (.B2(_06624_),
    .C1(_06617_),
    .B1(_06620_),
    .A1(_06611_),
    .Y(_06634_),
    .A2(_06618_));
 sg13g2_or3_1 _14790_ (.A(_06626_),
    .B(_06633_),
    .C(_06634_),
    .X(_06635_));
 sg13g2_o21ai_1 _14791_ (.B1(_06633_),
    .Y(_06636_),
    .A1(_06626_),
    .A2(_06634_));
 sg13g2_and2_1 _14792_ (.A(_06635_),
    .B(_06636_),
    .X(_00304_));
 sg13g2_a21oi_1 _14793_ (.A1(\TRNG.sha256.expand.dout2[6] ),
    .A2(_06630_),
    .Y(_06637_),
    .B1(_06629_));
 sg13g2_and2_1 _14794_ (.A(\TRNG.sha256.expand.dout1[7] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[7] ),
    .X(_06638_));
 sg13g2_xor2_1 _14795_ (.B(\TRNG.sha256.expand.sm0.sum_0[7] ),
    .A(\TRNG.sha256.expand.dout1[7] ),
    .X(_06639_));
 sg13g2_xnor2_1 _14796_ (.Y(_06640_),
    .A(\TRNG.sha256.expand.dout2[7] ),
    .B(_06639_));
 sg13g2_nor2_1 _14797_ (.A(_06637_),
    .B(_06640_),
    .Y(_06641_));
 sg13g2_xor2_1 _14798_ (.B(_06640_),
    .A(_06637_),
    .X(_06642_));
 sg13g2_inv_1 _14799_ (.Y(_06643_),
    .A(_06642_));
 sg13g2_a21oi_2 _14800_ (.B1(_06643_),
    .Y(_06644_),
    .A2(_06635_),
    .A1(_06632_));
 sg13g2_nand3_1 _14801_ (.B(_06635_),
    .C(_06643_),
    .A(_06632_),
    .Y(_06645_));
 sg13g2_nor2b_2 _14802_ (.A(_06644_),
    .B_N(_06645_),
    .Y(_00305_));
 sg13g2_nor2_1 _14803_ (.A(_06641_),
    .B(_06644_),
    .Y(_06646_));
 sg13g2_a21oi_1 _14804_ (.A1(\TRNG.sha256.expand.dout2[7] ),
    .A2(_06639_),
    .Y(_06647_),
    .B1(_06638_));
 sg13g2_nand2_1 _14805_ (.Y(_06648_),
    .A(\TRNG.sha256.expand.dout1[8] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[8] ));
 sg13g2_xor2_1 _14806_ (.B(\TRNG.sha256.expand.sm0.sum_0[8] ),
    .A(\TRNG.sha256.expand.dout1[8] ),
    .X(_06649_));
 sg13g2_nand2_1 _14807_ (.Y(_06650_),
    .A(\TRNG.sha256.expand.dout2[8] ),
    .B(_06649_));
 sg13g2_xnor2_1 _14808_ (.Y(_06651_),
    .A(\TRNG.sha256.expand.dout2[8] ),
    .B(_06649_));
 sg13g2_nor2_1 _14809_ (.A(_06647_),
    .B(_06651_),
    .Y(_06652_));
 sg13g2_inv_1 _14810_ (.Y(_06653_),
    .A(_06652_));
 sg13g2_xor2_1 _14811_ (.B(_06651_),
    .A(_06647_),
    .X(_06654_));
 sg13g2_o21ai_1 _14812_ (.B1(_06654_),
    .Y(_06655_),
    .A1(_06641_),
    .A2(_06644_));
 sg13g2_xnor2_1 _14813_ (.Y(_00306_),
    .A(_06646_),
    .B(_06654_));
 sg13g2_nand2_1 _14814_ (.Y(_06656_),
    .A(_06653_),
    .B(_06655_));
 sg13g2_and2_1 _14815_ (.A(\TRNG.sha256.expand.dout1[9] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[9] ),
    .X(_06657_));
 sg13g2_xor2_1 _14816_ (.B(\TRNG.sha256.expand.sm0.sum_0[9] ),
    .A(\TRNG.sha256.expand.dout1[9] ),
    .X(_06658_));
 sg13g2_xnor2_1 _14817_ (.Y(_06659_),
    .A(\TRNG.sha256.expand.dout2[9] ),
    .B(_06658_));
 sg13g2_a21oi_2 _14818_ (.B1(_06659_),
    .Y(_06660_),
    .A2(_06650_),
    .A1(_06648_));
 sg13g2_nand3_1 _14819_ (.B(_06650_),
    .C(_06659_),
    .A(_06648_),
    .Y(_06661_));
 sg13g2_inv_1 _14820_ (.Y(_06662_),
    .A(_06661_));
 sg13g2_nor2_1 _14821_ (.A(_06660_),
    .B(_06662_),
    .Y(_06663_));
 sg13g2_xor2_1 _14822_ (.B(_06663_),
    .A(_06656_),
    .X(_00307_));
 sg13g2_a21oi_1 _14823_ (.A1(\TRNG.sha256.expand.dout2[9] ),
    .A2(_06658_),
    .Y(_06664_),
    .B1(_06657_));
 sg13g2_nand2_1 _14824_ (.Y(_06665_),
    .A(\TRNG.sha256.expand.dout1[10] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[10] ));
 sg13g2_xor2_1 _14825_ (.B(\TRNG.sha256.expand.sm0.sum_0[10] ),
    .A(\TRNG.sha256.expand.dout1[10] ),
    .X(_06666_));
 sg13g2_nand2_1 _14826_ (.Y(_06667_),
    .A(\TRNG.sha256.expand.dout2[10] ),
    .B(_06666_));
 sg13g2_xnor2_1 _14827_ (.Y(_06668_),
    .A(\TRNG.sha256.expand.dout2[10] ),
    .B(_06666_));
 sg13g2_nor2_1 _14828_ (.A(_06664_),
    .B(_06668_),
    .Y(_06669_));
 sg13g2_inv_1 _14829_ (.Y(_06670_),
    .A(_06669_));
 sg13g2_xor2_1 _14830_ (.B(_06668_),
    .A(_06664_),
    .X(_06671_));
 sg13g2_a21oi_1 _14831_ (.A1(_06653_),
    .A2(_06655_),
    .Y(_06672_),
    .B1(_06662_));
 sg13g2_o21ai_1 _14832_ (.B1(_06671_),
    .Y(_06673_),
    .A1(_06660_),
    .A2(_06672_));
 sg13g2_or3_1 _14833_ (.A(_06660_),
    .B(_06671_),
    .C(_06672_),
    .X(_06674_));
 sg13g2_and2_1 _14834_ (.A(_06673_),
    .B(_06674_),
    .X(_00278_));
 sg13g2_nand2_1 _14835_ (.Y(_06675_),
    .A(_06670_),
    .B(_06673_));
 sg13g2_and2_1 _14836_ (.A(\TRNG.sha256.expand.dout1[11] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[11] ),
    .X(_06676_));
 sg13g2_xor2_1 _14837_ (.B(\TRNG.sha256.expand.sm0.sum_0[11] ),
    .A(\TRNG.sha256.expand.dout1[11] ),
    .X(_06677_));
 sg13g2_xnor2_1 _14838_ (.Y(_06678_),
    .A(\TRNG.sha256.expand.dout2[11] ),
    .B(_06677_));
 sg13g2_a21oi_2 _14839_ (.B1(_06678_),
    .Y(_06679_),
    .A2(_06667_),
    .A1(_06665_));
 sg13g2_nand3_1 _14840_ (.B(_06667_),
    .C(_06678_),
    .A(_06665_),
    .Y(_06680_));
 sg13g2_inv_1 _14841_ (.Y(_06681_),
    .A(_06680_));
 sg13g2_nor2_1 _14842_ (.A(_06679_),
    .B(_06681_),
    .Y(_06682_));
 sg13g2_xor2_1 _14843_ (.B(_06682_),
    .A(_06675_),
    .X(_00279_));
 sg13g2_a21oi_2 _14844_ (.B1(_06676_),
    .Y(_06683_),
    .A2(_06677_),
    .A1(\TRNG.sha256.expand.dout2[11] ));
 sg13g2_nand2_1 _14845_ (.Y(_06684_),
    .A(\TRNG.sha256.expand.dout1[12] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[12] ));
 sg13g2_xor2_1 _14846_ (.B(\TRNG.sha256.expand.sm0.sum_0[12] ),
    .A(\TRNG.sha256.expand.dout1[12] ),
    .X(_06685_));
 sg13g2_nand2_1 _14847_ (.Y(_06686_),
    .A(\TRNG.sha256.expand.dout2[12] ),
    .B(_06685_));
 sg13g2_xnor2_1 _14848_ (.Y(_06687_),
    .A(\TRNG.sha256.expand.dout2[12] ),
    .B(_06685_));
 sg13g2_nor2_1 _14849_ (.A(_06683_),
    .B(_06687_),
    .Y(_06688_));
 sg13g2_inv_1 _14850_ (.Y(_06689_),
    .A(_06688_));
 sg13g2_xor2_1 _14851_ (.B(_06687_),
    .A(_06683_),
    .X(_06690_));
 sg13g2_a21oi_2 _14852_ (.B1(_06681_),
    .Y(_06691_),
    .A2(_06673_),
    .A1(_06670_));
 sg13g2_or2_1 _14853_ (.X(_06692_),
    .B(_06691_),
    .A(_06679_));
 sg13g2_o21ai_1 _14854_ (.B1(_06690_),
    .Y(_06693_),
    .A1(_06679_),
    .A2(_06691_));
 sg13g2_xor2_1 _14855_ (.B(_06692_),
    .A(_06690_),
    .X(_00280_));
 sg13g2_and2_1 _14856_ (.A(_06689_),
    .B(_06693_),
    .X(_06694_));
 sg13g2_and2_1 _14857_ (.A(\TRNG.sha256.expand.dout1[13] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[13] ),
    .X(_06695_));
 sg13g2_xor2_1 _14858_ (.B(\TRNG.sha256.expand.sm0.sum_0[13] ),
    .A(\TRNG.sha256.expand.dout1[13] ),
    .X(_06696_));
 sg13g2_xnor2_1 _14859_ (.Y(_06697_),
    .A(\TRNG.sha256.expand.dout2[13] ),
    .B(_06696_));
 sg13g2_a21oi_1 _14860_ (.A1(_06684_),
    .A2(_06686_),
    .Y(_06698_),
    .B1(_06697_));
 sg13g2_nand3_1 _14861_ (.B(_06686_),
    .C(_06697_),
    .A(_06684_),
    .Y(_06699_));
 sg13g2_inv_1 _14862_ (.Y(_06700_),
    .A(_06699_));
 sg13g2_nor2_1 _14863_ (.A(_06698_),
    .B(_06700_),
    .Y(_06701_));
 sg13g2_xnor2_1 _14864_ (.Y(_00281_),
    .A(_06694_),
    .B(_06701_));
 sg13g2_a21oi_1 _14865_ (.A1(\TRNG.sha256.expand.dout2[13] ),
    .A2(_06696_),
    .Y(_06702_),
    .B1(_06695_));
 sg13g2_nand2_1 _14866_ (.Y(_06703_),
    .A(\TRNG.sha256.expand.dout1[14] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[14] ));
 sg13g2_xor2_1 _14867_ (.B(\TRNG.sha256.expand.sm0.sum_0[14] ),
    .A(\TRNG.sha256.expand.dout1[14] ),
    .X(_06704_));
 sg13g2_nand2_1 _14868_ (.Y(_06705_),
    .A(\TRNG.sha256.expand.dout2[14] ),
    .B(_06704_));
 sg13g2_xnor2_1 _14869_ (.Y(_06706_),
    .A(\TRNG.sha256.expand.dout2[14] ),
    .B(_06704_));
 sg13g2_nor2_1 _14870_ (.A(_06702_),
    .B(_06706_),
    .Y(_06707_));
 sg13g2_xor2_1 _14871_ (.B(_06706_),
    .A(_06702_),
    .X(_06708_));
 sg13g2_a21oi_1 _14872_ (.A1(_06689_),
    .A2(_06693_),
    .Y(_06709_),
    .B1(_06700_));
 sg13g2_or2_1 _14873_ (.X(_06710_),
    .B(_06709_),
    .A(_06698_));
 sg13g2_o21ai_1 _14874_ (.B1(_06708_),
    .Y(_06711_),
    .A1(_06698_),
    .A2(_06709_));
 sg13g2_xor2_1 _14875_ (.B(_06710_),
    .A(_06708_),
    .X(_00282_));
 sg13g2_nor2b_1 _14876_ (.A(_06707_),
    .B_N(_06711_),
    .Y(_06712_));
 sg13g2_and2_1 _14877_ (.A(\TRNG.sha256.expand.dout1[15] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[15] ),
    .X(_06713_));
 sg13g2_xor2_1 _14878_ (.B(\TRNG.sha256.expand.sm0.sum_0[15] ),
    .A(\TRNG.sha256.expand.dout1[15] ),
    .X(_06714_));
 sg13g2_xnor2_1 _14879_ (.Y(_06715_),
    .A(\TRNG.sha256.expand.dout2[15] ),
    .B(_06714_));
 sg13g2_a21o_1 _14880_ (.A2(_06705_),
    .A1(_06703_),
    .B1(_06715_),
    .X(_06716_));
 sg13g2_nand3_1 _14881_ (.B(_06705_),
    .C(_06715_),
    .A(_06703_),
    .Y(_06717_));
 sg13g2_and2_1 _14882_ (.A(_06716_),
    .B(_06717_),
    .X(_06718_));
 sg13g2_xnor2_1 _14883_ (.Y(_00283_),
    .A(_06712_),
    .B(_06718_));
 sg13g2_nand2_1 _14884_ (.Y(_06719_),
    .A(\TRNG.sha256.expand.dout1[16] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[16] ));
 sg13g2_xor2_1 _14885_ (.B(\TRNG.sha256.expand.sm0.sum_0[16] ),
    .A(\TRNG.sha256.expand.dout1[16] ),
    .X(_06720_));
 sg13g2_nand2_1 _14886_ (.Y(_06721_),
    .A(\TRNG.sha256.expand.dout2[16] ),
    .B(_06720_));
 sg13g2_xnor2_1 _14887_ (.Y(_06722_),
    .A(\TRNG.sha256.expand.dout2[16] ),
    .B(_06720_));
 sg13g2_a21oi_1 _14888_ (.A1(\TRNG.sha256.expand.dout2[15] ),
    .A2(_06714_),
    .Y(_06723_),
    .B1(_06713_));
 sg13g2_nor2_1 _14889_ (.A(_06722_),
    .B(_06723_),
    .Y(_06724_));
 sg13g2_xnor2_1 _14890_ (.Y(_06725_),
    .A(_06722_),
    .B(_06723_));
 sg13g2_inv_1 _14891_ (.Y(_06726_),
    .A(_06725_));
 sg13g2_nand3b_1 _14892_ (.B(_06711_),
    .C(_06716_),
    .Y(_06727_),
    .A_N(_06707_));
 sg13g2_and2_1 _14893_ (.A(_06717_),
    .B(_06727_),
    .X(_06728_));
 sg13g2_xnor2_1 _14894_ (.Y(_00284_),
    .A(_06725_),
    .B(_06728_));
 sg13g2_nand2_1 _14895_ (.Y(_06729_),
    .A(\TRNG.sha256.expand.dout1[17] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[17] ));
 sg13g2_xor2_1 _14896_ (.B(\TRNG.sha256.expand.sm0.sum_0[17] ),
    .A(\TRNG.sha256.expand.dout1[17] ),
    .X(_06730_));
 sg13g2_nand2_1 _14897_ (.Y(_06731_),
    .A(\TRNG.sha256.expand.dout2[17] ),
    .B(_06730_));
 sg13g2_xnor2_1 _14898_ (.Y(_06732_),
    .A(\TRNG.sha256.expand.dout2[17] ),
    .B(_06730_));
 sg13g2_a21oi_1 _14899_ (.A1(_06719_),
    .A2(_06721_),
    .Y(_06733_),
    .B1(_06732_));
 sg13g2_nand3_1 _14900_ (.B(_06721_),
    .C(_06732_),
    .A(_06719_),
    .Y(_06734_));
 sg13g2_nor2b_1 _14901_ (.A(_06733_),
    .B_N(_06734_),
    .Y(_06735_));
 sg13g2_a21oi_1 _14902_ (.A1(_06726_),
    .A2(_06728_),
    .Y(_06736_),
    .B1(_06724_));
 sg13g2_xnor2_1 _14903_ (.Y(_00285_),
    .A(_06735_),
    .B(_06736_));
 sg13g2_nand2_1 _14904_ (.Y(_06737_),
    .A(\TRNG.sha256.expand.dout1[18] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[18] ));
 sg13g2_xor2_1 _14905_ (.B(\TRNG.sha256.expand.sm0.sum_0[18] ),
    .A(\TRNG.sha256.expand.dout1[18] ),
    .X(_06738_));
 sg13g2_nand2_1 _14906_ (.Y(_06739_),
    .A(\TRNG.sha256.expand.dout2[18] ),
    .B(_06738_));
 sg13g2_xnor2_1 _14907_ (.Y(_06740_),
    .A(\TRNG.sha256.expand.dout2[18] ),
    .B(_06738_));
 sg13g2_a21oi_2 _14908_ (.B1(_06740_),
    .Y(_06741_),
    .A2(_06731_),
    .A1(_06729_));
 sg13g2_nand3_1 _14909_ (.B(_06731_),
    .C(_06740_),
    .A(_06729_),
    .Y(_06742_));
 sg13g2_nand2b_1 _14910_ (.Y(_06743_),
    .B(_06742_),
    .A_N(_06741_));
 sg13g2_nand2_1 _14911_ (.Y(_06744_),
    .A(_06724_),
    .B(_06734_));
 sg13g2_nand4_1 _14912_ (.B(_06726_),
    .C(_06727_),
    .A(_06717_),
    .Y(_06745_),
    .D(_06735_));
 sg13g2_nand3b_1 _14913_ (.B(_06744_),
    .C(_06745_),
    .Y(_06746_),
    .A_N(_06733_));
 sg13g2_nand2b_1 _14914_ (.Y(_06747_),
    .B(_06746_),
    .A_N(_06743_));
 sg13g2_xnor2_1 _14915_ (.Y(_00286_),
    .A(_06743_),
    .B(_06746_));
 sg13g2_and2_1 _14916_ (.A(\TRNG.sha256.expand.dout1[19] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[19] ),
    .X(_06748_));
 sg13g2_xor2_1 _14917_ (.B(\TRNG.sha256.expand.sm0.sum_0[19] ),
    .A(\TRNG.sha256.expand.dout1[19] ),
    .X(_06749_));
 sg13g2_xnor2_1 _14918_ (.Y(_06750_),
    .A(\TRNG.sha256.expand.dout2[19] ),
    .B(_06749_));
 sg13g2_a21oi_2 _14919_ (.B1(_06750_),
    .Y(_06751_),
    .A2(_06739_),
    .A1(_06737_));
 sg13g2_nand3_1 _14920_ (.B(_06739_),
    .C(_06750_),
    .A(_06737_),
    .Y(_06752_));
 sg13g2_inv_1 _14921_ (.Y(_06753_),
    .A(_06752_));
 sg13g2_nor2_1 _14922_ (.A(_06751_),
    .B(_06753_),
    .Y(_06754_));
 sg13g2_a21oi_1 _14923_ (.A1(_06742_),
    .A2(_06746_),
    .Y(_06755_),
    .B1(_06741_));
 sg13g2_xnor2_1 _14924_ (.Y(_00287_),
    .A(_06754_),
    .B(_06755_));
 sg13g2_nand2_1 _14925_ (.Y(_06756_),
    .A(\TRNG.sha256.expand.dout1[20] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[20] ));
 sg13g2_xor2_1 _14926_ (.B(\TRNG.sha256.expand.sm0.sum_0[20] ),
    .A(\TRNG.sha256.expand.dout1[20] ),
    .X(_06757_));
 sg13g2_nand2_1 _14927_ (.Y(_06758_),
    .A(\TRNG.sha256.expand.dout2[20] ),
    .B(_06757_));
 sg13g2_xnor2_1 _14928_ (.Y(_06759_),
    .A(\TRNG.sha256.expand.dout2[20] ),
    .B(_06757_));
 sg13g2_a21oi_1 _14929_ (.A1(\TRNG.sha256.expand.dout2[19] ),
    .A2(_06749_),
    .Y(_06760_),
    .B1(_06748_));
 sg13g2_nor2_1 _14930_ (.A(_06759_),
    .B(_06760_),
    .Y(_06761_));
 sg13g2_xnor2_1 _14931_ (.Y(_06762_),
    .A(_06759_),
    .B(_06760_));
 sg13g2_inv_1 _14932_ (.Y(_06763_),
    .A(_06762_));
 sg13g2_nor2_1 _14933_ (.A(_06741_),
    .B(_06751_),
    .Y(_06764_));
 sg13g2_nor3_1 _14934_ (.A(_06743_),
    .B(_06751_),
    .C(_06753_),
    .Y(_06765_));
 sg13g2_a21oi_1 _14935_ (.A1(_06747_),
    .A2(_06764_),
    .Y(_06766_),
    .B1(_06753_));
 sg13g2_a221oi_1 _14936_ (.B2(_06746_),
    .C1(_06751_),
    .B1(_06765_),
    .A1(_06741_),
    .Y(_06767_),
    .A2(_06752_));
 sg13g2_xnor2_1 _14937_ (.Y(_00288_),
    .A(_06763_),
    .B(_06767_));
 sg13g2_nand2_1 _14938_ (.Y(_06768_),
    .A(\TRNG.sha256.expand.dout1[21] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[21] ));
 sg13g2_xor2_1 _14939_ (.B(\TRNG.sha256.expand.sm0.sum_0[21] ),
    .A(\TRNG.sha256.expand.dout1[21] ),
    .X(_06769_));
 sg13g2_nand2_1 _14940_ (.Y(_06770_),
    .A(\TRNG.sha256.expand.dout2[21] ),
    .B(_06769_));
 sg13g2_xnor2_1 _14941_ (.Y(_06771_),
    .A(\TRNG.sha256.expand.dout2[21] ),
    .B(_06769_));
 sg13g2_nand3_1 _14942_ (.B(_06758_),
    .C(_06771_),
    .A(_06756_),
    .Y(_06772_));
 sg13g2_inv_1 _14943_ (.Y(_06773_),
    .A(_06772_));
 sg13g2_a21oi_1 _14944_ (.A1(_06756_),
    .A2(_06758_),
    .Y(_06774_),
    .B1(_06771_));
 sg13g2_nor2_1 _14945_ (.A(_06773_),
    .B(_06774_),
    .Y(_06775_));
 sg13g2_a21oi_1 _14946_ (.A1(_06763_),
    .A2(_06766_),
    .Y(_06776_),
    .B1(_06761_));
 sg13g2_xnor2_1 _14947_ (.Y(_00289_),
    .A(_06775_),
    .B(_06776_));
 sg13g2_nand2_1 _14948_ (.Y(_06777_),
    .A(\TRNG.sha256.expand.dout1[22] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[22] ));
 sg13g2_xor2_1 _14949_ (.B(\TRNG.sha256.expand.sm0.sum_0[22] ),
    .A(\TRNG.sha256.expand.dout1[22] ),
    .X(_06778_));
 sg13g2_nand2_1 _14950_ (.Y(_06779_),
    .A(\TRNG.sha256.expand.dout2[22] ),
    .B(_06778_));
 sg13g2_xnor2_1 _14951_ (.Y(_06780_),
    .A(\TRNG.sha256.expand.dout2[22] ),
    .B(_06778_));
 sg13g2_a21oi_1 _14952_ (.A1(_06768_),
    .A2(_06770_),
    .Y(_06781_),
    .B1(_06780_));
 sg13g2_nand3_1 _14953_ (.B(_06770_),
    .C(_06780_),
    .A(_06768_),
    .Y(_06782_));
 sg13g2_nor2b_1 _14954_ (.A(_06781_),
    .B_N(_06782_),
    .Y(_06783_));
 sg13g2_nor4_1 _14955_ (.A(_06762_),
    .B(_06767_),
    .C(_06773_),
    .D(_06774_),
    .Y(_06784_));
 sg13g2_a21oi_1 _14956_ (.A1(_06761_),
    .A2(_06772_),
    .Y(_06785_),
    .B1(_06774_));
 sg13g2_nor2b_1 _14957_ (.A(_06784_),
    .B_N(_06785_),
    .Y(_06786_));
 sg13g2_nor2b_1 _14958_ (.A(_06786_),
    .B_N(_06783_),
    .Y(_06787_));
 sg13g2_xnor2_1 _14959_ (.Y(_00290_),
    .A(_06783_),
    .B(_06786_));
 sg13g2_and2_1 _14960_ (.A(\TRNG.sha256.expand.dout1[23] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[23] ),
    .X(_06788_));
 sg13g2_xor2_1 _14961_ (.B(\TRNG.sha256.expand.sm0.sum_0[23] ),
    .A(\TRNG.sha256.expand.dout1[23] ),
    .X(_06789_));
 sg13g2_xnor2_1 _14962_ (.Y(_06790_),
    .A(\TRNG.sha256.expand.dout2[23] ),
    .B(_06789_));
 sg13g2_and3_1 _14963_ (.X(_06791_),
    .A(_06777_),
    .B(_06779_),
    .C(_06790_));
 sg13g2_a21oi_1 _14964_ (.A1(_06777_),
    .A2(_06779_),
    .Y(_06792_),
    .B1(_06790_));
 sg13g2_nor2_1 _14965_ (.A(_06791_),
    .B(_06792_),
    .Y(_06793_));
 sg13g2_nor2_1 _14966_ (.A(_06781_),
    .B(_06787_),
    .Y(_06794_));
 sg13g2_xnor2_1 _14967_ (.Y(_00291_),
    .A(_06793_),
    .B(_06794_));
 sg13g2_nor2_1 _14968_ (.A(_06781_),
    .B(_06792_),
    .Y(_06795_));
 sg13g2_o21ai_1 _14969_ (.B1(_06785_),
    .Y(_06796_),
    .A1(_06791_),
    .A2(_06795_));
 sg13g2_nor2_1 _14970_ (.A(_06782_),
    .B(_06792_),
    .Y(_06797_));
 sg13g2_nor2_1 _14971_ (.A(_06791_),
    .B(_06797_),
    .Y(_06798_));
 sg13g2_o21ai_1 _14972_ (.B1(_06798_),
    .Y(_06799_),
    .A1(_06784_),
    .A2(_06796_));
 sg13g2_nand2_1 _14973_ (.Y(_06800_),
    .A(\TRNG.sha256.expand.dout1[24] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[24] ));
 sg13g2_xor2_1 _14974_ (.B(\TRNG.sha256.expand.sm0.sum_0[24] ),
    .A(\TRNG.sha256.expand.dout1[24] ),
    .X(_06801_));
 sg13g2_nand2_1 _14975_ (.Y(_06802_),
    .A(\TRNG.sha256.expand.dout2[24] ),
    .B(_06801_));
 sg13g2_xnor2_1 _14976_ (.Y(_06803_),
    .A(\TRNG.sha256.expand.dout2[24] ),
    .B(_06801_));
 sg13g2_a21oi_1 _14977_ (.A1(\TRNG.sha256.expand.dout2[23] ),
    .A2(_06789_),
    .Y(_06804_),
    .B1(_06788_));
 sg13g2_nor2_1 _14978_ (.A(_06803_),
    .B(_06804_),
    .Y(_06805_));
 sg13g2_xnor2_1 _14979_ (.Y(_06806_),
    .A(_06803_),
    .B(_06804_));
 sg13g2_nor2_1 _14980_ (.A(_06799_),
    .B(_06806_),
    .Y(_06807_));
 sg13g2_xor2_1 _14981_ (.B(_06806_),
    .A(_06799_),
    .X(_00292_));
 sg13g2_and2_1 _14982_ (.A(\TRNG.sha256.expand.dout1[25] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[25] ),
    .X(_06808_));
 sg13g2_xor2_1 _14983_ (.B(\TRNG.sha256.expand.sm0.sum_0[25] ),
    .A(\TRNG.sha256.expand.dout1[25] ),
    .X(_06809_));
 sg13g2_xnor2_1 _14984_ (.Y(_06810_),
    .A(\TRNG.sha256.expand.dout2[25] ),
    .B(_06809_));
 sg13g2_a21oi_1 _14985_ (.A1(_06800_),
    .A2(_06802_),
    .Y(_06811_),
    .B1(_06810_));
 sg13g2_nand3_1 _14986_ (.B(_06802_),
    .C(_06810_),
    .A(_06800_),
    .Y(_06812_));
 sg13g2_nor2b_1 _14987_ (.A(_06811_),
    .B_N(_06812_),
    .Y(_06813_));
 sg13g2_nor2_1 _14988_ (.A(_06805_),
    .B(_06807_),
    .Y(_06814_));
 sg13g2_xnor2_1 _14989_ (.Y(_00293_),
    .A(_06813_),
    .B(_06814_));
 sg13g2_nand2b_1 _14990_ (.Y(_06815_),
    .B(_06813_),
    .A_N(_06806_));
 sg13g2_a21oi_1 _14991_ (.A1(_06805_),
    .A2(_06812_),
    .Y(_06816_),
    .B1(_06811_));
 sg13g2_o21ai_1 _14992_ (.B1(_06816_),
    .Y(_06817_),
    .A1(_06799_),
    .A2(_06815_));
 sg13g2_xor2_1 _14993_ (.B(\TRNG.sha256.expand.sm0.sum_0[26] ),
    .A(\TRNG.sha256.expand.dout1[26] ),
    .X(_06818_));
 sg13g2_and2_1 _14994_ (.A(\TRNG.sha256.expand.dout2[26] ),
    .B(_06818_),
    .X(_06819_));
 sg13g2_xnor2_1 _14995_ (.Y(_06820_),
    .A(\TRNG.sha256.expand.dout2[26] ),
    .B(_06818_));
 sg13g2_a21oi_2 _14996_ (.B1(_06808_),
    .Y(_06821_),
    .A2(_06809_),
    .A1(\TRNG.sha256.expand.dout2[25] ));
 sg13g2_nor2_1 _14997_ (.A(_06820_),
    .B(_06821_),
    .Y(_06822_));
 sg13g2_xnor2_1 _14998_ (.Y(_06823_),
    .A(_06820_),
    .B(_06821_));
 sg13g2_inv_1 _14999_ (.Y(_06824_),
    .A(_06823_));
 sg13g2_xnor2_1 _15000_ (.Y(_00294_),
    .A(_06817_),
    .B(_06823_));
 sg13g2_a21oi_2 _15001_ (.B1(_06819_),
    .Y(_06825_),
    .A2(\TRNG.sha256.expand.sm0.sum_0[26] ),
    .A1(\TRNG.sha256.expand.dout1[26] ));
 sg13g2_and2_1 _15002_ (.A(\TRNG.sha256.expand.dout1[27] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[27] ),
    .X(_06826_));
 sg13g2_xor2_1 _15003_ (.B(\TRNG.sha256.expand.sm0.sum_0[27] ),
    .A(\TRNG.sha256.expand.dout1[27] ),
    .X(_06827_));
 sg13g2_xnor2_1 _15004_ (.Y(_06828_),
    .A(\TRNG.sha256.expand.dout2[27] ),
    .B(_06827_));
 sg13g2_nand2_1 _15005_ (.Y(_06829_),
    .A(_06825_),
    .B(_06828_));
 sg13g2_xor2_1 _15006_ (.B(_06828_),
    .A(_06825_),
    .X(_06830_));
 sg13g2_a21oi_1 _15007_ (.A1(_06817_),
    .A2(_06824_),
    .Y(_06831_),
    .B1(_06822_));
 sg13g2_xnor2_1 _15008_ (.Y(_00295_),
    .A(_06830_),
    .B(_06831_));
 sg13g2_and2_1 _15009_ (.A(_06824_),
    .B(_06830_),
    .X(_06832_));
 sg13g2_nand2_1 _15010_ (.Y(_06833_),
    .A(_06822_),
    .B(_06829_));
 sg13g2_o21ai_1 _15011_ (.B1(_06833_),
    .Y(_06834_),
    .A1(_06825_),
    .A2(_06828_));
 sg13g2_a21o_1 _15012_ (.A2(_06832_),
    .A1(_06817_),
    .B1(_06834_),
    .X(_06835_));
 sg13g2_a21oi_1 _15013_ (.A1(\TRNG.sha256.expand.dout2[27] ),
    .A2(_06827_),
    .Y(_06836_),
    .B1(_06826_));
 sg13g2_nand2_1 _15014_ (.Y(_06837_),
    .A(\TRNG.sha256.expand.dout1[28] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[28] ));
 sg13g2_xor2_1 _15015_ (.B(\TRNG.sha256.expand.sm0.sum_0[28] ),
    .A(\TRNG.sha256.expand.dout1[28] ),
    .X(_06838_));
 sg13g2_nand2_1 _15016_ (.Y(_06839_),
    .A(\TRNG.sha256.expand.dout2[28] ),
    .B(_06838_));
 sg13g2_xnor2_1 _15017_ (.Y(_06840_),
    .A(\TRNG.sha256.expand.dout2[28] ),
    .B(_06838_));
 sg13g2_nor2_1 _15018_ (.A(_06836_),
    .B(_06840_),
    .Y(_06841_));
 sg13g2_xor2_1 _15019_ (.B(_06840_),
    .A(_06836_),
    .X(_06842_));
 sg13g2_xor2_1 _15020_ (.B(_06842_),
    .A(_06835_),
    .X(_00296_));
 sg13g2_a21oi_1 _15021_ (.A1(_06835_),
    .A2(_06842_),
    .Y(_06843_),
    .B1(_06841_));
 sg13g2_and2_1 _15022_ (.A(\TRNG.sha256.expand.dout1[29] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[29] ),
    .X(_06844_));
 sg13g2_xor2_1 _15023_ (.B(\TRNG.sha256.expand.sm0.sum_0[29] ),
    .A(\TRNG.sha256.expand.dout1[29] ),
    .X(_06845_));
 sg13g2_xnor2_1 _15024_ (.Y(_06846_),
    .A(\TRNG.sha256.expand.dout2[29] ),
    .B(_06845_));
 sg13g2_and3_1 _15025_ (.X(_06847_),
    .A(_06837_),
    .B(_06839_),
    .C(_06846_));
 sg13g2_a21o_1 _15026_ (.A2(_06839_),
    .A1(_06837_),
    .B1(_06846_),
    .X(_06848_));
 sg13g2_nor2b_1 _15027_ (.A(_06847_),
    .B_N(_06848_),
    .Y(_06849_));
 sg13g2_a21oi_1 _15028_ (.A1(_06843_),
    .A2(_06848_),
    .Y(_06850_),
    .B1(_06847_));
 sg13g2_xnor2_1 _15029_ (.Y(_00297_),
    .A(_06843_),
    .B(_06849_));
 sg13g2_a21oi_1 _15030_ (.A1(\TRNG.sha256.expand.dout2[29] ),
    .A2(_06845_),
    .Y(_06851_),
    .B1(_06844_));
 sg13g2_and2_1 _15031_ (.A(\TRNG.sha256.expand.dout1[30] ),
    .B(\TRNG.sha256.expand.sm0.sum_0[30] ),
    .X(_06852_));
 sg13g2_xor2_1 _15032_ (.B(\TRNG.sha256.expand.sm0.sum_0[30] ),
    .A(\TRNG.sha256.expand.dout1[30] ),
    .X(_06853_));
 sg13g2_xnor2_1 _15033_ (.Y(_06854_),
    .A(\TRNG.sha256.expand.dout2[30] ),
    .B(_06853_));
 sg13g2_nor2_1 _15034_ (.A(_06851_),
    .B(_06854_),
    .Y(_06855_));
 sg13g2_xor2_1 _15035_ (.B(_06854_),
    .A(_06851_),
    .X(_06856_));
 sg13g2_xor2_1 _15036_ (.B(_06856_),
    .A(_06850_),
    .X(_00299_));
 sg13g2_a21oi_1 _15037_ (.A1(_06850_),
    .A2(_06856_),
    .Y(_06857_),
    .B1(_06855_));
 sg13g2_a21oi_1 _15038_ (.A1(\TRNG.sha256.expand.dout2[30] ),
    .A2(_06853_),
    .Y(_06858_),
    .B1(_06852_));
 sg13g2_xnor2_1 _15039_ (.Y(_06859_),
    .A(\TRNG.sha256.expand.dout2[31] ),
    .B(\TRNG.sha256.expand.dout1[31] ));
 sg13g2_xnor2_1 _15040_ (.Y(_06860_),
    .A(\TRNG.sha256.expand.sm0.sum_0[31] ),
    .B(_06859_));
 sg13g2_xnor2_1 _15041_ (.Y(_06861_),
    .A(_06858_),
    .B(_06860_));
 sg13g2_xnor2_1 _15042_ (.Y(_00300_),
    .A(_06857_),
    .B(_06861_));
 sg13g2_xor2_1 _15043_ (.B(\TRNG.NOISE_SOURCE.Loop2.NOT2_OUT_TO_NAND1_IN2 ),
    .A(\TRNG.NOISE_SOURCE.Loop1.NOT2_OUT_TO_NAND1_IN2 ),
    .X(_06862_));
 sg13g2_xor2_1 _15044_ (.B(\TRNG.NOISE_SOURCE.Loop4.NOT2_OUT_TO_NAND1_IN2 ),
    .A(\TRNG.NOISE_SOURCE.Loop3.NOT2_OUT_TO_NAND1_IN2 ),
    .X(_06863_));
 sg13g2_xnor2_1 _15045_ (.Y(_06864_),
    .A(\TRNG.NOISE_SOURCE.Loop5.NOT2_OUT_TO_NAND1_IN2 ),
    .B(_06863_));
 sg13g2_xnor2_1 _15046_ (.Y(\TRNG.NOISE_SOURCE.Noise_Source_Out ),
    .A(_06862_),
    .B(_06864_));
 sg13g2_nor2_1 _15047_ (.A(net3392),
    .B(_05896_),
    .Y(_00308_));
 sg13g2_nand2_1 _15048_ (.Y(_06865_),
    .A(net1896),
    .B(_04831_));
 sg13g2_o21ai_1 _15049_ (.B1(_06865_),
    .Y(_00309_),
    .A1(_04884_),
    .A2(_05897_));
 sg13g2_nand2_1 _15050_ (.Y(_06866_),
    .A(net1210),
    .B(_04831_));
 sg13g2_o21ai_1 _15051_ (.B1(_06866_),
    .Y(_00310_),
    .A1(_04834_),
    .A2(_05896_));
 sg13g2_o21ai_1 _15052_ (.B1(_05917_),
    .Y(_00311_),
    .A1(net3292),
    .A2(_05897_));
 sg13g2_a21oi_1 _15053_ (.A1(_04887_),
    .A2(net2680),
    .Y(_00312_),
    .B1(_04885_));
 sg13g2_nor2_1 _15054_ (.A(net5873),
    .B(net5874),
    .Y(_06867_));
 sg13g2_or2_2 _15055_ (.X(_06868_),
    .B(net5874),
    .A(net5873));
 sg13g2_nor2_1 _15056_ (.A(\TRNG.sha256.compress.count[0] ),
    .B(\TRNG.sha256.compress.count[1] ),
    .Y(_06869_));
 sg13g2_or2_2 _15057_ (.X(_06870_),
    .B(\TRNG.sha256.compress.count[1] ),
    .A(\TRNG.sha256.compress.count[0] ));
 sg13g2_nor2_1 _15058_ (.A(_06868_),
    .B(_06870_),
    .Y(_06871_));
 sg13g2_and2_1 _15059_ (.A(_00118_),
    .B(_06871_),
    .X(_06872_));
 sg13g2_nand2_1 _15060_ (.Y(_06873_),
    .A(net3757),
    .B(_06871_));
 sg13g2_nor2_1 _15061_ (.A(net5520),
    .B(net5097),
    .Y(_06874_));
 sg13g2_nand2_2 _15062_ (.Y(_06875_),
    .A(net5472),
    .B(net5089));
 sg13g2_nor2_2 _15063_ (.A(net5847),
    .B(net4967),
    .Y(_06876_));
 sg13g2_nand2_2 _15064_ (.Y(_06877_),
    .A(net5491),
    .B(net4977));
 sg13g2_nor2_1 _15065_ (.A(net5491),
    .B(net4965),
    .Y(_06878_));
 sg13g2_a22oi_1 _15066_ (.Y(_06879_),
    .B1(net4744),
    .B2(net3521),
    .A2(_06876_),
    .A1(net3410));
 sg13g2_inv_1 _15067_ (.Y(_00313_),
    .A(_06879_));
 sg13g2_a22oi_1 _15068_ (.Y(_06880_),
    .B1(_06878_),
    .B2(net5554),
    .A2(_06876_),
    .A1(net3565));
 sg13g2_inv_1 _15069_ (.Y(_00314_),
    .A(net3566));
 sg13g2_a22oi_1 _15070_ (.Y(_06881_),
    .B1(net4745),
    .B2(net5555),
    .A2(_06876_),
    .A1(net3610));
 sg13g2_inv_1 _15071_ (.Y(_00315_),
    .A(net3611));
 sg13g2_a22oi_1 _15072_ (.Y(_06882_),
    .B1(net4744),
    .B2(net3410),
    .A2(_06876_),
    .A1(\TRNG.hash[128] ));
 sg13g2_inv_1 _15073_ (.Y(_00316_),
    .A(net3411));
 sg13g2_nand4_1 _15074_ (.B(_04277_),
    .C(\TRNG.sha256.expand.address1[2] ),
    .A(\TRNG.sha256.expand.exp_ctrl.write_en1 ),
    .Y(_06883_),
    .D(net5393));
 sg13g2_mux2_1 _15075_ (.A0(net5690),
    .A1(net3281),
    .S(net5194),
    .X(_00317_));
 sg13g2_mux2_1 _15076_ (.A0(net5687),
    .A1(net3244),
    .S(net5194),
    .X(_00318_));
 sg13g2_mux2_1 _15077_ (.A0(net5685),
    .A1(net3288),
    .S(net5196),
    .X(_00319_));
 sg13g2_nand2_1 _15078_ (.Y(_06884_),
    .A(net2413),
    .B(net5197));
 sg13g2_o21ai_1 _15079_ (.B1(_06884_),
    .Y(_00320_),
    .A1(net5494),
    .A2(net5197));
 sg13g2_mux2_1 _15080_ (.A0(net3204),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[4][4] ),
    .S(net5196),
    .X(_00321_));
 sg13g2_mux2_1 _15081_ (.A0(net5680),
    .A1(net3133),
    .S(net5196),
    .X(_00322_));
 sg13g2_mux2_1 _15082_ (.A0(net5677),
    .A1(net3322),
    .S(net5196),
    .X(_00323_));
 sg13g2_mux2_1 _15083_ (.A0(net5674),
    .A1(net3406),
    .S(net5195),
    .X(_00324_));
 sg13g2_mux2_1 _15084_ (.A0(net5672),
    .A1(net3359),
    .S(net5195),
    .X(_00325_));
 sg13g2_mux2_1 _15085_ (.A0(net5670),
    .A1(net3267),
    .S(net5196),
    .X(_00326_));
 sg13g2_mux2_1 _15086_ (.A0(net5668),
    .A1(net3324),
    .S(net5195),
    .X(_00327_));
 sg13g2_mux2_1 _15087_ (.A0(net5665),
    .A1(net3405),
    .S(net5194),
    .X(_00328_));
 sg13g2_mux2_1 _15088_ (.A0(net5662),
    .A1(net3407),
    .S(net5194),
    .X(_00329_));
 sg13g2_mux2_1 _15089_ (.A0(net5660),
    .A1(net3404),
    .S(net5194),
    .X(_00330_));
 sg13g2_mux2_1 _15090_ (.A0(net5659),
    .A1(net3328),
    .S(net5195),
    .X(_00331_));
 sg13g2_mux2_1 _15091_ (.A0(net5655),
    .A1(net3373),
    .S(net5193),
    .X(_00332_));
 sg13g2_mux2_1 _15092_ (.A0(net5654),
    .A1(net3319),
    .S(net5195),
    .X(_00333_));
 sg13g2_mux2_1 _15093_ (.A0(net5651),
    .A1(net3224),
    .S(net5197),
    .X(_00334_));
 sg13g2_mux2_1 _15094_ (.A0(net5650),
    .A1(net3335),
    .S(net5194),
    .X(_00335_));
 sg13g2_mux2_1 _15095_ (.A0(net5646),
    .A1(net3249),
    .S(net5194),
    .X(_00336_));
 sg13g2_mux2_1 _15096_ (.A0(net5643),
    .A1(net3374),
    .S(net5193),
    .X(_00337_));
 sg13g2_mux2_1 _15097_ (.A0(net5641),
    .A1(net3414),
    .S(net5193),
    .X(_00338_));
 sg13g2_mux2_1 _15098_ (.A0(net5638),
    .A1(net3368),
    .S(net5193),
    .X(_00339_));
 sg13g2_mux2_1 _15099_ (.A0(net5636),
    .A1(net3247),
    .S(net5193),
    .X(_00340_));
 sg13g2_mux2_1 _15100_ (.A0(net5633),
    .A1(net3306),
    .S(net5193),
    .X(_00341_));
 sg13g2_mux2_1 _15101_ (.A0(net5631),
    .A1(net3397),
    .S(net5193),
    .X(_00342_));
 sg13g2_mux2_1 _15102_ (.A0(net5629),
    .A1(net3261),
    .S(net5193),
    .X(_00343_));
 sg13g2_mux2_1 _15103_ (.A0(net5627),
    .A1(net3280),
    .S(net5196),
    .X(_00344_));
 sg13g2_mux2_1 _15104_ (.A0(net5624),
    .A1(net3246),
    .S(net5195),
    .X(_00345_));
 sg13g2_mux2_1 _15105_ (.A0(net5621),
    .A1(net3202),
    .S(net5195),
    .X(_00346_));
 sg13g2_mux2_1 _15106_ (.A0(net5619),
    .A1(net3332),
    .S(net5196),
    .X(_00347_));
 sg13g2_mux2_1 _15107_ (.A0(net5616),
    .A1(net3390),
    .S(net5195),
    .X(_00348_));
 sg13g2_nand2_2 _15108_ (.Y(_06885_),
    .A(\TRNG.sha256.expand.exp_ctrl.write_en1 ),
    .B(net5370));
 sg13g2_nor2_1 _15109_ (.A(net5202),
    .B(_06885_),
    .Y(_06886_));
 sg13g2_mux2_1 _15110_ (.A0(net3252),
    .A1(net5690),
    .S(net5084),
    .X(_00349_));
 sg13g2_mux2_1 _15111_ (.A0(net3137),
    .A1(net5687),
    .S(net5084),
    .X(_00350_));
 sg13g2_mux2_1 _15112_ (.A0(net3234),
    .A1(net5684),
    .S(net5085),
    .X(_00351_));
 sg13g2_nor2_1 _15113_ (.A(net2626),
    .B(net5086),
    .Y(_06887_));
 sg13g2_a21oi_1 _15114_ (.A1(net5494),
    .A2(net5086),
    .Y(_00352_),
    .B1(_06887_));
 sg13g2_mux2_1 _15115_ (.A0(net3111),
    .A1(net5683),
    .S(net5085),
    .X(_00353_));
 sg13g2_mux2_1 _15116_ (.A0(net3042),
    .A1(net5680),
    .S(net5085),
    .X(_00354_));
 sg13g2_mux2_1 _15117_ (.A0(net2973),
    .A1(net5676),
    .S(net5085),
    .X(_00355_));
 sg13g2_mux2_1 _15118_ (.A0(net3233),
    .A1(net5674),
    .S(net5087),
    .X(_00356_));
 sg13g2_mux2_1 _15119_ (.A0(net3072),
    .A1(net5672),
    .S(net5085),
    .X(_00357_));
 sg13g2_mux2_1 _15120_ (.A0(net2823),
    .A1(net5670),
    .S(net5088),
    .X(_00358_));
 sg13g2_mux2_1 _15121_ (.A0(net2919),
    .A1(net5667),
    .S(net5088),
    .X(_00359_));
 sg13g2_mux2_1 _15122_ (.A0(net3011),
    .A1(net5665),
    .S(net5084),
    .X(_00360_));
 sg13g2_mux2_1 _15123_ (.A0(net2951),
    .A1(net5662),
    .S(net5084),
    .X(_00361_));
 sg13g2_mux2_1 _15124_ (.A0(net3176),
    .A1(net5660),
    .S(net5084),
    .X(_00362_));
 sg13g2_mux2_1 _15125_ (.A0(net3376),
    .A1(\TRNG.sha256.expand.data1_to_ram[14] ),
    .S(net5087),
    .X(_00363_));
 sg13g2_mux2_1 _15126_ (.A0(net2851),
    .A1(net5655),
    .S(net5084),
    .X(_00364_));
 sg13g2_mux2_1 _15127_ (.A0(net3372),
    .A1(net5653),
    .S(net5087),
    .X(_00365_));
 sg13g2_mux2_1 _15128_ (.A0(net3016),
    .A1(net5651),
    .S(net5086),
    .X(_00366_));
 sg13g2_mux2_1 _15129_ (.A0(net2756),
    .A1(net5648),
    .S(net5084),
    .X(_00367_));
 sg13g2_mux2_1 _15130_ (.A0(net3387),
    .A1(net5646),
    .S(net5084),
    .X(_00368_));
 sg13g2_mux2_1 _15131_ (.A0(net3024),
    .A1(net5644),
    .S(net5086),
    .X(_00369_));
 sg13g2_mux2_1 _15132_ (.A0(net3113),
    .A1(net5640),
    .S(net5086),
    .X(_00370_));
 sg13g2_mux2_1 _15133_ (.A0(net3162),
    .A1(net5637),
    .S(net5086),
    .X(_00371_));
 sg13g2_mux2_1 _15134_ (.A0(net3226),
    .A1(net5635),
    .S(net5087),
    .X(_00372_));
 sg13g2_mux2_1 _15135_ (.A0(net3196),
    .A1(net5633),
    .S(net5087),
    .X(_00373_));
 sg13g2_mux2_1 _15136_ (.A0(net2848),
    .A1(net5632),
    .S(net5086),
    .X(_00374_));
 sg13g2_mux2_1 _15137_ (.A0(net2975),
    .A1(net5630),
    .S(net5086),
    .X(_00375_));
 sg13g2_mux2_1 _15138_ (.A0(net3061),
    .A1(net5627),
    .S(net5085),
    .X(_00376_));
 sg13g2_mux2_1 _15139_ (.A0(net2895),
    .A1(net5625),
    .S(net5087),
    .X(_00377_));
 sg13g2_mux2_1 _15140_ (.A0(net2955),
    .A1(net5622),
    .S(net5088),
    .X(_00378_));
 sg13g2_mux2_1 _15141_ (.A0(net2797),
    .A1(net5619),
    .S(net5085),
    .X(_00379_));
 sg13g2_mux2_1 _15142_ (.A0(net3187),
    .A1(net5616),
    .S(net5087),
    .X(_00380_));
 sg13g2_nor2_1 _15143_ (.A(net5360),
    .B(_06885_),
    .Y(_06888_));
 sg13g2_mux2_1 _15144_ (.A0(net3038),
    .A1(net5689),
    .S(net5075),
    .X(_00381_));
 sg13g2_nand2_1 _15145_ (.Y(_06889_),
    .A(net5688),
    .B(net5076));
 sg13g2_o21ai_1 _15146_ (.B1(_06889_),
    .Y(_00382_),
    .A1(_04344_),
    .A2(net5075));
 sg13g2_mux2_1 _15147_ (.A0(net3236),
    .A1(net5684),
    .S(net5077),
    .X(_00383_));
 sg13g2_nor2_1 _15148_ (.A(net3212),
    .B(net5079),
    .Y(_06890_));
 sg13g2_a21oi_1 _15149_ (.A1(net5496),
    .A2(net5079),
    .Y(_00384_),
    .B1(_06890_));
 sg13g2_mux2_1 _15150_ (.A0(net3142),
    .A1(net5683),
    .S(net5077),
    .X(_00385_));
 sg13g2_nand2_1 _15151_ (.Y(_06891_),
    .A(net5681),
    .B(net5077));
 sg13g2_o21ai_1 _15152_ (.B1(_06891_),
    .Y(_00386_),
    .A1(_04347_),
    .A2(net5077));
 sg13g2_nand2_1 _15153_ (.Y(_06892_),
    .A(net5676),
    .B(net5077));
 sg13g2_o21ai_1 _15154_ (.B1(_06892_),
    .Y(_00387_),
    .A1(_04348_),
    .A2(net5077));
 sg13g2_nand2_1 _15155_ (.Y(_06893_),
    .A(net5675),
    .B(net5082));
 sg13g2_o21ai_1 _15156_ (.B1(_06893_),
    .Y(_00388_),
    .A1(_04349_),
    .A2(net5082));
 sg13g2_mux2_1 _15157_ (.A0(net3303),
    .A1(net5671),
    .S(net5078),
    .X(_00389_));
 sg13g2_nand2_1 _15158_ (.Y(_06894_),
    .A(net5669),
    .B(net5081));
 sg13g2_o21ai_1 _15159_ (.B1(_06894_),
    .Y(_00390_),
    .A1(_04351_),
    .A2(net5081));
 sg13g2_mux2_1 _15160_ (.A0(net2965),
    .A1(net5667),
    .S(net5081),
    .X(_00391_));
 sg13g2_nand2_1 _15161_ (.Y(_06895_),
    .A(net5666),
    .B(net5076));
 sg13g2_o21ai_1 _15162_ (.B1(_06895_),
    .Y(_00392_),
    .A1(_04353_),
    .A2(net5076));
 sg13g2_nand2_1 _15163_ (.Y(_06896_),
    .A(net5663),
    .B(net5075));
 sg13g2_o21ai_1 _15164_ (.B1(_06896_),
    .Y(_00393_),
    .A1(_04354_),
    .A2(net5075));
 sg13g2_nand2_1 _15165_ (.Y(_06897_),
    .A(net5661),
    .B(net5075));
 sg13g2_o21ai_1 _15166_ (.B1(_06897_),
    .Y(_00394_),
    .A1(_04355_),
    .A2(net5075));
 sg13g2_mux2_1 _15167_ (.A0(net2821),
    .A1(net5658),
    .S(net5082),
    .X(_00395_));
 sg13g2_nand2_1 _15168_ (.Y(_06898_),
    .A(net5656),
    .B(net5076));
 sg13g2_o21ai_1 _15169_ (.B1(_06898_),
    .Y(_00396_),
    .A1(_04357_),
    .A2(net5076));
 sg13g2_mux2_1 _15170_ (.A0(net2981),
    .A1(net5653),
    .S(net5081),
    .X(_00397_));
 sg13g2_nand2_1 _15171_ (.Y(_06899_),
    .A(\TRNG.sha256.expand.data1_to_ram[17] ),
    .B(net5079));
 sg13g2_o21ai_1 _15172_ (.B1(_06899_),
    .Y(_00398_),
    .A1(_04359_),
    .A2(net5079));
 sg13g2_nand2_1 _15173_ (.Y(_06900_),
    .A(net5649),
    .B(net5076));
 sg13g2_o21ai_1 _15174_ (.B1(_06900_),
    .Y(_00399_),
    .A1(_04360_),
    .A2(net5076));
 sg13g2_nand2_1 _15175_ (.Y(_06901_),
    .A(net5647),
    .B(net5078));
 sg13g2_o21ai_1 _15176_ (.B1(_06901_),
    .Y(_00400_),
    .A1(_04361_),
    .A2(net5078));
 sg13g2_mux2_1 _15177_ (.A0(net3025),
    .A1(net5644),
    .S(net5080),
    .X(_00401_));
 sg13g2_nand2_1 _15178_ (.Y(_06902_),
    .A(net5641),
    .B(net5079));
 sg13g2_o21ai_1 _15179_ (.B1(_06902_),
    .Y(_00402_),
    .A1(_04363_),
    .A2(net5079));
 sg13g2_mux2_1 _15180_ (.A0(net3146),
    .A1(net5638),
    .S(net5080),
    .X(_00403_));
 sg13g2_nand2_1 _15181_ (.Y(_06903_),
    .A(net5636),
    .B(net5080));
 sg13g2_o21ai_1 _15182_ (.B1(_06903_),
    .Y(_00404_),
    .A1(_04365_),
    .A2(net5080));
 sg13g2_nand2_1 _15183_ (.Y(_06904_),
    .A(net5634),
    .B(net5080));
 sg13g2_o21ai_1 _15184_ (.B1(_06904_),
    .Y(_00405_),
    .A1(_04366_),
    .A2(net5080));
 sg13g2_nand2_1 _15185_ (.Y(_06905_),
    .A(net5632),
    .B(net5079));
 sg13g2_o21ai_1 _15186_ (.B1(_06905_),
    .Y(_00406_),
    .A1(_04367_),
    .A2(net5079));
 sg13g2_mux2_1 _15187_ (.A0(net2810),
    .A1(net5630),
    .S(net5081),
    .X(_00407_));
 sg13g2_nand2_1 _15188_ (.Y(_06906_),
    .A(net5627),
    .B(net5075));
 sg13g2_o21ai_1 _15189_ (.B1(_06906_),
    .Y(_00408_),
    .A1(_04369_),
    .A2(net5075));
 sg13g2_mux2_1 _15190_ (.A0(net2967),
    .A1(net5625),
    .S(net5082),
    .X(_00409_));
 sg13g2_nand2_1 _15191_ (.Y(_06907_),
    .A(net5621),
    .B(net5081));
 sg13g2_o21ai_1 _15192_ (.B1(_06907_),
    .Y(_00410_),
    .A1(_04371_),
    .A2(net5081));
 sg13g2_nand2_1 _15193_ (.Y(_06908_),
    .A(net5618),
    .B(net5077));
 sg13g2_o21ai_1 _15194_ (.B1(_06908_),
    .Y(_00411_),
    .A1(_04372_),
    .A2(net5077));
 sg13g2_nand2_1 _15195_ (.Y(_06909_),
    .A(net5617),
    .B(net5082));
 sg13g2_o21ai_1 _15196_ (.B1(_06909_),
    .Y(_00412_),
    .A1(_04373_),
    .A2(net5081));
 sg13g2_nand2_2 _15197_ (.Y(_06910_),
    .A(\TRNG.sha256.expand.exp_ctrl.write_en1 ),
    .B(net5417));
 sg13g2_nor2_1 _15198_ (.A(net5202),
    .B(_06910_),
    .Y(_06911_));
 sg13g2_mux2_1 _15199_ (.A0(net2804),
    .A1(net5690),
    .S(net5070),
    .X(_00413_));
 sg13g2_mux2_1 _15200_ (.A0(net2723),
    .A1(net5687),
    .S(net5070),
    .X(_00414_));
 sg13g2_mux2_1 _15201_ (.A0(net2565),
    .A1(net5684),
    .S(net5071),
    .X(_00415_));
 sg13g2_nor2_1 _15202_ (.A(net3002),
    .B(net5072),
    .Y(_06912_));
 sg13g2_a21oi_1 _15203_ (.A1(net5495),
    .A2(net5072),
    .Y(_00416_),
    .B1(_06912_));
 sg13g2_mux2_1 _15204_ (.A0(net2687),
    .A1(net5683),
    .S(net5071),
    .X(_00417_));
 sg13g2_mux2_1 _15205_ (.A0(net3172),
    .A1(net5679),
    .S(net5071),
    .X(_00418_));
 sg13g2_mux2_1 _15206_ (.A0(net3136),
    .A1(net5677),
    .S(net5071),
    .X(_00419_));
 sg13g2_mux2_1 _15207_ (.A0(net2979),
    .A1(net5674),
    .S(net5073),
    .X(_00420_));
 sg13g2_mux2_1 _15208_ (.A0(net2840),
    .A1(net5672),
    .S(net5071),
    .X(_00421_));
 sg13g2_mux2_1 _15209_ (.A0(net2731),
    .A1(net5670),
    .S(net5074),
    .X(_00422_));
 sg13g2_mux2_1 _15210_ (.A0(net2507),
    .A1(net5667),
    .S(net5074),
    .X(_00423_));
 sg13g2_mux2_1 _15211_ (.A0(net2829),
    .A1(net5665),
    .S(net5070),
    .X(_00424_));
 sg13g2_mux2_1 _15212_ (.A0(net3048),
    .A1(net5662),
    .S(net5070),
    .X(_00425_));
 sg13g2_mux2_1 _15213_ (.A0(net2852),
    .A1(net5660),
    .S(net5070),
    .X(_00426_));
 sg13g2_mux2_1 _15214_ (.A0(net2489),
    .A1(net5658),
    .S(net5073),
    .X(_00427_));
 sg13g2_mux2_1 _15215_ (.A0(net2816),
    .A1(net5655),
    .S(net5070),
    .X(_00428_));
 sg13g2_mux2_1 _15216_ (.A0(net2962),
    .A1(net5653),
    .S(net5073),
    .X(_00429_));
 sg13g2_mux2_1 _15217_ (.A0(net3052),
    .A1(net5651),
    .S(net5072),
    .X(_00430_));
 sg13g2_mux2_1 _15218_ (.A0(net3200),
    .A1(net5648),
    .S(net5070),
    .X(_00431_));
 sg13g2_mux2_1 _15219_ (.A0(net3004),
    .A1(net5646),
    .S(net5070),
    .X(_00432_));
 sg13g2_mux2_1 _15220_ (.A0(net2696),
    .A1(net5644),
    .S(net5072),
    .X(_00433_));
 sg13g2_mux2_1 _15221_ (.A0(net3240),
    .A1(net5640),
    .S(net5072),
    .X(_00434_));
 sg13g2_mux2_1 _15222_ (.A0(net2538),
    .A1(net5637),
    .S(net5072),
    .X(_00435_));
 sg13g2_mux2_1 _15223_ (.A0(net2906),
    .A1(net5635),
    .S(net5073),
    .X(_00436_));
 sg13g2_mux2_1 _15224_ (.A0(net3043),
    .A1(net5633),
    .S(net5073),
    .X(_00437_));
 sg13g2_mux2_1 _15225_ (.A0(net3156),
    .A1(net5631),
    .S(net5072),
    .X(_00438_));
 sg13g2_mux2_1 _15226_ (.A0(net2562),
    .A1(net5630),
    .S(net5072),
    .X(_00439_));
 sg13g2_mux2_1 _15227_ (.A0(net2833),
    .A1(\TRNG.sha256.expand.data1_to_ram[27] ),
    .S(net5071),
    .X(_00440_));
 sg13g2_mux2_1 _15228_ (.A0(net2515),
    .A1(net5625),
    .S(net5073),
    .X(_00441_));
 sg13g2_mux2_1 _15229_ (.A0(net3003),
    .A1(net5622),
    .S(net5074),
    .X(_00442_));
 sg13g2_mux2_1 _15230_ (.A0(net3144),
    .A1(net5619),
    .S(net5071),
    .X(_00443_));
 sg13g2_mux2_1 _15231_ (.A0(net2926),
    .A1(net5616),
    .S(net5073),
    .X(_00444_));
 sg13g2_nand2_2 _15232_ (.Y(_06913_),
    .A(\TRNG.sha256.expand.exp_ctrl.write_en1 ),
    .B(net5439));
 sg13g2_nor2_1 _15233_ (.A(net5202),
    .B(_06913_),
    .Y(_06914_));
 sg13g2_mux2_1 _15234_ (.A0(net2791),
    .A1(net5690),
    .S(net5065),
    .X(_00445_));
 sg13g2_mux2_1 _15235_ (.A0(net2946),
    .A1(net5687),
    .S(net5065),
    .X(_00446_));
 sg13g2_mux2_1 _15236_ (.A0(net2793),
    .A1(net5684),
    .S(net5066),
    .X(_00447_));
 sg13g2_nor2_1 _15237_ (.A(net2930),
    .B(net5067),
    .Y(_06915_));
 sg13g2_a21oi_1 _15238_ (.A1(net5494),
    .A2(net5067),
    .Y(_00448_),
    .B1(_06915_));
 sg13g2_mux2_1 _15239_ (.A0(net2705),
    .A1(net5683),
    .S(net5066),
    .X(_00449_));
 sg13g2_mux2_1 _15240_ (.A0(net2668),
    .A1(net5679),
    .S(net5066),
    .X(_00450_));
 sg13g2_mux2_1 _15241_ (.A0(net2887),
    .A1(net5677),
    .S(net5066),
    .X(_00451_));
 sg13g2_mux2_1 _15242_ (.A0(net2619),
    .A1(net5674),
    .S(net5068),
    .X(_00452_));
 sg13g2_mux2_1 _15243_ (.A0(net2945),
    .A1(net5672),
    .S(net5066),
    .X(_00453_));
 sg13g2_mux2_1 _15244_ (.A0(net3138),
    .A1(net5670),
    .S(net5069),
    .X(_00454_));
 sg13g2_mux2_1 _15245_ (.A0(net3084),
    .A1(net5667),
    .S(net5069),
    .X(_00455_));
 sg13g2_mux2_1 _15246_ (.A0(net3121),
    .A1(net5665),
    .S(net5065),
    .X(_00456_));
 sg13g2_mux2_1 _15247_ (.A0(net3075),
    .A1(net5662),
    .S(net5065),
    .X(_00457_));
 sg13g2_mux2_1 _15248_ (.A0(net2969),
    .A1(net5660),
    .S(net5065),
    .X(_00458_));
 sg13g2_mux2_1 _15249_ (.A0(net3086),
    .A1(net5658),
    .S(net5068),
    .X(_00459_));
 sg13g2_mux2_1 _15250_ (.A0(net3014),
    .A1(net5655),
    .S(net5065),
    .X(_00460_));
 sg13g2_mux2_1 _15251_ (.A0(net3053),
    .A1(net5653),
    .S(net5068),
    .X(_00461_));
 sg13g2_mux2_1 _15252_ (.A0(net2825),
    .A1(net5651),
    .S(net5067),
    .X(_00462_));
 sg13g2_mux2_1 _15253_ (.A0(net2942),
    .A1(net5648),
    .S(net5065),
    .X(_00463_));
 sg13g2_mux2_1 _15254_ (.A0(net3238),
    .A1(net5646),
    .S(net5065),
    .X(_00464_));
 sg13g2_mux2_1 _15255_ (.A0(net2722),
    .A1(net5643),
    .S(net5067),
    .X(_00465_));
 sg13g2_mux2_1 _15256_ (.A0(net2960),
    .A1(net5640),
    .S(net5067),
    .X(_00466_));
 sg13g2_mux2_1 _15257_ (.A0(net2904),
    .A1(net5637),
    .S(net5067),
    .X(_00467_));
 sg13g2_mux2_1 _15258_ (.A0(net2699),
    .A1(net5635),
    .S(net5068),
    .X(_00468_));
 sg13g2_mux2_1 _15259_ (.A0(net3012),
    .A1(net5633),
    .S(net5068),
    .X(_00469_));
 sg13g2_mux2_1 _15260_ (.A0(net2972),
    .A1(net5631),
    .S(net5067),
    .X(_00470_));
 sg13g2_mux2_1 _15261_ (.A0(net2801),
    .A1(net5630),
    .S(net5067),
    .X(_00471_));
 sg13g2_mux2_1 _15262_ (.A0(net2654),
    .A1(net5627),
    .S(net5066),
    .X(_00472_));
 sg13g2_mux2_1 _15263_ (.A0(net2977),
    .A1(net5624),
    .S(net5068),
    .X(_00473_));
 sg13g2_mux2_1 _15264_ (.A0(net2953),
    .A1(net5621),
    .S(net5069),
    .X(_00474_));
 sg13g2_mux2_1 _15265_ (.A0(net3022),
    .A1(net5619),
    .S(net5066),
    .X(_00475_));
 sg13g2_mux2_1 _15266_ (.A0(net2613),
    .A1(net5616),
    .S(net5068),
    .X(_00476_));
 sg13g2_nand2_1 _15267_ (.Y(_06916_),
    .A(net3563),
    .B(net4744));
 sg13g2_nand2_1 _15268_ (.Y(_06917_),
    .A(net5572),
    .B(\TRNG.hash[129] ));
 sg13g2_xor2_1 _15269_ (.B(_06917_),
    .A(\TRNG.hash[130] ),
    .X(_06918_));
 sg13g2_o21ai_1 _15270_ (.B1(_06916_),
    .Y(_00477_),
    .A1(net4746),
    .A2(_06918_));
 sg13g2_nor2_2 _15271_ (.A(_04228_),
    .B(net5844),
    .Y(_06919_));
 sg13g2_nand2_2 _15272_ (.Y(_06920_),
    .A(net5573),
    .B(net5490));
 sg13g2_and2_1 _15273_ (.A(\TRNG.hash[129] ),
    .B(\TRNG.hash[130] ),
    .X(_06921_));
 sg13g2_nor3_1 _15274_ (.A(\TRNG.hash[132] ),
    .B(\TRNG.hash[131] ),
    .C(_06921_),
    .Y(_06922_));
 sg13g2_nand2_1 _15275_ (.Y(_06923_),
    .A(net3643),
    .B(_06922_));
 sg13g2_xnor2_1 _15276_ (.Y(_06924_),
    .A(net3508),
    .B(_06923_));
 sg13g2_nand2_1 _15277_ (.Y(_06925_),
    .A(net5183),
    .B(net3509));
 sg13g2_nor2_2 _15278_ (.A(net5573),
    .B(net5857),
    .Y(_06926_));
 sg13g2_nand2_1 _15279_ (.Y(_06927_),
    .A(_04228_),
    .B(net5488));
 sg13g2_a22oi_1 _15280_ (.Y(_06928_),
    .B1(\TRNG.hash[134] ),
    .B2(net5345),
    .A2(net5831),
    .A1(\TRNG.hash[166] ));
 sg13g2_a21oi_1 _15281_ (.A1(_06925_),
    .A2(_06928_),
    .Y(_00478_),
    .B1(net4961));
 sg13g2_nand2_1 _15282_ (.Y(_06929_),
    .A(net3686),
    .B(net4744));
 sg13g2_nand2b_1 _15283_ (.Y(_06930_),
    .B(_06922_),
    .A_N(\TRNG.hash[133] ));
 sg13g2_and2_1 _15284_ (.A(\TRNG.hash[134] ),
    .B(_06930_),
    .X(_06931_));
 sg13g2_nand2_1 _15285_ (.Y(_06932_),
    .A(net5572),
    .B(_06931_));
 sg13g2_xnor2_1 _15286_ (.Y(_06933_),
    .A(_04300_),
    .B(_06932_));
 sg13g2_o21ai_1 _15287_ (.B1(_06929_),
    .Y(_00479_),
    .A1(net4747),
    .A2(_06933_));
 sg13g2_nand2_1 _15288_ (.Y(_06934_),
    .A(\TRNG.hash[135] ),
    .B(_06931_));
 sg13g2_a21oi_1 _15289_ (.A1(\TRNG.hash[135] ),
    .A2(_06931_),
    .Y(_06935_),
    .B1(\TRNG.hash[136] ));
 sg13g2_nor2_1 _15290_ (.A(_04228_),
    .B(_06935_),
    .Y(_06936_));
 sg13g2_xnor2_1 _15291_ (.Y(_06937_),
    .A(\TRNG.hash[137] ),
    .B(_06936_));
 sg13g2_nand2_1 _15292_ (.Y(_06938_),
    .A(net3497),
    .B(net4744));
 sg13g2_o21ai_1 _15293_ (.B1(_06938_),
    .Y(_00480_),
    .A1(net4747),
    .A2(_06937_));
 sg13g2_nand2b_1 _15294_ (.Y(_06939_),
    .B(\TRNG.hash[137] ),
    .A_N(_06935_));
 sg13g2_o21ai_1 _15295_ (.B1(_00136_),
    .Y(_06940_),
    .A1(\TRNG.hash[138] ),
    .A2(_06939_));
 sg13g2_nand2_1 _15296_ (.Y(_06941_),
    .A(\TRNG.hash[139] ),
    .B(_06940_));
 sg13g2_o21ai_1 _15297_ (.B1(net5183),
    .Y(_06942_),
    .A1(\TRNG.hash[139] ),
    .A2(_06940_));
 sg13g2_nand2b_1 _15298_ (.Y(_06943_),
    .B(_06941_),
    .A_N(_06942_));
 sg13g2_a22oi_1 _15299_ (.Y(_06944_),
    .B1(net3648),
    .B2(net5345),
    .A2(\TRNG.hash[171] ),
    .A1(net5829));
 sg13g2_a21oi_1 _15300_ (.A1(_06943_),
    .A2(net3649),
    .Y(_00481_),
    .B1(net4961));
 sg13g2_nand2b_1 _15301_ (.Y(_06945_),
    .B(_06939_),
    .A_N(\TRNG.hash[138] ));
 sg13g2_nand3b_1 _15302_ (.B(\TRNG.hash[139] ),
    .C(_06945_),
    .Y(_06946_),
    .A_N(\TRNG.hash[140] ));
 sg13g2_nand3_1 _15303_ (.B(_00138_),
    .C(_06946_),
    .A(_04233_),
    .Y(_06947_));
 sg13g2_nor3_2 _15304_ (.A(\TRNG.hash[143] ),
    .B(\TRNG.hash[142] ),
    .C(_06947_),
    .Y(_06948_));
 sg13g2_nor2b_1 _15305_ (.A(\TRNG.hash[144] ),
    .B_N(_06948_),
    .Y(_06949_));
 sg13g2_and2_1 _15306_ (.A(_04231_),
    .B(_06949_),
    .X(_06950_));
 sg13g2_and3_1 _15307_ (.X(_06951_),
    .A(_04229_),
    .B(_04230_),
    .C(_06950_));
 sg13g2_xor2_1 _15308_ (.B(_06951_),
    .A(net3482),
    .X(_06952_));
 sg13g2_nand2_1 _15309_ (.Y(_06953_),
    .A(net5185),
    .B(_06952_));
 sg13g2_a22oi_1 _15310_ (.Y(_06954_),
    .B1(\TRNG.hash[148] ),
    .B2(net5346),
    .A2(\TRNG.hash[180] ),
    .A1(net5833));
 sg13g2_a21oi_1 _15311_ (.A1(_06953_),
    .A2(_06954_),
    .Y(_00482_),
    .B1(net4960));
 sg13g2_nor2b_2 _15312_ (.A(_06951_),
    .B_N(\TRNG.hash[148] ),
    .Y(_06955_));
 sg13g2_xnor2_1 _15313_ (.Y(_06956_),
    .A(_00139_),
    .B(_06955_));
 sg13g2_nand2_1 _15314_ (.Y(_06957_),
    .A(net5185),
    .B(_06956_));
 sg13g2_a22oi_1 _15315_ (.Y(_06958_),
    .B1(net3616),
    .B2(net5348),
    .A2(net5841),
    .A1(\TRNG.hash[181] ));
 sg13g2_a21oi_1 _15316_ (.A1(_06957_),
    .A2(net3617),
    .Y(_00483_),
    .B1(net4963));
 sg13g2_nand2_1 _15317_ (.Y(_06959_),
    .A(\TRNG.hash[149] ),
    .B(_06955_));
 sg13g2_o21ai_1 _15318_ (.B1(net3645),
    .Y(_06960_),
    .A1(\TRNG.hash[150] ),
    .A2(_06959_));
 sg13g2_nand2_1 _15319_ (.Y(_06961_),
    .A(\TRNG.hash[151] ),
    .B(_06960_));
 sg13g2_o21ai_1 _15320_ (.B1(net5185),
    .Y(_06962_),
    .A1(\TRNG.hash[151] ),
    .A2(_06960_));
 sg13g2_nand2b_1 _15321_ (.Y(_06963_),
    .B(_06961_),
    .A_N(_06962_));
 sg13g2_a22oi_1 _15322_ (.Y(_06964_),
    .B1(net3854),
    .B2(net5348),
    .A2(net3805),
    .A1(net5841));
 sg13g2_a21oi_1 _15323_ (.A1(_06963_),
    .A2(_06964_),
    .Y(_00484_),
    .B1(net4963));
 sg13g2_a21oi_1 _15324_ (.A1(\TRNG.hash[149] ),
    .A2(_06955_),
    .Y(_06965_),
    .B1(\TRNG.hash[150] ));
 sg13g2_nand2b_1 _15325_ (.Y(_06966_),
    .B(\TRNG.hash[151] ),
    .A_N(\TRNG.hash[152] ));
 sg13g2_o21ai_1 _15326_ (.B1(_00141_),
    .Y(_06967_),
    .A1(_06965_),
    .A2(_06966_));
 sg13g2_and2_1 _15327_ (.A(\TRNG.hash[153] ),
    .B(_06967_),
    .X(_06968_));
 sg13g2_inv_1 _15328_ (.Y(_06969_),
    .A(_06968_));
 sg13g2_o21ai_1 _15329_ (.B1(net5185),
    .Y(_06970_),
    .A1(\TRNG.hash[153] ),
    .A2(_06967_));
 sg13g2_or2_1 _15330_ (.X(_06971_),
    .B(_06970_),
    .A(_06968_));
 sg13g2_a22oi_1 _15331_ (.Y(_06972_),
    .B1(net3793),
    .B2(net5348),
    .A2(\TRNG.hash[185] ),
    .A1(net5843));
 sg13g2_a21oi_1 _15332_ (.A1(_06971_),
    .A2(net3794),
    .Y(_00485_),
    .B1(net4962));
 sg13g2_o21ai_1 _15333_ (.B1(_00143_),
    .Y(_06973_),
    .A1(\TRNG.hash[154] ),
    .A2(_06969_));
 sg13g2_xnor2_1 _15334_ (.Y(_06974_),
    .A(net3541),
    .B(_06973_));
 sg13g2_nand2_1 _15335_ (.Y(_06975_),
    .A(net5183),
    .B(net3542));
 sg13g2_a22oi_1 _15336_ (.Y(_06976_),
    .B1(\TRNG.hash[155] ),
    .B2(net5346),
    .A2(net5835),
    .A1(\TRNG.hash[187] ));
 sg13g2_a21oi_1 _15337_ (.A1(_06975_),
    .A2(_06976_),
    .Y(_00486_),
    .B1(net4960));
 sg13g2_a21o_1 _15338_ (.A2(_06973_),
    .A1(\TRNG.hash[155] ),
    .B1(\TRNG.hash[156] ),
    .X(_06977_));
 sg13g2_and2_1 _15339_ (.A(\TRNG.hash[156] ),
    .B(\TRNG.hash[155] ),
    .X(_06978_));
 sg13g2_nand2_1 _15340_ (.Y(_06979_),
    .A(_06973_),
    .B(_06978_));
 sg13g2_nand3_1 _15341_ (.B(_06977_),
    .C(_06979_),
    .A(net5183),
    .Y(_06980_));
 sg13g2_a22oi_1 _15342_ (.Y(_06981_),
    .B1(\TRNG.hash[156] ),
    .B2(net5346),
    .A2(net5833),
    .A1(net2591));
 sg13g2_a21oi_1 _15343_ (.A1(_06980_),
    .A2(net2592),
    .Y(_00487_),
    .B1(net4960));
 sg13g2_o21ai_1 _15344_ (.B1(_06978_),
    .Y(_06982_),
    .A1(\TRNG.hash[154] ),
    .A2(_06968_));
 sg13g2_inv_1 _15345_ (.Y(_06983_),
    .A(_06982_));
 sg13g2_nand2_1 _15346_ (.Y(_06984_),
    .A(_00145_),
    .B(_06982_));
 sg13g2_xnor2_1 _15347_ (.Y(_06985_),
    .A(net3505),
    .B(_06984_));
 sg13g2_nand2_1 _15348_ (.Y(_06986_),
    .A(net5185),
    .B(net3506));
 sg13g2_a22oi_1 _15349_ (.Y(_06987_),
    .B1(\TRNG.hash[158] ),
    .B2(net5347),
    .A2(\TRNG.hash[190] ),
    .A1(net5843));
 sg13g2_a21oi_1 _15350_ (.A1(_06986_),
    .A2(_06987_),
    .Y(_00488_),
    .B1(net4962));
 sg13g2_a21oi_1 _15351_ (.A1(\TRNG.hash[0] ),
    .A2(net5177),
    .Y(_06988_),
    .B1(\TRNG.hash[1] ));
 sg13g2_and2_2 _15352_ (.A(\TRNG.hash[0] ),
    .B(\TRNG.hash[1] ),
    .X(_06989_));
 sg13g2_and2_1 _15353_ (.A(net5573),
    .B(_06989_),
    .X(_06990_));
 sg13g2_nor3_1 _15354_ (.A(net4748),
    .B(_06988_),
    .C(_06990_),
    .Y(_06991_));
 sg13g2_a21o_1 _15355_ (.A2(net4745),
    .A1(net3745),
    .B1(_06991_),
    .X(_00489_));
 sg13g2_nor3_1 _15356_ (.A(net5856),
    .B(\TRNG.hash[2] ),
    .C(_06990_),
    .Y(_06992_));
 sg13g2_nand3_1 _15357_ (.B(net5192),
    .C(_06989_),
    .A(\TRNG.hash[2] ),
    .Y(_06993_));
 sg13g2_o21ai_1 _15358_ (.B1(_06993_),
    .Y(_06994_),
    .A1(net5491),
    .A2(net3689));
 sg13g2_nor3_1 _15359_ (.A(net4966),
    .B(_06992_),
    .C(net3690),
    .Y(_00490_));
 sg13g2_a21oi_2 _15360_ (.B1(\TRNG.hash[3] ),
    .Y(_06995_),
    .A2(_06989_),
    .A1(\TRNG.hash[2] ));
 sg13g2_nand2_1 _15361_ (.Y(_06996_),
    .A(_00150_),
    .B(_06995_));
 sg13g2_xnor2_1 _15362_ (.Y(_06997_),
    .A(net3546),
    .B(_06996_));
 sg13g2_nand2_1 _15363_ (.Y(_06998_),
    .A(net5190),
    .B(net3547));
 sg13g2_a22oi_1 _15364_ (.Y(_06999_),
    .B1(\TRNG.hash[5] ),
    .B2(net5356),
    .A2(net5867),
    .A1(\TRNG.hash[37] ));
 sg13g2_a21oi_1 _15365_ (.A1(_06998_),
    .A2(_06999_),
    .Y(_00491_),
    .B1(net4970));
 sg13g2_nand2b_1 _15366_ (.Y(_07000_),
    .B(_06995_),
    .A_N(\TRNG.hash[4] ));
 sg13g2_and2_1 _15367_ (.A(\TRNG.hash[5] ),
    .B(_07000_),
    .X(_07001_));
 sg13g2_xnor2_1 _15368_ (.Y(_07002_),
    .A(net3583),
    .B(_07001_));
 sg13g2_nand2_1 _15369_ (.Y(_07003_),
    .A(net5190),
    .B(_07002_));
 sg13g2_a22oi_1 _15370_ (.Y(_07004_),
    .B1(\TRNG.hash[6] ),
    .B2(net5356),
    .A2(\TRNG.hash[38] ),
    .A1(net5869));
 sg13g2_a21oi_1 _15371_ (.A1(_07003_),
    .A2(_07004_),
    .Y(_00492_),
    .B1(net4970));
 sg13g2_nand2_1 _15372_ (.Y(_07005_),
    .A(net3461),
    .B(net4745));
 sg13g2_nand3_1 _15373_ (.B(\TRNG.hash[6] ),
    .C(_07001_),
    .A(net5573),
    .Y(_07006_));
 sg13g2_xor2_1 _15374_ (.B(_07006_),
    .A(\TRNG.hash[7] ),
    .X(_07007_));
 sg13g2_o21ai_1 _15375_ (.B1(_07005_),
    .Y(_00493_),
    .A1(_06877_),
    .A2(_07007_));
 sg13g2_nand3_1 _15376_ (.B(\TRNG.hash[6] ),
    .C(_07001_),
    .A(\TRNG.hash[7] ),
    .Y(_07008_));
 sg13g2_inv_1 _15377_ (.Y(_07009_),
    .A(_07008_));
 sg13g2_nand2_1 _15378_ (.Y(_07010_),
    .A(net3628),
    .B(_07008_));
 sg13g2_xnor2_1 _15379_ (.Y(_07011_),
    .A(_00152_),
    .B(_07010_));
 sg13g2_nand2_1 _15380_ (.Y(_07012_),
    .A(net5188),
    .B(_07011_));
 sg13g2_a22oi_1 _15381_ (.Y(_07013_),
    .B1(net3620),
    .B2(net5351),
    .A2(net3560),
    .A1(net5855));
 sg13g2_a21oi_1 _15382_ (.A1(_07012_),
    .A2(_07013_),
    .Y(_00494_),
    .B1(net4965));
 sg13g2_o21ai_1 _15383_ (.B1(\TRNG.hash[9] ),
    .Y(_07014_),
    .A1(\TRNG.hash[8] ),
    .A2(_07009_));
 sg13g2_nand2b_1 _15384_ (.Y(_07015_),
    .B(_07014_),
    .A_N(\TRNG.hash[10] ));
 sg13g2_or2_2 _15385_ (.X(_07016_),
    .B(_07015_),
    .A(\TRNG.hash[11] ));
 sg13g2_xnor2_1 _15386_ (.Y(_07017_),
    .A(net3574),
    .B(_07016_));
 sg13g2_nand2_1 _15387_ (.Y(_07018_),
    .A(net5190),
    .B(_07017_));
 sg13g2_a22oi_1 _15388_ (.Y(_07019_),
    .B1(\TRNG.hash[12] ),
    .B2(net5355),
    .A2(net5869),
    .A1(\TRNG.hash[44] ));
 sg13g2_a21oi_1 _15389_ (.A1(_07018_),
    .A2(_07019_),
    .Y(_00495_),
    .B1(net4970));
 sg13g2_nand3_1 _15390_ (.B(\TRNG.hash[12] ),
    .C(_07016_),
    .A(\TRNG.hash[13] ),
    .Y(_07020_));
 sg13g2_a21o_1 _15391_ (.A2(_07016_),
    .A1(\TRNG.hash[12] ),
    .B1(net3704),
    .X(_07021_));
 sg13g2_nand3_1 _15392_ (.B(_07020_),
    .C(_07021_),
    .A(net5190),
    .Y(_07022_));
 sg13g2_a22oi_1 _15393_ (.Y(_07023_),
    .B1(net3704),
    .B2(net5355),
    .A2(net3683),
    .A1(net5868));
 sg13g2_a21oi_1 _15394_ (.A1(_07022_),
    .A2(_07023_),
    .Y(_00496_),
    .B1(net4970));
 sg13g2_nor2_1 _15395_ (.A(\TRNG.hash[15] ),
    .B(\TRNG.hash[14] ),
    .Y(_07024_));
 sg13g2_a21oi_1 _15396_ (.A1(_07020_),
    .A2(_07024_),
    .Y(_07025_),
    .B1(_04297_));
 sg13g2_nand3_1 _15397_ (.B(_07020_),
    .C(_07024_),
    .A(_04297_),
    .Y(_07026_));
 sg13g2_nand3b_1 _15398_ (.B(_07026_),
    .C(net5190),
    .Y(_07027_),
    .A_N(_07025_));
 sg13g2_a22oi_1 _15399_ (.Y(_07028_),
    .B1(net3536),
    .B2(net5351),
    .A2(net5855),
    .A1(net3526));
 sg13g2_a21oi_1 _15400_ (.A1(_07027_),
    .A2(_07028_),
    .Y(_00497_),
    .B1(net4965));
 sg13g2_and2_1 _15401_ (.A(\TRNG.hash[17] ),
    .B(_07025_),
    .X(_07029_));
 sg13g2_o21ai_1 _15402_ (.B1(net5190),
    .Y(_07030_),
    .A1(\TRNG.hash[17] ),
    .A2(_07025_));
 sg13g2_a22oi_1 _15403_ (.Y(_07031_),
    .B1(net3856),
    .B2(net5355),
    .A2(net5867),
    .A1(net3679));
 sg13g2_o21ai_1 _15404_ (.B1(_07031_),
    .Y(_07032_),
    .A1(_07029_),
    .A2(_07030_));
 sg13g2_and2_1 _15405_ (.A(net4976),
    .B(_07032_),
    .X(_00498_));
 sg13g2_and2_1 _15406_ (.A(\TRNG.hash[18] ),
    .B(_07029_),
    .X(_07033_));
 sg13g2_nor2_1 _15407_ (.A(net5179),
    .B(_07033_),
    .Y(_07034_));
 sg13g2_o21ai_1 _15408_ (.B1(_07034_),
    .Y(_07035_),
    .A1(\TRNG.hash[18] ),
    .A2(_07029_));
 sg13g2_a22oi_1 _15409_ (.Y(_07036_),
    .B1(\TRNG.hash[18] ),
    .B2(net5355),
    .A2(net3576),
    .A1(net5867));
 sg13g2_a21oi_1 _15410_ (.A1(_07035_),
    .A2(net3577),
    .Y(_00499_),
    .B1(net4970));
 sg13g2_and2_1 _15411_ (.A(\TRNG.hash[19] ),
    .B(_07033_),
    .X(_07037_));
 sg13g2_o21ai_1 _15412_ (.B1(net5190),
    .Y(_07038_),
    .A1(\TRNG.hash[19] ),
    .A2(_07033_));
 sg13g2_a22oi_1 _15413_ (.Y(_07039_),
    .B1(net3874),
    .B2(net5355),
    .A2(net3587),
    .A1(net5867));
 sg13g2_o21ai_1 _15414_ (.B1(_07039_),
    .Y(_07040_),
    .A1(_07037_),
    .A2(_07038_));
 sg13g2_and2_1 _15415_ (.A(net4976),
    .B(_07040_),
    .X(_00500_));
 sg13g2_and2_1 _15416_ (.A(\TRNG.hash[20] ),
    .B(_07037_),
    .X(_07041_));
 sg13g2_inv_1 _15417_ (.Y(_07042_),
    .A(_07041_));
 sg13g2_nor2_1 _15418_ (.A(net5179),
    .B(_07041_),
    .Y(_07043_));
 sg13g2_o21ai_1 _15419_ (.B1(_07043_),
    .Y(_07044_),
    .A1(net3612),
    .A2(_07037_));
 sg13g2_a22oi_1 _15420_ (.Y(_07045_),
    .B1(net3612),
    .B2(net5355),
    .A2(\TRNG.hash[52] ),
    .A1(net5860));
 sg13g2_a21oi_1 _15421_ (.A1(_07044_),
    .A2(net3613),
    .Y(_00501_),
    .B1(net4970));
 sg13g2_nor4_2 _15422_ (.A(\TRNG.hash[23] ),
    .B(\TRNG.hash[22] ),
    .C(\TRNG.hash[21] ),
    .Y(_07046_),
    .D(_07041_));
 sg13g2_nor2b_1 _15423_ (.A(\TRNG.hash[24] ),
    .B_N(_07046_),
    .Y(_07047_));
 sg13g2_nor2b_1 _15424_ (.A(\TRNG.hash[25] ),
    .B_N(_07047_),
    .Y(_07048_));
 sg13g2_nor2b_2 _15425_ (.A(_07048_),
    .B_N(\TRNG.hash[26] ),
    .Y(_07049_));
 sg13g2_nand2b_1 _15426_ (.Y(_07050_),
    .B(_07048_),
    .A_N(net3761));
 sg13g2_nand3b_1 _15427_ (.B(_07050_),
    .C(net5191),
    .Y(_07051_),
    .A_N(_07049_));
 sg13g2_a22oi_1 _15428_ (.Y(_07052_),
    .B1(net3761),
    .B2(net5356),
    .A2(net5870),
    .A1(\TRNG.hash[58] ));
 sg13g2_a21oi_1 _15429_ (.A1(_07051_),
    .A2(net3762),
    .Y(_00502_),
    .B1(net4971));
 sg13g2_nor3_1 _15430_ (.A(\TRNG.hash[28] ),
    .B(\TRNG.hash[27] ),
    .C(_07049_),
    .Y(_07053_));
 sg13g2_nand2b_1 _15431_ (.Y(_07054_),
    .B(\TRNG.hash[29] ),
    .A_N(_07053_));
 sg13g2_nand2b_1 _15432_ (.Y(_07055_),
    .B(_07053_),
    .A_N(\TRNG.hash[29] ));
 sg13g2_nand3_1 _15433_ (.B(_07054_),
    .C(_07055_),
    .A(net5191),
    .Y(_07056_));
 sg13g2_a22oi_1 _15434_ (.Y(_07057_),
    .B1(\TRNG.hash[29] ),
    .B2(net5356),
    .A2(net3598),
    .A1(net5870));
 sg13g2_a21oi_1 _15435_ (.A1(_07056_),
    .A2(net3599),
    .Y(_00503_),
    .B1(net4971));
 sg13g2_nand2b_1 _15436_ (.Y(_07058_),
    .B(_07054_),
    .A_N(\TRNG.hash[30] ));
 sg13g2_a21oi_1 _15437_ (.A1(\TRNG.hash[31] ),
    .A2(_07058_),
    .Y(_07059_),
    .B1(net5179));
 sg13g2_o21ai_1 _15438_ (.B1(_07059_),
    .Y(_07060_),
    .A1(net3753),
    .A2(_07058_));
 sg13g2_a22oi_1 _15439_ (.Y(_07061_),
    .B1(net3753),
    .B2(net5356),
    .A2(\TRNG.hash[63] ),
    .A1(net5870));
 sg13g2_a21oi_1 _15440_ (.A1(_07060_),
    .A2(net3754),
    .Y(_00504_),
    .B1(net4971));
 sg13g2_nor2_1 _15441_ (.A(\TRNG.hash[33] ),
    .B(\TRNG.hash[32] ),
    .Y(_07062_));
 sg13g2_xor2_1 _15442_ (.B(_07062_),
    .A(net3517),
    .X(_07063_));
 sg13g2_nand2_1 _15443_ (.Y(_07064_),
    .A(net5192),
    .B(_07063_));
 sg13g2_a22oi_1 _15444_ (.Y(_07065_),
    .B1(\TRNG.hash[34] ),
    .B2(net5350),
    .A2(net5847),
    .A1(\TRNG.hash[66] ));
 sg13g2_a21oi_1 _15445_ (.A1(_07064_),
    .A2(_07065_),
    .Y(_00505_),
    .B1(net4965));
 sg13g2_o21ai_1 _15446_ (.B1(\TRNG.hash[34] ),
    .Y(_07066_),
    .A1(\TRNG.hash[33] ),
    .A2(\TRNG.hash[32] ));
 sg13g2_o21ai_1 _15447_ (.B1(_00162_),
    .Y(_07067_),
    .A1(\TRNG.hash[35] ),
    .A2(_07066_));
 sg13g2_xnor2_1 _15448_ (.Y(_07068_),
    .A(net3500),
    .B(_07067_));
 sg13g2_nand2_1 _15449_ (.Y(_07069_),
    .A(net5188),
    .B(net3501));
 sg13g2_a22oi_1 _15450_ (.Y(_07070_),
    .B1(\TRNG.hash[36] ),
    .B2(net5350),
    .A2(\TRNG.hash[68] ),
    .A1(net5857));
 sg13g2_a21oi_1 _15451_ (.A1(_07069_),
    .A2(_07070_),
    .Y(_00506_),
    .B1(net4965));
 sg13g2_nand2_2 _15452_ (.Y(_07071_),
    .A(\TRNG.hash[36] ),
    .B(_07067_));
 sg13g2_o21ai_1 _15453_ (.B1(_00164_),
    .Y(_07072_),
    .A1(\TRNG.hash[37] ),
    .A2(_07071_));
 sg13g2_xnor2_1 _15454_ (.Y(_07073_),
    .A(net3489),
    .B(_07072_));
 sg13g2_nand2_1 _15455_ (.Y(_07074_),
    .A(net5187),
    .B(net3490));
 sg13g2_a22oi_1 _15456_ (.Y(_07075_),
    .B1(\TRNG.hash[38] ),
    .B2(net5350),
    .A2(\TRNG.hash[70] ),
    .A1(net5848));
 sg13g2_a21oi_1 _15457_ (.A1(_07074_),
    .A2(_07075_),
    .Y(_00507_),
    .B1(net4967));
 sg13g2_nand2b_1 _15458_ (.Y(_07076_),
    .B(_07071_),
    .A_N(\TRNG.hash[37] ));
 sg13g2_a21o_1 _15459_ (.A2(_07076_),
    .A1(\TRNG.hash[38] ),
    .B1(\TRNG.hash[39] ),
    .X(_07077_));
 sg13g2_o21ai_1 _15460_ (.B1(\TRNG.hash[41] ),
    .Y(_07078_),
    .A1(\TRNG.hash[40] ),
    .A2(_07077_));
 sg13g2_or3_1 _15461_ (.A(\TRNG.hash[40] ),
    .B(\TRNG.hash[41] ),
    .C(_07077_),
    .X(_07079_));
 sg13g2_nand3_1 _15462_ (.B(_07078_),
    .C(_07079_),
    .A(net5192),
    .Y(_07080_));
 sg13g2_a22oi_1 _15463_ (.Y(_07081_),
    .B1(net3560),
    .B2(net5351),
    .A2(\TRNG.hash[73] ),
    .A1(net5855));
 sg13g2_a21oi_1 _15464_ (.A1(_07080_),
    .A2(net3561),
    .Y(_00508_),
    .B1(net4965));
 sg13g2_a21oi_1 _15465_ (.A1(net3412),
    .A2(_07078_),
    .Y(_07082_),
    .B1(net5180));
 sg13g2_o21ai_1 _15466_ (.B1(_07082_),
    .Y(_07083_),
    .A1(net3412),
    .A2(_07078_));
 sg13g2_a22oi_1 _15467_ (.Y(_07084_),
    .B1(\TRNG.hash[42] ),
    .B2(net5351),
    .A2(\TRNG.hash[74] ),
    .A1(net5854));
 sg13g2_a21oi_1 _15468_ (.A1(_07083_),
    .A2(_07084_),
    .Y(_00509_),
    .B1(net4965));
 sg13g2_nor2_1 _15469_ (.A(_04296_),
    .B(_07078_),
    .Y(_07085_));
 sg13g2_nor2_1 _15470_ (.A(\TRNG.hash[43] ),
    .B(_07085_),
    .Y(_07086_));
 sg13g2_inv_1 _15471_ (.Y(_07087_),
    .A(_07086_));
 sg13g2_nand2_1 _15472_ (.Y(_07088_),
    .A(_00167_),
    .B(_07086_));
 sg13g2_xnor2_1 _15473_ (.Y(_07089_),
    .A(net3486),
    .B(_07088_));
 sg13g2_nand2_1 _15474_ (.Y(_07090_),
    .A(net5188),
    .B(net3487));
 sg13g2_a22oi_1 _15475_ (.Y(_07091_),
    .B1(\TRNG.hash[45] ),
    .B2(net5351),
    .A2(net5854),
    .A1(net3447));
 sg13g2_a21oi_1 _15476_ (.A1(_07090_),
    .A2(_07091_),
    .Y(_00510_),
    .B1(net4966));
 sg13g2_o21ai_1 _15477_ (.B1(\TRNG.hash[45] ),
    .Y(_07092_),
    .A1(\TRNG.hash[44] ),
    .A2(_07087_));
 sg13g2_nand2b_1 _15478_ (.Y(_07093_),
    .B(_07092_),
    .A_N(\TRNG.hash[46] ));
 sg13g2_nor2_2 _15479_ (.A(\TRNG.hash[47] ),
    .B(_07093_),
    .Y(_07094_));
 sg13g2_or4_2 _15480_ (.A(\TRNG.hash[49] ),
    .B(\TRNG.hash[48] ),
    .C(\TRNG.hash[47] ),
    .D(_07093_),
    .X(_07095_));
 sg13g2_xnor2_1 _15481_ (.Y(_07096_),
    .A(net3480),
    .B(_07095_));
 sg13g2_nand2_1 _15482_ (.Y(_07097_),
    .A(net5190),
    .B(_07096_));
 sg13g2_a22oi_1 _15483_ (.Y(_07098_),
    .B1(\TRNG.hash[50] ),
    .B2(net5355),
    .A2(net5860),
    .A1(\TRNG.hash[82] ));
 sg13g2_a21oi_1 _15484_ (.A1(_07097_),
    .A2(_07098_),
    .Y(_00511_),
    .B1(net4970));
 sg13g2_and3_2 _15485_ (.X(_07099_),
    .A(\TRNG.hash[51] ),
    .B(\TRNG.hash[50] ),
    .C(_07095_));
 sg13g2_a21oi_1 _15486_ (.A1(net3576),
    .A2(_07095_),
    .Y(_07100_),
    .B1(net3587));
 sg13g2_nor3_1 _15487_ (.A(net5180),
    .B(_07099_),
    .C(_07100_),
    .Y(_07101_));
 sg13g2_a221oi_1 _15488_ (.B2(net5355),
    .C1(_07101_),
    .B1(net3587),
    .A1(net5860),
    .Y(_07102_),
    .A2(\TRNG.hash[83] ));
 sg13g2_nor2_1 _15489_ (.A(net4970),
    .B(net3588),
    .Y(_00512_));
 sg13g2_xnor2_1 _15490_ (.Y(_07103_),
    .A(net3549),
    .B(_07099_));
 sg13g2_nand2_1 _15491_ (.Y(_07104_),
    .A(net5189),
    .B(_07103_));
 sg13g2_a22oi_1 _15492_ (.Y(_07105_),
    .B1(\TRNG.hash[52] ),
    .B2(net5353),
    .A2(\TRNG.hash[84] ),
    .A1(net5860));
 sg13g2_a21oi_1 _15493_ (.A1(_07104_),
    .A2(_07105_),
    .Y(_00513_),
    .B1(net4968));
 sg13g2_nand3_1 _15494_ (.B(\TRNG.hash[52] ),
    .C(_07099_),
    .A(net3939),
    .Y(_07106_));
 sg13g2_a21o_1 _15495_ (.A2(_07099_),
    .A1(\TRNG.hash[52] ),
    .B1(net3571),
    .X(_07107_));
 sg13g2_nand3_1 _15496_ (.B(_07106_),
    .C(_07107_),
    .A(net5189),
    .Y(_07108_));
 sg13g2_a22oi_1 _15497_ (.Y(_07109_),
    .B1(net3571),
    .B2(net5353),
    .A2(\TRNG.hash[85] ),
    .A1(net5859));
 sg13g2_a21oi_1 _15498_ (.A1(_07108_),
    .A2(net3572),
    .Y(_00514_),
    .B1(net4968));
 sg13g2_or2_1 _15499_ (.X(_07110_),
    .B(_07106_),
    .A(_04295_));
 sg13g2_a21oi_1 _15500_ (.A1(_04295_),
    .A2(_07106_),
    .Y(_07111_),
    .B1(net5179));
 sg13g2_nand2_1 _15501_ (.Y(_07112_),
    .A(_07110_),
    .B(_07111_));
 sg13g2_a22oi_1 _15502_ (.Y(_07113_),
    .B1(net3558),
    .B2(net5353),
    .A2(\TRNG.hash[86] ),
    .A1(net5859));
 sg13g2_a21oi_1 _15503_ (.A1(_07112_),
    .A2(net3559),
    .Y(_00515_),
    .B1(net4968));
 sg13g2_o21ai_1 _15504_ (.B1(_00172_),
    .Y(_07114_),
    .A1(\TRNG.hash[55] ),
    .A2(_07110_));
 sg13g2_nor3_2 _15505_ (.A(\TRNG.hash[57] ),
    .B(\TRNG.hash[56] ),
    .C(_07114_),
    .Y(_07115_));
 sg13g2_nor2b_1 _15506_ (.A(\TRNG.hash[58] ),
    .B_N(_07115_),
    .Y(_07116_));
 sg13g2_nor2b_1 _15507_ (.A(\TRNG.hash[59] ),
    .B_N(_07116_),
    .Y(_07117_));
 sg13g2_nand2_1 _15508_ (.Y(_07118_),
    .A(_00171_),
    .B(_07117_));
 sg13g2_xnor2_1 _15509_ (.Y(_07119_),
    .A(net3469),
    .B(_07118_));
 sg13g2_nand2_1 _15510_ (.Y(_07120_),
    .A(net5189),
    .B(net3470));
 sg13g2_a22oi_1 _15511_ (.Y(_07121_),
    .B1(\TRNG.hash[61] ),
    .B2(net5354),
    .A2(\TRNG.hash[93] ),
    .A1(net5865));
 sg13g2_a21oi_1 _15512_ (.A1(_07120_),
    .A2(_07121_),
    .Y(_00516_),
    .B1(net4969));
 sg13g2_nor2b_1 _15513_ (.A(\TRNG.hash[60] ),
    .B_N(_07117_),
    .Y(_07122_));
 sg13g2_nor2b_1 _15514_ (.A(_07122_),
    .B_N(\TRNG.hash[61] ),
    .Y(_07123_));
 sg13g2_nand2_1 _15515_ (.Y(_07124_),
    .A(\TRNG.hash[62] ),
    .B(_07123_));
 sg13g2_o21ai_1 _15516_ (.B1(net5189),
    .Y(_07125_),
    .A1(\TRNG.hash[62] ),
    .A2(_07123_));
 sg13g2_nand2b_1 _15517_ (.Y(_07126_),
    .B(_07124_),
    .A_N(_07125_));
 sg13g2_a22oi_1 _15518_ (.Y(_07127_),
    .B1(net3722),
    .B2(net5356),
    .A2(\TRNG.hash[94] ),
    .A1(net5864));
 sg13g2_a21oi_1 _15519_ (.A1(_07126_),
    .A2(net3723),
    .Y(_00517_),
    .B1(net4968));
 sg13g2_xnor2_1 _15520_ (.Y(_07128_),
    .A(\TRNG.hash[63] ),
    .B(_07124_));
 sg13g2_nand2_1 _15521_ (.Y(_07129_),
    .A(net5191),
    .B(_07128_));
 sg13g2_a22oi_1 _15522_ (.Y(_07130_),
    .B1(\TRNG.hash[63] ),
    .B2(net5356),
    .A2(net5864),
    .A1(net3724));
 sg13g2_a21oi_1 _15523_ (.A1(_07129_),
    .A2(net3725),
    .Y(_00518_),
    .B1(net4971));
 sg13g2_or2_2 _15524_ (.X(_07131_),
    .B(\TRNG.hash[66] ),
    .A(\TRNG.hash[67] ));
 sg13g2_xnor2_1 _15525_ (.Y(_07132_),
    .A(net3457),
    .B(_07131_));
 sg13g2_nand2_1 _15526_ (.Y(_07133_),
    .A(net5188),
    .B(_07132_));
 sg13g2_a22oi_1 _15527_ (.Y(_07134_),
    .B1(\TRNG.hash[68] ),
    .B2(net5350),
    .A2(net5857),
    .A1(net5551));
 sg13g2_a21oi_1 _15528_ (.A1(_07133_),
    .A2(_07134_),
    .Y(_00519_),
    .B1(net4965));
 sg13g2_nand2_1 _15529_ (.Y(_07135_),
    .A(net5550),
    .B(net4745));
 sg13g2_nand3_1 _15530_ (.B(\TRNG.hash[68] ),
    .C(_07131_),
    .A(net5573),
    .Y(_07136_));
 sg13g2_nand4_1 _15531_ (.B(\TRNG.hash[69] ),
    .C(\TRNG.hash[68] ),
    .A(net5573),
    .Y(_07137_),
    .D(_07131_));
 sg13g2_xor2_1 _15532_ (.B(_07136_),
    .A(net3841),
    .X(_07138_));
 sg13g2_o21ai_1 _15533_ (.B1(_07135_),
    .Y(_00520_),
    .A1(net4748),
    .A2(_07138_));
 sg13g2_nand2_1 _15534_ (.Y(_07139_),
    .A(net5549),
    .B(net4745));
 sg13g2_nand4_1 _15535_ (.B(\TRNG.hash[69] ),
    .C(\TRNG.hash[68] ),
    .A(\TRNG.hash[70] ),
    .Y(_07140_),
    .D(_07131_));
 sg13g2_xor2_1 _15536_ (.B(_07137_),
    .A(net3824),
    .X(_07141_));
 sg13g2_o21ai_1 _15537_ (.B1(_07139_),
    .Y(_00521_),
    .A1(net4748),
    .A2(_07141_));
 sg13g2_o21ai_1 _15538_ (.B1(_00180_),
    .Y(_07142_),
    .A1(\TRNG.hash[71] ),
    .A2(_07140_));
 sg13g2_xnor2_1 _15539_ (.Y(_07143_),
    .A(net3492),
    .B(_07142_));
 sg13g2_nand2_1 _15540_ (.Y(_07144_),
    .A(net5186),
    .B(net3493));
 sg13g2_a22oi_1 _15541_ (.Y(_07145_),
    .B1(\TRNG.hash[72] ),
    .B2(net5352),
    .A2(net5896),
    .A1(net5851));
 sg13g2_a21oi_1 _15542_ (.A1(_07144_),
    .A2(_07145_),
    .Y(_00522_),
    .B1(net4967));
 sg13g2_a21o_1 _15543_ (.A2(_07142_),
    .A1(\TRNG.hash[72] ),
    .B1(\TRNG.hash[73] ),
    .X(_07146_));
 sg13g2_nand2_1 _15544_ (.Y(_07147_),
    .A(\TRNG.hash[73] ),
    .B(\TRNG.hash[72] ));
 sg13g2_nand2b_1 _15545_ (.Y(_07148_),
    .B(_07142_),
    .A_N(_07147_));
 sg13g2_nand3_1 _15546_ (.B(_07146_),
    .C(_07148_),
    .A(net5188),
    .Y(_07149_));
 sg13g2_a22oi_1 _15547_ (.Y(_07150_),
    .B1(net3809),
    .B2(net5352),
    .A2(net5851),
    .A1(\TRNG.hash[105] ));
 sg13g2_a21oi_1 _15548_ (.A1(_07149_),
    .A2(_07150_),
    .Y(_00523_),
    .B1(net4967));
 sg13g2_a21oi_1 _15549_ (.A1(_04220_),
    .A2(_07140_),
    .Y(_07151_),
    .B1(_07147_));
 sg13g2_nand2_1 _15550_ (.Y(_07152_),
    .A(net5573),
    .B(_07151_));
 sg13g2_xor2_1 _15551_ (.B(_07152_),
    .A(net3738),
    .X(_07153_));
 sg13g2_nand2_1 _15552_ (.Y(_07154_),
    .A(net5895),
    .B(net4745));
 sg13g2_o21ai_1 _15553_ (.B1(_07154_),
    .Y(_00524_),
    .A1(net4748),
    .A2(_07153_));
 sg13g2_nand2_1 _15554_ (.Y(_07155_),
    .A(\TRNG.hash[74] ),
    .B(_07151_));
 sg13g2_o21ai_1 _15555_ (.B1(_00182_),
    .Y(_07156_),
    .A1(\TRNG.hash[75] ),
    .A2(_07155_));
 sg13g2_xnor2_1 _15556_ (.Y(_07157_),
    .A(net3419),
    .B(_07156_));
 sg13g2_nand2_1 _15557_ (.Y(_07158_),
    .A(net5188),
    .B(_07157_));
 sg13g2_a22oi_1 _15558_ (.Y(_07159_),
    .B1(\TRNG.hash[76] ),
    .B2(net5351),
    .A2(net5854),
    .A1(net5548));
 sg13g2_a21oi_1 _15559_ (.A1(_07158_),
    .A2(_07159_),
    .Y(_00525_),
    .B1(net4966));
 sg13g2_nand2b_1 _15560_ (.Y(_07160_),
    .B(_07155_),
    .A_N(\TRNG.hash[75] ));
 sg13g2_a21oi_1 _15561_ (.A1(\TRNG.hash[76] ),
    .A2(_07160_),
    .Y(_07161_),
    .B1(\TRNG.hash[77] ));
 sg13g2_inv_1 _15562_ (.Y(_07162_),
    .A(_07161_));
 sg13g2_nand2_1 _15563_ (.Y(_07163_),
    .A(net3415),
    .B(_07161_));
 sg13g2_xnor2_1 _15564_ (.Y(_07164_),
    .A(_00183_),
    .B(_07163_));
 sg13g2_nand2_1 _15565_ (.Y(_07165_),
    .A(net5186),
    .B(net3416));
 sg13g2_a22oi_1 _15566_ (.Y(_07166_),
    .B1(\TRNG.hash[79] ),
    .B2(net5352),
    .A2(net5892),
    .A1(net5851));
 sg13g2_a21oi_1 _15567_ (.A1(_07165_),
    .A2(_07166_),
    .Y(_00526_),
    .B1(net4967));
 sg13g2_o21ai_1 _15568_ (.B1(\TRNG.hash[79] ),
    .Y(_07167_),
    .A1(\TRNG.hash[78] ),
    .A2(_07162_));
 sg13g2_nand2_1 _15569_ (.Y(_07168_),
    .A(net3601),
    .B(_07167_));
 sg13g2_a21oi_1 _15570_ (.A1(\TRNG.hash[81] ),
    .A2(_07168_),
    .Y(_07169_),
    .B1(net5180));
 sg13g2_o21ai_1 _15571_ (.B1(_07169_),
    .Y(_07170_),
    .A1(\TRNG.hash[81] ),
    .A2(_07168_));
 sg13g2_a22oi_1 _15572_ (.Y(_07171_),
    .B1(\TRNG.hash[81] ),
    .B2(net5351),
    .A2(net5852),
    .A1(net5546));
 sg13g2_a21oi_1 _15573_ (.A1(net3602),
    .A2(_07171_),
    .Y(_00527_),
    .B1(net4966));
 sg13g2_nand2b_1 _15574_ (.Y(_07172_),
    .B(_07167_),
    .A_N(\TRNG.hash[80] ));
 sg13g2_and2_2 _15575_ (.A(\TRNG.hash[81] ),
    .B(_07172_),
    .X(_07173_));
 sg13g2_nor2_1 _15576_ (.A(\TRNG.hash[82] ),
    .B(_07173_),
    .Y(_07174_));
 sg13g2_nor2b_1 _15577_ (.A(_07174_),
    .B_N(\TRNG.hash[83] ),
    .Y(_07175_));
 sg13g2_o21ai_1 _15578_ (.B1(\TRNG.hash[83] ),
    .Y(_07176_),
    .A1(\TRNG.hash[82] ),
    .A2(_07173_));
 sg13g2_nor3_1 _15579_ (.A(\TRNG.hash[82] ),
    .B(\TRNG.hash[83] ),
    .C(_07173_),
    .Y(_07177_));
 sg13g2_nor3_1 _15580_ (.A(net5179),
    .B(_07175_),
    .C(_07177_),
    .Y(_07178_));
 sg13g2_a221oi_1 _15581_ (.B2(net5353),
    .C1(_07178_),
    .B1(net3717),
    .A1(net5544),
    .Y(_07179_),
    .A2(net5860));
 sg13g2_nor2_1 _15582_ (.A(net4968),
    .B(_07179_),
    .Y(_00528_));
 sg13g2_a21oi_1 _15583_ (.A1(net3382),
    .A2(_07176_),
    .Y(_07180_),
    .B1(net5179));
 sg13g2_o21ai_1 _15584_ (.B1(_07180_),
    .Y(_07181_),
    .A1(net3382),
    .A2(_07176_));
 sg13g2_a22oi_1 _15585_ (.Y(_07182_),
    .B1(\TRNG.hash[84] ),
    .B2(net5353),
    .A2(\TRNG.hash[116] ),
    .A1(net5859));
 sg13g2_a21oi_1 _15586_ (.A1(_07181_),
    .A2(_07182_),
    .Y(_00529_),
    .B1(net4968));
 sg13g2_and3_2 _15587_ (.X(_07183_),
    .A(\TRNG.hash[85] ),
    .B(\TRNG.hash[84] ),
    .C(_07175_));
 sg13g2_a21oi_1 _15588_ (.A1(\TRNG.hash[84] ),
    .A2(_07175_),
    .Y(_07184_),
    .B1(net3581));
 sg13g2_nor3_1 _15589_ (.A(net5179),
    .B(_07183_),
    .C(_07184_),
    .Y(_07185_));
 sg13g2_a221oi_1 _15590_ (.B2(net5353),
    .C1(_07185_),
    .B1(net3581),
    .A1(net5860),
    .Y(_07186_),
    .A2(net5889));
 sg13g2_nor2_1 _15591_ (.A(net4968),
    .B(net3582),
    .Y(_00530_));
 sg13g2_xnor2_1 _15592_ (.Y(_07187_),
    .A(net3408),
    .B(_07183_));
 sg13g2_nand2_1 _15593_ (.Y(_07188_),
    .A(net5191),
    .B(_07187_));
 sg13g2_a22oi_1 _15594_ (.Y(_07189_),
    .B1(\TRNG.hash[86] ),
    .B2(net5354),
    .A2(\TRNG.hash[118] ),
    .A1(net5859));
 sg13g2_a21oi_1 _15595_ (.A1(_07188_),
    .A2(_07189_),
    .Y(_00531_),
    .B1(net4969));
 sg13g2_nand3_1 _15596_ (.B(\TRNG.hash[86] ),
    .C(_07183_),
    .A(\TRNG.hash[87] ),
    .Y(_07190_));
 sg13g2_a21o_1 _15597_ (.A2(_07183_),
    .A1(\TRNG.hash[86] ),
    .B1(net3608),
    .X(_07191_));
 sg13g2_nand3_1 _15598_ (.B(_07190_),
    .C(_07191_),
    .A(net5191),
    .Y(_07192_));
 sg13g2_a22oi_1 _15599_ (.Y(_07193_),
    .B1(net3608),
    .B2(net5353),
    .A2(\TRNG.hash[119] ),
    .A1(net5859));
 sg13g2_a21oi_1 _15600_ (.A1(_07192_),
    .A2(_07193_),
    .Y(_00532_),
    .B1(net4969));
 sg13g2_nor2_1 _15601_ (.A(\TRNG.hash[89] ),
    .B(\TRNG.hash[88] ),
    .Y(_07194_));
 sg13g2_nand2_1 _15602_ (.Y(_07195_),
    .A(_07190_),
    .B(_07194_));
 sg13g2_xnor2_1 _15603_ (.Y(_07196_),
    .A(net3472),
    .B(_07195_));
 sg13g2_nand2_1 _15604_ (.Y(_07197_),
    .A(net5189),
    .B(_07196_));
 sg13g2_a22oi_1 _15605_ (.Y(_07198_),
    .B1(\TRNG.hash[90] ),
    .B2(net5354),
    .A2(\TRNG.hash[122] ),
    .A1(net5862));
 sg13g2_a21oi_1 _15606_ (.A1(_07197_),
    .A2(_07198_),
    .Y(_00533_),
    .B1(net4969));
 sg13g2_nand2_1 _15607_ (.Y(_07199_),
    .A(\TRNG.hash[90] ),
    .B(_07195_));
 sg13g2_o21ai_1 _15608_ (.B1(_00190_),
    .Y(_07200_),
    .A1(\TRNG.hash[91] ),
    .A2(_07199_));
 sg13g2_nor2_1 _15609_ (.A(\TRNG.hash[92] ),
    .B(_07200_),
    .Y(_07201_));
 sg13g2_a21oi_1 _15610_ (.A1(net3463),
    .A2(_07201_),
    .Y(_07202_),
    .B1(net5179));
 sg13g2_o21ai_1 _15611_ (.B1(_07202_),
    .Y(_07203_),
    .A1(net3463),
    .A2(_07201_));
 sg13g2_a22oi_1 _15612_ (.Y(_07204_),
    .B1(\TRNG.hash[93] ),
    .B2(net5354),
    .A2(\TRNG.hash[125] ),
    .A1(net5861));
 sg13g2_a21oi_1 _15613_ (.A1(_07203_),
    .A2(_07204_),
    .Y(_00534_),
    .B1(net4969));
 sg13g2_nor2_1 _15614_ (.A(\TRNG.hash[92] ),
    .B(\TRNG.hash[91] ),
    .Y(_07205_));
 sg13g2_a21oi_1 _15615_ (.A1(_07199_),
    .A2(_07205_),
    .Y(_07206_),
    .B1(_04294_));
 sg13g2_nand2_1 _15616_ (.Y(_07207_),
    .A(\TRNG.hash[94] ),
    .B(_07206_));
 sg13g2_o21ai_1 _15617_ (.B1(net5189),
    .Y(_07208_),
    .A1(\TRNG.hash[94] ),
    .A2(_07206_));
 sg13g2_nand2b_1 _15618_ (.Y(_07209_),
    .B(_07207_),
    .A_N(_07208_));
 sg13g2_a22oi_1 _15619_ (.Y(_07210_),
    .B1(net3837),
    .B2(net5353),
    .A2(net5863),
    .A1(\TRNG.hash[126] ));
 sg13g2_a21oi_1 _15620_ (.A1(_07209_),
    .A2(_07210_),
    .Y(_00535_),
    .B1(net4969));
 sg13g2_nand2_1 _15621_ (.Y(_07211_),
    .A(\TRNG.sha256.W[3] ),
    .B(\TRNG.sha256.K[3] ));
 sg13g2_xor2_1 _15622_ (.B(\TRNG.sha256.K[3] ),
    .A(\TRNG.sha256.W[3] ),
    .X(_07212_));
 sg13g2_xnor2_1 _15623_ (.Y(_07213_),
    .A(_00156_),
    .B(_07212_));
 sg13g2_nand2_1 _15624_ (.Y(_07214_),
    .A(\TRNG.sha256.W[2] ),
    .B(\TRNG.sha256.K[2] ));
 sg13g2_o21ai_1 _15625_ (.B1(\TRNG.hash[2] ),
    .Y(_07215_),
    .A1(\TRNG.sha256.W[2] ),
    .A2(\TRNG.sha256.K[2] ));
 sg13g2_nand2_1 _15626_ (.Y(_07216_),
    .A(_07214_),
    .B(_07215_));
 sg13g2_and2_1 _15627_ (.A(_07213_),
    .B(_07216_),
    .X(_07217_));
 sg13g2_xnor2_1 _15628_ (.Y(_07218_),
    .A(\TRNG.hash[105] ),
    .B(_00200_));
 sg13g2_xnor2_1 _15629_ (.Y(_07219_),
    .A(net5547),
    .B(_07218_));
 sg13g2_xnor2_1 _15630_ (.Y(_07220_),
    .A(_07213_),
    .B(_07216_));
 sg13g2_nor2_1 _15631_ (.A(_07219_),
    .B(_07220_),
    .Y(_07221_));
 sg13g2_xnor2_1 _15632_ (.Y(_07222_),
    .A(net5895),
    .B(_00199_));
 sg13g2_xnor2_1 _15633_ (.Y(_07223_),
    .A(net5892),
    .B(_07222_));
 sg13g2_nand2_1 _15634_ (.Y(_07224_),
    .A(\TRNG.sha256.W[4] ),
    .B(\TRNG.sha256.K[4] ));
 sg13g2_xor2_1 _15635_ (.B(\TRNG.sha256.K[4] ),
    .A(\TRNG.sha256.W[4] ),
    .X(_07225_));
 sg13g2_xnor2_1 _15636_ (.Y(_07226_),
    .A(_00150_),
    .B(_07225_));
 sg13g2_o21ai_1 _15637_ (.B1(\TRNG.hash[3] ),
    .Y(_07227_),
    .A1(\TRNG.sha256.W[3] ),
    .A2(\TRNG.sha256.K[3] ));
 sg13g2_nand2_1 _15638_ (.Y(_07228_),
    .A(_07211_),
    .B(_07227_));
 sg13g2_nand2_1 _15639_ (.Y(_07229_),
    .A(_07226_),
    .B(_07228_));
 sg13g2_nor2_1 _15640_ (.A(_07226_),
    .B(_07228_),
    .Y(_07230_));
 sg13g2_xor2_1 _15641_ (.B(_07228_),
    .A(_07226_),
    .X(_07231_));
 sg13g2_xnor2_1 _15642_ (.Y(_07232_),
    .A(_07223_),
    .B(_07231_));
 sg13g2_o21ai_1 _15643_ (.B1(_07232_),
    .Y(_07233_),
    .A1(_07217_),
    .A2(_07221_));
 sg13g2_nor3_1 _15644_ (.A(_07217_),
    .B(_07221_),
    .C(_07232_),
    .Y(_07234_));
 sg13g2_or3_1 _15645_ (.A(_07217_),
    .B(_07221_),
    .C(_07232_),
    .X(_07235_));
 sg13g2_nand2_1 _15646_ (.Y(_07236_),
    .A(_07233_),
    .B(_07235_));
 sg13g2_mux2_1 _15647_ (.A0(_00161_),
    .A1(_00178_),
    .S(net5551),
    .X(_07237_));
 sg13g2_o21ai_1 _15648_ (.B1(_07233_),
    .Y(_07238_),
    .A1(_07234_),
    .A2(_07237_));
 sg13g2_o21ai_1 _15649_ (.B1(_07229_),
    .Y(_07239_),
    .A1(_07223_),
    .A2(_07230_));
 sg13g2_nand2_1 _15650_ (.Y(_07240_),
    .A(\TRNG.sha256.W[5] ),
    .B(\TRNG.sha256.K[5] ));
 sg13g2_xor2_1 _15651_ (.B(\TRNG.sha256.K[5] ),
    .A(\TRNG.sha256.W[5] ),
    .X(_07241_));
 sg13g2_xnor2_1 _15652_ (.Y(_07242_),
    .A(_00149_),
    .B(_07241_));
 sg13g2_o21ai_1 _15653_ (.B1(\TRNG.hash[4] ),
    .Y(_07243_),
    .A1(\TRNG.sha256.W[4] ),
    .A2(\TRNG.sha256.K[4] ));
 sg13g2_nand2_1 _15654_ (.Y(_07244_),
    .A(_07224_),
    .B(_07243_));
 sg13g2_and2_1 _15655_ (.A(_07242_),
    .B(_07244_),
    .X(_07245_));
 sg13g2_xor2_1 _15656_ (.B(_07244_),
    .A(_07242_),
    .X(_07246_));
 sg13g2_xnor2_1 _15657_ (.Y(_07247_),
    .A(\TRNG.hash[112] ),
    .B(net5894));
 sg13g2_xnor2_1 _15658_ (.Y(_07248_),
    .A(\TRNG.hash[126] ),
    .B(_07247_));
 sg13g2_xnor2_1 _15659_ (.Y(_07249_),
    .A(_07246_),
    .B(_07248_));
 sg13g2_nand2b_1 _15660_ (.Y(_07250_),
    .B(_07239_),
    .A_N(_07249_));
 sg13g2_xnor2_1 _15661_ (.Y(_07251_),
    .A(_07239_),
    .B(_07249_));
 sg13g2_mux2_1 _15662_ (.A0(\TRNG.hash[37] ),
    .A1(\TRNG.hash[69] ),
    .S(net5550),
    .X(_07252_));
 sg13g2_nand2_1 _15663_ (.Y(_07253_),
    .A(_07251_),
    .B(_07252_));
 sg13g2_xor2_1 _15664_ (.B(_07252_),
    .A(_07251_),
    .X(_07254_));
 sg13g2_nand2_1 _15665_ (.Y(_07255_),
    .A(_07238_),
    .B(_07254_));
 sg13g2_or2_1 _15666_ (.X(_07256_),
    .B(_07254_),
    .A(_07238_));
 sg13g2_nand2_1 _15667_ (.Y(_07257_),
    .A(_07255_),
    .B(_07256_));
 sg13g2_and2_1 _15668_ (.A(\TRNG.sha256.W[1] ),
    .B(\TRNG.sha256.K[1] ),
    .X(_07258_));
 sg13g2_xor2_1 _15669_ (.B(\TRNG.sha256.K[1] ),
    .A(\TRNG.sha256.W[1] ),
    .X(_07259_));
 sg13g2_a21oi_1 _15670_ (.A1(\TRNG.hash[1] ),
    .A2(_07259_),
    .Y(_07260_),
    .B1(_07258_));
 sg13g2_xor2_1 _15671_ (.B(\TRNG.sha256.K[2] ),
    .A(\TRNG.sha256.W[2] ),
    .X(_07261_));
 sg13g2_xnor2_1 _15672_ (.Y(_07262_),
    .A(_00157_),
    .B(_07261_));
 sg13g2_nand2b_1 _15673_ (.Y(_07263_),
    .B(_07262_),
    .A_N(_07260_));
 sg13g2_xnor2_1 _15674_ (.Y(_07264_),
    .A(\TRNG.hash[104] ),
    .B(_00201_));
 sg13g2_xnor2_1 _15675_ (.Y(_07265_),
    .A(net5893),
    .B(_07264_));
 sg13g2_nor2b_1 _15676_ (.A(_07262_),
    .B_N(_07260_),
    .Y(_07266_));
 sg13g2_xnor2_1 _15677_ (.Y(_07267_),
    .A(_07260_),
    .B(_07262_));
 sg13g2_o21ai_1 _15678_ (.B1(_07263_),
    .Y(_07268_),
    .A1(_07265_),
    .A2(_07266_));
 sg13g2_xor2_1 _15679_ (.B(_07220_),
    .A(_07219_),
    .X(_07269_));
 sg13g2_xnor2_1 _15680_ (.Y(_07270_),
    .A(_07268_),
    .B(_07269_));
 sg13g2_mux2_1 _15681_ (.A0(\TRNG.hash[35] ),
    .A1(\TRNG.hash[67] ),
    .S(net5552),
    .X(_07271_));
 sg13g2_nor2b_1 _15682_ (.A(_07270_),
    .B_N(_07271_),
    .Y(_07272_));
 sg13g2_a21oi_2 _15683_ (.B1(_07272_),
    .Y(_07273_),
    .A2(_07269_),
    .A1(_07268_));
 sg13g2_xnor2_1 _15684_ (.Y(_07274_),
    .A(_07236_),
    .B(_07237_));
 sg13g2_nor2_1 _15685_ (.A(_07273_),
    .B(_07274_),
    .Y(_07275_));
 sg13g2_xnor2_1 _15686_ (.Y(_07276_),
    .A(_07273_),
    .B(_07274_));
 sg13g2_and2_1 _15687_ (.A(\TRNG.sha256.W[0] ),
    .B(\TRNG.sha256.K[0] ),
    .X(_07277_));
 sg13g2_xor2_1 _15688_ (.B(\TRNG.sha256.K[0] ),
    .A(\TRNG.sha256.W[0] ),
    .X(_07278_));
 sg13g2_a21oi_1 _15689_ (.A1(\TRNG.hash[0] ),
    .A2(_07278_),
    .Y(_07279_),
    .B1(_07277_));
 sg13g2_xnor2_1 _15690_ (.Y(_07280_),
    .A(\TRNG.hash[1] ),
    .B(_07259_));
 sg13g2_nor2_1 _15691_ (.A(_07279_),
    .B(_07280_),
    .Y(_07281_));
 sg13g2_xor2_1 _15692_ (.B(_00202_),
    .A(net5897),
    .X(_07282_));
 sg13g2_xnor2_1 _15693_ (.Y(_07283_),
    .A(net5548),
    .B(_07282_));
 sg13g2_xor2_1 _15694_ (.B(_07280_),
    .A(_07279_),
    .X(_07284_));
 sg13g2_a21oi_1 _15695_ (.A1(_07283_),
    .A2(_07284_),
    .Y(_07285_),
    .B1(_07281_));
 sg13g2_xnor2_1 _15696_ (.Y(_07286_),
    .A(_07265_),
    .B(_07267_));
 sg13g2_nand2b_1 _15697_ (.Y(_07287_),
    .B(_07286_),
    .A_N(_07285_));
 sg13g2_xor2_1 _15698_ (.B(_07286_),
    .A(_07285_),
    .X(_07288_));
 sg13g2_mux2_1 _15699_ (.A0(_00160_),
    .A1(_00191_),
    .S(net5553),
    .X(_07289_));
 sg13g2_o21ai_1 _15700_ (.B1(_07287_),
    .Y(_07290_),
    .A1(_07288_),
    .A2(_07289_));
 sg13g2_xnor2_1 _15701_ (.Y(_07291_),
    .A(_07270_),
    .B(_07271_));
 sg13g2_nor2_1 _15702_ (.A(_07290_),
    .B(_07291_),
    .Y(_07292_));
 sg13g2_xnor2_1 _15703_ (.Y(_07293_),
    .A(\TRNG.hash[0] ),
    .B(_07278_));
 sg13g2_xnor2_1 _15704_ (.Y(_07294_),
    .A(net5894),
    .B(_00203_));
 sg13g2_xnor2_1 _15705_ (.Y(_07295_),
    .A(net5549),
    .B(_07294_));
 sg13g2_nor2_1 _15706_ (.A(_07293_),
    .B(_07295_),
    .Y(_07296_));
 sg13g2_xor2_1 _15707_ (.B(_07284_),
    .A(_07283_),
    .X(_07297_));
 sg13g2_and2_1 _15708_ (.A(_07296_),
    .B(_07297_),
    .X(_07298_));
 sg13g2_or2_1 _15709_ (.X(_07299_),
    .B(_07297_),
    .A(_07296_));
 sg13g2_xnor2_1 _15710_ (.Y(_07300_),
    .A(_07296_),
    .B(_07297_));
 sg13g2_mux2_1 _15711_ (.A0(\TRNG.hash[33] ),
    .A1(\TRNG.hash[65] ),
    .S(net5554),
    .X(_07301_));
 sg13g2_a21oi_1 _15712_ (.A1(_07299_),
    .A2(_07301_),
    .Y(_07302_),
    .B1(_07298_));
 sg13g2_xnor2_1 _15713_ (.Y(_07303_),
    .A(_07288_),
    .B(_07289_));
 sg13g2_nor2_1 _15714_ (.A(_07302_),
    .B(_07303_),
    .Y(_07304_));
 sg13g2_xnor2_1 _15715_ (.Y(_07305_),
    .A(_07300_),
    .B(_07301_));
 sg13g2_xnor2_1 _15716_ (.Y(_07306_),
    .A(_07293_),
    .B(_07295_));
 sg13g2_mux2_1 _15717_ (.A0(\TRNG.hash[32] ),
    .A1(\TRNG.hash[64] ),
    .S(net5555),
    .X(_07307_));
 sg13g2_nor2b_1 _15718_ (.A(_07306_),
    .B_N(_07307_),
    .Y(_07308_));
 sg13g2_and2_1 _15719_ (.A(_07305_),
    .B(_07308_),
    .X(_07309_));
 sg13g2_xor2_1 _15720_ (.B(_07303_),
    .A(_07302_),
    .X(_07310_));
 sg13g2_a21oi_1 _15721_ (.A1(_07309_),
    .A2(_07310_),
    .Y(_07311_),
    .B1(_07304_));
 sg13g2_a221oi_1 _15722_ (.B2(_07310_),
    .C1(_07304_),
    .B1(_07309_),
    .A1(_07290_),
    .Y(_07312_),
    .A2(_07291_));
 sg13g2_nor3_2 _15723_ (.A(_07276_),
    .B(_07292_),
    .C(_07312_),
    .Y(_07313_));
 sg13g2_nor2_1 _15724_ (.A(_07275_),
    .B(_07313_),
    .Y(_07314_));
 sg13g2_xnor2_1 _15725_ (.Y(_07315_),
    .A(_07257_),
    .B(_07314_));
 sg13g2_nand2b_1 _15726_ (.Y(_07316_),
    .B(\TRNG.hash[133] ),
    .A_N(_07315_));
 sg13g2_nor2b_1 _15727_ (.A(\TRNG.hash[133] ),
    .B_N(_07315_),
    .Y(_07317_));
 sg13g2_xnor2_1 _15728_ (.Y(_07318_),
    .A(\TRNG.hash[133] ),
    .B(_07315_));
 sg13g2_o21ai_1 _15729_ (.B1(_07276_),
    .Y(_07319_),
    .A1(_07292_),
    .A2(_07312_));
 sg13g2_nand2b_2 _15730_ (.Y(_07320_),
    .B(_07319_),
    .A_N(_07313_));
 sg13g2_nor2_1 _15731_ (.A(_04234_),
    .B(_07320_),
    .Y(_07321_));
 sg13g2_nand2_1 _15732_ (.Y(_07322_),
    .A(_04234_),
    .B(_07320_));
 sg13g2_nand2b_1 _15733_ (.Y(_07323_),
    .B(_07322_),
    .A_N(_07321_));
 sg13g2_xor2_1 _15734_ (.B(_07310_),
    .A(_07309_),
    .X(_07324_));
 sg13g2_and2_1 _15735_ (.A(\TRNG.hash[130] ),
    .B(_07324_),
    .X(_07325_));
 sg13g2_or2_1 _15736_ (.X(_07326_),
    .B(_07324_),
    .A(\TRNG.hash[130] ));
 sg13g2_nand2b_1 _15737_ (.Y(_07327_),
    .B(_07326_),
    .A_N(_07325_));
 sg13g2_xnor2_1 _15738_ (.Y(_07328_),
    .A(_07305_),
    .B(_07308_));
 sg13g2_or2_1 _15739_ (.X(_07329_),
    .B(_07328_),
    .A(_00146_));
 sg13g2_xnor2_1 _15740_ (.Y(_07330_),
    .A(_07306_),
    .B(_07307_));
 sg13g2_nand2_1 _15741_ (.Y(_07331_),
    .A(\TRNG.hash[128] ),
    .B(_07330_));
 sg13g2_and2_1 _15742_ (.A(_00146_),
    .B(_07328_),
    .X(_07332_));
 sg13g2_xor2_1 _15743_ (.B(_07328_),
    .A(_00146_),
    .X(_07333_));
 sg13g2_o21ai_1 _15744_ (.B1(_07329_),
    .Y(_07334_),
    .A1(_07331_),
    .A2(_07332_));
 sg13g2_a21oi_1 _15745_ (.A1(_07326_),
    .A2(_07334_),
    .Y(_07335_),
    .B1(_07325_));
 sg13g2_xnor2_1 _15746_ (.Y(_07336_),
    .A(_07290_),
    .B(_07291_));
 sg13g2_xor2_1 _15747_ (.B(_07336_),
    .A(_07311_),
    .X(_07337_));
 sg13g2_xnor2_1 _15748_ (.Y(_07338_),
    .A(\TRNG.hash[131] ),
    .B(_07337_));
 sg13g2_nor2_1 _15749_ (.A(_07335_),
    .B(_07338_),
    .Y(_07339_));
 sg13g2_nand2b_1 _15750_ (.Y(_07340_),
    .B(_07337_),
    .A_N(_00147_));
 sg13g2_o21ai_1 _15751_ (.B1(_07340_),
    .Y(_07341_),
    .A1(_07335_),
    .A2(_07338_));
 sg13g2_a21oi_1 _15752_ (.A1(_07322_),
    .A2(_07341_),
    .Y(_07342_),
    .B1(_07321_));
 sg13g2_o21ai_1 _15753_ (.B1(_07316_),
    .Y(_07343_),
    .A1(_07317_),
    .A2(_07342_));
 sg13g2_a21oi_2 _15754_ (.B1(_07245_),
    .Y(_07344_),
    .A2(_07248_),
    .A1(_07246_));
 sg13g2_xnor2_1 _15755_ (.Y(_07345_),
    .A(net5548),
    .B(_00198_));
 sg13g2_xnor2_1 _15756_ (.Y(_07346_),
    .A(net5546),
    .B(_07345_));
 sg13g2_nand2_1 _15757_ (.Y(_07347_),
    .A(\TRNG.sha256.W[6] ),
    .B(\TRNG.sha256.K[6] ));
 sg13g2_xor2_1 _15758_ (.B(\TRNG.sha256.K[6] ),
    .A(\TRNG.sha256.W[6] ),
    .X(_07348_));
 sg13g2_xnor2_1 _15759_ (.Y(_07349_),
    .A(_00151_),
    .B(_07348_));
 sg13g2_o21ai_1 _15760_ (.B1(\TRNG.hash[5] ),
    .Y(_07350_),
    .A1(\TRNG.sha256.W[5] ),
    .A2(\TRNG.sha256.K[5] ));
 sg13g2_nand2_1 _15761_ (.Y(_07351_),
    .A(_07240_),
    .B(_07350_));
 sg13g2_nand2_1 _15762_ (.Y(_07352_),
    .A(_07349_),
    .B(_07351_));
 sg13g2_nor2_1 _15763_ (.A(_07349_),
    .B(_07351_),
    .Y(_07353_));
 sg13g2_xor2_1 _15764_ (.B(_07351_),
    .A(_07349_),
    .X(_07354_));
 sg13g2_xnor2_1 _15765_ (.Y(_07355_),
    .A(_07346_),
    .B(_07354_));
 sg13g2_nor2b_1 _15766_ (.A(_07344_),
    .B_N(_07355_),
    .Y(_07356_));
 sg13g2_xnor2_1 _15767_ (.Y(_07357_),
    .A(_07344_),
    .B(_07355_));
 sg13g2_nor2_1 _15768_ (.A(net5549),
    .B(_00163_),
    .Y(_07358_));
 sg13g2_a21oi_2 _15769_ (.B1(_07358_),
    .Y(_07359_),
    .A2(_04378_),
    .A1(net5549));
 sg13g2_inv_1 _15770_ (.Y(_07360_),
    .A(_07359_));
 sg13g2_and2_1 _15771_ (.A(_07357_),
    .B(_07360_),
    .X(_07361_));
 sg13g2_xnor2_1 _15772_ (.Y(_07362_),
    .A(_07357_),
    .B(_07360_));
 sg13g2_a21oi_2 _15773_ (.B1(_07362_),
    .Y(_07363_),
    .A2(_07253_),
    .A1(_07250_));
 sg13g2_nand3_1 _15774_ (.B(_07253_),
    .C(_07362_),
    .A(_07250_),
    .Y(_07364_));
 sg13g2_nand2b_1 _15775_ (.Y(_07365_),
    .B(_07364_),
    .A_N(_07363_));
 sg13g2_o21ai_1 _15776_ (.B1(_07255_),
    .Y(_07366_),
    .A1(_07273_),
    .A2(_07274_));
 sg13g2_or4_2 _15777_ (.A(_07257_),
    .B(_07276_),
    .C(_07292_),
    .D(_07312_),
    .X(_07367_));
 sg13g2_o21ai_1 _15778_ (.B1(_07256_),
    .Y(_07368_),
    .A1(_07313_),
    .A2(_07366_));
 sg13g2_nor2_1 _15779_ (.A(_07365_),
    .B(_07368_),
    .Y(_07369_));
 sg13g2_xor2_1 _15780_ (.B(_07368_),
    .A(_07365_),
    .X(_07370_));
 sg13g2_xnor2_1 _15781_ (.Y(_07371_),
    .A(\TRNG.hash[134] ),
    .B(_07370_));
 sg13g2_inv_1 _15782_ (.Y(_07372_),
    .A(_07371_));
 sg13g2_a22oi_1 _15783_ (.Y(_07373_),
    .B1(_07372_),
    .B2(_07343_),
    .A2(_07370_),
    .A1(_04375_));
 sg13g2_o21ai_1 _15784_ (.B1(_07352_),
    .Y(_07374_),
    .A1(_07346_),
    .A2(_07353_));
 sg13g2_and2_1 _15785_ (.A(\TRNG.sha256.W[7] ),
    .B(\TRNG.sha256.K[7] ),
    .X(_07375_));
 sg13g2_xor2_1 _15786_ (.B(\TRNG.sha256.K[7] ),
    .A(\TRNG.sha256.W[7] ),
    .X(_07376_));
 sg13g2_xnor2_1 _15787_ (.Y(_07377_),
    .A(\TRNG.hash[7] ),
    .B(_07376_));
 sg13g2_o21ai_1 _15788_ (.B1(\TRNG.hash[6] ),
    .Y(_07378_),
    .A1(\TRNG.sha256.W[6] ),
    .A2(\TRNG.sha256.K[6] ));
 sg13g2_nand2_2 _15789_ (.Y(_07379_),
    .A(_07347_),
    .B(_07378_));
 sg13g2_nor2b_1 _15790_ (.A(_07377_),
    .B_N(_07379_),
    .Y(_07380_));
 sg13g2_nand2b_1 _15791_ (.Y(_07381_),
    .B(_07377_),
    .A_N(_07379_));
 sg13g2_xor2_1 _15792_ (.B(_07379_),
    .A(_07377_),
    .X(_07382_));
 sg13g2_xnor2_1 _15793_ (.Y(_07383_),
    .A(\TRNG.hash[96] ),
    .B(net5893));
 sg13g2_xnor2_1 _15794_ (.Y(_07384_),
    .A(net5545),
    .B(_07383_));
 sg13g2_xnor2_1 _15795_ (.Y(_07385_),
    .A(_07382_),
    .B(_07384_));
 sg13g2_nand2_1 _15796_ (.Y(_07386_),
    .A(_07374_),
    .B(_07385_));
 sg13g2_xnor2_1 _15797_ (.Y(_07387_),
    .A(_07374_),
    .B(_07385_));
 sg13g2_mux2_2 _15798_ (.A0(_00173_),
    .A1(_00180_),
    .S(net5897),
    .X(_07388_));
 sg13g2_xor2_1 _15799_ (.B(_07388_),
    .A(_07387_),
    .X(_07389_));
 sg13g2_o21ai_1 _15800_ (.B1(_07389_),
    .Y(_07390_),
    .A1(_07356_),
    .A2(_07361_));
 sg13g2_inv_1 _15801_ (.Y(_07391_),
    .A(_07390_));
 sg13g2_or3_1 _15802_ (.A(_07356_),
    .B(_07361_),
    .C(_07389_),
    .X(_07392_));
 sg13g2_nand2_1 _15803_ (.Y(_07393_),
    .A(_07390_),
    .B(_07392_));
 sg13g2_nor2_1 _15804_ (.A(_07363_),
    .B(_07369_),
    .Y(_07394_));
 sg13g2_xnor2_1 _15805_ (.Y(_07395_),
    .A(_07393_),
    .B(_07394_));
 sg13g2_or2_1 _15806_ (.X(_07396_),
    .B(_07395_),
    .A(_04300_));
 sg13g2_xnor2_1 _15807_ (.Y(_07397_),
    .A(_04300_),
    .B(_07395_));
 sg13g2_xnor2_1 _15808_ (.Y(_07398_),
    .A(_07373_),
    .B(_07397_));
 sg13g2_or2_1 _15809_ (.X(_07399_),
    .B(net5555),
    .A(net5554));
 sg13g2_nor2_1 _15810_ (.A(net5553),
    .B(_07399_),
    .Y(_07400_));
 sg13g2_nor3_1 _15811_ (.A(net5552),
    .B(net5553),
    .C(_07399_),
    .Y(_07401_));
 sg13g2_nor2b_1 _15812_ (.A(net5551),
    .B_N(_07401_),
    .Y(_07402_));
 sg13g2_nor2b_1 _15813_ (.A(net5550),
    .B_N(_07402_),
    .Y(_07403_));
 sg13g2_nor2b_1 _15814_ (.A(net5549),
    .B_N(_07403_),
    .Y(_07404_));
 sg13g2_nor2b_1 _15815_ (.A(_07404_),
    .B_N(net5897),
    .Y(_07405_));
 sg13g2_xor2_1 _15816_ (.B(_07404_),
    .A(net5897),
    .X(_07406_));
 sg13g2_o21ai_1 _15817_ (.B1(net4977),
    .Y(_07407_),
    .A1(net5897),
    .A2(net5177));
 sg13g2_a221oi_1 _15818_ (.B2(net5187),
    .C1(_07407_),
    .B1(_07406_),
    .A1(net5849),
    .Y(_00536_),
    .A2(_07398_));
 sg13g2_o21ai_1 _15819_ (.B1(_07396_),
    .Y(_07408_),
    .A1(_07373_),
    .A2(_07397_));
 sg13g2_a21oi_1 _15820_ (.A1(_07381_),
    .A2(_07384_),
    .Y(_07409_),
    .B1(_07380_));
 sg13g2_a21oi_2 _15821_ (.B1(_07375_),
    .Y(_07410_),
    .A2(_07376_),
    .A1(\TRNG.hash[7] ));
 sg13g2_and2_1 _15822_ (.A(\TRNG.sha256.W[8] ),
    .B(\TRNG.sha256.K[8] ),
    .X(_07411_));
 sg13g2_xor2_1 _15823_ (.B(\TRNG.sha256.K[8] ),
    .A(\TRNG.sha256.W[8] ),
    .X(_07412_));
 sg13g2_xnor2_1 _15824_ (.Y(_07413_),
    .A(\TRNG.hash[8] ),
    .B(_07412_));
 sg13g2_nor2_1 _15825_ (.A(_07410_),
    .B(_07413_),
    .Y(_07414_));
 sg13g2_xor2_1 _15826_ (.B(_07413_),
    .A(_07410_),
    .X(_07415_));
 sg13g2_xnor2_1 _15827_ (.Y(_07416_),
    .A(net5547),
    .B(net5554));
 sg13g2_xnor2_1 _15828_ (.Y(_07417_),
    .A(net5544),
    .B(_07416_));
 sg13g2_xnor2_1 _15829_ (.Y(_07418_),
    .A(_07415_),
    .B(_07417_));
 sg13g2_nor2_1 _15830_ (.A(_07409_),
    .B(_07418_),
    .Y(_07419_));
 sg13g2_xor2_1 _15831_ (.B(_07418_),
    .A(_07409_),
    .X(_07420_));
 sg13g2_mux2_1 _15832_ (.A0(_00174_),
    .A1(_00179_),
    .S(net5896),
    .X(_07421_));
 sg13g2_inv_1 _15833_ (.Y(_07422_),
    .A(_07421_));
 sg13g2_xnor2_1 _15834_ (.Y(_07423_),
    .A(_07420_),
    .B(_07421_));
 sg13g2_o21ai_1 _15835_ (.B1(_07386_),
    .Y(_07424_),
    .A1(_07387_),
    .A2(_07388_));
 sg13g2_nand2_1 _15836_ (.Y(_07425_),
    .A(_07423_),
    .B(_07424_));
 sg13g2_xnor2_1 _15837_ (.Y(_07426_),
    .A(_07423_),
    .B(_07424_));
 sg13g2_a21oi_1 _15838_ (.A1(_07363_),
    .A2(_07392_),
    .Y(_07427_),
    .B1(_07391_));
 sg13g2_or2_1 _15839_ (.X(_07428_),
    .B(_07393_),
    .A(_07365_));
 sg13g2_a221oi_1 _15840_ (.B2(_07363_),
    .C1(_07391_),
    .B1(_07392_),
    .A1(_07256_),
    .Y(_07429_),
    .A2(_07366_));
 sg13g2_a22oi_1 _15841_ (.Y(_07430_),
    .B1(_07429_),
    .B2(_07367_),
    .A2(_07428_),
    .A1(_07427_));
 sg13g2_nand2b_1 _15842_ (.Y(_07431_),
    .B(_07430_),
    .A_N(_07426_));
 sg13g2_xor2_1 _15843_ (.B(_07430_),
    .A(_07426_),
    .X(_07432_));
 sg13g2_xor2_1 _15844_ (.B(_07432_),
    .A(\TRNG.hash[136] ),
    .X(_07433_));
 sg13g2_inv_1 _15845_ (.Y(_07434_),
    .A(_07433_));
 sg13g2_xnor2_1 _15846_ (.Y(_07435_),
    .A(_07408_),
    .B(_07434_));
 sg13g2_nand2_1 _15847_ (.Y(_07436_),
    .A(net5896),
    .B(_07405_));
 sg13g2_xnor2_1 _15848_ (.Y(_07437_),
    .A(net5896),
    .B(_07405_));
 sg13g2_o21ai_1 _15849_ (.B1(net4977),
    .Y(_07438_),
    .A1(net5896),
    .A2(net5177));
 sg13g2_a221oi_1 _15850_ (.B2(net5187),
    .C1(_07438_),
    .B1(_07437_),
    .A1(net5846),
    .Y(_00537_),
    .A2(_07435_));
 sg13g2_a21o_1 _15851_ (.A2(_07422_),
    .A1(_07420_),
    .B1(_07419_),
    .X(_07439_));
 sg13g2_a21oi_2 _15852_ (.B1(_07414_),
    .Y(_07440_),
    .A2(_07417_),
    .A1(_07415_));
 sg13g2_a21oi_2 _15853_ (.B1(_07411_),
    .Y(_07441_),
    .A2(_07412_),
    .A1(\TRNG.hash[8] ));
 sg13g2_nand2_1 _15854_ (.Y(_07442_),
    .A(\TRNG.sha256.W[9] ),
    .B(\TRNG.sha256.K[9] ));
 sg13g2_xor2_1 _15855_ (.B(\TRNG.sha256.K[9] ),
    .A(\TRNG.sha256.W[9] ),
    .X(_07443_));
 sg13g2_xnor2_1 _15856_ (.Y(_07444_),
    .A(_00152_),
    .B(_07443_));
 sg13g2_nor2b_1 _15857_ (.A(_07441_),
    .B_N(_07444_),
    .Y(_07445_));
 sg13g2_xnor2_1 _15858_ (.Y(_07446_),
    .A(_07441_),
    .B(_07444_));
 sg13g2_xnor2_1 _15859_ (.Y(_07447_),
    .A(net5890),
    .B(net5892));
 sg13g2_xnor2_1 _15860_ (.Y(_07448_),
    .A(\TRNG.hash[98] ),
    .B(_07447_));
 sg13g2_xnor2_1 _15861_ (.Y(_07449_),
    .A(_07446_),
    .B(_07448_));
 sg13g2_nor2_1 _15862_ (.A(_07440_),
    .B(_07449_),
    .Y(_07450_));
 sg13g2_xor2_1 _15863_ (.B(_07449_),
    .A(_07440_),
    .X(_07451_));
 sg13g2_mux2_1 _15864_ (.A0(\TRNG.hash[41] ),
    .A1(\TRNG.hash[73] ),
    .S(\TRNG.hash[105] ),
    .X(_07452_));
 sg13g2_xor2_1 _15865_ (.B(_07452_),
    .A(_07451_),
    .X(_07453_));
 sg13g2_nor2_1 _15866_ (.A(_07439_),
    .B(_07453_),
    .Y(_07454_));
 sg13g2_nand2_1 _15867_ (.Y(_07455_),
    .A(_07439_),
    .B(_07453_));
 sg13g2_xnor2_1 _15868_ (.Y(_07456_),
    .A(_07439_),
    .B(_07453_));
 sg13g2_nand2_1 _15869_ (.Y(_07457_),
    .A(_07425_),
    .B(_07431_));
 sg13g2_xor2_1 _15870_ (.B(_07457_),
    .A(_07456_),
    .X(_07458_));
 sg13g2_nor2_1 _15871_ (.A(_04299_),
    .B(_07458_),
    .Y(_07459_));
 sg13g2_and2_1 _15872_ (.A(_04299_),
    .B(_07458_),
    .X(_07460_));
 sg13g2_nor2_1 _15873_ (.A(_00148_),
    .B(_07432_),
    .Y(_07461_));
 sg13g2_a21oi_1 _15874_ (.A1(_07408_),
    .A2(_07434_),
    .Y(_07462_),
    .B1(_07461_));
 sg13g2_or2_1 _15875_ (.X(_07463_),
    .B(_07461_),
    .A(_07459_));
 sg13g2_a21oi_1 _15876_ (.A1(_07408_),
    .A2(_07434_),
    .Y(_07464_),
    .B1(_07463_));
 sg13g2_or2_1 _15877_ (.X(_07465_),
    .B(_07460_),
    .A(_07459_));
 sg13g2_or2_1 _15878_ (.X(_07466_),
    .B(_07464_),
    .A(_07460_));
 sg13g2_a21oi_1 _15879_ (.A1(_07446_),
    .A2(_07448_),
    .Y(_07467_),
    .B1(_07445_));
 sg13g2_and2_1 _15880_ (.A(\TRNG.sha256.W[10] ),
    .B(\TRNG.sha256.K[10] ),
    .X(_07468_));
 sg13g2_xor2_1 _15881_ (.B(\TRNG.sha256.K[10] ),
    .A(\TRNG.sha256.W[10] ),
    .X(_07469_));
 sg13g2_xnor2_1 _15882_ (.Y(_07470_),
    .A(\TRNG.hash[10] ),
    .B(_07469_));
 sg13g2_o21ai_1 _15883_ (.B1(\TRNG.hash[9] ),
    .Y(_07471_),
    .A1(\TRNG.sha256.W[9] ),
    .A2(\TRNG.sha256.K[9] ));
 sg13g2_nand2_1 _15884_ (.Y(_07472_),
    .A(_07442_),
    .B(_07471_));
 sg13g2_nor2b_1 _15885_ (.A(_07470_),
    .B_N(_07472_),
    .Y(_07473_));
 sg13g2_nand2b_1 _15886_ (.Y(_07474_),
    .B(_07470_),
    .A_N(_07472_));
 sg13g2_xor2_1 _15887_ (.B(_07472_),
    .A(_07470_),
    .X(_07475_));
 sg13g2_xnor2_1 _15888_ (.Y(_07476_),
    .A(\TRNG.hash[117] ),
    .B(net5891));
 sg13g2_xnor2_1 _15889_ (.Y(_07477_),
    .A(net5552),
    .B(_07476_));
 sg13g2_xnor2_1 _15890_ (.Y(_07478_),
    .A(_07475_),
    .B(_07477_));
 sg13g2_nand2b_1 _15891_ (.Y(_07479_),
    .B(_07478_),
    .A_N(_07467_));
 sg13g2_xor2_1 _15892_ (.B(_07478_),
    .A(_07467_),
    .X(_07480_));
 sg13g2_mux2_2 _15893_ (.A0(_00165_),
    .A1(_00193_),
    .S(net5895),
    .X(_07481_));
 sg13g2_xnor2_1 _15894_ (.Y(_07482_),
    .A(_07480_),
    .B(_07481_));
 sg13g2_a21oi_1 _15895_ (.A1(_07451_),
    .A2(_07452_),
    .Y(_07483_),
    .B1(_07450_));
 sg13g2_or2_1 _15896_ (.X(_07484_),
    .B(_07483_),
    .A(_07482_));
 sg13g2_xnor2_1 _15897_ (.Y(_07485_),
    .A(_07482_),
    .B(_07483_));
 sg13g2_a21oi_1 _15898_ (.A1(_07425_),
    .A2(_07455_),
    .Y(_07486_),
    .B1(_07454_));
 sg13g2_nor2_1 _15899_ (.A(_07426_),
    .B(_07456_),
    .Y(_07487_));
 sg13g2_a21oi_1 _15900_ (.A1(_07430_),
    .A2(_07487_),
    .Y(_07488_),
    .B1(_07486_));
 sg13g2_xnor2_1 _15901_ (.Y(_07489_),
    .A(_07485_),
    .B(_07488_));
 sg13g2_xor2_1 _15902_ (.B(_07489_),
    .A(\TRNG.hash[138] ),
    .X(_07490_));
 sg13g2_nor2_1 _15903_ (.A(_07466_),
    .B(_07490_),
    .Y(_07491_));
 sg13g2_xnor2_1 _15904_ (.Y(_07492_),
    .A(_07466_),
    .B(_07490_));
 sg13g2_o21ai_1 _15905_ (.B1(_00206_),
    .Y(_07493_),
    .A1(\TRNG.hash[105] ),
    .A2(_07436_));
 sg13g2_xor2_1 _15906_ (.B(_07493_),
    .A(net3159),
    .X(_07494_));
 sg13g2_o21ai_1 _15907_ (.B1(net4977),
    .Y(_07495_),
    .A1(net5895),
    .A2(net5177));
 sg13g2_a221oi_1 _15908_ (.B2(net5187),
    .C1(_07495_),
    .B1(net3160),
    .A1(net5846),
    .Y(_00538_),
    .A2(_07492_));
 sg13g2_o21ai_1 _15909_ (.B1(_07484_),
    .Y(_07496_),
    .A1(_07485_),
    .A2(_07488_));
 sg13g2_o21ai_1 _15910_ (.B1(_07479_),
    .Y(_07497_),
    .A1(_07480_),
    .A2(_07481_));
 sg13g2_a21oi_1 _15911_ (.A1(_07474_),
    .A2(_07477_),
    .Y(_07498_),
    .B1(_07473_));
 sg13g2_a21oi_1 _15912_ (.A1(\TRNG.hash[10] ),
    .A2(_07469_),
    .Y(_07499_),
    .B1(_07468_));
 sg13g2_and2_1 _15913_ (.A(\TRNG.sha256.W[11] ),
    .B(\TRNG.sha256.K[11] ),
    .X(_07500_));
 sg13g2_xor2_1 _15914_ (.B(\TRNG.sha256.K[11] ),
    .A(\TRNG.sha256.W[11] ),
    .X(_07501_));
 sg13g2_xnor2_1 _15915_ (.Y(_07502_),
    .A(\TRNG.hash[11] ),
    .B(_07501_));
 sg13g2_nor2_1 _15916_ (.A(_07499_),
    .B(_07502_),
    .Y(_07503_));
 sg13g2_xor2_1 _15917_ (.B(_07502_),
    .A(_07499_),
    .X(_07504_));
 sg13g2_xnor2_1 _15918_ (.Y(_07505_),
    .A(net5551),
    .B(\TRNG.hash[118] ));
 sg13g2_xnor2_1 _15919_ (.Y(_07506_),
    .A(\TRNG.hash[113] ),
    .B(_07505_));
 sg13g2_xnor2_1 _15920_ (.Y(_07507_),
    .A(_07504_),
    .B(_07506_));
 sg13g2_or2_1 _15921_ (.X(_07508_),
    .B(_07507_),
    .A(_07498_));
 sg13g2_xnor2_1 _15922_ (.Y(_07509_),
    .A(_07498_),
    .B(_07507_));
 sg13g2_mux2_2 _15923_ (.A0(_00175_),
    .A1(_00182_),
    .S(net5894),
    .X(_07510_));
 sg13g2_xor2_1 _15924_ (.B(_07510_),
    .A(_07509_),
    .X(_07511_));
 sg13g2_nor2_1 _15925_ (.A(_07497_),
    .B(_07511_),
    .Y(_07512_));
 sg13g2_nand2_1 _15926_ (.Y(_07513_),
    .A(_07497_),
    .B(_07511_));
 sg13g2_xnor2_1 _15927_ (.Y(_07514_),
    .A(_07497_),
    .B(_07511_));
 sg13g2_xnor2_1 _15928_ (.Y(_07515_),
    .A(_07496_),
    .B(_07514_));
 sg13g2_nor2_1 _15929_ (.A(\TRNG.hash[139] ),
    .B(_07515_),
    .Y(_07516_));
 sg13g2_inv_1 _15930_ (.Y(_07517_),
    .A(_07516_));
 sg13g2_and2_1 _15931_ (.A(\TRNG.hash[139] ),
    .B(_07515_),
    .X(_07518_));
 sg13g2_or2_1 _15932_ (.X(_07519_),
    .B(_07518_),
    .A(_07516_));
 sg13g2_nor2_1 _15933_ (.A(_00136_),
    .B(_07489_),
    .Y(_07520_));
 sg13g2_nor3_1 _15934_ (.A(_07491_),
    .B(_07519_),
    .C(_07520_),
    .Y(_07521_));
 sg13g2_o21ai_1 _15935_ (.B1(_07519_),
    .Y(_07522_),
    .A1(_07491_),
    .A2(_07520_));
 sg13g2_nor2_1 _15936_ (.A(net5490),
    .B(_07521_),
    .Y(_07523_));
 sg13g2_nand2_1 _15937_ (.Y(_07524_),
    .A(net5895),
    .B(_07493_));
 sg13g2_xor2_1 _15938_ (.B(_07524_),
    .A(net5894),
    .X(_07525_));
 sg13g2_o21ai_1 _15939_ (.B1(net4977),
    .Y(_07526_),
    .A1(net5894),
    .A2(net5177));
 sg13g2_a221oi_1 _15940_ (.B2(net5187),
    .C1(_07526_),
    .B1(_07525_),
    .A1(_07522_),
    .Y(_00539_),
    .A2(_07523_));
 sg13g2_a21oi_1 _15941_ (.A1(_07517_),
    .A2(_07520_),
    .Y(_07527_),
    .B1(_07518_));
 sg13g2_o21ai_1 _15942_ (.B1(_07527_),
    .Y(_07528_),
    .A1(_07460_),
    .A2(_07464_));
 sg13g2_o21ai_1 _15943_ (.B1(_07527_),
    .Y(_07529_),
    .A1(_07490_),
    .A2(_07516_));
 sg13g2_a21oi_2 _15944_ (.B1(_07503_),
    .Y(_07530_),
    .A2(_07506_),
    .A1(_07504_));
 sg13g2_a21oi_1 _15945_ (.A1(\TRNG.hash[11] ),
    .A2(_07501_),
    .Y(_07531_),
    .B1(_07500_));
 sg13g2_nand2_1 _15946_ (.Y(_07532_),
    .A(\TRNG.sha256.W[12] ),
    .B(\TRNG.sha256.K[12] ));
 sg13g2_xor2_1 _15947_ (.B(\TRNG.sha256.K[12] ),
    .A(\TRNG.sha256.W[12] ),
    .X(_07533_));
 sg13g2_xnor2_1 _15948_ (.Y(_07534_),
    .A(_00154_),
    .B(_07533_));
 sg13g2_nor2b_1 _15949_ (.A(_07531_),
    .B_N(_07534_),
    .Y(_07535_));
 sg13g2_xnor2_1 _15950_ (.Y(_07536_),
    .A(_07531_),
    .B(_07534_));
 sg13g2_xnor2_1 _15951_ (.Y(_07537_),
    .A(\TRNG.hash[101] ),
    .B(\TRNG.hash[119] ));
 sg13g2_xnor2_1 _15952_ (.Y(_07538_),
    .A(net5545),
    .B(_07537_));
 sg13g2_xnor2_1 _15953_ (.Y(_07539_),
    .A(_07536_),
    .B(_07538_));
 sg13g2_or2_1 _15954_ (.X(_07540_),
    .B(_07539_),
    .A(_07530_));
 sg13g2_and2_1 _15955_ (.A(_07530_),
    .B(_07539_),
    .X(_07541_));
 sg13g2_xnor2_1 _15956_ (.Y(_07542_),
    .A(_07530_),
    .B(_07539_));
 sg13g2_mux2_1 _15957_ (.A0(_00167_),
    .A1(_00181_),
    .S(net5548),
    .X(_07543_));
 sg13g2_xnor2_1 _15958_ (.Y(_07544_),
    .A(_07542_),
    .B(_07543_));
 sg13g2_o21ai_1 _15959_ (.B1(_07508_),
    .Y(_07545_),
    .A1(_07509_),
    .A2(_07510_));
 sg13g2_nand2b_1 _15960_ (.Y(_07546_),
    .B(_07545_),
    .A_N(_07544_));
 sg13g2_xor2_1 _15961_ (.B(_07545_),
    .A(_07544_),
    .X(_07547_));
 sg13g2_nor2_1 _15962_ (.A(_07485_),
    .B(_07514_),
    .Y(_07548_));
 sg13g2_o21ai_1 _15963_ (.B1(_07513_),
    .Y(_07549_),
    .A1(_07484_),
    .A2(_07512_));
 sg13g2_a21o_1 _15964_ (.A2(_07548_),
    .A1(_07486_),
    .B1(_07549_),
    .X(_07550_));
 sg13g2_nand2_1 _15965_ (.Y(_07551_),
    .A(_07487_),
    .B(_07548_));
 sg13g2_a221oi_1 _15966_ (.B2(_07367_),
    .C1(_07551_),
    .B1(_07429_),
    .A1(_07427_),
    .Y(_07552_),
    .A2(_07428_));
 sg13g2_nor2_1 _15967_ (.A(_07550_),
    .B(_07552_),
    .Y(_07553_));
 sg13g2_xnor2_1 _15968_ (.Y(_07554_),
    .A(_07547_),
    .B(_07553_));
 sg13g2_xor2_1 _15969_ (.B(_07554_),
    .A(\TRNG.hash[140] ),
    .X(_07555_));
 sg13g2_inv_1 _15970_ (.Y(_07556_),
    .A(_07555_));
 sg13g2_and3_1 _15971_ (.X(_07557_),
    .A(_07528_),
    .B(_07529_),
    .C(_07556_));
 sg13g2_nand3_1 _15972_ (.B(_07529_),
    .C(_07556_),
    .A(_07528_),
    .Y(_07558_));
 sg13g2_nor2_1 _15973_ (.A(_00138_),
    .B(_07554_),
    .Y(_07559_));
 sg13g2_nor2_1 _15974_ (.A(_07557_),
    .B(_07559_),
    .Y(_07560_));
 sg13g2_o21ai_1 _15975_ (.B1(_07546_),
    .Y(_07561_),
    .A1(_07547_),
    .A2(_07553_));
 sg13g2_o21ai_1 _15976_ (.B1(_07540_),
    .Y(_07562_),
    .A1(_07541_),
    .A2(_07543_));
 sg13g2_a21oi_1 _15977_ (.A1(_07536_),
    .A2(_07538_),
    .Y(_07563_),
    .B1(_07535_));
 sg13g2_and2_1 _15978_ (.A(\TRNG.sha256.W[13] ),
    .B(\TRNG.sha256.K[13] ),
    .X(_07564_));
 sg13g2_xor2_1 _15979_ (.B(\TRNG.sha256.K[13] ),
    .A(\TRNG.sha256.W[13] ),
    .X(_07565_));
 sg13g2_xnor2_1 _15980_ (.Y(_07566_),
    .A(\TRNG.hash[13] ),
    .B(_07565_));
 sg13g2_o21ai_1 _15981_ (.B1(\TRNG.hash[12] ),
    .Y(_07567_),
    .A1(\TRNG.sha256.W[12] ),
    .A2(\TRNG.sha256.K[12] ));
 sg13g2_nand2_1 _15982_ (.Y(_07568_),
    .A(_07532_),
    .B(_07567_));
 sg13g2_nor2b_1 _15983_ (.A(_07566_),
    .B_N(_07568_),
    .Y(_07569_));
 sg13g2_xnor2_1 _15984_ (.Y(_07570_),
    .A(_07566_),
    .B(_07568_));
 sg13g2_xnor2_1 _15985_ (.Y(_07571_),
    .A(net5544),
    .B(\TRNG.hash[102] ));
 sg13g2_xnor2_1 _15986_ (.Y(_07572_),
    .A(\TRNG.hash[120] ),
    .B(_07571_));
 sg13g2_xor2_1 _15987_ (.B(_07572_),
    .A(_07570_),
    .X(_07573_));
 sg13g2_nand2b_1 _15988_ (.Y(_07574_),
    .B(_07573_),
    .A_N(_07563_));
 sg13g2_xor2_1 _15989_ (.B(_07573_),
    .A(_07563_),
    .X(_07575_));
 sg13g2_mux2_2 _15990_ (.A0(_00166_),
    .A1(_00194_),
    .S(net5893),
    .X(_07576_));
 sg13g2_xor2_1 _15991_ (.B(_07576_),
    .A(_07575_),
    .X(_07577_));
 sg13g2_nand2_1 _15992_ (.Y(_07578_),
    .A(_07562_),
    .B(_07577_));
 sg13g2_xnor2_1 _15993_ (.Y(_07579_),
    .A(_07562_),
    .B(_07577_));
 sg13g2_xor2_1 _15994_ (.B(_07579_),
    .A(_07561_),
    .X(_07580_));
 sg13g2_xnor2_1 _15995_ (.Y(_07581_),
    .A(_00207_),
    .B(_07580_));
 sg13g2_nor2b_1 _15996_ (.A(_07560_),
    .B_N(_07581_),
    .Y(_07582_));
 sg13g2_nor3_1 _15997_ (.A(_07557_),
    .B(_07559_),
    .C(_07581_),
    .Y(_07583_));
 sg13g2_nor3_1 _15998_ (.A(net5484),
    .B(_07582_),
    .C(_07583_),
    .Y(_07584_));
 sg13g2_nand2_1 _15999_ (.Y(_07585_),
    .A(net5894),
    .B(net5895));
 sg13g2_a21oi_2 _16000_ (.B1(_07585_),
    .Y(_07586_),
    .A2(_07436_),
    .A1(_04222_));
 sg13g2_o21ai_1 _16001_ (.B1(net5893),
    .Y(_07587_),
    .A1(net5548),
    .A2(_07586_));
 sg13g2_or3_1 _16002_ (.A(net5548),
    .B(net5893),
    .C(_07586_),
    .X(_07588_));
 sg13g2_a21oi_1 _16003_ (.A1(_07587_),
    .A2(_07588_),
    .Y(_07589_),
    .B1(net5180));
 sg13g2_o21ai_1 _16004_ (.B1(net4977),
    .Y(_07590_),
    .A1(net5893),
    .A2(net5177));
 sg13g2_nor3_1 _16005_ (.A(_07584_),
    .B(_07589_),
    .C(_07590_),
    .Y(_00540_));
 sg13g2_a21oi_1 _16006_ (.A1(\TRNG.hash[13] ),
    .A2(_07565_),
    .Y(_07591_),
    .B1(_07564_));
 sg13g2_and2_1 _16007_ (.A(\TRNG.sha256.W[14] ),
    .B(\TRNG.sha256.K[14] ),
    .X(_07592_));
 sg13g2_xor2_1 _16008_ (.B(\TRNG.sha256.K[14] ),
    .A(\TRNG.sha256.W[14] ),
    .X(_07593_));
 sg13g2_xnor2_1 _16009_ (.Y(_07594_),
    .A(\TRNG.hash[14] ),
    .B(_07593_));
 sg13g2_nor2_1 _16010_ (.A(_07591_),
    .B(_07594_),
    .Y(_07595_));
 sg13g2_xor2_1 _16011_ (.B(_07594_),
    .A(_07591_),
    .X(_07596_));
 sg13g2_xnor2_1 _16012_ (.Y(_07597_),
    .A(net5890),
    .B(net5897));
 sg13g2_xnor2_1 _16013_ (.Y(_07598_),
    .A(\TRNG.hash[121] ),
    .B(_07597_));
 sg13g2_a21oi_1 _16014_ (.A1(_07596_),
    .A2(_07598_),
    .Y(_07599_),
    .B1(_07595_));
 sg13g2_a21oi_2 _16015_ (.B1(_07592_),
    .Y(_07600_),
    .A2(_07593_),
    .A1(\TRNG.hash[14] ));
 sg13g2_and2_1 _16016_ (.A(\TRNG.sha256.W[15] ),
    .B(\TRNG.sha256.K[15] ),
    .X(_07601_));
 sg13g2_xor2_1 _16017_ (.B(\TRNG.sha256.K[15] ),
    .A(\TRNG.sha256.W[15] ),
    .X(_07602_));
 sg13g2_xnor2_1 _16018_ (.Y(_07603_),
    .A(\TRNG.hash[15] ),
    .B(_07602_));
 sg13g2_nor2_1 _16019_ (.A(_07600_),
    .B(_07603_),
    .Y(_07604_));
 sg13g2_xor2_1 _16020_ (.B(_07603_),
    .A(_07600_),
    .X(_07605_));
 sg13g2_xnor2_1 _16021_ (.Y(_07606_),
    .A(net5889),
    .B(net5896));
 sg13g2_xnor2_1 _16022_ (.Y(_07607_),
    .A(\TRNG.hash[122] ),
    .B(_07606_));
 sg13g2_xnor2_1 _16023_ (.Y(_07608_),
    .A(_07605_),
    .B(_07607_));
 sg13g2_nor2_1 _16024_ (.A(_07599_),
    .B(_07608_),
    .Y(_07609_));
 sg13g2_xor2_1 _16025_ (.B(_07608_),
    .A(_07599_),
    .X(_07610_));
 sg13g2_mux2_1 _16026_ (.A0(_00210_),
    .A1(_00183_),
    .S(net5892),
    .X(_07611_));
 sg13g2_inv_1 _16027_ (.Y(_07612_),
    .A(_07611_));
 sg13g2_xnor2_1 _16028_ (.Y(_07613_),
    .A(_07610_),
    .B(_07612_));
 sg13g2_a21oi_1 _16029_ (.A1(_07570_),
    .A2(_07572_),
    .Y(_07614_),
    .B1(_07569_));
 sg13g2_xnor2_1 _16030_ (.Y(_07615_),
    .A(_07596_),
    .B(_07598_));
 sg13g2_nor2_1 _16031_ (.A(_07614_),
    .B(_07615_),
    .Y(_07616_));
 sg13g2_xor2_1 _16032_ (.B(_07615_),
    .A(_07614_),
    .X(_07617_));
 sg13g2_mux2_2 _16033_ (.A0(\TRNG.hash[46] ),
    .A1(\TRNG.hash[78] ),
    .S(net5547),
    .X(_07618_));
 sg13g2_a21oi_2 _16034_ (.B1(_07616_),
    .Y(_07619_),
    .A2(_07618_),
    .A1(_07617_));
 sg13g2_nand2_1 _16035_ (.Y(_07620_),
    .A(_07613_),
    .B(_07619_));
 sg13g2_nor2_1 _16036_ (.A(_07613_),
    .B(_07619_),
    .Y(_07621_));
 sg13g2_xnor2_1 _16037_ (.Y(_07622_),
    .A(_07613_),
    .B(_07619_));
 sg13g2_xnor2_1 _16038_ (.Y(_07623_),
    .A(_07617_),
    .B(_07618_));
 sg13g2_o21ai_1 _16039_ (.B1(_07574_),
    .Y(_07624_),
    .A1(_07575_),
    .A2(_07576_));
 sg13g2_nor2b_1 _16040_ (.A(_07623_),
    .B_N(_07624_),
    .Y(_07625_));
 sg13g2_xor2_1 _16041_ (.B(_07624_),
    .A(_07623_),
    .X(_07626_));
 sg13g2_inv_1 _16042_ (.Y(_07627_),
    .A(_07626_));
 sg13g2_o21ai_1 _16043_ (.B1(_07578_),
    .Y(_07628_),
    .A1(_07546_),
    .A2(_07579_));
 sg13g2_nor2_1 _16044_ (.A(_07547_),
    .B(_07579_),
    .Y(_07629_));
 sg13g2_o21ai_1 _16045_ (.B1(_07629_),
    .Y(_07630_),
    .A1(_07550_),
    .A2(_07552_));
 sg13g2_nand2b_1 _16046_ (.Y(_07631_),
    .B(_07630_),
    .A_N(_07628_));
 sg13g2_a21oi_1 _16047_ (.A1(_07627_),
    .A2(_07631_),
    .Y(_07632_),
    .B1(_07625_));
 sg13g2_xnor2_1 _16048_ (.Y(_07633_),
    .A(_07622_),
    .B(_07632_));
 sg13g2_nand2b_1 _16049_ (.Y(_07634_),
    .B(\TRNG.hash[143] ),
    .A_N(_07633_));
 sg13g2_xnor2_1 _16050_ (.Y(_07635_),
    .A(\TRNG.hash[143] ),
    .B(_07633_));
 sg13g2_xnor2_1 _16051_ (.Y(_07636_),
    .A(_07627_),
    .B(_07631_));
 sg13g2_nor2_1 _16052_ (.A(_04232_),
    .B(_07636_),
    .Y(_07637_));
 sg13g2_xnor2_1 _16053_ (.Y(_07638_),
    .A(_04232_),
    .B(_07636_));
 sg13g2_or2_1 _16054_ (.X(_07639_),
    .B(_07580_),
    .A(_04233_));
 sg13g2_nor2b_1 _16055_ (.A(_07559_),
    .B_N(_07639_),
    .Y(_07640_));
 sg13g2_a22oi_1 _16056_ (.Y(_07641_),
    .B1(_07640_),
    .B2(_07558_),
    .A2(_07639_),
    .A1(_07581_));
 sg13g2_a221oi_1 _16057_ (.B2(_07558_),
    .C1(_07638_),
    .B1(_07640_),
    .A1(_07581_),
    .Y(_07642_),
    .A2(_07639_));
 sg13g2_o21ai_1 _16058_ (.B1(_07635_),
    .Y(_07643_),
    .A1(_07637_),
    .A2(_07642_));
 sg13g2_or3_1 _16059_ (.A(_07635_),
    .B(_07637_),
    .C(_07642_),
    .X(_07644_));
 sg13g2_nand2_1 _16060_ (.Y(_07645_),
    .A(_07643_),
    .B(_07644_));
 sg13g2_nand2b_1 _16061_ (.Y(_07646_),
    .B(_07587_),
    .A_N(net5547));
 sg13g2_xor2_1 _16062_ (.B(_07646_),
    .A(net3134),
    .X(_07647_));
 sg13g2_o21ai_1 _16063_ (.B1(net4975),
    .Y(_07648_),
    .A1(net5892),
    .A2(net5176));
 sg13g2_a221oi_1 _16064_ (.B2(net5186),
    .C1(_07648_),
    .B1(_07647_),
    .A1(net5850),
    .Y(_00541_),
    .A2(_07645_));
 sg13g2_nand2_2 _16065_ (.Y(_07649_),
    .A(_07634_),
    .B(_07643_));
 sg13g2_nor2_1 _16066_ (.A(_07622_),
    .B(_07626_),
    .Y(_07650_));
 sg13g2_nor4_2 _16067_ (.A(_07547_),
    .B(_07579_),
    .C(_07622_),
    .Y(_07651_),
    .D(_07626_));
 sg13g2_a21o_1 _16068_ (.A2(_07625_),
    .A1(_07620_),
    .B1(_07621_),
    .X(_07652_));
 sg13g2_a21o_1 _16069_ (.A2(_07650_),
    .A1(_07628_),
    .B1(_07652_),
    .X(_07653_));
 sg13g2_a21o_1 _16070_ (.A2(_07651_),
    .A1(_07550_),
    .B1(_07653_),
    .X(_07654_));
 sg13g2_nand3_1 _16071_ (.B(_07548_),
    .C(_07651_),
    .A(_07487_),
    .Y(_07655_));
 sg13g2_a221oi_1 _16072_ (.B2(_07367_),
    .C1(_07655_),
    .B1(_07429_),
    .A1(_07427_),
    .Y(_07656_),
    .A2(_07428_));
 sg13g2_nor2_2 _16073_ (.A(_07654_),
    .B(_07656_),
    .Y(_07657_));
 sg13g2_a21oi_1 _16074_ (.A1(_07605_),
    .A2(_07607_),
    .Y(_07658_),
    .B1(_07604_));
 sg13g2_a21oi_1 _16075_ (.A1(\TRNG.hash[15] ),
    .A2(_07602_),
    .Y(_07659_),
    .B1(_07601_));
 sg13g2_and2_1 _16076_ (.A(\TRNG.sha256.W[16] ),
    .B(\TRNG.sha256.K[16] ),
    .X(_07660_));
 sg13g2_xor2_1 _16077_ (.B(\TRNG.sha256.K[16] ),
    .A(\TRNG.sha256.W[16] ),
    .X(_07661_));
 sg13g2_xnor2_1 _16078_ (.Y(_07662_),
    .A(\TRNG.hash[16] ),
    .B(_07661_));
 sg13g2_nor2_1 _16079_ (.A(_07659_),
    .B(_07662_),
    .Y(_07663_));
 sg13g2_xor2_1 _16080_ (.B(_07662_),
    .A(_07659_),
    .X(_07664_));
 sg13g2_xnor2_1 _16081_ (.Y(_07665_),
    .A(\TRNG.hash[123] ),
    .B(\TRNG.hash[118] ));
 sg13g2_xnor2_1 _16082_ (.Y(_07666_),
    .A(\TRNG.hash[105] ),
    .B(_07665_));
 sg13g2_xnor2_1 _16083_ (.Y(_07667_),
    .A(_07664_),
    .B(_07666_));
 sg13g2_nor2_1 _16084_ (.A(_07658_),
    .B(_07667_),
    .Y(_07668_));
 sg13g2_xnor2_1 _16085_ (.Y(_07669_),
    .A(_07658_),
    .B(_07667_));
 sg13g2_mux2_1 _16086_ (.A0(_00176_),
    .A1(_00185_),
    .S(net5891),
    .X(_07670_));
 sg13g2_nor2_1 _16087_ (.A(_07669_),
    .B(_07670_),
    .Y(_07671_));
 sg13g2_xnor2_1 _16088_ (.Y(_07672_),
    .A(_07669_),
    .B(_07670_));
 sg13g2_a21oi_1 _16089_ (.A1(_07610_),
    .A2(_07612_),
    .Y(_07673_),
    .B1(_07609_));
 sg13g2_or2_1 _16090_ (.X(_07674_),
    .B(_07673_),
    .A(_07672_));
 sg13g2_xnor2_1 _16091_ (.Y(_07675_),
    .A(_07672_),
    .B(_07673_));
 sg13g2_xor2_1 _16092_ (.B(_07675_),
    .A(_07657_),
    .X(_07676_));
 sg13g2_and2_1 _16093_ (.A(\TRNG.hash[144] ),
    .B(_07676_),
    .X(_07677_));
 sg13g2_xnor2_1 _16094_ (.Y(_07678_),
    .A(\TRNG.hash[144] ),
    .B(_07676_));
 sg13g2_nand2b_1 _16095_ (.Y(_07679_),
    .B(_07649_),
    .A_N(_07678_));
 sg13g2_xor2_1 _16096_ (.B(_07678_),
    .A(_07649_),
    .X(_07680_));
 sg13g2_and3_1 _16097_ (.X(_07681_),
    .A(net5891),
    .B(net5892),
    .C(_07646_));
 sg13g2_a21oi_1 _16098_ (.A1(net5892),
    .A2(_07646_),
    .Y(_07682_),
    .B1(net5891));
 sg13g2_or2_1 _16099_ (.X(_07683_),
    .B(_07682_),
    .A(_07681_));
 sg13g2_o21ai_1 _16100_ (.B1(net4975),
    .Y(_07684_),
    .A1(net5891),
    .A2(net5176));
 sg13g2_a221oi_1 _16101_ (.B2(net5186),
    .C1(_07684_),
    .B1(_07683_),
    .A1(net5850),
    .Y(_00542_),
    .A2(_07680_));
 sg13g2_a21oi_1 _16102_ (.A1(\TRNG.hash[16] ),
    .A2(_07661_),
    .Y(_07685_),
    .B1(_07660_));
 sg13g2_and2_1 _16103_ (.A(\TRNG.sha256.W[17] ),
    .B(\TRNG.sha256.K[17] ),
    .X(_07686_));
 sg13g2_xor2_1 _16104_ (.B(\TRNG.sha256.K[17] ),
    .A(\TRNG.sha256.W[17] ),
    .X(_07687_));
 sg13g2_xnor2_1 _16105_ (.Y(_07688_),
    .A(\TRNG.hash[17] ),
    .B(_07687_));
 sg13g2_nor2_1 _16106_ (.A(_07685_),
    .B(_07688_),
    .Y(_07689_));
 sg13g2_xor2_1 _16107_ (.B(_07688_),
    .A(_07685_),
    .X(_07690_));
 sg13g2_xnor2_1 _16108_ (.Y(_07691_),
    .A(\TRNG.hash[119] ),
    .B(net5895));
 sg13g2_xnor2_1 _16109_ (.Y(_07692_),
    .A(\TRNG.hash[124] ),
    .B(_07691_));
 sg13g2_a21oi_1 _16110_ (.A1(_07690_),
    .A2(_07692_),
    .Y(_07693_),
    .B1(_07689_));
 sg13g2_a21oi_1 _16111_ (.A1(\TRNG.hash[17] ),
    .A2(_07687_),
    .Y(_07694_),
    .B1(_07686_));
 sg13g2_and2_1 _16112_ (.A(\TRNG.sha256.W[18] ),
    .B(\TRNG.sha256.K[18] ),
    .X(_07695_));
 sg13g2_xor2_1 _16113_ (.B(\TRNG.sha256.K[18] ),
    .A(\TRNG.sha256.W[18] ),
    .X(_07696_));
 sg13g2_xnor2_1 _16114_ (.Y(_07697_),
    .A(\TRNG.hash[18] ),
    .B(_07696_));
 sg13g2_nor2_1 _16115_ (.A(_07694_),
    .B(_07697_),
    .Y(_07698_));
 sg13g2_xor2_1 _16116_ (.B(_07697_),
    .A(_07694_),
    .X(_07699_));
 sg13g2_xnor2_1 _16117_ (.Y(_07700_),
    .A(\TRNG.hash[125] ),
    .B(net5894));
 sg13g2_xnor2_1 _16118_ (.Y(_07701_),
    .A(\TRNG.hash[120] ),
    .B(_07700_));
 sg13g2_xnor2_1 _16119_ (.Y(_07702_),
    .A(_07699_),
    .B(_07701_));
 sg13g2_nor2_1 _16120_ (.A(_07693_),
    .B(_07702_),
    .Y(_07703_));
 sg13g2_xnor2_1 _16121_ (.Y(_07704_),
    .A(_07693_),
    .B(_07702_));
 sg13g2_mux2_1 _16122_ (.A0(_00168_),
    .A1(_00195_),
    .S(\TRNG.hash[114] ),
    .X(_07705_));
 sg13g2_nor2_1 _16123_ (.A(_07704_),
    .B(_07705_),
    .Y(_07706_));
 sg13g2_a21oi_1 _16124_ (.A1(_07699_),
    .A2(_07701_),
    .Y(_07707_),
    .B1(_07698_));
 sg13g2_a21oi_1 _16125_ (.A1(\TRNG.hash[18] ),
    .A2(_07696_),
    .Y(_07708_),
    .B1(_07695_));
 sg13g2_and2_1 _16126_ (.A(\TRNG.sha256.W[19] ),
    .B(\TRNG.sha256.K[19] ),
    .X(_07709_));
 sg13g2_xor2_1 _16127_ (.B(\TRNG.sha256.K[19] ),
    .A(\TRNG.sha256.W[19] ),
    .X(_07710_));
 sg13g2_xnor2_1 _16128_ (.Y(_07711_),
    .A(\TRNG.hash[19] ),
    .B(_07710_));
 sg13g2_nor2_1 _16129_ (.A(_07708_),
    .B(_07711_),
    .Y(_07712_));
 sg13g2_xor2_1 _16130_ (.B(_07711_),
    .A(_07708_),
    .X(_07713_));
 sg13g2_xnor2_1 _16131_ (.Y(_07714_),
    .A(\TRNG.hash[108] ),
    .B(\TRNG.hash[121] ));
 sg13g2_xnor2_1 _16132_ (.Y(_07715_),
    .A(\TRNG.hash[126] ),
    .B(_07714_));
 sg13g2_xnor2_1 _16133_ (.Y(_07716_),
    .A(_07713_),
    .B(_07715_));
 sg13g2_nor2_1 _16134_ (.A(_07707_),
    .B(_07716_),
    .Y(_07717_));
 sg13g2_xor2_1 _16135_ (.B(_07716_),
    .A(_07707_),
    .X(_07718_));
 sg13g2_mux2_2 _16136_ (.A0(\TRNG.hash[51] ),
    .A1(\TRNG.hash[83] ),
    .S(\TRNG.hash[115] ),
    .X(_07719_));
 sg13g2_xor2_1 _16137_ (.B(_07719_),
    .A(_07718_),
    .X(_07720_));
 sg13g2_nor3_1 _16138_ (.A(_07703_),
    .B(_07706_),
    .C(_07720_),
    .Y(_07721_));
 sg13g2_o21ai_1 _16139_ (.B1(_07720_),
    .Y(_07722_),
    .A1(_07703_),
    .A2(_07706_));
 sg13g2_nand2b_1 _16140_ (.Y(_07723_),
    .B(_07722_),
    .A_N(_07721_));
 sg13g2_xnor2_1 _16141_ (.Y(_07724_),
    .A(_07704_),
    .B(_07705_));
 sg13g2_a21oi_1 _16142_ (.A1(_07664_),
    .A2(_07666_),
    .Y(_07725_),
    .B1(_07663_));
 sg13g2_xnor2_1 _16143_ (.Y(_07726_),
    .A(_07690_),
    .B(_07692_));
 sg13g2_xor2_1 _16144_ (.B(_07726_),
    .A(_07725_),
    .X(_07727_));
 sg13g2_mux2_1 _16145_ (.A0(\TRNG.hash[49] ),
    .A1(\TRNG.hash[81] ),
    .S(net5546),
    .X(_07728_));
 sg13g2_nand2_1 _16146_ (.Y(_07729_),
    .A(_07727_),
    .B(_07728_));
 sg13g2_o21ai_1 _16147_ (.B1(_07729_),
    .Y(_07730_),
    .A1(_07725_),
    .A2(_07726_));
 sg13g2_nor2b_1 _16148_ (.A(_07724_),
    .B_N(_07730_),
    .Y(_07731_));
 sg13g2_xor2_1 _16149_ (.B(_07730_),
    .A(_07724_),
    .X(_07732_));
 sg13g2_inv_1 _16150_ (.Y(_07733_),
    .A(_07732_));
 sg13g2_xor2_1 _16151_ (.B(_07728_),
    .A(_07727_),
    .X(_07734_));
 sg13g2_o21ai_1 _16152_ (.B1(_07734_),
    .Y(_07735_),
    .A1(_07668_),
    .A2(_07671_));
 sg13g2_or3_1 _16153_ (.A(_07668_),
    .B(_07671_),
    .C(_07734_),
    .X(_07736_));
 sg13g2_nand2_1 _16154_ (.Y(_07737_),
    .A(_07674_),
    .B(_07735_));
 sg13g2_nand2_1 _16155_ (.Y(_07738_),
    .A(_07736_),
    .B(_07737_));
 sg13g2_nand2_1 _16156_ (.Y(_07739_),
    .A(_07735_),
    .B(_07736_));
 sg13g2_nor2_1 _16157_ (.A(_07675_),
    .B(_07739_),
    .Y(_07740_));
 sg13g2_inv_1 _16158_ (.Y(_07741_),
    .A(_07740_));
 sg13g2_o21ai_1 _16159_ (.B1(_07738_),
    .Y(_07742_),
    .A1(_07657_),
    .A2(_07741_));
 sg13g2_a21oi_1 _16160_ (.A1(_07733_),
    .A2(_07742_),
    .Y(_07743_),
    .B1(_07731_));
 sg13g2_xnor2_1 _16161_ (.Y(_07744_),
    .A(_07723_),
    .B(_07743_));
 sg13g2_inv_1 _16162_ (.Y(_07745_),
    .A(_07744_));
 sg13g2_xnor2_1 _16163_ (.Y(_07746_),
    .A(\TRNG.hash[147] ),
    .B(_07744_));
 sg13g2_inv_1 _16164_ (.Y(_07747_),
    .A(_07746_));
 sg13g2_xnor2_1 _16165_ (.Y(_07748_),
    .A(_07733_),
    .B(_07742_));
 sg13g2_nor2_1 _16166_ (.A(_04230_),
    .B(_07748_),
    .Y(_07749_));
 sg13g2_xnor2_1 _16167_ (.Y(_07750_),
    .A(_04230_),
    .B(_07748_));
 sg13g2_nor2_1 _16168_ (.A(_07747_),
    .B(_07750_),
    .Y(_07751_));
 sg13g2_o21ai_1 _16169_ (.B1(_07674_),
    .Y(_07752_),
    .A1(_07657_),
    .A2(_07675_));
 sg13g2_xor2_1 _16170_ (.B(_07752_),
    .A(_07739_),
    .X(_07753_));
 sg13g2_inv_1 _16171_ (.Y(_07754_),
    .A(_07753_));
 sg13g2_a21oi_1 _16172_ (.A1(\TRNG.hash[145] ),
    .A2(_07754_),
    .Y(_07755_),
    .B1(_07677_));
 sg13g2_a21oi_1 _16173_ (.A1(_04231_),
    .A2(_07753_),
    .Y(_07756_),
    .B1(_07755_));
 sg13g2_a21oi_1 _16174_ (.A1(\TRNG.hash[147] ),
    .A2(_07745_),
    .Y(_07757_),
    .B1(_07749_));
 sg13g2_a21oi_1 _16175_ (.A1(_04229_),
    .A2(_07744_),
    .Y(_07758_),
    .B1(_07757_));
 sg13g2_a21oi_1 _16176_ (.A1(_07751_),
    .A2(_07756_),
    .Y(_07759_),
    .B1(_07758_));
 sg13g2_inv_1 _16177_ (.Y(_07760_),
    .A(_07759_));
 sg13g2_xnor2_1 _16178_ (.Y(_07761_),
    .A(\TRNG.hash[145] ),
    .B(_07753_));
 sg13g2_nand2b_1 _16179_ (.Y(_07762_),
    .B(_07761_),
    .A_N(_07678_));
 sg13g2_nor3_2 _16180_ (.A(_07747_),
    .B(_07750_),
    .C(_07762_),
    .Y(_07763_));
 sg13g2_a21oi_1 _16181_ (.A1(_07649_),
    .A2(_07763_),
    .Y(_07764_),
    .B1(_07760_));
 sg13g2_a21o_1 _16182_ (.A2(_07763_),
    .A1(_07649_),
    .B1(_07760_),
    .X(_07765_));
 sg13g2_nor2_1 _16183_ (.A(_07723_),
    .B(_07732_),
    .Y(_07766_));
 sg13g2_and2_1 _16184_ (.A(_07740_),
    .B(_07766_),
    .X(_07767_));
 sg13g2_o21ai_1 _16185_ (.B1(_07767_),
    .Y(_07768_),
    .A1(_07654_),
    .A2(_07656_));
 sg13g2_nand2b_1 _16186_ (.Y(_07769_),
    .B(_07766_),
    .A_N(_07738_));
 sg13g2_nand2b_1 _16187_ (.Y(_07770_),
    .B(_07731_),
    .A_N(_07721_));
 sg13g2_and3_2 _16188_ (.X(_07771_),
    .A(_07722_),
    .B(_07769_),
    .C(_07770_));
 sg13g2_nand2_1 _16189_ (.Y(_07772_),
    .A(_07768_),
    .B(_07771_));
 sg13g2_a21oi_2 _16190_ (.B1(_07712_),
    .Y(_07773_),
    .A2(_07715_),
    .A1(_07713_));
 sg13g2_a21oi_2 _16191_ (.B1(_07709_),
    .Y(_07774_),
    .A2(_07710_),
    .A1(\TRNG.hash[19] ));
 sg13g2_and2_1 _16192_ (.A(\TRNG.sha256.W[20] ),
    .B(\TRNG.sha256.K[20] ),
    .X(_07775_));
 sg13g2_xor2_1 _16193_ (.B(\TRNG.sha256.K[20] ),
    .A(\TRNG.sha256.W[20] ),
    .X(_07776_));
 sg13g2_xnor2_1 _16194_ (.Y(_07777_),
    .A(\TRNG.hash[20] ),
    .B(_07776_));
 sg13g2_nor2_1 _16195_ (.A(_07774_),
    .B(_07777_),
    .Y(_07778_));
 sg13g2_xor2_1 _16196_ (.B(_07777_),
    .A(_07774_),
    .X(_07779_));
 sg13g2_xnor2_1 _16197_ (.Y(_07780_),
    .A(\TRNG.hash[122] ),
    .B(\TRNG.hash[109] ));
 sg13g2_xnor2_1 _16198_ (.Y(_07781_),
    .A(\TRNG.hash[127] ),
    .B(_07780_));
 sg13g2_xnor2_1 _16199_ (.Y(_07782_),
    .A(_07779_),
    .B(_07781_));
 sg13g2_nor2_1 _16200_ (.A(_07773_),
    .B(_07782_),
    .Y(_07783_));
 sg13g2_xor2_1 _16201_ (.B(_07782_),
    .A(_07773_),
    .X(_07784_));
 sg13g2_mux2_1 _16202_ (.A0(_00169_),
    .A1(_00186_),
    .S(net5890),
    .X(_07785_));
 sg13g2_inv_1 _16203_ (.Y(_07786_),
    .A(_07785_));
 sg13g2_and2_1 _16204_ (.A(_07784_),
    .B(_07786_),
    .X(_07787_));
 sg13g2_xnor2_1 _16205_ (.Y(_07788_),
    .A(_07784_),
    .B(_07786_));
 sg13g2_a21oi_2 _16206_ (.B1(_07717_),
    .Y(_07789_),
    .A2(_07719_),
    .A1(_07718_));
 sg13g2_nor2_1 _16207_ (.A(_07788_),
    .B(_07789_),
    .Y(_07790_));
 sg13g2_xnor2_1 _16208_ (.Y(_07791_),
    .A(_07788_),
    .B(_07789_));
 sg13g2_inv_1 _16209_ (.Y(_07792_),
    .A(_07791_));
 sg13g2_xnor2_1 _16210_ (.Y(_07793_),
    .A(_07772_),
    .B(_07792_));
 sg13g2_xor2_1 _16211_ (.B(_07793_),
    .A(\TRNG.hash[148] ),
    .X(_07794_));
 sg13g2_xnor2_1 _16212_ (.Y(_07795_),
    .A(_07764_),
    .B(_07794_));
 sg13g2_or4_2 _16213_ (.A(net5544),
    .B(net5545),
    .C(net5546),
    .D(_07681_),
    .X(_07796_));
 sg13g2_xor2_1 _16214_ (.B(_07796_),
    .A(net3183),
    .X(_07797_));
 sg13g2_o21ai_1 _16215_ (.B1(net4975),
    .Y(_07798_),
    .A1(net5890),
    .A2(net5176));
 sg13g2_a221oi_1 _16216_ (.B2(net5186),
    .C1(_07798_),
    .B1(_07797_),
    .A1(net5835),
    .Y(_00543_),
    .A2(_07795_));
 sg13g2_a21oi_2 _16217_ (.B1(_07778_),
    .Y(_07799_),
    .A2(_07781_),
    .A1(_07779_));
 sg13g2_a21oi_1 _16218_ (.A1(\TRNG.hash[20] ),
    .A2(_07776_),
    .Y(_07800_),
    .B1(_07775_));
 sg13g2_and2_1 _16219_ (.A(\TRNG.sha256.W[21] ),
    .B(\TRNG.sha256.K[21] ),
    .X(_07801_));
 sg13g2_xor2_1 _16220_ (.B(\TRNG.sha256.K[21] ),
    .A(\TRNG.sha256.W[21] ),
    .X(_07802_));
 sg13g2_xnor2_1 _16221_ (.Y(_07803_),
    .A(\TRNG.hash[21] ),
    .B(_07802_));
 sg13g2_nor2_1 _16222_ (.A(_07800_),
    .B(_07803_),
    .Y(_07804_));
 sg13g2_xor2_1 _16223_ (.B(_07803_),
    .A(_07800_),
    .X(_07805_));
 sg13g2_xnor2_1 _16224_ (.Y(_07806_),
    .A(net5555),
    .B(\TRNG.hash[123] ));
 sg13g2_xnor2_1 _16225_ (.Y(_07807_),
    .A(\TRNG.hash[110] ),
    .B(_07806_));
 sg13g2_xnor2_1 _16226_ (.Y(_07808_),
    .A(_07805_),
    .B(_07807_));
 sg13g2_or2_1 _16227_ (.X(_07809_),
    .B(_07808_),
    .A(_07799_));
 sg13g2_and2_1 _16228_ (.A(_07799_),
    .B(_07808_),
    .X(_07810_));
 sg13g2_xor2_1 _16229_ (.B(_07808_),
    .A(_07799_),
    .X(_07811_));
 sg13g2_mux2_1 _16230_ (.A0(_00212_),
    .A1(_00213_),
    .S(net5889),
    .X(_07812_));
 sg13g2_xnor2_1 _16231_ (.Y(_07813_),
    .A(_07811_),
    .B(_07812_));
 sg13g2_or3_1 _16232_ (.A(_07783_),
    .B(_07787_),
    .C(_07813_),
    .X(_07814_));
 sg13g2_o21ai_1 _16233_ (.B1(_07813_),
    .Y(_07815_),
    .A1(_07783_),
    .A2(_07787_));
 sg13g2_nand2_1 _16234_ (.Y(_07816_),
    .A(_07814_),
    .B(_07815_));
 sg13g2_a21oi_1 _16235_ (.A1(_07772_),
    .A2(_07792_),
    .Y(_07817_),
    .B1(_07790_));
 sg13g2_xnor2_1 _16236_ (.Y(_07818_),
    .A(_07816_),
    .B(_07817_));
 sg13g2_inv_1 _16237_ (.Y(_07819_),
    .A(_07818_));
 sg13g2_xor2_1 _16238_ (.B(_07818_),
    .A(_00139_),
    .X(_07820_));
 sg13g2_nor2b_1 _16239_ (.A(_07794_),
    .B_N(_07820_),
    .Y(_07821_));
 sg13g2_inv_1 _16240_ (.Y(_07822_),
    .A(_07821_));
 sg13g2_nor2_1 _16241_ (.A(net3482),
    .B(_07793_),
    .Y(_07823_));
 sg13g2_nor2_1 _16242_ (.A(_07820_),
    .B(_07823_),
    .Y(_07824_));
 sg13g2_o21ai_1 _16243_ (.B1(_07824_),
    .Y(_07825_),
    .A1(_07764_),
    .A2(_07794_));
 sg13g2_nand2_1 _16244_ (.Y(_07826_),
    .A(_07820_),
    .B(_07823_));
 sg13g2_inv_1 _16245_ (.Y(_07827_),
    .A(_07826_));
 sg13g2_a221oi_1 _16246_ (.B2(_07820_),
    .C1(net5488),
    .B1(_07823_),
    .A1(_07765_),
    .Y(_07828_),
    .A2(_07821_));
 sg13g2_nand3_1 _16247_ (.B(net5890),
    .C(_07796_),
    .A(net5889),
    .Y(_07829_));
 sg13g2_a21o_1 _16248_ (.A2(_07796_),
    .A1(net5890),
    .B1(net5889),
    .X(_07830_));
 sg13g2_a21o_1 _16249_ (.A2(_07830_),
    .A1(_07829_),
    .B1(_04228_),
    .X(_07831_));
 sg13g2_a22oi_1 _16250_ (.Y(_07832_),
    .B1(_07831_),
    .B2(net5488),
    .A2(_07828_),
    .A1(_07825_));
 sg13g2_o21ai_1 _16251_ (.B1(net4975),
    .Y(_07833_),
    .A1(net5889),
    .A2(net5176));
 sg13g2_nor2_1 _16252_ (.A(_07832_),
    .B(_07833_),
    .Y(_00544_));
 sg13g2_a21oi_1 _16253_ (.A1(\TRNG.hash[149] ),
    .A2(_07819_),
    .Y(_07834_),
    .B1(_07827_));
 sg13g2_a221oi_1 _16254_ (.B2(_07765_),
    .C1(_07827_),
    .B1(_07821_),
    .A1(\TRNG.hash[149] ),
    .Y(_07835_),
    .A2(_07819_));
 sg13g2_a21oi_1 _16255_ (.A1(_07805_),
    .A2(_07807_),
    .Y(_07836_),
    .B1(_07804_));
 sg13g2_a21oi_2 _16256_ (.B1(_07801_),
    .Y(_07837_),
    .A2(_07802_),
    .A1(\TRNG.hash[21] ));
 sg13g2_and2_1 _16257_ (.A(\TRNG.sha256.W[22] ),
    .B(\TRNG.sha256.K[22] ),
    .X(_07838_));
 sg13g2_xor2_1 _16258_ (.B(\TRNG.sha256.K[22] ),
    .A(\TRNG.sha256.W[22] ),
    .X(_07839_));
 sg13g2_xnor2_1 _16259_ (.Y(_07840_),
    .A(\TRNG.hash[22] ),
    .B(_07839_));
 sg13g2_nor2_1 _16260_ (.A(_07837_),
    .B(_07840_),
    .Y(_07841_));
 sg13g2_xor2_1 _16261_ (.B(_07840_),
    .A(_07837_),
    .X(_07842_));
 sg13g2_xnor2_1 _16262_ (.Y(_07843_),
    .A(net5554),
    .B(\TRNG.hash[111] ));
 sg13g2_xnor2_1 _16263_ (.Y(_07844_),
    .A(\TRNG.hash[124] ),
    .B(_07843_));
 sg13g2_xnor2_1 _16264_ (.Y(_07845_),
    .A(_07842_),
    .B(_07844_));
 sg13g2_or2_1 _16265_ (.X(_07846_),
    .B(_07845_),
    .A(_07836_));
 sg13g2_and2_1 _16266_ (.A(_07836_),
    .B(_07845_),
    .X(_07847_));
 sg13g2_xnor2_1 _16267_ (.Y(_07848_),
    .A(_07836_),
    .B(_07845_));
 sg13g2_mux2_1 _16268_ (.A0(_00177_),
    .A1(_00187_),
    .S(\TRNG.hash[118] ),
    .X(_07849_));
 sg13g2_xnor2_1 _16269_ (.Y(_07850_),
    .A(_07848_),
    .B(_07849_));
 sg13g2_o21ai_1 _16270_ (.B1(_07809_),
    .Y(_07851_),
    .A1(_07810_),
    .A2(_07812_));
 sg13g2_nand2b_1 _16271_ (.Y(_07852_),
    .B(_07851_),
    .A_N(_07850_));
 sg13g2_xor2_1 _16272_ (.B(_07851_),
    .A(_07850_),
    .X(_07853_));
 sg13g2_nor2_1 _16273_ (.A(_07791_),
    .B(_07816_),
    .Y(_07854_));
 sg13g2_nand2_1 _16274_ (.Y(_07855_),
    .A(_07790_),
    .B(_07814_));
 sg13g2_nand2_1 _16275_ (.Y(_07856_),
    .A(_07815_),
    .B(_07855_));
 sg13g2_a21oi_1 _16276_ (.A1(_07772_),
    .A2(_07854_),
    .Y(_07857_),
    .B1(_07856_));
 sg13g2_xnor2_1 _16277_ (.Y(_07858_),
    .A(_07853_),
    .B(_07857_));
 sg13g2_xor2_1 _16278_ (.B(_07858_),
    .A(\TRNG.hash[150] ),
    .X(_07859_));
 sg13g2_xnor2_1 _16279_ (.Y(_07860_),
    .A(_07835_),
    .B(_07859_));
 sg13g2_nor2_1 _16280_ (.A(_04293_),
    .B(_07829_),
    .Y(_07861_));
 sg13g2_xnor2_1 _16281_ (.Y(_07862_),
    .A(\TRNG.hash[118] ),
    .B(_07829_));
 sg13g2_o21ai_1 _16282_ (.B1(net4975),
    .Y(_07863_),
    .A1(net5180),
    .A2(_07862_));
 sg13g2_a221oi_1 _16283_ (.B2(net5834),
    .C1(_07863_),
    .B1(_07860_),
    .A1(_04293_),
    .Y(_00545_),
    .A2(net5352));
 sg13g2_a21o_1 _16284_ (.A2(_07861_),
    .A1(net5574),
    .B1(\TRNG.hash[119] ),
    .X(_07864_));
 sg13g2_and2_1 _16285_ (.A(\TRNG.hash[119] ),
    .B(_07861_),
    .X(_07865_));
 sg13g2_a21oi_1 _16286_ (.A1(net5574),
    .A2(_07865_),
    .Y(_07866_),
    .B1(net5853));
 sg13g2_o21ai_1 _16287_ (.B1(_07852_),
    .Y(_07867_),
    .A1(_07853_),
    .A2(_07857_));
 sg13g2_o21ai_1 _16288_ (.B1(_07846_),
    .Y(_07868_),
    .A1(_07847_),
    .A2(_07849_));
 sg13g2_a21oi_1 _16289_ (.A1(_07842_),
    .A2(_07844_),
    .Y(_07869_),
    .B1(_07841_));
 sg13g2_a21oi_2 _16290_ (.B1(_07838_),
    .Y(_07870_),
    .A2(_07839_),
    .A1(\TRNG.hash[22] ));
 sg13g2_and2_1 _16291_ (.A(\TRNG.sha256.W[23] ),
    .B(\TRNG.sha256.K[23] ),
    .X(_07871_));
 sg13g2_xor2_1 _16292_ (.B(\TRNG.sha256.K[23] ),
    .A(\TRNG.sha256.W[23] ),
    .X(_07872_));
 sg13g2_xnor2_1 _16293_ (.Y(_07873_),
    .A(\TRNG.hash[23] ),
    .B(_07872_));
 sg13g2_nor2_1 _16294_ (.A(_07870_),
    .B(_07873_),
    .Y(_07874_));
 sg13g2_xor2_1 _16295_ (.B(_07873_),
    .A(_07870_),
    .X(_07875_));
 sg13g2_xnor2_1 _16296_ (.Y(_07876_),
    .A(\TRNG.hash[125] ),
    .B(net5891));
 sg13g2_xnor2_1 _16297_ (.Y(_07877_),
    .A(net5553),
    .B(_07876_));
 sg13g2_xnor2_1 _16298_ (.Y(_07878_),
    .A(_07875_),
    .B(_07877_));
 sg13g2_or2_1 _16299_ (.X(_07879_),
    .B(_07878_),
    .A(_07869_));
 sg13g2_xnor2_1 _16300_ (.Y(_07880_),
    .A(_07869_),
    .B(_07878_));
 sg13g2_mux2_1 _16301_ (.A0(_00172_),
    .A1(_00214_),
    .S(\TRNG.hash[119] ),
    .X(_07881_));
 sg13g2_xor2_1 _16302_ (.B(_07881_),
    .A(_07880_),
    .X(_07882_));
 sg13g2_nor2_1 _16303_ (.A(_07868_),
    .B(_07882_),
    .Y(_07883_));
 sg13g2_nand2_1 _16304_ (.Y(_07884_),
    .A(_07868_),
    .B(_07882_));
 sg13g2_nand2b_1 _16305_ (.Y(_07885_),
    .B(_07884_),
    .A_N(_07883_));
 sg13g2_xnor2_1 _16306_ (.Y(_07886_),
    .A(_07867_),
    .B(_07885_));
 sg13g2_nor2_1 _16307_ (.A(\TRNG.hash[151] ),
    .B(_07886_),
    .Y(_07887_));
 sg13g2_xnor2_1 _16308_ (.Y(_07888_),
    .A(\TRNG.hash[151] ),
    .B(_07886_));
 sg13g2_or2_1 _16309_ (.X(_07889_),
    .B(_07858_),
    .A(_00140_));
 sg13g2_o21ai_1 _16310_ (.B1(_07889_),
    .Y(_07890_),
    .A1(_07835_),
    .A2(_07859_));
 sg13g2_xnor2_1 _16311_ (.Y(_07891_),
    .A(_07888_),
    .B(_07890_));
 sg13g2_a22oi_1 _16312_ (.Y(_07892_),
    .B1(_07891_),
    .B2(net5853),
    .A2(_07866_),
    .A1(_07864_));
 sg13g2_nor2_1 _16313_ (.A(net4968),
    .B(_07892_),
    .Y(_00546_));
 sg13g2_a21oi_1 _16314_ (.A1(_07875_),
    .A2(_07877_),
    .Y(_07893_),
    .B1(_07874_));
 sg13g2_a21oi_1 _16315_ (.A1(\TRNG.hash[23] ),
    .A2(_07872_),
    .Y(_07894_),
    .B1(_07871_));
 sg13g2_and2_1 _16316_ (.A(\TRNG.sha256.W[24] ),
    .B(\TRNG.sha256.K[24] ),
    .X(_07895_));
 sg13g2_xor2_1 _16317_ (.B(\TRNG.sha256.K[24] ),
    .A(\TRNG.sha256.W[24] ),
    .X(_07896_));
 sg13g2_xnor2_1 _16318_ (.Y(_07897_),
    .A(\TRNG.hash[24] ),
    .B(_07896_));
 sg13g2_nor2_1 _16319_ (.A(_07894_),
    .B(_07897_),
    .Y(_07898_));
 sg13g2_xor2_1 _16320_ (.B(_07897_),
    .A(_07894_),
    .X(_07899_));
 sg13g2_xnor2_1 _16321_ (.Y(_07900_),
    .A(net5546),
    .B(net5552));
 sg13g2_xnor2_1 _16322_ (.Y(_07901_),
    .A(\TRNG.hash[126] ),
    .B(_07900_));
 sg13g2_xnor2_1 _16323_ (.Y(_07902_),
    .A(_07899_),
    .B(_07901_));
 sg13g2_nor2_1 _16324_ (.A(_07893_),
    .B(_07902_),
    .Y(_07903_));
 sg13g2_xor2_1 _16325_ (.B(_07902_),
    .A(_07893_),
    .X(_07904_));
 sg13g2_mux2_1 _16326_ (.A0(\TRNG.hash[56] ),
    .A1(\TRNG.hash[88] ),
    .S(\TRNG.hash[120] ),
    .X(_07905_));
 sg13g2_a21oi_2 _16327_ (.B1(_07903_),
    .Y(_07906_),
    .A2(_07905_),
    .A1(_07904_));
 sg13g2_a21oi_1 _16328_ (.A1(_07899_),
    .A2(_07901_),
    .Y(_07907_),
    .B1(_07898_));
 sg13g2_a21oi_1 _16329_ (.A1(\TRNG.hash[24] ),
    .A2(_07896_),
    .Y(_07908_),
    .B1(_07895_));
 sg13g2_and2_1 _16330_ (.A(\TRNG.sha256.W[25] ),
    .B(\TRNG.sha256.K[25] ),
    .X(_07909_));
 sg13g2_xor2_1 _16331_ (.B(\TRNG.sha256.K[25] ),
    .A(\TRNG.sha256.W[25] ),
    .X(_07910_));
 sg13g2_xnor2_1 _16332_ (.Y(_07911_),
    .A(\TRNG.hash[25] ),
    .B(_07910_));
 sg13g2_nor2_1 _16333_ (.A(_07908_),
    .B(_07911_),
    .Y(_07912_));
 sg13g2_xor2_1 _16334_ (.B(_07911_),
    .A(_07908_),
    .X(_07913_));
 sg13g2_xnor2_1 _16335_ (.Y(_07914_),
    .A(net5551),
    .B(\TRNG.hash[127] ));
 sg13g2_xnor2_1 _16336_ (.Y(_07915_),
    .A(net5545),
    .B(_07914_));
 sg13g2_xnor2_1 _16337_ (.Y(_07916_),
    .A(_07913_),
    .B(_07915_));
 sg13g2_or2_1 _16338_ (.X(_07917_),
    .B(_07916_),
    .A(_07907_));
 sg13g2_xnor2_1 _16339_ (.Y(_07918_),
    .A(_07907_),
    .B(_07916_));
 sg13g2_mux2_1 _16340_ (.A0(_00216_),
    .A1(_00217_),
    .S(\TRNG.hash[121] ),
    .X(_07919_));
 sg13g2_xnor2_1 _16341_ (.Y(_07920_),
    .A(_07918_),
    .B(_07919_));
 sg13g2_nor2_1 _16342_ (.A(_07906_),
    .B(_07920_),
    .Y(_07921_));
 sg13g2_xor2_1 _16343_ (.B(_07920_),
    .A(_07906_),
    .X(_07922_));
 sg13g2_xnor2_1 _16344_ (.Y(_07923_),
    .A(_07904_),
    .B(_07905_));
 sg13g2_o21ai_1 _16345_ (.B1(_07879_),
    .Y(_07924_),
    .A1(_07880_),
    .A2(_07881_));
 sg13g2_nor2b_1 _16346_ (.A(_07923_),
    .B_N(_07924_),
    .Y(_07925_));
 sg13g2_xor2_1 _16347_ (.B(_07924_),
    .A(_07923_),
    .X(_07926_));
 sg13g2_inv_1 _16348_ (.Y(_07927_),
    .A(_07926_));
 sg13g2_nor2_1 _16349_ (.A(_07853_),
    .B(_07885_),
    .Y(_07928_));
 sg13g2_nand2_1 _16350_ (.Y(_07929_),
    .A(_07854_),
    .B(_07928_));
 sg13g2_a21oi_2 _16351_ (.B1(_07929_),
    .Y(_07930_),
    .A2(_07771_),
    .A1(_07768_));
 sg13g2_o21ai_1 _16352_ (.B1(_07884_),
    .Y(_07931_),
    .A1(_07852_),
    .A2(_07883_));
 sg13g2_a21o_1 _16353_ (.A2(_07928_),
    .A1(_07856_),
    .B1(_07931_),
    .X(_07932_));
 sg13g2_nor2_1 _16354_ (.A(_07930_),
    .B(_07932_),
    .Y(_07933_));
 sg13g2_nor2_2 _16355_ (.A(_07926_),
    .B(_07933_),
    .Y(_07934_));
 sg13g2_o21ai_1 _16356_ (.B1(_07927_),
    .Y(_07935_),
    .A1(_07930_),
    .A2(_07932_));
 sg13g2_nor2_1 _16357_ (.A(_07925_),
    .B(_07934_),
    .Y(_07936_));
 sg13g2_xnor2_1 _16358_ (.Y(_07937_),
    .A(_07922_),
    .B(_07936_));
 sg13g2_nor2_1 _16359_ (.A(\TRNG.hash[153] ),
    .B(_07937_),
    .Y(_07938_));
 sg13g2_inv_1 _16360_ (.Y(_07939_),
    .A(_07938_));
 sg13g2_nor3_2 _16361_ (.A(_07927_),
    .B(_07930_),
    .C(_07932_),
    .Y(_07940_));
 sg13g2_nor2_2 _16362_ (.A(_07934_),
    .B(_07940_),
    .Y(_07941_));
 sg13g2_nor3_1 _16363_ (.A(_00141_),
    .B(_07934_),
    .C(_07940_),
    .Y(_07942_));
 sg13g2_nor2_1 _16364_ (.A(_07859_),
    .B(_07888_),
    .Y(_07943_));
 sg13g2_o21ai_1 _16365_ (.B1(_07834_),
    .Y(_07944_),
    .A1(_07759_),
    .A2(_07822_));
 sg13g2_a22oi_1 _16366_ (.Y(_07945_),
    .B1(_07943_),
    .B2(_07944_),
    .A2(_07886_),
    .A1(\TRNG.hash[151] ));
 sg13g2_o21ai_1 _16367_ (.B1(_07945_),
    .Y(_07946_),
    .A1(_07887_),
    .A2(_07889_));
 sg13g2_nand3_1 _16368_ (.B(_07821_),
    .C(_07943_),
    .A(_07763_),
    .Y(_07947_));
 sg13g2_a21oi_1 _16369_ (.A1(_07634_),
    .A2(_07643_),
    .Y(_07948_),
    .B1(_07947_));
 sg13g2_nor2_1 _16370_ (.A(_07946_),
    .B(_07948_),
    .Y(_07949_));
 sg13g2_xor2_1 _16371_ (.B(_07941_),
    .A(\TRNG.hash[152] ),
    .X(_07950_));
 sg13g2_o21ai_1 _16372_ (.B1(_07950_),
    .Y(_07951_),
    .A1(_07946_),
    .A2(_07948_));
 sg13g2_nor2b_1 _16373_ (.A(_07942_),
    .B_N(_07951_),
    .Y(_07952_));
 sg13g2_and2_1 _16374_ (.A(\TRNG.hash[153] ),
    .B(_07937_),
    .X(_07953_));
 sg13g2_nor2_1 _16375_ (.A(_07938_),
    .B(_07953_),
    .Y(_07954_));
 sg13g2_xor2_1 _16376_ (.B(_07954_),
    .A(_07952_),
    .X(_07955_));
 sg13g2_nor2b_1 _16377_ (.A(_07865_),
    .B_N(_00215_),
    .Y(_07956_));
 sg13g2_xnor2_1 _16378_ (.Y(_07957_),
    .A(net3591),
    .B(_07956_));
 sg13g2_o21ai_1 _16379_ (.B1(net4975),
    .Y(_07958_),
    .A1(\TRNG.hash[121] ),
    .A2(net5176));
 sg13g2_a221oi_1 _16380_ (.B2(net5186),
    .C1(_07958_),
    .B1(net3592),
    .A1(net5850),
    .Y(_00547_),
    .A2(_07955_));
 sg13g2_o21ai_1 _16381_ (.B1(_07939_),
    .Y(_07959_),
    .A1(_07942_),
    .A2(_07953_));
 sg13g2_o21ai_1 _16382_ (.B1(_07959_),
    .Y(_07960_),
    .A1(_07938_),
    .A2(_07951_));
 sg13g2_a21oi_1 _16383_ (.A1(_07913_),
    .A2(_07915_),
    .Y(_07961_),
    .B1(_07912_));
 sg13g2_a21oi_2 _16384_ (.B1(_07909_),
    .Y(_07962_),
    .A2(_07910_),
    .A1(\TRNG.hash[25] ));
 sg13g2_and2_1 _16385_ (.A(\TRNG.sha256.W[26] ),
    .B(\TRNG.sha256.K[26] ),
    .X(_07963_));
 sg13g2_xor2_1 _16386_ (.B(\TRNG.sha256.K[26] ),
    .A(\TRNG.sha256.W[26] ),
    .X(_07964_));
 sg13g2_xnor2_1 _16387_ (.Y(_07965_),
    .A(\TRNG.hash[26] ),
    .B(_07964_));
 sg13g2_nor2_1 _16388_ (.A(_07962_),
    .B(_07965_),
    .Y(_07966_));
 sg13g2_xor2_1 _16389_ (.B(_07965_),
    .A(_07962_),
    .X(_07967_));
 sg13g2_xnor2_1 _16390_ (.Y(_07968_),
    .A(net5550),
    .B(net5555));
 sg13g2_xnor2_1 _16391_ (.Y(_07969_),
    .A(net5544),
    .B(_07968_));
 sg13g2_xnor2_1 _16392_ (.Y(_07970_),
    .A(_07967_),
    .B(_07969_));
 sg13g2_nor2_1 _16393_ (.A(_07961_),
    .B(_07970_),
    .Y(_07971_));
 sg13g2_xor2_1 _16394_ (.B(_07970_),
    .A(_07961_),
    .X(_07972_));
 sg13g2_inv_1 _16395_ (.Y(_07973_),
    .A(_07972_));
 sg13g2_mux2_1 _16396_ (.A0(_00218_),
    .A1(_00188_),
    .S(\TRNG.hash[122] ),
    .X(_07974_));
 sg13g2_nor2_1 _16397_ (.A(_07973_),
    .B(_07974_),
    .Y(_07975_));
 sg13g2_xnor2_1 _16398_ (.Y(_07976_),
    .A(_07972_),
    .B(_07974_));
 sg13g2_o21ai_1 _16399_ (.B1(_07917_),
    .Y(_07977_),
    .A1(_07918_),
    .A2(_07919_));
 sg13g2_xnor2_1 _16400_ (.Y(_07978_),
    .A(_07976_),
    .B(_07977_));
 sg13g2_nor2_1 _16401_ (.A(_07921_),
    .B(_07925_),
    .Y(_07979_));
 sg13g2_a22oi_1 _16402_ (.Y(_07980_),
    .B1(_07935_),
    .B2(_07979_),
    .A2(_07920_),
    .A1(_07906_));
 sg13g2_a221oi_1 _16403_ (.B2(_07979_),
    .C1(_07978_),
    .B1(_07935_),
    .A1(_07906_),
    .Y(_07981_),
    .A2(_07920_));
 sg13g2_xnor2_1 _16404_ (.Y(_07982_),
    .A(_07978_),
    .B(_07980_));
 sg13g2_xnor2_1 _16405_ (.Y(_07983_),
    .A(\TRNG.hash[154] ),
    .B(_07982_));
 sg13g2_inv_1 _16406_ (.Y(_07984_),
    .A(_07983_));
 sg13g2_xnor2_1 _16407_ (.Y(_07985_),
    .A(_07960_),
    .B(_07984_));
 sg13g2_nor2_1 _16408_ (.A(\TRNG.hash[120] ),
    .B(_07865_),
    .Y(_07986_));
 sg13g2_nor2b_2 _16409_ (.A(_07986_),
    .B_N(\TRNG.hash[121] ),
    .Y(_07987_));
 sg13g2_xor2_1 _16410_ (.B(_07987_),
    .A(net3659),
    .X(_07988_));
 sg13g2_o21ai_1 _16411_ (.B1(net4975),
    .Y(_07989_),
    .A1(\TRNG.hash[122] ),
    .A2(net5176));
 sg13g2_a221oi_1 _16412_ (.B2(net5186),
    .C1(_07989_),
    .B1(_07988_),
    .A1(net5850),
    .Y(_00548_),
    .A2(_07985_));
 sg13g2_nor2b_1 _16413_ (.A(_00143_),
    .B_N(_07982_),
    .Y(_07990_));
 sg13g2_inv_1 _16414_ (.Y(_07991_),
    .A(_07990_));
 sg13g2_a21oi_1 _16415_ (.A1(_07960_),
    .A2(_07984_),
    .Y(_07992_),
    .B1(_07990_));
 sg13g2_a21oi_2 _16416_ (.B1(_07966_),
    .Y(_07993_),
    .A2(_07969_),
    .A1(_07967_));
 sg13g2_a21oi_2 _16417_ (.B1(_07963_),
    .Y(_07994_),
    .A2(_07964_),
    .A1(\TRNG.hash[26] ));
 sg13g2_and2_1 _16418_ (.A(\TRNG.sha256.W[27] ),
    .B(\TRNG.sha256.K[27] ),
    .X(_07995_));
 sg13g2_xor2_1 _16419_ (.B(\TRNG.sha256.K[27] ),
    .A(\TRNG.sha256.W[27] ),
    .X(_07996_));
 sg13g2_xnor2_1 _16420_ (.Y(_07997_),
    .A(\TRNG.hash[27] ),
    .B(_07996_));
 sg13g2_nor2_1 _16421_ (.A(_07994_),
    .B(_07997_),
    .Y(_07998_));
 sg13g2_xor2_1 _16422_ (.B(_07997_),
    .A(_07994_),
    .X(_07999_));
 sg13g2_xnor2_1 _16423_ (.Y(_08000_),
    .A(net5554),
    .B(net5890));
 sg13g2_xnor2_1 _16424_ (.Y(_08001_),
    .A(\TRNG.hash[102] ),
    .B(_08000_));
 sg13g2_xnor2_1 _16425_ (.Y(_08002_),
    .A(_07999_),
    .B(_08001_));
 sg13g2_or2_1 _16426_ (.X(_08003_),
    .B(_08002_),
    .A(_07993_));
 sg13g2_and2_1 _16427_ (.A(_07993_),
    .B(_08002_),
    .X(_08004_));
 sg13g2_xor2_1 _16428_ (.B(_08002_),
    .A(_07993_),
    .X(_08005_));
 sg13g2_mux2_1 _16429_ (.A0(_00219_),
    .A1(_00190_),
    .S(\TRNG.hash[123] ),
    .X(_08006_));
 sg13g2_xnor2_1 _16430_ (.Y(_08007_),
    .A(_08005_),
    .B(_08006_));
 sg13g2_nor3_1 _16431_ (.A(_07971_),
    .B(_07975_),
    .C(_08007_),
    .Y(_08008_));
 sg13g2_o21ai_1 _16432_ (.B1(_08007_),
    .Y(_08009_),
    .A1(_07971_),
    .A2(_07975_));
 sg13g2_nand2b_1 _16433_ (.Y(_08010_),
    .B(_08009_),
    .A_N(_08008_));
 sg13g2_a21oi_1 _16434_ (.A1(_07976_),
    .A2(_07977_),
    .Y(_08011_),
    .B1(_07981_));
 sg13g2_xnor2_1 _16435_ (.Y(_08012_),
    .A(_08010_),
    .B(_08011_));
 sg13g2_inv_1 _16436_ (.Y(_08013_),
    .A(_08012_));
 sg13g2_xor2_1 _16437_ (.B(_08012_),
    .A(_00142_),
    .X(_08014_));
 sg13g2_o21ai_1 _16438_ (.B1(net5835),
    .Y(_08015_),
    .A1(_07992_),
    .A2(_08014_));
 sg13g2_a21oi_2 _16439_ (.B1(_08015_),
    .Y(_08016_),
    .A2(_08014_),
    .A1(_07992_));
 sg13g2_nand3_1 _16440_ (.B(\TRNG.hash[122] ),
    .C(_07987_),
    .A(\TRNG.hash[123] ),
    .Y(_08017_));
 sg13g2_inv_1 _16441_ (.Y(_08018_),
    .A(_08017_));
 sg13g2_a21oi_1 _16442_ (.A1(\TRNG.hash[122] ),
    .A2(_07987_),
    .Y(_08019_),
    .B1(\TRNG.hash[123] ));
 sg13g2_o21ai_1 _16443_ (.B1(net5186),
    .Y(_08020_),
    .A1(_08018_),
    .A2(_08019_));
 sg13g2_o21ai_1 _16444_ (.B1(_08020_),
    .Y(_08021_),
    .A1(\TRNG.hash[123] ),
    .A2(net5176));
 sg13g2_nor3_1 _16445_ (.A(net4967),
    .B(_08016_),
    .C(_08021_),
    .Y(_00549_));
 sg13g2_o21ai_1 _16446_ (.B1(_08003_),
    .Y(_08022_),
    .A1(_08004_),
    .A2(_08006_));
 sg13g2_a21oi_1 _16447_ (.A1(_07999_),
    .A2(_08001_),
    .Y(_08023_),
    .B1(_07998_));
 sg13g2_a21oi_2 _16448_ (.B1(_07995_),
    .Y(_08024_),
    .A2(_07996_),
    .A1(\TRNG.hash[27] ));
 sg13g2_and2_1 _16449_ (.A(\TRNG.sha256.W[28] ),
    .B(\TRNG.sha256.K[28] ),
    .X(_08025_));
 sg13g2_xor2_1 _16450_ (.B(\TRNG.sha256.K[28] ),
    .A(\TRNG.sha256.W[28] ),
    .X(_08026_));
 sg13g2_xnor2_1 _16451_ (.Y(_08027_),
    .A(\TRNG.hash[28] ),
    .B(_08026_));
 sg13g2_nor2_1 _16452_ (.A(_08024_),
    .B(_08027_),
    .Y(_08028_));
 sg13g2_xor2_1 _16453_ (.B(_08027_),
    .A(_08024_),
    .X(_08029_));
 sg13g2_xnor2_1 _16454_ (.Y(_08030_),
    .A(net5889),
    .B(net5897));
 sg13g2_xnor2_1 _16455_ (.Y(_08031_),
    .A(net5553),
    .B(_08030_));
 sg13g2_xnor2_1 _16456_ (.Y(_08032_),
    .A(_08029_),
    .B(_08031_));
 sg13g2_nor2_1 _16457_ (.A(_08023_),
    .B(_08032_),
    .Y(_08033_));
 sg13g2_xor2_1 _16458_ (.B(_08032_),
    .A(_08023_),
    .X(_08034_));
 sg13g2_mux2_1 _16459_ (.A0(\TRNG.hash[60] ),
    .A1(\TRNG.hash[92] ),
    .S(\TRNG.hash[124] ),
    .X(_08035_));
 sg13g2_xnor2_1 _16460_ (.Y(_08036_),
    .A(_08034_),
    .B(_08035_));
 sg13g2_inv_1 _16461_ (.Y(_08037_),
    .A(_08036_));
 sg13g2_xor2_1 _16462_ (.B(_08036_),
    .A(_08022_),
    .X(_08038_));
 sg13g2_o21ai_1 _16463_ (.B1(_08009_),
    .Y(_08039_),
    .A1(_08008_),
    .A2(_08011_));
 sg13g2_nor2b_1 _16464_ (.A(_08038_),
    .B_N(_08039_),
    .Y(_08040_));
 sg13g2_xor2_1 _16465_ (.B(_08039_),
    .A(_08038_),
    .X(_08041_));
 sg13g2_nor2_1 _16466_ (.A(_04298_),
    .B(_08041_),
    .Y(_08042_));
 sg13g2_nand4_1 _16467_ (.B(_07954_),
    .C(_07984_),
    .A(_07950_),
    .Y(_08043_),
    .D(_08014_));
 sg13g2_o21ai_1 _16468_ (.B1(_07991_),
    .Y(_08044_),
    .A1(_07959_),
    .A2(_07983_));
 sg13g2_a22oi_1 _16469_ (.Y(_08045_),
    .B1(_08014_),
    .B2(_08044_),
    .A2(_08013_),
    .A1(\TRNG.hash[155] ));
 sg13g2_o21ai_1 _16470_ (.B1(_08045_),
    .Y(_08046_),
    .A1(_07949_),
    .A2(_08043_));
 sg13g2_xnor2_1 _16471_ (.Y(_08047_),
    .A(_04298_),
    .B(_08041_));
 sg13g2_inv_1 _16472_ (.Y(_08048_),
    .A(_08047_));
 sg13g2_a21oi_1 _16473_ (.A1(_08046_),
    .A2(_08048_),
    .Y(_08049_),
    .B1(_08042_));
 sg13g2_a21oi_1 _16474_ (.A1(_08022_),
    .A2(_08037_),
    .Y(_08050_),
    .B1(_08040_));
 sg13g2_a21oi_1 _16475_ (.A1(_08034_),
    .A2(_08035_),
    .Y(_08051_),
    .B1(_08033_));
 sg13g2_a21oi_1 _16476_ (.A1(_08029_),
    .A2(_08031_),
    .Y(_08052_),
    .B1(_08028_));
 sg13g2_a21oi_1 _16477_ (.A1(\TRNG.hash[28] ),
    .A2(_08026_),
    .Y(_08053_),
    .B1(_08025_));
 sg13g2_and2_1 _16478_ (.A(\TRNG.sha256.W[29] ),
    .B(\TRNG.sha256.K[29] ),
    .X(_08054_));
 sg13g2_xor2_1 _16479_ (.B(\TRNG.sha256.K[29] ),
    .A(\TRNG.sha256.W[29] ),
    .X(_08055_));
 sg13g2_xnor2_1 _16480_ (.Y(_08056_),
    .A(\TRNG.hash[29] ),
    .B(_08055_));
 sg13g2_nor2_1 _16481_ (.A(_08053_),
    .B(_08056_),
    .Y(_08057_));
 sg13g2_xor2_1 _16482_ (.B(_08056_),
    .A(_08053_),
    .X(_08058_));
 sg13g2_xnor2_1 _16483_ (.Y(_08059_),
    .A(\TRNG.hash[118] ),
    .B(net5896));
 sg13g2_xnor2_1 _16484_ (.Y(_08060_),
    .A(net5552),
    .B(_08059_));
 sg13g2_xnor2_1 _16485_ (.Y(_08061_),
    .A(_08058_),
    .B(_08060_));
 sg13g2_or2_1 _16486_ (.X(_08062_),
    .B(_08061_),
    .A(_08052_));
 sg13g2_xnor2_1 _16487_ (.Y(_08063_),
    .A(_08052_),
    .B(_08061_));
 sg13g2_mux2_1 _16488_ (.A0(_00170_),
    .A1(_00189_),
    .S(\TRNG.hash[125] ),
    .X(_08064_));
 sg13g2_xnor2_1 _16489_ (.Y(_08065_),
    .A(_08063_),
    .B(_08064_));
 sg13g2_nor2_1 _16490_ (.A(_08051_),
    .B(_08065_),
    .Y(_08066_));
 sg13g2_xor2_1 _16491_ (.B(_08065_),
    .A(_08051_),
    .X(_08067_));
 sg13g2_nor2b_1 _16492_ (.A(_08050_),
    .B_N(_08067_),
    .Y(_08068_));
 sg13g2_xor2_1 _16493_ (.B(_08067_),
    .A(_08050_),
    .X(_08069_));
 sg13g2_xnor2_1 _16494_ (.Y(_08070_),
    .A(\TRNG.hash[157] ),
    .B(_08069_));
 sg13g2_xor2_1 _16495_ (.B(_08070_),
    .A(_08049_),
    .X(_08071_));
 sg13g2_nand2_1 _16496_ (.Y(_08072_),
    .A(_00200_),
    .B(_08017_));
 sg13g2_xor2_1 _16497_ (.B(_08072_),
    .A(net3710),
    .X(_08073_));
 sg13g2_o21ai_1 _16498_ (.B1(net4976),
    .Y(_08074_),
    .A1(\TRNG.hash[125] ),
    .A2(net5176));
 sg13g2_a221oi_1 _16499_ (.B2(net5189),
    .C1(_08074_),
    .B1(net3711),
    .A1(net5859),
    .Y(_00550_),
    .A2(_08071_));
 sg13g2_and2_1 _16500_ (.A(_08048_),
    .B(_08070_),
    .X(_08075_));
 sg13g2_nand2_1 _16501_ (.Y(_08076_),
    .A(_08042_),
    .B(_08070_));
 sg13g2_o21ai_1 _16502_ (.B1(_08076_),
    .Y(_08077_),
    .A1(_00145_),
    .A2(_08069_));
 sg13g2_a21o_1 _16503_ (.A2(_08075_),
    .A1(_08046_),
    .B1(_08077_),
    .X(_08078_));
 sg13g2_nor2_1 _16504_ (.A(_08066_),
    .B(_08068_),
    .Y(_08079_));
 sg13g2_o21ai_1 _16505_ (.B1(_08062_),
    .Y(_08080_),
    .A1(_08063_),
    .A2(_08064_));
 sg13g2_a21oi_1 _16506_ (.A1(_08058_),
    .A2(_08060_),
    .Y(_08081_),
    .B1(_08057_));
 sg13g2_a21oi_1 _16507_ (.A1(\TRNG.hash[29] ),
    .A2(_08055_),
    .Y(_08082_),
    .B1(_08054_));
 sg13g2_and2_1 _16508_ (.A(\TRNG.sha256.W[30] ),
    .B(\TRNG.sha256.K[30] ),
    .X(_08083_));
 sg13g2_xor2_1 _16509_ (.B(\TRNG.sha256.K[30] ),
    .A(\TRNG.sha256.W[30] ),
    .X(_08084_));
 sg13g2_xnor2_1 _16510_ (.Y(_08085_),
    .A(\TRNG.hash[30] ),
    .B(_08084_));
 sg13g2_nor2_1 _16511_ (.A(_08082_),
    .B(_08085_),
    .Y(_08086_));
 sg13g2_xor2_1 _16512_ (.B(_08085_),
    .A(_08082_),
    .X(_08087_));
 sg13g2_xnor2_1 _16513_ (.Y(_08088_),
    .A(net5551),
    .B(\TRNG.hash[119] ));
 sg13g2_xnor2_1 _16514_ (.Y(_08089_),
    .A(\TRNG.hash[105] ),
    .B(_08088_));
 sg13g2_xnor2_1 _16515_ (.Y(_08090_),
    .A(_08087_),
    .B(_08089_));
 sg13g2_nor2_1 _16516_ (.A(_08081_),
    .B(_08090_),
    .Y(_08091_));
 sg13g2_xor2_1 _16517_ (.B(_08090_),
    .A(_08081_),
    .X(_08092_));
 sg13g2_mux2_1 _16518_ (.A0(\TRNG.hash[62] ),
    .A1(\TRNG.hash[94] ),
    .S(\TRNG.hash[126] ),
    .X(_08093_));
 sg13g2_xor2_1 _16519_ (.B(_08093_),
    .A(_08092_),
    .X(_08094_));
 sg13g2_nand2_1 _16520_ (.Y(_08095_),
    .A(_08080_),
    .B(_08094_));
 sg13g2_xnor2_1 _16521_ (.Y(_08096_),
    .A(_08080_),
    .B(_08094_));
 sg13g2_xor2_1 _16522_ (.B(_08096_),
    .A(_08079_),
    .X(_08097_));
 sg13g2_xnor2_1 _16523_ (.Y(_08098_),
    .A(\TRNG.hash[158] ),
    .B(_08097_));
 sg13g2_inv_1 _16524_ (.Y(_08099_),
    .A(_08098_));
 sg13g2_a22oi_1 _16525_ (.Y(_08100_),
    .B1(_08099_),
    .B2(_08078_),
    .A2(_08097_),
    .A1(_04376_));
 sg13g2_o21ai_1 _16526_ (.B1(_08095_),
    .Y(_08101_),
    .A1(_08079_),
    .A2(_08096_));
 sg13g2_a21oi_1 _16527_ (.A1(_08092_),
    .A2(_08093_),
    .Y(_08102_),
    .B1(_08091_));
 sg13g2_a21oi_1 _16528_ (.A1(_08087_),
    .A2(_08089_),
    .Y(_08103_),
    .B1(_08086_));
 sg13g2_nand2b_1 _16529_ (.Y(_08104_),
    .B(\TRNG.hash[127] ),
    .A_N(\TRNG.hash[95] ));
 sg13g2_o21ai_1 _16530_ (.B1(_08104_),
    .Y(_08105_),
    .A1(\TRNG.hash[127] ),
    .A2(\TRNG.hash[63] ));
 sg13g2_a21oi_1 _16531_ (.A1(\TRNG.hash[30] ),
    .A2(_08084_),
    .Y(_08106_),
    .B1(_08083_));
 sg13g2_xor2_1 _16532_ (.B(\TRNG.sha256.W[31] ),
    .A(\TRNG.hash[120] ),
    .X(_08107_));
 sg13g2_xnor2_1 _16533_ (.Y(_08108_),
    .A(\TRNG.hash[31] ),
    .B(\TRNG.sha256.K[31] ));
 sg13g2_xor2_1 _16534_ (.B(\TRNG.hash[106] ),
    .A(net5550),
    .X(_08109_));
 sg13g2_xnor2_1 _16535_ (.Y(_08110_),
    .A(_08107_),
    .B(_08108_));
 sg13g2_xnor2_1 _16536_ (.Y(_08111_),
    .A(_08105_),
    .B(_08110_));
 sg13g2_xnor2_1 _16537_ (.Y(_08112_),
    .A(_08106_),
    .B(_08109_));
 sg13g2_xnor2_1 _16538_ (.Y(_08113_),
    .A(_08111_),
    .B(_08112_));
 sg13g2_xnor2_1 _16539_ (.Y(_08114_),
    .A(_08103_),
    .B(_08113_));
 sg13g2_xnor2_1 _16540_ (.Y(_08115_),
    .A(_08102_),
    .B(_08114_));
 sg13g2_xnor2_1 _16541_ (.Y(_08116_),
    .A(_08101_),
    .B(_08115_));
 sg13g2_xor2_1 _16542_ (.B(_08116_),
    .A(\TRNG.hash[159] ),
    .X(_08117_));
 sg13g2_or2_1 _16543_ (.X(_08118_),
    .B(_08117_),
    .A(_08100_));
 sg13g2_a21oi_1 _16544_ (.A1(_08100_),
    .A2(_08117_),
    .Y(_08119_),
    .B1(net5492));
 sg13g2_o21ai_1 _16545_ (.B1(\TRNG.hash[125] ),
    .Y(_08120_),
    .A1(\TRNG.hash[124] ),
    .A2(_08018_));
 sg13g2_and2_1 _16546_ (.A(_04221_),
    .B(_08120_),
    .X(_08121_));
 sg13g2_xnor2_1 _16547_ (.Y(_08122_),
    .A(net3619),
    .B(_08121_));
 sg13g2_o21ai_1 _16548_ (.B1(net4975),
    .Y(_08123_),
    .A1(\TRNG.hash[127] ),
    .A2(net5178));
 sg13g2_a221oi_1 _16549_ (.B2(net5189),
    .C1(_08123_),
    .B1(_08122_),
    .A1(_08118_),
    .Y(_00551_),
    .A2(_08119_));
 sg13g2_and3_1 _16550_ (.X(_08124_),
    .A(\TRNG.hash[161] ),
    .B(net5571),
    .C(\TRNG.hash[162] ));
 sg13g2_a21oi_1 _16551_ (.A1(\TRNG.hash[161] ),
    .A2(net5175),
    .Y(_08125_),
    .B1(net3563));
 sg13g2_nor3_1 _16552_ (.A(net4746),
    .B(_08124_),
    .C(_08125_),
    .Y(_08126_));
 sg13g2_a21o_1 _16553_ (.A2(net4744),
    .A1(net3567),
    .B1(_08126_),
    .X(_00552_));
 sg13g2_nand2_1 _16554_ (.Y(_08127_),
    .A(net5828),
    .B(net3731));
 sg13g2_o21ai_1 _16555_ (.B1(net5484),
    .Y(_08128_),
    .A1(\TRNG.hash[163] ),
    .A2(_08124_));
 sg13g2_nand3_1 _16556_ (.B(\TRNG.hash[163] ),
    .C(\TRNG.hash[162] ),
    .A(\TRNG.hash[161] ),
    .Y(_08129_));
 sg13g2_o21ai_1 _16557_ (.B1(net4974),
    .Y(_08130_),
    .A1(net5181),
    .A2(_08129_));
 sg13g2_a21oi_1 _16558_ (.A1(_08127_),
    .A2(_08128_),
    .Y(_00553_),
    .B1(_08130_));
 sg13g2_nand2_1 _16559_ (.Y(_08131_),
    .A(net3513),
    .B(net4743));
 sg13g2_o21ai_1 _16560_ (.B1(_00221_),
    .Y(_08132_),
    .A1(\TRNG.hash[164] ),
    .A2(_08129_));
 sg13g2_nor2_1 _16561_ (.A(\TRNG.hash[165] ),
    .B(_08132_),
    .Y(_08133_));
 sg13g2_nor3_1 _16562_ (.A(\TRNG.hash[166] ),
    .B(\TRNG.hash[165] ),
    .C(_08132_),
    .Y(_08134_));
 sg13g2_inv_1 _16563_ (.Y(_08135_),
    .A(_08134_));
 sg13g2_nor2_1 _16564_ (.A(_04228_),
    .B(_08134_),
    .Y(_08136_));
 sg13g2_xnor2_1 _16565_ (.Y(_08137_),
    .A(\TRNG.hash[167] ),
    .B(_08136_));
 sg13g2_o21ai_1 _16566_ (.B1(_08131_),
    .Y(_00554_),
    .A1(net4746),
    .A2(_08137_));
 sg13g2_a21oi_2 _16567_ (.B1(\TRNG.hash[168] ),
    .Y(_08138_),
    .A2(_08135_),
    .A1(\TRNG.hash[167] ));
 sg13g2_nor2b_1 _16568_ (.A(\TRNG.hash[169] ),
    .B_N(_08138_),
    .Y(_08139_));
 sg13g2_nor2b_1 _16569_ (.A(_08139_),
    .B_N(\TRNG.hash[170] ),
    .Y(_08140_));
 sg13g2_nand2b_1 _16570_ (.Y(_08141_),
    .B(_08139_),
    .A_N(\TRNG.hash[170] ));
 sg13g2_nand3b_1 _16571_ (.B(_08141_),
    .C(net5182),
    .Y(_08142_),
    .A_N(_08140_));
 sg13g2_a22oi_1 _16572_ (.Y(_08143_),
    .B1(net3773),
    .B2(net5345),
    .A2(net5816),
    .A1(net3760));
 sg13g2_a21oi_1 _16573_ (.A1(_08142_),
    .A2(_08143_),
    .Y(_00555_),
    .B1(net4960));
 sg13g2_and2_1 _16574_ (.A(\TRNG.hash[171] ),
    .B(_08140_),
    .X(_08144_));
 sg13g2_o21ai_1 _16575_ (.B1(net5182),
    .Y(_08145_),
    .A1(\TRNG.hash[171] ),
    .A2(_08140_));
 sg13g2_a22oi_1 _16576_ (.Y(_08146_),
    .B1(net3888),
    .B2(net5345),
    .A2(net5818),
    .A1(net3845));
 sg13g2_o21ai_1 _16577_ (.B1(_08146_),
    .Y(_08147_),
    .A1(_08144_),
    .A2(_08145_));
 sg13g2_and2_1 _16578_ (.A(net4974),
    .B(_08147_),
    .X(_00556_));
 sg13g2_nor3_2 _16579_ (.A(\TRNG.hash[173] ),
    .B(\TRNG.hash[172] ),
    .C(_08144_),
    .Y(_08148_));
 sg13g2_nor2b_1 _16580_ (.A(\TRNG.hash[174] ),
    .B_N(_08148_),
    .Y(_08149_));
 sg13g2_nor2b_1 _16581_ (.A(\TRNG.hash[175] ),
    .B_N(_08149_),
    .Y(_08150_));
 sg13g2_nor2_2 _16582_ (.A(_04290_),
    .B(_08150_),
    .Y(_08151_));
 sg13g2_a21oi_1 _16583_ (.A1(_04290_),
    .A2(_08150_),
    .Y(_08152_),
    .B1(net5181));
 sg13g2_nand2b_1 _16584_ (.Y(_08153_),
    .B(_08152_),
    .A_N(_08151_));
 sg13g2_a22oi_1 _16585_ (.Y(_08154_),
    .B1(net3647),
    .B2(net5345),
    .A2(net5822),
    .A1(net3636));
 sg13g2_a21oi_1 _16586_ (.A1(_08153_),
    .A2(_08154_),
    .Y(_00557_),
    .B1(net4960));
 sg13g2_nor3_1 _16587_ (.A(\TRNG.hash[178] ),
    .B(\TRNG.hash[177] ),
    .C(_08151_),
    .Y(_08155_));
 sg13g2_nor2b_1 _16588_ (.A(\TRNG.hash[179] ),
    .B_N(_08155_),
    .Y(_08156_));
 sg13g2_nand2b_2 _16589_ (.Y(_08157_),
    .B(net3579),
    .A_N(_08156_));
 sg13g2_a21oi_1 _16590_ (.A1(_04289_),
    .A2(_08156_),
    .Y(_08158_),
    .B1(net5181));
 sg13g2_nand2_1 _16591_ (.Y(_08159_),
    .A(_08157_),
    .B(_08158_));
 sg13g2_a22oi_1 _16592_ (.Y(_08160_),
    .B1(net3579),
    .B2(net5346),
    .A2(\TRNG.hash[212] ),
    .A1(net5833));
 sg13g2_a21oi_1 _16593_ (.A1(_08159_),
    .A2(net3580),
    .Y(_00558_),
    .B1(net4961));
 sg13g2_nand2b_1 _16594_ (.Y(_08161_),
    .B(_08157_),
    .A_N(\TRNG.hash[181] ));
 sg13g2_nor2_1 _16595_ (.A(\TRNG.hash[182] ),
    .B(_08161_),
    .Y(_08162_));
 sg13g2_nor2b_1 _16596_ (.A(_08162_),
    .B_N(\TRNG.hash[183] ),
    .Y(_08163_));
 sg13g2_nor3_1 _16597_ (.A(\TRNG.hash[182] ),
    .B(\TRNG.hash[183] ),
    .C(_08161_),
    .Y(_08164_));
 sg13g2_or3_1 _16598_ (.A(net5181),
    .B(_08163_),
    .C(_08164_),
    .X(_08165_));
 sg13g2_a22oi_1 _16599_ (.Y(_08166_),
    .B1(net3805),
    .B2(net5348),
    .A2(\TRNG.hash[215] ),
    .A1(net5842));
 sg13g2_a21oi_1 _16600_ (.A1(_08165_),
    .A2(net3806),
    .Y(_00559_),
    .B1(net4963));
 sg13g2_and2_1 _16601_ (.A(\TRNG.hash[184] ),
    .B(_08163_),
    .X(_08167_));
 sg13g2_nor2_1 _16602_ (.A(net5181),
    .B(_08167_),
    .Y(_08168_));
 sg13g2_o21ai_1 _16603_ (.B1(_08168_),
    .Y(_08169_),
    .A1(net3823),
    .A2(_08163_));
 sg13g2_a22oi_1 _16604_ (.Y(_08170_),
    .B1(net3823),
    .B2(net5347),
    .A2(net5842),
    .A1(net3786));
 sg13g2_a21oi_1 _16605_ (.A1(_08169_),
    .A2(_08170_),
    .Y(_00560_),
    .B1(net4963));
 sg13g2_nand2_2 _16606_ (.Y(_08171_),
    .A(\TRNG.hash[185] ),
    .B(_08167_));
 sg13g2_o21ai_1 _16607_ (.B1(net5184),
    .Y(_08172_),
    .A1(\TRNG.hash[185] ),
    .A2(_08167_));
 sg13g2_nand2b_1 _16608_ (.Y(_08173_),
    .B(_08171_),
    .A_N(_08172_));
 sg13g2_a22oi_1 _16609_ (.Y(_08174_),
    .B1(net3861),
    .B2(net5347),
    .A2(net5839),
    .A1(net3814));
 sg13g2_a21oi_1 _16610_ (.A1(_08173_),
    .A2(_08174_),
    .Y(_00561_),
    .B1(net4962));
 sg13g2_nor3_1 _16611_ (.A(\TRNG.hash[188] ),
    .B(\TRNG.hash[187] ),
    .C(\TRNG.hash[186] ),
    .Y(_08175_));
 sg13g2_nand2_1 _16612_ (.Y(_08176_),
    .A(_08171_),
    .B(_08175_));
 sg13g2_or2_1 _16613_ (.X(_08177_),
    .B(_08176_),
    .A(\TRNG.hash[189] ));
 sg13g2_nand2_1 _16614_ (.Y(_08178_),
    .A(\TRNG.hash[190] ),
    .B(_08177_));
 sg13g2_o21ai_1 _16615_ (.B1(net5184),
    .Y(_08179_),
    .A1(\TRNG.hash[190] ),
    .A2(_08177_));
 sg13g2_nand2b_1 _16616_ (.Y(_08180_),
    .B(_08178_),
    .A_N(_08179_));
 sg13g2_a22oi_1 _16617_ (.Y(_08181_),
    .B1(\TRNG.hash[190] ),
    .B2(net5347),
    .A2(net3778),
    .A1(net5839));
 sg13g2_a21oi_1 _16618_ (.A1(_08180_),
    .A2(net3779),
    .Y(_00562_),
    .B1(net4962));
 sg13g2_xnor2_1 _16619_ (.Y(_08182_),
    .A(\TRNG.hash[191] ),
    .B(_08178_));
 sg13g2_nand2_1 _16620_ (.Y(_08183_),
    .A(net5184),
    .B(_08182_));
 sg13g2_a22oi_1 _16621_ (.Y(_08184_),
    .B1(net3801),
    .B2(net5347),
    .A2(net5844),
    .A1(\TRNG.hash[223] ));
 sg13g2_a21oi_1 _16622_ (.A1(_08183_),
    .A2(net3802),
    .Y(_00563_),
    .B1(net4962));
 sg13g2_nand2_1 _16623_ (.Y(_08185_),
    .A(net5569),
    .B(net4744));
 sg13g2_nand2_1 _16624_ (.Y(_08186_),
    .A(\TRNG.hash[192] ),
    .B(net5571));
 sg13g2_xor2_1 _16625_ (.B(_08186_),
    .A(net3897),
    .X(_08187_));
 sg13g2_o21ai_1 _16626_ (.B1(_08185_),
    .Y(_00564_),
    .A1(net4746),
    .A2(_08187_));
 sg13g2_a21o_1 _16627_ (.A2(\TRNG.hash[193] ),
    .A1(\TRNG.hash[192] ),
    .B1(\TRNG.hash[194] ),
    .X(_08188_));
 sg13g2_nand2_1 _16628_ (.Y(_08189_),
    .A(net5571),
    .B(_08188_));
 sg13g2_xor2_1 _16629_ (.B(_08189_),
    .A(net3731),
    .X(_08190_));
 sg13g2_nand2_1 _16630_ (.Y(_08191_),
    .A(net5888),
    .B(net4743));
 sg13g2_o21ai_1 _16631_ (.B1(_08191_),
    .Y(_00565_),
    .A1(net4746),
    .A2(_08190_));
 sg13g2_nand2_1 _16632_ (.Y(_08192_),
    .A(net5887),
    .B(net4743));
 sg13g2_and3_1 _16633_ (.X(_08193_),
    .A(\TRNG.hash[195] ),
    .B(net5175),
    .C(_08188_));
 sg13g2_nand3_1 _16634_ (.B(\TRNG.hash[195] ),
    .C(_08188_),
    .A(\TRNG.hash[196] ),
    .Y(_08194_));
 sg13g2_nor2_1 _16635_ (.A(_04228_),
    .B(_08194_),
    .Y(_08195_));
 sg13g2_o21ai_1 _16636_ (.B1(_06876_),
    .Y(_08196_),
    .A1(net3872),
    .A2(_08193_));
 sg13g2_o21ai_1 _16637_ (.B1(_08192_),
    .Y(_00566_),
    .A1(_08195_),
    .A2(_08196_));
 sg13g2_nand2_1 _16638_ (.Y(_08197_),
    .A(net5567),
    .B(net4743));
 sg13g2_and2_1 _16639_ (.A(\TRNG.hash[197] ),
    .B(_08195_),
    .X(_08198_));
 sg13g2_xnor2_1 _16640_ (.Y(_08199_),
    .A(net3863),
    .B(_08195_));
 sg13g2_o21ai_1 _16641_ (.B1(_08197_),
    .Y(_00567_),
    .A1(net4746),
    .A2(_08199_));
 sg13g2_nand2_1 _16642_ (.Y(_08200_),
    .A(\TRNG.hash[198] ),
    .B(\TRNG.hash[197] ));
 sg13g2_o21ai_1 _16643_ (.B1(_06876_),
    .Y(_08201_),
    .A1(\TRNG.hash[198] ),
    .A2(_08198_));
 sg13g2_a21oi_1 _16644_ (.A1(net3878),
    .A2(_08198_),
    .Y(_08202_),
    .B1(_08201_));
 sg13g2_a21o_1 _16645_ (.A2(net4743),
    .A1(net5566),
    .B1(_08202_),
    .X(_00568_));
 sg13g2_nand2_1 _16646_ (.Y(_08203_),
    .A(net5886),
    .B(net4743));
 sg13g2_o21ai_1 _16647_ (.B1(_04225_),
    .Y(_08204_),
    .A1(_08194_),
    .A2(_08200_));
 sg13g2_nand2_1 _16648_ (.Y(_08205_),
    .A(net5571),
    .B(_08204_));
 sg13g2_xor2_1 _16649_ (.B(_08205_),
    .A(\TRNG.hash[200] ),
    .X(_08206_));
 sg13g2_o21ai_1 _16650_ (.B1(_08203_),
    .Y(_00569_),
    .A1(net4746),
    .A2(_08206_));
 sg13g2_nand2_2 _16651_ (.Y(_08207_),
    .A(\TRNG.hash[200] ),
    .B(_08204_));
 sg13g2_nor3_1 _16652_ (.A(\TRNG.hash[203] ),
    .B(\TRNG.hash[202] ),
    .C(\TRNG.hash[201] ),
    .Y(_08208_));
 sg13g2_nand2_1 _16653_ (.Y(_08209_),
    .A(_08207_),
    .B(_08208_));
 sg13g2_nand2_1 _16654_ (.Y(_08210_),
    .A(\TRNG.hash[204] ),
    .B(_08209_));
 sg13g2_inv_1 _16655_ (.Y(_08211_),
    .A(_08210_));
 sg13g2_o21ai_1 _16656_ (.B1(net5182),
    .Y(_08212_),
    .A1(\TRNG.hash[204] ),
    .A2(_08209_));
 sg13g2_nand2b_1 _16657_ (.Y(_08213_),
    .B(_08210_),
    .A_N(_08212_));
 sg13g2_a22oi_1 _16658_ (.Y(_08214_),
    .B1(net3838),
    .B2(net5345),
    .A2(net5885),
    .A1(net5817));
 sg13g2_a21oi_1 _16659_ (.A1(_08213_),
    .A2(net3839),
    .Y(_00570_),
    .B1(net4960));
 sg13g2_o21ai_1 _16660_ (.B1(net3437),
    .Y(_08215_),
    .A1(\TRNG.hash[205] ),
    .A2(_08210_));
 sg13g2_nand2_1 _16661_ (.Y(_08216_),
    .A(\TRNG.hash[206] ),
    .B(_08215_));
 sg13g2_o21ai_1 _16662_ (.B1(net5182),
    .Y(_08217_),
    .A1(\TRNG.hash[206] ),
    .A2(_08215_));
 sg13g2_nand2b_1 _16663_ (.Y(_08218_),
    .B(_08216_),
    .A_N(_08217_));
 sg13g2_a22oi_1 _16664_ (.Y(_08219_),
    .B1(net3808),
    .B2(net5345),
    .A2(net5817),
    .A1(net5562));
 sg13g2_a21oi_1 _16665_ (.A1(_08218_),
    .A2(_08219_),
    .Y(_00571_),
    .B1(net4960));
 sg13g2_o21ai_1 _16666_ (.B1(\TRNG.hash[206] ),
    .Y(_08220_),
    .A1(\TRNG.hash[205] ),
    .A2(_08211_));
 sg13g2_nand2b_1 _16667_ (.Y(_08221_),
    .B(_08220_),
    .A_N(\TRNG.hash[207] ));
 sg13g2_nor3_2 _16668_ (.A(\TRNG.hash[209] ),
    .B(\TRNG.hash[208] ),
    .C(_08221_),
    .Y(_08222_));
 sg13g2_nand2b_1 _16669_ (.Y(_08223_),
    .B(_08222_),
    .A_N(\TRNG.hash[210] ));
 sg13g2_and2_2 _16670_ (.A(\TRNG.hash[211] ),
    .B(_08223_),
    .X(_08224_));
 sg13g2_nor2_1 _16671_ (.A(net5181),
    .B(_08224_),
    .Y(_08225_));
 sg13g2_o21ai_1 _16672_ (.B1(_08225_),
    .Y(_08226_),
    .A1(net3799),
    .A2(_08223_));
 sg13g2_a22oi_1 _16673_ (.Y(_08227_),
    .B1(net3799),
    .B2(net5345),
    .A2(net5825),
    .A1(net5560));
 sg13g2_a21oi_1 _16674_ (.A1(_08226_),
    .A2(net3800),
    .Y(_00572_),
    .B1(net4960));
 sg13g2_nand2_2 _16675_ (.Y(_08228_),
    .A(\TRNG.hash[212] ),
    .B(_08224_));
 sg13g2_o21ai_1 _16676_ (.B1(net5183),
    .Y(_08229_),
    .A1(\TRNG.hash[212] ),
    .A2(_08224_));
 sg13g2_nand2b_1 _16677_ (.Y(_08230_),
    .B(_08228_),
    .A_N(_08229_));
 sg13g2_a22oi_1 _16678_ (.Y(_08231_),
    .B1(\TRNG.hash[212] ),
    .B2(net5346),
    .A2(net3432),
    .A1(net5833));
 sg13g2_a21oi_1 _16679_ (.A1(_08230_),
    .A2(net3433),
    .Y(_00573_),
    .B1(net4961));
 sg13g2_o21ai_1 _16680_ (.B1(net3530),
    .Y(_08232_),
    .A1(\TRNG.hash[213] ),
    .A2(_08228_));
 sg13g2_nor2_1 _16681_ (.A(\TRNG.hash[214] ),
    .B(_08232_),
    .Y(_08233_));
 sg13g2_xnor2_1 _16682_ (.Y(_08234_),
    .A(\TRNG.hash[215] ),
    .B(_08233_));
 sg13g2_nand2_1 _16683_ (.Y(_08235_),
    .A(net5185),
    .B(_08234_));
 sg13g2_a22oi_1 _16684_ (.Y(_08236_),
    .B1(\TRNG.hash[215] ),
    .B2(net5348),
    .A2(net3395),
    .A1(net5842));
 sg13g2_a21oi_1 _16685_ (.A1(_08235_),
    .A2(net3396),
    .Y(_00574_),
    .B1(net4963));
 sg13g2_nand3_1 _16686_ (.B(_04224_),
    .C(_08228_),
    .A(_04223_),
    .Y(_08237_));
 sg13g2_a21oi_2 _16687_ (.B1(\TRNG.hash[216] ),
    .Y(_08238_),
    .A2(_08237_),
    .A1(\TRNG.hash[215] ));
 sg13g2_nor2b_1 _16688_ (.A(\TRNG.hash[217] ),
    .B_N(_08238_),
    .Y(_08239_));
 sg13g2_nand2b_1 _16689_ (.Y(_08240_),
    .B(\TRNG.hash[218] ),
    .A_N(_08239_));
 sg13g2_a21oi_1 _16690_ (.A1(_04286_),
    .A2(_08239_),
    .Y(_08241_),
    .B1(net5181));
 sg13g2_nand2_1 _16691_ (.Y(_08242_),
    .A(_08240_),
    .B(_08241_));
 sg13g2_a22oi_1 _16692_ (.Y(_08243_),
    .B1(\TRNG.hash[218] ),
    .B2(net5347),
    .A2(net3569),
    .A1(net5837));
 sg13g2_a21oi_1 _16693_ (.A1(_08242_),
    .A2(net3570),
    .Y(_00575_),
    .B1(net4962));
 sg13g2_o21ai_1 _16694_ (.B1(_00227_),
    .Y(_08244_),
    .A1(\TRNG.hash[219] ),
    .A2(_08240_));
 sg13g2_nor2_1 _16695_ (.A(\TRNG.hash[220] ),
    .B(_08244_),
    .Y(_08245_));
 sg13g2_nor3_1 _16696_ (.A(\TRNG.hash[221] ),
    .B(\TRNG.hash[220] ),
    .C(_08244_),
    .Y(_08246_));
 sg13g2_nand2b_1 _16697_ (.Y(_08247_),
    .B(\TRNG.hash[222] ),
    .A_N(_08246_));
 sg13g2_a21oi_1 _16698_ (.A1(_04285_),
    .A2(_08246_),
    .Y(_08248_),
    .B1(net5181));
 sg13g2_nand2_1 _16699_ (.Y(_08249_),
    .A(_08247_),
    .B(_08248_));
 sg13g2_a22oi_1 _16700_ (.Y(_08250_),
    .B1(\TRNG.hash[222] ),
    .B2(net5347),
    .A2(net5840),
    .A1(net3427));
 sg13g2_a21oi_1 _16701_ (.A1(_08249_),
    .A2(net3428),
    .Y(_00576_),
    .B1(net4962));
 sg13g2_xnor2_1 _16702_ (.Y(_08251_),
    .A(net5879),
    .B(\TRNG.hash[228] ));
 sg13g2_xnor2_1 _16703_ (.Y(_08252_),
    .A(\TRNG.hash[239] ),
    .B(_08251_));
 sg13g2_xnor2_1 _16704_ (.Y(_08253_),
    .A(_07324_),
    .B(_08252_));
 sg13g2_nor2_1 _16705_ (.A(net5568),
    .B(\TRNG.hash[162] ),
    .Y(_08254_));
 sg13g2_a21oi_1 _16706_ (.A1(net5568),
    .A2(\TRNG.hash[162] ),
    .Y(_08255_),
    .B1(\TRNG.hash[194] ));
 sg13g2_nor2_1 _16707_ (.A(_08254_),
    .B(_08255_),
    .Y(_08256_));
 sg13g2_nor2b_1 _16708_ (.A(_08253_),
    .B_N(_08256_),
    .Y(_08257_));
 sg13g2_xnor2_1 _16709_ (.Y(_08258_),
    .A(_08253_),
    .B(_08256_));
 sg13g2_xnor2_1 _16710_ (.Y(_08259_),
    .A(net5880),
    .B(\TRNG.hash[227] ));
 sg13g2_xnor2_1 _16711_ (.Y(_08260_),
    .A(\TRNG.hash[238] ),
    .B(_08259_));
 sg13g2_nor2b_1 _16712_ (.A(_07328_),
    .B_N(_08260_),
    .Y(_08261_));
 sg13g2_xnor2_1 _16713_ (.Y(_08262_),
    .A(_07328_),
    .B(_08260_));
 sg13g2_nor2_1 _16714_ (.A(net5569),
    .B(\TRNG.hash[193] ),
    .Y(_08263_));
 sg13g2_a21oi_1 _16715_ (.A1(net5569),
    .A2(\TRNG.hash[193] ),
    .Y(_08264_),
    .B1(\TRNG.hash[161] ));
 sg13g2_nor2_1 _16716_ (.A(_08263_),
    .B(_08264_),
    .Y(_08265_));
 sg13g2_a21oi_1 _16717_ (.A1(_08262_),
    .A2(_08265_),
    .Y(_08266_),
    .B1(_08261_));
 sg13g2_nor2b_1 _16718_ (.A(_08266_),
    .B_N(_08258_),
    .Y(_08267_));
 sg13g2_xnor2_1 _16719_ (.Y(_08268_),
    .A(\TRNG.hash[226] ),
    .B(\TRNG.hash[246] ));
 sg13g2_xnor2_1 _16720_ (.Y(_08269_),
    .A(\TRNG.hash[237] ),
    .B(_08268_));
 sg13g2_xnor2_1 _16721_ (.Y(_08270_),
    .A(_07330_),
    .B(_08269_));
 sg13g2_nor2_1 _16722_ (.A(net5570),
    .B(\TRNG.hash[160] ),
    .Y(_08271_));
 sg13g2_a21oi_1 _16723_ (.A1(net5570),
    .A2(\TRNG.hash[160] ),
    .Y(_08272_),
    .B1(\TRNG.hash[192] ));
 sg13g2_nor2_1 _16724_ (.A(_08271_),
    .B(_08272_),
    .Y(_08273_));
 sg13g2_nor2b_1 _16725_ (.A(_08270_),
    .B_N(_08273_),
    .Y(_08274_));
 sg13g2_a21oi_1 _16726_ (.A1(_07330_),
    .A2(_08269_),
    .Y(_08275_),
    .B1(_08274_));
 sg13g2_xnor2_1 _16727_ (.Y(_08276_),
    .A(_08262_),
    .B(_08265_));
 sg13g2_or2_1 _16728_ (.X(_08277_),
    .B(_08276_),
    .A(_08275_));
 sg13g2_inv_1 _16729_ (.Y(_08278_),
    .A(_08277_));
 sg13g2_xnor2_1 _16730_ (.Y(_08279_),
    .A(_08258_),
    .B(_08266_));
 sg13g2_a21oi_1 _16731_ (.A1(_08278_),
    .A2(_08279_),
    .Y(_08280_),
    .B1(_08267_));
 sg13g2_a21oi_1 _16732_ (.A1(_07324_),
    .A2(_08252_),
    .Y(_08281_),
    .B1(_08257_));
 sg13g2_xnor2_1 _16733_ (.Y(_08282_),
    .A(\TRNG.hash[240] ),
    .B(\TRNG.hash[229] ));
 sg13g2_xnor2_1 _16734_ (.Y(_08283_),
    .A(net5559),
    .B(_08282_));
 sg13g2_xnor2_1 _16735_ (.Y(_08284_),
    .A(_07337_),
    .B(_08283_));
 sg13g2_nor2_1 _16736_ (.A(\TRNG.hash[195] ),
    .B(\TRNG.hash[163] ),
    .Y(_08285_));
 sg13g2_a21oi_1 _16737_ (.A1(\TRNG.hash[195] ),
    .A2(\TRNG.hash[163] ),
    .Y(_08286_),
    .B1(net5888));
 sg13g2_nor2_1 _16738_ (.A(_08285_),
    .B(_08286_),
    .Y(_08287_));
 sg13g2_nor2b_1 _16739_ (.A(_08284_),
    .B_N(_08287_),
    .Y(_08288_));
 sg13g2_xnor2_1 _16740_ (.Y(_08289_),
    .A(_08284_),
    .B(_08287_));
 sg13g2_nand2b_1 _16741_ (.Y(_08290_),
    .B(_08289_),
    .A_N(_08281_));
 sg13g2_nor2b_1 _16742_ (.A(_08289_),
    .B_N(_08281_),
    .Y(_08291_));
 sg13g2_xor2_1 _16743_ (.B(_08289_),
    .A(_08281_),
    .X(_08292_));
 sg13g2_xnor2_1 _16744_ (.Y(_08293_),
    .A(_08280_),
    .B(_08292_));
 sg13g2_or2_1 _16745_ (.X(_08294_),
    .B(net5570),
    .A(net5569));
 sg13g2_nor2_1 _16746_ (.A(net5568),
    .B(_08294_),
    .Y(_08295_));
 sg13g2_nor2b_2 _16747_ (.A(_08295_),
    .B_N(net5888),
    .Y(_08296_));
 sg13g2_xor2_1 _16748_ (.B(_08295_),
    .A(net5888),
    .X(_08297_));
 sg13g2_o21ai_1 _16749_ (.B1(net4974),
    .Y(_08298_),
    .A1(net5888),
    .A2(net5175));
 sg13g2_a221oi_1 _16750_ (.B2(net5183),
    .C1(_08298_),
    .B1(_08297_),
    .A1(net5827),
    .Y(_00577_),
    .A2(_08293_));
 sg13g2_o21ai_1 _16751_ (.B1(_08290_),
    .Y(_08299_),
    .A1(_08280_),
    .A2(_08291_));
 sg13g2_a21oi_1 _16752_ (.A1(_07337_),
    .A2(_08283_),
    .Y(_08300_),
    .B1(_08288_));
 sg13g2_xnor2_1 _16753_ (.Y(_08301_),
    .A(net5878),
    .B(net5884));
 sg13g2_xnor2_1 _16754_ (.Y(_08302_),
    .A(net5566),
    .B(_08301_));
 sg13g2_nor2b_1 _16755_ (.A(_07320_),
    .B_N(_08302_),
    .Y(_08303_));
 sg13g2_xnor2_1 _16756_ (.Y(_08304_),
    .A(_07320_),
    .B(_08302_));
 sg13g2_nor2_1 _16757_ (.A(net5887),
    .B(\TRNG.hash[196] ),
    .Y(_08305_));
 sg13g2_a21oi_1 _16758_ (.A1(net5887),
    .A2(\TRNG.hash[196] ),
    .Y(_08306_),
    .B1(\TRNG.hash[164] ));
 sg13g2_nor2_1 _16759_ (.A(_08305_),
    .B(_08306_),
    .Y(_08307_));
 sg13g2_xnor2_1 _16760_ (.Y(_08308_),
    .A(_08304_),
    .B(_08307_));
 sg13g2_nor2_1 _16761_ (.A(_08300_),
    .B(_08308_),
    .Y(_08309_));
 sg13g2_xor2_1 _16762_ (.B(_08308_),
    .A(_08300_),
    .X(_08310_));
 sg13g2_xnor2_1 _16763_ (.Y(_08311_),
    .A(_08299_),
    .B(_08310_));
 sg13g2_nand2_2 _16764_ (.Y(_08312_),
    .A(net5887),
    .B(_08296_));
 sg13g2_xnor2_1 _16765_ (.Y(_08313_),
    .A(net5887),
    .B(_08296_));
 sg13g2_o21ai_1 _16766_ (.B1(net4974),
    .Y(_08314_),
    .A1(net5887),
    .A2(net5175));
 sg13g2_a221oi_1 _16767_ (.B2(net5182),
    .C1(_08314_),
    .B1(_08313_),
    .A1(net5820),
    .Y(_00578_),
    .A2(_08311_));
 sg13g2_xnor2_1 _16768_ (.Y(_08315_),
    .A(net5877),
    .B(\TRNG.hash[232] ));
 sg13g2_xnor2_1 _16769_ (.Y(_08316_),
    .A(net5560),
    .B(_08315_));
 sg13g2_and2_1 _16770_ (.A(_07370_),
    .B(_08316_),
    .X(_08317_));
 sg13g2_or2_1 _16771_ (.X(_08318_),
    .B(_08316_),
    .A(_07370_));
 sg13g2_nand2b_1 _16772_ (.Y(_08319_),
    .B(_08318_),
    .A_N(_08317_));
 sg13g2_nor2_1 _16773_ (.A(\TRNG.hash[230] ),
    .B(\TRNG.hash[198] ),
    .Y(_08320_));
 sg13g2_a21oi_1 _16774_ (.A1(\TRNG.hash[230] ),
    .A2(\TRNG.hash[198] ),
    .Y(_08321_),
    .B1(\TRNG.hash[166] ));
 sg13g2_nor2_1 _16775_ (.A(_08320_),
    .B(_08321_),
    .Y(_08322_));
 sg13g2_xnor2_1 _16776_ (.Y(_08323_),
    .A(_08319_),
    .B(_08322_));
 sg13g2_xnor2_1 _16777_ (.Y(_08324_),
    .A(net5883),
    .B(\TRNG.hash[231] ));
 sg13g2_xnor2_1 _16778_ (.Y(_08325_),
    .A(\TRNG.hash[251] ),
    .B(_08324_));
 sg13g2_nor2b_1 _16779_ (.A(_07315_),
    .B_N(_08325_),
    .Y(_08326_));
 sg13g2_xnor2_1 _16780_ (.Y(_08327_),
    .A(_07315_),
    .B(_08325_));
 sg13g2_nor2_1 _16781_ (.A(net5567),
    .B(\TRNG.hash[197] ),
    .Y(_08328_));
 sg13g2_a21oi_1 _16782_ (.A1(net5567),
    .A2(\TRNG.hash[197] ),
    .Y(_08329_),
    .B1(\TRNG.hash[165] ));
 sg13g2_nor2_1 _16783_ (.A(_08328_),
    .B(_08329_),
    .Y(_08330_));
 sg13g2_a21oi_1 _16784_ (.A1(_08327_),
    .A2(_08330_),
    .Y(_08331_),
    .B1(_08326_));
 sg13g2_nand2b_1 _16785_ (.Y(_08332_),
    .B(_08323_),
    .A_N(_08331_));
 sg13g2_xnor2_1 _16786_ (.Y(_08333_),
    .A(_08327_),
    .B(_08330_));
 sg13g2_a21o_1 _16787_ (.A2(_08307_),
    .A1(_08304_),
    .B1(_08303_),
    .X(_08334_));
 sg13g2_nor2b_1 _16788_ (.A(_08333_),
    .B_N(_08334_),
    .Y(_08335_));
 sg13g2_a21o_1 _16789_ (.A2(_08310_),
    .A1(_08299_),
    .B1(_08309_),
    .X(_08336_));
 sg13g2_nand2b_1 _16790_ (.Y(_08337_),
    .B(_08333_),
    .A_N(_08334_));
 sg13g2_nand2b_1 _16791_ (.Y(_08338_),
    .B(_08337_),
    .A_N(_08335_));
 sg13g2_a21oi_1 _16792_ (.A1(_08336_),
    .A2(_08337_),
    .Y(_08339_),
    .B1(_08335_));
 sg13g2_xor2_1 _16793_ (.B(_08331_),
    .A(_08323_),
    .X(_08340_));
 sg13g2_o21ai_1 _16794_ (.B1(_08332_),
    .Y(_08341_),
    .A1(_08339_),
    .A2(_08340_));
 sg13g2_a21oi_1 _16795_ (.A1(_08318_),
    .A2(_08322_),
    .Y(_08342_),
    .B1(_08317_));
 sg13g2_xnor2_1 _16796_ (.Y(_08343_),
    .A(\TRNG.hash[233] ),
    .B(net5882));
 sg13g2_xnor2_1 _16797_ (.Y(_08344_),
    .A(net5557),
    .B(_08343_));
 sg13g2_nand2b_1 _16798_ (.Y(_08345_),
    .B(_08344_),
    .A_N(_07395_));
 sg13g2_xnor2_1 _16799_ (.Y(_08346_),
    .A(_07395_),
    .B(_08344_));
 sg13g2_a21oi_1 _16800_ (.A1(\TRNG.hash[231] ),
    .A2(\TRNG.hash[167] ),
    .Y(_08347_),
    .B1(\TRNG.hash[199] ));
 sg13g2_a21oi_1 _16801_ (.A1(_04284_),
    .A2(_04292_),
    .Y(_08348_),
    .B1(_08347_));
 sg13g2_nand2_1 _16802_ (.Y(_08349_),
    .A(_08346_),
    .B(_08348_));
 sg13g2_xnor2_1 _16803_ (.Y(_08350_),
    .A(_08346_),
    .B(_08348_));
 sg13g2_nor2_1 _16804_ (.A(_08342_),
    .B(_08350_),
    .Y(_08351_));
 sg13g2_nand2_1 _16805_ (.Y(_08352_),
    .A(_08342_),
    .B(_08350_));
 sg13g2_nand2b_1 _16806_ (.Y(_08353_),
    .B(_08352_),
    .A_N(_08351_));
 sg13g2_xnor2_1 _16807_ (.Y(_08354_),
    .A(_08341_),
    .B(_08353_));
 sg13g2_nand2_1 _16808_ (.Y(_08355_),
    .A(net4743),
    .B(_08354_));
 sg13g2_o21ai_1 _16809_ (.B1(net3767),
    .Y(_08356_),
    .A1(net5567),
    .A2(_08312_));
 sg13g2_o21ai_1 _16810_ (.B1(net5571),
    .Y(_08357_),
    .A1(net5566),
    .A2(_08356_));
 sg13g2_xnor2_1 _16811_ (.Y(_08358_),
    .A(_04284_),
    .B(_08357_));
 sg13g2_o21ai_1 _16812_ (.B1(_08355_),
    .Y(_00579_),
    .A1(net4746),
    .A2(_08358_));
 sg13g2_xnor2_1 _16813_ (.Y(_08359_),
    .A(\TRNG.hash[234] ),
    .B(net5881));
 sg13g2_xnor2_1 _16814_ (.Y(_08360_),
    .A(net5556),
    .B(_08359_));
 sg13g2_nor2b_1 _16815_ (.A(_07432_),
    .B_N(_08360_),
    .Y(_08361_));
 sg13g2_xnor2_1 _16816_ (.Y(_08362_),
    .A(_07432_),
    .B(_08360_));
 sg13g2_nor2_1 _16817_ (.A(net5886),
    .B(\TRNG.hash[200] ),
    .Y(_08363_));
 sg13g2_a21oi_1 _16818_ (.A1(net5886),
    .A2(\TRNG.hash[200] ),
    .Y(_08364_),
    .B1(\TRNG.hash[168] ));
 sg13g2_nor2_1 _16819_ (.A(_08363_),
    .B(_08364_),
    .Y(_08365_));
 sg13g2_xnor2_1 _16820_ (.Y(_08366_),
    .A(_08362_),
    .B(_08365_));
 sg13g2_a21oi_1 _16821_ (.A1(_08345_),
    .A2(_08349_),
    .Y(_08367_),
    .B1(_08366_));
 sg13g2_nand3_1 _16822_ (.B(_08349_),
    .C(_08366_),
    .A(_08345_),
    .Y(_08368_));
 sg13g2_nand2b_1 _16823_ (.Y(_08369_),
    .B(_08368_),
    .A_N(_08367_));
 sg13g2_a21oi_2 _16824_ (.B1(_08351_),
    .Y(_08370_),
    .A2(_08352_),
    .A1(_08341_));
 sg13g2_nor2_1 _16825_ (.A(_08369_),
    .B(_08370_),
    .Y(_08371_));
 sg13g2_xnor2_1 _16826_ (.Y(_08372_),
    .A(_08369_),
    .B(_08370_));
 sg13g2_nor2_1 _16827_ (.A(net5566),
    .B(net5567),
    .Y(_08373_));
 sg13g2_a21oi_2 _16828_ (.B1(_04284_),
    .Y(_08374_),
    .A2(_08373_),
    .A1(_08312_));
 sg13g2_nand2_2 _16829_ (.Y(_08375_),
    .A(net5886),
    .B(_08374_));
 sg13g2_xnor2_1 _16830_ (.Y(_08376_),
    .A(net5886),
    .B(_08374_));
 sg13g2_o21ai_1 _16831_ (.B1(net4974),
    .Y(_08377_),
    .A1(net5886),
    .A2(net5175));
 sg13g2_a221oi_1 _16832_ (.B2(net5182),
    .C1(_08377_),
    .B1(_08376_),
    .A1(net5820),
    .Y(_00580_),
    .A2(_08372_));
 sg13g2_xnor2_1 _16833_ (.Y(_08378_),
    .A(net5880),
    .B(net5885));
 sg13g2_xnor2_1 _16834_ (.Y(_08379_),
    .A(net5570),
    .B(_08378_));
 sg13g2_nor2b_1 _16835_ (.A(_07489_),
    .B_N(_08379_),
    .Y(_08380_));
 sg13g2_xnor2_1 _16836_ (.Y(_08381_),
    .A(_07489_),
    .B(_08379_));
 sg13g2_nor2_1 _16837_ (.A(net5564),
    .B(\TRNG.hash[170] ),
    .Y(_08382_));
 sg13g2_a21oi_1 _16838_ (.A1(net5564),
    .A2(\TRNG.hash[170] ),
    .Y(_08383_),
    .B1(\TRNG.hash[202] ));
 sg13g2_nor2_1 _16839_ (.A(_08382_),
    .B(_08383_),
    .Y(_08384_));
 sg13g2_xnor2_1 _16840_ (.Y(_08385_),
    .A(_08381_),
    .B(_08384_));
 sg13g2_xnor2_1 _16841_ (.Y(_08386_),
    .A(\TRNG.hash[246] ),
    .B(\TRNG.hash[235] ));
 sg13g2_xnor2_1 _16842_ (.Y(_08387_),
    .A(\TRNG.hash[255] ),
    .B(_08386_));
 sg13g2_nor2b_1 _16843_ (.A(_07458_),
    .B_N(_08387_),
    .Y(_08388_));
 sg13g2_xnor2_1 _16844_ (.Y(_08389_),
    .A(_07458_),
    .B(_08387_));
 sg13g2_nor2_1 _16845_ (.A(\TRNG.hash[201] ),
    .B(net5565),
    .Y(_08390_));
 sg13g2_a21oi_1 _16846_ (.A1(\TRNG.hash[201] ),
    .A2(net5565),
    .Y(_08391_),
    .B1(\TRNG.hash[169] ));
 sg13g2_nor2_1 _16847_ (.A(_08390_),
    .B(_08391_),
    .Y(_08392_));
 sg13g2_a21oi_1 _16848_ (.A1(_08389_),
    .A2(_08392_),
    .Y(_08393_),
    .B1(_08388_));
 sg13g2_nor2_1 _16849_ (.A(_08385_),
    .B(_08393_),
    .Y(_08394_));
 sg13g2_xnor2_1 _16850_ (.Y(_08395_),
    .A(_08385_),
    .B(_08393_));
 sg13g2_a21oi_1 _16851_ (.A1(_08362_),
    .A2(_08365_),
    .Y(_08396_),
    .B1(_08361_));
 sg13g2_xnor2_1 _16852_ (.Y(_08397_),
    .A(_08389_),
    .B(_08392_));
 sg13g2_and2_1 _16853_ (.A(_08396_),
    .B(_08397_),
    .X(_08398_));
 sg13g2_inv_1 _16854_ (.Y(_08399_),
    .A(_08398_));
 sg13g2_or2_1 _16855_ (.X(_08400_),
    .B(_08397_),
    .A(_08396_));
 sg13g2_nor2_1 _16856_ (.A(_08367_),
    .B(_08371_),
    .Y(_08401_));
 sg13g2_nor2b_1 _16857_ (.A(_08367_),
    .B_N(_08400_),
    .Y(_08402_));
 sg13g2_o21ai_1 _16858_ (.B1(_08402_),
    .Y(_08403_),
    .A1(_08369_),
    .A2(_08370_));
 sg13g2_nand2_1 _16859_ (.Y(_08404_),
    .A(_08399_),
    .B(_08403_));
 sg13g2_nor2_1 _16860_ (.A(_08395_),
    .B(_08404_),
    .Y(_08405_));
 sg13g2_nor2_1 _16861_ (.A(_08394_),
    .B(_08405_),
    .Y(_08406_));
 sg13g2_a21o_1 _16862_ (.A2(_08384_),
    .A1(_08381_),
    .B1(_08380_),
    .X(_08407_));
 sg13g2_xnor2_1 _16863_ (.Y(_08408_),
    .A(\TRNG.hash[225] ),
    .B(net5879));
 sg13g2_xnor2_1 _16864_ (.Y(_08409_),
    .A(\TRNG.hash[237] ),
    .B(_08408_));
 sg13g2_nand2_1 _16865_ (.Y(_08410_),
    .A(_07515_),
    .B(_08409_));
 sg13g2_xor2_1 _16866_ (.B(_08409_),
    .A(_07515_),
    .X(_08411_));
 sg13g2_a21oi_1 _16867_ (.A1(\TRNG.hash[235] ),
    .A2(\TRNG.hash[171] ),
    .Y(_08412_),
    .B1(\TRNG.hash[203] ));
 sg13g2_a21oi_1 _16868_ (.A1(_04283_),
    .A2(_04291_),
    .Y(_08413_),
    .B1(_08412_));
 sg13g2_nand2_1 _16869_ (.Y(_08414_),
    .A(_08411_),
    .B(_08413_));
 sg13g2_xnor2_1 _16870_ (.Y(_08415_),
    .A(_08411_),
    .B(_08413_));
 sg13g2_nand2b_1 _16871_ (.Y(_08416_),
    .B(_08415_),
    .A_N(_08407_));
 sg13g2_nor2b_1 _16872_ (.A(_08415_),
    .B_N(_08407_),
    .Y(_08417_));
 sg13g2_inv_1 _16873_ (.Y(_08418_),
    .A(_08417_));
 sg13g2_xnor2_1 _16874_ (.Y(_08419_),
    .A(_08407_),
    .B(_08415_));
 sg13g2_o21ai_1 _16875_ (.B1(net5818),
    .Y(_08420_),
    .A1(_08406_),
    .A2(_08419_));
 sg13g2_a21oi_1 _16876_ (.A1(_08406_),
    .A2(_08419_),
    .Y(_08421_),
    .B1(_08420_));
 sg13g2_o21ai_1 _16877_ (.B1(net3940),
    .Y(_08422_),
    .A1(net5565),
    .A2(_08375_));
 sg13g2_o21ai_1 _16878_ (.B1(net5571),
    .Y(_08423_),
    .A1(net5564),
    .A2(_08422_));
 sg13g2_xnor2_1 _16879_ (.Y(_08424_),
    .A(\TRNG.hash[235] ),
    .B(_08423_));
 sg13g2_o21ai_1 _16880_ (.B1(net4974),
    .Y(_08425_),
    .A1(net5819),
    .A2(_08424_));
 sg13g2_nor2_1 _16881_ (.A(_08421_),
    .B(_08425_),
    .Y(_00581_));
 sg13g2_nor2_1 _16882_ (.A(net5564),
    .B(net5565),
    .Y(_08426_));
 sg13g2_a21oi_1 _16883_ (.A1(_08375_),
    .A2(_08426_),
    .Y(_08427_),
    .B1(_04283_));
 sg13g2_nand2_1 _16884_ (.Y(_08428_),
    .A(net5571),
    .B(_08427_));
 sg13g2_xor2_1 _16885_ (.B(_08428_),
    .A(net5885),
    .X(_08429_));
 sg13g2_xnor2_1 _16886_ (.Y(_08430_),
    .A(\TRNG.hash[238] ),
    .B(net5568));
 sg13g2_xnor2_1 _16887_ (.Y(_08431_),
    .A(net5559),
    .B(_08430_));
 sg13g2_nor2b_1 _16888_ (.A(_07554_),
    .B_N(_08431_),
    .Y(_08432_));
 sg13g2_xnor2_1 _16889_ (.Y(_08433_),
    .A(_07554_),
    .B(_08431_));
 sg13g2_nor2_1 _16890_ (.A(\TRNG.hash[236] ),
    .B(\TRNG.hash[204] ),
    .Y(_08434_));
 sg13g2_a21oi_1 _16891_ (.A1(net5885),
    .A2(\TRNG.hash[204] ),
    .Y(_08435_),
    .B1(\TRNG.hash[172] ));
 sg13g2_nor2_1 _16892_ (.A(_08434_),
    .B(_08435_),
    .Y(_08436_));
 sg13g2_xnor2_1 _16893_ (.Y(_08437_),
    .A(_08433_),
    .B(_08436_));
 sg13g2_nand2_1 _16894_ (.Y(_08438_),
    .A(_08410_),
    .B(_08414_));
 sg13g2_a21oi_1 _16895_ (.A1(_08410_),
    .A2(_08414_),
    .Y(_08439_),
    .B1(_08437_));
 sg13g2_xor2_1 _16896_ (.B(_08438_),
    .A(_08437_),
    .X(_08440_));
 sg13g2_nand2_1 _16897_ (.Y(_08441_),
    .A(_08394_),
    .B(_08416_));
 sg13g2_nor2b_1 _16898_ (.A(_08395_),
    .B_N(_08419_),
    .Y(_08442_));
 sg13g2_nand3_1 _16899_ (.B(_08403_),
    .C(_08442_),
    .A(_08399_),
    .Y(_08443_));
 sg13g2_and3_1 _16900_ (.X(_08444_),
    .A(_08418_),
    .B(_08441_),
    .C(_08443_));
 sg13g2_nand3_1 _16901_ (.B(_08441_),
    .C(_08443_),
    .A(_08418_),
    .Y(_08445_));
 sg13g2_nand2_1 _16902_ (.Y(_08446_),
    .A(_08440_),
    .B(_08444_));
 sg13g2_nor2_1 _16903_ (.A(_08440_),
    .B(_08444_),
    .Y(_08447_));
 sg13g2_nand3b_1 _16904_ (.B(net4743),
    .C(_08446_),
    .Y(_08448_),
    .A_N(_08447_));
 sg13g2_o21ai_1 _16905_ (.B1(_08448_),
    .Y(_00582_),
    .A1(net4747),
    .A2(_08429_));
 sg13g2_xnor2_1 _16906_ (.Y(_08449_),
    .A(\TRNG.hash[230] ),
    .B(net5883));
 sg13g2_xnor2_1 _16907_ (.Y(_08450_),
    .A(net5557),
    .B(_08449_));
 sg13g2_xnor2_1 _16908_ (.Y(_08451_),
    .A(_07676_),
    .B(_08450_));
 sg13g2_a21oi_1 _16909_ (.A1(\TRNG.hash[240] ),
    .A2(\TRNG.hash[176] ),
    .Y(_08452_),
    .B1(\TRNG.hash[208] ));
 sg13g2_a21oi_1 _16910_ (.A1(_04226_),
    .A2(_04290_),
    .Y(_08453_),
    .B1(_08452_));
 sg13g2_nor2b_1 _16911_ (.A(_08451_),
    .B_N(_08453_),
    .Y(_08454_));
 sg13g2_a21o_1 _16912_ (.A2(_08450_),
    .A1(_07676_),
    .B1(_08454_),
    .X(_08455_));
 sg13g2_xnor2_1 _16913_ (.Y(_08456_),
    .A(net5560),
    .B(\TRNG.hash[231] ));
 sg13g2_xnor2_1 _16914_ (.Y(_08457_),
    .A(net5556),
    .B(_08456_));
 sg13g2_nand2_1 _16915_ (.Y(_08458_),
    .A(_07754_),
    .B(_08457_));
 sg13g2_nor2_1 _16916_ (.A(_07754_),
    .B(_08457_),
    .Y(_08459_));
 sg13g2_xor2_1 _16917_ (.B(_08457_),
    .A(_07753_),
    .X(_08460_));
 sg13g2_a21o_1 _16918_ (.A2(\TRNG.hash[241] ),
    .A1(\TRNG.hash[209] ),
    .B1(\TRNG.hash[177] ),
    .X(_08461_));
 sg13g2_o21ai_1 _16919_ (.B1(_08461_),
    .Y(_08462_),
    .A1(\TRNG.hash[209] ),
    .A2(\TRNG.hash[241] ));
 sg13g2_xnor2_1 _16920_ (.Y(_08463_),
    .A(_08460_),
    .B(_08462_));
 sg13g2_nor2b_1 _16921_ (.A(_08455_),
    .B_N(_08463_),
    .Y(_08464_));
 sg13g2_nand2b_1 _16922_ (.Y(_08465_),
    .B(_08455_),
    .A_N(_08463_));
 sg13g2_nor2b_1 _16923_ (.A(_08464_),
    .B_N(_08465_),
    .Y(_08466_));
 sg13g2_xnor2_1 _16924_ (.Y(_08467_),
    .A(_08451_),
    .B(_08453_));
 sg13g2_xnor2_1 _16925_ (.Y(_08468_),
    .A(net5877),
    .B(net5884));
 sg13g2_xnor2_1 _16926_ (.Y(_08469_),
    .A(\TRNG.hash[229] ),
    .B(_08468_));
 sg13g2_nor2b_1 _16927_ (.A(_07633_),
    .B_N(_08469_),
    .Y(_08470_));
 sg13g2_xnor2_1 _16928_ (.Y(_08471_),
    .A(_07633_),
    .B(_08469_));
 sg13g2_nor2_1 _16929_ (.A(\TRNG.hash[207] ),
    .B(net5561),
    .Y(_08472_));
 sg13g2_a21oi_1 _16930_ (.A1(\TRNG.hash[207] ),
    .A2(net5561),
    .Y(_08473_),
    .B1(\TRNG.hash[175] ));
 sg13g2_nor2_1 _16931_ (.A(_08472_),
    .B(_08473_),
    .Y(_08474_));
 sg13g2_a21oi_1 _16932_ (.A1(_08471_),
    .A2(_08474_),
    .Y(_08475_),
    .B1(_08470_));
 sg13g2_nand2b_1 _16933_ (.Y(_08476_),
    .B(_08467_),
    .A_N(_08475_));
 sg13g2_xnor2_1 _16934_ (.Y(_08477_),
    .A(\TRNG.hash[240] ),
    .B(\TRNG.hash[228] ));
 sg13g2_xnor2_1 _16935_ (.Y(_08478_),
    .A(net5558),
    .B(_08477_));
 sg13g2_nor2b_1 _16936_ (.A(_07636_),
    .B_N(_08478_),
    .Y(_08479_));
 sg13g2_xnor2_1 _16937_ (.Y(_08480_),
    .A(_07636_),
    .B(_08478_));
 sg13g2_nor2_1 _16938_ (.A(net5562),
    .B(\TRNG.hash[206] ),
    .Y(_08481_));
 sg13g2_a21oi_1 _16939_ (.A1(net5562),
    .A2(\TRNG.hash[206] ),
    .Y(_08482_),
    .B1(\TRNG.hash[174] ));
 sg13g2_nor2_1 _16940_ (.A(_08481_),
    .B(_08482_),
    .Y(_08483_));
 sg13g2_xnor2_1 _16941_ (.Y(_08484_),
    .A(_08480_),
    .B(_08483_));
 sg13g2_xnor2_1 _16942_ (.Y(_08485_),
    .A(net5878),
    .B(net5888));
 sg13g2_xnor2_1 _16943_ (.Y(_08486_),
    .A(\TRNG.hash[239] ),
    .B(_08485_));
 sg13g2_nand2b_1 _16944_ (.Y(_08487_),
    .B(_08486_),
    .A_N(_07580_));
 sg13g2_xnor2_1 _16945_ (.Y(_08488_),
    .A(_07580_),
    .B(_08486_));
 sg13g2_nor2_1 _16946_ (.A(\TRNG.hash[205] ),
    .B(net5563),
    .Y(_08489_));
 sg13g2_a21oi_1 _16947_ (.A1(\TRNG.hash[205] ),
    .A2(net5563),
    .Y(_08490_),
    .B1(\TRNG.hash[173] ));
 sg13g2_nor2_1 _16948_ (.A(_08489_),
    .B(_08490_),
    .Y(_08491_));
 sg13g2_nand2_1 _16949_ (.Y(_08492_),
    .A(_08488_),
    .B(_08491_));
 sg13g2_a21oi_1 _16950_ (.A1(_08487_),
    .A2(_08492_),
    .Y(_08493_),
    .B1(_08484_));
 sg13g2_inv_1 _16951_ (.Y(_08494_),
    .A(_08493_));
 sg13g2_nand3_1 _16952_ (.B(_08487_),
    .C(_08492_),
    .A(_08484_),
    .Y(_08495_));
 sg13g2_nand2_1 _16953_ (.Y(_08496_),
    .A(_08494_),
    .B(_08495_));
 sg13g2_a21o_1 _16954_ (.A2(_08483_),
    .A1(_08480_),
    .B1(_08479_),
    .X(_08497_));
 sg13g2_xnor2_1 _16955_ (.Y(_08498_),
    .A(_08471_),
    .B(_08474_));
 sg13g2_nor2b_1 _16956_ (.A(_08497_),
    .B_N(_08498_),
    .Y(_08499_));
 sg13g2_nand2b_1 _16957_ (.Y(_08500_),
    .B(_08497_),
    .A_N(_08498_));
 sg13g2_nand2b_1 _16958_ (.Y(_08501_),
    .B(_08500_),
    .A_N(_08499_));
 sg13g2_nor2_1 _16959_ (.A(_08496_),
    .B(_08501_),
    .Y(_08502_));
 sg13g2_a21o_1 _16960_ (.A2(_08436_),
    .A1(_08433_),
    .B1(_08432_),
    .X(_08503_));
 sg13g2_xnor2_1 _16961_ (.Y(_08504_),
    .A(_08488_),
    .B(_08491_));
 sg13g2_nor2b_1 _16962_ (.A(_08504_),
    .B_N(_08503_),
    .Y(_08505_));
 sg13g2_nand2b_1 _16963_ (.Y(_08506_),
    .B(_08504_),
    .A_N(_08503_));
 sg13g2_nor2b_1 _16964_ (.A(_08505_),
    .B_N(_08506_),
    .Y(_08507_));
 sg13g2_nor2b_1 _16965_ (.A(_08440_),
    .B_N(_08507_),
    .Y(_08508_));
 sg13g2_and2_1 _16966_ (.A(_08502_),
    .B(_08508_),
    .X(_08509_));
 sg13g2_nand2_1 _16967_ (.Y(_08510_),
    .A(_08502_),
    .B(_08508_));
 sg13g2_a21o_1 _16968_ (.A2(_08506_),
    .A1(_08439_),
    .B1(_08505_),
    .X(_08511_));
 sg13g2_a21oi_1 _16969_ (.A1(_08494_),
    .A2(_08500_),
    .Y(_08512_),
    .B1(_08499_));
 sg13g2_a21oi_1 _16970_ (.A1(_08502_),
    .A2(_08511_),
    .Y(_08513_),
    .B1(_08512_));
 sg13g2_a221oi_1 _16971_ (.B2(_08502_),
    .C1(_08512_),
    .B1(_08511_),
    .A1(_08445_),
    .Y(_08514_),
    .A2(_08509_));
 sg13g2_o21ai_1 _16972_ (.B1(_08513_),
    .Y(_08515_),
    .A1(_08444_),
    .A2(_08510_));
 sg13g2_xor2_1 _16973_ (.B(_08475_),
    .A(_08467_),
    .X(_08516_));
 sg13g2_inv_1 _16974_ (.Y(_08517_),
    .A(_08516_));
 sg13g2_o21ai_1 _16975_ (.B1(_08476_),
    .Y(_08518_),
    .A1(_08514_),
    .A2(_08516_));
 sg13g2_xnor2_1 _16976_ (.Y(_08519_),
    .A(_08466_),
    .B(_08518_));
 sg13g2_nand2_2 _16977_ (.Y(_08520_),
    .A(net5885),
    .B(_08427_));
 sg13g2_nor3_1 _16978_ (.A(net5561),
    .B(net5562),
    .C(net5563),
    .Y(_08521_));
 sg13g2_nand2_1 _16979_ (.Y(_08522_),
    .A(_08520_),
    .B(_08521_));
 sg13g2_nand3_1 _16980_ (.B(_08520_),
    .C(_08521_),
    .A(_04226_),
    .Y(_08523_));
 sg13g2_xnor2_1 _16981_ (.Y(_08524_),
    .A(net5884),
    .B(_08523_));
 sg13g2_o21ai_1 _16982_ (.B1(net4973),
    .Y(_08525_),
    .A1(net5884),
    .A2(net5174));
 sg13g2_a221oi_1 _16983_ (.B2(net5182),
    .C1(_08525_),
    .B1(_08524_),
    .A1(net5823),
    .Y(_00583_),
    .A2(_08519_));
 sg13g2_xnor2_1 _16984_ (.Y(_08526_),
    .A(net5882),
    .B(\TRNG.hash[232] ));
 sg13g2_xnor2_1 _16985_ (.Y(_08527_),
    .A(\TRNG.hash[255] ),
    .B(_08526_));
 sg13g2_nor2b_1 _16986_ (.A(_07748_),
    .B_N(_08527_),
    .Y(_08528_));
 sg13g2_xnor2_1 _16987_ (.Y(_08529_),
    .A(_07748_),
    .B(_08527_));
 sg13g2_nor2_1 _16988_ (.A(\TRNG.hash[210] ),
    .B(\TRNG.hash[242] ),
    .Y(_08530_));
 sg13g2_a21oi_1 _16989_ (.A1(\TRNG.hash[210] ),
    .A2(\TRNG.hash[242] ),
    .Y(_08531_),
    .B1(\TRNG.hash[178] ));
 sg13g2_nor2_1 _16990_ (.A(_08530_),
    .B(_08531_),
    .Y(_08532_));
 sg13g2_xnor2_1 _16991_ (.Y(_08533_),
    .A(_08529_),
    .B(_08532_));
 sg13g2_o21ai_1 _16992_ (.B1(_08458_),
    .Y(_08534_),
    .A1(_08459_),
    .A2(_08462_));
 sg13g2_nor2b_1 _16993_ (.A(_08533_),
    .B_N(_08534_),
    .Y(_08535_));
 sg13g2_xor2_1 _16994_ (.B(_08534_),
    .A(_08533_),
    .X(_08536_));
 sg13g2_o21ai_1 _16995_ (.B1(_08465_),
    .Y(_08537_),
    .A1(_08464_),
    .A2(_08476_));
 sg13g2_inv_1 _16996_ (.Y(_08538_),
    .A(_08537_));
 sg13g2_nand2_1 _16997_ (.Y(_08539_),
    .A(_08466_),
    .B(_08517_));
 sg13g2_o21ai_1 _16998_ (.B1(_08538_),
    .Y(_08540_),
    .A1(_08514_),
    .A2(_08539_));
 sg13g2_nor2b_1 _16999_ (.A(_08536_),
    .B_N(_08540_),
    .Y(_08541_));
 sg13g2_xor2_1 _17000_ (.B(_08540_),
    .A(_08536_),
    .X(_08542_));
 sg13g2_nand3_1 _17001_ (.B(net5884),
    .C(_08523_),
    .A(net5883),
    .Y(_08543_));
 sg13g2_a21o_1 _17002_ (.A2(_08523_),
    .A1(net5884),
    .B1(net5883),
    .X(_08544_));
 sg13g2_nand2_1 _17003_ (.Y(_08545_),
    .A(_08543_),
    .B(_08544_));
 sg13g2_o21ai_1 _17004_ (.B1(net4973),
    .Y(_08546_),
    .A1(net5883),
    .A2(net5174));
 sg13g2_a221oi_1 _17005_ (.B2(net5182),
    .C1(_08546_),
    .B1(_08545_),
    .A1(net5825),
    .Y(_00584_),
    .A2(_08542_));
 sg13g2_xnor2_1 _17006_ (.Y(_08547_),
    .A(net5569),
    .B(\TRNG.hash[246] ));
 sg13g2_xnor2_1 _17007_ (.Y(_08548_),
    .A(\TRNG.hash[234] ),
    .B(_08547_));
 sg13g2_nor2b_1 _17008_ (.A(_07793_),
    .B_N(_08548_),
    .Y(_08549_));
 sg13g2_xnor2_1 _17009_ (.Y(_08550_),
    .A(_07793_),
    .B(_08548_));
 sg13g2_a21oi_1 _17010_ (.A1(\TRNG.hash[212] ),
    .A2(\TRNG.hash[180] ),
    .Y(_08551_),
    .B1(net5882));
 sg13g2_a21oi_1 _17011_ (.A1(_04287_),
    .A2(_04289_),
    .Y(_08552_),
    .B1(_08551_));
 sg13g2_xnor2_1 _17012_ (.Y(_08553_),
    .A(_08550_),
    .B(_08552_));
 sg13g2_xnor2_1 _17013_ (.Y(_08554_),
    .A(\TRNG.hash[224] ),
    .B(net5881));
 sg13g2_xnor2_1 _17014_ (.Y(_08555_),
    .A(\TRNG.hash[233] ),
    .B(_08554_));
 sg13g2_nor2b_1 _17015_ (.A(_07744_),
    .B_N(_08555_),
    .Y(_08556_));
 sg13g2_xnor2_1 _17016_ (.Y(_08557_),
    .A(_07744_),
    .B(_08555_));
 sg13g2_nor2_1 _17017_ (.A(\TRNG.hash[243] ),
    .B(\TRNG.hash[211] ),
    .Y(_08558_));
 sg13g2_a21oi_1 _17018_ (.A1(net5560),
    .A2(\TRNG.hash[211] ),
    .Y(_08559_),
    .B1(\TRNG.hash[179] ));
 sg13g2_nor2_1 _17019_ (.A(_08558_),
    .B(_08559_),
    .Y(_08560_));
 sg13g2_a21o_1 _17020_ (.A2(_08560_),
    .A1(_08557_),
    .B1(_08556_),
    .X(_08561_));
 sg13g2_nand2b_1 _17021_ (.Y(_08562_),
    .B(_08561_),
    .A_N(_08553_));
 sg13g2_xnor2_1 _17022_ (.Y(_08563_),
    .A(_08553_),
    .B(_08561_));
 sg13g2_a21o_1 _17023_ (.A2(_08532_),
    .A1(_08529_),
    .B1(_08528_),
    .X(_08564_));
 sg13g2_xnor2_1 _17024_ (.Y(_08565_),
    .A(_08557_),
    .B(_08560_));
 sg13g2_nor2b_1 _17025_ (.A(_08565_),
    .B_N(_08564_),
    .Y(_08566_));
 sg13g2_nand2b_1 _17026_ (.Y(_08567_),
    .B(_08565_),
    .A_N(_08564_));
 sg13g2_nor2b_1 _17027_ (.A(_08566_),
    .B_N(_08567_),
    .Y(_08568_));
 sg13g2_nor2b_1 _17028_ (.A(_08536_),
    .B_N(_08568_),
    .Y(_08569_));
 sg13g2_a221oi_1 _17029_ (.B2(_08537_),
    .C1(_08566_),
    .B1(_08569_),
    .A1(_08535_),
    .Y(_08570_),
    .A2(_08567_));
 sg13g2_nand3_1 _17030_ (.B(_08517_),
    .C(_08569_),
    .A(_08466_),
    .Y(_08571_));
 sg13g2_o21ai_1 _17031_ (.B1(_08570_),
    .Y(_08572_),
    .A1(_08514_),
    .A2(_08571_));
 sg13g2_nand2_1 _17032_ (.Y(_08573_),
    .A(_08563_),
    .B(_08572_));
 sg13g2_xnor2_1 _17033_ (.Y(_08574_),
    .A(_08563_),
    .B(_08572_));
 sg13g2_o21ai_1 _17034_ (.B1(net3795),
    .Y(_08575_),
    .A1(net5560),
    .A2(_08543_));
 sg13g2_and2_1 _17035_ (.A(net5882),
    .B(_08575_),
    .X(_08576_));
 sg13g2_xnor2_1 _17036_ (.Y(_08577_),
    .A(net5882),
    .B(_08575_));
 sg13g2_o21ai_1 _17037_ (.B1(net4973),
    .Y(_08578_),
    .A1(net5882),
    .A2(net5174));
 sg13g2_a221oi_1 _17038_ (.B2(net5183),
    .C1(_08578_),
    .B1(_08577_),
    .A1(net5826),
    .Y(_00585_),
    .A2(_08574_));
 sg13g2_a21o_1 _17039_ (.A2(_08552_),
    .A1(_08550_),
    .B1(_08549_),
    .X(_08579_));
 sg13g2_xnor2_1 _17040_ (.Y(_08580_),
    .A(net5880),
    .B(\TRNG.hash[235] ));
 sg13g2_xnor2_1 _17041_ (.Y(_08581_),
    .A(net5568),
    .B(_08580_));
 sg13g2_xor2_1 _17042_ (.B(_08581_),
    .A(_07818_),
    .X(_08582_));
 sg13g2_a21oi_1 _17043_ (.A1(\TRNG.hash[213] ),
    .A2(net5881),
    .Y(_08583_),
    .B1(\TRNG.hash[181] ));
 sg13g2_a21oi_1 _17044_ (.A1(_04224_),
    .A2(_04282_),
    .Y(_08584_),
    .B1(_08583_));
 sg13g2_nor2b_1 _17045_ (.A(_08582_),
    .B_N(_08584_),
    .Y(_08585_));
 sg13g2_xor2_1 _17046_ (.B(_08584_),
    .A(_08582_),
    .X(_08586_));
 sg13g2_nor2b_1 _17047_ (.A(_08579_),
    .B_N(_08586_),
    .Y(_08587_));
 sg13g2_nand2b_1 _17048_ (.Y(_08588_),
    .B(_08586_),
    .A_N(_08579_));
 sg13g2_nand2b_1 _17049_ (.Y(_08589_),
    .B(_08579_),
    .A_N(_08586_));
 sg13g2_and2_1 _17050_ (.A(_08588_),
    .B(_08589_),
    .X(_08590_));
 sg13g2_nand2_1 _17051_ (.Y(_08591_),
    .A(_08562_),
    .B(_08573_));
 sg13g2_xnor2_1 _17052_ (.Y(_08592_),
    .A(_08590_),
    .B(_08591_));
 sg13g2_nand2_1 _17053_ (.Y(_08593_),
    .A(net5881),
    .B(_08576_));
 sg13g2_xnor2_1 _17054_ (.Y(_08594_),
    .A(net3499),
    .B(_08576_));
 sg13g2_o21ai_1 _17055_ (.B1(net4973),
    .Y(_08595_),
    .A1(net3499),
    .A2(net5174));
 sg13g2_a221oi_1 _17056_ (.B2(net5184),
    .C1(_08595_),
    .B1(_08594_),
    .A1(net5839),
    .Y(_00586_),
    .A2(_08592_));
 sg13g2_xnor2_1 _17057_ (.Y(_08596_),
    .A(net5885),
    .B(net5888));
 sg13g2_xnor2_1 _17058_ (.Y(_08597_),
    .A(net5879),
    .B(_08596_));
 sg13g2_nor2b_1 _17059_ (.A(_07858_),
    .B_N(_08597_),
    .Y(_08598_));
 sg13g2_xnor2_1 _17060_ (.Y(_08599_),
    .A(_07858_),
    .B(_08597_));
 sg13g2_a21oi_1 _17061_ (.A1(\TRNG.hash[214] ),
    .A2(\TRNG.hash[246] ),
    .Y(_08600_),
    .B1(\TRNG.hash[182] ));
 sg13g2_a21oi_2 _17062_ (.B1(_08600_),
    .Y(_08601_),
    .A2(_04281_),
    .A1(_04223_));
 sg13g2_xnor2_1 _17063_ (.Y(_08602_),
    .A(_08599_),
    .B(_08601_));
 sg13g2_a21oi_1 _17064_ (.A1(_07819_),
    .A2(_08581_),
    .Y(_08603_),
    .B1(_08585_));
 sg13g2_nor2_1 _17065_ (.A(_08602_),
    .B(_08603_),
    .Y(_08604_));
 sg13g2_inv_1 _17066_ (.Y(_08605_),
    .A(_08604_));
 sg13g2_xnor2_1 _17067_ (.Y(_08606_),
    .A(_08602_),
    .B(_08603_));
 sg13g2_and3_1 _17068_ (.X(_08607_),
    .A(_08563_),
    .B(_08588_),
    .C(_08589_));
 sg13g2_a21oi_1 _17069_ (.A1(_08562_),
    .A2(_08589_),
    .Y(_08608_),
    .B1(_08587_));
 sg13g2_a21oi_1 _17070_ (.A1(_08572_),
    .A2(_08607_),
    .Y(_08609_),
    .B1(_08608_));
 sg13g2_xnor2_1 _17071_ (.Y(_08610_),
    .A(_08606_),
    .B(_08609_));
 sg13g2_nor2_1 _17072_ (.A(_04281_),
    .B(_08593_),
    .Y(_08611_));
 sg13g2_xnor2_1 _17073_ (.Y(_08612_),
    .A(_04281_),
    .B(_08593_));
 sg13g2_o21ai_1 _17074_ (.B1(net4974),
    .Y(_08613_),
    .A1(net3901),
    .A2(net5174));
 sg13g2_a221oi_1 _17075_ (.B2(net5184),
    .C1(_08613_),
    .B1(_08612_),
    .A1(net5839),
    .Y(_00587_),
    .A2(_08610_));
 sg13g2_and2_1 _17076_ (.A(net5880),
    .B(_08611_),
    .X(_08614_));
 sg13g2_o21ai_1 _17077_ (.B1(net5572),
    .Y(_08615_),
    .A1(net5880),
    .A2(_08611_));
 sg13g2_o21ai_1 _17078_ (.B1(net5486),
    .Y(_08616_),
    .A1(_08614_),
    .A2(_08615_));
 sg13g2_a21oi_2 _17079_ (.B1(_08598_),
    .Y(_08617_),
    .A2(_08601_),
    .A1(_08599_));
 sg13g2_xnor2_1 _17080_ (.Y(_08618_),
    .A(net5563),
    .B(net5887));
 sg13g2_xnor2_1 _17081_ (.Y(_08619_),
    .A(net5559),
    .B(_08618_));
 sg13g2_and2_1 _17082_ (.A(_07886_),
    .B(_08619_),
    .X(_08620_));
 sg13g2_xor2_1 _17083_ (.B(_08619_),
    .A(_07886_),
    .X(_08621_));
 sg13g2_nor2_1 _17084_ (.A(\TRNG.hash[215] ),
    .B(\TRNG.hash[183] ),
    .Y(_08622_));
 sg13g2_a21oi_1 _17085_ (.A1(\TRNG.hash[215] ),
    .A2(\TRNG.hash[183] ),
    .Y(_08623_),
    .B1(net5880));
 sg13g2_nor2_1 _17086_ (.A(_08622_),
    .B(_08623_),
    .Y(_08624_));
 sg13g2_xnor2_1 _17087_ (.Y(_08625_),
    .A(_08621_),
    .B(_08624_));
 sg13g2_nand2_1 _17088_ (.Y(_08626_),
    .A(_08617_),
    .B(_08625_));
 sg13g2_nor2_1 _17089_ (.A(_08617_),
    .B(_08625_),
    .Y(_08627_));
 sg13g2_xor2_1 _17090_ (.B(_08625_),
    .A(_08617_),
    .X(_08628_));
 sg13g2_o21ai_1 _17091_ (.B1(_08605_),
    .Y(_08629_),
    .A1(_08606_),
    .A2(_08609_));
 sg13g2_xor2_1 _17092_ (.B(_08629_),
    .A(_08628_),
    .X(_08630_));
 sg13g2_o21ai_1 _17093_ (.B1(_08616_),
    .Y(_08631_),
    .A1(net5486),
    .A2(_08630_));
 sg13g2_nand2_1 _17094_ (.Y(_08632_),
    .A(net5880),
    .B(net5347));
 sg13g2_a21oi_1 _17095_ (.A1(_08631_),
    .A2(_08632_),
    .Y(_00588_),
    .B1(net4962));
 sg13g2_nor2b_1 _17096_ (.A(_08606_),
    .B_N(_08628_),
    .Y(_08633_));
 sg13g2_nand2_1 _17097_ (.Y(_08634_),
    .A(_08607_),
    .B(_08633_));
 sg13g2_nor2_1 _17098_ (.A(_08571_),
    .B(_08634_),
    .Y(_08635_));
 sg13g2_a221oi_1 _17099_ (.B2(_08608_),
    .C1(_08627_),
    .B1(_08633_),
    .A1(_08604_),
    .Y(_08636_),
    .A2(_08626_));
 sg13g2_o21ai_1 _17100_ (.B1(_08636_),
    .Y(_08637_),
    .A1(_08570_),
    .A2(_08634_));
 sg13g2_a21oi_2 _17101_ (.B1(_08637_),
    .Y(_08638_),
    .A2(_08635_),
    .A1(_08515_));
 sg13g2_a21o_1 _17102_ (.A2(_08635_),
    .A1(_08515_),
    .B1(_08637_),
    .X(_08639_));
 sg13g2_xnor2_1 _17103_ (.Y(_08640_),
    .A(net5567),
    .B(net5878));
 sg13g2_xnor2_1 _17104_ (.Y(_08641_),
    .A(\TRNG.hash[238] ),
    .B(_08640_));
 sg13g2_xnor2_1 _17105_ (.Y(_08642_),
    .A(_07941_),
    .B(_08641_));
 sg13g2_nor2_1 _17106_ (.A(\TRNG.hash[248] ),
    .B(\TRNG.hash[184] ),
    .Y(_08643_));
 sg13g2_a21oi_1 _17107_ (.A1(\TRNG.hash[248] ),
    .A2(\TRNG.hash[184] ),
    .Y(_08644_),
    .B1(\TRNG.hash[216] ));
 sg13g2_nor2_1 _17108_ (.A(_08643_),
    .B(_08644_),
    .Y(_08645_));
 sg13g2_nor2b_1 _17109_ (.A(_08642_),
    .B_N(_08645_),
    .Y(_08646_));
 sg13g2_xnor2_1 _17110_ (.Y(_08647_),
    .A(_08642_),
    .B(_08645_));
 sg13g2_a21oi_1 _17111_ (.A1(_08621_),
    .A2(_08624_),
    .Y(_08648_),
    .B1(_08620_));
 sg13g2_nor2b_1 _17112_ (.A(_08648_),
    .B_N(_08647_),
    .Y(_08649_));
 sg13g2_xor2_1 _17113_ (.B(_08648_),
    .A(_08647_),
    .X(_08650_));
 sg13g2_nor2_1 _17114_ (.A(_08638_),
    .B(_08650_),
    .Y(_08651_));
 sg13g2_xnor2_1 _17115_ (.Y(_08652_),
    .A(_08638_),
    .B(_08650_));
 sg13g2_and2_1 _17116_ (.A(net5879),
    .B(_08614_),
    .X(_08653_));
 sg13g2_inv_1 _17117_ (.Y(_08654_),
    .A(_08653_));
 sg13g2_xnor2_1 _17118_ (.Y(_08655_),
    .A(net5879),
    .B(_08614_));
 sg13g2_o21ai_1 _17119_ (.B1(net4973),
    .Y(_08656_),
    .A1(net5879),
    .A2(net5175));
 sg13g2_a221oi_1 _17120_ (.B2(net5184),
    .C1(_08656_),
    .B1(_08655_),
    .A1(net5839),
    .Y(_00589_),
    .A2(_08652_));
 sg13g2_xnor2_1 _17121_ (.Y(_08657_),
    .A(net5877),
    .B(\TRNG.hash[231] ));
 sg13g2_xnor2_1 _17122_ (.Y(_08658_),
    .A(\TRNG.hash[240] ),
    .B(_08657_));
 sg13g2_xnor2_1 _17123_ (.Y(_08659_),
    .A(_07982_),
    .B(_08658_));
 sg13g2_a21oi_1 _17124_ (.A1(\TRNG.hash[250] ),
    .A2(\TRNG.hash[218] ),
    .Y(_08660_),
    .B1(\TRNG.hash[186] ));
 sg13g2_a21oi_1 _17125_ (.A1(_04280_),
    .A2(_04286_),
    .Y(_08661_),
    .B1(_08660_));
 sg13g2_nor2b_1 _17126_ (.A(_08659_),
    .B_N(_08661_),
    .Y(_08662_));
 sg13g2_xnor2_1 _17127_ (.Y(_08663_),
    .A(_08659_),
    .B(_08661_));
 sg13g2_xnor2_1 _17128_ (.Y(_08664_),
    .A(net5561),
    .B(net5566));
 sg13g2_xnor2_1 _17129_ (.Y(_08665_),
    .A(net5558),
    .B(_08664_));
 sg13g2_nand2_1 _17130_ (.Y(_08666_),
    .A(_07937_),
    .B(_08665_));
 sg13g2_xnor2_1 _17131_ (.Y(_08667_),
    .A(_07937_),
    .B(_08665_));
 sg13g2_nor2_1 _17132_ (.A(\TRNG.hash[249] ),
    .B(\TRNG.hash[185] ),
    .Y(_08668_));
 sg13g2_a21oi_1 _17133_ (.A1(\TRNG.hash[249] ),
    .A2(\TRNG.hash[185] ),
    .Y(_08669_),
    .B1(\TRNG.hash[217] ));
 sg13g2_nor2_1 _17134_ (.A(_08668_),
    .B(_08669_),
    .Y(_08670_));
 sg13g2_inv_1 _17135_ (.Y(_08671_),
    .A(_08670_));
 sg13g2_o21ai_1 _17136_ (.B1(_08666_),
    .Y(_08672_),
    .A1(_08667_),
    .A2(_08671_));
 sg13g2_and2_1 _17137_ (.A(_08663_),
    .B(_08672_),
    .X(_08673_));
 sg13g2_xor2_1 _17138_ (.B(_08672_),
    .A(_08663_),
    .X(_08674_));
 sg13g2_a21oi_2 _17139_ (.B1(_08646_),
    .Y(_08675_),
    .A2(_08641_),
    .A1(_07941_));
 sg13g2_xnor2_1 _17140_ (.Y(_08676_),
    .A(_08667_),
    .B(_08670_));
 sg13g2_nand2b_1 _17141_ (.Y(_08677_),
    .B(_08675_),
    .A_N(_08676_));
 sg13g2_nor2b_1 _17142_ (.A(_08675_),
    .B_N(_08676_),
    .Y(_08678_));
 sg13g2_a21oi_1 _17143_ (.A1(_08649_),
    .A2(_08677_),
    .Y(_08679_),
    .B1(_08678_));
 sg13g2_xor2_1 _17144_ (.B(_08676_),
    .A(_08675_),
    .X(_08680_));
 sg13g2_or2_1 _17145_ (.X(_08681_),
    .B(_08680_),
    .A(_08650_));
 sg13g2_o21ai_1 _17146_ (.B1(_08679_),
    .Y(_08682_),
    .A1(_08638_),
    .A2(_08681_));
 sg13g2_xnor2_1 _17147_ (.Y(_08683_),
    .A(_08674_),
    .B(_08682_));
 sg13g2_o21ai_1 _17148_ (.B1(net3741),
    .Y(_08684_),
    .A1(net5559),
    .A2(_08654_));
 sg13g2_nand2_1 _17149_ (.Y(_08685_),
    .A(net5878),
    .B(_08684_));
 sg13g2_xnor2_1 _17150_ (.Y(_08686_),
    .A(net5878),
    .B(_08684_));
 sg13g2_o21ai_1 _17151_ (.B1(net4973),
    .Y(_08687_),
    .A1(net5878),
    .A2(net5174));
 sg13g2_a221oi_1 _17152_ (.B2(net5184),
    .C1(_08687_),
    .B1(_08686_),
    .A1(net5838),
    .Y(_00590_),
    .A2(_08683_));
 sg13g2_a21oi_2 _17153_ (.B1(_08662_),
    .Y(_08688_),
    .A2(_08658_),
    .A1(_07982_));
 sg13g2_xnor2_1 _17154_ (.Y(_08689_),
    .A(net5884),
    .B(net5886));
 sg13g2_xnor2_1 _17155_ (.Y(_08690_),
    .A(net5557),
    .B(_08689_));
 sg13g2_nor2b_1 _17156_ (.A(_08012_),
    .B_N(_08690_),
    .Y(_08691_));
 sg13g2_xnor2_1 _17157_ (.Y(_08692_),
    .A(_08012_),
    .B(_08690_));
 sg13g2_nor2_1 _17158_ (.A(\TRNG.hash[219] ),
    .B(net5558),
    .Y(_08693_));
 sg13g2_a21oi_1 _17159_ (.A1(\TRNG.hash[219] ),
    .A2(net5558),
    .Y(_08694_),
    .B1(\TRNG.hash[187] ));
 sg13g2_nor2_1 _17160_ (.A(_08693_),
    .B(_08694_),
    .Y(_08695_));
 sg13g2_xnor2_1 _17161_ (.Y(_08696_),
    .A(_08692_),
    .B(_08695_));
 sg13g2_or2_1 _17162_ (.X(_08697_),
    .B(_08696_),
    .A(_08688_));
 sg13g2_nand2_1 _17163_ (.Y(_08698_),
    .A(_08688_),
    .B(_08696_));
 sg13g2_xor2_1 _17164_ (.B(_08696_),
    .A(_08688_),
    .X(_08699_));
 sg13g2_inv_1 _17165_ (.Y(_08700_),
    .A(_08699_));
 sg13g2_nand2_1 _17166_ (.Y(_08701_),
    .A(_08674_),
    .B(_08699_));
 sg13g2_nor2_1 _17167_ (.A(_08681_),
    .B(_08701_),
    .Y(_08702_));
 sg13g2_or2_1 _17168_ (.X(_08703_),
    .B(_08701_),
    .A(_08681_));
 sg13g2_o21ai_1 _17169_ (.B1(_08697_),
    .Y(_08704_),
    .A1(_08679_),
    .A2(_08701_));
 sg13g2_a21oi_1 _17170_ (.A1(_08673_),
    .A2(_08698_),
    .Y(_08705_),
    .B1(_08704_));
 sg13g2_a221oi_1 _17171_ (.B2(_08639_),
    .C1(_08704_),
    .B1(_08702_),
    .A1(_08673_),
    .Y(_08706_),
    .A2(_08698_));
 sg13g2_o21ai_1 _17172_ (.B1(_08705_),
    .Y(_08707_),
    .A1(_08638_),
    .A2(_08703_));
 sg13g2_xnor2_1 _17173_ (.Y(_08708_),
    .A(net5565),
    .B(net5883));
 sg13g2_xnor2_1 _17174_ (.Y(_08709_),
    .A(net5556),
    .B(_08708_));
 sg13g2_nor2b_1 _17175_ (.A(_08041_),
    .B_N(_08709_),
    .Y(_08710_));
 sg13g2_xor2_1 _17176_ (.B(_08709_),
    .A(_08041_),
    .X(_08711_));
 sg13g2_a21o_1 _17177_ (.A2(net5877),
    .A1(\TRNG.hash[220] ),
    .B1(\TRNG.hash[188] ),
    .X(_08712_));
 sg13g2_o21ai_1 _17178_ (.B1(_08712_),
    .Y(_08713_),
    .A1(\TRNG.hash[220] ),
    .A2(net5877));
 sg13g2_nor2_1 _17179_ (.A(_08711_),
    .B(_08713_),
    .Y(_08714_));
 sg13g2_xnor2_1 _17180_ (.Y(_08715_),
    .A(_08711_),
    .B(_08713_));
 sg13g2_a21oi_2 _17181_ (.B1(_08691_),
    .Y(_08716_),
    .A2(_08695_),
    .A1(_08692_));
 sg13g2_nor2_1 _17182_ (.A(_08715_),
    .B(_08716_),
    .Y(_08717_));
 sg13g2_xor2_1 _17183_ (.B(_08716_),
    .A(_08715_),
    .X(_08718_));
 sg13g2_xnor2_1 _17184_ (.Y(_08719_),
    .A(_08707_),
    .B(_08718_));
 sg13g2_nor2b_1 _17185_ (.A(net5558),
    .B_N(net5878),
    .Y(_08720_));
 sg13g2_o21ai_1 _17186_ (.B1(_08720_),
    .Y(_08721_),
    .A1(net5559),
    .A2(_08653_));
 sg13g2_nand2_1 _17187_ (.Y(_08722_),
    .A(_00235_),
    .B(_08721_));
 sg13g2_nand2_1 _17188_ (.Y(_08723_),
    .A(\TRNG.hash[252] ),
    .B(_08722_));
 sg13g2_xnor2_1 _17189_ (.Y(_08724_),
    .A(net5877),
    .B(_08722_));
 sg13g2_o21ai_1 _17190_ (.B1(net4973),
    .Y(_08725_),
    .A1(net3440),
    .A2(net5174));
 sg13g2_a221oi_1 _17191_ (.B2(net5184),
    .C1(_08725_),
    .B1(_08724_),
    .A1(net5837),
    .Y(_00591_),
    .A2(_08719_));
 sg13g2_xnor2_1 _17192_ (.Y(_08726_),
    .A(net5882),
    .B(\TRNG.hash[235] ));
 sg13g2_xnor2_1 _17193_ (.Y(_08727_),
    .A(net5570),
    .B(_08726_));
 sg13g2_xnor2_1 _17194_ (.Y(_08728_),
    .A(_08097_),
    .B(_08727_));
 sg13g2_a21oi_1 _17195_ (.A1(\TRNG.hash[222] ),
    .A2(\TRNG.hash[190] ),
    .Y(_08729_),
    .B1(net5556));
 sg13g2_a21oi_1 _17196_ (.A1(_04285_),
    .A2(_04288_),
    .Y(_08730_),
    .B1(_08729_));
 sg13g2_nor2b_1 _17197_ (.A(_08728_),
    .B_N(_08730_),
    .Y(_08731_));
 sg13g2_xor2_1 _17198_ (.B(_08730_),
    .A(_08728_),
    .X(_08732_));
 sg13g2_xnor2_1 _17199_ (.Y(_08733_),
    .A(\TRNG.hash[234] ),
    .B(\TRNG.hash[255] ));
 sg13g2_xnor2_1 _17200_ (.Y(_08734_),
    .A(net5560),
    .B(_08733_));
 sg13g2_nor2b_1 _17201_ (.A(_08069_),
    .B_N(_08734_),
    .Y(_08735_));
 sg13g2_xnor2_1 _17202_ (.Y(_08736_),
    .A(_08069_),
    .B(_08734_));
 sg13g2_nor2_1 _17203_ (.A(\TRNG.hash[221] ),
    .B(\TRNG.hash[253] ),
    .Y(_08737_));
 sg13g2_a21oi_1 _17204_ (.A1(\TRNG.hash[221] ),
    .A2(net5557),
    .Y(_08738_),
    .B1(\TRNG.hash[189] ));
 sg13g2_nor2_1 _17205_ (.A(_08737_),
    .B(_08738_),
    .Y(_08739_));
 sg13g2_a21oi_2 _17206_ (.B1(_08735_),
    .Y(_08740_),
    .A2(_08739_),
    .A1(_08736_));
 sg13g2_nor2_1 _17207_ (.A(_08732_),
    .B(_08740_),
    .Y(_08741_));
 sg13g2_nor2_1 _17208_ (.A(_08710_),
    .B(_08714_),
    .Y(_08742_));
 sg13g2_xnor2_1 _17209_ (.Y(_08743_),
    .A(_08736_),
    .B(_08739_));
 sg13g2_nor2_1 _17210_ (.A(_08742_),
    .B(_08743_),
    .Y(_08744_));
 sg13g2_nand2_1 _17211_ (.Y(_08745_),
    .A(_08742_),
    .B(_08743_));
 sg13g2_xor2_1 _17212_ (.B(_08743_),
    .A(_08742_),
    .X(_08746_));
 sg13g2_nand2_1 _17213_ (.Y(_08747_),
    .A(_08718_),
    .B(_08746_));
 sg13g2_a21oi_1 _17214_ (.A1(_08717_),
    .A2(_08745_),
    .Y(_08748_),
    .B1(_08744_));
 sg13g2_o21ai_1 _17215_ (.B1(_08748_),
    .Y(_08749_),
    .A1(_08706_),
    .A2(_08747_));
 sg13g2_nand2_1 _17216_ (.Y(_08750_),
    .A(_08732_),
    .B(_08740_));
 sg13g2_xnor2_1 _17217_ (.Y(_08751_),
    .A(_08732_),
    .B(_08740_));
 sg13g2_a21oi_1 _17218_ (.A1(_08749_),
    .A2(_08750_),
    .Y(_08752_),
    .B1(_08741_));
 sg13g2_a21oi_1 _17219_ (.A1(_08097_),
    .A2(_08727_),
    .Y(_08753_),
    .B1(_08731_));
 sg13g2_xor2_1 _17220_ (.B(net5885),
    .A(net5881),
    .X(_08754_));
 sg13g2_xnor2_1 _17221_ (.Y(_08755_),
    .A(\TRNG.hash[225] ),
    .B(_08754_));
 sg13g2_a21o_1 _17222_ (.A2(\TRNG.hash[191] ),
    .A1(\TRNG.hash[223] ),
    .B1(\TRNG.hash[255] ),
    .X(_08756_));
 sg13g2_o21ai_1 _17223_ (.B1(_08756_),
    .Y(_08757_),
    .A1(\TRNG.hash[223] ),
    .A2(\TRNG.hash[191] ));
 sg13g2_xnor2_1 _17224_ (.Y(_08758_),
    .A(_08755_),
    .B(_08757_));
 sg13g2_xnor2_1 _17225_ (.Y(_08759_),
    .A(_08116_),
    .B(_08758_));
 sg13g2_xnor2_1 _17226_ (.Y(_08760_),
    .A(_08753_),
    .B(_08759_));
 sg13g2_or2_1 _17227_ (.X(_08761_),
    .B(_08760_),
    .A(_08752_));
 sg13g2_a21oi_1 _17228_ (.A1(_08752_),
    .A2(_08760_),
    .Y(_08762_),
    .B1(net5487));
 sg13g2_o21ai_1 _17229_ (.B1(net3788),
    .Y(_08763_),
    .A1(net5557),
    .A2(_08723_));
 sg13g2_nor2_1 _17230_ (.A(net5556),
    .B(_08763_),
    .Y(_08764_));
 sg13g2_xor2_1 _17231_ (.B(_08764_),
    .A(\TRNG.hash[255] ),
    .X(_08765_));
 sg13g2_o21ai_1 _17232_ (.B1(net4973),
    .Y(_08766_),
    .A1(\TRNG.hash[255] ),
    .A2(net5174));
 sg13g2_a221oi_1 _17233_ (.B2(net5185),
    .C1(_08766_),
    .B1(_08765_),
    .A1(_08761_),
    .Y(_00592_),
    .A2(_08762_));
 sg13g2_nor2_2 _17234_ (.A(net5360),
    .B(_06910_),
    .Y(_08767_));
 sg13g2_mux2_1 _17235_ (.A0(net2550),
    .A1(net5689),
    .S(net5060),
    .X(_00593_));
 sg13g2_mux2_1 _17236_ (.A0(net3186),
    .A1(net5688),
    .S(net5060),
    .X(_00594_));
 sg13g2_mux2_1 _17237_ (.A0(net2571),
    .A1(net5684),
    .S(net5061),
    .X(_00595_));
 sg13g2_nor2_1 _17238_ (.A(net2682),
    .B(net5062),
    .Y(_08768_));
 sg13g2_a21oi_1 _17239_ (.A1(net5495),
    .A2(net5062),
    .Y(_00596_),
    .B1(_08768_));
 sg13g2_mux2_1 _17240_ (.A0(net2475),
    .A1(net5682),
    .S(net5061),
    .X(_00597_));
 sg13g2_mux2_1 _17241_ (.A0(net3218),
    .A1(net5681),
    .S(net5061),
    .X(_00598_));
 sg13g2_mux2_1 _17242_ (.A0(net3194),
    .A1(net5677),
    .S(net5061),
    .X(_00599_));
 sg13g2_mux2_1 _17243_ (.A0(net3019),
    .A1(\TRNG.sha256.expand.data1_to_ram[7] ),
    .S(net5063),
    .X(_00600_));
 sg13g2_mux2_1 _17244_ (.A0(net3188),
    .A1(net5671),
    .S(net5061),
    .X(_00601_));
 sg13g2_mux2_1 _17245_ (.A0(net3104),
    .A1(net5669),
    .S(net5063),
    .X(_00602_));
 sg13g2_mux2_1 _17246_ (.A0(net2745),
    .A1(net5667),
    .S(net5063),
    .X(_00603_));
 sg13g2_mux2_1 _17247_ (.A0(net2940),
    .A1(net5666),
    .S(net5060),
    .X(_00604_));
 sg13g2_mux2_1 _17248_ (.A0(net3117),
    .A1(net5663),
    .S(net5060),
    .X(_00605_));
 sg13g2_mux2_1 _17249_ (.A0(net3195),
    .A1(net5661),
    .S(net5060),
    .X(_00606_));
 sg13g2_mux2_1 _17250_ (.A0(net2527),
    .A1(net5658),
    .S(net5063),
    .X(_00607_));
 sg13g2_mux2_1 _17251_ (.A0(net2811),
    .A1(net5656),
    .S(net5060),
    .X(_00608_));
 sg13g2_mux2_1 _17252_ (.A0(net2646),
    .A1(net5653),
    .S(net5063),
    .X(_00609_));
 sg13g2_mux2_1 _17253_ (.A0(net3021),
    .A1(net5652),
    .S(net5062),
    .X(_00610_));
 sg13g2_mux2_1 _17254_ (.A0(net3110),
    .A1(net5649),
    .S(net5060),
    .X(_00611_));
 sg13g2_mux2_1 _17255_ (.A0(net2963),
    .A1(net5647),
    .S(net5061),
    .X(_00612_));
 sg13g2_mux2_1 _17256_ (.A0(net2620),
    .A1(net5644),
    .S(net5062),
    .X(_00613_));
 sg13g2_mux2_1 _17257_ (.A0(net2826),
    .A1(net5641),
    .S(net5062),
    .X(_00614_));
 sg13g2_mux2_1 _17258_ (.A0(net2552),
    .A1(net5637),
    .S(net5062),
    .X(_00615_));
 sg13g2_mux2_1 _17259_ (.A0(net3307),
    .A1(\TRNG.sha256.expand.data1_to_ram[23] ),
    .S(net5064),
    .X(_00616_));
 sg13g2_mux2_1 _17260_ (.A0(net2928),
    .A1(net5634),
    .S(net5062),
    .X(_00617_));
 sg13g2_mux2_1 _17261_ (.A0(net3026),
    .A1(net5632),
    .S(net5062),
    .X(_00618_));
 sg13g2_mux2_1 _17262_ (.A0(net2794),
    .A1(net5630),
    .S(net5064),
    .X(_00619_));
 sg13g2_mux2_1 _17263_ (.A0(net3277),
    .A1(net5628),
    .S(net5060),
    .X(_00620_));
 sg13g2_mux2_1 _17264_ (.A0(net2609),
    .A1(net5625),
    .S(net5063),
    .X(_00621_));
 sg13g2_mux2_1 _17265_ (.A0(net3037),
    .A1(net5621),
    .S(net5063),
    .X(_00622_));
 sg13g2_mux2_1 _17266_ (.A0(net3358),
    .A1(net5619),
    .S(net5061),
    .X(_00623_));
 sg13g2_mux2_1 _17267_ (.A0(net3102),
    .A1(\TRNG.sha256.expand.data1_to_ram[31] ),
    .S(net5063),
    .X(_00624_));
 sg13g2_nor2_1 _17268_ (.A(net5213),
    .B(_06913_),
    .Y(_08769_));
 sg13g2_mux2_1 _17269_ (.A0(net3153),
    .A1(net5690),
    .S(net5056),
    .X(_00625_));
 sg13g2_mux2_1 _17270_ (.A0(net2855),
    .A1(net5687),
    .S(net5056),
    .X(_00626_));
 sg13g2_mux2_1 _17271_ (.A0(net3114),
    .A1(net5685),
    .S(net5057),
    .X(_00627_));
 sg13g2_nor2_1 _17272_ (.A(net3299),
    .B(net5059),
    .Y(_08770_));
 sg13g2_a21oi_1 _17273_ (.A1(net5494),
    .A2(net5059),
    .Y(_00628_),
    .B1(_08770_));
 sg13g2_mux2_1 _17274_ (.A0(net2882),
    .A1(\TRNG.sha256.expand.data1_to_ram[4] ),
    .S(net5057),
    .X(_00629_));
 sg13g2_mux2_1 _17275_ (.A0(net2649),
    .A1(net5679),
    .S(net5057),
    .X(_00630_));
 sg13g2_mux2_1 _17276_ (.A0(net3082),
    .A1(net5677),
    .S(net5057),
    .X(_00631_));
 sg13g2_mux2_1 _17277_ (.A0(net3302),
    .A1(net5674),
    .S(net5057),
    .X(_00632_));
 sg13g2_mux2_1 _17278_ (.A0(net3178),
    .A1(net5672),
    .S(net5057),
    .X(_00633_));
 sg13g2_mux2_1 _17279_ (.A0(net2740),
    .A1(net5670),
    .S(net5058),
    .X(_00634_));
 sg13g2_mux2_1 _17280_ (.A0(net2719),
    .A1(net5668),
    .S(net5058),
    .X(_00635_));
 sg13g2_mux2_1 _17281_ (.A0(net3167),
    .A1(net5665),
    .S(net5056),
    .X(_00636_));
 sg13g2_mux2_1 _17282_ (.A0(net3115),
    .A1(net5662),
    .S(net5056),
    .X(_00637_));
 sg13g2_mux2_1 _17283_ (.A0(net3088),
    .A1(net5660),
    .S(net5056),
    .X(_00638_));
 sg13g2_mux2_1 _17284_ (.A0(net2784),
    .A1(net5659),
    .S(net5058),
    .X(_00639_));
 sg13g2_mux2_1 _17285_ (.A0(net3100),
    .A1(net5655),
    .S(net5055),
    .X(_00640_));
 sg13g2_mux2_1 _17286_ (.A0(net3227),
    .A1(net5653),
    .S(net5058),
    .X(_00641_));
 sg13g2_mux2_1 _17287_ (.A0(net2738),
    .A1(net5651),
    .S(net5059),
    .X(_00642_));
 sg13g2_mux2_1 _17288_ (.A0(net2771),
    .A1(net5648),
    .S(net5056),
    .X(_00643_));
 sg13g2_mux2_1 _17289_ (.A0(net3364),
    .A1(net5646),
    .S(net5056),
    .X(_00644_));
 sg13g2_mux2_1 _17290_ (.A0(net2644),
    .A1(net5643),
    .S(net5055),
    .X(_00645_));
 sg13g2_mux2_1 _17291_ (.A0(net3326),
    .A1(net5640),
    .S(net5055),
    .X(_00646_));
 sg13g2_mux2_1 _17292_ (.A0(net2660),
    .A1(net5638),
    .S(net5055),
    .X(_00647_));
 sg13g2_mux2_1 _17293_ (.A0(net2884),
    .A1(net5635),
    .S(net5055),
    .X(_00648_));
 sg13g2_mux2_1 _17294_ (.A0(net3177),
    .A1(net5633),
    .S(net5055),
    .X(_00649_));
 sg13g2_mux2_1 _17295_ (.A0(net3154),
    .A1(net5631),
    .S(net5055),
    .X(_00650_));
 sg13g2_mux2_1 _17296_ (.A0(net2878),
    .A1(net5629),
    .S(net5055),
    .X(_00651_));
 sg13g2_mux2_1 _17297_ (.A0(net3106),
    .A1(net5627),
    .S(net5057),
    .X(_00652_));
 sg13g2_mux2_1 _17298_ (.A0(net2728),
    .A1(net5624),
    .S(net5058),
    .X(_00653_));
 sg13g2_mux2_1 _17299_ (.A0(net2921),
    .A1(net5621),
    .S(net5058),
    .X(_00654_));
 sg13g2_mux2_1 _17300_ (.A0(net3066),
    .A1(net5619),
    .S(net5057),
    .X(_00655_));
 sg13g2_mux2_1 _17301_ (.A0(net2980),
    .A1(net5616),
    .S(net5058),
    .X(_00656_));
 sg13g2_nand4_1 _17302_ (.B(_04277_),
    .C(_04278_),
    .A(\TRNG.sha256.expand.exp_ctrl.write_en1 ),
    .Y(_08771_),
    .D(net5393));
 sg13g2_mux2_1 _17303_ (.A0(net5690),
    .A1(net3320),
    .S(net5169),
    .X(_00657_));
 sg13g2_mux2_1 _17304_ (.A0(net5687),
    .A1(net3124),
    .S(net5169),
    .X(_00658_));
 sg13g2_mux2_1 _17305_ (.A0(net5685),
    .A1(net3325),
    .S(net5170),
    .X(_00659_));
 sg13g2_nand2_1 _17306_ (.Y(_08772_),
    .A(net2301),
    .B(net5171));
 sg13g2_o21ai_1 _17307_ (.B1(_08772_),
    .Y(_00660_),
    .A1(net5496),
    .A2(net5171));
 sg13g2_mux2_1 _17308_ (.A0(net5683),
    .A1(net3369),
    .S(net5170),
    .X(_00661_));
 sg13g2_mux2_1 _17309_ (.A0(net5679),
    .A1(net3293),
    .S(net5170),
    .X(_00662_));
 sg13g2_mux2_1 _17310_ (.A0(net5678),
    .A1(net3348),
    .S(net5170),
    .X(_00663_));
 sg13g2_mux2_1 _17311_ (.A0(net5674),
    .A1(net3351),
    .S(net5172),
    .X(_00664_));
 sg13g2_mux2_1 _17312_ (.A0(net5673),
    .A1(net3197),
    .S(net5170),
    .X(_00665_));
 sg13g2_mux2_1 _17313_ (.A0(net5670),
    .A1(net3366),
    .S(net5173),
    .X(_00666_));
 sg13g2_mux2_1 _17314_ (.A0(net5667),
    .A1(net3272),
    .S(net5173),
    .X(_00667_));
 sg13g2_mux2_1 _17315_ (.A0(net5665),
    .A1(net3357),
    .S(net5169),
    .X(_00668_));
 sg13g2_mux2_1 _17316_ (.A0(net5662),
    .A1(net3330),
    .S(net5169),
    .X(_00669_));
 sg13g2_mux2_1 _17317_ (.A0(net5660),
    .A1(net3327),
    .S(net5169),
    .X(_00670_));
 sg13g2_mux2_1 _17318_ (.A0(net5658),
    .A1(net3360),
    .S(net5172),
    .X(_00671_));
 sg13g2_mux2_1 _17319_ (.A0(net5655),
    .A1(net3305),
    .S(net5169),
    .X(_00672_));
 sg13g2_mux2_1 _17320_ (.A0(net5653),
    .A1(net3403),
    .S(net5172),
    .X(_00673_));
 sg13g2_mux2_1 _17321_ (.A0(net5651),
    .A1(net3287),
    .S(net5171),
    .X(_00674_));
 sg13g2_mux2_1 _17322_ (.A0(net5648),
    .A1(net3321),
    .S(net5169),
    .X(_00675_));
 sg13g2_mux2_1 _17323_ (.A0(net5646),
    .A1(net3294),
    .S(net5169),
    .X(_00676_));
 sg13g2_mux2_1 _17324_ (.A0(net5643),
    .A1(net3301),
    .S(net5171),
    .X(_00677_));
 sg13g2_mux2_1 _17325_ (.A0(net5640),
    .A1(net3429),
    .S(net5171),
    .X(_00678_));
 sg13g2_mux2_1 _17326_ (.A0(net5637),
    .A1(net3210),
    .S(net5171),
    .X(_00679_));
 sg13g2_mux2_1 _17327_ (.A0(net5635),
    .A1(net3237),
    .S(net5172),
    .X(_00680_));
 sg13g2_mux2_1 _17328_ (.A0(net5633),
    .A1(net3312),
    .S(net5172),
    .X(_00681_));
 sg13g2_mux2_1 _17329_ (.A0(net5631),
    .A1(net3385),
    .S(net5171),
    .X(_00682_));
 sg13g2_mux2_1 _17330_ (.A0(net5630),
    .A1(net3304),
    .S(net5171),
    .X(_00683_));
 sg13g2_mux2_1 _17331_ (.A0(net3345),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[0][27] ),
    .S(net5170),
    .X(_00684_));
 sg13g2_mux2_1 _17332_ (.A0(net5625),
    .A1(net3329),
    .S(net5172),
    .X(_00685_));
 sg13g2_mux2_1 _17333_ (.A0(net5623),
    .A1(net3166),
    .S(net5173),
    .X(_00686_));
 sg13g2_mux2_1 _17334_ (.A0(net5620),
    .A1(net3259),
    .S(net5170),
    .X(_00687_));
 sg13g2_mux2_1 _17335_ (.A0(net5616),
    .A1(net3340),
    .S(net5172),
    .X(_00688_));
 sg13g2_nor2_2 _17336_ (.A(net5213),
    .B(_06885_),
    .Y(_08773_));
 sg13g2_mux2_1 _17337_ (.A0(net2988),
    .A1(net5690),
    .S(net5050),
    .X(_00689_));
 sg13g2_mux2_1 _17338_ (.A0(net2986),
    .A1(net5687),
    .S(net5050),
    .X(_00690_));
 sg13g2_nand2_1 _17339_ (.Y(_08774_),
    .A(net5684),
    .B(net5051));
 sg13g2_o21ai_1 _17340_ (.B1(_08774_),
    .Y(_00691_),
    .A1(_04345_),
    .A2(net5051));
 sg13g2_nor2_1 _17341_ (.A(net2692),
    .B(net5049),
    .Y(_08775_));
 sg13g2_a21oi_1 _17342_ (.A1(net5494),
    .A2(net5049),
    .Y(_00692_),
    .B1(_08775_));
 sg13g2_nand2_1 _17343_ (.Y(_08776_),
    .A(net5683),
    .B(net5051));
 sg13g2_o21ai_1 _17344_ (.B1(_08776_),
    .Y(_00693_),
    .A1(_04346_),
    .A2(net5051));
 sg13g2_mux2_1 _17345_ (.A0(net2998),
    .A1(net5680),
    .S(net5054),
    .X(_00694_));
 sg13g2_mux2_1 _17346_ (.A0(net3118),
    .A1(net5677),
    .S(net5051),
    .X(_00695_));
 sg13g2_mux2_1 _17347_ (.A0(net3201),
    .A1(net5674),
    .S(net5053),
    .X(_00696_));
 sg13g2_nand2_1 _17348_ (.Y(_08777_),
    .A(net5672),
    .B(net5054));
 sg13g2_o21ai_1 _17349_ (.B1(_08777_),
    .Y(_00697_),
    .A1(_04350_),
    .A2(net5051));
 sg13g2_mux2_1 _17350_ (.A0(net2828),
    .A1(net5670),
    .S(net5053),
    .X(_00698_));
 sg13g2_nand2_1 _17351_ (.Y(_08778_),
    .A(\TRNG.sha256.expand.data1_to_ram[10] ),
    .B(net5052));
 sg13g2_o21ai_1 _17352_ (.B1(_08778_),
    .Y(_00699_),
    .A1(_04352_),
    .A2(net5052));
 sg13g2_mux2_1 _17353_ (.A0(net3266),
    .A1(net5665),
    .S(net5050),
    .X(_00700_));
 sg13g2_mux2_1 _17354_ (.A0(net3219),
    .A1(net5662),
    .S(net5050),
    .X(_00701_));
 sg13g2_mux2_1 _17355_ (.A0(net3257),
    .A1(net5660),
    .S(net5050),
    .X(_00702_));
 sg13g2_nand2_1 _17356_ (.Y(_08779_),
    .A(net5658),
    .B(net5053));
 sg13g2_o21ai_1 _17357_ (.B1(_08779_),
    .Y(_00703_),
    .A1(_04356_),
    .A2(net5053));
 sg13g2_mux2_1 _17358_ (.A0(net3062),
    .A1(net5655),
    .S(net5048),
    .X(_00704_));
 sg13g2_nand2_1 _17359_ (.Y(_08780_),
    .A(net5654),
    .B(net5052));
 sg13g2_o21ai_1 _17360_ (.B1(_08780_),
    .Y(_00705_),
    .A1(_04358_),
    .A2(net5052));
 sg13g2_mux2_1 _17361_ (.A0(net2966),
    .A1(net5651),
    .S(net5049),
    .X(_00706_));
 sg13g2_mux2_1 _17362_ (.A0(net2983),
    .A1(net5648),
    .S(net5050),
    .X(_00707_));
 sg13g2_mux2_1 _17363_ (.A0(net3297),
    .A1(net5646),
    .S(net5050),
    .X(_00708_));
 sg13g2_nand2_1 _17364_ (.Y(_08781_),
    .A(net5643),
    .B(net5049));
 sg13g2_o21ai_1 _17365_ (.B1(_08781_),
    .Y(_00709_),
    .A1(_04362_),
    .A2(net5049));
 sg13g2_mux2_1 _17366_ (.A0(net3250),
    .A1(net5640),
    .S(net5048),
    .X(_00710_));
 sg13g2_nand2_1 _17367_ (.Y(_08782_),
    .A(net5637),
    .B(net5048));
 sg13g2_o21ai_1 _17368_ (.B1(_08782_),
    .Y(_00711_),
    .A1(_04364_),
    .A2(net5048));
 sg13g2_mux2_1 _17369_ (.A0(net3109),
    .A1(net5635),
    .S(net5048),
    .X(_00712_));
 sg13g2_mux2_1 _17370_ (.A0(net3217),
    .A1(net5633),
    .S(net5048),
    .X(_00713_));
 sg13g2_mux2_1 _17371_ (.A0(net3152),
    .A1(net5631),
    .S(net5048),
    .X(_00714_));
 sg13g2_nand2_1 _17372_ (.Y(_08783_),
    .A(net5629),
    .B(net5048));
 sg13g2_o21ai_1 _17373_ (.B1(_08783_),
    .Y(_00715_),
    .A1(_04368_),
    .A2(net5049));
 sg13g2_mux2_1 _17374_ (.A0(net3058),
    .A1(net5627),
    .S(net5051),
    .X(_00716_));
 sg13g2_nand2_1 _17375_ (.Y(_08784_),
    .A(net5624),
    .B(net5052));
 sg13g2_o21ai_1 _17376_ (.B1(_08784_),
    .Y(_00717_),
    .A1(_04370_),
    .A2(net5052));
 sg13g2_mux2_1 _17377_ (.A0(net2935),
    .A1(net5622),
    .S(net5052),
    .X(_00718_));
 sg13g2_mux2_1 _17378_ (.A0(net3049),
    .A1(net5619),
    .S(net5051),
    .X(_00719_));
 sg13g2_mux2_1 _17379_ (.A0(net3000),
    .A1(net5616),
    .S(net5052),
    .X(_00720_));
 sg13g2_nand4_1 _17380_ (.B(\TRNG.sha256.expand.address1[3] ),
    .C(_04278_),
    .A(\TRNG.sha256.expand.exp_ctrl.write_en1 ),
    .Y(_08785_),
    .D(net5393));
 sg13g2_mux2_1 _17381_ (.A0(net3063),
    .A1(\TRNG.sha256.expand.msg_schdl.RAM[8][0] ),
    .S(net5164),
    .X(_00721_));
 sg13g2_mux2_1 _17382_ (.A0(net5688),
    .A1(net3339),
    .S(net5164),
    .X(_00722_));
 sg13g2_mux2_1 _17383_ (.A0(net5686),
    .A1(net3316),
    .S(net5165),
    .X(_00723_));
 sg13g2_nand2_1 _17384_ (.Y(_08786_),
    .A(net2674),
    .B(net5166));
 sg13g2_o21ai_1 _17385_ (.B1(_08786_),
    .Y(_00724_),
    .A1(net5495),
    .A2(net5166));
 sg13g2_mux2_1 _17386_ (.A0(net5682),
    .A1(net3352),
    .S(net5165),
    .X(_00725_));
 sg13g2_mux2_1 _17387_ (.A0(net5679),
    .A1(net3331),
    .S(net5165),
    .X(_00726_));
 sg13g2_mux2_1 _17388_ (.A0(net5676),
    .A1(net3353),
    .S(net5165),
    .X(_00727_));
 sg13g2_mux2_1 _17389_ (.A0(net5675),
    .A1(net3251),
    .S(net5167),
    .X(_00728_));
 sg13g2_mux2_1 _17390_ (.A0(net5671),
    .A1(net3361),
    .S(net5167),
    .X(_00729_));
 sg13g2_mux2_1 _17391_ (.A0(net5669),
    .A1(net3350),
    .S(net5167),
    .X(_00730_));
 sg13g2_mux2_1 _17392_ (.A0(net5668),
    .A1(net3231),
    .S(net5168),
    .X(_00731_));
 sg13g2_mux2_1 _17393_ (.A0(net5666),
    .A1(net3274),
    .S(net5164),
    .X(_00732_));
 sg13g2_mux2_1 _17394_ (.A0(net5664),
    .A1(net3333),
    .S(net5164),
    .X(_00733_));
 sg13g2_mux2_1 _17395_ (.A0(net5661),
    .A1(net3323),
    .S(net5164),
    .X(_00734_));
 sg13g2_mux2_1 _17396_ (.A0(net5659),
    .A1(net3235),
    .S(net5167),
    .X(_00735_));
 sg13g2_mux2_1 _17397_ (.A0(net5657),
    .A1(net3317),
    .S(net5166),
    .X(_00736_));
 sg13g2_mux2_1 _17398_ (.A0(net5654),
    .A1(net3262),
    .S(net5167),
    .X(_00737_));
 sg13g2_mux2_1 _17399_ (.A0(net5652),
    .A1(net3221),
    .S(net5166),
    .X(_00738_));
 sg13g2_mux2_1 _17400_ (.A0(net5650),
    .A1(net3228),
    .S(net5164),
    .X(_00739_));
 sg13g2_mux2_1 _17401_ (.A0(net5647),
    .A1(net3239),
    .S(net5164),
    .X(_00740_));
 sg13g2_mux2_1 _17402_ (.A0(net5645),
    .A1(net3268),
    .S(net5166),
    .X(_00741_));
 sg13g2_mux2_1 _17403_ (.A0(net5642),
    .A1(net3275),
    .S(net5166),
    .X(_00742_));
 sg13g2_mux2_1 _17404_ (.A0(net5639),
    .A1(net3242),
    .S(net5166),
    .X(_00743_));
 sg13g2_mux2_1 _17405_ (.A0(net5636),
    .A1(net3258),
    .S(net5168),
    .X(_00744_));
 sg13g2_mux2_1 _17406_ (.A0(net5634),
    .A1(net3341),
    .S(net5168),
    .X(_00745_));
 sg13g2_mux2_1 _17407_ (.A0(net5632),
    .A1(net3190),
    .S(net5166),
    .X(_00746_));
 sg13g2_mux2_1 _17408_ (.A0(net5629),
    .A1(net3289),
    .S(net5168),
    .X(_00747_));
 sg13g2_mux2_1 _17409_ (.A0(net5628),
    .A1(net3342),
    .S(net5165),
    .X(_00748_));
 sg13g2_mux2_1 _17410_ (.A0(net5626),
    .A1(net3362),
    .S(net5167),
    .X(_00749_));
 sg13g2_mux2_1 _17411_ (.A0(net5623),
    .A1(net3284),
    .S(net5167),
    .X(_00750_));
 sg13g2_mux2_1 _17412_ (.A0(net5618),
    .A1(net3367),
    .S(net5164),
    .X(_00751_));
 sg13g2_mux2_1 _17413_ (.A0(net5617),
    .A1(net3286),
    .S(net5167),
    .X(_00752_));
 sg13g2_nor2_1 _17414_ (.A(net5213),
    .B(_06910_),
    .Y(_08787_));
 sg13g2_mux2_1 _17415_ (.A0(net2697),
    .A1(net5690),
    .S(net5044),
    .X(_00753_));
 sg13g2_mux2_1 _17416_ (.A0(net2736),
    .A1(net5687),
    .S(net5044),
    .X(_00754_));
 sg13g2_mux2_1 _17417_ (.A0(net3248),
    .A1(net5685),
    .S(net5045),
    .X(_00755_));
 sg13g2_nor2_1 _17418_ (.A(net2676),
    .B(net5047),
    .Y(_08788_));
 sg13g2_a21oi_1 _17419_ (.A1(net5494),
    .A2(net5047),
    .Y(_00756_),
    .B1(_08788_));
 sg13g2_mux2_1 _17420_ (.A0(net2970),
    .A1(net5683),
    .S(net5045),
    .X(_00757_));
 sg13g2_mux2_1 _17421_ (.A0(net2471),
    .A1(net5680),
    .S(net5045),
    .X(_00758_));
 sg13g2_mux2_1 _17422_ (.A0(net2567),
    .A1(net5677),
    .S(net5045),
    .X(_00759_));
 sg13g2_mux2_1 _17423_ (.A0(net2925),
    .A1(net5674),
    .S(net5045),
    .X(_00760_));
 sg13g2_mux2_1 _17424_ (.A0(net2968),
    .A1(net5672),
    .S(net5045),
    .X(_00761_));
 sg13g2_mux2_1 _17425_ (.A0(net2517),
    .A1(net5670),
    .S(net5046),
    .X(_00762_));
 sg13g2_mux2_1 _17426_ (.A0(net3253),
    .A1(net5668),
    .S(net5046),
    .X(_00763_));
 sg13g2_mux2_1 _17427_ (.A0(net2559),
    .A1(net5665),
    .S(net5044),
    .X(_00764_));
 sg13g2_mux2_1 _17428_ (.A0(net2704),
    .A1(net5662),
    .S(net5044),
    .X(_00765_));
 sg13g2_mux2_1 _17429_ (.A0(net2553),
    .A1(net5660),
    .S(net5044),
    .X(_00766_));
 sg13g2_mux2_1 _17430_ (.A0(net2867),
    .A1(net5659),
    .S(net5046),
    .X(_00767_));
 sg13g2_mux2_1 _17431_ (.A0(net3076),
    .A1(net5655),
    .S(net5043),
    .X(_00768_));
 sg13g2_mux2_1 _17432_ (.A0(net3173),
    .A1(\TRNG.sha256.expand.data1_to_ram[16] ),
    .S(net5046),
    .X(_00769_));
 sg13g2_mux2_1 _17433_ (.A0(net2498),
    .A1(net5651),
    .S(net5047),
    .X(_00770_));
 sg13g2_mux2_1 _17434_ (.A0(net2604),
    .A1(net5648),
    .S(net5044),
    .X(_00771_));
 sg13g2_mux2_1 _17435_ (.A0(net2647),
    .A1(net5646),
    .S(net5044),
    .X(_00772_));
 sg13g2_mux2_1 _17436_ (.A0(net2744),
    .A1(net5643),
    .S(net5043),
    .X(_00773_));
 sg13g2_mux2_1 _17437_ (.A0(net3241),
    .A1(net5641),
    .S(net5043),
    .X(_00774_));
 sg13g2_mux2_1 _17438_ (.A0(net2915),
    .A1(net5638),
    .S(net5043),
    .X(_00775_));
 sg13g2_mux2_1 _17439_ (.A0(net2695),
    .A1(net5635),
    .S(net5043),
    .X(_00776_));
 sg13g2_mux2_1 _17440_ (.A0(net2877),
    .A1(net5633),
    .S(net5043),
    .X(_00777_));
 sg13g2_mux2_1 _17441_ (.A0(net3126),
    .A1(net5631),
    .S(net5043),
    .X(_00778_));
 sg13g2_mux2_1 _17442_ (.A0(net2827),
    .A1(net5629),
    .S(net5043),
    .X(_00779_));
 sg13g2_mux2_1 _17443_ (.A0(net2628),
    .A1(net5627),
    .S(net5045),
    .X(_00780_));
 sg13g2_mux2_1 _17444_ (.A0(net3045),
    .A1(net5624),
    .S(net5046),
    .X(_00781_));
 sg13g2_mux2_1 _17445_ (.A0(net2577),
    .A1(net5622),
    .S(net5046),
    .X(_00782_));
 sg13g2_mux2_1 _17446_ (.A0(net2518),
    .A1(net5618),
    .S(net5045),
    .X(_00783_));
 sg13g2_mux2_1 _17447_ (.A0(net2714),
    .A1(net5616),
    .S(net5046),
    .X(_00784_));
 sg13g2_nor2_2 _17448_ (.A(net5207),
    .B(_06910_),
    .Y(_08789_));
 sg13g2_mux2_1 _17449_ (.A0(net3081),
    .A1(net5689),
    .S(net5038),
    .X(_00785_));
 sg13g2_mux2_1 _17450_ (.A0(net3029),
    .A1(net5688),
    .S(net5038),
    .X(_00786_));
 sg13g2_mux2_1 _17451_ (.A0(net2523),
    .A1(net5686),
    .S(net5039),
    .X(_00787_));
 sg13g2_nor2_1 _17452_ (.A(net2753),
    .B(net5040),
    .Y(_08790_));
 sg13g2_a21oi_1 _17453_ (.A1(net5494),
    .A2(net5040),
    .Y(_00788_),
    .B1(_08790_));
 sg13g2_mux2_1 _17454_ (.A0(net2847),
    .A1(net5682),
    .S(net5039),
    .X(_00789_));
 sg13g2_mux2_1 _17455_ (.A0(net2954),
    .A1(net5679),
    .S(net5039),
    .X(_00790_));
 sg13g2_mux2_1 _17456_ (.A0(net2751),
    .A1(net5676),
    .S(net5039),
    .X(_00791_));
 sg13g2_mux2_1 _17457_ (.A0(net2992),
    .A1(net5675),
    .S(net5041),
    .X(_00792_));
 sg13g2_mux2_1 _17458_ (.A0(net3245),
    .A1(net5671),
    .S(net5041),
    .X(_00793_));
 sg13g2_mux2_1 _17459_ (.A0(net2866),
    .A1(net5669),
    .S(net5041),
    .X(_00794_));
 sg13g2_mux2_1 _17460_ (.A0(net2822),
    .A1(net5668),
    .S(net5042),
    .X(_00795_));
 sg13g2_mux2_1 _17461_ (.A0(net2941),
    .A1(net5666),
    .S(net5038),
    .X(_00796_));
 sg13g2_mux2_1 _17462_ (.A0(net3035),
    .A1(net5664),
    .S(net5038),
    .X(_00797_));
 sg13g2_mux2_1 _17463_ (.A0(net3089),
    .A1(net5661),
    .S(net5038),
    .X(_00798_));
 sg13g2_mux2_1 _17464_ (.A0(net2964),
    .A1(net5659),
    .S(net5041),
    .X(_00799_));
 sg13g2_mux2_1 _17465_ (.A0(net3215),
    .A1(net5657),
    .S(net5040),
    .X(_00800_));
 sg13g2_mux2_1 _17466_ (.A0(net2835),
    .A1(net5654),
    .S(net5041),
    .X(_00801_));
 sg13g2_mux2_1 _17467_ (.A0(net3065),
    .A1(net5652),
    .S(net5040),
    .X(_00802_));
 sg13g2_mux2_1 _17468_ (.A0(net2802),
    .A1(net5650),
    .S(net5038),
    .X(_00803_));
 sg13g2_mux2_1 _17469_ (.A0(net2995),
    .A1(net5647),
    .S(net5038),
    .X(_00804_));
 sg13g2_mux2_1 _17470_ (.A0(net2959),
    .A1(net5643),
    .S(net5040),
    .X(_00805_));
 sg13g2_mux2_1 _17471_ (.A0(net2993),
    .A1(net5642),
    .S(net5040),
    .X(_00806_));
 sg13g2_mux2_1 _17472_ (.A0(net2767),
    .A1(net5638),
    .S(net5040),
    .X(_00807_));
 sg13g2_mux2_1 _17473_ (.A0(net2729),
    .A1(net5636),
    .S(net5042),
    .X(_00808_));
 sg13g2_mux2_1 _17474_ (.A0(net3083),
    .A1(net5634),
    .S(net5042),
    .X(_00809_));
 sg13g2_mux2_1 _17475_ (.A0(net3145),
    .A1(net5632),
    .S(net5040),
    .X(_00810_));
 sg13g2_mux2_1 _17476_ (.A0(net3057),
    .A1(net5629),
    .S(net5042),
    .X(_00811_));
 sg13g2_mux2_1 _17477_ (.A0(net2746),
    .A1(net5628),
    .S(net5039),
    .X(_00812_));
 sg13g2_mux2_1 _17478_ (.A0(net3059),
    .A1(net5626),
    .S(net5041),
    .X(_00813_));
 sg13g2_mux2_1 _17479_ (.A0(net2678),
    .A1(net5623),
    .S(net5041),
    .X(_00814_));
 sg13g2_mux2_1 _17480_ (.A0(net2839),
    .A1(net5618),
    .S(net5038),
    .X(_00815_));
 sg13g2_mux2_1 _17481_ (.A0(net3163),
    .A1(net5617),
    .S(net5041),
    .X(_00816_));
 sg13g2_nor3_2 _17482_ (.A(_05952_),
    .B(_06001_),
    .C(net5358),
    .Y(_08791_));
 sg13g2_nor2b_2 _17483_ (.A(\TRNG.sha256.control.iteration[6] ),
    .B_N(_08791_),
    .Y(_08792_));
 sg13g2_nand3_1 _17484_ (.B(net3336),
    .C(_08792_),
    .A(\TRNG.sha256.control.iteration[7] ),
    .Y(_08793_));
 sg13g2_nand3_1 _17485_ (.B(\TRNG.sha256.control.iteration[6] ),
    .C(_08791_),
    .A(net5575),
    .Y(_08794_));
 sg13g2_nand4_1 _17486_ (.B(\TRNG.sha256.control.iteration[6] ),
    .C(_00117_),
    .A(net5575),
    .Y(_08795_),
    .D(_08791_));
 sg13g2_nor2b_1 _17487_ (.A(net5575),
    .B_N(\TRNG.sha256.control.iteration[8] ),
    .Y(_08796_));
 sg13g2_nand3_1 _17488_ (.B(_08791_),
    .C(_08796_),
    .A(\TRNG.sha256.control.iteration[6] ),
    .Y(_08797_));
 sg13g2_nand2_1 _17489_ (.Y(_08798_),
    .A(_08795_),
    .B(_08797_));
 sg13g2_nand2_1 _17490_ (.Y(_08799_),
    .A(_08792_),
    .B(_08796_));
 sg13g2_nand2_1 _17491_ (.Y(_08800_),
    .A(_00117_),
    .B(_08792_));
 sg13g2_nand3_1 _17492_ (.B(_00117_),
    .C(_08792_),
    .A(net5575),
    .Y(_08801_));
 sg13g2_and2_2 _17493_ (.A(_08799_),
    .B(_08801_),
    .X(_08802_));
 sg13g2_nand2_2 _17494_ (.Y(_08803_),
    .A(\TRNG.sha256.compress.count[0] ),
    .B(net3817));
 sg13g2_nand3_1 _17495_ (.B(net3817),
    .C(net5874),
    .A(\TRNG.sha256.compress.count[0] ),
    .Y(_08804_));
 sg13g2_nor2b_2 _17496_ (.A(net5876),
    .B_N(net5873),
    .Y(_08805_));
 sg13g2_nand2_2 _17497_ (.Y(_08806_),
    .A(net5873),
    .B(net5874));
 sg13g2_nor2b_1 _17498_ (.A(net5876),
    .B_N(\TRNG.sha256.compress.count[1] ),
    .Y(_08807_));
 sg13g2_nand2_2 _17499_ (.Y(_08808_),
    .A(\TRNG.sha256.compress.count[0] ),
    .B(_08807_));
 sg13g2_nor2_2 _17500_ (.A(_08806_),
    .B(_08808_),
    .Y(_08809_));
 sg13g2_nand2b_2 _17501_ (.Y(_08810_),
    .B(_08805_),
    .A_N(_08804_));
 sg13g2_nand2_2 _17502_ (.Y(_08811_),
    .A(net5876),
    .B(_06867_));
 sg13g2_o21ai_1 _17503_ (.B1(_08810_),
    .Y(_08812_),
    .A1(_06869_),
    .A2(_08811_));
 sg13g2_nand2b_2 _17504_ (.Y(_08813_),
    .B(net5874),
    .A_N(net5873));
 sg13g2_nand3b_1 _17505_ (.B(\TRNG.sha256.compress.count[2] ),
    .C(net5876),
    .Y(_08814_),
    .A_N(net5873));
 sg13g2_nand2b_1 _17506_ (.Y(_08815_),
    .B(_06871_),
    .A_N(_00118_));
 sg13g2_o21ai_1 _17507_ (.B1(_08815_),
    .Y(_08816_),
    .A1(_06870_),
    .A2(net5344));
 sg13g2_o21ai_1 _17508_ (.B1(_08802_),
    .Y(_08817_),
    .A1(_08812_),
    .A2(_08816_));
 sg13g2_nor2_1 _17509_ (.A(_08798_),
    .B(_08817_),
    .Y(_08818_));
 sg13g2_nand2_1 _17510_ (.Y(_08819_),
    .A(_08793_),
    .B(_08818_));
 sg13g2_o21ai_1 _17511_ (.B1(_08819_),
    .Y(_08820_),
    .A1(_00117_),
    .A2(_08793_));
 sg13g2_nor2b_1 _17512_ (.A(_00133_),
    .B_N(_08791_),
    .Y(_08821_));
 sg13g2_xor2_1 _17513_ (.B(_08791_),
    .A(_00133_),
    .X(_08822_));
 sg13g2_o21ai_1 _17514_ (.B1(_08802_),
    .Y(_08823_),
    .A1(_08798_),
    .A2(_08822_));
 sg13g2_nor2_1 _17515_ (.A(_08820_),
    .B(_08823_),
    .Y(_08824_));
 sg13g2_o21ai_1 _17516_ (.B1(net5473),
    .Y(_08825_),
    .A1(net5575),
    .A2(_08800_));
 sg13g2_nor2b_1 _17517_ (.A(net3451),
    .B_N(_08820_),
    .Y(_08826_));
 sg13g2_nor3_1 _17518_ (.A(_08824_),
    .B(_08825_),
    .C(_08826_),
    .Y(_00817_));
 sg13g2_nor2b_1 _17519_ (.A(_00117_),
    .B_N(_08794_),
    .Y(_08827_));
 sg13g2_nor3_1 _17520_ (.A(_08798_),
    .B(_08820_),
    .C(_08827_),
    .Y(_08828_));
 sg13g2_nor2_1 _17521_ (.A(net3336),
    .B(_08819_),
    .Y(_08829_));
 sg13g2_nor3_1 _17522_ (.A(_08825_),
    .B(_08828_),
    .C(net3337),
    .Y(_00818_));
 sg13g2_nor2_2 _17523_ (.A(net5207),
    .B(_06885_),
    .Y(_08830_));
 sg13g2_mux2_1 _17524_ (.A0(net2885),
    .A1(net5689),
    .S(net5033),
    .X(_00819_));
 sg13g2_mux2_1 _17525_ (.A0(net2765),
    .A1(net5688),
    .S(net5033),
    .X(_00820_));
 sg13g2_mux2_1 _17526_ (.A0(net3207),
    .A1(net5686),
    .S(net5034),
    .X(_00821_));
 sg13g2_nor2_1 _17527_ (.A(net2974),
    .B(net5035),
    .Y(_08831_));
 sg13g2_a21oi_1 _17528_ (.A1(net5494),
    .A2(net5035),
    .Y(_00822_),
    .B1(_08831_));
 sg13g2_mux2_1 _17529_ (.A0(net2863),
    .A1(net5682),
    .S(net5034),
    .X(_00823_));
 sg13g2_mux2_1 _17530_ (.A0(net3155),
    .A1(net5679),
    .S(net5034),
    .X(_00824_));
 sg13g2_mux2_1 _17531_ (.A0(net2990),
    .A1(net5676),
    .S(net5034),
    .X(_00825_));
 sg13g2_mux2_1 _17532_ (.A0(net3031),
    .A1(net5675),
    .S(net5036),
    .X(_00826_));
 sg13g2_mux2_1 _17533_ (.A0(net3097),
    .A1(net5671),
    .S(net5036),
    .X(_00827_));
 sg13g2_mux2_1 _17534_ (.A0(net2933),
    .A1(net5669),
    .S(net5036),
    .X(_00828_));
 sg13g2_mux2_1 _17535_ (.A0(net2901),
    .A1(net5668),
    .S(net5037),
    .X(_00829_));
 sg13g2_mux2_1 _17536_ (.A0(net2845),
    .A1(net5666),
    .S(net5033),
    .X(_00830_));
 sg13g2_mux2_1 _17537_ (.A0(net3017),
    .A1(net5664),
    .S(net5033),
    .X(_00831_));
 sg13g2_mux2_1 _17538_ (.A0(net2824),
    .A1(net5661),
    .S(net5033),
    .X(_00832_));
 sg13g2_mux2_1 _17539_ (.A0(net3077),
    .A1(net5659),
    .S(net5036),
    .X(_00833_));
 sg13g2_mux2_1 _17540_ (.A0(net2761),
    .A1(net5657),
    .S(net5035),
    .X(_00834_));
 sg13g2_mux2_1 _17541_ (.A0(net2961),
    .A1(net5654),
    .S(net5036),
    .X(_00835_));
 sg13g2_mux2_1 _17542_ (.A0(net2799),
    .A1(net5652),
    .S(net5035),
    .X(_00836_));
 sg13g2_mux2_1 _17543_ (.A0(net3015),
    .A1(net5649),
    .S(net5033),
    .X(_00837_));
 sg13g2_mux2_1 _17544_ (.A0(net3131),
    .A1(net5647),
    .S(net5033),
    .X(_00838_));
 sg13g2_mux2_1 _17545_ (.A0(net2768),
    .A1(net5643),
    .S(net5035),
    .X(_00839_));
 sg13g2_mux2_1 _17546_ (.A0(net2889),
    .A1(net5641),
    .S(net5035),
    .X(_00840_));
 sg13g2_mux2_1 _17547_ (.A0(net2861),
    .A1(net5638),
    .S(net5035),
    .X(_00841_));
 sg13g2_mux2_1 _17548_ (.A0(net2732),
    .A1(net5636),
    .S(net5037),
    .X(_00842_));
 sg13g2_mux2_1 _17549_ (.A0(net2703),
    .A1(net5634),
    .S(net5037),
    .X(_00843_));
 sg13g2_mux2_1 _17550_ (.A0(net2812),
    .A1(net5632),
    .S(net5035),
    .X(_00844_));
 sg13g2_mux2_1 _17551_ (.A0(net2846),
    .A1(net5629),
    .S(net5037),
    .X(_00845_));
 sg13g2_mux2_1 _17552_ (.A0(net2787),
    .A1(net5627),
    .S(net5034),
    .X(_00846_));
 sg13g2_mux2_1 _17553_ (.A0(net3067),
    .A1(net5625),
    .S(net5036),
    .X(_00847_));
 sg13g2_mux2_1 _17554_ (.A0(net3033),
    .A1(net5621),
    .S(net5036),
    .X(_00848_));
 sg13g2_mux2_1 _17555_ (.A0(net3139),
    .A1(net5618),
    .S(net5033),
    .X(_00849_));
 sg13g2_mux2_1 _17556_ (.A0(net2913),
    .A1(net5617),
    .S(net5036),
    .X(_00850_));
 sg13g2_o21ai_1 _17557_ (.B1(net5875),
    .Y(_08832_),
    .A1(_08803_),
    .A2(_08806_));
 sg13g2_a21oi_1 _17558_ (.A1(_08810_),
    .A2(_08832_),
    .Y(_00851_),
    .B1(net5536));
 sg13g2_nor2_1 _17559_ (.A(\TRNG.sha256.compress.count[1] ),
    .B(net5344),
    .Y(_08833_));
 sg13g2_nand2b_1 _17560_ (.Y(_08834_),
    .B(\TRNG.sha256.compress.count[0] ),
    .A_N(\TRNG.sha256.compress.count[1] ));
 sg13g2_nor2_1 _17561_ (.A(net5344),
    .B(net5342),
    .Y(_08835_));
 sg13g2_nor3_1 _17562_ (.A(net5536),
    .B(_04827_),
    .C(net5156),
    .Y(_00852_));
 sg13g2_nand2_1 _17563_ (.Y(_08836_),
    .A(_06870_),
    .B(_08803_));
 sg13g2_nor3_1 _17564_ (.A(net5536),
    .B(net5156),
    .C(_08836_),
    .Y(_00853_));
 sg13g2_xor2_1 _17565_ (.B(_08803_),
    .A(net5874),
    .X(_08837_));
 sg13g2_nor3_1 _17566_ (.A(net5536),
    .B(net5156),
    .C(_08837_),
    .Y(_00854_));
 sg13g2_xor2_1 _17567_ (.B(_08804_),
    .A(net5873),
    .X(_08838_));
 sg13g2_nor3_1 _17568_ (.A(net5536),
    .B(net5156),
    .C(_08838_),
    .Y(_00855_));
 sg13g2_nand3_1 _17569_ (.B(_04885_),
    .C(_05896_),
    .A(net1142),
    .Y(_08839_));
 sg13g2_o21ai_1 _17570_ (.B1(_08839_),
    .Y(_00856_),
    .A1(_04301_),
    .A2(_04885_));
 sg13g2_and3_1 _17571_ (.X(_08840_),
    .A(\TRNG.uart_tx_inst.ticks_counter[0] ),
    .B(net2385),
    .C(_04885_));
 sg13g2_a21oi_1 _17572_ (.A1(\TRNG.uart_tx_inst.ticks_counter[0] ),
    .A2(_04885_),
    .Y(_08841_),
    .B1(net2385));
 sg13g2_nor2b_1 _17573_ (.A(_05896_),
    .B_N(_04885_),
    .Y(_08842_));
 sg13g2_nand2_1 _17574_ (.Y(_08843_),
    .A(_04885_),
    .B(_05897_));
 sg13g2_nor3_1 _17575_ (.A(_08840_),
    .B(net2386),
    .C(_08842_),
    .Y(_00857_));
 sg13g2_xor2_1 _17576_ (.B(_08840_),
    .A(net3354),
    .X(_00858_));
 sg13g2_nand3_1 _17577_ (.B(net3354),
    .C(_08840_),
    .A(net3696),
    .Y(_08844_));
 sg13g2_a21o_1 _17578_ (.A2(_08840_),
    .A1(net3354),
    .B1(net3696),
    .X(_08845_));
 sg13g2_and2_1 _17579_ (.A(_08844_),
    .B(_08845_),
    .X(_00859_));
 sg13g2_nor2_2 _17580_ (.A(_04303_),
    .B(_08844_),
    .Y(_08846_));
 sg13g2_a21oi_1 _17581_ (.A1(_04303_),
    .A2(_08844_),
    .Y(_08847_),
    .B1(_08842_));
 sg13g2_nor2b_1 _17582_ (.A(_08846_),
    .B_N(_08847_),
    .Y(_00860_));
 sg13g2_a21oi_1 _17583_ (.A1(net3169),
    .A2(_08843_),
    .Y(_08848_),
    .B1(_08846_));
 sg13g2_a21oi_1 _17584_ (.A1(net3169),
    .A2(_08846_),
    .Y(_00861_),
    .B1(_08848_));
 sg13g2_and3_1 _17585_ (.X(_08849_),
    .A(net3169),
    .B(net2400),
    .C(_08846_));
 sg13g2_a21oi_1 _17586_ (.A1(\TRNG.uart_tx_inst.ticks_counter[5] ),
    .A2(_08846_),
    .Y(_08850_),
    .B1(net2400));
 sg13g2_nor2_1 _17587_ (.A(_08849_),
    .B(net2401),
    .Y(_00862_));
 sg13g2_o21ai_1 _17588_ (.B1(_08843_),
    .Y(_08851_),
    .A1(net3418),
    .A2(_08849_));
 sg13g2_nand2_1 _17589_ (.Y(_08852_),
    .A(net3418),
    .B(_08849_));
 sg13g2_nor2b_1 _17590_ (.A(_08851_),
    .B_N(_08852_),
    .Y(_00863_));
 sg13g2_xor2_1 _17591_ (.B(_08852_),
    .A(net3269),
    .X(_08853_));
 sg13g2_nor2_1 _17592_ (.A(_08842_),
    .B(net3270),
    .Y(_00864_));
 sg13g2_nor2_2 _17593_ (.A(net5207),
    .B(_06913_),
    .Y(_08854_));
 sg13g2_mux2_1 _17594_ (.A0(net2817),
    .A1(net5689),
    .S(net5028),
    .X(_00865_));
 sg13g2_mux2_1 _17595_ (.A0(net2841),
    .A1(net5688),
    .S(net5028),
    .X(_00866_));
 sg13g2_mux2_1 _17596_ (.A0(net2642),
    .A1(net5686),
    .S(net5029),
    .X(_00867_));
 sg13g2_nor2_1 _17597_ (.A(net2874),
    .B(net5030),
    .Y(_08855_));
 sg13g2_a21oi_1 _17598_ (.A1(net5495),
    .A2(net5030),
    .Y(_00868_),
    .B1(_08855_));
 sg13g2_mux2_1 _17599_ (.A0(net2927),
    .A1(net5682),
    .S(net5029),
    .X(_00869_));
 sg13g2_mux2_1 _17600_ (.A0(net2677),
    .A1(net5679),
    .S(net5029),
    .X(_00870_));
 sg13g2_mux2_1 _17601_ (.A0(net2741),
    .A1(net5676),
    .S(net5029),
    .X(_00871_));
 sg13g2_mux2_1 _17602_ (.A0(net2645),
    .A1(net5675),
    .S(net5031),
    .X(_00872_));
 sg13g2_mux2_1 _17603_ (.A0(net2929),
    .A1(net5671),
    .S(net5031),
    .X(_00873_));
 sg13g2_mux2_1 _17604_ (.A0(net2796),
    .A1(net5669),
    .S(net5031),
    .X(_00874_));
 sg13g2_mux2_1 _17605_ (.A0(net2780),
    .A1(net5668),
    .S(net5032),
    .X(_00875_));
 sg13g2_mux2_1 _17606_ (.A0(net2777),
    .A1(net5666),
    .S(net5028),
    .X(_00876_));
 sg13g2_mux2_1 _17607_ (.A0(net2726),
    .A1(net5664),
    .S(net5028),
    .X(_00877_));
 sg13g2_mux2_1 _17608_ (.A0(net2764),
    .A1(net5661),
    .S(net5028),
    .X(_00878_));
 sg13g2_mux2_1 _17609_ (.A0(net2621),
    .A1(net5659),
    .S(net5031),
    .X(_00879_));
 sg13g2_mux2_1 _17610_ (.A0(net2672),
    .A1(net5657),
    .S(net5030),
    .X(_00880_));
 sg13g2_mux2_1 _17611_ (.A0(net2707),
    .A1(net5654),
    .S(net5031),
    .X(_00881_));
 sg13g2_mux2_1 _17612_ (.A0(net2815),
    .A1(net5652),
    .S(net5030),
    .X(_00882_));
 sg13g2_mux2_1 _17613_ (.A0(net2857),
    .A1(net5650),
    .S(net5028),
    .X(_00883_));
 sg13g2_mux2_1 _17614_ (.A0(net2600),
    .A1(net5647),
    .S(net5028),
    .X(_00884_));
 sg13g2_mux2_1 _17615_ (.A0(net2739),
    .A1(net5645),
    .S(net5030),
    .X(_00885_));
 sg13g2_mux2_1 _17616_ (.A0(net2788),
    .A1(net5641),
    .S(net5032),
    .X(_00886_));
 sg13g2_mux2_1 _17617_ (.A0(net2601),
    .A1(net5639),
    .S(net5030),
    .X(_00887_));
 sg13g2_mux2_1 _17618_ (.A0(net2665),
    .A1(net5636),
    .S(net5030),
    .X(_00888_));
 sg13g2_mux2_1 _17619_ (.A0(net2783),
    .A1(net5634),
    .S(net5032),
    .X(_00889_));
 sg13g2_mux2_1 _17620_ (.A0(net2650),
    .A1(net5632),
    .S(net5030),
    .X(_00890_));
 sg13g2_mux2_1 _17621_ (.A0(net2836),
    .A1(net5629),
    .S(net5032),
    .X(_00891_));
 sg13g2_mux2_1 _17622_ (.A0(net2806),
    .A1(net5628),
    .S(net5029),
    .X(_00892_));
 sg13g2_mux2_1 _17623_ (.A0(net2693),
    .A1(net5624),
    .S(net5031),
    .X(_00893_));
 sg13g2_mux2_1 _17624_ (.A0(net2894),
    .A1(net5623),
    .S(net5031),
    .X(_00894_));
 sg13g2_mux2_1 _17625_ (.A0(net2813),
    .A1(net5618),
    .S(net5028),
    .X(_00895_));
 sg13g2_mux2_1 _17626_ (.A0(net2871),
    .A1(net5617),
    .S(net5031),
    .X(_00896_));
 sg13g2_nand2b_2 _17627_ (.Y(_08856_),
    .B(_08805_),
    .A_N(net5874));
 sg13g2_nor2_1 _17628_ (.A(_08803_),
    .B(_08856_),
    .Y(_08857_));
 sg13g2_nor3_1 _17629_ (.A(net5875),
    .B(_08813_),
    .C(_08834_),
    .Y(_08858_));
 sg13g2_nor2_1 _17630_ (.A(_08808_),
    .B(_08813_),
    .Y(_08859_));
 sg13g2_nand3_1 _17631_ (.B(net5874),
    .C(_00118_),
    .A(net5873),
    .Y(_08860_));
 sg13g2_nor2_2 _17632_ (.A(net5342),
    .B(_08860_),
    .Y(_08861_));
 sg13g2_nor3_1 _17633_ (.A(net5875),
    .B(_06870_),
    .C(_08813_),
    .Y(_08862_));
 sg13g2_nor2_1 _17634_ (.A(_06870_),
    .B(_08856_),
    .Y(_08863_));
 sg13g2_nor2_1 _17635_ (.A(_06868_),
    .B(_08808_),
    .Y(_08864_));
 sg13g2_nand2b_2 _17636_ (.Y(_08865_),
    .B(\TRNG.sha256.compress.count[1] ),
    .A_N(\TRNG.sha256.compress.count[0] ));
 sg13g2_nor3_1 _17637_ (.A(net5875),
    .B(_06868_),
    .C(_08865_),
    .Y(_08866_));
 sg13g2_nor2_1 _17638_ (.A(_08856_),
    .B(_08865_),
    .Y(_08867_));
 sg13g2_nor3_1 _17639_ (.A(net5875),
    .B(_06870_),
    .C(_08806_),
    .Y(_08868_));
 sg13g2_nor3_2 _17640_ (.A(net5875),
    .B(_08813_),
    .C(_08865_),
    .Y(_08869_));
 sg13g2_nand2_1 _17641_ (.Y(_08870_),
    .A(net3737),
    .B(net5126));
 sg13g2_nor3_1 _17642_ (.A(net5875),
    .B(_06868_),
    .C(net5342),
    .Y(_08871_));
 sg13g2_inv_1 _17643_ (.Y(_08872_),
    .A(net5123));
 sg13g2_nor2_1 _17644_ (.A(_08834_),
    .B(_08856_),
    .Y(_08873_));
 sg13g2_a22oi_1 _17645_ (.Y(_08874_),
    .B1(net5135),
    .B2(\TRNG.Padded_Out[416] ),
    .A2(net5141),
    .A1(\TRNG.Padded_Out[352] ));
 sg13g2_a22oi_1 _17646_ (.Y(_08875_),
    .B1(net5004),
    .B2(\TRNG.Padded_Out[160] ),
    .A2(net5010),
    .A1(\TRNG.Padded_Out[384] ));
 sg13g2_a22oi_1 _17647_ (.Y(_08876_),
    .B1(net5131),
    .B2(\TRNG.Padded_Out[96] ),
    .A2(net5024),
    .A1(\TRNG.Padded_Out[128] ));
 sg13g2_a22oi_1 _17648_ (.Y(_08877_),
    .B1(net5146),
    .B2(\TRNG.Padded_Out[64] ),
    .A2(net5150),
    .A1(\TRNG.Padded_Out[320] ));
 sg13g2_a22oi_1 _17649_ (.Y(_08878_),
    .B1(net5121),
    .B2(\TRNG.Padded_Out[448] ),
    .A2(net5022),
    .A1(\TRNG.Padded_Out[256] ));
 sg13g2_a22oi_1 _17650_ (.Y(_08879_),
    .B1(net4998),
    .B2(\TRNG.Padded_Out[192] ),
    .A2(net5014),
    .A1(\TRNG.Padded_Out[224] ));
 sg13g2_nand3_1 _17651_ (.B(_08878_),
    .C(_08879_),
    .A(_08874_),
    .Y(_08880_));
 sg13g2_nand4_1 _17652_ (.B(_08875_),
    .C(_08876_),
    .A(_08870_),
    .Y(_08881_),
    .D(_08877_));
 sg13g2_nor2_2 _17653_ (.A(_08880_),
    .B(_08881_),
    .Y(_08882_));
 sg13g2_nor2_1 _17654_ (.A(_06869_),
    .B(_08806_),
    .Y(_08883_));
 sg13g2_nor3_1 _17655_ (.A(net5875),
    .B(_06871_),
    .C(_08883_),
    .Y(_08884_));
 sg13g2_nor2_1 _17656_ (.A(_08836_),
    .B(_08860_),
    .Y(_08885_));
 sg13g2_nor2_1 _17657_ (.A(_08884_),
    .B(_08885_),
    .Y(_08886_));
 sg13g2_nand3_1 _17658_ (.B(_08810_),
    .C(net4959),
    .A(net5090),
    .Y(_08887_));
 sg13g2_nor2_1 _17659_ (.A(_08809_),
    .B(net5156),
    .Y(_08888_));
 sg13g2_nand2_1 _17660_ (.Y(_08889_),
    .A(net4959),
    .B(net4958));
 sg13g2_nor2_1 _17661_ (.A(net5093),
    .B(_08889_),
    .Y(_08890_));
 sg13g2_nand3_1 _17662_ (.B(net4959),
    .C(net4958),
    .A(net5090),
    .Y(_08891_));
 sg13g2_nor3_1 _17663_ (.A(_04271_),
    .B(net5343),
    .C(net5341),
    .Y(_08892_));
 sg13g2_a221oi_1 _17664_ (.B2(\TRNG.sha256.W[0] ),
    .C1(_08892_),
    .B1(net4567),
    .A1(net2539),
    .Y(_08893_),
    .A2(net5091));
 sg13g2_a21oi_1 _17665_ (.A1(_08882_),
    .A2(_08893_),
    .Y(_00897_),
    .B1(net5531));
 sg13g2_a22oi_1 _17666_ (.Y(_08894_),
    .B1(net5004),
    .B2(\TRNG.Padded_Out[161] ),
    .A2(net5010),
    .A1(\TRNG.Padded_Out[385] ));
 sg13g2_nand2_1 _17667_ (.Y(_08895_),
    .A(\TRNG.Padded_Out[225] ),
    .B(net5014));
 sg13g2_a22oi_1 _17668_ (.Y(_08896_),
    .B1(net5126),
    .B2(\TRNG.Padded_Out[289] ),
    .A2(net5135),
    .A1(\TRNG.Padded_Out[417] ));
 sg13g2_a22oi_1 _17669_ (.Y(_08897_),
    .B1(net5121),
    .B2(\TRNG.Padded_Out[449] ),
    .A2(net5019),
    .A1(\TRNG.Padded_Out[257] ));
 sg13g2_a22oi_1 _17670_ (.Y(_08898_),
    .B1(net4998),
    .B2(\TRNG.Padded_Out[193] ),
    .A2(net5150),
    .A1(\TRNG.Padded_Out[321] ));
 sg13g2_a22oi_1 _17671_ (.Y(_08899_),
    .B1(net5131),
    .B2(\TRNG.Padded_Out[97] ),
    .A2(net5146),
    .A1(\TRNG.Padded_Out[65] ));
 sg13g2_nand3_1 _17672_ (.B(_08895_),
    .C(_08899_),
    .A(_08894_),
    .Y(_08900_));
 sg13g2_a221oi_1 _17673_ (.B2(\TRNG.Padded_Out[353] ),
    .C1(_08900_),
    .B1(net5144),
    .A1(\TRNG.Padded_Out[129] ),
    .Y(_08901_),
    .A2(net5024));
 sg13g2_nand4_1 _17674_ (.B(_08897_),
    .C(_08898_),
    .A(_08896_),
    .Y(_08902_),
    .D(_08901_));
 sg13g2_a22oi_1 _17675_ (.Y(_08903_),
    .B1(net4568),
    .B2(net3371),
    .A2(net5091),
    .A1(net2354));
 sg13g2_a21oi_1 _17676_ (.A1(net2352),
    .A2(net5155),
    .Y(_08904_),
    .B1(_08902_));
 sg13g2_a21oi_1 _17677_ (.A1(_08903_),
    .A2(_08904_),
    .Y(_00898_),
    .B1(net5531));
 sg13g2_nand2_1 _17678_ (.Y(_08905_),
    .A(\TRNG.Padded_Out[322] ),
    .B(net5150));
 sg13g2_a22oi_1 _17679_ (.Y(_08906_),
    .B1(net5146),
    .B2(\TRNG.Padded_Out[66] ),
    .A2(net5024),
    .A1(\TRNG.Padded_Out[130] ));
 sg13g2_a22oi_1 _17680_ (.Y(_08907_),
    .B1(net5121),
    .B2(\TRNG.Padded_Out[450] ),
    .A2(net5004),
    .A1(\TRNG.Padded_Out[162] ));
 sg13g2_a22oi_1 _17681_ (.Y(_08908_),
    .B1(net5135),
    .B2(\TRNG.Padded_Out[418] ),
    .A2(net5010),
    .A1(\TRNG.Padded_Out[386] ));
 sg13g2_a22oi_1 _17682_ (.Y(_08909_),
    .B1(net5131),
    .B2(\TRNG.Padded_Out[98] ),
    .A2(net5019),
    .A1(\TRNG.Padded_Out[258] ));
 sg13g2_a22oi_1 _17683_ (.Y(_08910_),
    .B1(net4998),
    .B2(\TRNG.Padded_Out[194] ),
    .A2(net5126),
    .A1(\TRNG.Padded_Out[290] ));
 sg13g2_nand3_1 _17684_ (.B(_08907_),
    .C(_08908_),
    .A(_08905_),
    .Y(_08911_));
 sg13g2_a221oi_1 _17685_ (.B2(\TRNG.Padded_Out[226] ),
    .C1(_08911_),
    .B1(net5014),
    .A1(\TRNG.Padded_Out[354] ),
    .Y(_08912_),
    .A2(net5141));
 sg13g2_nand4_1 _17686_ (.B(_08909_),
    .C(_08910_),
    .A(_08906_),
    .Y(_08913_),
    .D(_08912_));
 sg13g2_a221oi_1 _17687_ (.B2(net4958),
    .C1(_08913_),
    .B1(net4959),
    .A1(net2265),
    .Y(_08914_),
    .A2(net5157));
 sg13g2_a21oi_1 _17688_ (.A1(_04311_),
    .A2(net5093),
    .Y(_08915_),
    .B1(net5534));
 sg13g2_o21ai_1 _17689_ (.B1(_08915_),
    .Y(_08916_),
    .A1(\TRNG.sha256.W[2] ),
    .A2(_08891_));
 sg13g2_nor2_1 _17690_ (.A(_08914_),
    .B(_08916_),
    .Y(_00899_));
 sg13g2_a22oi_1 _17691_ (.Y(_08917_),
    .B1(net5126),
    .B2(\TRNG.Padded_Out[291] ),
    .A2(net5131),
    .A1(\TRNG.Padded_Out[99] ));
 sg13g2_a22oi_1 _17692_ (.Y(_08918_),
    .B1(net5010),
    .B2(\TRNG.Padded_Out[387] ),
    .A2(net5150),
    .A1(\TRNG.Padded_Out[323] ));
 sg13g2_a22oi_1 _17693_ (.Y(_08919_),
    .B1(net5121),
    .B2(\TRNG.Padded_Out[451] ),
    .A2(net5135),
    .A1(\TRNG.Padded_Out[419] ));
 sg13g2_a22oi_1 _17694_ (.Y(_08920_),
    .B1(net4998),
    .B2(\TRNG.Padded_Out[195] ),
    .A2(net5024),
    .A1(\TRNG.Padded_Out[131] ));
 sg13g2_a22oi_1 _17695_ (.Y(_08921_),
    .B1(net5004),
    .B2(\TRNG.Padded_Out[163] ),
    .A2(net5141),
    .A1(\TRNG.Padded_Out[355] ));
 sg13g2_a22oi_1 _17696_ (.Y(_08922_),
    .B1(net5014),
    .B2(\TRNG.Padded_Out[227] ),
    .A2(net5019),
    .A1(\TRNG.Padded_Out[259] ));
 sg13g2_nand2_1 _17697_ (.Y(_08923_),
    .A(_08919_),
    .B(_08922_));
 sg13g2_nand4_1 _17698_ (.B(_08918_),
    .C(_08920_),
    .A(_08917_),
    .Y(_08924_),
    .D(_08921_));
 sg13g2_nor2_2 _17699_ (.A(_08923_),
    .B(_08924_),
    .Y(_08925_));
 sg13g2_a22oi_1 _17700_ (.Y(_08926_),
    .B1(net5149),
    .B2(net3589),
    .A2(net5157),
    .A1(net2403));
 sg13g2_and2_1 _17701_ (.A(_08889_),
    .B(_08926_),
    .X(_08927_));
 sg13g2_a21oi_1 _17702_ (.A1(_04312_),
    .A2(net5093),
    .Y(_08928_),
    .B1(net5535));
 sg13g2_o21ai_1 _17703_ (.B1(_08928_),
    .Y(_08929_),
    .A1(\TRNG.sha256.W[3] ),
    .A2(_08891_));
 sg13g2_a21oi_1 _17704_ (.A1(_08925_),
    .A2(_08927_),
    .Y(_00900_),
    .B1(_08929_));
 sg13g2_a22oi_1 _17705_ (.Y(_08930_),
    .B1(net5126),
    .B2(\TRNG.Padded_Out[292] ),
    .A2(net5150),
    .A1(\TRNG.Padded_Out[324] ));
 sg13g2_a22oi_1 _17706_ (.Y(_08931_),
    .B1(net5135),
    .B2(\TRNG.Padded_Out[420] ),
    .A2(net5022),
    .A1(\TRNG.Padded_Out[260] ));
 sg13g2_a22oi_1 _17707_ (.Y(_08932_),
    .B1(net5141),
    .B2(\TRNG.Padded_Out[356] ),
    .A2(net5027),
    .A1(\TRNG.Padded_Out[132] ));
 sg13g2_nand3_1 _17708_ (.B(_08931_),
    .C(_08932_),
    .A(_08930_),
    .Y(_08933_));
 sg13g2_nand2_1 _17709_ (.Y(_08934_),
    .A(\TRNG.Padded_Out[228] ),
    .B(net5014));
 sg13g2_a22oi_1 _17710_ (.Y(_08935_),
    .B1(net4998),
    .B2(\TRNG.Padded_Out[196] ),
    .A2(net5131),
    .A1(\TRNG.Padded_Out[100] ));
 sg13g2_a22oi_1 _17711_ (.Y(_08936_),
    .B1(net5011),
    .B2(\TRNG.Padded_Out[388] ),
    .A2(net5146),
    .A1(\TRNG.Padded_Out[68] ));
 sg13g2_a22oi_1 _17712_ (.Y(_08937_),
    .B1(net5121),
    .B2(\TRNG.Padded_Out[452] ),
    .A2(net5004),
    .A1(\TRNG.Padded_Out[164] ));
 sg13g2_nand4_1 _17713_ (.B(_08935_),
    .C(_08936_),
    .A(_08934_),
    .Y(_08938_),
    .D(_08937_));
 sg13g2_nor2_2 _17714_ (.A(_08933_),
    .B(_08938_),
    .Y(_08939_));
 sg13g2_nand2_1 _17715_ (.Y(_08940_),
    .A(net2307),
    .B(net5157));
 sg13g2_and2_1 _17716_ (.A(_08939_),
    .B(_08940_),
    .X(_08941_));
 sg13g2_a22oi_1 _17717_ (.Y(_08942_),
    .B1(net4569),
    .B2(net3478),
    .A2(net5094),
    .A1(net2809));
 sg13g2_a21oi_1 _17718_ (.A1(_08941_),
    .A2(_08942_),
    .Y(_00901_),
    .B1(net5535));
 sg13g2_nand2_1 _17719_ (.Y(_08943_),
    .A(\TRNG.Padded_Out[421] ),
    .B(net5135));
 sg13g2_a22oi_1 _17720_ (.Y(_08944_),
    .B1(net5011),
    .B2(\TRNG.Padded_Out[389] ),
    .A2(net5154),
    .A1(\TRNG.Padded_Out[325] ));
 sg13g2_a22oi_1 _17721_ (.Y(_08945_),
    .B1(net5014),
    .B2(\TRNG.Padded_Out[229] ),
    .A2(net5024),
    .A1(\TRNG.Padded_Out[133] ));
 sg13g2_a22oi_1 _17722_ (.Y(_08946_),
    .B1(net4998),
    .B2(\TRNG.Padded_Out[197] ),
    .A2(net5019),
    .A1(\TRNG.Padded_Out[261] ));
 sg13g2_a22oi_1 _17723_ (.Y(_08947_),
    .B1(net5121),
    .B2(\TRNG.Padded_Out[453] ),
    .A2(net5004),
    .A1(\TRNG.Padded_Out[165] ));
 sg13g2_a22oi_1 _17724_ (.Y(_08948_),
    .B1(net5126),
    .B2(\TRNG.Padded_Out[293] ),
    .A2(net5146),
    .A1(\TRNG.Padded_Out[69] ));
 sg13g2_nand3_1 _17725_ (.B(_08947_),
    .C(_08948_),
    .A(_08943_),
    .Y(_08949_));
 sg13g2_a221oi_1 _17726_ (.B2(\TRNG.Padded_Out[101] ),
    .C1(_08949_),
    .B1(net5131),
    .A1(\TRNG.Padded_Out[357] ),
    .Y(_08950_),
    .A2(net5141));
 sg13g2_nand4_1 _17727_ (.B(_08945_),
    .C(_08946_),
    .A(_08944_),
    .Y(_08951_),
    .D(_08950_));
 sg13g2_a22oi_1 _17728_ (.Y(_08952_),
    .B1(net4570),
    .B2(net3375),
    .A2(net5094),
    .A1(net2860));
 sg13g2_a21oi_1 _17729_ (.A1(net2038),
    .A2(net5157),
    .Y(_08953_),
    .B1(_08951_));
 sg13g2_a21oi_1 _17730_ (.A1(_08952_),
    .A2(_08953_),
    .Y(_00902_),
    .B1(net5537));
 sg13g2_a22oi_1 _17731_ (.Y(_08954_),
    .B1(net5004),
    .B2(\TRNG.Padded_Out[166] ),
    .A2(net5135),
    .A1(\TRNG.Padded_Out[422] ));
 sg13g2_a22oi_1 _17732_ (.Y(_08955_),
    .B1(net5014),
    .B2(\TRNG.Padded_Out[230] ),
    .A2(net5146),
    .A1(\TRNG.Padded_Out[70] ));
 sg13g2_a22oi_1 _17733_ (.Y(_08956_),
    .B1(net5131),
    .B2(\TRNG.Padded_Out[102] ),
    .A2(net5150),
    .A1(\TRNG.Padded_Out[326] ));
 sg13g2_a22oi_1 _17734_ (.Y(_08957_),
    .B1(net5002),
    .B2(\TRNG.Padded_Out[198] ),
    .A2(net5010),
    .A1(\TRNG.Padded_Out[390] ));
 sg13g2_a22oi_1 _17735_ (.Y(_08958_),
    .B1(net5122),
    .B2(\TRNG.Padded_Out[454] ),
    .A2(net5019),
    .A1(\TRNG.Padded_Out[262] ));
 sg13g2_a22oi_1 _17736_ (.Y(_08959_),
    .B1(net5126),
    .B2(\TRNG.Padded_Out[294] ),
    .A2(net5141),
    .A1(\TRNG.Padded_Out[358] ));
 sg13g2_nand3_1 _17737_ (.B(_08955_),
    .C(_08959_),
    .A(_08954_),
    .Y(_08960_));
 sg13g2_a221oi_1 _17738_ (.B2(\TRNG.Padded_Out[134] ),
    .C1(_08960_),
    .B1(net5024),
    .A1(\TRNG.Padded_Out[64] ),
    .Y(_08961_),
    .A2(_08809_));
 sg13g2_nand4_1 _17739_ (.B(_08957_),
    .C(_08958_),
    .A(_08956_),
    .Y(_08962_),
    .D(_08961_));
 sg13g2_a221oi_1 _17740_ (.B2(net4958),
    .C1(_08962_),
    .B1(net4959),
    .A1(net2299),
    .Y(_08963_),
    .A2(net5156));
 sg13g2_a21oi_1 _17741_ (.A1(_04315_),
    .A2(net5093),
    .Y(_08964_),
    .B1(net5537));
 sg13g2_o21ai_1 _17742_ (.B1(_08964_),
    .Y(_08965_),
    .A1(\TRNG.sha256.W[6] ),
    .A2(_08891_));
 sg13g2_nor2_1 _17743_ (.A(_08963_),
    .B(_08965_),
    .Y(_00903_));
 sg13g2_a22oi_1 _17744_ (.Y(_08966_),
    .B1(net4998),
    .B2(\TRNG.Padded_Out[199] ),
    .A2(net5010),
    .A1(\TRNG.Padded_Out[391] ));
 sg13g2_a22oi_1 _17745_ (.Y(_08967_),
    .B1(net5121),
    .B2(\TRNG.Padded_Out[455] ),
    .A2(net5126),
    .A1(\TRNG.Padded_Out[295] ));
 sg13g2_a22oi_1 _17746_ (.Y(_08968_),
    .B1(net5134),
    .B2(\TRNG.Padded_Out[103] ),
    .A2(net5016),
    .A1(\TRNG.Padded_Out[231] ));
 sg13g2_a22oi_1 _17747_ (.Y(_08969_),
    .B1(net5027),
    .B2(\TRNG.Padded_Out[135] ),
    .A2(_08809_),
    .A1(\TRNG.Padded_Out[64] ));
 sg13g2_a22oi_1 _17748_ (.Y(_08970_),
    .B1(net5143),
    .B2(\TRNG.Padded_Out[359] ),
    .A2(net5021),
    .A1(\TRNG.Padded_Out[263] ));
 sg13g2_nand3_1 _17749_ (.B(_08969_),
    .C(_08970_),
    .A(_08968_),
    .Y(_08971_));
 sg13g2_a22oi_1 _17750_ (.Y(_08972_),
    .B1(net5135),
    .B2(\TRNG.Padded_Out[423] ),
    .A2(net5148),
    .A1(\TRNG.Padded_Out[71] ));
 sg13g2_a22oi_1 _17751_ (.Y(_08973_),
    .B1(net5006),
    .B2(\TRNG.Padded_Out[167] ),
    .A2(net5150),
    .A1(\TRNG.Padded_Out[327] ));
 sg13g2_nand4_1 _17752_ (.B(_08967_),
    .C(_08972_),
    .A(_08966_),
    .Y(_08974_),
    .D(_08973_));
 sg13g2_or2_2 _17753_ (.X(_08975_),
    .B(_08974_),
    .A(_08971_));
 sg13g2_a221oi_1 _17754_ (.B2(net4958),
    .C1(_08975_),
    .B1(net4959),
    .A1(net2226),
    .Y(_08976_),
    .A2(net5156));
 sg13g2_a21oi_1 _17755_ (.A1(_04316_),
    .A2(net5093),
    .Y(_08977_),
    .B1(net5537));
 sg13g2_o21ai_1 _17756_ (.B1(_08977_),
    .Y(_08978_),
    .A1(\TRNG.sha256.W[7] ),
    .A2(_08891_));
 sg13g2_nor2_1 _17757_ (.A(_08976_),
    .B(_08978_),
    .Y(_00904_));
 sg13g2_a22oi_1 _17758_ (.Y(_08979_),
    .B1(net5138),
    .B2(\TRNG.Padded_Out[424] ),
    .A2(net5012),
    .A1(\TRNG.Padded_Out[392] ));
 sg13g2_a22oi_1 _17759_ (.Y(_08980_),
    .B1(net5144),
    .B2(\TRNG.Padded_Out[360] ),
    .A2(net5026),
    .A1(\TRNG.Padded_Out[136] ));
 sg13g2_a22oi_1 _17760_ (.Y(_08981_),
    .B1(net5133),
    .B2(\TRNG.Padded_Out[104] ),
    .A2(_08809_),
    .A1(\TRNG.Padded_Out[64] ));
 sg13g2_a22oi_1 _17761_ (.Y(_08982_),
    .B1(net5129),
    .B2(\TRNG.Padded_Out[296] ),
    .A2(net5148),
    .A1(\TRNG.Padded_Out[72] ));
 sg13g2_nand3_1 _17762_ (.B(_08981_),
    .C(_08982_),
    .A(_08980_),
    .Y(_08983_));
 sg13g2_a22oi_1 _17763_ (.Y(_08984_),
    .B1(net5002),
    .B2(\TRNG.Padded_Out[200] ),
    .A2(net5006),
    .A1(\TRNG.Padded_Out[168] ));
 sg13g2_a22oi_1 _17764_ (.Y(_08985_),
    .B1(net5122),
    .B2(\TRNG.Padded_Out[456] ),
    .A2(net5153),
    .A1(\TRNG.Padded_Out[328] ));
 sg13g2_a22oi_1 _17765_ (.Y(_08986_),
    .B1(net5017),
    .B2(\TRNG.Padded_Out[232] ),
    .A2(net5021),
    .A1(\TRNG.Padded_Out[264] ));
 sg13g2_nand4_1 _17766_ (.B(_08984_),
    .C(_08985_),
    .A(_08979_),
    .Y(_08987_),
    .D(_08986_));
 sg13g2_or2_2 _17767_ (.X(_08988_),
    .B(_08987_),
    .A(_08983_));
 sg13g2_a221oi_1 _17768_ (.B2(net4958),
    .C1(_08988_),
    .B1(net4959),
    .A1(net2415),
    .Y(_08989_),
    .A2(net5156));
 sg13g2_a21oi_1 _17769_ (.A1(_04317_),
    .A2(net5093),
    .Y(_08990_),
    .B1(net5537));
 sg13g2_o21ai_1 _17770_ (.B1(_08990_),
    .Y(_08991_),
    .A1(\TRNG.sha256.W[8] ),
    .A2(_08891_));
 sg13g2_nor2_1 _17771_ (.A(_08989_),
    .B(_08991_),
    .Y(_00905_));
 sg13g2_a22oi_1 _17772_ (.Y(_08992_),
    .B1(net5001),
    .B2(net3708),
    .A2(net5148),
    .A1(\TRNG.Padded_Out[73] ));
 sg13g2_a22oi_1 _17773_ (.Y(_08993_),
    .B1(net5016),
    .B2(\TRNG.Padded_Out[233] ),
    .A2(net5153),
    .A1(\TRNG.Padded_Out[329] ));
 sg13g2_a22oi_1 _17774_ (.Y(_08994_),
    .B1(net5138),
    .B2(\TRNG.Padded_Out[425] ),
    .A2(net5026),
    .A1(\TRNG.Padded_Out[137] ));
 sg13g2_nand3_1 _17775_ (.B(_08993_),
    .C(_08994_),
    .A(_08992_),
    .Y(_08995_));
 sg13g2_nand2_1 _17776_ (.Y(_08996_),
    .A(\TRNG.Padded_Out[457] ),
    .B(net5124));
 sg13g2_a22oi_1 _17777_ (.Y(_08997_),
    .B1(net5011),
    .B2(\TRNG.Padded_Out[393] ),
    .A2(net5143),
    .A1(\TRNG.Padded_Out[361] ));
 sg13g2_a22oi_1 _17778_ (.Y(_08998_),
    .B1(net5006),
    .B2(\TRNG.Padded_Out[169] ),
    .A2(net5021),
    .A1(\TRNG.Padded_Out[265] ));
 sg13g2_a22oi_1 _17779_ (.Y(_08999_),
    .B1(net5129),
    .B2(\TRNG.Padded_Out[297] ),
    .A2(net5133),
    .A1(\TRNG.Padded_Out[105] ));
 sg13g2_nand4_1 _17780_ (.B(_08997_),
    .C(_08998_),
    .A(_08996_),
    .Y(_09000_),
    .D(_08999_));
 sg13g2_nor2_2 _17781_ (.A(_08995_),
    .B(_09000_),
    .Y(_09001_));
 sg13g2_nor3_1 _17782_ (.A(_04262_),
    .B(net5344),
    .C(net5342),
    .Y(_09002_));
 sg13g2_a221oi_1 _17783_ (.B2(\TRNG.sha256.W[9] ),
    .C1(_09002_),
    .B1(net4570),
    .A1(net2582),
    .Y(_09003_),
    .A2(net5093));
 sg13g2_a21oi_1 _17784_ (.A1(net3709),
    .A2(_09003_),
    .Y(_00906_),
    .B1(net5543));
 sg13g2_nand2_1 _17785_ (.Y(_09004_),
    .A(\TRNG.Padded_Out[394] ),
    .B(net5011));
 sg13g2_a22oi_1 _17786_ (.Y(_09005_),
    .B1(net5001),
    .B2(net1408),
    .A2(net5153),
    .A1(\TRNG.Padded_Out[330] ));
 sg13g2_a22oi_1 _17787_ (.Y(_09006_),
    .B1(net5006),
    .B2(\TRNG.Padded_Out[170] ),
    .A2(net5138),
    .A1(\TRNG.Padded_Out[426] ));
 sg13g2_a22oi_1 _17788_ (.Y(_09007_),
    .B1(net5016),
    .B2(\TRNG.Padded_Out[234] ),
    .A2(net5143),
    .A1(\TRNG.Padded_Out[362] ));
 sg13g2_a22oi_1 _17789_ (.Y(_09008_),
    .B1(net5124),
    .B2(\TRNG.Padded_Out[458] ),
    .A2(net5148),
    .A1(\TRNG.Padded_Out[74] ));
 sg13g2_nand3_1 _17790_ (.B(_09007_),
    .C(_09008_),
    .A(_09005_),
    .Y(_09009_));
 sg13g2_a22oi_1 _17791_ (.Y(_09010_),
    .B1(net5021),
    .B2(\TRNG.Padded_Out[266] ),
    .A2(net5026),
    .A1(\TRNG.Padded_Out[138] ));
 sg13g2_a22oi_1 _17792_ (.Y(_09011_),
    .B1(net5128),
    .B2(\TRNG.Padded_Out[298] ),
    .A2(net5133),
    .A1(\TRNG.Padded_Out[106] ));
 sg13g2_nand4_1 _17793_ (.B(_09006_),
    .C(_09010_),
    .A(_09004_),
    .Y(_09012_),
    .D(_09011_));
 sg13g2_nor2_2 _17794_ (.A(_09009_),
    .B(_09012_),
    .Y(_09013_));
 sg13g2_nor3_1 _17795_ (.A(_04261_),
    .B(net5344),
    .C(net5342),
    .Y(_09014_));
 sg13g2_a221oi_1 _17796_ (.B2(\TRNG.sha256.W[10] ),
    .C1(_09014_),
    .B1(net4569),
    .A1(net2480),
    .Y(_09015_),
    .A2(net5095));
 sg13g2_a21oi_1 _17797_ (.A1(_09013_),
    .A2(_09015_),
    .Y(_00907_),
    .B1(net5534));
 sg13g2_nand2_1 _17798_ (.Y(_09016_),
    .A(net1810),
    .B(net5021));
 sg13g2_a22oi_1 _17799_ (.Y(_09017_),
    .B1(net5133),
    .B2(\TRNG.Padded_Out[107] ),
    .A2(net5011),
    .A1(\TRNG.Padded_Out[395] ));
 sg13g2_a22oi_1 _17800_ (.Y(_09018_),
    .B1(net5006),
    .B2(net1849),
    .A2(net5143),
    .A1(\TRNG.Padded_Out[363] ));
 sg13g2_a22oi_1 _17801_ (.Y(_09019_),
    .B1(net5121),
    .B2(\TRNG.Padded_Out[459] ),
    .A2(net5153),
    .A1(\TRNG.Padded_Out[331] ));
 sg13g2_a22oi_1 _17802_ (.Y(_09020_),
    .B1(net5138),
    .B2(\TRNG.Padded_Out[427] ),
    .A2(net5026),
    .A1(\TRNG.Padded_Out[139] ));
 sg13g2_a22oi_1 _17803_ (.Y(_09021_),
    .B1(net5001),
    .B2(net3697),
    .A2(net5016),
    .A1(\TRNG.Padded_Out[235] ));
 sg13g2_a22oi_1 _17804_ (.Y(_09022_),
    .B1(net5129),
    .B2(\TRNG.Padded_Out[299] ),
    .A2(net5149),
    .A1(\TRNG.Padded_Out[75] ));
 sg13g2_nand3_1 _17805_ (.B(_09021_),
    .C(_09022_),
    .A(_09017_),
    .Y(_09023_));
 sg13g2_nand4_1 _17806_ (.B(_09018_),
    .C(_09019_),
    .A(_09016_),
    .Y(_09024_),
    .D(_09020_));
 sg13g2_nor2_2 _17807_ (.A(_09023_),
    .B(_09024_),
    .Y(_09025_));
 sg13g2_nor3_1 _17808_ (.A(_04260_),
    .B(net5343),
    .C(net5341),
    .Y(_09026_));
 sg13g2_a221oi_1 _17809_ (.B2(\TRNG.sha256.W[11] ),
    .C1(_09026_),
    .B1(net4569),
    .A1(net2442),
    .Y(_09027_),
    .A2(net5095));
 sg13g2_a21oi_1 _17810_ (.A1(_09025_),
    .A2(_09027_),
    .Y(_00908_),
    .B1(net5534));
 sg13g2_nand2_1 _17811_ (.Y(_09028_),
    .A(\TRNG.Padded_Out[76] ),
    .B(net5148));
 sg13g2_a22oi_1 _17812_ (.Y(_09029_),
    .B1(net5133),
    .B2(\TRNG.Padded_Out[108] ),
    .A2(net5143),
    .A1(\TRNG.Padded_Out[364] ));
 sg13g2_a22oi_1 _17813_ (.Y(_09030_),
    .B1(net5129),
    .B2(\TRNG.Padded_Out[300] ),
    .A2(net5026),
    .A1(\TRNG.Padded_Out[140] ));
 sg13g2_a22oi_1 _17814_ (.Y(_09031_),
    .B1(net5021),
    .B2(\TRNG.Padded_Out[268] ),
    .A2(net5153),
    .A1(\TRNG.Padded_Out[332] ));
 sg13g2_a22oi_1 _17815_ (.Y(_09032_),
    .B1(net5124),
    .B2(\TRNG.Padded_Out[460] ),
    .A2(net5012),
    .A1(\TRNG.Padded_Out[396] ));
 sg13g2_a22oi_1 _17816_ (.Y(_09033_),
    .B1(net5001),
    .B2(\TRNG.Padded_Out[204] ),
    .A2(net5138),
    .A1(\TRNG.Padded_Out[428] ));
 sg13g2_nand3_1 _17817_ (.B(_09032_),
    .C(_09033_),
    .A(_09028_),
    .Y(_09034_));
 sg13g2_a221oi_1 _17818_ (.B2(\TRNG.Padded_Out[172] ),
    .C1(_09034_),
    .B1(net5007),
    .A1(\TRNG.Padded_Out[236] ),
    .Y(_09035_),
    .A2(net5016));
 sg13g2_nand4_1 _17819_ (.B(_09030_),
    .C(_09031_),
    .A(_09029_),
    .Y(_09036_),
    .D(_09035_));
 sg13g2_a21oi_1 _17820_ (.A1(net2342),
    .A2(net5155),
    .Y(_09037_),
    .B1(_09036_));
 sg13g2_a22oi_1 _17821_ (.Y(_09038_),
    .B1(net4569),
    .B2(net3300),
    .A2(net5095),
    .A1(net2441));
 sg13g2_a21oi_1 _17822_ (.A1(_09037_),
    .A2(_09038_),
    .Y(_00909_),
    .B1(net5534));
 sg13g2_nand2_1 _17823_ (.Y(_09039_),
    .A(\TRNG.Padded_Out[173] ),
    .B(net5006));
 sg13g2_a22oi_1 _17824_ (.Y(_09040_),
    .B1(net5133),
    .B2(\TRNG.Padded_Out[109] ),
    .A2(net5026),
    .A1(net1247));
 sg13g2_a22oi_1 _17825_ (.Y(_09041_),
    .B1(net5138),
    .B2(\TRNG.Padded_Out[429] ),
    .A2(net5143),
    .A1(\TRNG.Padded_Out[365] ));
 sg13g2_a22oi_1 _17826_ (.Y(_09042_),
    .B1(net5001),
    .B2(\TRNG.Padded_Out[205] ),
    .A2(net5129),
    .A1(\TRNG.Padded_Out[301] ));
 sg13g2_a22oi_1 _17827_ (.Y(_09043_),
    .B1(net5148),
    .B2(\TRNG.Padded_Out[77] ),
    .A2(net5153),
    .A1(\TRNG.Padded_Out[333] ));
 sg13g2_a22oi_1 _17828_ (.Y(_09044_),
    .B1(net5122),
    .B2(\TRNG.Padded_Out[461] ),
    .A2(net5018),
    .A1(\TRNG.Padded_Out[269] ));
 sg13g2_nand3_1 _17829_ (.B(_09043_),
    .C(_09044_),
    .A(_09039_),
    .Y(_09045_));
 sg13g2_a221oi_1 _17830_ (.B2(\TRNG.Padded_Out[397] ),
    .C1(_09045_),
    .B1(net5011),
    .A1(\TRNG.Padded_Out[237] ),
    .Y(_09046_),
    .A2(net5016));
 sg13g2_nand4_1 _17831_ (.B(_09041_),
    .C(_09042_),
    .A(_09040_),
    .Y(_09047_),
    .D(_09046_));
 sg13g2_a21oi_1 _17832_ (.A1(net2229),
    .A2(net5158),
    .Y(_09048_),
    .B1(_09047_));
 sg13g2_a22oi_1 _17833_ (.Y(_09049_),
    .B1(net4568),
    .B2(net3094),
    .A2(net5095),
    .A1(net2293));
 sg13g2_a21oi_1 _17834_ (.A1(_09048_),
    .A2(_09049_),
    .Y(_00910_),
    .B1(net5531));
 sg13g2_nand2_1 _17835_ (.Y(_09050_),
    .A(\TRNG.Padded_Out[270] ),
    .B(net5018));
 sg13g2_a22oi_1 _17836_ (.Y(_09051_),
    .B1(net5000),
    .B2(net1826),
    .A2(net5153),
    .A1(\TRNG.Padded_Out[334] ));
 sg13g2_a22oi_1 _17837_ (.Y(_09052_),
    .B1(net5129),
    .B2(\TRNG.Padded_Out[302] ),
    .A2(net5133),
    .A1(\TRNG.Padded_Out[110] ));
 sg13g2_a22oi_1 _17838_ (.Y(_09053_),
    .B1(net5138),
    .B2(\TRNG.Padded_Out[430] ),
    .A2(net5011),
    .A1(\TRNG.Padded_Out[398] ));
 sg13g2_a22oi_1 _17839_ (.Y(_09054_),
    .B1(net5147),
    .B2(\TRNG.Padded_Out[78] ),
    .A2(net5025),
    .A1(\TRNG.Padded_Out[142] ));
 sg13g2_a22oi_1 _17840_ (.Y(_09055_),
    .B1(net5120),
    .B2(\TRNG.Padded_Out[462] ),
    .A2(net5015),
    .A1(\TRNG.Padded_Out[238] ));
 sg13g2_nand3_1 _17841_ (.B(_09054_),
    .C(_09055_),
    .A(_09050_),
    .Y(_09056_));
 sg13g2_a221oi_1 _17842_ (.B2(\TRNG.Padded_Out[174] ),
    .C1(_09056_),
    .B1(net5005),
    .A1(\TRNG.Padded_Out[366] ),
    .Y(_09057_),
    .A2(net5142));
 sg13g2_nand4_1 _17843_ (.B(_09052_),
    .C(_09053_),
    .A(_09051_),
    .Y(_09058_),
    .D(_09057_));
 sg13g2_a22oi_1 _17844_ (.Y(_09059_),
    .B1(net5155),
    .B2(net2467),
    .A2(net5095),
    .A1(net2472));
 sg13g2_a21oi_1 _17845_ (.A1(net2636),
    .A2(net4568),
    .Y(_09060_),
    .B1(_09058_));
 sg13g2_a21oi_1 _17846_ (.A1(_09059_),
    .A2(_09060_),
    .Y(_00911_),
    .B1(net5533));
 sg13g2_and2_1 _17847_ (.A(\TRNG.Padded_Out[335] ),
    .B(net5152),
    .X(_09061_));
 sg13g2_a22oi_1 _17848_ (.Y(_09062_),
    .B1(net5123),
    .B2(\TRNG.Padded_Out[463] ),
    .A2(net5132),
    .A1(\TRNG.Padded_Out[111] ));
 sg13g2_a22oi_1 _17849_ (.Y(_09063_),
    .B1(net5005),
    .B2(\TRNG.Padded_Out[175] ),
    .A2(net5147),
    .A1(\TRNG.Padded_Out[79] ));
 sg13g2_a22oi_1 _17850_ (.Y(_09064_),
    .B1(net5137),
    .B2(\TRNG.Padded_Out[431] ),
    .A2(net5142),
    .A1(\TRNG.Padded_Out[367] ));
 sg13g2_nand2_1 _17851_ (.Y(_09065_),
    .A(_09063_),
    .B(_09064_));
 sg13g2_a221oi_1 _17852_ (.B2(\TRNG.Padded_Out[303] ),
    .C1(_09065_),
    .B1(net5128),
    .A1(\TRNG.Padded_Out[399] ),
    .Y(_09066_),
    .A2(net5009));
 sg13g2_a221oi_1 _17853_ (.B2(\TRNG.Padded_Out[271] ),
    .C1(_09061_),
    .B1(net5020),
    .A1(\TRNG.Padded_Out[143] ),
    .Y(_09067_),
    .A2(net5025));
 sg13g2_a22oi_1 _17854_ (.Y(_09068_),
    .B1(net5000),
    .B2(\TRNG.Padded_Out[207] ),
    .A2(net5015),
    .A1(\TRNG.Padded_Out[239] ));
 sg13g2_nand4_1 _17855_ (.B(_09066_),
    .C(_09067_),
    .A(_09062_),
    .Y(_09069_),
    .D(_09068_));
 sg13g2_a21oi_1 _17856_ (.A1(net2476),
    .A2(net5155),
    .Y(_09070_),
    .B1(_09069_));
 sg13g2_a22oi_1 _17857_ (.Y(_09071_),
    .B1(net4568),
    .B2(net3442),
    .A2(net5095),
    .A1(net2666));
 sg13g2_a21oi_1 _17858_ (.A1(_09070_),
    .A2(_09071_),
    .Y(_00912_),
    .B1(net5531));
 sg13g2_a22oi_1 _17859_ (.Y(_09072_),
    .B1(net5123),
    .B2(\TRNG.Padded_Out[464] ),
    .A2(net5005),
    .A1(\TRNG.Padded_Out[176] ));
 sg13g2_nand2_1 _17860_ (.Y(_09073_),
    .A(net1547),
    .B(net5137));
 sg13g2_a22oi_1 _17861_ (.Y(_09074_),
    .B1(net5001),
    .B2(\TRNG.Padded_Out[208] ),
    .A2(net5132),
    .A1(\TRNG.Padded_Out[112] ));
 sg13g2_a22oi_1 _17862_ (.Y(_09075_),
    .B1(net5128),
    .B2(\TRNG.Padded_Out[304] ),
    .A2(net5025),
    .A1(\TRNG.Padded_Out[144] ));
 sg13g2_a22oi_1 _17863_ (.Y(_09076_),
    .B1(net5142),
    .B2(\TRNG.Padded_Out[368] ),
    .A2(net5152),
    .A1(\TRNG.Padded_Out[336] ));
 sg13g2_nand3_1 _17864_ (.B(_09074_),
    .C(_09076_),
    .A(_09072_),
    .Y(_09077_));
 sg13g2_a22oi_1 _17865_ (.Y(_09078_),
    .B1(net5009),
    .B2(\TRNG.Padded_Out[400] ),
    .A2(net5016),
    .A1(\TRNG.Padded_Out[240] ));
 sg13g2_a22oi_1 _17866_ (.Y(_09079_),
    .B1(net5147),
    .B2(\TRNG.Padded_Out[80] ),
    .A2(net5020),
    .A1(\TRNG.Padded_Out[272] ));
 sg13g2_nand4_1 _17867_ (.B(_09075_),
    .C(_09078_),
    .A(_09073_),
    .Y(_09080_),
    .D(_09079_));
 sg13g2_nor2_2 _17868_ (.A(_09077_),
    .B(_09080_),
    .Y(_09081_));
 sg13g2_nor3_1 _17869_ (.A(_04255_),
    .B(net5343),
    .C(net5341),
    .Y(_09082_));
 sg13g2_a221oi_1 _17870_ (.B2(\TRNG.sha256.W[16] ),
    .C1(_09082_),
    .B1(net4568),
    .A1(net2511),
    .Y(_09083_),
    .A2(net5091));
 sg13g2_a21oi_1 _17871_ (.A1(_09081_),
    .A2(_09083_),
    .Y(_00913_),
    .B1(net5531));
 sg13g2_nand2_1 _17872_ (.Y(_09084_),
    .A(net1840),
    .B(net5015));
 sg13g2_a22oi_1 _17873_ (.Y(_09085_),
    .B1(net5000),
    .B2(net3797),
    .A2(net5025),
    .A1(\TRNG.Padded_Out[145] ));
 sg13g2_a22oi_1 _17874_ (.Y(_09086_),
    .B1(net5143),
    .B2(\TRNG.Padded_Out[369] ),
    .A2(net5147),
    .A1(\TRNG.Padded_Out[81] ));
 sg13g2_a22oi_1 _17875_ (.Y(_09087_),
    .B1(net5128),
    .B2(\TRNG.Padded_Out[305] ),
    .A2(net5137),
    .A1(\TRNG.Padded_Out[433] ));
 sg13g2_a22oi_1 _17876_ (.Y(_09088_),
    .B1(net5123),
    .B2(\TRNG.Padded_Out[465] ),
    .A2(net5020),
    .A1(\TRNG.Padded_Out[273] ));
 sg13g2_a22oi_1 _17877_ (.Y(_09089_),
    .B1(net5009),
    .B2(\TRNG.Padded_Out[401] ),
    .A2(net5152),
    .A1(\TRNG.Padded_Out[337] ));
 sg13g2_nand3_1 _17878_ (.B(_09088_),
    .C(_09089_),
    .A(_09087_),
    .Y(_09090_));
 sg13g2_a22oi_1 _17879_ (.Y(_09091_),
    .B1(net5132),
    .B2(\TRNG.Padded_Out[113] ),
    .A2(net5006),
    .A1(\TRNG.Padded_Out[177] ));
 sg13g2_nand4_1 _17880_ (.B(_09085_),
    .C(_09086_),
    .A(_09084_),
    .Y(_09092_),
    .D(_09091_));
 sg13g2_nor2_2 _17881_ (.A(_09090_),
    .B(_09092_),
    .Y(_09093_));
 sg13g2_nor3_1 _17882_ (.A(_04254_),
    .B(net5343),
    .C(net5341),
    .Y(_09094_));
 sg13g2_a221oi_1 _17883_ (.B2(\TRNG.sha256.W[17] ),
    .C1(_09094_),
    .B1(net4567),
    .A1(net2733),
    .Y(_09095_),
    .A2(net5092));
 sg13g2_a21oi_1 _17884_ (.A1(_09093_),
    .A2(_09095_),
    .Y(_00914_),
    .B1(net5531));
 sg13g2_nand2_1 _17885_ (.Y(_09096_),
    .A(\TRNG.Padded_Out[402] ),
    .B(net5009));
 sg13g2_a22oi_1 _17886_ (.Y(_09097_),
    .B1(net5128),
    .B2(\TRNG.Padded_Out[306] ),
    .A2(net5015),
    .A1(\TRNG.Padded_Out[242] ));
 sg13g2_a22oi_1 _17887_ (.Y(_09098_),
    .B1(net5000),
    .B2(\TRNG.Padded_Out[210] ),
    .A2(net5025),
    .A1(\TRNG.Padded_Out[146] ));
 sg13g2_a22oi_1 _17888_ (.Y(_09099_),
    .B1(net5123),
    .B2(\TRNG.Padded_Out[466] ),
    .A2(net5132),
    .A1(\TRNG.Padded_Out[114] ));
 sg13g2_a22oi_1 _17889_ (.Y(_09100_),
    .B1(net5142),
    .B2(\TRNG.Padded_Out[370] ),
    .A2(net5152),
    .A1(\TRNG.Padded_Out[338] ));
 sg13g2_a22oi_1 _17890_ (.Y(_09101_),
    .B1(net5005),
    .B2(\TRNG.Padded_Out[178] ),
    .A2(net5149),
    .A1(\TRNG.Padded_Out[82] ));
 sg13g2_nand3_1 _17891_ (.B(_09100_),
    .C(_09101_),
    .A(_09096_),
    .Y(_09102_));
 sg13g2_a221oi_1 _17892_ (.B2(\TRNG.Padded_Out[434] ),
    .C1(_09102_),
    .B1(net5137),
    .A1(\TRNG.Padded_Out[274] ),
    .Y(_09103_),
    .A2(net5020));
 sg13g2_nand4_1 _17893_ (.B(_09098_),
    .C(_09099_),
    .A(_09097_),
    .Y(_09104_),
    .D(_09103_));
 sg13g2_a21oi_1 _17894_ (.A1(net2269),
    .A2(net5155),
    .Y(_09105_),
    .B1(_09104_));
 sg13g2_a22oi_1 _17895_ (.Y(_09106_),
    .B1(net4567),
    .B2(net3347),
    .A2(net5092),
    .A1(net2526));
 sg13g2_a21oi_1 _17896_ (.A1(_09105_),
    .A2(_09106_),
    .Y(_00915_),
    .B1(net5531));
 sg13g2_a22oi_1 _17897_ (.Y(_09107_),
    .B1(net5152),
    .B2(\TRNG.Padded_Out[339] ),
    .A2(net5025),
    .A1(\TRNG.Padded_Out[147] ));
 sg13g2_nand2_1 _17898_ (.Y(_09108_),
    .A(\TRNG.Padded_Out[403] ),
    .B(net5009));
 sg13g2_a22oi_1 _17899_ (.Y(_09109_),
    .B1(net5123),
    .B2(\TRNG.Padded_Out[467] ),
    .A2(net5128),
    .A1(\TRNG.Padded_Out[307] ));
 sg13g2_a22oi_1 _17900_ (.Y(_09110_),
    .B1(net5005),
    .B2(\TRNG.Padded_Out[179] ),
    .A2(net5020),
    .A1(\TRNG.Padded_Out[275] ));
 sg13g2_a22oi_1 _17901_ (.Y(_09111_),
    .B1(net5000),
    .B2(\TRNG.Padded_Out[211] ),
    .A2(net5137),
    .A1(\TRNG.Padded_Out[435] ));
 sg13g2_a22oi_1 _17902_ (.Y(_09112_),
    .B1(net5015),
    .B2(\TRNG.Padded_Out[243] ),
    .A2(net5142),
    .A1(\TRNG.Padded_Out[371] ));
 sg13g2_nand3_1 _17903_ (.B(_09111_),
    .C(_09112_),
    .A(_09109_),
    .Y(_09113_));
 sg13g2_a22oi_1 _17904_ (.Y(_09114_),
    .B1(net5132),
    .B2(\TRNG.Padded_Out[115] ),
    .A2(net5147),
    .A1(\TRNG.Padded_Out[83] ));
 sg13g2_nand4_1 _17905_ (.B(_09108_),
    .C(_09110_),
    .A(_09107_),
    .Y(_09115_),
    .D(_09114_));
 sg13g2_nor2_2 _17906_ (.A(_09113_),
    .B(_09115_),
    .Y(_09116_));
 sg13g2_nor3_1 _17907_ (.A(_04252_),
    .B(net5343),
    .C(net5341),
    .Y(_09117_));
 sg13g2_a221oi_1 _17908_ (.B2(\TRNG.sha256.W[19] ),
    .C1(_09117_),
    .B1(net4567),
    .A1(net2685),
    .Y(_09118_),
    .A2(net5091));
 sg13g2_a21oi_1 _17909_ (.A1(_09116_),
    .A2(_09118_),
    .Y(_00916_),
    .B1(net5530));
 sg13g2_a22oi_1 _17910_ (.Y(_09119_),
    .B1(net5123),
    .B2(\TRNG.Padded_Out[468] ),
    .A2(net5137),
    .A1(\TRNG.Padded_Out[436] ));
 sg13g2_a22oi_1 _17911_ (.Y(_09120_),
    .B1(net5009),
    .B2(\TRNG.Padded_Out[404] ),
    .A2(net5152),
    .A1(\TRNG.Padded_Out[340] ));
 sg13g2_a22oi_1 _17912_ (.Y(_09121_),
    .B1(net5128),
    .B2(\TRNG.Padded_Out[308] ),
    .A2(net5020),
    .A1(\TRNG.Padded_Out[276] ));
 sg13g2_nand3_1 _17913_ (.B(_09120_),
    .C(_09121_),
    .A(_09119_),
    .Y(_09122_));
 sg13g2_nand2_1 _17914_ (.Y(_09123_),
    .A(\TRNG.Padded_Out[148] ),
    .B(net5026));
 sg13g2_a22oi_1 _17915_ (.Y(_09124_),
    .B1(net5000),
    .B2(\TRNG.Padded_Out[212] ),
    .A2(net5005),
    .A1(\TRNG.Padded_Out[180] ));
 sg13g2_a22oi_1 _17916_ (.Y(_09125_),
    .B1(net5015),
    .B2(\TRNG.Padded_Out[244] ),
    .A2(net5147),
    .A1(\TRNG.Padded_Out[84] ));
 sg13g2_a22oi_1 _17917_ (.Y(_09126_),
    .B1(net5132),
    .B2(\TRNG.Padded_Out[116] ),
    .A2(net5142),
    .A1(\TRNG.Padded_Out[372] ));
 sg13g2_nand4_1 _17918_ (.B(_09124_),
    .C(_09125_),
    .A(_09123_),
    .Y(_09127_),
    .D(_09126_));
 sg13g2_nor2_2 _17919_ (.A(_09122_),
    .B(_09127_),
    .Y(_09128_));
 sg13g2_a22oi_1 _17920_ (.Y(_09129_),
    .B1(net5155),
    .B2(net1886),
    .A2(net5092),
    .A1(net3356));
 sg13g2_nand2_2 _17921_ (.Y(_09130_),
    .A(_09128_),
    .B(_09129_));
 sg13g2_a21oi_1 _17922_ (.A1(net3819),
    .A2(net4569),
    .Y(_09131_),
    .B1(_09130_));
 sg13g2_nor2_1 _17923_ (.A(net5543),
    .B(_09131_),
    .Y(_00917_));
 sg13g2_nand2_1 _17924_ (.Y(_09132_),
    .A(\TRNG.Padded_Out[341] ),
    .B(net5152));
 sg13g2_a22oi_1 _17925_ (.Y(_09133_),
    .B1(net5005),
    .B2(net3811),
    .A2(net5025),
    .A1(\TRNG.Padded_Out[149] ));
 sg13g2_a22oi_1 _17926_ (.Y(_09134_),
    .B1(net5137),
    .B2(\TRNG.Padded_Out[437] ),
    .A2(net5015),
    .A1(\TRNG.Padded_Out[245] ));
 sg13g2_a22oi_1 _17927_ (.Y(_09135_),
    .B1(net5123),
    .B2(\TRNG.Padded_Out[469] ),
    .A2(net5147),
    .A1(\TRNG.Padded_Out[85] ));
 sg13g2_a22oi_1 _17928_ (.Y(_09136_),
    .B1(net5132),
    .B2(\TRNG.Padded_Out[117] ),
    .A2(net5020),
    .A1(\TRNG.Padded_Out[277] ));
 sg13g2_nand3_1 _17929_ (.B(_09135_),
    .C(_09136_),
    .A(_09133_),
    .Y(_09137_));
 sg13g2_a22oi_1 _17930_ (.Y(_09138_),
    .B1(net5000),
    .B2(\TRNG.Padded_Out[213] ),
    .A2(net5128),
    .A1(\TRNG.Padded_Out[309] ));
 sg13g2_a22oi_1 _17931_ (.Y(_09139_),
    .B1(net5008),
    .B2(\TRNG.Padded_Out[405] ),
    .A2(net5142),
    .A1(\TRNG.Padded_Out[373] ));
 sg13g2_nand4_1 _17932_ (.B(_09134_),
    .C(_09138_),
    .A(_09132_),
    .Y(_09140_),
    .D(_09139_));
 sg13g2_nor2_2 _17933_ (.A(net3812),
    .B(_09140_),
    .Y(_09141_));
 sg13g2_nor3_1 _17934_ (.A(_04250_),
    .B(net5343),
    .C(net5341),
    .Y(_09142_));
 sg13g2_a221oi_1 _17935_ (.B2(\TRNG.sha256.W[21] ),
    .C1(_09142_),
    .B1(net4567),
    .A1(net2997),
    .Y(_09143_),
    .A2(net5091));
 sg13g2_a21oi_1 _17936_ (.A1(_09141_),
    .A2(_09143_),
    .Y(_00918_),
    .B1(net5529));
 sg13g2_a22oi_1 _17937_ (.Y(_09144_),
    .B1(net5000),
    .B2(\TRNG.Padded_Out[214] ),
    .A2(net5020),
    .A1(\TRNG.Padded_Out[278] ));
 sg13g2_nand2_1 _17938_ (.Y(_09145_),
    .A(\TRNG.Padded_Out[438] ),
    .B(net5137));
 sg13g2_a22oi_1 _17939_ (.Y(_09146_),
    .B1(net5125),
    .B2(\TRNG.Padded_Out[310] ),
    .A2(net5025),
    .A1(\TRNG.Padded_Out[150] ));
 sg13g2_a22oi_1 _17940_ (.Y(_09147_),
    .B1(net5132),
    .B2(\TRNG.Padded_Out[118] ),
    .A2(net5005),
    .A1(\TRNG.Padded_Out[182] ));
 sg13g2_a22oi_1 _17941_ (.Y(_09148_),
    .B1(net5009),
    .B2(\TRNG.Padded_Out[406] ),
    .A2(net5152),
    .A1(\TRNG.Padded_Out[342] ));
 sg13g2_a22oi_1 _17942_ (.Y(_09149_),
    .B1(net5122),
    .B2(\TRNG.Padded_Out[470] ),
    .A2(net5147),
    .A1(\TRNG.Padded_Out[86] ));
 sg13g2_nand3_1 _17943_ (.B(_09148_),
    .C(_09149_),
    .A(_09145_),
    .Y(_09150_));
 sg13g2_a221oi_1 _17944_ (.B2(\TRNG.Padded_Out[246] ),
    .C1(_09150_),
    .B1(net5015),
    .A1(\TRNG.Padded_Out[374] ),
    .Y(_09151_),
    .A2(net5142));
 sg13g2_nand4_1 _17945_ (.B(_09146_),
    .C(_09147_),
    .A(_09144_),
    .Y(_09152_),
    .D(_09151_));
 sg13g2_a21oi_1 _17946_ (.A1(net1853),
    .A2(net5155),
    .Y(_09153_),
    .B1(_09152_));
 sg13g2_a22oi_1 _17947_ (.Y(_09154_),
    .B1(net4567),
    .B2(\TRNG.sha256.W[22] ),
    .A2(net5091),
    .A1(net2700));
 sg13g2_a21oi_1 _17948_ (.A1(_09153_),
    .A2(_09154_),
    .Y(_00919_),
    .B1(net5532));
 sg13g2_a22oi_1 _17949_ (.Y(_09155_),
    .B1(net5003),
    .B2(\TRNG.Padded_Out[183] ),
    .A2(net5145),
    .A1(\TRNG.Padded_Out[87] ));
 sg13g2_nand2_1 _17950_ (.Y(_09156_),
    .A(\TRNG.Padded_Out[439] ),
    .B(net5136));
 sg13g2_a22oi_1 _17951_ (.Y(_09157_),
    .B1(net5008),
    .B2(\TRNG.Padded_Out[407] ),
    .A2(net5151),
    .A1(\TRNG.Padded_Out[343] ));
 sg13g2_a22oi_1 _17952_ (.Y(_09158_),
    .B1(net4999),
    .B2(net1965),
    .A2(net5019),
    .A1(\TRNG.Padded_Out[279] ));
 sg13g2_a22oi_1 _17953_ (.Y(_09159_),
    .B1(net5130),
    .B2(\TRNG.Padded_Out[119] ),
    .A2(net5013),
    .A1(\TRNG.Padded_Out[247] ));
 sg13g2_a22oi_1 _17954_ (.Y(_09160_),
    .B1(net5120),
    .B2(\TRNG.Padded_Out[471] ),
    .A2(net5140),
    .A1(\TRNG.Padded_Out[375] ));
 sg13g2_a22oi_1 _17955_ (.Y(_09161_),
    .B1(net5127),
    .B2(net1966),
    .A2(net5024),
    .A1(net3664));
 sg13g2_nand3_1 _17956_ (.B(_09160_),
    .C(_09161_),
    .A(_09158_),
    .Y(_09162_));
 sg13g2_nand4_1 _17957_ (.B(_09156_),
    .C(_09157_),
    .A(_09155_),
    .Y(_09163_),
    .D(_09159_));
 sg13g2_nor2_2 _17958_ (.A(_09162_),
    .B(_09163_),
    .Y(_09164_));
 sg13g2_nor3_1 _17959_ (.A(_04248_),
    .B(net5343),
    .C(net5341),
    .Y(_09165_));
 sg13g2_a221oi_1 _17960_ (.B2(\TRNG.sha256.W[23] ),
    .C1(_09165_),
    .B1(net4567),
    .A1(net2464),
    .Y(_09166_),
    .A2(net5091));
 sg13g2_a21oi_1 _17961_ (.A1(_09164_),
    .A2(_09166_),
    .Y(_00920_),
    .B1(net5530));
 sg13g2_a22oi_1 _17962_ (.Y(_09167_),
    .B1(net5136),
    .B2(\TRNG.Padded_Out[440] ),
    .A2(net5013),
    .A1(\TRNG.Padded_Out[248] ));
 sg13g2_nand2_1 _17963_ (.Y(_09168_),
    .A(net3726),
    .B(net5023));
 sg13g2_a22oi_1 _17964_ (.Y(_09169_),
    .B1(net5122),
    .B2(\TRNG.Padded_Out[472] ),
    .A2(net5151),
    .A1(\TRNG.Padded_Out[344] ));
 sg13g2_a22oi_1 _17965_ (.Y(_09170_),
    .B1(net5125),
    .B2(net1908),
    .A2(net5130),
    .A1(\TRNG.Padded_Out[120] ));
 sg13g2_a22oi_1 _17966_ (.Y(_09171_),
    .B1(net5008),
    .B2(\TRNG.Padded_Out[408] ),
    .A2(net5145),
    .A1(\TRNG.Padded_Out[88] ));
 sg13g2_a22oi_1 _17967_ (.Y(_09172_),
    .B1(net5141),
    .B2(\TRNG.Padded_Out[376] ),
    .A2(net5019),
    .A1(\TRNG.Padded_Out[280] ));
 sg13g2_nand3_1 _17968_ (.B(_09170_),
    .C(_09172_),
    .A(_09169_),
    .Y(_09173_));
 sg13g2_a22oi_1 _17969_ (.Y(_09174_),
    .B1(net4999),
    .B2(\TRNG.Padded_Out[216] ),
    .A2(net5003),
    .A1(\TRNG.Padded_Out[184] ));
 sg13g2_nand4_1 _17970_ (.B(_09168_),
    .C(_09171_),
    .A(_09167_),
    .Y(_02168_),
    .D(_09174_));
 sg13g2_nor2_2 _17971_ (.A(_09173_),
    .B(_02168_),
    .Y(_02169_));
 sg13g2_nor3_1 _17972_ (.A(_04247_),
    .B(net5343),
    .C(net5341),
    .Y(_02170_));
 sg13g2_a221oi_1 _17973_ (.B2(\TRNG.sha256.W[24] ),
    .C1(_02170_),
    .B1(net4567),
    .A1(net2575),
    .Y(_02171_),
    .A2(net5091));
 sg13g2_a21oi_1 _17974_ (.A1(_02169_),
    .A2(_02171_),
    .Y(_00921_),
    .B1(net5532));
 sg13g2_nand2_1 _17975_ (.Y(_02172_),
    .A(\TRNG.Padded_Out[441] ),
    .B(net5136));
 sg13g2_a22oi_1 _17976_ (.Y(_02173_),
    .B1(net4999),
    .B2(\TRNG.Padded_Out[217] ),
    .A2(net5013),
    .A1(\TRNG.Padded_Out[249] ));
 sg13g2_a22oi_1 _17977_ (.Y(_02174_),
    .B1(net5125),
    .B2(\TRNG.Padded_Out[313] ),
    .A2(net5023),
    .A1(\TRNG.Padded_Out[153] ));
 sg13g2_a22oi_1 _17978_ (.Y(_02175_),
    .B1(net5120),
    .B2(\TRNG.Padded_Out[473] ),
    .A2(net5003),
    .A1(\TRNG.Padded_Out[185] ));
 sg13g2_a22oi_1 _17979_ (.Y(_02176_),
    .B1(net5145),
    .B2(\TRNG.Padded_Out[89] ),
    .A2(net5018),
    .A1(\TRNG.Padded_Out[281] ));
 sg13g2_a22oi_1 _17980_ (.Y(_02177_),
    .B1(net5140),
    .B2(\TRNG.Padded_Out[377] ),
    .A2(net5151),
    .A1(\TRNG.Padded_Out[345] ));
 sg13g2_a22oi_1 _17981_ (.Y(_02178_),
    .B1(net5130),
    .B2(\TRNG.Padded_Out[121] ),
    .A2(net5008),
    .A1(\TRNG.Padded_Out[409] ));
 sg13g2_nand3_1 _17982_ (.B(_02177_),
    .C(_02178_),
    .A(_02173_),
    .Y(_02179_));
 sg13g2_nand4_1 _17983_ (.B(_02174_),
    .C(_02175_),
    .A(_02172_),
    .Y(_02180_),
    .D(_02176_));
 sg13g2_nor2_2 _17984_ (.A(_02179_),
    .B(_02180_),
    .Y(_02181_));
 sg13g2_nand2_1 _17985_ (.Y(_02182_),
    .A(net2623),
    .B(net5155));
 sg13g2_and2_1 _17986_ (.A(_02181_),
    .B(_02182_),
    .X(_02183_));
 sg13g2_a22oi_1 _17987_ (.Y(_02184_),
    .B1(net4568),
    .B2(net3426),
    .A2(net5095),
    .A1(net2378));
 sg13g2_a21oi_1 _17988_ (.A1(_02183_),
    .A2(_02184_),
    .Y(_00922_),
    .B1(net5532));
 sg13g2_a22oi_1 _17989_ (.Y(_02185_),
    .B1(net5120),
    .B2(\TRNG.Padded_Out[474] ),
    .A2(net5151),
    .A1(\TRNG.Padded_Out[346] ));
 sg13g2_a22oi_1 _17990_ (.Y(_02186_),
    .B1(net5003),
    .B2(\TRNG.Padded_Out[186] ),
    .A2(net5008),
    .A1(\TRNG.Padded_Out[410] ));
 sg13g2_a22oi_1 _17991_ (.Y(_02187_),
    .B1(net5125),
    .B2(\TRNG.Padded_Out[314] ),
    .A2(net5140),
    .A1(\TRNG.Padded_Out[378] ));
 sg13g2_nand3_1 _17992_ (.B(_02186_),
    .C(_02187_),
    .A(_02185_),
    .Y(_02188_));
 sg13g2_nand2_1 _17993_ (.Y(_02189_),
    .A(\TRNG.Padded_Out[154] ),
    .B(net5023));
 sg13g2_a22oi_1 _17994_ (.Y(_02190_),
    .B1(net5013),
    .B2(\TRNG.Padded_Out[250] ),
    .A2(net5145),
    .A1(\TRNG.Padded_Out[90] ));
 sg13g2_a22oi_1 _17995_ (.Y(_02191_),
    .B1(net5130),
    .B2(\TRNG.Padded_Out[122] ),
    .A2(net5136),
    .A1(\TRNG.Padded_Out[442] ));
 sg13g2_a22oi_1 _17996_ (.Y(_02192_),
    .B1(net4999),
    .B2(\TRNG.Padded_Out[218] ),
    .A2(net5018),
    .A1(\TRNG.Padded_Out[282] ));
 sg13g2_nand4_1 _17997_ (.B(_02190_),
    .C(_02191_),
    .A(_02189_),
    .Y(_02193_),
    .D(_02192_));
 sg13g2_nor2_2 _17998_ (.A(_02188_),
    .B(_02193_),
    .Y(_02194_));
 sg13g2_nor3_1 _17999_ (.A(_04245_),
    .B(net5344),
    .C(net5342),
    .Y(_02195_));
 sg13g2_a221oi_1 _18000_ (.B2(\TRNG.sha256.W[26] ),
    .C1(_02195_),
    .B1(net4569),
    .A1(net2580),
    .Y(_02196_),
    .A2(net5095));
 sg13g2_a21oi_1 _18001_ (.A1(_02194_),
    .A2(_02196_),
    .Y(_00923_),
    .B1(net5542));
 sg13g2_a22oi_1 _18002_ (.Y(_02197_),
    .B1(net5003),
    .B2(\TRNG.Padded_Out[187] ),
    .A2(net5140),
    .A1(\TRNG.Padded_Out[379] ));
 sg13g2_nand2_1 _18003_ (.Y(_02198_),
    .A(\TRNG.Padded_Out[91] ),
    .B(net5145));
 sg13g2_a22oi_1 _18004_ (.Y(_02199_),
    .B1(net4999),
    .B2(\TRNG.Padded_Out[219] ),
    .A2(net5008),
    .A1(\TRNG.Padded_Out[411] ));
 sg13g2_a22oi_1 _18005_ (.Y(_02200_),
    .B1(net5013),
    .B2(\TRNG.Padded_Out[251] ),
    .A2(net5018),
    .A1(\TRNG.Padded_Out[283] ));
 sg13g2_a22oi_1 _18006_ (.Y(_02201_),
    .B1(net5120),
    .B2(\TRNG.Padded_Out[475] ),
    .A2(net5125),
    .A1(\TRNG.Padded_Out[315] ));
 sg13g2_a22oi_1 _18007_ (.Y(_02202_),
    .B1(net5151),
    .B2(\TRNG.Padded_Out[347] ),
    .A2(net5023),
    .A1(\TRNG.Padded_Out[155] ));
 sg13g2_nand3_1 _18008_ (.B(_02198_),
    .C(_02202_),
    .A(_02197_),
    .Y(_02203_));
 sg13g2_a221oi_1 _18009_ (.B2(\TRNG.Padded_Out[123] ),
    .C1(_02203_),
    .B1(net5130),
    .A1(\TRNG.Padded_Out[443] ),
    .Y(_02204_),
    .A2(net5136));
 sg13g2_nand4_1 _18010_ (.B(_02200_),
    .C(_02201_),
    .A(_02199_),
    .Y(_02205_),
    .D(_02204_));
 sg13g2_a221oi_1 _18011_ (.B2(net4958),
    .C1(_02205_),
    .B1(net4959),
    .A1(net2134),
    .Y(_02206_),
    .A2(net5157));
 sg13g2_a21oi_1 _18012_ (.A1(_04336_),
    .A2(net5094),
    .Y(_02207_),
    .B1(net5542));
 sg13g2_o21ai_1 _18013_ (.B1(_02207_),
    .Y(_02208_),
    .A1(net3590),
    .A2(_08891_));
 sg13g2_nor2_1 _18014_ (.A(_02206_),
    .B(_02208_),
    .Y(_00924_));
 sg13g2_nand2_1 _18015_ (.Y(_02209_),
    .A(\TRNG.Padded_Out[380] ),
    .B(net5140));
 sg13g2_a22oi_1 _18016_ (.Y(_02210_),
    .B1(net5003),
    .B2(\TRNG.Padded_Out[188] ),
    .A2(net5023),
    .A1(\TRNG.Padded_Out[156] ));
 sg13g2_a22oi_1 _18017_ (.Y(_02211_),
    .B1(net5130),
    .B2(\TRNG.Padded_Out[124] ),
    .A2(net5018),
    .A1(\TRNG.Padded_Out[284] ));
 sg13g2_a22oi_1 _18018_ (.Y(_02212_),
    .B1(net5125),
    .B2(\TRNG.Padded_Out[316] ),
    .A2(net5008),
    .A1(\TRNG.Padded_Out[412] ));
 sg13g2_a22oi_1 _18019_ (.Y(_02213_),
    .B1(net5120),
    .B2(\TRNG.Padded_Out[476] ),
    .A2(net5013),
    .A1(\TRNG.Padded_Out[252] ));
 sg13g2_a22oi_1 _18020_ (.Y(_02214_),
    .B1(net5136),
    .B2(\TRNG.Padded_Out[444] ),
    .A2(net5151),
    .A1(\TRNG.Padded_Out[348] ));
 sg13g2_nand3_1 _18021_ (.B(_02213_),
    .C(_02214_),
    .A(_02209_),
    .Y(_02215_));
 sg13g2_a221oi_1 _18022_ (.B2(\TRNG.Padded_Out[220] ),
    .C1(_02215_),
    .B1(net4999),
    .A1(\TRNG.Padded_Out[92] ),
    .Y(_02216_),
    .A2(net5145));
 sg13g2_nand4_1 _18023_ (.B(_02211_),
    .C(_02212_),
    .A(_02210_),
    .Y(_02217_),
    .D(_02216_));
 sg13g2_a22oi_1 _18024_ (.Y(_02218_),
    .B1(net5157),
    .B2(net2271),
    .A2(net5094),
    .A1(net2364));
 sg13g2_a21oi_1 _18025_ (.A1(\TRNG.sha256.W[28] ),
    .A2(net4570),
    .Y(_02219_),
    .B1(_02217_));
 sg13g2_a21oi_1 _18026_ (.A1(_02218_),
    .A2(_02219_),
    .Y(_00925_),
    .B1(net5543));
 sg13g2_nand2_1 _18027_ (.Y(_02220_),
    .A(\TRNG.Padded_Out[125] ),
    .B(net5130));
 sg13g2_a22oi_1 _18028_ (.Y(_02221_),
    .B1(net5003),
    .B2(\TRNG.Padded_Out[189] ),
    .A2(net5023),
    .A1(\TRNG.Padded_Out[157] ));
 sg13g2_a22oi_1 _18029_ (.Y(_02222_),
    .B1(net5013),
    .B2(\TRNG.Padded_Out[253] ),
    .A2(net5018),
    .A1(\TRNG.Padded_Out[285] ));
 sg13g2_a22oi_1 _18030_ (.Y(_02223_),
    .B1(net4999),
    .B2(\TRNG.Padded_Out[221] ),
    .A2(net5008),
    .A1(\TRNG.Padded_Out[413] ));
 sg13g2_a22oi_1 _18031_ (.Y(_02224_),
    .B1(net5125),
    .B2(\TRNG.Padded_Out[317] ),
    .A2(net5140),
    .A1(\TRNG.Padded_Out[381] ));
 sg13g2_a22oi_1 _18032_ (.Y(_02225_),
    .B1(net5120),
    .B2(\TRNG.Padded_Out[477] ),
    .A2(net5145),
    .A1(\TRNG.Padded_Out[93] ));
 sg13g2_nand3_1 _18033_ (.B(_02221_),
    .C(_02225_),
    .A(_02220_),
    .Y(_02226_));
 sg13g2_a221oi_1 _18034_ (.B2(\TRNG.Padded_Out[445] ),
    .C1(_02226_),
    .B1(net5136),
    .A1(\TRNG.Padded_Out[349] ),
    .Y(_02227_),
    .A2(net5151));
 sg13g2_nand4_1 _18035_ (.B(_02223_),
    .C(_02224_),
    .A(_02222_),
    .Y(_02228_),
    .D(_02227_));
 sg13g2_a22oi_1 _18036_ (.Y(_02229_),
    .B1(net5157),
    .B2(net1931),
    .A2(net5093),
    .A1(net2357));
 sg13g2_a21oi_1 _18037_ (.A1(net2778),
    .A2(net4569),
    .Y(_02230_),
    .B1(_02228_));
 sg13g2_a21oi_1 _18038_ (.A1(_02229_),
    .A2(_02230_),
    .Y(_00926_),
    .B1(net5543));
 sg13g2_nand2_1 _18039_ (.Y(_02231_),
    .A(\TRNG.Padded_Out[350] ),
    .B(net5151));
 sg13g2_a22oi_1 _18040_ (.Y(_02232_),
    .B1(net5145),
    .B2(\TRNG.Padded_Out[94] ),
    .A2(net5018),
    .A1(\TRNG.Padded_Out[286] ));
 sg13g2_a22oi_1 _18041_ (.Y(_02233_),
    .B1(net5013),
    .B2(\TRNG.Padded_Out[254] ),
    .A2(net5140),
    .A1(\TRNG.Padded_Out[382] ));
 sg13g2_a22oi_1 _18042_ (.Y(_02234_),
    .B1(net5130),
    .B2(\TRNG.Padded_Out[126] ),
    .A2(net5136),
    .A1(\TRNG.Padded_Out[446] ));
 sg13g2_a22oi_1 _18043_ (.Y(_02235_),
    .B1(net5010),
    .B2(\TRNG.Padded_Out[414] ),
    .A2(net5023),
    .A1(\TRNG.Padded_Out[158] ));
 sg13g2_a22oi_1 _18044_ (.Y(_02236_),
    .B1(net4999),
    .B2(\TRNG.Padded_Out[222] ),
    .A2(net5125),
    .A1(\TRNG.Padded_Out[318] ));
 sg13g2_nand3_1 _18045_ (.B(_02235_),
    .C(_02236_),
    .A(_02231_),
    .Y(_02237_));
 sg13g2_a221oi_1 _18046_ (.B2(\TRNG.Padded_Out[478] ),
    .C1(_02237_),
    .B1(net5120),
    .A1(\TRNG.Padded_Out[190] ),
    .Y(_02238_),
    .A2(net5003));
 sg13g2_nand4_1 _18047_ (.B(_02233_),
    .C(_02234_),
    .A(_02232_),
    .Y(_02239_),
    .D(_02238_));
 sg13g2_a221oi_1 _18048_ (.B2(_08888_),
    .C1(_02239_),
    .B1(_08886_),
    .A1(net2512),
    .Y(_02240_),
    .A2(net5158));
 sg13g2_a21oi_1 _18049_ (.A1(_04339_),
    .A2(net5094),
    .Y(_02241_),
    .B1(net5540));
 sg13g2_o21ai_1 _18050_ (.B1(_02241_),
    .Y(_02242_),
    .A1(net3524),
    .A2(_08891_));
 sg13g2_nor2_1 _18051_ (.A(_02240_),
    .B(_02242_),
    .Y(_00927_));
 sg13g2_a22oi_1 _18052_ (.Y(_02243_),
    .B1(net5122),
    .B2(\TRNG.Padded_Out[479] ),
    .A2(net5140),
    .A1(\TRNG.Padded_Out[383] ));
 sg13g2_nand2_1 _18053_ (.Y(_02244_),
    .A(\TRNG.Padded_Out[415] ),
    .B(net5010));
 sg13g2_a22oi_1 _18054_ (.Y(_02245_),
    .B1(net4998),
    .B2(\TRNG.Padded_Out[223] ),
    .A2(net5004),
    .A1(\TRNG.Padded_Out[191] ));
 sg13g2_a22oi_1 _18055_ (.Y(_02246_),
    .B1(net5127),
    .B2(\TRNG.Padded_Out[319] ),
    .A2(net5150),
    .A1(\TRNG.Padded_Out[351] ));
 sg13g2_a22oi_1 _18056_ (.Y(_02247_),
    .B1(net5131),
    .B2(\TRNG.Padded_Out[127] ),
    .A2(net5014),
    .A1(\TRNG.Padded_Out[255] ));
 sg13g2_a22oi_1 _18057_ (.Y(_02248_),
    .B1(net5146),
    .B2(\TRNG.Padded_Out[95] ),
    .A2(net5023),
    .A1(\TRNG.Padded_Out[159] ));
 sg13g2_nand3_1 _18058_ (.B(_02244_),
    .C(_02248_),
    .A(_02243_),
    .Y(_02249_));
 sg13g2_a221oi_1 _18059_ (.B2(\TRNG.Padded_Out[447] ),
    .C1(_02249_),
    .B1(net5139),
    .A1(\TRNG.Padded_Out[287] ),
    .Y(_02250_),
    .A2(net5022));
 sg13g2_nand4_1 _18060_ (.B(_02246_),
    .C(_02247_),
    .A(_02245_),
    .Y(_02251_),
    .D(_02250_));
 sg13g2_a21oi_1 _18061_ (.A1(net2478),
    .A2(net5157),
    .Y(_02252_),
    .B1(_02251_));
 sg13g2_a22oi_1 _18062_ (.Y(_02253_),
    .B1(net4569),
    .B2(\TRNG.sha256.W[31] ),
    .A2(net5094),
    .A1(net3309));
 sg13g2_a21oi_1 _18063_ (.A1(_02252_),
    .A2(net3310),
    .Y(_00928_),
    .B1(net5540));
 sg13g2_a21oi_2 _18064_ (.B1(net5161),
    .Y(_02254_),
    .A2(_06867_),
    .A1(net5876));
 sg13g2_nor2b_2 _18065_ (.A(_08887_),
    .B_N(net4996),
    .Y(_02255_));
 sg13g2_nand2b_1 _18066_ (.Y(_02256_),
    .B(net4996),
    .A_N(_08887_));
 sg13g2_nand3_1 _18067_ (.B(net4958),
    .C(_02256_),
    .A(_08811_),
    .Y(_02257_));
 sg13g2_a21oi_1 _18068_ (.A1(net3807),
    .A2(net4565),
    .Y(_02258_),
    .B1(net5543));
 sg13g2_nand2_1 _18069_ (.Y(_00929_),
    .A(_02257_),
    .B(_02258_));
 sg13g2_nor2_1 _18070_ (.A(_06870_),
    .B(_08811_),
    .Y(_02259_));
 sg13g2_nor2_2 _18071_ (.A(_08811_),
    .B(net5342),
    .Y(_02260_));
 sg13g2_nor3_2 _18072_ (.A(_08887_),
    .B(net4987),
    .C(_02260_),
    .Y(_02261_));
 sg13g2_o21ai_1 _18073_ (.B1(_02261_),
    .Y(_02262_),
    .A1(_06868_),
    .A2(_08865_));
 sg13g2_nor2_2 _18074_ (.A(_08811_),
    .B(_08865_),
    .Y(_02263_));
 sg13g2_nor2_2 _18075_ (.A(_08811_),
    .B(_08836_),
    .Y(_02264_));
 sg13g2_nand2b_1 _18076_ (.Y(_02265_),
    .B(net4987),
    .A_N(_00270_));
 sg13g2_nor3_2 _18077_ (.A(net5153),
    .B(net5149),
    .C(net5001),
    .Y(_02266_));
 sg13g2_nand4_1 _18078_ (.B(_08872_),
    .C(_02265_),
    .A(_08808_),
    .Y(_02267_),
    .D(_02266_));
 sg13g2_a21oi_1 _18079_ (.A1(net3661),
    .A2(_02264_),
    .Y(_02268_),
    .B1(_02267_));
 sg13g2_o21ai_1 _18080_ (.B1(net5478),
    .Y(_02269_),
    .A1(\TRNG.sha256.expand.address1[0] ),
    .A2(_02262_));
 sg13g2_a21oi_1 _18081_ (.A1(_02262_),
    .A2(net3662),
    .Y(_00930_),
    .B1(_02269_));
 sg13g2_o21ai_1 _18082_ (.B1(_08807_),
    .Y(_02270_),
    .A1(\TRNG.sha256.compress.count[0] ),
    .A2(_08806_));
 sg13g2_o21ai_1 _18083_ (.B1(_02270_),
    .Y(_02271_),
    .A1(_08860_),
    .A2(_08865_));
 sg13g2_a221oi_1 _18084_ (.B2(net2494),
    .C1(_02271_),
    .B1(_02264_),
    .A1(net2655),
    .Y(_02272_),
    .A2(net4987));
 sg13g2_o21ai_1 _18085_ (.B1(net5478),
    .Y(_02273_),
    .A1(net3653),
    .A2(_02262_));
 sg13g2_a21oi_1 _18086_ (.A1(_02262_),
    .A2(_02272_),
    .Y(_00931_),
    .B1(_02273_));
 sg13g2_a221oi_1 _18087_ (.B2(net3459),
    .C1(net3651),
    .B1(_02264_),
    .A1(net3430),
    .Y(_02274_),
    .A2(net4987));
 sg13g2_o21ai_1 _18088_ (.B1(net5478),
    .Y(_02275_),
    .A1(\TRNG.sha256.expand.address1[2] ),
    .A2(_02262_));
 sg13g2_a21oi_1 _18089_ (.A1(_02262_),
    .A2(_02274_),
    .Y(_00932_),
    .B1(_02275_));
 sg13g2_a221oi_1 _18090_ (.B2(net3398),
    .C1(net3596),
    .B1(_02264_),
    .A1(net3450),
    .Y(_02276_),
    .A2(net4987));
 sg13g2_o21ai_1 _18091_ (.B1(net5478),
    .Y(_02277_),
    .A1(\TRNG.sha256.expand.address1[3] ),
    .A2(_02262_));
 sg13g2_a21oi_1 _18092_ (.A1(_02262_),
    .A2(_02276_),
    .Y(_00933_),
    .B1(_02277_));
 sg13g2_nand2_1 _18093_ (.Y(_02278_),
    .A(_04274_),
    .B(_02259_));
 sg13g2_a22oi_1 _18094_ (.Y(_02279_),
    .B1(_02261_),
    .B2(net5779),
    .A2(_02260_),
    .A1(net2311));
 sg13g2_a21oi_1 _18095_ (.A1(_02278_),
    .A2(_02279_),
    .Y(_00934_),
    .B1(net5538));
 sg13g2_nand2_1 _18096_ (.Y(_02280_),
    .A(net3386),
    .B(_02259_));
 sg13g2_a22oi_1 _18097_ (.Y(_02281_),
    .B1(_02261_),
    .B2(net5737),
    .A2(_02260_),
    .A1(net2388));
 sg13g2_a21oi_1 _18098_ (.A1(_02280_),
    .A2(_02281_),
    .Y(_00935_),
    .B1(net5538));
 sg13g2_nand2_1 _18099_ (.Y(_02282_),
    .A(net3285),
    .B(net4987));
 sg13g2_a22oi_1 _18100_ (.Y(_02283_),
    .B1(_02261_),
    .B2(net5706),
    .A2(_02260_),
    .A1(net2532));
 sg13g2_a21oi_1 _18101_ (.A1(_02282_),
    .A2(_02283_),
    .Y(_00936_),
    .B1(net5538));
 sg13g2_nand2_1 _18102_ (.Y(_02284_),
    .A(net2064),
    .B(net4987));
 sg13g2_a22oi_1 _18103_ (.Y(_02285_),
    .B1(_02261_),
    .B2(net5694),
    .A2(_02260_),
    .A1(net2289));
 sg13g2_a21oi_1 _18104_ (.A1(_02284_),
    .A2(_02285_),
    .Y(_00937_),
    .B1(net5538));
 sg13g2_nor3_1 _18105_ (.A(net5876),
    .B(_08806_),
    .C(_08865_),
    .Y(_02286_));
 sg13g2_or4_1 _18106_ (.A(net5161),
    .B(net5148),
    .C(net4987),
    .D(_02286_),
    .X(_02287_));
 sg13g2_nor3_1 _18107_ (.A(_08812_),
    .B(_08884_),
    .C(_02287_),
    .Y(_02288_));
 sg13g2_a21oi_1 _18108_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[0] ),
    .A2(net5159),
    .Y(_02289_),
    .B1(net4734));
 sg13g2_a221oi_1 _18109_ (.B2(_08882_),
    .C1(net4561),
    .B1(_02289_),
    .A1(_04309_),
    .Y(_02290_),
    .A2(net4734));
 sg13g2_a21oi_1 _18110_ (.A1(net5689),
    .A2(net4558),
    .Y(_02291_),
    .B1(_02290_));
 sg13g2_nor2_1 _18111_ (.A(net5529),
    .B(_02291_),
    .Y(_00938_));
 sg13g2_a21oi_1 _18112_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[1] ),
    .A2(net5160),
    .Y(_02292_),
    .B1(net4736));
 sg13g2_nand2b_1 _18113_ (.Y(_02293_),
    .B(_02292_),
    .A_N(_08902_));
 sg13g2_a21oi_1 _18114_ (.A1(_04310_),
    .A2(net4735),
    .Y(_02294_),
    .B1(net4560));
 sg13g2_a22oi_1 _18115_ (.Y(_02295_),
    .B1(_02293_),
    .B2(_02294_),
    .A2(net4560),
    .A1(net3068));
 sg13g2_nor2_1 _18116_ (.A(net5532),
    .B(net3069),
    .Y(_00939_));
 sg13g2_a21oi_1 _18117_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[2] ),
    .A2(net5162),
    .Y(_02296_),
    .B1(net4738));
 sg13g2_nand2b_1 _18118_ (.Y(_02297_),
    .B(_02296_),
    .A_N(_08913_));
 sg13g2_a21oi_1 _18119_ (.A1(_04311_),
    .A2(net4737),
    .Y(_02298_),
    .B1(net4563));
 sg13g2_a22oi_1 _18120_ (.Y(_02299_),
    .B1(_02297_),
    .B2(_02298_),
    .A2(net4563),
    .A1(net3079));
 sg13g2_nor2_1 _18121_ (.A(net5534),
    .B(net3080),
    .Y(_00940_));
 sg13g2_a221oi_1 _18122_ (.B2(\TRNG.Padded_Out[67] ),
    .C1(net4737),
    .B1(net5148),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[3] ),
    .Y(_02300_),
    .A2(net5162));
 sg13g2_a22oi_1 _18123_ (.Y(_02301_),
    .B1(_02300_),
    .B2(_08925_),
    .A2(net4737),
    .A1(_04312_));
 sg13g2_o21ai_1 _18124_ (.B1(net5475),
    .Y(_02302_),
    .A1(net4560),
    .A2(_02301_));
 sg13g2_a21oi_1 _18125_ (.A1(_04276_),
    .A2(net4560),
    .Y(_00941_),
    .B1(_02302_));
 sg13g2_a21oi_1 _18126_ (.A1(net3847),
    .A2(net5162),
    .Y(_02303_),
    .B1(net4740));
 sg13g2_a221oi_1 _18127_ (.B2(_08939_),
    .C1(net4564),
    .B1(_02303_),
    .A1(_04313_),
    .Y(_02304_),
    .A2(net4740));
 sg13g2_a21oi_1 _18128_ (.A1(net5682),
    .A2(net4564),
    .Y(_02305_),
    .B1(_02304_));
 sg13g2_nor2_1 _18129_ (.A(net5535),
    .B(_02305_),
    .Y(_00942_));
 sg13g2_a21oi_1 _18130_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[5] ),
    .A2(net5161),
    .Y(_02306_),
    .B1(net4740));
 sg13g2_nand2b_1 _18131_ (.Y(_02307_),
    .B(_02306_),
    .A_N(_08951_));
 sg13g2_a21oi_1 _18132_ (.A1(_04314_),
    .A2(net4740),
    .Y(_02308_),
    .B1(net4564));
 sg13g2_a22oi_1 _18133_ (.Y(_02309_),
    .B1(_02307_),
    .B2(_02308_),
    .A2(net4564),
    .A1(net2439));
 sg13g2_nor2_1 _18134_ (.A(net5540),
    .B(net2440),
    .Y(_00943_));
 sg13g2_a21oi_1 _18135_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[6] ),
    .A2(net5161),
    .Y(_02310_),
    .B1(net4739));
 sg13g2_nand2b_1 _18136_ (.Y(_02311_),
    .B(_02310_),
    .A_N(_08962_));
 sg13g2_a21oi_1 _18137_ (.A1(_04315_),
    .A2(net4739),
    .Y(_02312_),
    .B1(net4565));
 sg13g2_a22oi_1 _18138_ (.Y(_02313_),
    .B1(_02311_),
    .B2(_02312_),
    .A2(net4565),
    .A1(net5678));
 sg13g2_nor2_1 _18139_ (.A(net5537),
    .B(net3702),
    .Y(_00944_));
 sg13g2_a21oi_1 _18140_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[7] ),
    .A2(net5161),
    .Y(_02314_),
    .B1(net4739));
 sg13g2_nand2b_1 _18141_ (.Y(_02315_),
    .B(_02314_),
    .A_N(_08975_));
 sg13g2_a21oi_1 _18142_ (.A1(_04316_),
    .A2(net4739),
    .Y(_02316_),
    .B1(net4565));
 sg13g2_a22oi_1 _18143_ (.Y(_02317_),
    .B1(_02315_),
    .B2(_02316_),
    .A2(net4565),
    .A1(net3622));
 sg13g2_nor2_1 _18144_ (.A(net5537),
    .B(net3623),
    .Y(_00945_));
 sg13g2_a21oi_1 _18145_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[8] ),
    .A2(net5161),
    .Y(_02318_),
    .B1(net4739));
 sg13g2_nand2b_1 _18146_ (.Y(_02319_),
    .B(_02318_),
    .A_N(_08988_));
 sg13g2_a21oi_1 _18147_ (.A1(_04317_),
    .A2(net4739),
    .Y(_02320_),
    .B1(net4565));
 sg13g2_a22oi_1 _18148_ (.Y(_02321_),
    .B1(_02319_),
    .B2(_02320_),
    .A2(net4565),
    .A1(net5673));
 sg13g2_nor2_1 _18149_ (.A(net5537),
    .B(net3658),
    .Y(_00946_));
 sg13g2_a21oi_1 _18150_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[9] ),
    .A2(net5161),
    .Y(_02322_),
    .B1(net4739));
 sg13g2_a221oi_1 _18151_ (.B2(_09001_),
    .C1(net4565),
    .B1(_02322_),
    .A1(_04318_),
    .Y(_02323_),
    .A2(net4739));
 sg13g2_a21oi_1 _18152_ (.A1(net3626),
    .A2(net4564),
    .Y(_02324_),
    .B1(_02323_));
 sg13g2_nor2_1 _18153_ (.A(net5540),
    .B(net3627),
    .Y(_00947_));
 sg13g2_a21oi_1 _18154_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[10] ),
    .A2(net5162),
    .Y(_02325_),
    .B1(net4737));
 sg13g2_a221oi_1 _18155_ (.B2(_09013_),
    .C1(net4563),
    .B1(_02325_),
    .A1(_04319_),
    .Y(_02326_),
    .A2(net4737));
 sg13g2_a21oi_1 _18156_ (.A1(net3641),
    .A2(net4562),
    .Y(_02327_),
    .B1(_02326_));
 sg13g2_nor2_1 _18157_ (.A(net5534),
    .B(net3642),
    .Y(_00948_));
 sg13g2_a21oi_1 _18158_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[11] ),
    .A2(net5160),
    .Y(_02328_),
    .B1(net4737));
 sg13g2_a221oi_1 _18159_ (.B2(_09025_),
    .C1(net4563),
    .B1(_02328_),
    .A1(_04320_),
    .Y(_02329_),
    .A2(net4737));
 sg13g2_a21oi_1 _18160_ (.A1(net3528),
    .A2(net4557),
    .Y(_02330_),
    .B1(_02329_));
 sg13g2_nor2_1 _18161_ (.A(net5530),
    .B(_02330_),
    .Y(_00949_));
 sg13g2_a21oi_1 _18162_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[12] ),
    .A2(net5160),
    .Y(_02331_),
    .B1(net4737));
 sg13g2_nand2b_1 _18163_ (.Y(_02332_),
    .B(_02331_),
    .A_N(_09036_));
 sg13g2_a21oi_1 _18164_ (.A1(_04321_),
    .A2(net4735),
    .Y(_02333_),
    .B1(net4563));
 sg13g2_a22oi_1 _18165_ (.Y(_02334_),
    .B1(_02332_),
    .B2(_02333_),
    .A2(net4563),
    .A1(net3532));
 sg13g2_nor2_1 _18166_ (.A(net5534),
    .B(net3533),
    .Y(_00950_));
 sg13g2_a21oi_1 _18167_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[13] ),
    .A2(net5163),
    .Y(_02335_),
    .B1(net4736));
 sg13g2_nand2b_1 _18168_ (.Y(_02336_),
    .B(_02335_),
    .A_N(_09047_));
 sg13g2_a21oi_1 _18169_ (.A1(_04322_),
    .A2(net4736),
    .Y(_02337_),
    .B1(net4560));
 sg13g2_a22oi_1 _18170_ (.Y(_02338_),
    .B1(_02336_),
    .B2(_02337_),
    .A2(net4561),
    .A1(net3519));
 sg13g2_nor2_1 _18171_ (.A(net5532),
    .B(net3520),
    .Y(_00951_));
 sg13g2_a21oi_1 _18172_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[14] ),
    .A2(net5163),
    .Y(_02339_),
    .B1(net4735));
 sg13g2_nand2b_1 _18173_ (.Y(_02340_),
    .B(_02339_),
    .A_N(_09058_));
 sg13g2_a21oi_1 _18174_ (.A1(_04323_),
    .A2(net4735),
    .Y(_02341_),
    .B1(net4563));
 sg13g2_a22oi_1 _18175_ (.Y(_02342_),
    .B1(_02340_),
    .B2(_02341_),
    .A2(net4563),
    .A1(net3743));
 sg13g2_nor2_1 _18176_ (.A(net5534),
    .B(net3744),
    .Y(_00952_));
 sg13g2_a21oi_1 _18177_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[15] ),
    .A2(net5159),
    .Y(_02343_),
    .B1(net4735));
 sg13g2_nand2b_1 _18178_ (.Y(_02344_),
    .B(_02343_),
    .A_N(_09069_));
 sg13g2_a21oi_1 _18179_ (.A1(_04324_),
    .A2(net4735),
    .Y(_02345_),
    .B1(net4561));
 sg13g2_a22oi_1 _18180_ (.Y(_02346_),
    .B1(_02344_),
    .B2(_02345_),
    .A2(net4561),
    .A1(net3421));
 sg13g2_nor2_1 _18181_ (.A(net5531),
    .B(net3422),
    .Y(_00953_));
 sg13g2_a21oi_1 _18182_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[16] ),
    .A2(net5159),
    .Y(_02347_),
    .B1(net4735));
 sg13g2_a221oi_1 _18183_ (.B2(_09081_),
    .C1(net4560),
    .B1(_02347_),
    .A1(_04325_),
    .Y(_02348_),
    .A2(net4735));
 sg13g2_a21oi_1 _18184_ (.A1(net3698),
    .A2(net4564),
    .Y(_02349_),
    .B1(_02348_));
 sg13g2_nor2_1 _18185_ (.A(net5540),
    .B(_02349_),
    .Y(_00954_));
 sg13g2_a21oi_1 _18186_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[17] ),
    .A2(net5159),
    .Y(_02350_),
    .B1(net4734));
 sg13g2_a221oi_1 _18187_ (.B2(_09093_),
    .C1(net4559),
    .B1(_02350_),
    .A1(_04326_),
    .Y(_02351_),
    .A2(net4734));
 sg13g2_a21oi_1 _18188_ (.A1(net3511),
    .A2(net4558),
    .Y(_02352_),
    .B1(_02351_));
 sg13g2_nor2_1 _18189_ (.A(net5532),
    .B(net3512),
    .Y(_00955_));
 sg13g2_a21oi_1 _18190_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[18] ),
    .A2(net5159),
    .Y(_02353_),
    .B1(net4732));
 sg13g2_nand2b_1 _18191_ (.Y(_02354_),
    .B(_02353_),
    .A_N(_09104_));
 sg13g2_a21oi_1 _18192_ (.A1(_04327_),
    .A2(net4732),
    .Y(_02355_),
    .B1(net4559));
 sg13g2_a22oi_1 _18193_ (.Y(_02356_),
    .B1(_02354_),
    .B2(_02355_),
    .A2(net4558),
    .A1(net2418));
 sg13g2_nor2_1 _18194_ (.A(net5529),
    .B(net2419),
    .Y(_00956_));
 sg13g2_a21oi_1 _18195_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[19] ),
    .A2(net5160),
    .Y(_02357_),
    .B1(net4732));
 sg13g2_a221oi_1 _18196_ (.B2(_09116_),
    .C1(net4557),
    .B1(_02357_),
    .A1(_04328_),
    .Y(_02358_),
    .A2(net4732));
 sg13g2_a21oi_1 _18197_ (.A1(net3453),
    .A2(net4557),
    .Y(_02359_),
    .B1(_02358_));
 sg13g2_nor2_1 _18198_ (.A(net5529),
    .B(net3454),
    .Y(_00957_));
 sg13g2_a21oi_1 _18199_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[20] ),
    .A2(net5159),
    .Y(_02360_),
    .B1(net4733));
 sg13g2_a221oi_1 _18200_ (.B2(_09128_),
    .C1(net4558),
    .B1(_02360_),
    .A1(_04329_),
    .Y(_02361_),
    .A2(net4733));
 sg13g2_a21oi_1 _18201_ (.A1(net2631),
    .A2(net4558),
    .Y(_02362_),
    .B1(_02361_));
 sg13g2_nor2_1 _18202_ (.A(net5532),
    .B(net2632),
    .Y(_00958_));
 sg13g2_a21oi_1 _18203_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[21] ),
    .A2(net5159),
    .Y(_02363_),
    .B1(net4733));
 sg13g2_a221oi_1 _18204_ (.B2(_09141_),
    .C1(net4557),
    .B1(_02363_),
    .A1(_04330_),
    .Y(_02364_),
    .A2(net4733));
 sg13g2_a21oi_1 _18205_ (.A1(net5642),
    .A2(net4557),
    .Y(_02365_),
    .B1(_02364_));
 sg13g2_nor2_1 _18206_ (.A(net5529),
    .B(net3721),
    .Y(_00959_));
 sg13g2_a21oi_1 _18207_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[22] ),
    .A2(net5159),
    .Y(_02366_),
    .B1(net4732));
 sg13g2_nand2b_1 _18208_ (.Y(_02367_),
    .B(_02366_),
    .A_N(_09152_));
 sg13g2_a21oi_1 _18209_ (.A1(_04331_),
    .A2(net4732),
    .Y(_02368_),
    .B1(net4558));
 sg13g2_a22oi_1 _18210_ (.Y(_02369_),
    .B1(_02367_),
    .B2(_02368_),
    .A2(net4558),
    .A1(net5639));
 sg13g2_nor2_1 _18211_ (.A(net5529),
    .B(net3633),
    .Y(_00960_));
 sg13g2_a21oi_1 _18212_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[23] ),
    .A2(net5160),
    .Y(_02370_),
    .B1(net4732));
 sg13g2_a221oi_1 _18213_ (.B2(_09164_),
    .C1(net4557),
    .B1(_02370_),
    .A1(_04332_),
    .Y(_02371_),
    .A2(net4732));
 sg13g2_a21oi_1 _18214_ (.A1(net3671),
    .A2(net4557),
    .Y(_02372_),
    .B1(_02371_));
 sg13g2_nor2_1 _18215_ (.A(net5530),
    .B(net3672),
    .Y(_00961_));
 sg13g2_a21oi_1 _18216_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[24] ),
    .A2(net5160),
    .Y(_02373_),
    .B1(net4733));
 sg13g2_a221oi_1 _18217_ (.B2(_02169_),
    .C1(net4560),
    .B1(_02373_),
    .A1(_04333_),
    .Y(_02374_),
    .A2(net4733));
 sg13g2_a21oi_1 _18218_ (.A1(net3706),
    .A2(net4559),
    .Y(_02375_),
    .B1(_02374_));
 sg13g2_nor2_1 _18219_ (.A(net5529),
    .B(net3707),
    .Y(_00962_));
 sg13g2_a21oi_1 _18220_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[25] ),
    .A2(net5163),
    .Y(_02376_),
    .B1(net4736));
 sg13g2_a221oi_1 _18221_ (.B2(_02181_),
    .C1(net4560),
    .B1(_02376_),
    .A1(_04334_),
    .Y(_02377_),
    .A2(net4736));
 sg13g2_a21oi_1 _18222_ (.A1(net3529),
    .A2(net4557),
    .Y(_02378_),
    .B1(_02377_));
 sg13g2_nor2_1 _18223_ (.A(net5529),
    .B(_02378_),
    .Y(_00963_));
 sg13g2_a21oi_1 _18224_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[26] ),
    .A2(net5160),
    .Y(_02379_),
    .B1(net4741));
 sg13g2_a221oi_1 _18225_ (.B2(_02194_),
    .C1(net4562),
    .B1(_02379_),
    .A1(_04335_),
    .Y(_02380_),
    .A2(net4741));
 sg13g2_a21oi_1 _18226_ (.A1(net3673),
    .A2(net4562),
    .Y(_02381_),
    .B1(_02380_));
 sg13g2_nor2_1 _18227_ (.A(net5535),
    .B(net3674),
    .Y(_00964_));
 sg13g2_a21oi_1 _18228_ (.A1(net3816),
    .A2(net5162),
    .Y(_02382_),
    .B1(net4738));
 sg13g2_nand2b_1 _18229_ (.Y(_02383_),
    .B(_02382_),
    .A_N(_02205_));
 sg13g2_a21oi_1 _18230_ (.A1(_04336_),
    .A2(net4738),
    .Y(_02384_),
    .B1(net4562));
 sg13g2_a22oi_1 _18231_ (.Y(_02385_),
    .B1(_02383_),
    .B2(_02384_),
    .A2(net4562),
    .A1(net5628));
 sg13g2_nor2_1 _18232_ (.A(net5535),
    .B(_02385_),
    .Y(_00965_));
 sg13g2_a21oi_1 _18233_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[28] ),
    .A2(net5162),
    .Y(_02386_),
    .B1(net4738));
 sg13g2_nand2b_1 _18234_ (.Y(_02387_),
    .B(_02386_),
    .A_N(_02217_));
 sg13g2_a21oi_1 _18235_ (.A1(_04337_),
    .A2(net4738),
    .Y(_02388_),
    .B1(net4562));
 sg13g2_a22oi_1 _18236_ (.Y(_02389_),
    .B1(_02387_),
    .B2(_02388_),
    .A2(net4562),
    .A1(net3467));
 sg13g2_nor2_1 _18237_ (.A(net5535),
    .B(net3468),
    .Y(_00966_));
 sg13g2_a21oi_1 _18238_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[29] ),
    .A2(net5162),
    .Y(_02390_),
    .B1(net4738));
 sg13g2_nand2b_1 _18239_ (.Y(_02391_),
    .B(_02390_),
    .A_N(_02228_));
 sg13g2_a21oi_1 _18240_ (.A1(_04338_),
    .A2(net4738),
    .Y(_02392_),
    .B1(net4566));
 sg13g2_a22oi_1 _18241_ (.Y(_02393_),
    .B1(_02391_),
    .B2(_02392_),
    .A2(net4562),
    .A1(net2492));
 sg13g2_nor2_1 _18242_ (.A(net5535),
    .B(net2493),
    .Y(_00967_));
 sg13g2_a21oi_1 _18243_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[30] ),
    .A2(net5161),
    .Y(_02394_),
    .B1(net4740));
 sg13g2_nand2b_1 _18244_ (.Y(_02395_),
    .B(_02394_),
    .A_N(_02239_));
 sg13g2_a21oi_1 _18245_ (.A1(_04339_),
    .A2(net4740),
    .Y(_02396_),
    .B1(net4566));
 sg13g2_a22oi_1 _18246_ (.Y(_02397_),
    .B1(_02395_),
    .B2(_02396_),
    .A2(net4566),
    .A1(net5620));
 sg13g2_nor2_1 _18247_ (.A(net5540),
    .B(net3688),
    .Y(_00968_));
 sg13g2_a21oi_1 _18248_ (.A1(\TRNG.sha256.expand.exp_ctrl.final_sum[31] ),
    .A2(net5163),
    .Y(_02398_),
    .B1(net4740));
 sg13g2_nand2b_1 _18249_ (.Y(_02399_),
    .B(_02398_),
    .A_N(_02251_));
 sg13g2_a21oi_1 _18250_ (.A1(_04340_),
    .A2(net4740),
    .Y(_02400_),
    .B1(net4564));
 sg13g2_a22oi_1 _18251_ (.Y(_02401_),
    .B1(_02399_),
    .B2(_02400_),
    .A2(net4564),
    .A1(net3638));
 sg13g2_nor2_1 _18252_ (.A(net5540),
    .B(net3639),
    .Y(_00969_));
 sg13g2_o21ai_1 _18253_ (.B1(_08811_),
    .Y(_02402_),
    .A1(\TRNG.sha256.expand.exp_ctrl.write_en1 ),
    .A2(_02256_));
 sg13g2_o21ai_1 _18254_ (.B1(net5478),
    .Y(_00970_),
    .A1(net5158),
    .A2(_02402_));
 sg13g2_o21ai_1 _18255_ (.B1(net5478),
    .Y(_02403_),
    .A1(\TRNG.sha256.expand.exp_ctrl.j[0] ),
    .A2(net4986));
 sg13g2_a21oi_1 _18256_ (.A1(_04275_),
    .A2(net4986),
    .Y(_00971_),
    .B1(_02403_));
 sg13g2_a21oi_1 _18257_ (.A1(\TRNG.sha256.expand.exp_ctrl.j[0] ),
    .A2(net4986),
    .Y(_02404_),
    .B1(net2494));
 sg13g2_and3_1 _18258_ (.X(_02405_),
    .A(net2494),
    .B(\TRNG.sha256.expand.exp_ctrl.j[0] ),
    .C(net4986));
 sg13g2_nor3_1 _18259_ (.A(net5541),
    .B(net2495),
    .C(_02405_),
    .Y(_00972_));
 sg13g2_and2_1 _18260_ (.A(net3459),
    .B(_02405_),
    .X(_02406_));
 sg13g2_o21ai_1 _18261_ (.B1(net5478),
    .Y(_02407_),
    .A1(net3459),
    .A2(_02405_));
 sg13g2_nor2_1 _18262_ (.A(_02406_),
    .B(net3460),
    .Y(_00973_));
 sg13g2_a21oi_1 _18263_ (.A1(net3398),
    .A2(_02406_),
    .Y(_02408_),
    .B1(net5541));
 sg13g2_o21ai_1 _18264_ (.B1(_02408_),
    .Y(_02409_),
    .A1(net3398),
    .A2(_02406_));
 sg13g2_inv_1 _18265_ (.Y(_00974_),
    .A(net3399));
 sg13g2_o21ai_1 _18266_ (.B1(net5479),
    .Y(_02410_),
    .A1(\TRNG.sha256.expand.exp_ctrl.j_2[0] ),
    .A2(net4985));
 sg13g2_a21oi_1 _18267_ (.A1(_04274_),
    .A2(net4985),
    .Y(_00975_),
    .B1(_02410_));
 sg13g2_nand3_1 _18268_ (.B(net3749),
    .C(net4985),
    .A(net3386),
    .Y(_02411_));
 sg13g2_a21o_1 _18269_ (.A2(net4985),
    .A1(net3749),
    .B1(net3386),
    .X(_02412_));
 sg13g2_a21o_1 _18270_ (.A2(_02412_),
    .A1(_02411_),
    .B1(net5539),
    .X(_00976_));
 sg13g2_nand4_1 _18271_ (.B(net3386),
    .C(net3749),
    .A(net3285),
    .Y(_02413_),
    .D(net4985));
 sg13g2_nand2b_1 _18272_ (.Y(_02414_),
    .B(_02411_),
    .A_N(net3285));
 sg13g2_a21o_1 _18273_ (.A2(_02414_),
    .A1(_02413_),
    .B1(net5538),
    .X(_00977_));
 sg13g2_a21oi_1 _18274_ (.A1(net2064),
    .A2(_02413_),
    .Y(_02415_),
    .B1(net5538));
 sg13g2_o21ai_1 _18275_ (.B1(_02415_),
    .Y(_00978_),
    .A1(net2064),
    .A2(_02413_));
 sg13g2_a21oi_1 _18276_ (.A1(net1532),
    .A2(net4985),
    .Y(_02416_),
    .B1(net5539));
 sg13g2_o21ai_1 _18277_ (.B1(_02416_),
    .Y(_00979_),
    .A1(_04273_),
    .A2(_02263_));
 sg13g2_a21oi_1 _18278_ (.A1(net2311),
    .A2(net4985),
    .Y(_02417_),
    .B1(net2388));
 sg13g2_and3_1 _18279_ (.X(_02418_),
    .A(net2388),
    .B(net2311),
    .C(net4985));
 sg13g2_nor3_1 _18280_ (.A(net5538),
    .B(_02417_),
    .C(_02418_),
    .Y(_00980_));
 sg13g2_or2_1 _18281_ (.X(_02419_),
    .B(_02418_),
    .A(net2532));
 sg13g2_nand2_1 _18282_ (.Y(_02420_),
    .A(net2532),
    .B(_02418_));
 sg13g2_and3_1 _18283_ (.X(_00981_),
    .A(net5478),
    .B(_02419_),
    .C(_02420_));
 sg13g2_a21oi_1 _18284_ (.A1(net2289),
    .A2(_02420_),
    .Y(_02421_),
    .B1(net5538));
 sg13g2_o21ai_1 _18285_ (.B1(_02421_),
    .Y(_00982_),
    .A1(net2289),
    .A2(_02420_));
 sg13g2_a21oi_1 _18286_ (.A1(net2376),
    .A2(net4986),
    .Y(_02422_),
    .B1(net5536));
 sg13g2_o21ai_1 _18287_ (.B1(_02422_),
    .Y(_00983_),
    .A1(_04272_),
    .A2(net4986));
 sg13g2_a21oi_1 _18288_ (.A1(\TRNG.sha256.expand.exp_ctrl.j_15[0] ),
    .A2(net4986),
    .Y(_02423_),
    .B1(net2655));
 sg13g2_and3_1 _18289_ (.X(_02424_),
    .A(net2655),
    .B(\TRNG.sha256.expand.exp_ctrl.j_15[0] ),
    .C(net4986));
 sg13g2_nor3_1 _18290_ (.A(net5536),
    .B(net2656),
    .C(_02424_),
    .Y(_00984_));
 sg13g2_and2_1 _18291_ (.A(net3430),
    .B(_02424_),
    .X(_02425_));
 sg13g2_o21ai_1 _18292_ (.B1(net5480),
    .Y(_02426_),
    .A1(net3430),
    .A2(_02424_));
 sg13g2_nor2_1 _18293_ (.A(_02425_),
    .B(net3431),
    .Y(_00985_));
 sg13g2_a21oi_1 _18294_ (.A1(net3450),
    .A2(_02425_),
    .Y(_02427_),
    .B1(net5536));
 sg13g2_o21ai_1 _18295_ (.B1(_02427_),
    .Y(_02428_),
    .A1(net3450),
    .A2(_02425_));
 sg13g2_inv_1 _18296_ (.Y(_00986_),
    .A(_02428_));
 sg13g2_o21ai_1 _18297_ (.B1(net5476),
    .Y(_02429_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[0] ),
    .A2(net4990));
 sg13g2_a21oi_1 _18298_ (.A1(_04271_),
    .A2(net4990),
    .Y(_00987_),
    .B1(_02429_));
 sg13g2_o21ai_1 _18299_ (.B1(net5476),
    .Y(_02430_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[1] ),
    .A2(net4991));
 sg13g2_a21oi_1 _18300_ (.A1(_04270_),
    .A2(net4991),
    .Y(_00988_),
    .B1(_02430_));
 sg13g2_o21ai_1 _18301_ (.B1(net5481),
    .Y(_02431_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[2] ),
    .A2(net4994));
 sg13g2_a21oi_1 _18302_ (.A1(_04269_),
    .A2(net4994),
    .Y(_00989_),
    .B1(_02431_));
 sg13g2_o21ai_1 _18303_ (.B1(net5477),
    .Y(_02432_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[3] ),
    .A2(net4994));
 sg13g2_a21oi_1 _18304_ (.A1(_04268_),
    .A2(net4994),
    .Y(_00990_),
    .B1(_02432_));
 sg13g2_o21ai_1 _18305_ (.B1(net5477),
    .Y(_02433_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[4] ),
    .A2(net4993));
 sg13g2_a21oi_1 _18306_ (.A1(_04267_),
    .A2(net4996),
    .Y(_00991_),
    .B1(_02433_));
 sg13g2_o21ai_1 _18307_ (.B1(net5479),
    .Y(_02434_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[5] ),
    .A2(net4996));
 sg13g2_a21oi_1 _18308_ (.A1(_04266_),
    .A2(net4997),
    .Y(_00992_),
    .B1(_02434_));
 sg13g2_o21ai_1 _18309_ (.B1(net5480),
    .Y(_02435_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[6] ),
    .A2(net4995));
 sg13g2_a21oi_1 _18310_ (.A1(_04265_),
    .A2(net4995),
    .Y(_00993_),
    .B1(_02435_));
 sg13g2_o21ai_1 _18311_ (.B1(net5480),
    .Y(_02436_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[7] ),
    .A2(net4995));
 sg13g2_a21oi_1 _18312_ (.A1(_04264_),
    .A2(net4995),
    .Y(_00994_),
    .B1(_02436_));
 sg13g2_o21ai_1 _18313_ (.B1(net5480),
    .Y(_02437_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[8] ),
    .A2(net4995));
 sg13g2_a21oi_1 _18314_ (.A1(_04263_),
    .A2(net4995),
    .Y(_00995_),
    .B1(_02437_));
 sg13g2_o21ai_1 _18315_ (.B1(net5477),
    .Y(_02438_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[9] ),
    .A2(net4995));
 sg13g2_a21oi_1 _18316_ (.A1(_04262_),
    .A2(net4995),
    .Y(_00996_),
    .B1(_02438_));
 sg13g2_o21ai_1 _18317_ (.B1(net5477),
    .Y(_02439_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[10] ),
    .A2(net4994));
 sg13g2_a21oi_1 _18318_ (.A1(_04261_),
    .A2(net4994),
    .Y(_00997_),
    .B1(_02439_));
 sg13g2_o21ai_1 _18319_ (.B1(net5477),
    .Y(_02440_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[11] ),
    .A2(net4991));
 sg13g2_a21oi_1 _18320_ (.A1(_04260_),
    .A2(net4991),
    .Y(_00998_),
    .B1(_02440_));
 sg13g2_o21ai_1 _18321_ (.B1(net5477),
    .Y(_02441_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[12] ),
    .A2(net4994));
 sg13g2_a21oi_1 _18322_ (.A1(_04259_),
    .A2(net4994),
    .Y(_00999_),
    .B1(_02441_));
 sg13g2_o21ai_1 _18323_ (.B1(net5475),
    .Y(_02442_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[13] ),
    .A2(net4991));
 sg13g2_a21oi_1 _18324_ (.A1(_04258_),
    .A2(net4992),
    .Y(_01000_),
    .B1(_02442_));
 sg13g2_o21ai_1 _18325_ (.B1(net5476),
    .Y(_02443_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[14] ),
    .A2(net4991));
 sg13g2_a21oi_1 _18326_ (.A1(_04257_),
    .A2(net4991),
    .Y(_01001_),
    .B1(_02443_));
 sg13g2_o21ai_1 _18327_ (.B1(net5476),
    .Y(_02444_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[15] ),
    .A2(net4990));
 sg13g2_a21oi_1 _18328_ (.A1(_04256_),
    .A2(net4991),
    .Y(_01002_),
    .B1(_02444_));
 sg13g2_o21ai_1 _18329_ (.B1(net5475),
    .Y(_02445_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[16] ),
    .A2(net4989));
 sg13g2_a21oi_1 _18330_ (.A1(_04255_),
    .A2(net4989),
    .Y(_01003_),
    .B1(_02445_));
 sg13g2_o21ai_1 _18331_ (.B1(net5476),
    .Y(_02446_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[17] ),
    .A2(net4990));
 sg13g2_a21oi_1 _18332_ (.A1(_04254_),
    .A2(net4990),
    .Y(_01004_),
    .B1(_02446_));
 sg13g2_o21ai_1 _18333_ (.B1(net5475),
    .Y(_02447_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[18] ),
    .A2(net4990));
 sg13g2_a21oi_1 _18334_ (.A1(_04253_),
    .A2(net4990),
    .Y(_01005_),
    .B1(_02447_));
 sg13g2_o21ai_1 _18335_ (.B1(net5475),
    .Y(_02448_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[19] ),
    .A2(net4988));
 sg13g2_a21oi_1 _18336_ (.A1(_04252_),
    .A2(net4988),
    .Y(_01006_),
    .B1(_02448_));
 sg13g2_o21ai_1 _18337_ (.B1(net5475),
    .Y(_02449_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[20] ),
    .A2(net4988));
 sg13g2_a21oi_1 _18338_ (.A1(_04251_),
    .A2(net4988),
    .Y(_01007_),
    .B1(_02449_));
 sg13g2_o21ai_1 _18339_ (.B1(net5482),
    .Y(_02450_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[21] ),
    .A2(net4988));
 sg13g2_a21oi_1 _18340_ (.A1(_04250_),
    .A2(net4989),
    .Y(_01008_),
    .B1(_02450_));
 sg13g2_o21ai_1 _18341_ (.B1(net5475),
    .Y(_02451_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[22] ),
    .A2(net4988));
 sg13g2_a21oi_1 _18342_ (.A1(_04249_),
    .A2(net4988),
    .Y(_01009_),
    .B1(_02451_));
 sg13g2_o21ai_1 _18343_ (.B1(net5482),
    .Y(_02452_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[23] ),
    .A2(net4989));
 sg13g2_a21oi_1 _18344_ (.A1(_04248_),
    .A2(net4988),
    .Y(_01010_),
    .B1(_02452_));
 sg13g2_o21ai_1 _18345_ (.B1(net5475),
    .Y(_02453_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[24] ),
    .A2(net4989));
 sg13g2_a21oi_1 _18346_ (.A1(_04247_),
    .A2(net4989),
    .Y(_01011_),
    .B1(_02453_));
 sg13g2_o21ai_1 _18347_ (.B1(net5476),
    .Y(_02454_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[25] ),
    .A2(net4992));
 sg13g2_a21oi_1 _18348_ (.A1(_04246_),
    .A2(net4992),
    .Y(_01012_),
    .B1(_02454_));
 sg13g2_o21ai_1 _18349_ (.B1(net5481),
    .Y(_02455_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[26] ),
    .A2(net4993));
 sg13g2_a21oi_1 _18350_ (.A1(_04245_),
    .A2(net4993),
    .Y(_01013_),
    .B1(_02455_));
 sg13g2_o21ai_1 _18351_ (.B1(net5481),
    .Y(_02456_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[27] ),
    .A2(net4993));
 sg13g2_a21oi_1 _18352_ (.A1(_04244_),
    .A2(net4993),
    .Y(_01014_),
    .B1(_02456_));
 sg13g2_o21ai_1 _18353_ (.B1(net5477),
    .Y(_02457_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[28] ),
    .A2(net4993));
 sg13g2_a21oi_1 _18354_ (.A1(_04243_),
    .A2(net4993),
    .Y(_01015_),
    .B1(_02457_));
 sg13g2_o21ai_1 _18355_ (.B1(net5477),
    .Y(_02458_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[29] ),
    .A2(net4997));
 sg13g2_a21oi_1 _18356_ (.A1(_04242_),
    .A2(net4993),
    .Y(_01016_),
    .B1(_02458_));
 sg13g2_o21ai_1 _18357_ (.B1(net5479),
    .Y(_02459_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[30] ),
    .A2(net4996));
 sg13g2_a21oi_1 _18358_ (.A1(_04241_),
    .A2(net4997),
    .Y(_01017_),
    .B1(_02459_));
 sg13g2_o21ai_1 _18359_ (.B1(net5479),
    .Y(_02460_),
    .A1(\TRNG.sha256.expand.exp_ctrl.final_sum[31] ),
    .A2(net4996));
 sg13g2_a21oi_1 _18360_ (.A1(_04240_),
    .A2(net4996),
    .Y(_01018_),
    .B1(_02460_));
 sg13g2_and4_2 _18361_ (.A(\TRNG.sha256.expand.exp_ctrl.write_en1 ),
    .B(\TRNG.sha256.expand.address1[3] ),
    .C(\TRNG.sha256.expand.address1[2] ),
    .D(net5393),
    .X(_02461_));
 sg13g2_mux2_1 _18362_ (.A0(net2595),
    .A1(net5689),
    .S(net5115),
    .X(_01019_));
 sg13g2_mux2_1 _18363_ (.A0(net2607),
    .A1(net5688),
    .S(net5115),
    .X(_01020_));
 sg13g2_mux2_1 _18364_ (.A0(net2844),
    .A1(net5684),
    .S(net5116),
    .X(_01021_));
 sg13g2_nor2_1 _18365_ (.A(net2858),
    .B(net5117),
    .Y(_02462_));
 sg13g2_a21oi_1 _18366_ (.A1(net5496),
    .A2(net5117),
    .Y(_01022_),
    .B1(_02462_));
 sg13g2_mux2_1 _18367_ (.A0(net2663),
    .A1(net5682),
    .S(net5116),
    .X(_01023_));
 sg13g2_mux2_1 _18368_ (.A0(net2748),
    .A1(net5681),
    .S(net5116),
    .X(_01024_));
 sg13g2_mux2_1 _18369_ (.A0(net2803),
    .A1(net5676),
    .S(net5116),
    .X(_01025_));
 sg13g2_mux2_1 _18370_ (.A0(net2808),
    .A1(net5675),
    .S(net5118),
    .X(_01026_));
 sg13g2_mux2_1 _18371_ (.A0(net2789),
    .A1(net5671),
    .S(net5115),
    .X(_01027_));
 sg13g2_mux2_1 _18372_ (.A0(net2785),
    .A1(net5669),
    .S(net5118),
    .X(_01028_));
 sg13g2_mux2_1 _18373_ (.A0(net2800),
    .A1(net5667),
    .S(net5118),
    .X(_01029_));
 sg13g2_mux2_1 _18374_ (.A0(net2694),
    .A1(net5666),
    .S(net5115),
    .X(_01030_));
 sg13g2_mux2_1 _18375_ (.A0(net2772),
    .A1(net5663),
    .S(net5115),
    .X(_01031_));
 sg13g2_mux2_1 _18376_ (.A0(net2779),
    .A1(net5661),
    .S(net5115),
    .X(_01032_));
 sg13g2_mux2_1 _18377_ (.A0(net3168),
    .A1(net5658),
    .S(net5118),
    .X(_01033_));
 sg13g2_mux2_1 _18378_ (.A0(net2625),
    .A1(net5656),
    .S(net5117),
    .X(_01034_));
 sg13g2_mux2_1 _18379_ (.A0(net2888),
    .A1(net5654),
    .S(net5118),
    .X(_01035_));
 sg13g2_mux2_1 _18380_ (.A0(net2996),
    .A1(net5652),
    .S(net5117),
    .X(_01036_));
 sg13g2_mux2_1 _18381_ (.A0(net3056),
    .A1(net5648),
    .S(net5115),
    .X(_01037_));
 sg13g2_mux2_1 _18382_ (.A0(net2566),
    .A1(net5647),
    .S(net5115),
    .X(_01038_));
 sg13g2_mux2_1 _18383_ (.A0(net2832),
    .A1(net5644),
    .S(net5117),
    .X(_01039_));
 sg13g2_mux2_1 _18384_ (.A0(net2900),
    .A1(net5640),
    .S(net5119),
    .X(_01040_));
 sg13g2_mux2_1 _18385_ (.A0(net2814),
    .A1(net5637),
    .S(net5117),
    .X(_01041_));
 sg13g2_mux2_1 _18386_ (.A0(net2721),
    .A1(net5635),
    .S(net5119),
    .X(_01042_));
 sg13g2_mux2_1 _18387_ (.A0(net2750),
    .A1(net5634),
    .S(net5117),
    .X(_01043_));
 sg13g2_mux2_1 _18388_ (.A0(net2781),
    .A1(net5631),
    .S(net5117),
    .X(_01044_));
 sg13g2_mux2_1 _18389_ (.A0(net2949),
    .A1(net5630),
    .S(net5119),
    .X(_01045_));
 sg13g2_mux2_1 _18390_ (.A0(net2569),
    .A1(net5628),
    .S(net5116),
    .X(_01046_));
 sg13g2_mux2_1 _18391_ (.A0(net2720),
    .A1(net5624),
    .S(net5118),
    .X(_01047_));
 sg13g2_mux2_1 _18392_ (.A0(net2563),
    .A1(net5621),
    .S(net5118),
    .X(_01048_));
 sg13g2_mux2_1 _18393_ (.A0(net2637),
    .A1(net5618),
    .S(net5116),
    .X(_01049_));
 sg13g2_mux2_1 _18394_ (.A0(net2713),
    .A1(net5617),
    .S(net5118),
    .X(_01050_));
 sg13g2_nand2_1 _18395_ (.Y(_02463_),
    .A(_08795_),
    .B(_08799_));
 sg13g2_and2_1 _18396_ (.A(_08797_),
    .B(_08800_),
    .X(_02464_));
 sg13g2_nor2b_2 _18397_ (.A(_02463_),
    .B_N(_02464_),
    .Y(_02465_));
 sg13g2_nor2_1 _18398_ (.A(net5526),
    .B(_02465_),
    .Y(_01051_));
 sg13g2_o21ai_1 _18399_ (.B1(_08820_),
    .Y(_02466_),
    .A1(net5575),
    .A2(_08800_));
 sg13g2_nand2_1 _18400_ (.Y(_02467_),
    .A(_02465_),
    .B(_02466_));
 sg13g2_nor2_1 _18401_ (.A(net5614),
    .B(_02466_),
    .Y(_02468_));
 sg13g2_o21ai_1 _18402_ (.B1(net5473),
    .Y(_02469_),
    .A1(net3855),
    .A2(_02467_));
 sg13g2_nor2_1 _18403_ (.A(_02468_),
    .B(_02469_),
    .Y(_01052_));
 sg13g2_nor2_1 _18404_ (.A(net5611),
    .B(_02466_),
    .Y(_02470_));
 sg13g2_o21ai_1 _18405_ (.B1(net5473),
    .Y(_02471_),
    .A1(net5099),
    .A2(_02467_));
 sg13g2_nor2_1 _18406_ (.A(_02470_),
    .B(_02471_),
    .Y(_01053_));
 sg13g2_nor2_1 _18407_ (.A(net5608),
    .B(_02466_),
    .Y(_02472_));
 sg13g2_o21ai_1 _18408_ (.B1(net5473),
    .Y(_02473_),
    .A1(_06205_),
    .A2(_02467_));
 sg13g2_nor2_1 _18409_ (.A(_02472_),
    .B(_02473_),
    .Y(_01054_));
 sg13g2_nand3b_1 _18410_ (.B(_05983_),
    .C(_02466_),
    .Y(_02474_),
    .A_N(net5603));
 sg13g2_o21ai_1 _18411_ (.B1(_02465_),
    .Y(_02475_),
    .A1(net5601),
    .A2(_02474_));
 sg13g2_a21oi_1 _18412_ (.A1(net5601),
    .A2(_02474_),
    .Y(_02476_),
    .B1(_02475_));
 sg13g2_nor2_1 _18413_ (.A(net5526),
    .B(_02476_),
    .Y(_01055_));
 sg13g2_nand3_1 _18414_ (.B(_06000_),
    .C(_02466_),
    .A(_05951_),
    .Y(_02477_));
 sg13g2_xnor2_1 _18415_ (.Y(_02478_),
    .A(net5504),
    .B(_02477_));
 sg13g2_a21oi_1 _18416_ (.A1(_02465_),
    .A2(_02478_),
    .Y(_01056_),
    .B1(net5526));
 sg13g2_nor2_1 _18417_ (.A(net3384),
    .B(_02477_),
    .Y(_02479_));
 sg13g2_xnor2_1 _18418_ (.Y(_02480_),
    .A(net5579),
    .B(_02479_));
 sg13g2_a21oi_1 _18419_ (.A1(_02465_),
    .A2(_02480_),
    .Y(_01057_),
    .B1(net5526));
 sg13g2_xnor2_1 _18420_ (.Y(_02481_),
    .A(net5575),
    .B(_08821_));
 sg13g2_a22oi_1 _18421_ (.Y(_02482_),
    .B1(_02464_),
    .B2(_02481_),
    .A2(_02463_),
    .A1(_08800_));
 sg13g2_a22oi_1 _18422_ (.Y(_02483_),
    .B1(_02466_),
    .B2(_02482_),
    .A2(_08820_),
    .A1(net5575));
 sg13g2_nor2_1 _18423_ (.A(net5526),
    .B(net3827),
    .Y(_01058_));
 sg13g2_and2_1 _18424_ (.A(net1184),
    .B(net1135),
    .X(_01059_));
 sg13g2_and2_1 _18425_ (.A(net1135),
    .B(net1149),
    .X(_01060_));
 sg13g2_and2_1 _18426_ (.A(net1135),
    .B(net1148),
    .X(_01061_));
 sg13g2_and2_1 _18427_ (.A(net1135),
    .B(net1703),
    .X(_01062_));
 sg13g2_and2_1 _18428_ (.A(\TRNG.hash[161] ),
    .B(net5831),
    .X(_02484_));
 sg13g2_a221oi_1 _18429_ (.B2(\TRNG.hash[129] ),
    .C1(_02484_),
    .B1(net5352),
    .A1(net3765),
    .Y(_02485_),
    .A2(net5187));
 sg13g2_a21oi_1 _18430_ (.A1(net5089),
    .A2(net3766),
    .Y(_01063_),
    .B1(net5521));
 sg13g2_nor2_2 _18431_ (.A(net5097),
    .B(net5352),
    .Y(_02486_));
 sg13g2_nand2_1 _18432_ (.Y(_02487_),
    .A(net5090),
    .B(net5177));
 sg13g2_nand2b_1 _18433_ (.Y(_02488_),
    .B(_00147_),
    .A_N(_06921_));
 sg13g2_xnor2_1 _18434_ (.Y(_02489_),
    .A(_00147_),
    .B(_06921_));
 sg13g2_nor2_1 _18435_ (.A(net5830),
    .B(_02489_),
    .Y(_02490_));
 sg13g2_a21oi_1 _18436_ (.A1(net5830),
    .A2(\TRNG.hash[163] ),
    .Y(_02491_),
    .B1(_02490_));
 sg13g2_nor2_1 _18437_ (.A(net5097),
    .B(net5177),
    .Y(_02492_));
 sg13g2_nand2_1 _18438_ (.Y(_02493_),
    .A(net5089),
    .B(net5350));
 sg13g2_o21ai_1 _18439_ (.B1(net5465),
    .Y(_02494_),
    .A1(net3630),
    .A2(net4920));
 sg13g2_a21oi_1 _18440_ (.A1(net4956),
    .A2(_02491_),
    .Y(_01064_),
    .B1(_02494_));
 sg13g2_xnor2_1 _18441_ (.Y(_02495_),
    .A(_04234_),
    .B(_02488_));
 sg13g2_nor2_1 _18442_ (.A(net5830),
    .B(_02495_),
    .Y(_02496_));
 sg13g2_a21oi_1 _18443_ (.A1(\TRNG.hash[164] ),
    .A2(net5830),
    .Y(_02497_),
    .B1(_02496_));
 sg13g2_a221oi_1 _18444_ (.B2(net4956),
    .C1(net5521),
    .B1(_02497_),
    .A1(_04234_),
    .Y(_01065_),
    .A2(net4934));
 sg13g2_or2_1 _18445_ (.X(_02498_),
    .B(_06922_),
    .A(net3643));
 sg13g2_a21o_1 _18446_ (.A2(_02498_),
    .A1(_06923_),
    .B1(net5830),
    .X(_02499_));
 sg13g2_a21oi_1 _18447_ (.A1(\TRNG.hash[165] ),
    .A2(net5827),
    .Y(_02500_),
    .B1(net4939));
 sg13g2_o21ai_1 _18448_ (.B1(net5464),
    .Y(_02501_),
    .A1(\TRNG.hash[133] ),
    .A2(net4919));
 sg13g2_a21oi_1 _18449_ (.A1(_02499_),
    .A2(_02500_),
    .Y(_01066_),
    .B1(_02501_));
 sg13g2_xor2_1 _18450_ (.B(_06934_),
    .A(_00148_),
    .X(_02502_));
 sg13g2_nor2_1 _18451_ (.A(net5831),
    .B(_02502_),
    .Y(_02503_));
 sg13g2_a21oi_1 _18452_ (.A1(\TRNG.hash[168] ),
    .A2(net5831),
    .Y(_02504_),
    .B1(_02503_));
 sg13g2_o21ai_1 _18453_ (.B1(net5464),
    .Y(_02505_),
    .A1(net3515),
    .A2(net4920));
 sg13g2_a21oi_1 _18454_ (.A1(net4956),
    .A2(_02504_),
    .Y(_01067_),
    .B1(_02505_));
 sg13g2_xor2_1 _18455_ (.B(_06939_),
    .A(_00136_),
    .X(_02506_));
 sg13g2_nor2_1 _18456_ (.A(net5829),
    .B(_02506_),
    .Y(_02507_));
 sg13g2_a21oi_1 _18457_ (.A1(net5829),
    .A2(\TRNG.hash[170] ),
    .Y(_02508_),
    .B1(_02507_));
 sg13g2_o21ai_1 _18458_ (.B1(net5464),
    .Y(_02509_),
    .A1(net3665),
    .A2(net4920));
 sg13g2_a21oi_1 _18459_ (.A1(net4953),
    .A2(_02508_),
    .Y(_01068_),
    .B1(_02509_));
 sg13g2_xor2_1 _18460_ (.B(_06941_),
    .A(_00138_),
    .X(_02510_));
 sg13g2_a21oi_1 _18461_ (.A1(\TRNG.hash[172] ),
    .A2(net5836),
    .Y(_02511_),
    .B1(net4939));
 sg13g2_o21ai_1 _18462_ (.B1(_02511_),
    .Y(_02512_),
    .A1(net5829),
    .A2(_02510_));
 sg13g2_o21ai_1 _18463_ (.B1(_02512_),
    .Y(_02513_),
    .A1(net3624),
    .A2(net4920));
 sg13g2_nor2_1 _18464_ (.A(net5520),
    .B(net3625),
    .Y(_01069_));
 sg13g2_a21o_1 _18465_ (.A2(_06946_),
    .A1(_00138_),
    .B1(_04233_),
    .X(_02514_));
 sg13g2_a21o_1 _18466_ (.A2(_02514_),
    .A1(_06947_),
    .B1(net5829),
    .X(_02515_));
 sg13g2_a21oi_1 _18467_ (.A1(\TRNG.hash[173] ),
    .A2(net5829),
    .Y(_02516_),
    .B1(net4939));
 sg13g2_a221oi_1 _18468_ (.B2(_02516_),
    .C1(net5520),
    .B1(_02515_),
    .A1(_04233_),
    .Y(_01070_),
    .A2(net4934));
 sg13g2_xnor2_1 _18469_ (.Y(_02517_),
    .A(net3842),
    .B(_06947_));
 sg13g2_nand2_1 _18470_ (.Y(_02518_),
    .A(net5485),
    .B(_02517_));
 sg13g2_a21oi_1 _18471_ (.A1(\TRNG.hash[174] ),
    .A2(net5832),
    .Y(_02519_),
    .B1(net4940));
 sg13g2_a221oi_1 _18472_ (.B2(_02519_),
    .C1(net5520),
    .B1(_02518_),
    .A1(_04232_),
    .Y(_01071_),
    .A2(net4934));
 sg13g2_o21ai_1 _18473_ (.B1(\TRNG.hash[143] ),
    .Y(_02520_),
    .A1(\TRNG.hash[142] ),
    .A2(_06947_));
 sg13g2_nor2b_1 _18474_ (.A(_06948_),
    .B_N(_02520_),
    .Y(_02521_));
 sg13g2_a21oi_1 _18475_ (.A1(\TRNG.hash[175] ),
    .A2(net5832),
    .Y(_02522_),
    .B1(net4939));
 sg13g2_o21ai_1 _18476_ (.B1(_02522_),
    .Y(_02523_),
    .A1(net5832),
    .A2(_02521_));
 sg13g2_o21ai_1 _18477_ (.B1(_02523_),
    .Y(_02524_),
    .A1(net3759),
    .A2(net4920));
 sg13g2_nor2_1 _18478_ (.A(net5520),
    .B(_02524_),
    .Y(_01072_));
 sg13g2_xnor2_1 _18479_ (.Y(_02525_),
    .A(\TRNG.hash[144] ),
    .B(_06948_));
 sg13g2_a21oi_1 _18480_ (.A1(net5832),
    .A2(\TRNG.hash[176] ),
    .Y(_02526_),
    .B1(net4940));
 sg13g2_o21ai_1 _18481_ (.B1(_02526_),
    .Y(_02527_),
    .A1(net5832),
    .A2(_02525_));
 sg13g2_o21ai_1 _18482_ (.B1(_02527_),
    .Y(_02528_),
    .A1(net3718),
    .A2(net4920));
 sg13g2_nor2_1 _18483_ (.A(net5522),
    .B(net3719),
    .Y(_01073_));
 sg13g2_nor2_1 _18484_ (.A(_04231_),
    .B(_06949_),
    .Y(_02529_));
 sg13g2_o21ai_1 _18485_ (.B1(net5484),
    .Y(_02530_),
    .A1(_06950_),
    .A2(_02529_));
 sg13g2_a21oi_1 _18486_ (.A1(\TRNG.hash[177] ),
    .A2(net5832),
    .Y(_02531_),
    .B1(net4940));
 sg13g2_a221oi_1 _18487_ (.B2(_02531_),
    .C1(net5522),
    .B1(_02530_),
    .A1(_04231_),
    .Y(_01074_),
    .A2(net4935));
 sg13g2_xnor2_1 _18488_ (.Y(_02532_),
    .A(_04230_),
    .B(_06950_));
 sg13g2_nand2_1 _18489_ (.Y(_02533_),
    .A(net5484),
    .B(_02532_));
 sg13g2_a21oi_1 _18490_ (.A1(\TRNG.hash[178] ),
    .A2(net5832),
    .Y(_02534_),
    .B1(net4940));
 sg13g2_a221oi_1 _18491_ (.B2(_02534_),
    .C1(net5521),
    .B1(_02533_),
    .A1(_04230_),
    .Y(_01075_),
    .A2(net4935));
 sg13g2_a21oi_1 _18492_ (.A1(_04230_),
    .A2(_06950_),
    .Y(_02535_),
    .B1(_04229_));
 sg13g2_o21ai_1 _18493_ (.B1(net5484),
    .Y(_02536_),
    .A1(_06951_),
    .A2(_02535_));
 sg13g2_a21oi_1 _18494_ (.A1(\TRNG.hash[179] ),
    .A2(net5833),
    .Y(_02537_),
    .B1(net4940));
 sg13g2_a221oi_1 _18495_ (.B2(_02537_),
    .C1(net5521),
    .B1(_02536_),
    .A1(_04229_),
    .Y(_01076_),
    .A2(net4934));
 sg13g2_xnor2_1 _18496_ (.Y(_02538_),
    .A(net3645),
    .B(_06959_));
 sg13g2_nand2_1 _18497_ (.Y(_02539_),
    .A(net5489),
    .B(_02538_));
 sg13g2_a21oi_1 _18498_ (.A1(\TRNG.hash[182] ),
    .A2(net5842),
    .Y(_02540_),
    .B1(net4942));
 sg13g2_o21ai_1 _18499_ (.B1(net5467),
    .Y(_02541_),
    .A1(\TRNG.hash[150] ),
    .A2(net4923));
 sg13g2_a21oi_1 _18500_ (.A1(_02539_),
    .A2(_02540_),
    .Y(_01077_),
    .B1(_02541_));
 sg13g2_xor2_1 _18501_ (.B(_06961_),
    .A(_00141_),
    .X(_02542_));
 sg13g2_a21oi_1 _18502_ (.A1(net5841),
    .A2(\TRNG.hash[184] ),
    .Y(_02543_),
    .B1(net4942));
 sg13g2_o21ai_1 _18503_ (.B1(_02543_),
    .Y(_02544_),
    .A1(net5841),
    .A2(_02542_));
 sg13g2_o21ai_1 _18504_ (.B1(_02544_),
    .Y(_02545_),
    .A1(net3699),
    .A2(net4923));
 sg13g2_nor2_1 _18505_ (.A(net5524),
    .B(net3700),
    .Y(_01078_));
 sg13g2_xnor2_1 _18506_ (.Y(_02546_),
    .A(_00143_),
    .B(_06968_));
 sg13g2_a21oi_1 _18507_ (.A1(\TRNG.hash[186] ),
    .A2(net5833),
    .Y(_02547_),
    .B1(net4942));
 sg13g2_o21ai_1 _18508_ (.B1(_02547_),
    .Y(_02548_),
    .A1(net5832),
    .A2(_02546_));
 sg13g2_o21ai_1 _18509_ (.B1(_02548_),
    .Y(_02549_),
    .A1(net3712),
    .A2(net4923));
 sg13g2_nor2_1 _18510_ (.A(net5521),
    .B(net3713),
    .Y(_01079_));
 sg13g2_xor2_1 _18511_ (.B(_06982_),
    .A(_00145_),
    .X(_02550_));
 sg13g2_a21oi_1 _18512_ (.A1(\TRNG.hash[189] ),
    .A2(net5843),
    .Y(_02551_),
    .B1(net4942));
 sg13g2_o21ai_1 _18513_ (.B1(_02551_),
    .Y(_02552_),
    .A1(net5843),
    .A2(_02550_));
 sg13g2_o21ai_1 _18514_ (.B1(_02552_),
    .Y(_02553_),
    .A1(net3681),
    .A2(net4923));
 sg13g2_nor2_1 _18515_ (.A(net5524),
    .B(net3682),
    .Y(_01080_));
 sg13g2_o21ai_1 _18516_ (.B1(\TRNG.hash[158] ),
    .Y(_02554_),
    .A1(\TRNG.hash[157] ),
    .A2(_06983_));
 sg13g2_xnor2_1 _18517_ (.Y(_02555_),
    .A(\TRNG.hash[159] ),
    .B(_02554_));
 sg13g2_a21oi_1 _18518_ (.A1(net5842),
    .A2(\TRNG.hash[191] ),
    .Y(_02556_),
    .B1(net4943));
 sg13g2_o21ai_1 _18519_ (.B1(_02556_),
    .Y(_02557_),
    .A1(net5842),
    .A2(_02555_));
 sg13g2_o21ai_1 _18520_ (.B1(net5467),
    .Y(_02558_),
    .A1(net3772),
    .A2(net4923));
 sg13g2_nor2b_1 _18521_ (.A(_02558_),
    .B_N(_02557_),
    .Y(_01081_));
 sg13g2_a21oi_1 _18522_ (.A1(_04227_),
    .A2(_04228_),
    .Y(_01083_),
    .B1(_06877_));
 sg13g2_xnor2_1 _18523_ (.Y(_02559_),
    .A(_08270_),
    .B(_08273_));
 sg13g2_o21ai_1 _18524_ (.B1(net4956),
    .Y(_02560_),
    .A1(net5830),
    .A2(_04379_));
 sg13g2_a21oi_1 _18525_ (.A1(net5830),
    .A2(_02559_),
    .Y(_02561_),
    .B1(_02560_));
 sg13g2_o21ai_1 _18526_ (.B1(net5464),
    .Y(_02562_),
    .A1(net5570),
    .A2(net4919));
 sg13g2_nor2_1 _18527_ (.A(_02561_),
    .B(_02562_),
    .Y(_01084_));
 sg13g2_nand2_1 _18528_ (.Y(_02563_),
    .A(_08275_),
    .B(_08276_));
 sg13g2_nand3_1 _18529_ (.B(_08277_),
    .C(_02563_),
    .A(net5828),
    .Y(_02564_));
 sg13g2_nand2_1 _18530_ (.Y(_02565_),
    .A(net5569),
    .B(net5570));
 sg13g2_a21oi_1 _18531_ (.A1(_08294_),
    .A2(_02565_),
    .Y(_02566_),
    .B1(net5828));
 sg13g2_nor2_1 _18532_ (.A(net4939),
    .B(_02566_),
    .Y(_02567_));
 sg13g2_o21ai_1 _18533_ (.B1(net5464),
    .Y(_02568_),
    .A1(net5569),
    .A2(net4919));
 sg13g2_a21oi_1 _18534_ (.A1(_02564_),
    .A2(_02567_),
    .Y(_01085_),
    .B1(_02568_));
 sg13g2_xnor2_1 _18535_ (.Y(_02569_),
    .A(_08277_),
    .B(_08279_));
 sg13g2_xor2_1 _18536_ (.B(_08294_),
    .A(net5568),
    .X(_02570_));
 sg13g2_o21ai_1 _18537_ (.B1(net4953),
    .Y(_02571_),
    .A1(net5828),
    .A2(_02570_));
 sg13g2_a21oi_1 _18538_ (.A1(net5828),
    .A2(_02569_),
    .Y(_02572_),
    .B1(_02571_));
 sg13g2_o21ai_1 _18539_ (.B1(net5464),
    .Y(_02573_),
    .A1(net5568),
    .A2(net4919));
 sg13g2_nor2_1 _18540_ (.A(_02572_),
    .B(_02573_),
    .Y(_01086_));
 sg13g2_xnor2_1 _18541_ (.Y(_02574_),
    .A(_08336_),
    .B(_08338_));
 sg13g2_xor2_1 _18542_ (.B(_08312_),
    .A(net3767),
    .X(_02575_));
 sg13g2_o21ai_1 _18543_ (.B1(net4953),
    .Y(_02576_),
    .A1(net5820),
    .A2(_02575_));
 sg13g2_a21oi_1 _18544_ (.A1(net5820),
    .A2(_02574_),
    .Y(_02577_),
    .B1(_02576_));
 sg13g2_o21ai_1 _18545_ (.B1(net5462),
    .Y(_02578_),
    .A1(net5567),
    .A2(net4916));
 sg13g2_nor2_1 _18546_ (.A(_02577_),
    .B(_02578_),
    .Y(_01087_));
 sg13g2_o21ai_1 _18547_ (.B1(net5820),
    .Y(_02579_),
    .A1(_08339_),
    .A2(_08340_));
 sg13g2_a21o_1 _18548_ (.A2(_08340_),
    .A1(_08339_),
    .B1(_02579_),
    .X(_02580_));
 sg13g2_xnor2_1 _18549_ (.Y(_02581_),
    .A(net5566),
    .B(_08356_));
 sg13g2_a21oi_1 _18550_ (.A1(net5483),
    .A2(_02581_),
    .Y(_02582_),
    .B1(net4936));
 sg13g2_o21ai_1 _18551_ (.B1(net5462),
    .Y(_02583_),
    .A1(net5566),
    .A2(net4916));
 sg13g2_a21oi_1 _18552_ (.A1(_02580_),
    .A2(_02582_),
    .Y(_01088_),
    .B1(_02583_));
 sg13g2_nand2_1 _18553_ (.Y(_02584_),
    .A(_08399_),
    .B(_08400_));
 sg13g2_a21oi_1 _18554_ (.A1(_08401_),
    .A2(_02584_),
    .Y(_02585_),
    .B1(net5483));
 sg13g2_o21ai_1 _18555_ (.B1(_02585_),
    .Y(_02586_),
    .A1(_08401_),
    .A2(_02584_));
 sg13g2_xnor2_1 _18556_ (.Y(_02587_),
    .A(net3716),
    .B(_08375_));
 sg13g2_a21oi_1 _18557_ (.A1(net5483),
    .A2(_02587_),
    .Y(_02588_),
    .B1(net4936));
 sg13g2_o21ai_1 _18558_ (.B1(net5461),
    .Y(_02589_),
    .A1(net5565),
    .A2(net4915));
 sg13g2_a21oi_1 _18559_ (.A1(_02586_),
    .A2(_02588_),
    .Y(_01089_),
    .B1(_02589_));
 sg13g2_xor2_1 _18560_ (.B(_08404_),
    .A(_08395_),
    .X(_02590_));
 sg13g2_xor2_1 _18561_ (.B(_08422_),
    .A(net5564),
    .X(_02591_));
 sg13g2_o21ai_1 _18562_ (.B1(net4953),
    .Y(_02592_),
    .A1(net5816),
    .A2(_02591_));
 sg13g2_a21oi_1 _18563_ (.A1(net5816),
    .A2(_02590_),
    .Y(_02593_),
    .B1(_02592_));
 sg13g2_o21ai_1 _18564_ (.B1(net5461),
    .Y(_02594_),
    .A1(net5564),
    .A2(net4915));
 sg13g2_nor2_1 _18565_ (.A(_02593_),
    .B(_02594_),
    .Y(_01090_));
 sg13g2_nor2_1 _18566_ (.A(_08439_),
    .B(_08447_),
    .Y(_02595_));
 sg13g2_xnor2_1 _18567_ (.Y(_02596_),
    .A(_08507_),
    .B(_02595_));
 sg13g2_xor2_1 _18568_ (.B(_08520_),
    .A(net3833),
    .X(_02597_));
 sg13g2_o21ai_1 _18569_ (.B1(net4953),
    .Y(_02598_),
    .A1(net5818),
    .A2(_02597_));
 sg13g2_a21oi_1 _18570_ (.A1(net5817),
    .A2(_02596_),
    .Y(_02599_),
    .B1(_02598_));
 sg13g2_o21ai_1 _18571_ (.B1(net5461),
    .Y(_02600_),
    .A1(net5563),
    .A2(net4916));
 sg13g2_nor2_1 _18572_ (.A(_02599_),
    .B(_02600_),
    .Y(_01091_));
 sg13g2_a21o_1 _18573_ (.A2(_08508_),
    .A1(_08445_),
    .B1(_08511_),
    .X(_02601_));
 sg13g2_nand2b_1 _18574_ (.Y(_02602_),
    .B(_02601_),
    .A_N(_08496_));
 sg13g2_xnor2_1 _18575_ (.Y(_02603_),
    .A(_08496_),
    .B(_02601_));
 sg13g2_o21ai_1 _18576_ (.B1(net3924),
    .Y(_02604_),
    .A1(net5563),
    .A2(_08520_));
 sg13g2_nor2_1 _18577_ (.A(net5562),
    .B(_02604_),
    .Y(_02605_));
 sg13g2_xor2_1 _18578_ (.B(_02604_),
    .A(net5562),
    .X(_02606_));
 sg13g2_o21ai_1 _18579_ (.B1(net4953),
    .Y(_02607_),
    .A1(net5818),
    .A2(_02606_));
 sg13g2_a21oi_1 _18580_ (.A1(net5823),
    .A2(_02603_),
    .Y(_02608_),
    .B1(_02607_));
 sg13g2_o21ai_1 _18581_ (.B1(net5461),
    .Y(_02609_),
    .A1(net5562),
    .A2(net4917));
 sg13g2_nor2_1 _18582_ (.A(_02608_),
    .B(_02609_),
    .Y(_01092_));
 sg13g2_a21oi_1 _18583_ (.A1(_08494_),
    .A2(_02602_),
    .Y(_02610_),
    .B1(_08501_));
 sg13g2_nand3_1 _18584_ (.B(_08501_),
    .C(_02602_),
    .A(_08494_),
    .Y(_02611_));
 sg13g2_nor2_1 _18585_ (.A(net5483),
    .B(_02610_),
    .Y(_02612_));
 sg13g2_xor2_1 _18586_ (.B(_02605_),
    .A(net5561),
    .X(_02613_));
 sg13g2_a221oi_1 _18587_ (.B2(net5483),
    .C1(net4937),
    .B1(_02613_),
    .A1(_02611_),
    .Y(_02614_),
    .A2(_02612_));
 sg13g2_o21ai_1 _18588_ (.B1(net5468),
    .Y(_02615_),
    .A1(net5561),
    .A2(net4917));
 sg13g2_nor2_1 _18589_ (.A(_02614_),
    .B(_02615_),
    .Y(_01093_));
 sg13g2_o21ai_1 _18590_ (.B1(net5823),
    .Y(_02616_),
    .A1(_08514_),
    .A2(_08516_));
 sg13g2_a21oi_1 _18591_ (.A1(_08514_),
    .A2(_08516_),
    .Y(_02617_),
    .B1(_02616_));
 sg13g2_xnor2_1 _18592_ (.Y(_02618_),
    .A(_04226_),
    .B(_08522_));
 sg13g2_o21ai_1 _18593_ (.B1(net4954),
    .Y(_02619_),
    .A1(net5823),
    .A2(_02618_));
 sg13g2_o21ai_1 _18594_ (.B1(net5463),
    .Y(_02620_),
    .A1(_02617_),
    .A2(_02619_));
 sg13g2_a21oi_1 _18595_ (.A1(_04226_),
    .A2(net4934),
    .Y(_01094_),
    .B1(_02620_));
 sg13g2_nor2_1 _18596_ (.A(_08535_),
    .B(_08541_),
    .Y(_02621_));
 sg13g2_xnor2_1 _18597_ (.Y(_02622_),
    .A(_08568_),
    .B(_02621_));
 sg13g2_xor2_1 _18598_ (.B(_08543_),
    .A(net3795),
    .X(_02623_));
 sg13g2_o21ai_1 _18599_ (.B1(net4954),
    .Y(_02624_),
    .A1(net5825),
    .A2(_02623_));
 sg13g2_a21oi_1 _18600_ (.A1(net5825),
    .A2(_02622_),
    .Y(_02625_),
    .B1(_02624_));
 sg13g2_o21ai_1 _18601_ (.B1(net5463),
    .Y(_02626_),
    .A1(net5560),
    .A2(net4921));
 sg13g2_nor2_1 _18602_ (.A(_02625_),
    .B(_02626_),
    .Y(_01095_));
 sg13g2_nor2_1 _18603_ (.A(_08649_),
    .B(_08651_),
    .Y(_02627_));
 sg13g2_xor2_1 _18604_ (.B(_02627_),
    .A(_08680_),
    .X(_02628_));
 sg13g2_xnor2_1 _18605_ (.Y(_02629_),
    .A(net3741),
    .B(_08653_));
 sg13g2_o21ai_1 _18606_ (.B1(net4954),
    .Y(_02630_),
    .A1(net5838),
    .A2(_02629_));
 sg13g2_a21oi_1 _18607_ (.A1(net5837),
    .A2(_02628_),
    .Y(_02631_),
    .B1(_02630_));
 sg13g2_o21ai_1 _18608_ (.B1(net5466),
    .Y(_02632_),
    .A1(net5559),
    .A2(net4922));
 sg13g2_nor2_1 _18609_ (.A(_02631_),
    .B(_02632_),
    .Y(_01096_));
 sg13g2_a21oi_1 _18610_ (.A1(_08674_),
    .A2(_08682_),
    .Y(_02633_),
    .B1(_08673_));
 sg13g2_a21oi_1 _18611_ (.A1(_08700_),
    .A2(_02633_),
    .Y(_02634_),
    .B1(net5486));
 sg13g2_o21ai_1 _18612_ (.B1(_02634_),
    .Y(_02635_),
    .A1(_08700_),
    .A2(_02633_));
 sg13g2_xnor2_1 _18613_ (.Y(_02636_),
    .A(net3783),
    .B(_08685_));
 sg13g2_a21oi_1 _18614_ (.A1(net5486),
    .A2(_02636_),
    .Y(_02637_),
    .B1(net4941));
 sg13g2_o21ai_1 _18615_ (.B1(net5463),
    .Y(_02638_),
    .A1(net5558),
    .A2(net4921));
 sg13g2_a21oi_1 _18616_ (.A1(_02635_),
    .A2(_02637_),
    .Y(_01097_),
    .B1(_02638_));
 sg13g2_a21oi_1 _18617_ (.A1(_08707_),
    .A2(_08718_),
    .Y(_02639_),
    .B1(_08717_));
 sg13g2_xnor2_1 _18618_ (.Y(_02640_),
    .A(_08746_),
    .B(_02639_));
 sg13g2_xor2_1 _18619_ (.B(_08723_),
    .A(net3788),
    .X(_02641_));
 sg13g2_o21ai_1 _18620_ (.B1(net4953),
    .Y(_02642_),
    .A1(net5838),
    .A2(_02641_));
 sg13g2_a21oi_1 _18621_ (.A1(net5840),
    .A2(_02640_),
    .Y(_02643_),
    .B1(_02642_));
 sg13g2_o21ai_1 _18622_ (.B1(net5466),
    .Y(_02644_),
    .A1(net5557),
    .A2(net4921));
 sg13g2_nor2_1 _18623_ (.A(_02643_),
    .B(_02644_),
    .Y(_01098_));
 sg13g2_xor2_1 _18624_ (.B(_08751_),
    .A(_08749_),
    .X(_02645_));
 sg13g2_xnor2_1 _18625_ (.Y(_02646_),
    .A(net5556),
    .B(_08763_));
 sg13g2_a21oi_1 _18626_ (.A1(net5487),
    .A2(_02646_),
    .Y(_02647_),
    .B1(net4941));
 sg13g2_o21ai_1 _18627_ (.B1(_02647_),
    .Y(_02648_),
    .A1(net5487),
    .A2(_02645_));
 sg13g2_o21ai_1 _18628_ (.B1(net5466),
    .Y(_02649_),
    .A1(net5556),
    .A2(net4922));
 sg13g2_nor2b_1 _18629_ (.A(_02649_),
    .B_N(_02648_),
    .Y(_01099_));
 sg13g2_or2_1 _18630_ (.X(_02650_),
    .B(net5571),
    .A(\TRNG.hash[192] ));
 sg13g2_nand3_1 _18631_ (.B(_08186_),
    .C(_02650_),
    .A(net5484),
    .Y(_02651_));
 sg13g2_a21oi_1 _18632_ (.A1(net5830),
    .A2(_04379_),
    .Y(_02652_),
    .B1(net5097));
 sg13g2_a21oi_1 _18633_ (.A1(_02651_),
    .A2(_02652_),
    .Y(_01100_),
    .B1(net5521));
 sg13g2_nand3_1 _18634_ (.B(\TRNG.hash[192] ),
    .C(\TRNG.hash[193] ),
    .A(net3703),
    .Y(_02653_));
 sg13g2_a21oi_1 _18635_ (.A1(_08188_),
    .A2(_02653_),
    .Y(_02654_),
    .B1(net5827));
 sg13g2_a21oi_1 _18636_ (.A1(net5568),
    .A2(net5827),
    .Y(_02655_),
    .B1(_02654_));
 sg13g2_o21ai_1 _18637_ (.B1(net5462),
    .Y(_02656_),
    .A1(net3567),
    .A2(net4919));
 sg13g2_a21oi_1 _18638_ (.A1(net4953),
    .A2(_02655_),
    .Y(_01101_),
    .B1(_02656_));
 sg13g2_or3_1 _18639_ (.A(_04225_),
    .B(_08194_),
    .C(_08200_),
    .X(_02657_));
 sg13g2_a21o_1 _18640_ (.A2(_02657_),
    .A1(_08204_),
    .B1(net5820),
    .X(_02658_));
 sg13g2_a21oi_1 _18641_ (.A1(net5820),
    .A2(\TRNG.hash[231] ),
    .Y(_02659_),
    .B1(net4938));
 sg13g2_a221oi_1 _18642_ (.B2(_02659_),
    .C1(net5518),
    .B1(_02658_),
    .A1(_04225_),
    .Y(_01102_),
    .A2(net4934));
 sg13g2_xnor2_1 _18643_ (.Y(_02660_),
    .A(net3474),
    .B(_08207_));
 sg13g2_nand2_1 _18644_ (.Y(_02661_),
    .A(net5483),
    .B(_02660_));
 sg13g2_a21oi_1 _18645_ (.A1(net5565),
    .A2(net5816),
    .Y(_02662_),
    .B1(net4936));
 sg13g2_o21ai_1 _18646_ (.B1(net5461),
    .Y(_02663_),
    .A1(\TRNG.hash[201] ),
    .A2(net4915));
 sg13g2_a21oi_1 _18647_ (.A1(_02661_),
    .A2(_02662_),
    .Y(_01103_),
    .B1(_02663_));
 sg13g2_o21ai_1 _18648_ (.B1(net3474),
    .Y(_02664_),
    .A1(\TRNG.hash[201] ),
    .A2(_08207_));
 sg13g2_nor2_1 _18649_ (.A(\TRNG.hash[202] ),
    .B(_02664_),
    .Y(_02665_));
 sg13g2_and2_1 _18650_ (.A(\TRNG.hash[202] ),
    .B(_02664_),
    .X(_02666_));
 sg13g2_o21ai_1 _18651_ (.B1(net5483),
    .Y(_02667_),
    .A1(_02665_),
    .A2(_02666_));
 sg13g2_a21oi_1 _18652_ (.A1(net5564),
    .A2(net5816),
    .Y(_02668_),
    .B1(net4936));
 sg13g2_o21ai_1 _18653_ (.B1(net5461),
    .Y(_02669_),
    .A1(net3760),
    .A2(net4915));
 sg13g2_a21oi_1 _18654_ (.A1(_02667_),
    .A2(_02668_),
    .Y(_01104_),
    .B1(_02669_));
 sg13g2_xnor2_1 _18655_ (.Y(_02670_),
    .A(\TRNG.hash[203] ),
    .B(_02665_));
 sg13g2_a21oi_1 _18656_ (.A1(net5816),
    .A2(\TRNG.hash[235] ),
    .Y(_02671_),
    .B1(net4936));
 sg13g2_o21ai_1 _18657_ (.B1(_02671_),
    .Y(_02672_),
    .A1(net5816),
    .A2(_02670_));
 sg13g2_o21ai_1 _18658_ (.B1(_02672_),
    .Y(_02673_),
    .A1(net3845),
    .A2(net4915));
 sg13g2_nor2_1 _18659_ (.A(net5518),
    .B(_02673_),
    .Y(_01105_));
 sg13g2_a21oi_1 _18660_ (.A1(net3437),
    .A2(_08211_),
    .Y(_02674_),
    .B1(net5817));
 sg13g2_o21ai_1 _18661_ (.B1(_02674_),
    .Y(_02675_),
    .A1(net3437),
    .A2(_08211_));
 sg13g2_a21oi_1 _18662_ (.A1(net5563),
    .A2(net5817),
    .Y(_02676_),
    .B1(net4936));
 sg13g2_o21ai_1 _18663_ (.B1(net5461),
    .Y(_02677_),
    .A1(\TRNG.hash[205] ),
    .A2(net4915));
 sg13g2_a21oi_1 _18664_ (.A1(_02675_),
    .A2(_02676_),
    .Y(_01106_),
    .B1(_02677_));
 sg13g2_xnor2_1 _18665_ (.Y(_02678_),
    .A(\TRNG.hash[207] ),
    .B(_08216_));
 sg13g2_a21oi_1 _18666_ (.A1(net5561),
    .A2(net5822),
    .Y(_02679_),
    .B1(net4937));
 sg13g2_o21ai_1 _18667_ (.B1(_02679_),
    .Y(_02680_),
    .A1(net5822),
    .A2(_02678_));
 sg13g2_o21ai_1 _18668_ (.B1(_02680_),
    .Y(_02681_),
    .A1(net3832),
    .A2(net4917));
 sg13g2_nor2_1 _18669_ (.A(net5518),
    .B(_02681_),
    .Y(_01107_));
 sg13g2_nor2_1 _18670_ (.A(_04380_),
    .B(_08221_),
    .Y(_02682_));
 sg13g2_and2_1 _18671_ (.A(_04380_),
    .B(_08221_),
    .X(_02683_));
 sg13g2_o21ai_1 _18672_ (.B1(net5485),
    .Y(_02684_),
    .A1(_02682_),
    .A2(_02683_));
 sg13g2_a21oi_1 _18673_ (.A1(\TRNG.hash[240] ),
    .A2(net5823),
    .Y(_02685_),
    .B1(net4937));
 sg13g2_o21ai_1 _18674_ (.B1(net5463),
    .Y(_02686_),
    .A1(net3636),
    .A2(net4917));
 sg13g2_a21oi_1 _18675_ (.A1(_02684_),
    .A2(_02685_),
    .Y(_01108_),
    .B1(_02686_));
 sg13g2_xnor2_1 _18676_ (.Y(_02687_),
    .A(\TRNG.hash[209] ),
    .B(_02682_));
 sg13g2_a21oi_1 _18677_ (.A1(net5823),
    .A2(net5884),
    .Y(_02688_),
    .B1(net4937));
 sg13g2_o21ai_1 _18678_ (.B1(_02688_),
    .Y(_02689_),
    .A1(net5822),
    .A2(_02687_));
 sg13g2_o21ai_1 _18679_ (.B1(_02689_),
    .Y(_02690_),
    .A1(net3844),
    .A2(net4917));
 sg13g2_nor2_1 _18680_ (.A(net5519),
    .B(_02690_),
    .Y(_01109_));
 sg13g2_xnor2_1 _18681_ (.Y(_02691_),
    .A(\TRNG.hash[210] ),
    .B(_08222_));
 sg13g2_a21oi_1 _18682_ (.A1(net5824),
    .A2(net5883),
    .Y(_02692_),
    .B1(net4937));
 sg13g2_o21ai_1 _18683_ (.B1(_02692_),
    .Y(_02693_),
    .A1(net5824),
    .A2(_02691_));
 sg13g2_o21ai_1 _18684_ (.B1(_02693_),
    .Y(_02694_),
    .A1(net3792),
    .A2(net4918));
 sg13g2_nor2_1 _18685_ (.A(net5519),
    .B(_02694_),
    .Y(_01110_));
 sg13g2_xnor2_1 _18686_ (.Y(_02695_),
    .A(net3530),
    .B(_08228_));
 sg13g2_nand2_1 _18687_ (.Y(_02696_),
    .A(net5489),
    .B(_02695_));
 sg13g2_a21oi_1 _18688_ (.A1(net5841),
    .A2(net5881),
    .Y(_02697_),
    .B1(net4942));
 sg13g2_a221oi_1 _18689_ (.B2(_02697_),
    .C1(net5524),
    .B1(_02696_),
    .A1(_04224_),
    .Y(_01111_),
    .A2(net4935));
 sg13g2_and2_1 _18690_ (.A(net3828),
    .B(_08232_),
    .X(_02698_));
 sg13g2_o21ai_1 _18691_ (.B1(net5488),
    .Y(_02699_),
    .A1(_08233_),
    .A2(_02698_));
 sg13g2_a21oi_1 _18692_ (.A1(net5841),
    .A2(\TRNG.hash[246] ),
    .Y(_02700_),
    .B1(net4942));
 sg13g2_a221oi_1 _18693_ (.B2(_02700_),
    .C1(net5523),
    .B1(_02699_),
    .A1(_04223_),
    .Y(_01112_),
    .A2(net4935));
 sg13g2_and3_1 _18694_ (.X(_02701_),
    .A(\TRNG.hash[216] ),
    .B(\TRNG.hash[215] ),
    .C(_08237_));
 sg13g2_o21ai_1 _18695_ (.B1(net5486),
    .Y(_02702_),
    .A1(_08238_),
    .A2(_02701_));
 sg13g2_a21oi_1 _18696_ (.A1(net5839),
    .A2(net5879),
    .Y(_02703_),
    .B1(net4942));
 sg13g2_o21ai_1 _18697_ (.B1(net5466),
    .Y(_02704_),
    .A1(net3786),
    .A2(net4924));
 sg13g2_a21oi_1 _18698_ (.A1(_02702_),
    .A2(_02703_),
    .Y(_01113_),
    .B1(_02704_));
 sg13g2_xnor2_1 _18699_ (.Y(_02705_),
    .A(\TRNG.hash[217] ),
    .B(_08238_));
 sg13g2_a21oi_1 _18700_ (.A1(net5559),
    .A2(net5837),
    .Y(_02706_),
    .B1(net4941));
 sg13g2_o21ai_1 _18701_ (.B1(_02706_),
    .Y(_02707_),
    .A1(net5837),
    .A2(_02705_));
 sg13g2_o21ai_1 _18702_ (.B1(_02707_),
    .Y(_02708_),
    .A1(net3814),
    .A2(net4921));
 sg13g2_nor2_1 _18703_ (.A(net5523),
    .B(_02708_),
    .Y(_01114_));
 sg13g2_xnor2_1 _18704_ (.Y(_02709_),
    .A(net3476),
    .B(_08240_));
 sg13g2_nand2_1 _18705_ (.Y(_02710_),
    .A(net5486),
    .B(_02709_));
 sg13g2_a21oi_1 _18706_ (.A1(net5558),
    .A2(net5837),
    .Y(_02711_),
    .B1(net4941));
 sg13g2_o21ai_1 _18707_ (.B1(net5463),
    .Y(_02712_),
    .A1(\TRNG.hash[219] ),
    .A2(net4921));
 sg13g2_a21oi_1 _18708_ (.A1(_02710_),
    .A2(_02711_),
    .Y(_01115_),
    .B1(_02712_));
 sg13g2_and2_1 _18709_ (.A(\TRNG.hash[220] ),
    .B(_08244_),
    .X(_02713_));
 sg13g2_o21ai_1 _18710_ (.B1(net5487),
    .Y(_02714_),
    .A1(_08245_),
    .A2(_02713_));
 sg13g2_a21oi_1 _18711_ (.A1(net5838),
    .A2(net5877),
    .Y(_02715_),
    .B1(net4943));
 sg13g2_o21ai_1 _18712_ (.B1(net5466),
    .Y(_02716_),
    .A1(net3866),
    .A2(net4922));
 sg13g2_a21oi_1 _18713_ (.A1(_02714_),
    .A2(_02715_),
    .Y(_01116_),
    .B1(_02716_));
 sg13g2_xnor2_1 _18714_ (.Y(_02717_),
    .A(\TRNG.hash[221] ),
    .B(_08245_));
 sg13g2_a21oi_1 _18715_ (.A1(net5557),
    .A2(net5840),
    .Y(_02718_),
    .B1(net4943));
 sg13g2_o21ai_1 _18716_ (.B1(_02718_),
    .Y(_02719_),
    .A1(net5838),
    .A2(_02717_));
 sg13g2_o21ai_1 _18717_ (.B1(_02719_),
    .Y(_02720_),
    .A1(net3887),
    .A2(net4922));
 sg13g2_nor2_1 _18718_ (.A(net5523),
    .B(_02720_),
    .Y(_01117_));
 sg13g2_xnor2_1 _18719_ (.Y(_02721_),
    .A(\TRNG.hash[223] ),
    .B(_08247_));
 sg13g2_a21oi_1 _18720_ (.A1(net5840),
    .A2(\TRNG.hash[255] ),
    .Y(_02722_),
    .B1(net4941));
 sg13g2_o21ai_1 _18721_ (.B1(_02722_),
    .Y(_02723_),
    .A1(net5844),
    .A2(_02721_));
 sg13g2_o21ai_1 _18722_ (.B1(_02723_),
    .Y(_02724_),
    .A1(net3846),
    .A2(net4922));
 sg13g2_nor2_1 _18723_ (.A(net5523),
    .B(_02724_),
    .Y(_01118_));
 sg13g2_and2_1 _18724_ (.A(net5831),
    .B(\TRNG.hash[193] ),
    .X(_02725_));
 sg13g2_a221oi_1 _18725_ (.B2(\TRNG.hash[161] ),
    .C1(_02725_),
    .B1(net5352),
    .A1(net3423),
    .Y(_02726_),
    .A2(net5187));
 sg13g2_a21oi_1 _18726_ (.A1(net5089),
    .A2(net3424),
    .Y(_01119_),
    .B1(net5520));
 sg13g2_xnor2_1 _18727_ (.Y(_02727_),
    .A(net3503),
    .B(_08129_));
 sg13g2_nand2_1 _18728_ (.Y(_02728_),
    .A(net5484),
    .B(_02727_));
 sg13g2_a21oi_1 _18729_ (.A1(net5827),
    .A2(\TRNG.hash[196] ),
    .Y(_02729_),
    .B1(net4939));
 sg13g2_o21ai_1 _18730_ (.B1(net5462),
    .Y(_02730_),
    .A1(\TRNG.hash[164] ),
    .A2(net4919));
 sg13g2_a21oi_1 _18731_ (.A1(_02728_),
    .A2(_02729_),
    .Y(_01120_),
    .B1(_02730_));
 sg13g2_and2_1 _18732_ (.A(\TRNG.hash[165] ),
    .B(_08132_),
    .X(_02731_));
 sg13g2_o21ai_1 _18733_ (.B1(net5484),
    .Y(_02732_),
    .A1(_08133_),
    .A2(_02731_));
 sg13g2_a21oi_1 _18734_ (.A1(net5827),
    .A2(\TRNG.hash[197] ),
    .Y(_02733_),
    .B1(net4939));
 sg13g2_o21ai_1 _18735_ (.B1(net5462),
    .Y(_02734_),
    .A1(net3729),
    .A2(net4919));
 sg13g2_a21oi_1 _18736_ (.A1(_02732_),
    .A2(_02733_),
    .Y(_01121_),
    .B1(_02734_));
 sg13g2_xnor2_1 _18737_ (.Y(_02735_),
    .A(\TRNG.hash[166] ),
    .B(_08133_));
 sg13g2_a21oi_1 _18738_ (.A1(net5827),
    .A2(\TRNG.hash[198] ),
    .Y(_02736_),
    .B1(net4939));
 sg13g2_o21ai_1 _18739_ (.B1(_02736_),
    .Y(_02737_),
    .A1(net5827),
    .A2(_02735_));
 sg13g2_o21ai_1 _18740_ (.B1(_02737_),
    .Y(_02738_),
    .A1(net3848),
    .A2(net4919));
 sg13g2_nor2_1 _18741_ (.A(net5520),
    .B(_02738_),
    .Y(_01122_));
 sg13g2_nand3_1 _18742_ (.B(\TRNG.hash[167] ),
    .C(_08135_),
    .A(\TRNG.hash[168] ),
    .Y(_02739_));
 sg13g2_nor2b_1 _18743_ (.A(_08138_),
    .B_N(_02739_),
    .Y(_02740_));
 sg13g2_a21oi_1 _18744_ (.A1(net5821),
    .A2(\TRNG.hash[200] ),
    .Y(_02741_),
    .B1(net4938));
 sg13g2_o21ai_1 _18745_ (.B1(_02741_),
    .Y(_02742_),
    .A1(net5821),
    .A2(_02740_));
 sg13g2_o21ai_1 _18746_ (.B1(_02742_),
    .Y(_02743_),
    .A1(net3818),
    .A2(net4916));
 sg13g2_nor2_1 _18747_ (.A(net5518),
    .B(_02743_),
    .Y(_01123_));
 sg13g2_xnor2_1 _18748_ (.Y(_02744_),
    .A(\TRNG.hash[169] ),
    .B(_08138_));
 sg13g2_a21oi_1 _18749_ (.A1(\TRNG.hash[201] ),
    .A2(net5820),
    .Y(_02745_),
    .B1(net4938));
 sg13g2_o21ai_1 _18750_ (.B1(_02745_),
    .Y(_02746_),
    .A1(net5816),
    .A2(_02744_));
 sg13g2_o21ai_1 _18751_ (.B1(_02746_),
    .Y(_02747_),
    .A1(net3497),
    .A2(net4916));
 sg13g2_nor2_1 _18752_ (.A(net5518),
    .B(_02747_),
    .Y(_01124_));
 sg13g2_xnor2_1 _18753_ (.Y(_02748_),
    .A(\TRNG.hash[172] ),
    .B(_08144_));
 sg13g2_nand2_1 _18754_ (.Y(_02749_),
    .A(net5483),
    .B(_02748_));
 sg13g2_a21oi_1 _18755_ (.A1(net5817),
    .A2(net3838),
    .Y(_02750_),
    .B1(net4936));
 sg13g2_o21ai_1 _18756_ (.B1(net5461),
    .Y(_02751_),
    .A1(net3849),
    .A2(net4915));
 sg13g2_a21oi_1 _18757_ (.A1(_02749_),
    .A2(_02750_),
    .Y(_01125_),
    .B1(_02751_));
 sg13g2_o21ai_1 _18758_ (.B1(\TRNG.hash[173] ),
    .Y(_02752_),
    .A1(\TRNG.hash[172] ),
    .A2(_08144_));
 sg13g2_nor2b_1 _18759_ (.A(_08148_),
    .B_N(_02752_),
    .Y(_02753_));
 sg13g2_a21oi_1 _18760_ (.A1(\TRNG.hash[205] ),
    .A2(net5817),
    .Y(_02754_),
    .B1(net4936));
 sg13g2_o21ai_1 _18761_ (.B1(_02754_),
    .Y(_02755_),
    .A1(net5817),
    .A2(_02753_));
 sg13g2_o21ai_1 _18762_ (.B1(_02755_),
    .Y(_02756_),
    .A1(net3798),
    .A2(net4915));
 sg13g2_nor2_1 _18763_ (.A(net5518),
    .B(_02756_),
    .Y(_01126_));
 sg13g2_xnor2_1 _18764_ (.Y(_02757_),
    .A(\TRNG.hash[174] ),
    .B(_08148_));
 sg13g2_a21oi_1 _18765_ (.A1(net5822),
    .A2(\TRNG.hash[206] ),
    .Y(_02758_),
    .B1(net4937));
 sg13g2_o21ai_1 _18766_ (.B1(_02758_),
    .Y(_02759_),
    .A1(net5822),
    .A2(_02757_));
 sg13g2_o21ai_1 _18767_ (.B1(_02759_),
    .Y(_02760_),
    .A1(net3857),
    .A2(net4917));
 sg13g2_nor2_1 _18768_ (.A(net5518),
    .B(_02760_),
    .Y(_01127_));
 sg13g2_xnor2_1 _18769_ (.Y(_02761_),
    .A(\TRNG.hash[175] ),
    .B(_08149_));
 sg13g2_a21oi_1 _18770_ (.A1(\TRNG.hash[207] ),
    .A2(net5822),
    .Y(_02762_),
    .B1(net4937));
 sg13g2_o21ai_1 _18771_ (.B1(_02762_),
    .Y(_02763_),
    .A1(net5822),
    .A2(_02761_));
 sg13g2_o21ai_1 _18772_ (.B1(_02763_),
    .Y(_02764_),
    .A1(net3840),
    .A2(net4917));
 sg13g2_nor2_1 _18773_ (.A(net5518),
    .B(_02764_),
    .Y(_01128_));
 sg13g2_nor2b_1 _18774_ (.A(_08151_),
    .B_N(_00223_),
    .Y(_02765_));
 sg13g2_xnor2_1 _18775_ (.Y(_02766_),
    .A(_00223_),
    .B(_08151_));
 sg13g2_nor2_1 _18776_ (.A(net5824),
    .B(_02766_),
    .Y(_02767_));
 sg13g2_a21oi_1 _18777_ (.A1(\TRNG.hash[209] ),
    .A2(net5824),
    .Y(_02768_),
    .B1(_02767_));
 sg13g2_o21ai_1 _18778_ (.B1(net5463),
    .Y(_02769_),
    .A1(net3684),
    .A2(net4918));
 sg13g2_a21oi_1 _18779_ (.A1(net4954),
    .A2(_02768_),
    .Y(_01129_),
    .B1(_02769_));
 sg13g2_xnor2_1 _18780_ (.Y(_02770_),
    .A(\TRNG.hash[178] ),
    .B(_02765_));
 sg13g2_a21oi_1 _18781_ (.A1(\TRNG.hash[210] ),
    .A2(net5824),
    .Y(_02771_),
    .B1(net4938));
 sg13g2_o21ai_1 _18782_ (.B1(_02771_),
    .Y(_02772_),
    .A1(net5824),
    .A2(_02770_));
 sg13g2_o21ai_1 _18783_ (.B1(_02772_),
    .Y(_02773_),
    .A1(net3860),
    .A2(net4918));
 sg13g2_nor2_1 _18784_ (.A(net5519),
    .B(_02773_),
    .Y(_01130_));
 sg13g2_xnor2_1 _18785_ (.Y(_02774_),
    .A(\TRNG.hash[179] ),
    .B(_08155_));
 sg13g2_a21oi_1 _18786_ (.A1(net5824),
    .A2(\TRNG.hash[211] ),
    .Y(_02775_),
    .B1(net4937));
 sg13g2_o21ai_1 _18787_ (.B1(_02775_),
    .Y(_02776_),
    .A1(net5824),
    .A2(_02774_));
 sg13g2_o21ai_1 _18788_ (.B1(_02776_),
    .Y(_02777_),
    .A1(net3777),
    .A2(net4917));
 sg13g2_nor2_1 _18789_ (.A(net5519),
    .B(_02777_),
    .Y(_01131_));
 sg13g2_xnor2_1 _18790_ (.Y(_02778_),
    .A(net3692),
    .B(_08157_));
 sg13g2_a21oi_1 _18791_ (.A1(\TRNG.hash[213] ),
    .A2(net5841),
    .Y(_02779_),
    .B1(net4942));
 sg13g2_o21ai_1 _18792_ (.B1(_02779_),
    .Y(_02780_),
    .A1(net5841),
    .A2(_02778_));
 sg13g2_o21ai_1 _18793_ (.B1(_02780_),
    .Y(_02781_),
    .A1(net3692),
    .A2(net4923));
 sg13g2_nor2_1 _18794_ (.A(net5524),
    .B(net3693),
    .Y(_01132_));
 sg13g2_and2_1 _18795_ (.A(\TRNG.hash[182] ),
    .B(_08161_),
    .X(_02782_));
 sg13g2_o21ai_1 _18796_ (.B1(net5488),
    .Y(_02783_),
    .A1(_08162_),
    .A2(_02782_));
 sg13g2_a21oi_1 _18797_ (.A1(net3784),
    .A2(net5842),
    .Y(_02784_),
    .B1(net4943));
 sg13g2_o21ai_1 _18798_ (.B1(net5467),
    .Y(_02785_),
    .A1(\TRNG.hash[182] ),
    .A2(net4923));
 sg13g2_a21oi_1 _18799_ (.A1(_02783_),
    .A2(_02784_),
    .Y(_01133_),
    .B1(_02785_));
 sg13g2_xnor2_1 _18800_ (.Y(_02786_),
    .A(net3495),
    .B(_08171_));
 sg13g2_nand2_1 _18801_ (.Y(_02787_),
    .A(net5486),
    .B(_02786_));
 sg13g2_a21oi_1 _18802_ (.A1(net5837),
    .A2(\TRNG.hash[218] ),
    .Y(_02788_),
    .B1(net4941));
 sg13g2_o21ai_1 _18803_ (.B1(net5466),
    .Y(_02789_),
    .A1(\TRNG.hash[186] ),
    .A2(net4921));
 sg13g2_a21oi_1 _18804_ (.A1(_02787_),
    .A2(_02788_),
    .Y(_01134_),
    .B1(_02789_));
 sg13g2_o21ai_1 _18805_ (.B1(net3495),
    .Y(_02790_),
    .A1(\TRNG.hash[186] ),
    .A2(_08171_));
 sg13g2_nor2_1 _18806_ (.A(\TRNG.hash[187] ),
    .B(_02790_),
    .Y(_02791_));
 sg13g2_and2_1 _18807_ (.A(\TRNG.hash[187] ),
    .B(_02790_),
    .X(_02792_));
 sg13g2_o21ai_1 _18808_ (.B1(net5486),
    .Y(_02793_),
    .A1(_02791_),
    .A2(_02792_));
 sg13g2_a21oi_1 _18809_ (.A1(net3868),
    .A2(net5837),
    .Y(_02794_),
    .B1(net4941));
 sg13g2_o21ai_1 _18810_ (.B1(net5466),
    .Y(_02795_),
    .A1(\TRNG.hash[187] ),
    .A2(net4921));
 sg13g2_a21oi_1 _18811_ (.A1(_02793_),
    .A2(_02794_),
    .Y(_01135_),
    .B1(_02795_));
 sg13g2_xnor2_1 _18812_ (.Y(_02796_),
    .A(\TRNG.hash[188] ),
    .B(_02791_));
 sg13g2_a21oi_1 _18813_ (.A1(\TRNG.hash[220] ),
    .A2(net5838),
    .Y(_02797_),
    .B1(net4941));
 sg13g2_o21ai_1 _18814_ (.B1(_02797_),
    .Y(_02798_),
    .A1(net5838),
    .A2(_02796_));
 sg13g2_o21ai_1 _18815_ (.B1(_02798_),
    .Y(_02799_),
    .A1(net2591),
    .A2(net4921));
 sg13g2_nor2_1 _18816_ (.A(net5523),
    .B(_02799_),
    .Y(_01136_));
 sg13g2_nand2_1 _18817_ (.Y(_02800_),
    .A(\TRNG.hash[189] ),
    .B(_08176_));
 sg13g2_a21o_1 _18818_ (.A2(_02800_),
    .A1(_08177_),
    .B1(net5839),
    .X(_02801_));
 sg13g2_a21oi_1 _18819_ (.A1(\TRNG.hash[221] ),
    .A2(net5839),
    .Y(_02802_),
    .B1(net4943));
 sg13g2_o21ai_1 _18820_ (.B1(net5466),
    .Y(_02803_),
    .A1(net3830),
    .A2(net4922));
 sg13g2_a21oi_1 _18821_ (.A1(_02801_),
    .A2(_02802_),
    .Y(_01137_),
    .B1(_02803_));
 sg13g2_xor2_1 _18822_ (.B(_07330_),
    .A(\TRNG.hash[128] ),
    .X(_02804_));
 sg13g2_o21ai_1 _18823_ (.B1(net5089),
    .Y(_02805_),
    .A1(net5555),
    .A2(net5845));
 sg13g2_a221oi_1 _18824_ (.B2(net5845),
    .C1(_02805_),
    .B1(_02804_),
    .A1(net5089),
    .Y(_02806_),
    .A2(net5352));
 sg13g2_nor4_1 _18825_ (.A(net5555),
    .B(net5573),
    .C(net5845),
    .D(net5097),
    .Y(_02807_));
 sg13g2_nor3_1 _18826_ (.A(net5527),
    .B(_02806_),
    .C(_02807_),
    .Y(_01138_));
 sg13g2_xnor2_1 _18827_ (.Y(_02808_),
    .A(_07331_),
    .B(_07333_));
 sg13g2_xor2_1 _18828_ (.B(net5555),
    .A(net5554),
    .X(_02809_));
 sg13g2_o21ai_1 _18829_ (.B1(net4955),
    .Y(_02810_),
    .A1(net5845),
    .A2(_02809_));
 sg13g2_a21oi_1 _18830_ (.A1(net5845),
    .A2(_02808_),
    .Y(_02811_),
    .B1(_02810_));
 sg13g2_o21ai_1 _18831_ (.B1(net5469),
    .Y(_02812_),
    .A1(net5554),
    .A2(net4925));
 sg13g2_nor2_1 _18832_ (.A(_02811_),
    .B(_02812_),
    .Y(_01139_));
 sg13g2_xnor2_1 _18833_ (.Y(_02813_),
    .A(_07327_),
    .B(_07334_));
 sg13g2_xor2_1 _18834_ (.B(_07399_),
    .A(net5553),
    .X(_02814_));
 sg13g2_o21ai_1 _18835_ (.B1(net4955),
    .Y(_02815_),
    .A1(net5845),
    .A2(_02814_));
 sg13g2_a21oi_1 _18836_ (.A1(net5846),
    .A2(_02813_),
    .Y(_02816_),
    .B1(_02815_));
 sg13g2_o21ai_1 _18837_ (.B1(net5469),
    .Y(_02817_),
    .A1(net5553),
    .A2(net4925));
 sg13g2_nor2_1 _18838_ (.A(_02816_),
    .B(_02817_),
    .Y(_01140_));
 sg13g2_nand2_1 _18839_ (.Y(_02818_),
    .A(_07335_),
    .B(_07338_));
 sg13g2_nor2_1 _18840_ (.A(net5490),
    .B(_07339_),
    .Y(_02819_));
 sg13g2_xor2_1 _18841_ (.B(_07400_),
    .A(net5552),
    .X(_02820_));
 sg13g2_a221oi_1 _18842_ (.B2(net5490),
    .C1(net4947),
    .B1(_02820_),
    .A1(_02818_),
    .Y(_02821_),
    .A2(_02819_));
 sg13g2_o21ai_1 _18843_ (.B1(net5469),
    .Y(_02822_),
    .A1(net5552),
    .A2(net4925));
 sg13g2_nor2_1 _18844_ (.A(_02821_),
    .B(_02822_),
    .Y(_01141_));
 sg13g2_xnor2_1 _18845_ (.Y(_02823_),
    .A(_07323_),
    .B(_07341_));
 sg13g2_xnor2_1 _18846_ (.Y(_02824_),
    .A(net5551),
    .B(_07401_));
 sg13g2_o21ai_1 _18847_ (.B1(net4955),
    .Y(_02825_),
    .A1(net5845),
    .A2(_02824_));
 sg13g2_a21oi_1 _18848_ (.A1(net5845),
    .A2(_02823_),
    .Y(_02826_),
    .B1(_02825_));
 sg13g2_o21ai_1 _18849_ (.B1(net5469),
    .Y(_02827_),
    .A1(net5551),
    .A2(net4925));
 sg13g2_nor2_1 _18850_ (.A(_02826_),
    .B(_02827_),
    .Y(_01142_));
 sg13g2_xnor2_1 _18851_ (.Y(_02828_),
    .A(_07318_),
    .B(_07342_));
 sg13g2_xnor2_1 _18852_ (.Y(_02829_),
    .A(net5550),
    .B(_07402_));
 sg13g2_o21ai_1 _18853_ (.B1(net4956),
    .Y(_02830_),
    .A1(net5846),
    .A2(_02829_));
 sg13g2_a21oi_1 _18854_ (.A1(net5846),
    .A2(_02828_),
    .Y(_02831_),
    .B1(_02830_));
 sg13g2_o21ai_1 _18855_ (.B1(net5464),
    .Y(_02832_),
    .A1(net5550),
    .A2(net4925));
 sg13g2_nor2_1 _18856_ (.A(_02831_),
    .B(_02832_),
    .Y(_01143_));
 sg13g2_xnor2_1 _18857_ (.Y(_02833_),
    .A(_07343_),
    .B(_07371_));
 sg13g2_xnor2_1 _18858_ (.Y(_02834_),
    .A(net5549),
    .B(_07403_));
 sg13g2_o21ai_1 _18859_ (.B1(net4955),
    .Y(_02835_),
    .A1(net5849),
    .A2(_02834_));
 sg13g2_a21oi_1 _18860_ (.A1(net5846),
    .A2(_02833_),
    .Y(_02836_),
    .B1(_02835_));
 sg13g2_o21ai_1 _18861_ (.B1(net5469),
    .Y(_02837_),
    .A1(net5549),
    .A2(net4925));
 sg13g2_nor2_1 _18862_ (.A(_02836_),
    .B(_02837_),
    .Y(_01144_));
 sg13g2_xor2_1 _18863_ (.B(_07465_),
    .A(_07462_),
    .X(_02838_));
 sg13g2_nand2_1 _18864_ (.Y(_02839_),
    .A(net5846),
    .B(_02838_));
 sg13g2_nand2b_1 _18865_ (.Y(_02840_),
    .B(_07405_),
    .A_N(_00204_));
 sg13g2_xnor2_1 _18866_ (.Y(_02841_),
    .A(net3750),
    .B(_02840_));
 sg13g2_a21oi_1 _18867_ (.A1(net5490),
    .A2(net3751),
    .Y(_02842_),
    .B1(net4947));
 sg13g2_a221oi_1 _18868_ (.B2(_02842_),
    .C1(net5520),
    .B1(_02839_),
    .A1(_04222_),
    .Y(_01145_),
    .A2(net4934));
 sg13g2_a21oi_1 _18869_ (.A1(_07528_),
    .A2(_07529_),
    .Y(_02843_),
    .B1(_07556_));
 sg13g2_nand3b_1 _18870_ (.B(net5834),
    .C(_07558_),
    .Y(_02844_),
    .A_N(_02843_));
 sg13g2_xor2_1 _18871_ (.B(_07586_),
    .A(net3551),
    .X(_02845_));
 sg13g2_a21oi_1 _18872_ (.A1(net5490),
    .A2(_02845_),
    .Y(_02846_),
    .B1(net4947));
 sg13g2_o21ai_1 _18873_ (.B1(net5464),
    .Y(_02847_),
    .A1(net5548),
    .A2(net4926));
 sg13g2_a21oi_1 _18874_ (.A1(_02844_),
    .A2(_02846_),
    .Y(_01146_),
    .B1(_02847_));
 sg13g2_xnor2_1 _18875_ (.Y(_02848_),
    .A(_07638_),
    .B(_07641_));
 sg13g2_xnor2_1 _18876_ (.Y(_02849_),
    .A(net5547),
    .B(_07587_));
 sg13g2_o21ai_1 _18877_ (.B1(net4956),
    .Y(_02850_),
    .A1(net5850),
    .A2(_02849_));
 sg13g2_a21oi_1 _18878_ (.A1(net5850),
    .A2(_02848_),
    .Y(_02851_),
    .B1(_02850_));
 sg13g2_o21ai_1 _18879_ (.B1(net5465),
    .Y(_02852_),
    .A1(net5547),
    .A2(net4926));
 sg13g2_nor2_1 _18880_ (.A(_02851_),
    .B(_02852_),
    .Y(_01147_));
 sg13g2_nand2b_1 _18881_ (.Y(_02853_),
    .B(_07679_),
    .A_N(_07677_));
 sg13g2_xor2_1 _18882_ (.B(_02853_),
    .A(_07761_),
    .X(_02854_));
 sg13g2_xnor2_1 _18883_ (.Y(_02855_),
    .A(net3714),
    .B(_07681_));
 sg13g2_o21ai_1 _18884_ (.B1(net4957),
    .Y(_02856_),
    .A1(net5834),
    .A2(_02855_));
 sg13g2_a21oi_1 _18885_ (.A1(net5834),
    .A2(_02854_),
    .Y(_02857_),
    .B1(_02856_));
 sg13g2_o21ai_1 _18886_ (.B1(net5465),
    .Y(_02858_),
    .A1(net5546),
    .A2(net4926));
 sg13g2_nor2_1 _18887_ (.A(_02857_),
    .B(_02858_),
    .Y(_01148_));
 sg13g2_a22oi_1 _18888_ (.Y(_02859_),
    .B1(_07755_),
    .B2(_07679_),
    .A2(_07753_),
    .A1(_04231_));
 sg13g2_a221oi_1 _18889_ (.B2(_07679_),
    .C1(_07750_),
    .B1(_07755_),
    .A1(_04231_),
    .Y(_02860_),
    .A2(_07753_));
 sg13g2_xnor2_1 _18890_ (.Y(_02861_),
    .A(_07750_),
    .B(_02859_));
 sg13g2_nand2b_1 _18891_ (.Y(_02862_),
    .B(_07681_),
    .A_N(net5546));
 sg13g2_nand2_1 _18892_ (.Y(_02863_),
    .A(net3923),
    .B(_02862_));
 sg13g2_nor2_1 _18893_ (.A(net5545),
    .B(_02863_),
    .Y(_02864_));
 sg13g2_xor2_1 _18894_ (.B(_02863_),
    .A(net5545),
    .X(_02865_));
 sg13g2_o21ai_1 _18895_ (.B1(net4957),
    .Y(_02866_),
    .A1(net5834),
    .A2(_02865_));
 sg13g2_a21oi_1 _18896_ (.A1(net5834),
    .A2(_02861_),
    .Y(_02867_),
    .B1(_02866_));
 sg13g2_o21ai_1 _18897_ (.B1(net5465),
    .Y(_02868_),
    .A1(net5545),
    .A2(net4926));
 sg13g2_nor2_1 _18898_ (.A(_02867_),
    .B(_02868_),
    .Y(_01149_));
 sg13g2_nor2_1 _18899_ (.A(_07749_),
    .B(_02860_),
    .Y(_02869_));
 sg13g2_xnor2_1 _18900_ (.Y(_02870_),
    .A(_07746_),
    .B(_02869_));
 sg13g2_xnor2_1 _18901_ (.Y(_02871_),
    .A(net5544),
    .B(_02864_));
 sg13g2_o21ai_1 _18902_ (.B1(net4957),
    .Y(_02872_),
    .A1(net5834),
    .A2(_02871_));
 sg13g2_a21oi_1 _18903_ (.A1(net5834),
    .A2(_02870_),
    .Y(_02873_),
    .B1(_02872_));
 sg13g2_o21ai_1 _18904_ (.B1(net5465),
    .Y(_02874_),
    .A1(net5544),
    .A2(net4926));
 sg13g2_nor2_1 _18905_ (.A(_02873_),
    .B(_02874_),
    .Y(_01150_));
 sg13g2_xnor2_1 _18906_ (.Y(_02875_),
    .A(_07949_),
    .B(_07950_));
 sg13g2_xnor2_1 _18907_ (.Y(_02876_),
    .A(net3740),
    .B(_07865_));
 sg13g2_o21ai_1 _18908_ (.B1(net4957),
    .Y(_02877_),
    .A1(net5850),
    .A2(_02876_));
 sg13g2_a21oi_1 _18909_ (.A1(net5850),
    .A2(_02875_),
    .Y(_02878_),
    .B1(_02877_));
 sg13g2_o21ai_1 _18910_ (.B1(net5465),
    .Y(_02879_),
    .A1(\TRNG.hash[120] ),
    .A2(net4930));
 sg13g2_nor2_1 _18911_ (.A(_02878_),
    .B(_02879_),
    .Y(_01151_));
 sg13g2_a21oi_1 _18912_ (.A1(_08046_),
    .A2(_08048_),
    .Y(_02880_),
    .B1(net5488));
 sg13g2_o21ai_1 _18913_ (.B1(_02880_),
    .Y(_02881_),
    .A1(_08046_),
    .A2(_08048_));
 sg13g2_xnor2_1 _18914_ (.Y(_02882_),
    .A(_00200_),
    .B(_08017_));
 sg13g2_a21oi_1 _18915_ (.A1(net5492),
    .A2(_02882_),
    .Y(_02883_),
    .B1(net4949));
 sg13g2_o21ai_1 _18916_ (.B1(net5465),
    .Y(_02884_),
    .A1(net3919),
    .A2(net4930));
 sg13g2_a21oi_1 _18917_ (.A1(_02881_),
    .A2(_02883_),
    .Y(_01152_),
    .B1(_02884_));
 sg13g2_xnor2_1 _18918_ (.Y(_02885_),
    .A(_08078_),
    .B(_08099_));
 sg13g2_xnor2_1 _18919_ (.Y(_02886_),
    .A(_04221_),
    .B(_08120_));
 sg13g2_a21oi_1 _18920_ (.A1(net5492),
    .A2(_02886_),
    .Y(_02887_),
    .B1(net4949));
 sg13g2_o21ai_1 _18921_ (.B1(_02887_),
    .Y(_02888_),
    .A1(net5492),
    .A2(_02885_));
 sg13g2_a21oi_1 _18922_ (.A1(_04221_),
    .A2(net4934),
    .Y(_02889_),
    .B1(net5521));
 sg13g2_and2_1 _18923_ (.A(_02888_),
    .B(_02889_),
    .X(_01153_));
 sg13g2_and2_1 _18924_ (.A(net5553),
    .B(net5847),
    .X(_02890_));
 sg13g2_a221oi_1 _18925_ (.B2(\TRNG.hash[66] ),
    .C1(_02890_),
    .B1(net5350),
    .A1(net3445),
    .Y(_02891_),
    .A2(net5187));
 sg13g2_a21oi_1 _18926_ (.A1(net5089),
    .A2(net3446),
    .Y(_01154_),
    .B1(net5527));
 sg13g2_nand2_1 _18927_ (.Y(_02892_),
    .A(\TRNG.hash[67] ),
    .B(\TRNG.hash[66] ));
 sg13g2_a21oi_1 _18928_ (.A1(_07131_),
    .A2(_02892_),
    .Y(_02893_),
    .B1(net5847));
 sg13g2_a21oi_1 _18929_ (.A1(net5552),
    .A2(net5847),
    .Y(_02894_),
    .B1(_02893_));
 sg13g2_o21ai_1 _18930_ (.B1(net5469),
    .Y(_02895_),
    .A1(net3835),
    .A2(net4928));
 sg13g2_a21oi_1 _18931_ (.A1(net4955),
    .A2(_02894_),
    .Y(_01155_),
    .B1(_02895_));
 sg13g2_and4_1 _18932_ (.A(\TRNG.hash[69] ),
    .B(\TRNG.hash[68] ),
    .C(_04378_),
    .D(_07131_),
    .X(_02896_));
 sg13g2_xnor2_1 _18933_ (.Y(_02897_),
    .A(_00180_),
    .B(_02896_));
 sg13g2_a21oi_1 _18934_ (.A1(net5848),
    .A2(net5897),
    .Y(_02898_),
    .B1(net4946));
 sg13g2_o21ai_1 _18935_ (.B1(_02898_),
    .Y(_02899_),
    .A1(net5848),
    .A2(_02897_));
 sg13g2_o21ai_1 _18936_ (.B1(_02899_),
    .Y(_02900_),
    .A1(net3733),
    .A2(net4925));
 sg13g2_nor2_1 _18937_ (.A(net5527),
    .B(net3734),
    .Y(_01156_));
 sg13g2_nor2b_1 _18938_ (.A(_00193_),
    .B_N(_07151_),
    .Y(_02901_));
 sg13g2_xnor2_1 _18939_ (.Y(_02902_),
    .A(_00182_),
    .B(_02901_));
 sg13g2_nor2_1 _18940_ (.A(net5852),
    .B(_02902_),
    .Y(_02903_));
 sg13g2_a21oi_1 _18941_ (.A1(net5852),
    .A2(net3434),
    .Y(_02904_),
    .B1(_02903_));
 sg13g2_o21ai_1 _18942_ (.B1(net5469),
    .Y(_02905_),
    .A1(\TRNG.hash[75] ),
    .A2(net4927));
 sg13g2_a21oi_1 _18943_ (.A1(net4956),
    .A2(net3435),
    .Y(_01157_),
    .B1(_02905_));
 sg13g2_a21oi_1 _18944_ (.A1(\TRNG.hash[76] ),
    .A2(_07156_),
    .Y(_02906_),
    .B1(_00194_));
 sg13g2_nand3_1 _18945_ (.B(_00194_),
    .C(_07156_),
    .A(\TRNG.hash[76] ),
    .Y(_02907_));
 sg13g2_nor2_1 _18946_ (.A(net5851),
    .B(_02906_),
    .Y(_02908_));
 sg13g2_a22oi_1 _18947_ (.Y(_02909_),
    .B1(_02907_),
    .B2(_02908_),
    .A2(net5893),
    .A1(net5851));
 sg13g2_o21ai_1 _18948_ (.B1(net5470),
    .Y(_02910_),
    .A1(net3447),
    .A2(net4927));
 sg13g2_a21oi_1 _18949_ (.A1(net4955),
    .A2(_02909_),
    .Y(_01158_),
    .B1(_02910_));
 sg13g2_or2_1 _18950_ (.X(_02911_),
    .B(_07161_),
    .A(net3415));
 sg13g2_a21o_1 _18951_ (.A2(_02911_),
    .A1(_07163_),
    .B1(net5851),
    .X(_02912_));
 sg13g2_a21oi_1 _18952_ (.A1(net5547),
    .A2(net5851),
    .Y(_02913_),
    .B1(net4947));
 sg13g2_o21ai_1 _18953_ (.B1(net5470),
    .Y(_02914_),
    .A1(net3604),
    .A2(net4926));
 sg13g2_a21oi_1 _18954_ (.A1(_02912_),
    .A2(_02913_),
    .Y(_01159_),
    .B1(_02914_));
 sg13g2_xnor2_1 _18955_ (.Y(_02915_),
    .A(net3553),
    .B(_07167_));
 sg13g2_nor2_1 _18956_ (.A(net5853),
    .B(_02915_),
    .Y(_02916_));
 sg13g2_a21oi_1 _18957_ (.A1(net5852),
    .A2(net5891),
    .Y(_02917_),
    .B1(_02916_));
 sg13g2_o21ai_1 _18958_ (.B1(net5470),
    .Y(_02918_),
    .A1(net3553),
    .A2(net4925));
 sg13g2_a21oi_1 _18959_ (.A1(net4957),
    .A2(_02917_),
    .Y(_01160_),
    .B1(_02918_));
 sg13g2_a21oi_1 _18960_ (.A1(net3455),
    .A2(_07173_),
    .Y(_02919_),
    .B1(net5866));
 sg13g2_o21ai_1 _18961_ (.B1(_02919_),
    .Y(_02920_),
    .A1(net3455),
    .A2(_07173_));
 sg13g2_a21oi_1 _18962_ (.A1(\TRNG.hash[114] ),
    .A2(net5866),
    .Y(_02921_),
    .B1(net4951));
 sg13g2_o21ai_1 _18963_ (.B1(net5470),
    .Y(_02922_),
    .A1(\TRNG.hash[82] ),
    .A2(net4930));
 sg13g2_a21oi_1 _18964_ (.A1(_02920_),
    .A2(_02921_),
    .Y(_01161_),
    .B1(_02922_));
 sg13g2_nand2_1 _18965_ (.Y(_02923_),
    .A(net3667),
    .B(_07190_));
 sg13g2_or2_1 _18966_ (.X(_02924_),
    .B(_07190_),
    .A(net3667));
 sg13g2_a21o_1 _18967_ (.A2(_02924_),
    .A1(_02923_),
    .B1(net5861),
    .X(_02925_));
 sg13g2_a21oi_1 _18968_ (.A1(\TRNG.hash[120] ),
    .A2(net5861),
    .Y(_02926_),
    .B1(net4948));
 sg13g2_o21ai_1 _18969_ (.B1(net5467),
    .Y(_02927_),
    .A1(\TRNG.hash[88] ),
    .A2(net4929));
 sg13g2_a21oi_1 _18970_ (.A1(_02925_),
    .A2(_02926_),
    .Y(_01162_),
    .B1(_02927_));
 sg13g2_xor2_1 _18971_ (.B(_02923_),
    .A(\TRNG.hash[89] ),
    .X(_02928_));
 sg13g2_a21oi_1 _18972_ (.A1(net5861),
    .A2(\TRNG.hash[121] ),
    .Y(_02929_),
    .B1(net4948));
 sg13g2_o21ai_1 _18973_ (.B1(_02929_),
    .Y(_02930_),
    .A1(net5861),
    .A2(_02928_));
 sg13g2_o21ai_1 _18974_ (.B1(_02930_),
    .Y(_02931_),
    .A1(net3815),
    .A2(net4929));
 sg13g2_nor2_1 _18975_ (.A(net5523),
    .B(_02931_),
    .Y(_01163_));
 sg13g2_xor2_1 _18976_ (.B(_07199_),
    .A(_00190_),
    .X(_02932_));
 sg13g2_a21oi_1 _18977_ (.A1(net5862),
    .A2(\TRNG.hash[123] ),
    .Y(_02933_),
    .B1(net4948));
 sg13g2_o21ai_1 _18978_ (.B1(_02933_),
    .Y(_02934_),
    .A1(net5862),
    .A2(_02932_));
 sg13g2_o21ai_1 _18979_ (.B1(_02934_),
    .Y(_02935_),
    .A1(net3781),
    .A2(net4930));
 sg13g2_nor2_1 _18980_ (.A(net5525),
    .B(net3782),
    .Y(_01164_));
 sg13g2_and2_1 _18981_ (.A(\TRNG.hash[92] ),
    .B(_07200_),
    .X(_02936_));
 sg13g2_o21ai_1 _18982_ (.B1(net5492),
    .Y(_02937_),
    .A1(_07201_),
    .A2(_02936_));
 sg13g2_a21oi_1 _18983_ (.A1(\TRNG.hash[124] ),
    .A2(net5862),
    .Y(_02938_),
    .B1(net4948));
 sg13g2_o21ai_1 _18984_ (.B1(net5467),
    .Y(_02939_),
    .A1(net3821),
    .A2(net4929));
 sg13g2_a21oi_1 _18985_ (.A1(_02937_),
    .A2(_02938_),
    .Y(_01165_),
    .B1(_02939_));
 sg13g2_xnor2_1 _18986_ (.Y(_02940_),
    .A(net3388),
    .B(_07207_));
 sg13g2_nand2_1 _18987_ (.Y(_02941_),
    .A(net5492),
    .B(_02940_));
 sg13g2_a21oi_1 _18988_ (.A1(net5863),
    .A2(\TRNG.hash[127] ),
    .Y(_02942_),
    .B1(net4950));
 sg13g2_o21ai_1 _18989_ (.B1(net5473),
    .Y(_02943_),
    .A1(\TRNG.hash[95] ),
    .A2(net4929));
 sg13g2_a21oi_1 _18990_ (.A1(_02941_),
    .A2(_02942_),
    .Y(_01166_),
    .B1(_02943_));
 sg13g2_nor2_1 _18991_ (.A(_04377_),
    .B(net5180),
    .Y(_02944_));
 sg13g2_a221oi_1 _18992_ (.B2(\TRNG.hash[32] ),
    .C1(_02944_),
    .B1(net5350),
    .A1(net5847),
    .Y(_02945_),
    .A2(net3610));
 sg13g2_a21oi_1 _18993_ (.A1(net5090),
    .A2(_02945_),
    .Y(_01167_),
    .B1(net5527));
 sg13g2_xor2_1 _18994_ (.B(\TRNG.hash[32] ),
    .A(\TRNG.hash[33] ),
    .X(_02946_));
 sg13g2_nor2_1 _18995_ (.A(net5847),
    .B(_02946_),
    .Y(_02947_));
 sg13g2_a21oi_1 _18996_ (.A1(net5847),
    .A2(net3565),
    .Y(_02948_),
    .B1(_02947_));
 sg13g2_o21ai_1 _18997_ (.B1(net5469),
    .Y(_02949_),
    .A1(net3745),
    .A2(net4928));
 sg13g2_a21oi_1 _18998_ (.A1(net4955),
    .A2(_02948_),
    .Y(_01168_),
    .B1(_02949_));
 sg13g2_xnor2_1 _18999_ (.Y(_02950_),
    .A(net3537),
    .B(_07066_));
 sg13g2_nand2_1 _19000_ (.Y(_02951_),
    .A(net5491),
    .B(_02950_));
 sg13g2_a21oi_1 _19001_ (.A1(\TRNG.hash[67] ),
    .A2(net5857),
    .Y(_02952_),
    .B1(net4946));
 sg13g2_o21ai_1 _19002_ (.B1(net5471),
    .Y(_02953_),
    .A1(\TRNG.hash[35] ),
    .A2(net4928));
 sg13g2_a21oi_1 _19003_ (.A1(_02951_),
    .A2(_02952_),
    .Y(_01169_),
    .B1(_02953_));
 sg13g2_xor2_1 _19004_ (.B(_07071_),
    .A(net3769),
    .X(_02954_));
 sg13g2_nor2_1 _19005_ (.A(net5857),
    .B(_02954_),
    .Y(_02955_));
 sg13g2_a21oi_1 _19006_ (.A1(net5857),
    .A2(\TRNG.hash[69] ),
    .Y(_02956_),
    .B1(_02955_));
 sg13g2_o21ai_1 _19007_ (.B1(net5471),
    .Y(_02957_),
    .A1(\TRNG.hash[37] ),
    .A2(net4928));
 sg13g2_a21oi_1 _19008_ (.A1(net4955),
    .A2(net3770),
    .Y(_01170_),
    .B1(_02957_));
 sg13g2_a21oi_1 _19009_ (.A1(\TRNG.hash[38] ),
    .A2(_07072_),
    .Y(_02958_),
    .B1(net3522));
 sg13g2_nand3_1 _19010_ (.B(net3522),
    .C(_07072_),
    .A(\TRNG.hash[38] ),
    .Y(_02959_));
 sg13g2_nor2_1 _19011_ (.A(net5848),
    .B(_02958_),
    .Y(_02960_));
 sg13g2_a22oi_1 _19012_ (.Y(_02961_),
    .B1(_02959_),
    .B2(_02960_),
    .A2(net5848),
    .A1(\TRNG.hash[71] ));
 sg13g2_o21ai_1 _19013_ (.B1(net5471),
    .Y(_02962_),
    .A1(net3461),
    .A2(net4928));
 sg13g2_a21oi_1 _19014_ (.A1(net4957),
    .A2(net3523),
    .Y(_01171_),
    .B1(_02962_));
 sg13g2_xnor2_1 _19015_ (.Y(_02963_),
    .A(_00174_),
    .B(_07077_));
 sg13g2_a21oi_1 _19016_ (.A1(net5851),
    .A2(\TRNG.hash[72] ),
    .Y(_02964_),
    .B1(net4945));
 sg13g2_o21ai_1 _19017_ (.B1(_02964_),
    .Y(_02965_),
    .A1(net5848),
    .A2(_02963_));
 sg13g2_o21ai_1 _19018_ (.B1(_02965_),
    .Y(_02966_),
    .A1(net3669),
    .A2(net4927));
 sg13g2_nor2_1 _19019_ (.A(net5527),
    .B(net3670),
    .Y(_01172_));
 sg13g2_xnor2_1 _19020_ (.Y(_02967_),
    .A(_00175_),
    .B(_07085_));
 sg13g2_a21oi_1 _19021_ (.A1(\TRNG.hash[75] ),
    .A2(net5854),
    .Y(_02968_),
    .B1(net4946));
 sg13g2_o21ai_1 _19022_ (.B1(_02968_),
    .Y(_02969_),
    .A1(net5854),
    .A2(_02967_));
 sg13g2_o21ai_1 _19023_ (.B1(net5470),
    .Y(_02970_),
    .A1(net3585),
    .A2(net4928));
 sg13g2_nor2b_1 _19024_ (.A(_02970_),
    .B_N(_02969_),
    .Y(_01173_));
 sg13g2_or2_1 _19025_ (.X(_02971_),
    .B(_07086_),
    .A(_00167_));
 sg13g2_a21o_1 _19026_ (.A2(_02971_),
    .A1(_07088_),
    .B1(net5854),
    .X(_02972_));
 sg13g2_a21oi_1 _19027_ (.A1(net5854),
    .A2(\TRNG.hash[76] ),
    .Y(_02973_),
    .B1(net4945));
 sg13g2_o21ai_1 _19028_ (.B1(net5471),
    .Y(_02974_),
    .A1(net3594),
    .A2(net4927));
 sg13g2_a21oi_1 _19029_ (.A1(_02972_),
    .A2(_02973_),
    .Y(_01174_),
    .B1(_02974_));
 sg13g2_xnor2_1 _19030_ (.Y(_02975_),
    .A(net3614),
    .B(_07092_));
 sg13g2_a21oi_1 _19031_ (.A1(net3604),
    .A2(net5855),
    .Y(_02976_),
    .B1(net4945));
 sg13g2_o21ai_1 _19032_ (.B1(_02976_),
    .Y(_02977_),
    .A1(net5855),
    .A2(_02975_));
 sg13g2_o21ai_1 _19033_ (.B1(_02977_),
    .Y(_02978_),
    .A1(net3614),
    .A2(net4931));
 sg13g2_nor2_1 _19034_ (.A(net5527),
    .B(_02978_),
    .Y(_01175_));
 sg13g2_and2_1 _19035_ (.A(\TRNG.hash[47] ),
    .B(_07093_),
    .X(_02979_));
 sg13g2_o21ai_1 _19036_ (.B1(net5491),
    .Y(_02980_),
    .A1(_07094_),
    .A2(_02979_));
 sg13g2_a21oi_1 _19037_ (.A1(net5852),
    .A2(net3606),
    .Y(_02981_),
    .B1(net4945));
 sg13g2_o21ai_1 _19038_ (.B1(net5470),
    .Y(_02982_),
    .A1(\TRNG.hash[47] ),
    .A2(net4927));
 sg13g2_a21oi_1 _19039_ (.A1(_02980_),
    .A2(_02981_),
    .Y(_01176_),
    .B1(_02982_));
 sg13g2_xnor2_1 _19040_ (.Y(_02983_),
    .A(_00176_),
    .B(_07094_));
 sg13g2_nand2_1 _19041_ (.Y(_02984_),
    .A(net5490),
    .B(_02983_));
 sg13g2_a21oi_1 _19042_ (.A1(\TRNG.hash[80] ),
    .A2(net5853),
    .Y(_02985_),
    .B1(net4945));
 sg13g2_o21ai_1 _19043_ (.B1(net5470),
    .Y(_02986_),
    .A1(net3526),
    .A2(net4927));
 sg13g2_a21oi_1 _19044_ (.A1(_02984_),
    .A2(_02985_),
    .Y(_01177_),
    .B1(_02986_));
 sg13g2_nand3_1 _19045_ (.B(_00176_),
    .C(_07094_),
    .A(net3679),
    .Y(_02987_));
 sg13g2_a21oi_1 _19046_ (.A1(_00176_),
    .A2(_07094_),
    .Y(_02988_),
    .B1(\TRNG.hash[49] ));
 sg13g2_nor2_1 _19047_ (.A(net5852),
    .B(_02988_),
    .Y(_02989_));
 sg13g2_a221oi_1 _19048_ (.B2(_02989_),
    .C1(net4945),
    .B1(_02987_),
    .A1(net5852),
    .Y(_02990_),
    .A2(\TRNG.hash[81] ));
 sg13g2_o21ai_1 _19049_ (.B1(net5470),
    .Y(_02991_),
    .A1(net3679),
    .A2(net4931));
 sg13g2_nor2_1 _19050_ (.A(_02990_),
    .B(_02991_),
    .Y(_01178_));
 sg13g2_nor2_1 _19051_ (.A(_00177_),
    .B(_07106_),
    .Y(_02992_));
 sg13g2_xnor2_1 _19052_ (.Y(_02993_),
    .A(_00172_),
    .B(_02992_));
 sg13g2_a21oi_1 _19053_ (.A1(net5859),
    .A2(net3608),
    .Y(_02994_),
    .B1(net4948));
 sg13g2_o21ai_1 _19054_ (.B1(_02994_),
    .Y(_02995_),
    .A1(net5859),
    .A2(_02993_));
 sg13g2_o21ai_1 _19055_ (.B1(_02995_),
    .Y(_02996_),
    .A1(net3694),
    .A2(net4929));
 sg13g2_nor2_1 _19056_ (.A(net5523),
    .B(net3695),
    .Y(_01179_));
 sg13g2_xnor2_1 _19057_ (.Y(_02997_),
    .A(\TRNG.hash[56] ),
    .B(_07114_));
 sg13g2_nand2_1 _19058_ (.Y(_02998_),
    .A(net5492),
    .B(_02997_));
 sg13g2_a21oi_1 _19059_ (.A1(net3803),
    .A2(net5861),
    .Y(_02999_),
    .B1(net4948));
 sg13g2_o21ai_1 _19060_ (.B1(net5467),
    .Y(_03000_),
    .A1(\TRNG.hash[56] ),
    .A2(net4929));
 sg13g2_a21oi_1 _19061_ (.A1(_02998_),
    .A2(_02999_),
    .Y(_01180_),
    .B1(_03000_));
 sg13g2_o21ai_1 _19062_ (.B1(\TRNG.hash[57] ),
    .Y(_03001_),
    .A1(\TRNG.hash[56] ),
    .A2(_07114_));
 sg13g2_nor2b_1 _19063_ (.A(_07115_),
    .B_N(_03001_),
    .Y(_03002_));
 sg13g2_a21oi_1 _19064_ (.A1(\TRNG.hash[89] ),
    .A2(net5861),
    .Y(_03003_),
    .B1(net4948));
 sg13g2_o21ai_1 _19065_ (.B1(_03003_),
    .Y(_03004_),
    .A1(net5861),
    .A2(_03002_));
 sg13g2_o21ai_1 _19066_ (.B1(_03004_),
    .Y(_03005_),
    .A1(net3850),
    .A2(net4929));
 sg13g2_nor2_1 _19067_ (.A(net5523),
    .B(net3851),
    .Y(_01181_));
 sg13g2_xnor2_1 _19068_ (.Y(_03006_),
    .A(\TRNG.hash[58] ),
    .B(_07115_));
 sg13g2_a21oi_1 _19069_ (.A1(net5863),
    .A2(\TRNG.hash[90] ),
    .Y(_03007_),
    .B1(net4949));
 sg13g2_o21ai_1 _19070_ (.B1(_03007_),
    .Y(_03008_),
    .A1(net5863),
    .A2(_03006_));
 sg13g2_o21ai_1 _19071_ (.B1(_03008_),
    .Y(_03009_),
    .A1(net3763),
    .A2(net4929));
 sg13g2_nor2_1 _19072_ (.A(net5525),
    .B(net3764),
    .Y(_01182_));
 sg13g2_xnor2_1 _19073_ (.Y(_03010_),
    .A(\TRNG.hash[59] ),
    .B(_07116_));
 sg13g2_a21oi_1 _19074_ (.A1(\TRNG.hash[91] ),
    .A2(net5863),
    .Y(_03011_),
    .B1(net4949));
 sg13g2_o21ai_1 _19075_ (.B1(_03011_),
    .Y(_03012_),
    .A1(net5863),
    .A2(_03010_));
 sg13g2_o21ai_1 _19076_ (.B1(_03012_),
    .Y(_03013_),
    .A1(net3775),
    .A2(net4930));
 sg13g2_nor2_1 _19077_ (.A(net5525),
    .B(net3776),
    .Y(_01183_));
 sg13g2_or2_1 _19078_ (.X(_03014_),
    .B(_07117_),
    .A(_00171_));
 sg13g2_a21o_1 _19079_ (.A2(_03014_),
    .A1(_07118_),
    .B1(net5864),
    .X(_03015_));
 sg13g2_a21oi_1 _19080_ (.A1(\TRNG.hash[92] ),
    .A2(net5863),
    .Y(_03016_),
    .B1(net4948));
 sg13g2_o21ai_1 _19081_ (.B1(net5473),
    .Y(_03017_),
    .A1(net3634),
    .A2(net4930));
 sg13g2_a21oi_1 _19082_ (.A1(_03015_),
    .A2(_03016_),
    .Y(_01184_),
    .B1(_03017_));
 sg13g2_nor2_1 _19083_ (.A(\TRNG.hash[0] ),
    .B(net5180),
    .Y(_03018_));
 sg13g2_a221oi_1 _19084_ (.B2(\TRNG.hash[0] ),
    .C1(_03018_),
    .B1(net5350),
    .A1(net5857),
    .Y(_03019_),
    .A2(_04377_));
 sg13g2_a21oi_1 _19085_ (.A1(net5089),
    .A2(_03019_),
    .Y(_01185_),
    .B1(net5527));
 sg13g2_nand2b_1 _19086_ (.Y(_03020_),
    .B(_06989_),
    .A_N(_00157_));
 sg13g2_xnor2_1 _19087_ (.Y(_03021_),
    .A(net3555),
    .B(_03020_));
 sg13g2_nand2_1 _19088_ (.Y(_03022_),
    .A(net5490),
    .B(net3556));
 sg13g2_a21oi_1 _19089_ (.A1(\TRNG.hash[35] ),
    .A2(net5854),
    .Y(_03023_),
    .B1(net4946));
 sg13g2_o21ai_1 _19090_ (.B1(net5472),
    .Y(_03024_),
    .A1(\TRNG.hash[3] ),
    .A2(net4927));
 sg13g2_a21oi_1 _19091_ (.A1(_03022_),
    .A2(_03023_),
    .Y(_01186_),
    .B1(_03024_));
 sg13g2_or2_1 _19092_ (.X(_03025_),
    .B(_06995_),
    .A(_00150_));
 sg13g2_a21o_1 _19093_ (.A2(_03025_),
    .A1(_06996_),
    .B1(net5869),
    .X(_03026_));
 sg13g2_a21oi_1 _19094_ (.A1(net5867),
    .A2(\TRNG.hash[36] ),
    .Y(_03027_),
    .B1(net4951));
 sg13g2_o21ai_1 _19095_ (.B1(net5474),
    .Y(_03028_),
    .A1(net3539),
    .A2(net4931));
 sg13g2_a21oi_1 _19096_ (.A1(_03026_),
    .A2(_03027_),
    .Y(_01187_),
    .B1(_03028_));
 sg13g2_or2_1 _19097_ (.X(_03029_),
    .B(_07008_),
    .A(net3628));
 sg13g2_a21o_1 _19098_ (.A2(_03029_),
    .A1(_07010_),
    .B1(net5856),
    .X(_03030_));
 sg13g2_a21oi_1 _19099_ (.A1(\TRNG.hash[40] ),
    .A2(net5855),
    .Y(_03031_),
    .B1(net4945));
 sg13g2_o21ai_1 _19100_ (.B1(net5472),
    .Y(_03032_),
    .A1(\TRNG.hash[8] ),
    .A2(net4927));
 sg13g2_a21oi_1 _19101_ (.A1(_03030_),
    .A2(_03031_),
    .Y(_01188_),
    .B1(_03032_));
 sg13g2_xnor2_1 _19102_ (.Y(_03033_),
    .A(\TRNG.hash[10] ),
    .B(_07014_));
 sg13g2_a21oi_1 _19103_ (.A1(net5856),
    .A2(\TRNG.hash[42] ),
    .Y(_03034_),
    .B1(net4945));
 sg13g2_o21ai_1 _19104_ (.B1(_03034_),
    .Y(_03035_),
    .A1(net5856),
    .A2(_03033_));
 sg13g2_o21ai_1 _19105_ (.B1(_03035_),
    .Y(_03036_),
    .A1(net3747),
    .A2(net4931));
 sg13g2_nor2_1 _19106_ (.A(net5527),
    .B(net3748),
    .Y(_01189_));
 sg13g2_nand2_1 _19107_ (.Y(_03037_),
    .A(\TRNG.hash[11] ),
    .B(_07015_));
 sg13g2_a21o_1 _19108_ (.A2(_03037_),
    .A1(_07016_),
    .B1(net5869),
    .X(_03038_));
 sg13g2_a21oi_1 _19109_ (.A1(net3585),
    .A2(net5855),
    .Y(_03039_),
    .B1(net4951));
 sg13g2_o21ai_1 _19110_ (.B1(net5472),
    .Y(_03040_),
    .A1(net3768),
    .A2(net4931));
 sg13g2_a21oi_1 _19111_ (.A1(_03038_),
    .A2(_03039_),
    .Y(_01190_),
    .B1(_03040_));
 sg13g2_nand2_1 _19112_ (.Y(_03041_),
    .A(_00158_),
    .B(_07020_));
 sg13g2_or2_1 _19113_ (.X(_03042_),
    .B(_07020_),
    .A(_00158_));
 sg13g2_a21o_1 _19114_ (.A2(_03042_),
    .A1(_03041_),
    .B1(net5868),
    .X(_03043_));
 sg13g2_a21oi_1 _19115_ (.A1(net3614),
    .A2(net5867),
    .Y(_03044_),
    .B1(net4951));
 sg13g2_o21ai_1 _19116_ (.B1(net5474),
    .Y(_03045_),
    .A1(\TRNG.hash[14] ),
    .A2(net4931));
 sg13g2_a21oi_1 _19117_ (.A1(_03043_),
    .A2(_03044_),
    .Y(_01191_),
    .B1(_03045_));
 sg13g2_xor2_1 _19118_ (.B(_03041_),
    .A(\TRNG.hash[15] ),
    .X(_03046_));
 sg13g2_a21oi_1 _19119_ (.A1(\TRNG.hash[47] ),
    .A2(net5867),
    .Y(_03047_),
    .B1(net4951));
 sg13g2_o21ai_1 _19120_ (.B1(_03047_),
    .Y(_03048_),
    .A1(net5867),
    .A2(_03046_));
 sg13g2_o21ai_1 _19121_ (.B1(_03048_),
    .Y(_03049_),
    .A1(net3858),
    .A2(net4931));
 sg13g2_nor2_1 _19122_ (.A(net5525),
    .B(net3859),
    .Y(_01192_));
 sg13g2_xnor2_1 _19123_ (.Y(_03050_),
    .A(net3677),
    .B(_07041_));
 sg13g2_a21oi_1 _19124_ (.A1(net5868),
    .A2(net3571),
    .Y(_03051_),
    .B1(net4950));
 sg13g2_o21ai_1 _19125_ (.B1(_03051_),
    .Y(_03052_),
    .A1(net5868),
    .A2(_03050_));
 sg13g2_o21ai_1 _19126_ (.B1(_03052_),
    .Y(_03053_),
    .A1(\TRNG.hash[21] ),
    .A2(net4932));
 sg13g2_nor2_1 _19127_ (.A(net5526),
    .B(net3678),
    .Y(_01193_));
 sg13g2_o21ai_1 _19128_ (.B1(net3677),
    .Y(_03054_),
    .A1(\TRNG.hash[21] ),
    .A2(_07042_));
 sg13g2_nor2_1 _19129_ (.A(\TRNG.hash[22] ),
    .B(_03054_),
    .Y(_03055_));
 sg13g2_and2_1 _19130_ (.A(\TRNG.hash[22] ),
    .B(_03054_),
    .X(_03056_));
 sg13g2_o21ai_1 _19131_ (.B1(net5493),
    .Y(_03057_),
    .A1(_03055_),
    .A2(_03056_));
 sg13g2_a21oi_1 _19132_ (.A1(net5860),
    .A2(net3558),
    .Y(_03058_),
    .B1(net4950));
 sg13g2_o21ai_1 _19133_ (.B1(net5473),
    .Y(_03059_),
    .A1(net3728),
    .A2(net4932));
 sg13g2_a21oi_1 _19134_ (.A1(_03057_),
    .A2(_03058_),
    .Y(_01194_),
    .B1(_03059_));
 sg13g2_xnor2_1 _19135_ (.Y(_03060_),
    .A(\TRNG.hash[23] ),
    .B(_03055_));
 sg13g2_a21oi_1 _19136_ (.A1(net3694),
    .A2(net5868),
    .Y(_03061_),
    .B1(net4950));
 sg13g2_o21ai_1 _19137_ (.B1(_03061_),
    .Y(_03062_),
    .A1(net5868),
    .A2(_03060_));
 sg13g2_o21ai_1 _19138_ (.B1(_03062_),
    .Y(_03063_),
    .A1(net3813),
    .A2(net4932));
 sg13g2_nor2_1 _19139_ (.A(net5525),
    .B(_03063_),
    .Y(_01195_));
 sg13g2_xnor2_1 _19140_ (.Y(_03064_),
    .A(\TRNG.hash[24] ),
    .B(_07046_));
 sg13g2_a21oi_1 _19141_ (.A1(\TRNG.hash[56] ),
    .A2(net5868),
    .Y(_03065_),
    .B1(net4950));
 sg13g2_o21ai_1 _19142_ (.B1(_03065_),
    .Y(_03066_),
    .A1(net5869),
    .A2(_03064_));
 sg13g2_o21ai_1 _19143_ (.B1(_03066_),
    .Y(_03067_),
    .A1(net3829),
    .A2(net4932));
 sg13g2_nor2_1 _19144_ (.A(net5525),
    .B(_03067_),
    .Y(_01196_));
 sg13g2_xnor2_1 _19145_ (.Y(_03068_),
    .A(\TRNG.hash[25] ),
    .B(_07047_));
 sg13g2_a21oi_1 _19146_ (.A1(\TRNG.hash[57] ),
    .A2(net5870),
    .Y(_03069_),
    .B1(net4950));
 sg13g2_o21ai_1 _19147_ (.B1(_03069_),
    .Y(_03070_),
    .A1(net5871),
    .A2(_03068_));
 sg13g2_o21ai_1 _19148_ (.B1(_03070_),
    .Y(_03071_),
    .A1(net3834),
    .A2(net4931));
 sg13g2_nor2_1 _19149_ (.A(net5525),
    .B(_03071_),
    .Y(_01197_));
 sg13g2_xnor2_1 _19150_ (.Y(_03072_),
    .A(\TRNG.hash[27] ),
    .B(_07049_));
 sg13g2_nand2_1 _19151_ (.Y(_03073_),
    .A(net5492),
    .B(_03072_));
 sg13g2_a21oi_1 _19152_ (.A1(net3775),
    .A2(net5870),
    .Y(_03074_),
    .B1(net4951));
 sg13g2_o21ai_1 _19153_ (.B1(net5473),
    .Y(_03075_),
    .A1(net3820),
    .A2(net4932));
 sg13g2_a21oi_1 _19154_ (.A1(_03073_),
    .A2(_03074_),
    .Y(_01198_),
    .B1(_03075_));
 sg13g2_o21ai_1 _19155_ (.B1(\TRNG.hash[28] ),
    .Y(_03076_),
    .A1(\TRNG.hash[27] ),
    .A2(_07049_));
 sg13g2_nor2b_1 _19156_ (.A(_07053_),
    .B_N(_03076_),
    .Y(_03077_));
 sg13g2_a21oi_1 _19157_ (.A1(net3634),
    .A2(net5870),
    .Y(_03078_),
    .B1(net4950));
 sg13g2_o21ai_1 _19158_ (.B1(_03078_),
    .Y(_03079_),
    .A1(net5870),
    .A2(_03077_));
 sg13g2_o21ai_1 _19159_ (.B1(_03079_),
    .Y(_03080_),
    .A1(net3735),
    .A2(net4932));
 sg13g2_nor2_1 _19160_ (.A(net5525),
    .B(_03080_),
    .Y(_01199_));
 sg13g2_xnor2_1 _19161_ (.Y(_03081_),
    .A(\TRNG.hash[30] ),
    .B(_07054_));
 sg13g2_a21oi_1 _19162_ (.A1(net5863),
    .A2(net3722),
    .Y(_03082_),
    .B1(net4950));
 sg13g2_o21ai_1 _19163_ (.B1(_03082_),
    .Y(_03083_),
    .A1(net5864),
    .A2(_03081_));
 sg13g2_o21ai_1 _19164_ (.B1(_03083_),
    .Y(_03084_),
    .A1(net3862),
    .A2(net4932));
 sg13g2_nor2_1 _19165_ (.A(net5526),
    .B(_03084_),
    .Y(_01200_));
 sg13g2_nor2_2 _19166_ (.A(net5360),
    .B(_06913_),
    .Y(_03085_));
 sg13g2_mux2_1 _19167_ (.A0(net2837),
    .A1(net5689),
    .S(net4980),
    .X(_01201_));
 sg13g2_mux2_1 _19168_ (.A0(net2774),
    .A1(net5688),
    .S(net4980),
    .X(_01202_));
 sg13g2_mux2_1 _19169_ (.A0(net2790),
    .A1(net5684),
    .S(net4981),
    .X(_01203_));
 sg13g2_nor2_1 _19170_ (.A(net2617),
    .B(net4982),
    .Y(_03086_));
 sg13g2_a21oi_1 _19171_ (.A1(net5496),
    .A2(net4982),
    .Y(_01204_),
    .B1(_03086_));
 sg13g2_mux2_1 _19172_ (.A0(net2664),
    .A1(net5682),
    .S(net4981),
    .X(_01205_));
 sg13g2_mux2_1 _19173_ (.A0(net2715),
    .A1(net5681),
    .S(net4981),
    .X(_01206_));
 sg13g2_mux2_1 _19174_ (.A0(net2798),
    .A1(net5676),
    .S(net4981),
    .X(_01207_));
 sg13g2_mux2_1 _19175_ (.A0(net2742),
    .A1(net5675),
    .S(net4983),
    .X(_01208_));
 sg13g2_mux2_1 _19176_ (.A0(net3122),
    .A1(net5671),
    .S(net4981),
    .X(_01209_));
 sg13g2_mux2_1 _19177_ (.A0(net3055),
    .A1(net5669),
    .S(net4983),
    .X(_01210_));
 sg13g2_mux2_1 _19178_ (.A0(net2897),
    .A1(net5667),
    .S(net4983),
    .X(_01211_));
 sg13g2_mux2_1 _19179_ (.A0(net2675),
    .A1(net5666),
    .S(net4980),
    .X(_01212_));
 sg13g2_mux2_1 _19180_ (.A0(net2931),
    .A1(net5663),
    .S(net4980),
    .X(_01213_));
 sg13g2_mux2_1 _19181_ (.A0(net2752),
    .A1(net5661),
    .S(net4980),
    .X(_01214_));
 sg13g2_mux2_1 _19182_ (.A0(net2922),
    .A1(net5658),
    .S(net4983),
    .X(_01215_));
 sg13g2_mux2_1 _19183_ (.A0(net2952),
    .A1(net5656),
    .S(net4980),
    .X(_01216_));
 sg13g2_mux2_1 _19184_ (.A0(net2923),
    .A1(net5653),
    .S(net4983),
    .X(_01217_));
 sg13g2_mux2_1 _19185_ (.A0(net2920),
    .A1(net5652),
    .S(net4982),
    .X(_01218_));
 sg13g2_mux2_1 _19186_ (.A0(net2849),
    .A1(net5649),
    .S(net4980),
    .X(_01219_));
 sg13g2_mux2_1 _19187_ (.A0(net2892),
    .A1(net5647),
    .S(net4981),
    .X(_01220_));
 sg13g2_mux2_1 _19188_ (.A0(net2911),
    .A1(net5644),
    .S(net4982),
    .X(_01221_));
 sg13g2_mux2_1 _19189_ (.A0(net2893),
    .A1(net5640),
    .S(net4982),
    .X(_01222_));
 sg13g2_mux2_1 _19190_ (.A0(net2872),
    .A1(net5637),
    .S(net4982),
    .X(_01223_));
 sg13g2_mux2_1 _19191_ (.A0(net3001),
    .A1(net5636),
    .S(net4984),
    .X(_01224_));
 sg13g2_mux2_1 _19192_ (.A0(net2667),
    .A1(net5634),
    .S(net4982),
    .X(_01225_));
 sg13g2_mux2_1 _19193_ (.A0(net2716),
    .A1(\TRNG.sha256.expand.data1_to_ram[25] ),
    .S(net4982),
    .X(_01226_));
 sg13g2_mux2_1 _19194_ (.A0(net3013),
    .A1(net5630),
    .S(net4984),
    .X(_01227_));
 sg13g2_mux2_1 _19195_ (.A0(net3255),
    .A1(net5628),
    .S(net4980),
    .X(_01228_));
 sg13g2_mux2_1 _19196_ (.A0(net2782),
    .A1(net5624),
    .S(net4983),
    .X(_01229_));
 sg13g2_mux2_1 _19197_ (.A0(net2743),
    .A1(net5621),
    .S(net4983),
    .X(_01230_));
 sg13g2_mux2_1 _19198_ (.A0(net2918),
    .A1(net5618),
    .S(net4981),
    .X(_01231_));
 sg13g2_mux2_1 _19199_ (.A0(net2924),
    .A1(net5617),
    .S(net4983),
    .X(_01232_));
 sg13g2_nor2_1 _19200_ (.A(net3149),
    .B(\TRNG.Repetition_Count_Test.failure ),
    .Y(_03087_));
 sg13g2_nor2_1 _19201_ (.A(_06328_),
    .B(net3150),
    .Y(_01233_));
 sg13g2_nor2_2 _19202_ (.A(_04838_),
    .B(_04888_),
    .Y(_03088_));
 sg13g2_nand2_1 _19203_ (.Y(_03089_),
    .A(_04838_),
    .B(_04883_));
 sg13g2_mux2_1 _19204_ (.A0(net2999),
    .A1(_04889_),
    .S(_03089_),
    .X(_01234_));
 sg13g2_o21ai_1 _19205_ (.B1(net5524),
    .Y(_03090_),
    .A1(net3870),
    .A2(_04837_));
 sg13g2_o21ai_1 _19206_ (.B1(net4606),
    .Y(_01235_),
    .A1(_04853_),
    .A2(_03090_));
 sg13g2_nand2_1 _19207_ (.Y(_03091_),
    .A(net5899),
    .B(_03088_));
 sg13g2_and2_1 _19208_ (.A(\TRNG.chunk_index[0] ),
    .B(\TRNG.chunk_index[1] ),
    .X(_03092_));
 sg13g2_nor2_2 _19209_ (.A(_04343_),
    .B(\TRNG.chunk_index[1] ),
    .Y(_03093_));
 sg13g2_nor2_2 _19210_ (.A(\TRNG.chunk_index[0] ),
    .B(\TRNG.chunk_index[1] ),
    .Y(_03094_));
 sg13g2_a22oi_1 _19211_ (.Y(_03095_),
    .B1(net5320),
    .B2(\TRNG.hash[128] ),
    .A2(net5107),
    .A1(\TRNG.hash[136] ));
 sg13g2_nor2b_1 _19212_ (.A(\TRNG.chunk_index[0] ),
    .B_N(\TRNG.chunk_index[1] ),
    .Y(_03096_));
 sg13g2_a221oi_1 _19213_ (.B2(\TRNG.hash[144] ),
    .C1(net5512),
    .B1(net5309),
    .A1(\TRNG.hash[152] ),
    .Y(_03097_),
    .A2(net5333));
 sg13g2_a22oi_1 _19214_ (.Y(_03098_),
    .B1(net5316),
    .B2(\TRNG.hash[160] ),
    .A2(net5107),
    .A1(\TRNG.hash[168] ));
 sg13g2_a221oi_1 _19215_ (.B2(\TRNG.hash[176] ),
    .C1(net5459),
    .B1(net5307),
    .A1(\TRNG.hash[184] ),
    .Y(_03099_),
    .A2(net5332));
 sg13g2_a221oi_1 _19216_ (.B2(_03099_),
    .C1(net5509),
    .B1(_03098_),
    .A1(_03095_),
    .Y(_03100_),
    .A2(_03097_));
 sg13g2_nand2_1 _19217_ (.Y(_03101_),
    .A(net5510),
    .B(net5514));
 sg13g2_a22oi_1 _19218_ (.Y(_03102_),
    .B1(net5305),
    .B2(\TRNG.hash[240] ),
    .A2(net5317),
    .A1(net5570));
 sg13g2_a22oi_1 _19219_ (.Y(_03103_),
    .B1(net5103),
    .B2(net5886),
    .A2(net5328),
    .A1(net5879));
 sg13g2_a21oi_1 _19220_ (.A1(_03102_),
    .A2(_03103_),
    .Y(_03104_),
    .B1(net5303));
 sg13g2_nand2_1 _19221_ (.Y(_03105_),
    .A(net5510),
    .B(net5460));
 sg13g2_a22oi_1 _19222_ (.Y(_03106_),
    .B1(net5305),
    .B2(\TRNG.hash[208] ),
    .A2(net5103),
    .A1(\TRNG.hash[200] ));
 sg13g2_a22oi_1 _19223_ (.Y(_03107_),
    .B1(net5318),
    .B2(\TRNG.hash[192] ),
    .A2(net5330),
    .A1(\TRNG.hash[216] ));
 sg13g2_a21oi_1 _19224_ (.A1(_03106_),
    .A2(_03107_),
    .Y(_03108_),
    .B1(net5101));
 sg13g2_nor4_2 _19225_ (.A(_04341_),
    .B(_03100_),
    .C(_03104_),
    .Y(_03109_),
    .D(_03108_));
 sg13g2_a22oi_1 _19226_ (.Y(_03110_),
    .B1(net5324),
    .B2(\TRNG.hash[0] ),
    .A2(net5339),
    .A1(\TRNG.hash[24] ));
 sg13g2_a221oi_1 _19227_ (.B2(\TRNG.hash[16] ),
    .C1(net5513),
    .B1(net5314),
    .A1(\TRNG.hash[8] ),
    .Y(_03111_),
    .A2(net5111));
 sg13g2_a21oi_1 _19228_ (.A1(\TRNG.hash[56] ),
    .A2(net5337),
    .Y(_03112_),
    .B1(_04342_));
 sg13g2_nand2_1 _19229_ (.Y(_03113_),
    .A(\TRNG.hash[32] ),
    .B(net5327));
 sg13g2_a22oi_1 _19230_ (.Y(_03114_),
    .B1(net5314),
    .B2(\TRNG.hash[48] ),
    .A2(net5111),
    .A1(\TRNG.hash[40] ));
 sg13g2_and2_1 _19231_ (.A(_03112_),
    .B(_03114_),
    .X(_03115_));
 sg13g2_a221oi_1 _19232_ (.B2(_03115_),
    .C1(\TRNG.chunk_index[3] ),
    .B1(_03113_),
    .A1(_03110_),
    .Y(_03116_),
    .A2(_03111_));
 sg13g2_a22oi_1 _19233_ (.Y(_03117_),
    .B1(net5327),
    .B2(\TRNG.hash[64] ),
    .A2(net5334),
    .A1(\TRNG.hash[88] ));
 sg13g2_a22oi_1 _19234_ (.Y(_03118_),
    .B1(net5310),
    .B2(\TRNG.hash[80] ),
    .A2(net5114),
    .A1(\TRNG.hash[72] ));
 sg13g2_a21oi_1 _19235_ (.A1(_03117_),
    .A2(_03118_),
    .Y(_03119_),
    .B1(net5102));
 sg13g2_a22oi_1 _19236_ (.Y(_03120_),
    .B1(net5310),
    .B2(net5891),
    .A2(net5334),
    .A1(\TRNG.hash[120] ));
 sg13g2_a22oi_1 _19237_ (.Y(_03121_),
    .B1(net5322),
    .B2(\TRNG.hash[96] ),
    .A2(net5109),
    .A1(net5896));
 sg13g2_a21oi_1 _19238_ (.A1(_03120_),
    .A2(_03121_),
    .Y(_03122_),
    .B1(net5304));
 sg13g2_nor4_2 _19239_ (.A(\TRNG.chunk_index[4] ),
    .B(_03116_),
    .C(_03119_),
    .Y(_03123_),
    .D(_03122_));
 sg13g2_nor3_2 _19240_ (.A(net4556),
    .B(_03109_),
    .C(_03123_),
    .Y(_03124_));
 sg13g2_a21o_1 _19241_ (.A2(net4556),
    .A1(net3108),
    .B1(_03124_),
    .X(_01236_));
 sg13g2_a22oi_1 _19242_ (.Y(_03125_),
    .B1(net5316),
    .B2(\TRNG.hash[161] ),
    .A2(net5106),
    .A1(\TRNG.hash[169] ));
 sg13g2_a221oi_1 _19243_ (.B2(\TRNG.hash[177] ),
    .C1(net5459),
    .B1(net5315),
    .A1(\TRNG.hash[185] ),
    .Y(_03126_),
    .A2(net5332));
 sg13g2_a22oi_1 _19244_ (.Y(_03127_),
    .B1(net5316),
    .B2(\TRNG.hash[129] ),
    .A2(net5107),
    .A1(\TRNG.hash[137] ));
 sg13g2_a221oi_1 _19245_ (.B2(\TRNG.hash[145] ),
    .C1(net5512),
    .B1(net5309),
    .A1(\TRNG.hash[153] ),
    .Y(_03128_),
    .A2(net5332));
 sg13g2_a221oi_1 _19246_ (.B2(_03128_),
    .C1(net5509),
    .B1(_03127_),
    .A1(_03125_),
    .Y(_03129_),
    .A2(_03126_));
 sg13g2_a22oi_1 _19247_ (.Y(_03130_),
    .B1(net5318),
    .B2(net5569),
    .A2(net5103),
    .A1(net5565));
 sg13g2_a22oi_1 _19248_ (.Y(_03131_),
    .B1(net5305),
    .B2(\TRNG.hash[241] ),
    .A2(net5328),
    .A1(net5559));
 sg13g2_a21oi_1 _19249_ (.A1(_03130_),
    .A2(_03131_),
    .Y(_03132_),
    .B1(net5303));
 sg13g2_a22oi_1 _19250_ (.Y(_03133_),
    .B1(net5318),
    .B2(\TRNG.hash[193] ),
    .A2(net5330),
    .A1(\TRNG.hash[217] ));
 sg13g2_a22oi_1 _19251_ (.Y(_03134_),
    .B1(net5305),
    .B2(\TRNG.hash[209] ),
    .A2(net5104),
    .A1(\TRNG.hash[201] ));
 sg13g2_a21oi_1 _19252_ (.A1(_03133_),
    .A2(_03134_),
    .Y(_03135_),
    .B1(net5101));
 sg13g2_nor4_2 _19253_ (.A(_04341_),
    .B(_03129_),
    .C(_03132_),
    .Y(_03136_),
    .D(_03135_));
 sg13g2_a22oi_1 _19254_ (.Y(_03137_),
    .B1(net5324),
    .B2(\TRNG.hash[1] ),
    .A2(net5111),
    .A1(\TRNG.hash[9] ));
 sg13g2_a221oi_1 _19255_ (.B2(\TRNG.hash[17] ),
    .C1(net5513),
    .B1(net5314),
    .A1(\TRNG.hash[25] ),
    .Y(_03138_),
    .A2(net5339));
 sg13g2_a22oi_1 _19256_ (.Y(_03139_),
    .B1(net5327),
    .B2(\TRNG.hash[33] ),
    .A2(net5114),
    .A1(\TRNG.hash[41] ));
 sg13g2_a221oi_1 _19257_ (.B2(\TRNG.hash[49] ),
    .C1(_04342_),
    .B1(net5314),
    .A1(\TRNG.hash[57] ),
    .Y(_03140_),
    .A2(net5339));
 sg13g2_a221oi_1 _19258_ (.B2(_03140_),
    .C1(\TRNG.chunk_index[3] ),
    .B1(_03139_),
    .A1(_03137_),
    .Y(_03141_),
    .A2(_03138_));
 sg13g2_a22oi_1 _19259_ (.Y(_03142_),
    .B1(net5109),
    .B2(\TRNG.hash[105] ),
    .A2(net5334),
    .A1(\TRNG.hash[121] ));
 sg13g2_a22oi_1 _19260_ (.Y(_03143_),
    .B1(net5310),
    .B2(net5546),
    .A2(net5322),
    .A1(\TRNG.hash[97] ));
 sg13g2_a21oi_1 _19261_ (.A1(_03142_),
    .A2(_03143_),
    .Y(_03144_),
    .B1(net5304));
 sg13g2_a22oi_1 _19262_ (.Y(_03145_),
    .B1(net5310),
    .B2(\TRNG.hash[81] ),
    .A2(net5327),
    .A1(\TRNG.hash[65] ));
 sg13g2_a22oi_1 _19263_ (.Y(_03146_),
    .B1(net5114),
    .B2(\TRNG.hash[73] ),
    .A2(net5334),
    .A1(\TRNG.hash[89] ));
 sg13g2_a21oi_1 _19264_ (.A1(_03145_),
    .A2(_03146_),
    .Y(_03147_),
    .B1(net5102));
 sg13g2_nor4_2 _19265_ (.A(\TRNG.chunk_index[4] ),
    .B(_03141_),
    .C(_03144_),
    .Y(_03148_),
    .D(_03147_));
 sg13g2_nor3_2 _19266_ (.A(net4556),
    .B(_03136_),
    .C(_03148_),
    .Y(_03149_));
 sg13g2_a21o_1 _19267_ (.A2(net4556),
    .A1(net2862),
    .B1(_03149_),
    .X(_01237_));
 sg13g2_a22oi_1 _19268_ (.Y(_03150_),
    .B1(net5327),
    .B2(\TRNG.hash[34] ),
    .A2(net5111),
    .A1(\TRNG.hash[42] ));
 sg13g2_a221oi_1 _19269_ (.B2(\TRNG.hash[50] ),
    .C1(net5460),
    .B1(net5312),
    .A1(\TRNG.hash[58] ),
    .Y(_03151_),
    .A2(net5336));
 sg13g2_a22oi_1 _19270_ (.Y(_03152_),
    .B1(net5324),
    .B2(\TRNG.hash[2] ),
    .A2(net5111),
    .A1(\TRNG.hash[10] ));
 sg13g2_a221oi_1 _19271_ (.B2(\TRNG.hash[18] ),
    .C1(net5513),
    .B1(net5312),
    .A1(\TRNG.hash[26] ),
    .Y(_03153_),
    .A2(net5336));
 sg13g2_a221oi_1 _19272_ (.B2(_03153_),
    .C1(net5511),
    .B1(_03152_),
    .A1(_03150_),
    .Y(_03154_),
    .A2(_03151_));
 sg13g2_a22oi_1 _19273_ (.Y(_03155_),
    .B1(net5310),
    .B2(\TRNG.hash[82] ),
    .A2(net5109),
    .A1(\TRNG.hash[74] ));
 sg13g2_a22oi_1 _19274_ (.Y(_03156_),
    .B1(net5322),
    .B2(\TRNG.hash[66] ),
    .A2(net5339),
    .A1(\TRNG.hash[90] ));
 sg13g2_a21oi_1 _19275_ (.A1(_03155_),
    .A2(_03156_),
    .Y(_03157_),
    .B1(net5102));
 sg13g2_a22oi_1 _19276_ (.Y(_03158_),
    .B1(net5322),
    .B2(\TRNG.hash[98] ),
    .A2(net5109),
    .A1(net5895));
 sg13g2_a22oi_1 _19277_ (.Y(_03159_),
    .B1(net5310),
    .B2(net5545),
    .A2(net5334),
    .A1(\TRNG.hash[122] ));
 sg13g2_a21oi_1 _19278_ (.A1(_03158_),
    .A2(_03159_),
    .Y(_03160_),
    .B1(net5304));
 sg13g2_nor4_2 _19279_ (.A(net5508),
    .B(_03154_),
    .C(_03157_),
    .Y(_03161_),
    .D(_03160_));
 sg13g2_a22oi_1 _19280_ (.Y(_03162_),
    .B1(net5307),
    .B2(\TRNG.hash[178] ),
    .A2(net5105),
    .A1(\TRNG.hash[170] ));
 sg13g2_a221oi_1 _19281_ (.B2(\TRNG.hash[162] ),
    .C1(net5459),
    .B1(net5319),
    .A1(\TRNG.hash[186] ),
    .Y(_03163_),
    .A2(net5332));
 sg13g2_a22oi_1 _19282_ (.Y(_03164_),
    .B1(net5316),
    .B2(\TRNG.hash[130] ),
    .A2(net5107),
    .A1(\TRNG.hash[138] ));
 sg13g2_a221oi_1 _19283_ (.B2(\TRNG.hash[146] ),
    .C1(net5512),
    .B1(net5309),
    .A1(\TRNG.hash[154] ),
    .Y(_03165_),
    .A2(net5332));
 sg13g2_a221oi_1 _19284_ (.B2(_03165_),
    .C1(net5509),
    .B1(_03164_),
    .A1(_03162_),
    .Y(_03166_),
    .A2(_03163_));
 sg13g2_a22oi_1 _19285_ (.Y(_03167_),
    .B1(net5316),
    .B2(\TRNG.hash[194] ),
    .A2(net5106),
    .A1(\TRNG.hash[202] ));
 sg13g2_a22oi_1 _19286_ (.Y(_03168_),
    .B1(net5305),
    .B2(\TRNG.hash[210] ),
    .A2(net5328),
    .A1(\TRNG.hash[218] ));
 sg13g2_a21oi_1 _19287_ (.A1(_03167_),
    .A2(_03168_),
    .Y(_03169_),
    .B1(net5101));
 sg13g2_a22oi_1 _19288_ (.Y(_03170_),
    .B1(net5305),
    .B2(net5883),
    .A2(net5328),
    .A1(net5878));
 sg13g2_a22oi_1 _19289_ (.Y(_03171_),
    .B1(net5317),
    .B2(\TRNG.hash[226] ),
    .A2(net5103),
    .A1(net5564));
 sg13g2_a21oi_1 _19290_ (.A1(_03170_),
    .A2(_03171_),
    .Y(_03172_),
    .B1(net5303));
 sg13g2_nor4_2 _19291_ (.A(_04341_),
    .B(_03166_),
    .C(_03169_),
    .Y(_03173_),
    .D(_03172_));
 sg13g2_nor3_2 _19292_ (.A(net4556),
    .B(_03161_),
    .C(_03173_),
    .Y(_03174_));
 sg13g2_a21o_1 _19293_ (.A2(net4555),
    .A1(net2763),
    .B1(_03174_),
    .X(_01238_));
 sg13g2_a22oi_1 _19294_ (.Y(_03175_),
    .B1(net5327),
    .B2(\TRNG.hash[35] ),
    .A2(net5114),
    .A1(\TRNG.hash[43] ));
 sg13g2_a221oi_1 _19295_ (.B2(\TRNG.hash[51] ),
    .C1(net5460),
    .B1(net5312),
    .A1(\TRNG.hash[59] ),
    .Y(_03176_),
    .A2(net5336));
 sg13g2_a22oi_1 _19296_ (.Y(_03177_),
    .B1(net5324),
    .B2(\TRNG.hash[3] ),
    .A2(net5111),
    .A1(\TRNG.hash[11] ));
 sg13g2_a221oi_1 _19297_ (.B2(\TRNG.hash[19] ),
    .C1(net5513),
    .B1(net5312),
    .A1(\TRNG.hash[27] ),
    .Y(_03178_),
    .A2(net5336));
 sg13g2_a221oi_1 _19298_ (.B2(_03178_),
    .C1(net5511),
    .B1(_03177_),
    .A1(_03175_),
    .Y(_03179_),
    .A2(_03176_));
 sg13g2_a22oi_1 _19299_ (.Y(_03180_),
    .B1(net5322),
    .B2(\TRNG.hash[99] ),
    .A2(net5109),
    .A1(net5894));
 sg13g2_a22oi_1 _19300_ (.Y(_03181_),
    .B1(net5310),
    .B2(net5544),
    .A2(net5334),
    .A1(\TRNG.hash[123] ));
 sg13g2_a21oi_1 _19301_ (.A1(_03180_),
    .A2(_03181_),
    .Y(_03182_),
    .B1(net5304));
 sg13g2_a22oi_1 _19302_ (.Y(_03183_),
    .B1(net5109),
    .B2(\TRNG.hash[75] ),
    .A2(net5339),
    .A1(\TRNG.hash[91] ));
 sg13g2_a22oi_1 _19303_ (.Y(_03184_),
    .B1(net5313),
    .B2(\TRNG.hash[83] ),
    .A2(net5322),
    .A1(\TRNG.hash[67] ));
 sg13g2_a21oi_1 _19304_ (.A1(_03183_),
    .A2(_03184_),
    .Y(_03185_),
    .B1(net5102));
 sg13g2_nor4_2 _19305_ (.A(net5508),
    .B(_03179_),
    .C(_03182_),
    .Y(_03186_),
    .D(_03185_));
 sg13g2_a22oi_1 _19306_ (.Y(_03187_),
    .B1(net5320),
    .B2(\TRNG.hash[131] ),
    .A2(net5107),
    .A1(\TRNG.hash[139] ));
 sg13g2_a221oi_1 _19307_ (.B2(\TRNG.hash[147] ),
    .C1(net5512),
    .B1(net5309),
    .A1(\TRNG.hash[155] ),
    .Y(_03188_),
    .A2(net5332));
 sg13g2_a22oi_1 _19308_ (.Y(_03189_),
    .B1(net5316),
    .B2(\TRNG.hash[163] ),
    .A2(net5106),
    .A1(\TRNG.hash[171] ));
 sg13g2_a221oi_1 _19309_ (.B2(\TRNG.hash[179] ),
    .C1(net5459),
    .B1(net5307),
    .A1(\TRNG.hash[187] ),
    .Y(_03190_),
    .A2(net5330));
 sg13g2_a21o_1 _19310_ (.A2(_03188_),
    .A1(_03187_),
    .B1(net5509),
    .X(_03191_));
 sg13g2_a21oi_1 _19311_ (.A1(_03189_),
    .A2(_03190_),
    .Y(_03192_),
    .B1(_03191_));
 sg13g2_a22oi_1 _19312_ (.Y(_03193_),
    .B1(net5305),
    .B2(\TRNG.hash[211] ),
    .A2(net5317),
    .A1(\TRNG.hash[195] ));
 sg13g2_a22oi_1 _19313_ (.Y(_03194_),
    .B1(net5103),
    .B2(\TRNG.hash[203] ),
    .A2(net5328),
    .A1(\TRNG.hash[219] ));
 sg13g2_a21oi_1 _19314_ (.A1(_03193_),
    .A2(_03194_),
    .Y(_03195_),
    .B1(net5101));
 sg13g2_a22oi_1 _19315_ (.Y(_03196_),
    .B1(net5305),
    .B2(net5560),
    .A2(net5104),
    .A1(\TRNG.hash[235] ));
 sg13g2_a22oi_1 _19316_ (.Y(_03197_),
    .B1(net5318),
    .B2(net5888),
    .A2(net5329),
    .A1(net5558));
 sg13g2_a21oi_1 _19317_ (.A1(_03196_),
    .A2(_03197_),
    .Y(_03198_),
    .B1(net5303));
 sg13g2_nor4_2 _19318_ (.A(_04341_),
    .B(_03192_),
    .C(_03195_),
    .Y(_03199_),
    .D(_03198_));
 sg13g2_nor3_2 _19319_ (.A(net4556),
    .B(_03186_),
    .C(_03199_),
    .Y(_03200_));
 sg13g2_a21o_1 _19320_ (.A2(net4555),
    .A1(net2948),
    .B1(_03200_),
    .X(_01239_));
 sg13g2_a22oi_1 _19321_ (.Y(_03201_),
    .B1(net5316),
    .B2(\TRNG.hash[164] ),
    .A2(net5106),
    .A1(\TRNG.hash[172] ));
 sg13g2_a221oi_1 _19322_ (.B2(\TRNG.hash[180] ),
    .C1(net5459),
    .B1(net5307),
    .A1(\TRNG.hash[188] ),
    .Y(_03202_),
    .A2(net5330));
 sg13g2_and2_1 _19323_ (.A(\TRNG.hash[132] ),
    .B(net5320),
    .X(_03203_));
 sg13g2_a21oi_1 _19324_ (.A1(\TRNG.hash[156] ),
    .A2(net5332),
    .Y(_03204_),
    .B1(net5512));
 sg13g2_a221oi_1 _19325_ (.B2(\TRNG.hash[148] ),
    .C1(_03203_),
    .B1(net5309),
    .A1(\TRNG.hash[140] ),
    .Y(_03205_),
    .A2(net5107));
 sg13g2_a221oi_1 _19326_ (.B2(_03205_),
    .C1(net5509),
    .B1(_03204_),
    .A1(_03201_),
    .Y(_03206_),
    .A2(_03202_));
 sg13g2_a22oi_1 _19327_ (.Y(_03207_),
    .B1(net5317),
    .B2(\TRNG.hash[196] ),
    .A2(net5329),
    .A1(\TRNG.hash[220] ));
 sg13g2_a22oi_1 _19328_ (.Y(_03208_),
    .B1(net5306),
    .B2(\TRNG.hash[212] ),
    .A2(net5104),
    .A1(\TRNG.hash[204] ));
 sg13g2_a21oi_1 _19329_ (.A1(_03207_),
    .A2(_03208_),
    .Y(_03209_),
    .B1(net5101));
 sg13g2_a22oi_1 _19330_ (.Y(_03210_),
    .B1(net5317),
    .B2(net5887),
    .A2(net5103),
    .A1(net5885));
 sg13g2_a22oi_1 _19331_ (.Y(_03211_),
    .B1(net5306),
    .B2(net5882),
    .A2(net5329),
    .A1(net5877));
 sg13g2_a21oi_1 _19332_ (.A1(_03210_),
    .A2(_03211_),
    .Y(_03212_),
    .B1(net5303));
 sg13g2_nor4_2 _19333_ (.A(_04341_),
    .B(_03206_),
    .C(_03209_),
    .Y(_03213_),
    .D(_03212_));
 sg13g2_a22oi_1 _19334_ (.Y(_03214_),
    .B1(net5325),
    .B2(\TRNG.hash[36] ),
    .A2(net5112),
    .A1(\TRNG.hash[44] ));
 sg13g2_a221oi_1 _19335_ (.B2(\TRNG.hash[52] ),
    .C1(net5460),
    .B1(net5313),
    .A1(\TRNG.hash[60] ),
    .Y(_03215_),
    .A2(net5337));
 sg13g2_a22oi_1 _19336_ (.Y(_03216_),
    .B1(net5313),
    .B2(\TRNG.hash[20] ),
    .A2(net5337),
    .A1(\TRNG.hash[28] ));
 sg13g2_a221oi_1 _19337_ (.B2(\TRNG.hash[4] ),
    .C1(net5514),
    .B1(net5325),
    .A1(\TRNG.hash[12] ),
    .Y(_03217_),
    .A2(net5112));
 sg13g2_a221oi_1 _19338_ (.B2(_03217_),
    .C1(net5511),
    .B1(_03216_),
    .A1(_03214_),
    .Y(_03218_),
    .A2(_03215_));
 sg13g2_a22oi_1 _19339_ (.Y(_03219_),
    .B1(net5311),
    .B2(\TRNG.hash[84] ),
    .A2(net5335),
    .A1(\TRNG.hash[92] ));
 sg13g2_a22oi_1 _19340_ (.Y(_03220_),
    .B1(net5327),
    .B2(\TRNG.hash[68] ),
    .A2(net5114),
    .A1(\TRNG.hash[76] ));
 sg13g2_a21oi_1 _19341_ (.A1(_03219_),
    .A2(_03220_),
    .Y(_03221_),
    .B1(net5102));
 sg13g2_a22oi_1 _19342_ (.Y(_03222_),
    .B1(net5110),
    .B2(net5548),
    .A2(net5335),
    .A1(\TRNG.hash[124] ));
 sg13g2_a22oi_1 _19343_ (.Y(_03223_),
    .B1(net5311),
    .B2(net5890),
    .A2(net5323),
    .A1(\TRNG.hash[100] ));
 sg13g2_a21oi_1 _19344_ (.A1(_03222_),
    .A2(_03223_),
    .Y(_03224_),
    .B1(net5304));
 sg13g2_nor4_2 _19345_ (.A(net5508),
    .B(_03218_),
    .C(_03221_),
    .Y(_03225_),
    .D(_03224_));
 sg13g2_nor3_2 _19346_ (.A(net4556),
    .B(_03213_),
    .C(_03225_),
    .Y(_03226_));
 sg13g2_a21o_1 _19347_ (.A2(net4555),
    .A1(net2658),
    .B1(_03226_),
    .X(_01240_));
 sg13g2_a22oi_1 _19348_ (.Y(_03227_),
    .B1(net5313),
    .B2(\TRNG.hash[53] ),
    .A2(net5337),
    .A1(\TRNG.hash[61] ));
 sg13g2_a22oi_1 _19349_ (.Y(_03228_),
    .B1(net5325),
    .B2(\TRNG.hash[37] ),
    .A2(net5112),
    .A1(\TRNG.hash[45] ));
 sg13g2_nand3_1 _19350_ (.B(_03227_),
    .C(_03228_),
    .A(net5513),
    .Y(_03229_));
 sg13g2_a22oi_1 _19351_ (.Y(_03230_),
    .B1(net5324),
    .B2(\TRNG.hash[5] ),
    .A2(net5336),
    .A1(\TRNG.hash[29] ));
 sg13g2_a221oi_1 _19352_ (.B2(\TRNG.hash[21] ),
    .C1(net5513),
    .B1(net5312),
    .A1(\TRNG.hash[13] ),
    .Y(_03231_),
    .A2(net5111));
 sg13g2_a21oi_1 _19353_ (.A1(_03230_),
    .A2(_03231_),
    .Y(_03232_),
    .B1(net5511));
 sg13g2_nand2_2 _19354_ (.Y(_03233_),
    .A(_03229_),
    .B(_03232_));
 sg13g2_a22oi_1 _19355_ (.Y(_03234_),
    .B1(net5311),
    .B2(\TRNG.hash[85] ),
    .A2(net5335),
    .A1(\TRNG.hash[93] ));
 sg13g2_a22oi_1 _19356_ (.Y(_03235_),
    .B1(net5327),
    .B2(\TRNG.hash[69] ),
    .A2(net5114),
    .A1(\TRNG.hash[77] ));
 sg13g2_a21oi_1 _19357_ (.A1(_03234_),
    .A2(_03235_),
    .Y(_03236_),
    .B1(net5102));
 sg13g2_a22oi_1 _19358_ (.Y(_03237_),
    .B1(net5110),
    .B2(net5893),
    .A2(net5334),
    .A1(\TRNG.hash[125] ));
 sg13g2_a22oi_1 _19359_ (.Y(_03238_),
    .B1(net5311),
    .B2(net5889),
    .A2(net5323),
    .A1(net5550));
 sg13g2_a21oi_1 _19360_ (.A1(_03237_),
    .A2(_03238_),
    .Y(_03239_),
    .B1(net5304));
 sg13g2_nor3_1 _19361_ (.A(net5508),
    .B(_03236_),
    .C(_03239_),
    .Y(_03240_));
 sg13g2_a22oi_1 _19362_ (.Y(_03241_),
    .B1(net5319),
    .B2(\TRNG.hash[165] ),
    .A2(net5106),
    .A1(\TRNG.hash[173] ));
 sg13g2_a221oi_1 _19363_ (.B2(\TRNG.hash[181] ),
    .C1(net5460),
    .B1(net5309),
    .A1(\TRNG.hash[189] ),
    .Y(_03242_),
    .A2(net5333));
 sg13g2_a22oi_1 _19364_ (.Y(_03243_),
    .B1(net5320),
    .B2(\TRNG.hash[133] ),
    .A2(net5107),
    .A1(\TRNG.hash[141] ));
 sg13g2_a22oi_1 _19365_ (.Y(_03244_),
    .B1(net5309),
    .B2(\TRNG.hash[149] ),
    .A2(net5340),
    .A1(\TRNG.hash[157] ));
 sg13g2_nand3_1 _19366_ (.B(_03243_),
    .C(_03244_),
    .A(net5459),
    .Y(_03245_));
 sg13g2_a21oi_1 _19367_ (.A1(_03241_),
    .A2(_03242_),
    .Y(_03246_),
    .B1(net5510));
 sg13g2_nand2_1 _19368_ (.Y(_03247_),
    .A(_03245_),
    .B(_03246_));
 sg13g2_a22oi_1 _19369_ (.Y(_03248_),
    .B1(net5306),
    .B2(\TRNG.hash[213] ),
    .A2(net5108),
    .A1(\TRNG.hash[205] ));
 sg13g2_a22oi_1 _19370_ (.Y(_03249_),
    .B1(net5321),
    .B2(\TRNG.hash[197] ),
    .A2(net5329),
    .A1(\TRNG.hash[221] ));
 sg13g2_a21oi_1 _19371_ (.A1(_03248_),
    .A2(_03249_),
    .Y(_03250_),
    .B1(net5101));
 sg13g2_a22oi_1 _19372_ (.Y(_03251_),
    .B1(net5306),
    .B2(net5881),
    .A2(net5328),
    .A1(net5557));
 sg13g2_a22oi_1 _19373_ (.Y(_03252_),
    .B1(net5317),
    .B2(net5567),
    .A2(net5103),
    .A1(net5563));
 sg13g2_a21oi_1 _19374_ (.A1(_03251_),
    .A2(_03252_),
    .Y(_03253_),
    .B1(net5303));
 sg13g2_nor3_2 _19375_ (.A(_04341_),
    .B(_03250_),
    .C(_03253_),
    .Y(_03254_));
 sg13g2_a22oi_1 _19376_ (.Y(_03255_),
    .B1(_03247_),
    .B2(_03254_),
    .A2(_03240_),
    .A1(_03233_));
 sg13g2_mux2_1 _19377_ (.A0(_03255_),
    .A1(net2760),
    .S(net4555),
    .X(_01241_));
 sg13g2_a22oi_1 _19378_ (.Y(_03256_),
    .B1(net5324),
    .B2(\TRNG.hash[6] ),
    .A2(net5111),
    .A1(\TRNG.hash[14] ));
 sg13g2_a221oi_1 _19379_ (.B2(\TRNG.hash[22] ),
    .C1(net5513),
    .B1(net5312),
    .A1(\TRNG.hash[30] ),
    .Y(_03257_),
    .A2(net5336));
 sg13g2_and2_1 _19380_ (.A(\TRNG.hash[62] ),
    .B(net5338),
    .X(_03258_));
 sg13g2_a21oi_1 _19381_ (.A1(\TRNG.hash[46] ),
    .A2(net5112),
    .Y(_03259_),
    .B1(net5460));
 sg13g2_a221oi_1 _19382_ (.B2(\TRNG.hash[54] ),
    .C1(_03258_),
    .B1(net5313),
    .A1(\TRNG.hash[38] ),
    .Y(_03260_),
    .A2(net5324));
 sg13g2_a221oi_1 _19383_ (.B2(_03260_),
    .C1(net5511),
    .B1(_03259_),
    .A1(_03256_),
    .Y(_03261_),
    .A2(_03257_));
 sg13g2_a22oi_1 _19384_ (.Y(_03262_),
    .B1(net5310),
    .B2(\TRNG.hash[86] ),
    .A2(net5110),
    .A1(\TRNG.hash[78] ));
 sg13g2_a22oi_1 _19385_ (.Y(_03263_),
    .B1(net5322),
    .B2(\TRNG.hash[70] ),
    .A2(net5338),
    .A1(\TRNG.hash[94] ));
 sg13g2_a21oi_1 _19386_ (.A1(_03262_),
    .A2(_03263_),
    .Y(_03264_),
    .B1(net5102));
 sg13g2_a22oi_1 _19387_ (.Y(_03265_),
    .B1(net5323),
    .B2(net5549),
    .A2(net5335),
    .A1(\TRNG.hash[126] ));
 sg13g2_a22oi_1 _19388_ (.Y(_03266_),
    .B1(net5311),
    .B2(\TRNG.hash[118] ),
    .A2(net5109),
    .A1(net5547));
 sg13g2_a21oi_1 _19389_ (.A1(_03265_),
    .A2(_03266_),
    .Y(_03267_),
    .B1(net5304));
 sg13g2_nor4_2 _19390_ (.A(net5508),
    .B(_03261_),
    .C(_03264_),
    .Y(_03268_),
    .D(_03267_));
 sg13g2_and2_1 _19391_ (.A(\TRNG.hash[182] ),
    .B(net5308),
    .X(_03269_));
 sg13g2_a21oi_1 _19392_ (.A1(\TRNG.hash[174] ),
    .A2(net5105),
    .Y(_03270_),
    .B1(net5459));
 sg13g2_a221oi_1 _19393_ (.B2(\TRNG.hash[166] ),
    .C1(_03269_),
    .B1(net5321),
    .A1(\TRNG.hash[190] ),
    .Y(_03271_),
    .A2(net5331));
 sg13g2_a22oi_1 _19394_ (.Y(_03272_),
    .B1(net5320),
    .B2(\TRNG.hash[134] ),
    .A2(net5332),
    .A1(\TRNG.hash[158] ));
 sg13g2_a221oi_1 _19395_ (.B2(\TRNG.hash[150] ),
    .C1(net5512),
    .B1(net5307),
    .A1(\TRNG.hash[142] ),
    .Y(_03273_),
    .A2(net5108));
 sg13g2_a221oi_1 _19396_ (.B2(_03273_),
    .C1(net5509),
    .B1(_03272_),
    .A1(_03270_),
    .Y(_03274_),
    .A2(_03271_));
 sg13g2_a22oi_1 _19397_ (.Y(_03275_),
    .B1(net5317),
    .B2(net5566),
    .A2(net5328),
    .A1(net5556));
 sg13g2_a22oi_1 _19398_ (.Y(_03276_),
    .B1(net5307),
    .B2(\TRNG.hash[246] ),
    .A2(net5103),
    .A1(net5562));
 sg13g2_a21oi_1 _19399_ (.A1(_03275_),
    .A2(_03276_),
    .Y(_03277_),
    .B1(net5303));
 sg13g2_a22oi_1 _19400_ (.Y(_03278_),
    .B1(net5308),
    .B2(\TRNG.hash[214] ),
    .A2(net5331),
    .A1(\TRNG.hash[222] ));
 sg13g2_a22oi_1 _19401_ (.Y(_03279_),
    .B1(net5316),
    .B2(\TRNG.hash[198] ),
    .A2(net5106),
    .A1(\TRNG.hash[206] ));
 sg13g2_a21oi_1 _19402_ (.A1(_03278_),
    .A2(_03279_),
    .Y(_03280_),
    .B1(net5101));
 sg13g2_nor4_2 _19403_ (.A(_04341_),
    .B(_03274_),
    .C(_03277_),
    .Y(_03281_),
    .D(_03280_));
 sg13g2_nor3_2 _19404_ (.A(net4555),
    .B(_03268_),
    .C(_03281_),
    .Y(_03282_));
 sg13g2_a21o_1 _19405_ (.A2(net4555),
    .A1(net2560),
    .B1(_03282_),
    .X(_01242_));
 sg13g2_a21oi_1 _19406_ (.A1(\TRNG.hash[183] ),
    .A2(net5308),
    .Y(_03283_),
    .B1(net5459));
 sg13g2_and2_1 _19407_ (.A(\TRNG.hash[191] ),
    .B(net5331),
    .X(_03284_));
 sg13g2_a221oi_1 _19408_ (.B2(\TRNG.hash[167] ),
    .C1(_03284_),
    .B1(net5321),
    .A1(\TRNG.hash[175] ),
    .Y(_03285_),
    .A2(net5108));
 sg13g2_a22oi_1 _19409_ (.Y(_03286_),
    .B1(net5321),
    .B2(\TRNG.hash[135] ),
    .A2(net5333),
    .A1(\TRNG.hash[159] ));
 sg13g2_a221oi_1 _19410_ (.B2(\TRNG.hash[151] ),
    .C1(net5512),
    .B1(net5307),
    .A1(\TRNG.hash[143] ),
    .Y(_03287_),
    .A2(net5108));
 sg13g2_a221oi_1 _19411_ (.B2(_03287_),
    .C1(net5509),
    .B1(_03286_),
    .A1(_03283_),
    .Y(_03288_),
    .A2(_03285_));
 sg13g2_a22oi_1 _19412_ (.Y(_03289_),
    .B1(net5306),
    .B2(\TRNG.hash[215] ),
    .A2(net5321),
    .A1(\TRNG.hash[199] ));
 sg13g2_a22oi_1 _19413_ (.Y(_03290_),
    .B1(net5108),
    .B2(\TRNG.hash[207] ),
    .A2(net5329),
    .A1(\TRNG.hash[223] ));
 sg13g2_a21oi_1 _19414_ (.A1(_03289_),
    .A2(_03290_),
    .Y(_03291_),
    .B1(net5101));
 sg13g2_a22oi_1 _19415_ (.Y(_03292_),
    .B1(net5306),
    .B2(net5880),
    .A2(net5104),
    .A1(net5561));
 sg13g2_a22oi_1 _19416_ (.Y(_03293_),
    .B1(net5317),
    .B2(\TRNG.hash[231] ),
    .A2(net5328),
    .A1(\TRNG.hash[255] ));
 sg13g2_a21oi_1 _19417_ (.A1(_03292_),
    .A2(_03293_),
    .Y(_03294_),
    .B1(net5303));
 sg13g2_nor4_2 _19418_ (.A(_04341_),
    .B(_03288_),
    .C(_03291_),
    .Y(_03295_),
    .D(_03294_));
 sg13g2_a21oi_1 _19419_ (.A1(\TRNG.hash[47] ),
    .A2(net5112),
    .Y(_03296_),
    .B1(net5460));
 sg13g2_and2_1 _19420_ (.A(\TRNG.hash[39] ),
    .B(net5325),
    .X(_03297_));
 sg13g2_a221oi_1 _19421_ (.B2(\TRNG.hash[55] ),
    .C1(_03297_),
    .B1(net5312),
    .A1(\TRNG.hash[63] ),
    .Y(_03298_),
    .A2(net5336));
 sg13g2_a22oi_1 _19422_ (.Y(_03299_),
    .B1(net5324),
    .B2(\TRNG.hash[7] ),
    .A2(net5336),
    .A1(\TRNG.hash[31] ));
 sg13g2_a221oi_1 _19423_ (.B2(\TRNG.hash[23] ),
    .C1(net5513),
    .B1(net5312),
    .A1(\TRNG.hash[15] ),
    .Y(_03300_),
    .A2(net5112));
 sg13g2_a221oi_1 _19424_ (.B2(_03300_),
    .C1(net5511),
    .B1(_03299_),
    .A1(_03296_),
    .Y(_03301_),
    .A2(_03298_));
 sg13g2_a22oi_1 _19425_ (.Y(_03302_),
    .B1(net5311),
    .B2(\TRNG.hash[119] ),
    .A2(net5322),
    .A1(\TRNG.hash[103] ));
 sg13g2_a22oi_1 _19426_ (.Y(_03303_),
    .B1(net5109),
    .B2(net5892),
    .A2(net5334),
    .A1(\TRNG.hash[127] ));
 sg13g2_a21oi_1 _19427_ (.A1(_03302_),
    .A2(_03303_),
    .Y(_03304_),
    .B1(net5304));
 sg13g2_a22oi_1 _19428_ (.Y(_03305_),
    .B1(net5311),
    .B2(\TRNG.hash[87] ),
    .A2(net5110),
    .A1(\TRNG.hash[79] ));
 sg13g2_a22oi_1 _19429_ (.Y(_03306_),
    .B1(net5323),
    .B2(\TRNG.hash[71] ),
    .A2(net5338),
    .A1(\TRNG.hash[95] ));
 sg13g2_a21oi_1 _19430_ (.A1(_03305_),
    .A2(_03306_),
    .Y(_03307_),
    .B1(net5102));
 sg13g2_nor4_2 _19431_ (.A(net5508),
    .B(_03301_),
    .C(_03304_),
    .Y(_03308_),
    .D(_03307_));
 sg13g2_nor3_2 _19432_ (.A(net4555),
    .B(_03295_),
    .C(_03308_),
    .Y(_03309_));
 sg13g2_a21o_1 _19433_ (.A2(net4555),
    .A1(net2830),
    .B1(_03309_),
    .X(_01243_));
 sg13g2_nand2b_1 _19434_ (.Y(_03310_),
    .B(_04891_),
    .A_N(_04853_));
 sg13g2_nand3_1 _19435_ (.B(net5237),
    .C(net4790),
    .A(net2880),
    .Y(_03311_));
 sg13g2_o21ai_1 _19436_ (.B1(_03311_),
    .Y(_01244_),
    .A1(_04381_),
    .A2(net4770));
 sg13g2_nand3_1 _19437_ (.B(net5232),
    .C(net4770),
    .A(net1864),
    .Y(_03312_));
 sg13g2_o21ai_1 _19438_ (.B1(_03312_),
    .Y(_01245_),
    .A1(_04382_),
    .A2(net4770));
 sg13g2_nand3_1 _19439_ (.B(net5233),
    .C(net4789),
    .A(net3085),
    .Y(_03313_));
 sg13g2_o21ai_1 _19440_ (.B1(_03313_),
    .Y(_01246_),
    .A1(_04383_),
    .A2(net4780));
 sg13g2_nand3_1 _19441_ (.B(net5233),
    .C(net4780),
    .A(net2611),
    .Y(_03314_));
 sg13g2_o21ai_1 _19442_ (.B1(_03314_),
    .Y(_01247_),
    .A1(_04384_),
    .A2(net4781));
 sg13g2_nand3_1 _19443_ (.B(net5234),
    .C(net4782),
    .A(net3209),
    .Y(_03315_));
 sg13g2_o21ai_1 _19444_ (.B1(_03315_),
    .Y(_01248_),
    .A1(_04385_),
    .A2(net4880));
 sg13g2_nand3_1 _19445_ (.B(net5285),
    .C(net4880),
    .A(net1937),
    .Y(_03316_));
 sg13g2_o21ai_1 _19446_ (.B1(_03316_),
    .Y(_01249_),
    .A1(_04386_),
    .A2(net4880));
 sg13g2_nand3_1 _19447_ (.B(net5283),
    .C(net4879),
    .A(net2606),
    .Y(_03317_));
 sg13g2_o21ai_1 _19448_ (.B1(_03317_),
    .Y(_01250_),
    .A1(_04387_),
    .A2(net4886));
 sg13g2_nand3_1 _19449_ (.B(net5287),
    .C(net4885),
    .A(net1820),
    .Y(_03318_));
 sg13g2_o21ai_1 _19450_ (.B1(_03318_),
    .Y(_01251_),
    .A1(_04388_),
    .A2(net4886));
 sg13g2_nand3_1 _19451_ (.B(net5288),
    .C(net4887),
    .A(net1193),
    .Y(_03319_));
 sg13g2_o21ai_1 _19452_ (.B1(_03319_),
    .Y(_01252_),
    .A1(_04389_),
    .A2(net4887));
 sg13g2_nand3_1 _19453_ (.B(net5288),
    .C(net4887),
    .A(net2909),
    .Y(_03320_));
 sg13g2_o21ai_1 _19454_ (.B1(_03320_),
    .Y(_01253_),
    .A1(_04390_),
    .A2(net4871));
 sg13g2_nand3_1 _19455_ (.B(net5281),
    .C(net4873),
    .A(net1718),
    .Y(_03321_));
 sg13g2_o21ai_1 _19456_ (.B1(_03321_),
    .Y(_01254_),
    .A1(_04391_),
    .A2(net4873));
 sg13g2_nand3_1 _19457_ (.B(net5281),
    .C(net4872),
    .A(net2615),
    .Y(_03322_));
 sg13g2_o21ai_1 _19458_ (.B1(_03322_),
    .Y(_01255_),
    .A1(_04392_),
    .A2(net4869));
 sg13g2_nand3_1 _19459_ (.B(net5278),
    .C(net4866),
    .A(net2690),
    .Y(_03323_));
 sg13g2_o21ai_1 _19460_ (.B1(_03323_),
    .Y(_01256_),
    .A1(_04393_),
    .A2(net4824));
 sg13g2_nand3_1 _19461_ (.B(net5254),
    .C(net4821),
    .A(net3087),
    .Y(_03324_));
 sg13g2_o21ai_1 _19462_ (.B1(_03324_),
    .Y(_01257_),
    .A1(_04394_),
    .A2(net4821));
 sg13g2_nand3_1 _19463_ (.B(net5252),
    .C(net4820),
    .A(net1229),
    .Y(_03325_));
 sg13g2_o21ai_1 _19464_ (.B1(_03325_),
    .Y(_01258_),
    .A1(_04395_),
    .A2(net4818));
 sg13g2_nand3_1 _19465_ (.B(net5253),
    .C(net4819),
    .A(net1601),
    .Y(_03326_));
 sg13g2_o21ai_1 _19466_ (.B1(_03326_),
    .Y(_01259_),
    .A1(_04396_),
    .A2(net4846));
 sg13g2_nand3_1 _19467_ (.B(net5269),
    .C(net4846),
    .A(net1362),
    .Y(_03327_));
 sg13g2_o21ai_1 _19468_ (.B1(_03327_),
    .Y(_01260_),
    .A1(_04397_),
    .A2(net4848));
 sg13g2_nand3_1 _19469_ (.B(net5262),
    .C(net4835),
    .A(net1984),
    .Y(_03328_));
 sg13g2_o21ai_1 _19470_ (.B1(_03328_),
    .Y(_01261_),
    .A1(_04398_),
    .A2(net4834));
 sg13g2_nand3_1 _19471_ (.B(net5259),
    .C(net4830),
    .A(net1978),
    .Y(_03329_));
 sg13g2_o21ai_1 _19472_ (.B1(_03329_),
    .Y(_01262_),
    .A1(_04399_),
    .A2(net4831));
 sg13g2_nand3_1 _19473_ (.B(net5260),
    .C(net4830),
    .A(net2469),
    .Y(_03330_));
 sg13g2_o21ai_1 _19474_ (.B1(_03330_),
    .Y(_01263_),
    .A1(_04400_),
    .A2(net4828));
 sg13g2_nand3_1 _19475_ (.B(net5260),
    .C(net4831),
    .A(net3116),
    .Y(_03331_));
 sg13g2_o21ai_1 _19476_ (.B1(_03331_),
    .Y(_01264_),
    .A1(_04401_),
    .A2(net4802));
 sg13g2_nand3_1 _19477_ (.B(net5243),
    .C(net4802),
    .A(net2757),
    .Y(_03332_));
 sg13g2_o21ai_1 _19478_ (.B1(_03332_),
    .Y(_01265_),
    .A1(_04402_),
    .A2(net4800));
 sg13g2_nand3_1 _19479_ (.B(net5244),
    .C(net4800),
    .A(net2548),
    .Y(_03333_));
 sg13g2_o21ai_1 _19480_ (.B1(_03333_),
    .Y(_01266_),
    .A1(_04403_),
    .A2(net4792));
 sg13g2_nand3_1 _19481_ (.B(net5240),
    .C(net4793),
    .A(net2129),
    .Y(_03334_));
 sg13g2_o21ai_1 _19482_ (.B1(_03334_),
    .Y(_01267_),
    .A1(_04404_),
    .A2(net4791));
 sg13g2_nand3_1 _19483_ (.B(net5239),
    .C(net4793),
    .A(net2622),
    .Y(_03335_));
 sg13g2_o21ai_1 _19484_ (.B1(_03335_),
    .Y(_01268_),
    .A1(_04405_),
    .A2(net4794));
 sg13g2_nand3_1 _19485_ (.B(net5241),
    .C(net4794),
    .A(net1150),
    .Y(_03336_));
 sg13g2_o21ai_1 _19486_ (.B1(_03336_),
    .Y(_01269_),
    .A1(_04406_),
    .A2(net4795));
 sg13g2_nand3_1 _19487_ (.B(net5221),
    .C(net4754),
    .A(net3182),
    .Y(_03337_));
 sg13g2_o21ai_1 _19488_ (.B1(_03337_),
    .Y(_01270_),
    .A1(_04407_),
    .A2(net4758));
 sg13g2_nand3_1 _19489_ (.B(net5223),
    .C(net4758),
    .A(net2280),
    .Y(_03338_));
 sg13g2_o21ai_1 _19490_ (.B1(_03338_),
    .Y(_01271_),
    .A1(_04408_),
    .A2(net4758));
 sg13g2_nand3_1 _19491_ (.B(net5223),
    .C(net4762),
    .A(net2819),
    .Y(_03339_));
 sg13g2_o21ai_1 _19492_ (.B1(_03339_),
    .Y(_01272_),
    .A1(_04409_),
    .A2(net4763));
 sg13g2_nand3_1 _19493_ (.B(net5224),
    .C(net4763),
    .A(net3189),
    .Y(_03340_));
 sg13g2_o21ai_1 _19494_ (.B1(_03340_),
    .Y(_01273_),
    .A1(_04410_),
    .A2(net4764));
 sg13g2_nand3_1 _19495_ (.B(net5227),
    .C(net4771),
    .A(net1231),
    .Y(_03341_));
 sg13g2_o21ai_1 _19496_ (.B1(_03341_),
    .Y(_01274_),
    .A1(_04411_),
    .A2(net4771));
 sg13g2_nand3_1 _19497_ (.B(net5227),
    .C(net4768),
    .A(net1191),
    .Y(_03342_));
 sg13g2_o21ai_1 _19498_ (.B1(_03342_),
    .Y(_01275_),
    .A1(_04412_),
    .A2(net4768));
 sg13g2_nand3_1 _19499_ (.B(net5229),
    .C(net4770),
    .A(net2486),
    .Y(_03343_));
 sg13g2_o21ai_1 _19500_ (.B1(_03343_),
    .Y(_01276_),
    .A1(_04413_),
    .A2(net4770));
 sg13g2_nand3_1 _19501_ (.B(net5229),
    .C(net4776),
    .A(net2573),
    .Y(_03344_));
 sg13g2_o21ai_1 _19502_ (.B1(_03344_),
    .Y(_01277_),
    .A1(_04414_),
    .A2(net4776));
 sg13g2_nand3_1 _19503_ (.B(net5233),
    .C(net4780),
    .A(net2709),
    .Y(_03345_));
 sg13g2_o21ai_1 _19504_ (.B1(_03345_),
    .Y(_01278_),
    .A1(_04415_),
    .A2(net4781));
 sg13g2_nand3_1 _19505_ (.B(net5235),
    .C(net4784),
    .A(net3199),
    .Y(_03346_));
 sg13g2_o21ai_1 _19506_ (.B1(_03346_),
    .Y(_01279_),
    .A1(_04416_),
    .A2(net4784));
 sg13g2_nand3_1 _19507_ (.B(net5236),
    .C(net4787),
    .A(net2113),
    .Y(_03347_));
 sg13g2_o21ai_1 _19508_ (.B1(_03347_),
    .Y(_01280_),
    .A1(_04417_),
    .A2(net4787));
 sg13g2_nand3_1 _19509_ (.B(net5285),
    .C(net4881),
    .A(net1223),
    .Y(_03348_));
 sg13g2_o21ai_1 _19510_ (.B1(_03348_),
    .Y(_01281_),
    .A1(_04418_),
    .A2(net4881));
 sg13g2_nand3_1 _19511_ (.B(net5289),
    .C(net4890),
    .A(net2549),
    .Y(_03349_));
 sg13g2_o21ai_1 _19512_ (.B1(_03349_),
    .Y(_01282_),
    .A1(_04419_),
    .A2(net4890));
 sg13g2_nand3_1 _19513_ (.B(net5290),
    .C(net4892),
    .A(net1239),
    .Y(_03350_));
 sg13g2_o21ai_1 _19514_ (.B1(_03350_),
    .Y(_01283_),
    .A1(_04420_),
    .A2(net4892));
 sg13g2_nand3_1 _19515_ (.B(net5298),
    .C(net4910),
    .A(net2510),
    .Y(_03351_));
 sg13g2_o21ai_1 _19516_ (.B1(_03351_),
    .Y(_01284_),
    .A1(_04421_),
    .A2(net4912));
 sg13g2_nand3_1 _19517_ (.B(net5299),
    .C(net4910),
    .A(net1653),
    .Y(_03352_));
 sg13g2_o21ai_1 _19518_ (.B1(_03352_),
    .Y(_01285_),
    .A1(_04422_),
    .A2(net4910));
 sg13g2_nand3_1 _19519_ (.B(net5299),
    .C(net4910),
    .A(net3120),
    .Y(_03353_));
 sg13g2_o21ai_1 _19520_ (.B1(_03353_),
    .Y(_01286_),
    .A1(_04423_),
    .A2(net4906));
 sg13g2_nand3_1 _19521_ (.B(net5300),
    .C(net4906),
    .A(net2850),
    .Y(_03354_));
 sg13g2_o21ai_1 _19522_ (.B1(_03354_),
    .Y(_01287_),
    .A1(_04424_),
    .A2(net4900));
 sg13g2_nand3_1 _19523_ (.B(net5295),
    .C(net4900),
    .A(net2586),
    .Y(_03355_));
 sg13g2_o21ai_1 _19524_ (.B1(_03355_),
    .Y(_01288_),
    .A1(_04425_),
    .A2(net4896));
 sg13g2_nand3_1 _19525_ (.B(net5295),
    .C(net4896),
    .A(net2268),
    .Y(_03356_));
 sg13g2_o21ai_1 _19526_ (.B1(_03356_),
    .Y(_01289_),
    .A1(_04426_),
    .A2(net4896));
 sg13g2_nand3_1 _19527_ (.B(net5270),
    .C(net4852),
    .A(net2112),
    .Y(_03357_));
 sg13g2_o21ai_1 _19528_ (.B1(_03357_),
    .Y(_01290_),
    .A1(_04427_),
    .A2(net4852));
 sg13g2_nand3_1 _19529_ (.B(net5271),
    .C(net4853),
    .A(net1821),
    .Y(_03358_));
 sg13g2_o21ai_1 _19530_ (.B1(_03358_),
    .Y(_01291_),
    .A1(_04428_),
    .A2(net4852));
 sg13g2_nand3_1 _19531_ (.B(net5271),
    .C(net4852),
    .A(net2462),
    .Y(_03359_));
 sg13g2_o21ai_1 _19532_ (.B1(_03359_),
    .Y(_01292_),
    .A1(_04429_),
    .A2(net4849));
 sg13g2_nand3_1 _19533_ (.B(net5273),
    .C(net4854),
    .A(net2939),
    .Y(_03360_));
 sg13g2_o21ai_1 _19534_ (.B1(_03360_),
    .Y(_01293_),
    .A1(_04430_),
    .A2(net4842));
 sg13g2_nand3_1 _19535_ (.B(net5262),
    .C(net4834),
    .A(net2351),
    .Y(_03361_));
 sg13g2_o21ai_1 _19536_ (.B1(_03361_),
    .Y(_01294_),
    .A1(_04431_),
    .A2(net4835));
 sg13g2_nand3_1 _19537_ (.B(net5262),
    .C(net4834),
    .A(net2108),
    .Y(_03362_));
 sg13g2_o21ai_1 _19538_ (.B1(_03362_),
    .Y(_01295_),
    .A1(_04432_),
    .A2(net4832));
 sg13g2_nand3_1 _19539_ (.B(net5261),
    .C(net4832),
    .A(net3093),
    .Y(_03363_));
 sg13g2_o21ai_1 _19540_ (.B1(_03363_),
    .Y(_01296_),
    .A1(_04433_),
    .A2(net4805));
 sg13g2_nand3_1 _19541_ (.B(net5246),
    .C(net4805),
    .A(net2244),
    .Y(_03364_));
 sg13g2_o21ai_1 _19542_ (.B1(_03364_),
    .Y(_01297_),
    .A1(_04434_),
    .A2(net4803));
 sg13g2_nand3_1 _19543_ (.B(net5245),
    .C(net4803),
    .A(net1941),
    .Y(_03365_));
 sg13g2_o21ai_1 _19544_ (.B1(_03365_),
    .Y(_01298_),
    .A1(_04435_),
    .A2(net4804));
 sg13g2_nand3_1 _19545_ (.B(net5245),
    .C(net4804),
    .A(net2506),
    .Y(_03366_));
 sg13g2_o21ai_1 _19546_ (.B1(_03366_),
    .Y(_01299_),
    .A1(_04436_),
    .A2(net4796));
 sg13g2_nand3_1 _19547_ (.B(net5241),
    .C(net4796),
    .A(net1722),
    .Y(_03367_));
 sg13g2_o21ai_1 _19548_ (.B1(_03367_),
    .Y(_01300_),
    .A1(_04437_),
    .A2(net4753));
 sg13g2_nand3_1 _19549_ (.B(net5220),
    .C(net4754),
    .A(net2235),
    .Y(_03368_));
 sg13g2_o21ai_1 _19550_ (.B1(_03368_),
    .Y(_01301_),
    .A1(_04438_),
    .A2(net4753));
 sg13g2_nand3_1 _19551_ (.B(net5223),
    .C(net4760),
    .A(net2938),
    .Y(_03369_));
 sg13g2_o21ai_1 _19552_ (.B1(_03369_),
    .Y(_01302_),
    .A1(_04439_),
    .A2(net4760));
 sg13g2_nand3_1 _19553_ (.B(net5223),
    .C(net4760),
    .A(net2578),
    .Y(_03370_));
 sg13g2_o21ai_1 _19554_ (.B1(_03370_),
    .Y(_01303_),
    .A1(_04440_),
    .A2(net4763));
 sg13g2_nand3_1 _19555_ (.B(net5224),
    .C(net4763),
    .A(net3298),
    .Y(_03371_));
 sg13g2_o21ai_1 _19556_ (.B1(_03371_),
    .Y(_01304_),
    .A1(_04441_),
    .A2(net4764));
 sg13g2_nand3_1 _19557_ (.B(net5228),
    .C(net4771),
    .A(net1215),
    .Y(_03372_));
 sg13g2_o21ai_1 _19558_ (.B1(_03372_),
    .Y(_01305_),
    .A1(_04442_),
    .A2(net4772));
 sg13g2_nand3_1 _19559_ (.B(net5228),
    .C(net4772),
    .A(net2457),
    .Y(_03373_));
 sg13g2_o21ai_1 _19560_ (.B1(_03373_),
    .Y(_01306_),
    .A1(_04443_),
    .A2(net4773));
 sg13g2_nand3_1 _19561_ (.B(net5227),
    .C(net4774),
    .A(net2106),
    .Y(_03374_));
 sg13g2_o21ai_1 _19562_ (.B1(_03374_),
    .Y(_01307_),
    .A1(_04444_),
    .A2(net4774));
 sg13g2_nand3_1 _19563_ (.B(net5229),
    .C(net4775),
    .A(net1170),
    .Y(_03375_));
 sg13g2_o21ai_1 _19564_ (.B1(_03375_),
    .Y(_01308_),
    .A1(_04445_),
    .A2(net4775));
 sg13g2_nand3_1 _19565_ (.B(net5229),
    .C(net4776),
    .A(net2890),
    .Y(_03376_));
 sg13g2_o21ai_1 _19566_ (.B1(_03376_),
    .Y(_01309_),
    .A1(_04446_),
    .A2(net4789));
 sg13g2_nand3_1 _19567_ (.B(net5233),
    .C(net4781),
    .A(net3165),
    .Y(_03377_));
 sg13g2_o21ai_1 _19568_ (.B1(_03377_),
    .Y(_01310_),
    .A1(_04447_),
    .A2(net4784));
 sg13g2_nand3_1 _19569_ (.B(net5235),
    .C(net4784),
    .A(net1857),
    .Y(_03378_));
 sg13g2_o21ai_1 _19570_ (.B1(_03378_),
    .Y(_01311_),
    .A1(_04448_),
    .A2(net4785));
 sg13g2_nand3_1 _19571_ (.B(net5235),
    .C(net4785),
    .A(net2123),
    .Y(_03379_));
 sg13g2_o21ai_1 _19572_ (.B1(_03379_),
    .Y(_01312_),
    .A1(_04449_),
    .A2(net4785));
 sg13g2_nand3_1 _19573_ (.B(net5235),
    .C(net4787),
    .A(net2773),
    .Y(_03380_));
 sg13g2_o21ai_1 _19574_ (.B1(_03380_),
    .Y(_01313_),
    .A1(_04450_),
    .A2(net4883));
 sg13g2_nand3_1 _19575_ (.B(net5289),
    .C(net4890),
    .A(net2189),
    .Y(_03381_));
 sg13g2_o21ai_1 _19576_ (.B1(_03381_),
    .Y(_01314_),
    .A1(_04451_),
    .A2(net4890));
 sg13g2_nand3_1 _19577_ (.B(net5290),
    .C(net4891),
    .A(net1206),
    .Y(_03382_));
 sg13g2_o21ai_1 _19578_ (.B1(_03382_),
    .Y(_01315_),
    .A1(_04452_),
    .A2(net4892));
 sg13g2_nand3_1 _19579_ (.B(net5298),
    .C(net4909),
    .A(net1577),
    .Y(_03383_));
 sg13g2_o21ai_1 _19580_ (.B1(_03383_),
    .Y(_01316_),
    .A1(_04453_),
    .A2(net4909));
 sg13g2_nand3_1 _19581_ (.B(net5298),
    .C(net4909),
    .A(net1724),
    .Y(_03384_));
 sg13g2_o21ai_1 _19582_ (.B1(_03384_),
    .Y(_01317_),
    .A1(_04454_),
    .A2(net4909));
 sg13g2_nand3_1 _19583_ (.B(net5300),
    .C(net4907),
    .A(net2958),
    .Y(_03385_));
 sg13g2_o21ai_1 _19584_ (.B1(_03385_),
    .Y(_01318_),
    .A1(_04455_),
    .A2(net4900));
 sg13g2_nand3_1 _19585_ (.B(net5294),
    .C(net4900),
    .A(net2153),
    .Y(_03386_));
 sg13g2_o21ai_1 _19586_ (.B1(_03386_),
    .Y(_01319_),
    .A1(_04456_),
    .A2(net4903));
 sg13g2_nand3_1 _19587_ (.B(net5293),
    .C(net4896),
    .A(net3214),
    .Y(_03387_));
 sg13g2_o21ai_1 _19588_ (.B1(_03387_),
    .Y(_01320_),
    .A1(_04457_),
    .A2(net4896));
 sg13g2_nand3_1 _19589_ (.B(net5293),
    .C(net4895),
    .A(net3193),
    .Y(_03388_));
 sg13g2_o21ai_1 _19590_ (.B1(_03388_),
    .Y(_01321_),
    .A1(_04458_),
    .A2(net4822));
 sg13g2_nand3_1 _19591_ (.B(net5254),
    .C(net4822),
    .A(net2474),
    .Y(_03389_));
 sg13g2_o21ai_1 _19592_ (.B1(_03389_),
    .Y(_01322_),
    .A1(_04459_),
    .A2(net4846));
 sg13g2_nand3_1 _19593_ (.B(net5269),
    .C(net4846),
    .A(net1200),
    .Y(_03390_));
 sg13g2_o21ai_1 _19594_ (.B1(_03390_),
    .Y(_01323_),
    .A1(_04460_),
    .A2(net4849));
 sg13g2_nand3_1 _19595_ (.B(net5269),
    .C(net4848),
    .A(net1943),
    .Y(_03391_));
 sg13g2_o21ai_1 _19596_ (.B1(_03391_),
    .Y(_01324_),
    .A1(_04461_),
    .A2(net4848));
 sg13g2_nand3_1 _19597_ (.B(net5273),
    .C(net4854),
    .A(net2099),
    .Y(_03392_));
 sg13g2_o21ai_1 _19598_ (.B1(_03392_),
    .Y(_01325_),
    .A1(_04462_),
    .A2(net4854));
 sg13g2_nand3_1 _19599_ (.B(net5269),
    .C(net4848),
    .A(net2373),
    .Y(_03393_));
 sg13g2_o21ai_1 _19600_ (.B1(_03393_),
    .Y(_01326_),
    .A1(_04463_),
    .A2(net4834));
 sg13g2_nand3_1 _19601_ (.B(net5261),
    .C(net4832),
    .A(net2433),
    .Y(_03394_));
 sg13g2_o21ai_1 _19602_ (.B1(_03394_),
    .Y(_01327_),
    .A1(_04464_),
    .A2(net4833));
 sg13g2_nand3_1 _19603_ (.B(net5261),
    .C(net4846),
    .A(net3158),
    .Y(_03395_));
 sg13g2_o21ai_1 _19604_ (.B1(_03395_),
    .Y(_01328_),
    .A1(_04465_),
    .A2(net4819));
 sg13g2_nand3_1 _19605_ (.B(net5253),
    .C(net4819),
    .A(net2284),
    .Y(_03396_));
 sg13g2_o21ai_1 _19606_ (.B1(_03396_),
    .Y(_01329_),
    .A1(_04466_),
    .A2(net4818));
 sg13g2_nand3_1 _19607_ (.B(net5245),
    .C(net4804),
    .A(net2558),
    .Y(_03397_));
 sg13g2_o21ai_1 _19608_ (.B1(_03397_),
    .Y(_01330_),
    .A1(_04467_),
    .A2(net4804));
 sg13g2_nand3_1 _19609_ (.B(net5245),
    .C(net4797),
    .A(net2211),
    .Y(_03398_));
 sg13g2_o21ai_1 _19610_ (.B1(_03398_),
    .Y(_01331_),
    .A1(_04468_),
    .A2(net4797));
 sg13g2_nand3_1 _19611_ (.B(net5241),
    .C(net4797),
    .A(net1341),
    .Y(_03399_));
 sg13g2_o21ai_1 _19612_ (.B1(_03399_),
    .Y(_01332_),
    .A1(_04469_),
    .A2(net4794));
 sg13g2_nand3_1 _19613_ (.B(net5241),
    .C(net4795),
    .A(net1241),
    .Y(_03400_));
 sg13g2_o21ai_1 _19614_ (.B1(_03400_),
    .Y(_01333_),
    .A1(_04470_),
    .A2(net4795));
 sg13g2_nand3_1 _19615_ (.B(net5247),
    .C(net4809),
    .A(net3344),
    .Y(_03401_));
 sg13g2_o21ai_1 _19616_ (.B1(_03401_),
    .Y(_01334_),
    .A1(_04471_),
    .A2(net4758));
 sg13g2_nand3_1 _19617_ (.B(net5226),
    .C(net4758),
    .A(net2202),
    .Y(_03402_));
 sg13g2_o21ai_1 _19618_ (.B1(_03402_),
    .Y(_01335_),
    .A1(_04472_),
    .A2(net4758));
 sg13g2_nand3_1 _19619_ (.B(net5226),
    .C(net4759),
    .A(net2701),
    .Y(_03403_));
 sg13g2_o21ai_1 _19620_ (.B1(_03403_),
    .Y(_01336_),
    .A1(_04473_),
    .A2(net4759));
 sg13g2_nand3_1 _19621_ (.B(net5224),
    .C(net4764),
    .A(net2978),
    .Y(_03404_));
 sg13g2_o21ai_1 _19622_ (.B1(_03404_),
    .Y(_01337_),
    .A1(_04474_),
    .A2(net4763));
 sg13g2_nand3_1 _19623_ (.B(net5227),
    .C(net4771),
    .A(net1176),
    .Y(_03405_));
 sg13g2_o21ai_1 _19624_ (.B1(_03405_),
    .Y(_01338_),
    .A1(_04475_),
    .A2(net4771));
 sg13g2_nand3_1 _19625_ (.B(net5227),
    .C(net4771),
    .A(net1763),
    .Y(_03406_));
 sg13g2_o21ai_1 _19626_ (.B1(_03406_),
    .Y(_01339_),
    .A1(_04476_),
    .A2(net4771));
 sg13g2_nand3_1 _19627_ (.B(net5227),
    .C(net4772),
    .A(net2058),
    .Y(_03407_));
 sg13g2_o21ai_1 _19628_ (.B1(_03407_),
    .Y(_01340_),
    .A1(_04477_),
    .A2(net4773));
 sg13g2_nand3_1 _19629_ (.B(net5230),
    .C(net4777),
    .A(net2169),
    .Y(_03408_));
 sg13g2_o21ai_1 _19630_ (.B1(_03408_),
    .Y(_01341_),
    .A1(_04478_),
    .A2(net4777));
 sg13g2_nand3_1 _19631_ (.B(net5229),
    .C(net4777),
    .A(net2075),
    .Y(_03409_));
 sg13g2_o21ai_1 _19632_ (.B1(_03409_),
    .Y(_01342_),
    .A1(_04479_),
    .A2(net4778));
 sg13g2_nand3_1 _19633_ (.B(net5234),
    .C(net4782),
    .A(net1816),
    .Y(_03410_));
 sg13g2_o21ai_1 _19634_ (.B1(_03410_),
    .Y(_01343_),
    .A1(_04480_),
    .A2(net4782));
 sg13g2_nand3_1 _19635_ (.B(net5284),
    .C(net4876),
    .A(net3054),
    .Y(_03411_));
 sg13g2_o21ai_1 _19636_ (.B1(_03411_),
    .Y(_01344_),
    .A1(_04481_),
    .A2(net4876));
 sg13g2_nand3_1 _19637_ (.B(net5283),
    .C(net4878),
    .A(net1879),
    .Y(_03412_));
 sg13g2_o21ai_1 _19638_ (.B1(_03412_),
    .Y(_01345_),
    .A1(_04482_),
    .A2(net4878));
 sg13g2_nand3_1 _19639_ (.B(net5283),
    .C(net4878),
    .A(net2253),
    .Y(_03413_));
 sg13g2_o21ai_1 _19640_ (.B1(_03413_),
    .Y(_01346_),
    .A1(_04483_),
    .A2(net4885));
 sg13g2_nand3_1 _19641_ (.B(net5287),
    .C(net4885),
    .A(net1736),
    .Y(_03414_));
 sg13g2_o21ai_1 _19642_ (.B1(_03414_),
    .Y(_01347_),
    .A1(_04484_),
    .A2(net4888));
 sg13g2_nand3_1 _19643_ (.B(net5288),
    .C(net4888),
    .A(net1182),
    .Y(_03415_));
 sg13g2_o21ai_1 _19644_ (.B1(_03415_),
    .Y(_01348_),
    .A1(_04485_),
    .A2(net4888));
 sg13g2_nand3_1 _19645_ (.B(net5297),
    .C(net4904),
    .A(net1643),
    .Y(_03416_));
 sg13g2_o21ai_1 _19646_ (.B1(_03416_),
    .Y(_01349_),
    .A1(_04486_),
    .A2(net4904));
 sg13g2_nand3_1 _19647_ (.B(net5294),
    .C(net4899),
    .A(net2032),
    .Y(_03417_));
 sg13g2_o21ai_1 _19648_ (.B1(_03417_),
    .Y(_01350_),
    .A1(_04487_),
    .A2(net4898));
 sg13g2_nand3_1 _19649_ (.B(net5294),
    .C(net4898),
    .A(net2982),
    .Y(_03418_));
 sg13g2_o21ai_1 _19650_ (.B1(_03418_),
    .Y(_01351_),
    .A1(_04488_),
    .A2(net4869));
 sg13g2_nand3_1 _19651_ (.B(net5279),
    .C(net4869),
    .A(net1832),
    .Y(_03419_));
 sg13g2_o21ai_1 _19652_ (.B1(_03419_),
    .Y(_01352_),
    .A1(_04489_),
    .A2(net4868));
 sg13g2_nand3_1 _19653_ (.B(net5255),
    .C(net4823),
    .A(net2530),
    .Y(_03420_));
 sg13g2_o21ai_1 _19654_ (.B1(_03420_),
    .Y(_01353_),
    .A1(_04490_),
    .A2(net4824));
 sg13g2_nand3_1 _19655_ (.B(net5255),
    .C(net4822),
    .A(net2917),
    .Y(_03421_));
 sg13g2_o21ai_1 _19656_ (.B1(_03421_),
    .Y(_01354_),
    .A1(_04491_),
    .A2(net4822));
 sg13g2_nand3_1 _19657_ (.B(net5252),
    .C(net4820),
    .A(net1964),
    .Y(_03422_));
 sg13g2_o21ai_1 _19658_ (.B1(_03422_),
    .Y(_01355_),
    .A1(_04492_),
    .A2(net4847));
 sg13g2_nand3_1 _19659_ (.B(net5269),
    .C(net4847),
    .A(net1506),
    .Y(_03423_));
 sg13g2_o21ai_1 _19660_ (.B1(_03423_),
    .Y(_01356_),
    .A1(_04493_),
    .A2(net4848));
 sg13g2_nand3_1 _19661_ (.B(net5271),
    .C(net4848),
    .A(net1225),
    .Y(_03424_));
 sg13g2_o21ai_1 _19662_ (.B1(_03424_),
    .Y(_01357_),
    .A1(_04494_),
    .A2(net4834));
 sg13g2_nand3_1 _19663_ (.B(net5262),
    .C(net4835),
    .A(net1461),
    .Y(_03425_));
 sg13g2_o21ai_1 _19664_ (.B1(_03425_),
    .Y(_01358_),
    .A1(_04495_),
    .A2(net4835));
 sg13g2_nand3_1 _19665_ (.B(net5261),
    .C(net4833),
    .A(net3157),
    .Y(_03426_));
 sg13g2_o21ai_1 _19666_ (.B1(_03426_),
    .Y(_01359_),
    .A1(_04496_),
    .A2(net4833));
 sg13g2_nand3_1 _19667_ (.B(net5261),
    .C(net4833),
    .A(net2267),
    .Y(_03427_));
 sg13g2_o21ai_1 _19668_ (.B1(_03427_),
    .Y(_01360_),
    .A1(_04497_),
    .A2(net4806));
 sg13g2_nand3_1 _19669_ (.B(net5246),
    .C(net4806),
    .A(net2240),
    .Y(_03428_));
 sg13g2_o21ai_1 _19670_ (.B1(_03428_),
    .Y(_01361_),
    .A1(_04498_),
    .A2(net4805));
 sg13g2_nand3_1 _19671_ (.B(net5245),
    .C(net4803),
    .A(net2708),
    .Y(_03429_));
 sg13g2_o21ai_1 _19672_ (.B1(_03429_),
    .Y(_01362_),
    .A1(_04499_),
    .A2(net4796));
 sg13g2_nand3_1 _19673_ (.B(net5239),
    .C(net4792),
    .A(net2014),
    .Y(_03430_));
 sg13g2_o21ai_1 _19674_ (.B1(_03430_),
    .Y(_01363_),
    .A1(_04500_),
    .A2(net4796));
 sg13g2_nand3_1 _19675_ (.B(net5239),
    .C(net4751),
    .A(net2505),
    .Y(_03431_));
 sg13g2_o21ai_1 _19676_ (.B1(_03431_),
    .Y(_01364_),
    .A1(_04501_),
    .A2(net4751));
 sg13g2_nand3_1 _19677_ (.B(net5221),
    .C(net4753),
    .A(net1549),
    .Y(_03432_));
 sg13g2_o21ai_1 _19678_ (.B1(_03432_),
    .Y(_01365_),
    .A1(_04502_),
    .A2(net4757));
 sg13g2_nand3_1 _19679_ (.B(net5238),
    .C(net4757),
    .A(net1681),
    .Y(_03433_));
 sg13g2_o21ai_1 _19680_ (.B1(_03433_),
    .Y(_01366_),
    .A1(_04503_),
    .A2(net4757));
 sg13g2_nand3_1 _19681_ (.B(net5226),
    .C(net4758),
    .A(net2070),
    .Y(_03434_));
 sg13g2_o21ai_1 _19682_ (.B1(_03434_),
    .Y(_01367_),
    .A1(_04504_),
    .A2(net4758));
 sg13g2_nand3_1 _19683_ (.B(net5226),
    .C(net4759),
    .A(net2287),
    .Y(_03435_));
 sg13g2_o21ai_1 _19684_ (.B1(_03435_),
    .Y(_01368_),
    .A1(_04505_),
    .A2(net4759));
 sg13g2_nand3_1 _19685_ (.B(net5226),
    .C(net4759),
    .A(net2242),
    .Y(_03436_));
 sg13g2_o21ai_1 _19686_ (.B1(_03436_),
    .Y(_01369_),
    .A1(_04506_),
    .A2(net4759));
 sg13g2_nand3_1 _19687_ (.B(net5232),
    .C(net4768),
    .A(net1217),
    .Y(_03437_));
 sg13g2_o21ai_1 _19688_ (.B1(_03437_),
    .Y(_01370_),
    .A1(_04507_),
    .A2(net4768));
 sg13g2_nand3_1 _19689_ (.B(net5232),
    .C(net4768),
    .A(net2868),
    .Y(_03438_));
 sg13g2_o21ai_1 _19690_ (.B1(_03438_),
    .Y(_01371_),
    .A1(_04508_),
    .A2(net4769));
 sg13g2_nand3_1 _19691_ (.B(net5227),
    .C(net4774),
    .A(net1152),
    .Y(_03439_));
 sg13g2_o21ai_1 _19692_ (.B1(_03439_),
    .Y(_01372_),
    .A1(_04509_),
    .A2(net4775));
 sg13g2_nand3_1 _19693_ (.B(net5229),
    .C(net4775),
    .A(net1927),
    .Y(_03440_));
 sg13g2_o21ai_1 _19694_ (.B1(_03440_),
    .Y(_01373_),
    .A1(_04510_),
    .A2(net4775));
 sg13g2_nand3_1 _19695_ (.B(net5233),
    .C(net4780),
    .A(net3273),
    .Y(_03441_));
 sg13g2_o21ai_1 _19696_ (.B1(_03441_),
    .Y(_01374_),
    .A1(_04511_),
    .A2(net4781));
 sg13g2_nand3_1 _19697_ (.B(net5235),
    .C(net4784),
    .A(net2786),
    .Y(_03442_));
 sg13g2_o21ai_1 _19698_ (.B1(_03442_),
    .Y(_01375_),
    .A1(_04512_),
    .A2(net4784));
 sg13g2_nand3_1 _19699_ (.B(net5236),
    .C(net4786),
    .A(net1367),
    .Y(_03443_));
 sg13g2_o21ai_1 _19700_ (.B1(_03443_),
    .Y(_01376_),
    .A1(_04513_),
    .A2(net4786));
 sg13g2_nand3_1 _19701_ (.B(net5285),
    .C(net4786),
    .A(net2910),
    .Y(_03444_));
 sg13g2_o21ai_1 _19702_ (.B1(_03444_),
    .Y(_01377_),
    .A1(_04514_),
    .A2(net4879));
 sg13g2_nand3_1 _19703_ (.B(net5283),
    .C(net4879),
    .A(net1160),
    .Y(_03445_));
 sg13g2_o21ai_1 _19704_ (.B1(_03445_),
    .Y(_01378_),
    .A1(_04515_),
    .A2(net4886));
 sg13g2_nand3_1 _19705_ (.B(net5287),
    .C(net4886),
    .A(net2914),
    .Y(_03446_));
 sg13g2_o21ai_1 _19706_ (.B1(_03446_),
    .Y(_01379_),
    .A1(_04516_),
    .A2(net4885));
 sg13g2_nand3_1 _19707_ (.B(net5288),
    .C(net4887),
    .A(net1221),
    .Y(_03447_));
 sg13g2_o21ai_1 _19708_ (.B1(_03447_),
    .Y(_01380_),
    .A1(_04517_),
    .A2(net4887));
 sg13g2_nand3_1 _19709_ (.B(net5280),
    .C(net4873),
    .A(net3028),
    .Y(_03448_));
 sg13g2_o21ai_1 _19710_ (.B1(_03448_),
    .Y(_01381_),
    .A1(_04518_),
    .A2(net4872));
 sg13g2_nand3_1 _19711_ (.B(net5280),
    .C(net4873),
    .A(net2118),
    .Y(_03449_));
 sg13g2_o21ai_1 _19712_ (.B1(_03449_),
    .Y(_01382_),
    .A1(_04519_),
    .A2(net4872));
 sg13g2_nand3_1 _19713_ (.B(net5294),
    .C(net4898),
    .A(net1144),
    .Y(_03450_));
 sg13g2_o21ai_1 _19714_ (.B1(_03450_),
    .Y(_01383_),
    .A1(_04520_),
    .A2(net4898));
 sg13g2_nand3_1 _19715_ (.B(net5293),
    .C(net4897),
    .A(net2248),
    .Y(_03451_));
 sg13g2_o21ai_1 _19716_ (.B1(_03451_),
    .Y(_01384_),
    .A1(_04521_),
    .A2(net4895));
 sg13g2_nand3_1 _19717_ (.B(net5293),
    .C(net4895),
    .A(net3271),
    .Y(_03452_));
 sg13g2_o21ai_1 _19718_ (.B1(_03452_),
    .Y(_01385_),
    .A1(_04522_),
    .A2(net4895));
 sg13g2_nand3_1 _19719_ (.B(net5293),
    .C(net4895),
    .A(net1162),
    .Y(_03453_));
 sg13g2_o21ai_1 _19720_ (.B1(_03453_),
    .Y(_01386_),
    .A1(_04523_),
    .A2(net4851));
 sg13g2_nand3_1 _19721_ (.B(net5271),
    .C(net4852),
    .A(net2261),
    .Y(_03454_));
 sg13g2_o21ai_1 _19722_ (.B1(_03454_),
    .Y(_01387_),
    .A1(_04524_),
    .A2(net4853));
 sg13g2_nand3_1 _19723_ (.B(net5272),
    .C(net4855),
    .A(net2317),
    .Y(_03455_));
 sg13g2_o21ai_1 _19724_ (.B1(_03455_),
    .Y(_01388_),
    .A1(_04525_),
    .A2(net4854));
 sg13g2_nand3_1 _19725_ (.B(net5273),
    .C(net4854),
    .A(net2503),
    .Y(_03456_));
 sg13g2_o21ai_1 _19726_ (.B1(_03456_),
    .Y(_01389_),
    .A1(_04526_),
    .A2(net4854));
 sg13g2_nand3_1 _19727_ (.B(net5265),
    .C(net4842),
    .A(net2544),
    .Y(_03457_));
 sg13g2_o21ai_1 _19728_ (.B1(_03457_),
    .Y(_01390_),
    .A1(_04527_),
    .A2(net4842));
 sg13g2_nand3_1 _19729_ (.B(net5265),
    .C(net4842),
    .A(net3254),
    .Y(_03458_));
 sg13g2_o21ai_1 _19730_ (.B1(_03458_),
    .Y(_01391_),
    .A1(_04528_),
    .A2(net4832));
 sg13g2_nand3_1 _19731_ (.B(net5246),
    .C(net4805),
    .A(net2396),
    .Y(_03459_));
 sg13g2_o21ai_1 _19732_ (.B1(_03459_),
    .Y(_01392_),
    .A1(_04529_),
    .A2(net4805));
 sg13g2_nand3_1 _19733_ (.B(net5253),
    .C(net4819),
    .A(net2957),
    .Y(_03460_));
 sg13g2_o21ai_1 _19734_ (.B1(_03460_),
    .Y(_01393_),
    .A1(_04530_),
    .A2(net4818));
 sg13g2_nand3_1 _19735_ (.B(net5252),
    .C(net4818),
    .A(net1541),
    .Y(_03461_));
 sg13g2_o21ai_1 _19736_ (.B1(_03461_),
    .Y(_01394_),
    .A1(_04531_),
    .A2(net4818));
 sg13g2_nand3_1 _19737_ (.B(net5248),
    .C(net4810),
    .A(net1866),
    .Y(_03462_));
 sg13g2_o21ai_1 _19738_ (.B1(_03462_),
    .Y(_01395_),
    .A1(_04532_),
    .A2(net4810));
 sg13g2_nand3_1 _19739_ (.B(net5248),
    .C(net4810),
    .A(net1921),
    .Y(_03463_));
 sg13g2_o21ai_1 _19740_ (.B1(_03463_),
    .Y(_01396_),
    .A1(_04533_),
    .A2(net4810));
 sg13g2_nand3_1 _19741_ (.B(net5251),
    .C(net4810),
    .A(net2422),
    .Y(_03464_));
 sg13g2_o21ai_1 _19742_ (.B1(_03464_),
    .Y(_01397_),
    .A1(_04534_),
    .A2(net4809));
 sg13g2_nand3_1 _19743_ (.B(net5247),
    .C(net4809),
    .A(net2603),
    .Y(_03465_));
 sg13g2_o21ai_1 _19744_ (.B1(_03465_),
    .Y(_01398_),
    .A1(_04535_),
    .A2(net4761));
 sg13g2_nand3_1 _19745_ (.B(net5223),
    .C(net4761),
    .A(net1189),
    .Y(_03466_));
 sg13g2_o21ai_1 _19746_ (.B1(_03466_),
    .Y(_01399_),
    .A1(_04536_),
    .A2(net4760));
 sg13g2_nand3_1 _19747_ (.B(net5224),
    .C(net4763),
    .A(net2686),
    .Y(_03467_));
 sg13g2_o21ai_1 _19748_ (.B1(_03467_),
    .Y(_01400_),
    .A1(_04537_),
    .A2(net4764));
 sg13g2_nand3_1 _19749_ (.B(net5226),
    .C(net4759),
    .A(net2454),
    .Y(_03468_));
 sg13g2_o21ai_1 _19750_ (.B1(_03468_),
    .Y(_01401_),
    .A1(_04538_),
    .A2(net4768));
 sg13g2_nand3_1 _19751_ (.B(net5232),
    .C(net4768),
    .A(net1236),
    .Y(_03469_));
 sg13g2_o21ai_1 _19752_ (.B1(_03469_),
    .Y(_01402_),
    .A1(_04539_),
    .A2(net4769));
 sg13g2_nand3_1 _19753_ (.B(net5232),
    .C(net4768),
    .A(net1960),
    .Y(_03470_));
 sg13g2_o21ai_1 _19754_ (.B1(_03470_),
    .Y(_01403_),
    .A1(_04540_),
    .A2(net4769));
 sg13g2_nand3_1 _19755_ (.B(net5232),
    .C(net4770),
    .A(net2408),
    .Y(_03471_));
 sg13g2_o21ai_1 _19756_ (.B1(_03471_),
    .Y(_01404_),
    .A1(_04541_),
    .A2(net4770));
 sg13g2_nand3_1 _19757_ (.B(net5229),
    .C(net4776),
    .A(net2651),
    .Y(_03472_));
 sg13g2_o21ai_1 _19758_ (.B1(_03472_),
    .Y(_01405_),
    .A1(_04542_),
    .A2(net4775));
 sg13g2_nand3_1 _19759_ (.B(net5233),
    .C(net4780),
    .A(net2410),
    .Y(_03473_));
 sg13g2_o21ai_1 _19760_ (.B1(_03473_),
    .Y(_01406_),
    .A1(_04543_),
    .A2(net4780));
 sg13g2_nand3_1 _19761_ (.B(net5233),
    .C(net4781),
    .A(net3128),
    .Y(_03474_));
 sg13g2_o21ai_1 _19762_ (.B1(_03474_),
    .Y(_01407_),
    .A1(_04544_),
    .A2(net4784));
 sg13g2_nand3_1 _19763_ (.B(net5235),
    .C(net4784),
    .A(net1823),
    .Y(_03475_));
 sg13g2_o21ai_1 _19764_ (.B1(_03475_),
    .Y(_01408_),
    .A1(_04545_),
    .A2(net4785));
 sg13g2_nand3_1 _19765_ (.B(net5235),
    .C(net4786),
    .A(net1579),
    .Y(_03476_));
 sg13g2_o21ai_1 _19766_ (.B1(_03476_),
    .Y(_01409_),
    .A1(_04546_),
    .A2(net4881));
 sg13g2_nand3_1 _19767_ (.B(net5289),
    .C(net4890),
    .A(net2831),
    .Y(_03477_));
 sg13g2_o21ai_1 _19768_ (.B1(_03477_),
    .Y(_01410_),
    .A1(_04547_),
    .A2(net4890));
 sg13g2_nand3_1 _19769_ (.B(net5289),
    .C(net4889),
    .A(net1493),
    .Y(_03478_));
 sg13g2_o21ai_1 _19770_ (.B1(_03478_),
    .Y(_01411_),
    .A1(_04548_),
    .A2(net4889));
 sg13g2_nand3_1 _19771_ (.B(net5288),
    .C(net4888),
    .A(net2902),
    .Y(_03479_));
 sg13g2_o21ai_1 _19772_ (.B1(_03479_),
    .Y(_01412_),
    .A1(_04549_),
    .A2(net4887));
 sg13g2_nand3_1 _19773_ (.B(net5287),
    .C(net4887),
    .A(net3090),
    .Y(_03480_));
 sg13g2_o21ai_1 _19774_ (.B1(_03480_),
    .Y(_01413_),
    .A1(_04550_),
    .A2(net4872));
 sg13g2_nand3_1 _19775_ (.B(net5280),
    .C(net4872),
    .A(net1569),
    .Y(_03481_));
 sg13g2_o21ai_1 _19776_ (.B1(_03481_),
    .Y(_01414_),
    .A1(_04551_),
    .A2(net4872));
 sg13g2_nand3_1 _19777_ (.B(net5281),
    .C(net4872),
    .A(net2405),
    .Y(_03482_));
 sg13g2_o21ai_1 _19778_ (.B1(_03482_),
    .Y(_01415_),
    .A1(_04552_),
    .A2(net4868));
 sg13g2_nand3_1 _19779_ (.B(net5279),
    .C(net4868),
    .A(net2429),
    .Y(_03483_));
 sg13g2_o21ai_1 _19780_ (.B1(_03483_),
    .Y(_01416_),
    .A1(_04553_),
    .A2(net4868));
 sg13g2_nand3_1 _19781_ (.B(net5255),
    .C(net4823),
    .A(net2233),
    .Y(_03484_));
 sg13g2_o21ai_1 _19782_ (.B1(_03484_),
    .Y(_01417_),
    .A1(_04554_),
    .A2(net4823));
 sg13g2_nand3_1 _19783_ (.B(net5254),
    .C(net4822),
    .A(net2239),
    .Y(_03485_));
 sg13g2_o21ai_1 _19784_ (.B1(_03485_),
    .Y(_01418_),
    .A1(_04555_),
    .A2(net4850));
 sg13g2_nand3_1 _19785_ (.B(net5270),
    .C(net4850),
    .A(net1156),
    .Y(_03486_));
 sg13g2_o21ai_1 _19786_ (.B1(_03486_),
    .Y(_01419_),
    .A1(_04556_),
    .A2(net4852));
 sg13g2_nand3_1 _19787_ (.B(net5269),
    .C(net4848),
    .A(net2711),
    .Y(_03487_));
 sg13g2_o21ai_1 _19788_ (.B1(_03487_),
    .Y(_01420_),
    .A1(_04557_),
    .A2(net4854));
 sg13g2_nand3_1 _19789_ (.B(net5263),
    .C(net4837),
    .A(net3107),
    .Y(_03488_));
 sg13g2_o21ai_1 _19790_ (.B1(_03488_),
    .Y(_01421_),
    .A1(_04558_),
    .A2(net4837));
 sg13g2_nand3_1 _19791_ (.B(net5263),
    .C(net4837),
    .A(net2103),
    .Y(_03489_));
 sg13g2_o21ai_1 _19792_ (.B1(_03489_),
    .Y(_01422_),
    .A1(_04559_),
    .A2(net4837));
 sg13g2_nand3_1 _19793_ (.B(net5258),
    .C(net4827),
    .A(net2590),
    .Y(_03490_));
 sg13g2_o21ai_1 _19794_ (.B1(_03490_),
    .Y(_01423_),
    .A1(_04560_),
    .A2(net4827));
 sg13g2_nand3_1 _19795_ (.B(net5258),
    .C(net4827),
    .A(net2465),
    .Y(_03491_));
 sg13g2_o21ai_1 _19796_ (.B1(_03491_),
    .Y(_01424_),
    .A1(_04561_),
    .A2(net4801));
 sg13g2_nand3_1 _19797_ (.B(net5244),
    .C(net4802),
    .A(net3092),
    .Y(_03492_));
 sg13g2_o21ai_1 _19798_ (.B1(_03492_),
    .Y(_01425_),
    .A1(_04562_),
    .A2(net4800));
 sg13g2_nand3_1 _19799_ (.B(net5244),
    .C(net4800),
    .A(net2054),
    .Y(_03493_));
 sg13g2_o21ai_1 _19800_ (.B1(_03493_),
    .Y(_01426_),
    .A1(_04563_),
    .A2(net4800));
 sg13g2_nand3_1 _19801_ (.B(net5242),
    .C(net4796),
    .A(net2516),
    .Y(_03494_));
 sg13g2_o21ai_1 _19802_ (.B1(_03494_),
    .Y(_01427_),
    .A1(_04564_),
    .A2(net4796));
 sg13g2_nand3_1 _19803_ (.B(net5241),
    .C(net4797),
    .A(net2219),
    .Y(_03495_));
 sg13g2_o21ai_1 _19804_ (.B1(_03495_),
    .Y(_01428_),
    .A1(_04565_),
    .A2(net4794));
 sg13g2_nand3_1 _19805_ (.B(net5247),
    .C(net4809),
    .A(net2438),
    .Y(_03496_));
 sg13g2_o21ai_1 _19806_ (.B1(_03496_),
    .Y(_01429_),
    .A1(_04566_),
    .A2(net4809));
 sg13g2_nand3_1 _19807_ (.B(net5247),
    .C(net4809),
    .A(net1954),
    .Y(_03497_));
 sg13g2_o21ai_1 _19808_ (.B1(_03497_),
    .Y(_01430_),
    .A1(_04567_),
    .A2(net4809));
 sg13g2_nand3_1 _19809_ (.B(net5247),
    .C(net4808),
    .A(net2178),
    .Y(_03498_));
 sg13g2_o21ai_1 _19810_ (.B1(_03498_),
    .Y(_01431_),
    .A1(_04568_),
    .A2(net4808));
 sg13g2_nand3_1 _19811_ (.B(net5249),
    .C(net4813),
    .A(net2427),
    .Y(_03499_));
 sg13g2_o21ai_1 _19812_ (.B1(_03499_),
    .Y(_01432_),
    .A1(_04569_),
    .A2(net4813));
 sg13g2_nand3_1 _19813_ (.B(net5249),
    .C(net4814),
    .A(net2448),
    .Y(_03500_));
 sg13g2_o21ai_1 _19814_ (.B1(_03500_),
    .Y(_01433_),
    .A1(_04570_),
    .A2(net4814));
 sg13g2_nand3_1 _19815_ (.B(net5275),
    .C(net4859),
    .A(net1202),
    .Y(_03501_));
 sg13g2_o21ai_1 _19816_ (.B1(_03501_),
    .Y(_01434_),
    .A1(_04571_),
    .A2(net4859));
 sg13g2_nand3_1 _19817_ (.B(net5275),
    .C(net4860),
    .A(net2083),
    .Y(_03502_));
 sg13g2_o21ai_1 _19818_ (.B1(_03502_),
    .Y(_01435_),
    .A1(_04572_),
    .A2(net4860));
 sg13g2_nand3_1 _19819_ (.B(net5275),
    .C(net4860),
    .A(net3211),
    .Y(_03503_));
 sg13g2_o21ai_1 _19820_ (.B1(_03503_),
    .Y(_01436_),
    .A1(_04573_),
    .A2(net4863));
 sg13g2_nand3_1 _19821_ (.B(net5230),
    .C(net4777),
    .A(net1133),
    .Y(_03504_));
 sg13g2_o21ai_1 _19822_ (.B1(_03504_),
    .Y(_01437_),
    .A1(_04574_),
    .A2(net4777));
 sg13g2_nand3_1 _19823_ (.B(net5230),
    .C(net4778),
    .A(\TRNG.Word_Out[193] ),
    .Y(_03505_));
 sg13g2_o21ai_1 _19824_ (.B1(_03505_),
    .Y(_01438_),
    .A1(_04575_),
    .A2(net4782));
 sg13g2_nand3_1 _19825_ (.B(net5234),
    .C(net4783),
    .A(net2875),
    .Y(_03506_));
 sg13g2_o21ai_1 _19826_ (.B1(_03506_),
    .Y(_01439_),
    .A1(_04576_),
    .A2(net4786));
 sg13g2_nand3_1 _19827_ (.B(net5236),
    .C(net4786),
    .A(net1962),
    .Y(_03507_));
 sg13g2_o21ai_1 _19828_ (.B1(_03507_),
    .Y(_01440_),
    .A1(_04577_),
    .A2(net4786));
 sg13g2_nand3_1 _19829_ (.B(net5285),
    .C(net4880),
    .A(net2417),
    .Y(_03508_));
 sg13g2_o21ai_1 _19830_ (.B1(_03508_),
    .Y(_01441_),
    .A1(_04578_),
    .A2(net4882));
 sg13g2_nand3_1 _19831_ (.B(net5289),
    .C(net4889),
    .A(net1573),
    .Y(_03509_));
 sg13g2_o21ai_1 _19832_ (.B1(_03509_),
    .Y(_01442_),
    .A1(_04579_),
    .A2(net4889));
 sg13g2_nand3_1 _19833_ (.B(net5290),
    .C(net4891),
    .A(net1749),
    .Y(_03510_));
 sg13g2_o21ai_1 _19834_ (.B1(_03510_),
    .Y(_01443_),
    .A1(_04580_),
    .A2(net4888));
 sg13g2_nand3_1 _19835_ (.B(net5287),
    .C(net4888),
    .A(net2252),
    .Y(_03511_));
 sg13g2_o21ai_1 _19836_ (.B1(_03511_),
    .Y(_01444_),
    .A1(_04581_),
    .A2(net4905));
 sg13g2_nand3_1 _19837_ (.B(net5297),
    .C(net4904),
    .A(net1280),
    .Y(_03512_));
 sg13g2_o21ai_1 _19838_ (.B1(_03512_),
    .Y(_01445_),
    .A1(_04582_),
    .A2(net4905));
 sg13g2_nand3_1 _19839_ (.B(net5297),
    .C(net4904),
    .A(net2984),
    .Y(_03513_));
 sg13g2_o21ai_1 _19840_ (.B1(_03513_),
    .Y(_01446_),
    .A1(_04583_),
    .A2(net4898));
 sg13g2_nand3_1 _19841_ (.B(net5278),
    .C(net4866),
    .A(net3171),
    .Y(_03514_));
 sg13g2_o21ai_1 _19842_ (.B1(_03514_),
    .Y(_01447_),
    .A1(_04584_),
    .A2(net4867));
 sg13g2_nand3_1 _19843_ (.B(net5278),
    .C(net4866),
    .A(net3044),
    .Y(_03515_));
 sg13g2_o21ai_1 _19844_ (.B1(_03515_),
    .Y(_01448_),
    .A1(_04585_),
    .A2(net4821));
 sg13g2_nand3_1 _19845_ (.B(net5254),
    .C(net4821),
    .A(net2648),
    .Y(_03516_));
 sg13g2_o21ai_1 _19846_ (.B1(_03516_),
    .Y(_01449_),
    .A1(_04586_),
    .A2(net4821));
 sg13g2_nand3_1 _19847_ (.B(net5252),
    .C(net4818),
    .A(net2105),
    .Y(_03517_));
 sg13g2_o21ai_1 _19848_ (.B1(_03517_),
    .Y(_01450_),
    .A1(_04587_),
    .A2(net4820));
 sg13g2_nand3_1 _19849_ (.B(net5252),
    .C(net4819),
    .A(net2005),
    .Y(_03518_));
 sg13g2_o21ai_1 _19850_ (.B1(_03518_),
    .Y(_01451_),
    .A1(_04588_),
    .A2(net4846));
 sg13g2_nand3_1 _19851_ (.B(net5261),
    .C(net4832),
    .A(net2238),
    .Y(_03519_));
 sg13g2_o21ai_1 _19852_ (.B1(_03519_),
    .Y(_01452_),
    .A1(_04589_),
    .A2(net4834));
 sg13g2_nand3_1 _19853_ (.B(net5265),
    .C(net4841),
    .A(net1891),
    .Y(_03520_));
 sg13g2_o21ai_1 _19854_ (.B1(_03520_),
    .Y(_01453_),
    .A1(_04590_),
    .A2(net4841));
 sg13g2_nand3_1 _19855_ (.B(net5262),
    .C(net4834),
    .A(net1973),
    .Y(_03521_));
 sg13g2_o21ai_1 _19856_ (.B1(_03521_),
    .Y(_01454_),
    .A1(_04591_),
    .A2(net4834));
 sg13g2_nand3_1 _19857_ (.B(net5261),
    .C(net4832),
    .A(net2114),
    .Y(_03522_));
 sg13g2_o21ai_1 _19858_ (.B1(_03522_),
    .Y(_01455_),
    .A1(_04592_),
    .A2(net4832));
 sg13g2_nand3_1 _19859_ (.B(net5261),
    .C(net4832),
    .A(net3296),
    .Y(_03523_));
 sg13g2_o21ai_1 _19860_ (.B1(_03523_),
    .Y(_01456_),
    .A1(_04593_),
    .A2(net4805));
 sg13g2_nand3_1 _19861_ (.B(net5253),
    .C(net4819),
    .A(net2564),
    .Y(_03524_));
 sg13g2_o21ai_1 _19862_ (.B1(_03524_),
    .Y(_01457_),
    .A1(_04594_),
    .A2(net4818));
 sg13g2_nand3_1 _19863_ (.B(net5252),
    .C(net4820),
    .A(net2446),
    .Y(_03525_));
 sg13g2_o21ai_1 _19864_ (.B1(_03525_),
    .Y(_01458_),
    .A1(_04595_),
    .A2(net4820));
 sg13g2_nand3_1 _19865_ (.B(net5248),
    .C(net4810),
    .A(net2540),
    .Y(_03526_));
 sg13g2_o21ai_1 _19866_ (.B1(_03526_),
    .Y(_01459_),
    .A1(_04596_),
    .A2(net4810));
 sg13g2_nand3_1 _19867_ (.B(net5248),
    .C(net4811),
    .A(net1904),
    .Y(_03527_));
 sg13g2_o21ai_1 _19868_ (.B1(_03527_),
    .Y(_01460_),
    .A1(_04597_),
    .A2(net4811));
 sg13g2_nand3_1 _19869_ (.B(net5248),
    .C(net4811),
    .A(net2225),
    .Y(_03528_));
 sg13g2_o21ai_1 _19870_ (.B1(_03528_),
    .Y(_01461_),
    .A1(_04598_),
    .A2(net4808));
 sg13g2_nand3_1 _19871_ (.B(net5247),
    .C(net4808),
    .A(net2017),
    .Y(_03529_));
 sg13g2_o21ai_1 _19872_ (.B1(_03529_),
    .Y(_01462_),
    .A1(_04599_),
    .A2(net4808));
 sg13g2_nand3_1 _19873_ (.B(net5247),
    .C(net4808),
    .A(net1994),
    .Y(_03530_));
 sg13g2_o21ai_1 _19874_ (.B1(_03530_),
    .Y(_01463_),
    .A1(_04600_),
    .A2(net4813));
 sg13g2_nand3_1 _19875_ (.B(net5249),
    .C(net4813),
    .A(net2407),
    .Y(_03531_));
 sg13g2_o21ai_1 _19876_ (.B1(_03531_),
    .Y(_01464_),
    .A1(_04601_),
    .A2(net4813));
 sg13g2_nand3_1 _19877_ (.B(net5249),
    .C(net4814),
    .A(net2366),
    .Y(_03532_));
 sg13g2_o21ai_1 _19878_ (.B1(_03532_),
    .Y(_01465_),
    .A1(_04602_),
    .A2(net4814));
 sg13g2_nand3_1 _19879_ (.B(net5250),
    .C(net4816),
    .A(net2445),
    .Y(_03533_));
 sg13g2_o21ai_1 _19880_ (.B1(_03533_),
    .Y(_01466_),
    .A1(_04603_),
    .A2(net4861));
 sg13g2_nand3_1 _19881_ (.B(net5276),
    .C(net4861),
    .A(net1947),
    .Y(_03534_));
 sg13g2_o21ai_1 _19882_ (.B1(_03534_),
    .Y(_01467_),
    .A1(_04604_),
    .A2(net4861));
 sg13g2_nand3_1 _19883_ (.B(net5276),
    .C(net4862),
    .A(net2769),
    .Y(_03535_));
 sg13g2_o21ai_1 _19884_ (.B1(_03535_),
    .Y(_01468_),
    .A1(_04605_),
    .A2(net4864));
 sg13g2_nand3_1 _19885_ (.B(net5230),
    .C(net4778),
    .A(net1158),
    .Y(_03536_));
 sg13g2_o21ai_1 _19886_ (.B1(_03536_),
    .Y(_01469_),
    .A1(_04606_),
    .A2(net4778));
 sg13g2_nand3_1 _19887_ (.B(net5234),
    .C(net4782),
    .A(\TRNG.Word_Out[225] ),
    .Y(_03537_));
 sg13g2_o21ai_1 _19888_ (.B1(_03537_),
    .Y(_01470_),
    .A1(_04607_),
    .A2(net4782));
 sg13g2_nand3_1 _19889_ (.B(net5234),
    .C(net4783),
    .A(net3229),
    .Y(_03538_));
 sg13g2_o21ai_1 _19890_ (.B1(_03538_),
    .Y(_01471_),
    .A1(_04608_),
    .A2(net4787));
 sg13g2_nand3_1 _19891_ (.B(net5285),
    .C(net4881),
    .A(net1956),
    .Y(_03539_));
 sg13g2_o21ai_1 _19892_ (.B1(_03539_),
    .Y(_01472_),
    .A1(_04609_),
    .A2(net4881));
 sg13g2_nand3_1 _19893_ (.B(net5286),
    .C(net4882),
    .A(net1208),
    .Y(_03540_));
 sg13g2_o21ai_1 _19894_ (.B1(_03540_),
    .Y(_01473_),
    .A1(_04610_),
    .A2(net4883));
 sg13g2_nand3_1 _19895_ (.B(net5285),
    .C(net4882),
    .A(net1741),
    .Y(_03541_));
 sg13g2_o21ai_1 _19896_ (.B1(_03541_),
    .Y(_01474_),
    .A1(_04611_),
    .A2(net4882));
 sg13g2_nand3_1 _19897_ (.B(net5290),
    .C(net4891),
    .A(net2283),
    .Y(_03542_));
 sg13g2_o21ai_1 _19898_ (.B1(_03542_),
    .Y(_01475_),
    .A1(_04612_),
    .A2(net4908));
 sg13g2_nand3_1 _19899_ (.B(net5298),
    .C(net4908),
    .A(net1836),
    .Y(_03543_));
 sg13g2_o21ai_1 _19900_ (.B1(_03543_),
    .Y(_01476_),
    .A1(_04613_),
    .A2(net4908));
 sg13g2_nand3_1 _19901_ (.B(net5299),
    .C(net4910),
    .A(net2204),
    .Y(_03544_));
 sg13g2_o21ai_1 _19902_ (.B1(_03544_),
    .Y(_01477_),
    .A1(_04614_),
    .A2(net4910));
 sg13g2_nand3_1 _19903_ (.B(net5299),
    .C(net4910),
    .A(net3311),
    .Y(_03545_));
 sg13g2_o21ai_1 _19904_ (.B1(_03545_),
    .Y(_01478_),
    .A1(_04615_),
    .A2(net4906));
 sg13g2_nand3_1 _19905_ (.B(net5295),
    .C(net4900),
    .A(net2274),
    .Y(_03546_));
 sg13g2_o21ai_1 _19906_ (.B1(_03546_),
    .Y(_01479_),
    .A1(_04616_),
    .A2(net4900));
 sg13g2_nand3_1 _19907_ (.B(net5294),
    .C(net4900),
    .A(net2383),
    .Y(_03547_));
 sg13g2_o21ai_1 _19908_ (.B1(_03547_),
    .Y(_01480_),
    .A1(_04617_),
    .A2(net4896));
 sg13g2_nand3_1 _19909_ (.B(net5295),
    .C(net4897),
    .A(net2659),
    .Y(_03548_));
 sg13g2_o21ai_1 _19910_ (.B1(_03548_),
    .Y(_01481_),
    .A1(_04618_),
    .A2(net4896));
 sg13g2_nand3_1 _19911_ (.B(net5295),
    .C(net4896),
    .A(net2243),
    .Y(_03549_));
 sg13g2_o21ai_1 _19912_ (.B1(_03549_),
    .Y(_01482_),
    .A1(_04619_),
    .A2(net4852));
 sg13g2_nand3_1 _19913_ (.B(net5270),
    .C(net4852),
    .A(net2094),
    .Y(_03550_));
 sg13g2_o21ai_1 _19914_ (.B1(_03550_),
    .Y(_01483_),
    .A1(_04620_),
    .A2(net4855));
 sg13g2_nand3_1 _19915_ (.B(net5265),
    .C(net4841),
    .A(net3220),
    .Y(_03551_));
 sg13g2_o21ai_1 _19916_ (.B1(_03551_),
    .Y(_01484_),
    .A1(_04621_),
    .A2(net4841));
 sg13g2_nand3_1 _19917_ (.B(net5264),
    .C(net4839),
    .A(net1428),
    .Y(_03552_));
 sg13g2_o21ai_1 _19918_ (.B1(_03552_),
    .Y(_01485_),
    .A1(_04622_),
    .A2(net4839));
 sg13g2_nand3_1 _19919_ (.B(net5263),
    .C(net4840),
    .A(net2339),
    .Y(_03553_));
 sg13g2_o21ai_1 _19920_ (.B1(_03553_),
    .Y(_01486_),
    .A1(_04623_),
    .A2(net4840));
 sg13g2_nand3_1 _19921_ (.B(net5264),
    .C(net4839),
    .A(net3203),
    .Y(_03554_));
 sg13g2_o21ai_1 _19922_ (.B1(_03554_),
    .Y(_01487_),
    .A1(_04624_),
    .A2(net4828));
 sg13g2_nand3_1 _19923_ (.B(net5258),
    .C(net4828),
    .A(net3127),
    .Y(_03555_));
 sg13g2_o21ai_1 _19924_ (.B1(_03555_),
    .Y(_01488_),
    .A1(_04625_),
    .A2(net4805));
 sg13g2_nand3_1 _19925_ (.B(net5245),
    .C(net4805),
    .A(net2488),
    .Y(_03556_));
 sg13g2_o21ai_1 _19926_ (.B1(_03556_),
    .Y(_01489_),
    .A1(_04626_),
    .A2(net4803));
 sg13g2_nand3_1 _19927_ (.B(net5245),
    .C(net4803),
    .A(net2425),
    .Y(_03557_));
 sg13g2_o21ai_1 _19928_ (.B1(_03557_),
    .Y(_01490_),
    .A1(_04627_),
    .A2(net4818));
 sg13g2_nand3_1 _19929_ (.B(net5248),
    .C(net4810),
    .A(net2485),
    .Y(_03558_));
 sg13g2_o21ai_1 _19930_ (.B1(_03558_),
    .Y(_01491_),
    .A1(_04628_),
    .A2(net4797));
 sg13g2_nand3_1 _19931_ (.B(net5242),
    .C(net4795),
    .A(net1560),
    .Y(_03559_));
 sg13g2_o21ai_1 _19932_ (.B1(_03559_),
    .Y(_01492_),
    .A1(_04629_),
    .A2(net4794));
 sg13g2_nand3_1 _19933_ (.B(net5241),
    .C(net4794),
    .A(net2583),
    .Y(_03560_));
 sg13g2_o21ai_1 _19934_ (.B1(_03560_),
    .Y(_01493_),
    .A1(_04630_),
    .A2(net4753));
 sg13g2_nand3_1 _19935_ (.B(net5220),
    .C(net4754),
    .A(net1348),
    .Y(_03561_));
 sg13g2_o21ai_1 _19936_ (.B1(_03561_),
    .Y(_01494_),
    .A1(_04631_),
    .A2(net4754));
 sg13g2_nand3_1 _19937_ (.B(net5225),
    .C(net4761),
    .A(net3290),
    .Y(_03562_));
 sg13g2_o21ai_1 _19938_ (.B1(_03562_),
    .Y(_01495_),
    .A1(_04632_),
    .A2(net4761));
 sg13g2_nand3_1 _19939_ (.B(net5247),
    .C(net4808),
    .A(net2431),
    .Y(_03563_));
 sg13g2_o21ai_1 _19940_ (.B1(_03563_),
    .Y(_01496_),
    .A1(_04633_),
    .A2(net4811));
 sg13g2_nand3_1 _19941_ (.B(net5250),
    .C(net4815),
    .A(net2605),
    .Y(_03564_));
 sg13g2_o21ai_1 _19942_ (.B1(_03564_),
    .Y(_01497_),
    .A1(_04634_),
    .A2(net4815));
 sg13g2_nand3_1 _19943_ (.B(net5250),
    .C(net4816),
    .A(net2254),
    .Y(_03565_));
 sg13g2_o21ai_1 _19944_ (.B1(_03565_),
    .Y(_01498_),
    .A1(_04635_),
    .A2(net4816));
 sg13g2_nand3_1 _19945_ (.B(net5276),
    .C(net4861),
    .A(net1195),
    .Y(_03566_));
 sg13g2_o21ai_1 _19946_ (.B1(_03566_),
    .Y(_01499_),
    .A1(_04636_),
    .A2(net4861));
 sg13g2_nand3_1 _19947_ (.B(net5276),
    .C(net4861),
    .A(net3046),
    .Y(_03567_));
 sg13g2_o21ai_1 _19948_ (.B1(_03567_),
    .Y(_01500_),
    .A1(_04637_),
    .A2(net4863));
 sg13g2_nand3_1 _19949_ (.B(net5277),
    .C(net4863),
    .A(net2206),
    .Y(_03568_));
 sg13g2_o21ai_1 _19950_ (.B1(_03568_),
    .Y(_01501_),
    .A1(_04638_),
    .A2(net4865));
 sg13g2_nand3_1 _19951_ (.B(net5282),
    .C(net4865),
    .A(net2398),
    .Y(_03569_));
 sg13g2_o21ai_1 _19952_ (.B1(_03569_),
    .Y(_01502_),
    .A1(_04639_),
    .A2(net4876));
 sg13g2_nand3_1 _19953_ (.B(net5284),
    .C(net4876),
    .A(net1851),
    .Y(_03570_));
 sg13g2_o21ai_1 _19954_ (.B1(_03570_),
    .Y(_01503_),
    .A1(_04640_),
    .A2(net4877));
 sg13g2_nand3_1 _19955_ (.B(net5284),
    .C(net4877),
    .A(net1920),
    .Y(_03571_));
 sg13g2_o21ai_1 _19956_ (.B1(_03571_),
    .Y(_01504_),
    .A1(_04641_),
    .A2(net4877));
 sg13g2_nand3_1 _19957_ (.B(net5284),
    .C(net4876),
    .A(net1759),
    .Y(_03572_));
 sg13g2_o21ai_1 _19958_ (.B1(_03572_),
    .Y(_01505_),
    .A1(_04642_),
    .A2(net4878));
 sg13g2_nand3_1 _19959_ (.B(net5283),
    .C(net4878),
    .A(net2546),
    .Y(_03573_));
 sg13g2_o21ai_1 _19960_ (.B1(_03573_),
    .Y(_01506_),
    .A1(_04643_),
    .A2(net4864));
 sg13g2_nand3_1 _19961_ (.B(net5277),
    .C(net4864),
    .A(net1788),
    .Y(_03574_));
 sg13g2_o21ai_1 _19962_ (.B1(_03574_),
    .Y(_01507_),
    .A1(_04644_),
    .A2(net4864));
 sg13g2_nand3_1 _19963_ (.B(net5280),
    .C(net4871),
    .A(net1371),
    .Y(_03575_));
 sg13g2_o21ai_1 _19964_ (.B1(_03575_),
    .Y(_01508_),
    .A1(_04645_),
    .A2(net4871));
 sg13g2_nand3_1 _19965_ (.B(net5280),
    .C(net4871),
    .A(net2188),
    .Y(_03576_));
 sg13g2_o21ai_1 _19966_ (.B1(_03576_),
    .Y(_01509_),
    .A1(_04646_),
    .A2(net4871));
 sg13g2_nand3_1 _19967_ (.B(net5280),
    .C(net4871),
    .A(net1253),
    .Y(_03577_));
 sg13g2_o21ai_1 _19968_ (.B1(_03577_),
    .Y(_01510_),
    .A1(_04647_),
    .A2(net4867));
 sg13g2_nand3_1 _19969_ (.B(net5278),
    .C(net4866),
    .A(net1623),
    .Y(_03578_));
 sg13g2_o21ai_1 _19970_ (.B1(_03578_),
    .Y(_01511_),
    .A1(_04648_),
    .A2(net4867));
 sg13g2_nand3_1 _19971_ (.B(net5278),
    .C(net4866),
    .A(net1732),
    .Y(_03579_));
 sg13g2_o21ai_1 _19972_ (.B1(_03579_),
    .Y(_01512_),
    .A1(_04649_),
    .A2(net4866));
 sg13g2_nand3_1 _19973_ (.B(net5255),
    .C(net4823),
    .A(net3050),
    .Y(_03580_));
 sg13g2_o21ai_1 _19974_ (.B1(_03580_),
    .Y(_01513_),
    .A1(_04650_),
    .A2(net4823));
 sg13g2_nand3_1 _19975_ (.B(net5255),
    .C(net4822),
    .A(net3091),
    .Y(_03581_));
 sg13g2_o21ai_1 _19976_ (.B1(_03581_),
    .Y(_01514_),
    .A1(_04651_),
    .A2(net4820));
 sg13g2_nand3_1 _19977_ (.B(net5252),
    .C(net4819),
    .A(net1998),
    .Y(_03582_));
 sg13g2_o21ai_1 _19978_ (.B1(_03582_),
    .Y(_01515_),
    .A1(_04652_),
    .A2(net4846));
 sg13g2_nand3_1 _19979_ (.B(net5258),
    .C(net4828),
    .A(net2177),
    .Y(_03583_));
 sg13g2_o21ai_1 _19980_ (.B1(_03583_),
    .Y(_01516_),
    .A1(_04653_),
    .A2(net4830));
 sg13g2_nand3_1 _19981_ (.B(net5259),
    .C(net4830),
    .A(net2081),
    .Y(_03584_));
 sg13g2_o21ai_1 _19982_ (.B1(_03584_),
    .Y(_01517_),
    .A1(_04654_),
    .A2(net4829));
 sg13g2_nand3_1 _19983_ (.B(net5259),
    .C(net4829),
    .A(net2296),
    .Y(_03585_));
 sg13g2_o21ai_1 _19984_ (.B1(_03585_),
    .Y(_01518_),
    .A1(_04655_),
    .A2(net4830));
 sg13g2_nand3_1 _19985_ (.B(net5259),
    .C(net4829),
    .A(net2436),
    .Y(_03586_));
 sg13g2_o21ai_1 _19986_ (.B1(_03586_),
    .Y(_01519_),
    .A1(_04656_),
    .A2(net4827));
 sg13g2_nand3_1 _19987_ (.B(net5258),
    .C(net4827),
    .A(net2639),
    .Y(_03587_));
 sg13g2_o21ai_1 _19988_ (.B1(_03587_),
    .Y(_01520_),
    .A1(_04657_),
    .A2(net4827));
 sg13g2_nand3_1 _19989_ (.B(net5243),
    .C(net4801),
    .A(net3180),
    .Y(_03588_));
 sg13g2_o21ai_1 _19990_ (.B1(_03588_),
    .Y(_01521_),
    .A1(_04658_),
    .A2(net4800));
 sg13g2_nand3_1 _19991_ (.B(net5244),
    .C(net4799),
    .A(net2865),
    .Y(_03589_));
 sg13g2_o21ai_1 _19992_ (.B1(_03589_),
    .Y(_01522_),
    .A1(_04659_),
    .A2(net4792));
 sg13g2_nand3_1 _19993_ (.B(net5240),
    .C(net4792),
    .A(net2380),
    .Y(_03590_));
 sg13g2_o21ai_1 _19994_ (.B1(_03590_),
    .Y(_01523_),
    .A1(_04660_),
    .A2(net4791));
 sg13g2_nand3_1 _19995_ (.B(net5239),
    .C(net4791),
    .A(net2424),
    .Y(_03591_));
 sg13g2_o21ai_1 _19996_ (.B1(_03591_),
    .Y(_01524_),
    .A1(_04661_),
    .A2(net4751));
 sg13g2_nand3_1 _19997_ (.B(net5222),
    .C(net4751),
    .A(net1138),
    .Y(_03592_));
 sg13g2_o21ai_1 _19998_ (.B1(_03592_),
    .Y(_01525_),
    .A1(_04662_),
    .A2(net4751));
 sg13g2_nand3_1 _19999_ (.B(net5220),
    .C(net4752),
    .A(net3425),
    .Y(_03593_));
 sg13g2_o21ai_1 _20000_ (.B1(_03593_),
    .Y(_01526_),
    .A1(_04663_),
    .A2(net4755));
 sg13g2_nand3_1 _20001_ (.B(net5223),
    .C(net4760),
    .A(net2669),
    .Y(_03594_));
 sg13g2_o21ai_1 _20002_ (.B1(_03594_),
    .Y(_01527_),
    .A1(_04664_),
    .A2(net4760));
 sg13g2_nand3_1 _20003_ (.B(net5224),
    .C(net4763),
    .A(net1935),
    .Y(_03595_));
 sg13g2_o21ai_1 _20004_ (.B1(_03595_),
    .Y(_01528_),
    .A1(_04665_),
    .A2(net4763));
 sg13g2_nand3_1 _20005_ (.B(net5225),
    .C(net4766),
    .A(net3225),
    .Y(_03596_));
 sg13g2_o21ai_1 _20006_ (.B1(_03596_),
    .Y(_01529_),
    .A1(_04666_),
    .A2(net4765));
 sg13g2_nand3_1 _20007_ (.B(net5228),
    .C(net4772),
    .A(net1410),
    .Y(_03597_));
 sg13g2_o21ai_1 _20008_ (.B1(_03597_),
    .Y(_01530_),
    .A1(_04667_),
    .A2(net4772));
 sg13g2_nand3_1 _20009_ (.B(net5228),
    .C(net4772),
    .A(net2165),
    .Y(_03598_));
 sg13g2_o21ai_1 _20010_ (.B1(_03598_),
    .Y(_01531_),
    .A1(_04668_),
    .A2(net4773));
 sg13g2_nand3_1 _20011_ (.B(net5227),
    .C(net4773),
    .A(net2382),
    .Y(_03599_));
 sg13g2_o21ai_1 _20012_ (.B1(_03599_),
    .Y(_01532_),
    .A1(_04669_),
    .A2(net4771));
 sg13g2_nand3_1 _20013_ (.B(net5229),
    .C(net4775),
    .A(net2286),
    .Y(_03600_));
 sg13g2_o21ai_1 _20014_ (.B1(_03600_),
    .Y(_01533_),
    .A1(_04670_),
    .A2(net4775));
 sg13g2_nand3_1 _20015_ (.B(net5233),
    .C(net4780),
    .A(net1751),
    .Y(_03601_));
 sg13g2_o21ai_1 _20016_ (.B1(_03601_),
    .Y(_01534_),
    .A1(_04671_),
    .A2(net4780));
 sg13g2_nand3_1 _20017_ (.B(net5234),
    .C(net4783),
    .A(net3078),
    .Y(_03602_));
 sg13g2_o21ai_1 _20018_ (.B1(_03602_),
    .Y(_01535_),
    .A1(_04672_),
    .A2(net4787));
 sg13g2_nand3_1 _20019_ (.B(net5235),
    .C(net4787),
    .A(net1212),
    .Y(_03603_));
 sg13g2_o21ai_1 _20020_ (.B1(_03603_),
    .Y(_01536_),
    .A1(_04673_),
    .A2(net4786));
 sg13g2_nand3_1 _20021_ (.B(net5285),
    .C(net4881),
    .A(net2290),
    .Y(_03604_));
 sg13g2_o21ai_1 _20022_ (.B1(_03604_),
    .Y(_01537_),
    .A1(_04674_),
    .A2(net4880));
 sg13g2_nand3_1 _20023_ (.B(net5289),
    .C(net4890),
    .A(net2519),
    .Y(_03605_));
 sg13g2_o21ai_1 _20024_ (.B1(_03605_),
    .Y(_01538_),
    .A1(_04675_),
    .A2(net4890));
 sg13g2_nand3_1 _20025_ (.B(net5290),
    .C(net4891),
    .A(net1245),
    .Y(_03606_));
 sg13g2_o21ai_1 _20026_ (.B1(_03606_),
    .Y(_01539_),
    .A1(_04676_),
    .A2(net4892));
 sg13g2_nand3_1 _20027_ (.B(net5298),
    .C(net4908),
    .A(net1911),
    .Y(_03607_));
 sg13g2_o21ai_1 _20028_ (.B1(_03607_),
    .Y(_01540_),
    .A1(_04677_),
    .A2(net4908));
 sg13g2_nand3_1 _20029_ (.B(net5298),
    .C(net4908),
    .A(net3282),
    .Y(_03608_));
 sg13g2_o21ai_1 _20030_ (.B1(_03608_),
    .Y(_01541_),
    .A1(_04678_),
    .A2(net4904));
 sg13g2_nand3_1 _20031_ (.B(net5294),
    .C(net4899),
    .A(net2121),
    .Y(_03609_));
 sg13g2_o21ai_1 _20032_ (.B1(_03609_),
    .Y(_01542_),
    .A1(_04679_),
    .A2(net4899));
 sg13g2_nand3_1 _20033_ (.B(net5294),
    .C(net4898),
    .A(net2347),
    .Y(_03610_));
 sg13g2_o21ai_1 _20034_ (.B1(_03610_),
    .Y(_01543_),
    .A1(_04680_),
    .A2(net4898));
 sg13g2_nand3_1 _20035_ (.B(net5293),
    .C(net4895),
    .A(net2508),
    .Y(_03611_));
 sg13g2_o21ai_1 _20036_ (.B1(_03611_),
    .Y(_01544_),
    .A1(_04681_),
    .A2(net4897));
 sg13g2_nand3_1 _20037_ (.B(net5279),
    .C(net4868),
    .A(net3365),
    .Y(_03612_));
 sg13g2_o21ai_1 _20038_ (.B1(_03612_),
    .Y(_01545_),
    .A1(_04682_),
    .A2(net4823));
 sg13g2_nand3_1 _20039_ (.B(net5254),
    .C(net4822),
    .A(net2730),
    .Y(_03613_));
 sg13g2_o21ai_1 _20040_ (.B1(_03613_),
    .Y(_01546_),
    .A1(_04683_),
    .A2(net4822));
 sg13g2_nand3_1 _20041_ (.B(net5252),
    .C(net4819),
    .A(net2237),
    .Y(_03614_));
 sg13g2_o21ai_1 _20042_ (.B1(_03614_),
    .Y(_01547_),
    .A1(_04684_),
    .A2(net4847));
 sg13g2_nand3_1 _20043_ (.B(net5269),
    .C(net4846),
    .A(net1298),
    .Y(_03615_));
 sg13g2_o21ai_1 _20044_ (.B1(_03615_),
    .Y(_01548_),
    .A1(_04685_),
    .A2(net4848));
 sg13g2_nand3_1 _20045_ (.B(net5265),
    .C(net4842),
    .A(net2533),
    .Y(_03616_));
 sg13g2_o21ai_1 _20046_ (.B1(_03616_),
    .Y(_01549_),
    .A1(_04686_),
    .A2(net4838));
 sg13g2_nand3_1 _20047_ (.B(net5263),
    .C(net4837),
    .A(net2349),
    .Y(_03617_));
 sg13g2_o21ai_1 _20048_ (.B1(_03617_),
    .Y(_01550_),
    .A1(_04687_),
    .A2(net4838));
 sg13g2_nand3_1 _20049_ (.B(net5258),
    .C(net4828),
    .A(net2991),
    .Y(_03618_));
 sg13g2_o21ai_1 _20050_ (.B1(_03618_),
    .Y(_01551_),
    .A1(_04688_),
    .A2(net4828));
 sg13g2_nand3_1 _20051_ (.B(net5243),
    .C(net4802),
    .A(net2916),
    .Y(_03619_));
 sg13g2_o21ai_1 _20052_ (.B1(_03619_),
    .Y(_01552_),
    .A1(_04689_),
    .A2(net4807));
 sg13g2_nand3_1 _20053_ (.B(net5243),
    .C(net4802),
    .A(net2683),
    .Y(_03620_));
 sg13g2_o21ai_1 _20054_ (.B1(_03620_),
    .Y(_01553_),
    .A1(_04690_),
    .A2(net4803));
 sg13g2_nand3_1 _20055_ (.B(net5245),
    .C(net4803),
    .A(net2034),
    .Y(_03621_));
 sg13g2_o21ai_1 _20056_ (.B1(_03621_),
    .Y(_01554_),
    .A1(_04691_),
    .A2(net4803));
 sg13g2_nand3_1 _20057_ (.B(net5242),
    .C(net4796),
    .A(net2136),
    .Y(_03622_));
 sg13g2_o21ai_1 _20058_ (.B1(_03622_),
    .Y(_01555_),
    .A1(_04692_),
    .A2(net4796));
 sg13g2_nand3_1 _20059_ (.B(net5241),
    .C(net4794),
    .A(net2435),
    .Y(_03623_));
 sg13g2_o21ai_1 _20060_ (.B1(_03623_),
    .Y(_01556_),
    .A1(_04693_),
    .A2(net4753));
 sg13g2_nand3_1 _20061_ (.B(net5220),
    .C(net4753),
    .A(net1198),
    .Y(_03624_));
 sg13g2_o21ai_1 _20062_ (.B1(_03624_),
    .Y(_01557_),
    .A1(_04694_),
    .A2(net4752));
 sg13g2_nand3_1 _20063_ (.B(net5220),
    .C(net4752),
    .A(net1286),
    .Y(_03625_));
 sg13g2_o21ai_1 _20064_ (.B1(_03625_),
    .Y(_01558_),
    .A1(_04695_),
    .A2(net4752));
 sg13g2_nand3_1 _20065_ (.B(net5220),
    .C(net4755),
    .A(net2255),
    .Y(_03626_));
 sg13g2_o21ai_1 _20066_ (.B1(_03626_),
    .Y(_01559_),
    .A1(_04696_),
    .A2(net4760));
 sg13g2_nand3_1 _20067_ (.B(net5248),
    .C(net4808),
    .A(net2356),
    .Y(_03627_));
 sg13g2_o21ai_1 _20068_ (.B1(_03627_),
    .Y(_01560_),
    .A1(_04697_),
    .A2(net4812));
 sg13g2_nand3_1 _20069_ (.B(net5249),
    .C(net4813),
    .A(net2627),
    .Y(_03628_));
 sg13g2_o21ai_1 _20070_ (.B1(_03628_),
    .Y(_01561_),
    .A1(_04698_),
    .A2(net4813));
 sg13g2_nand3_1 _20071_ (.B(net5250),
    .C(net4815),
    .A(net1959),
    .Y(_03629_));
 sg13g2_o21ai_1 _20072_ (.B1(_03629_),
    .Y(_01562_),
    .A1(_04699_),
    .A2(net4816));
 sg13g2_nand3_1 _20073_ (.B(net5249),
    .C(net4815),
    .A(net1290),
    .Y(_03630_));
 sg13g2_o21ai_1 _20074_ (.B1(_03630_),
    .Y(_01563_),
    .A1(_04700_),
    .A2(net4861));
 sg13g2_nand3_1 _20075_ (.B(net5275),
    .C(net4859),
    .A(net2554),
    .Y(_03631_));
 sg13g2_o21ai_1 _20076_ (.B1(_03631_),
    .Y(_01564_),
    .A1(_04701_),
    .A2(net4773));
 sg13g2_nand3_1 _20077_ (.B(net5230),
    .C(net4777),
    .A(net3027),
    .Y(_03632_));
 sg13g2_o21ai_1 _20078_ (.B1(_03632_),
    .Y(_01565_),
    .A1(_04702_),
    .A2(net4777));
 sg13g2_nand3_1 _20079_ (.B(net5230),
    .C(net4777),
    .A(net1140),
    .Y(_03633_));
 sg13g2_o21ai_1 _20080_ (.B1(_03633_),
    .Y(_01566_),
    .A1(_04703_),
    .A2(net4778));
 sg13g2_nand3_1 _20081_ (.B(net5234),
    .C(net4782),
    .A(net1166),
    .Y(_03634_));
 sg13g2_o21ai_1 _20082_ (.B1(_03634_),
    .Y(_01567_),
    .A1(_04704_),
    .A2(net4782));
 sg13g2_nand3_1 _20083_ (.B(net5284),
    .C(net4877),
    .A(net1197),
    .Y(_03635_));
 sg13g2_o21ai_1 _20084_ (.B1(_03635_),
    .Y(_01568_),
    .A1(_04705_),
    .A2(net4877));
 sg13g2_nand3_1 _20085_ (.B(net5286),
    .C(net4880),
    .A(net1172),
    .Y(_03636_));
 sg13g2_o21ai_1 _20086_ (.B1(_03636_),
    .Y(_01569_),
    .A1(_04706_),
    .A2(net4882));
 sg13g2_nand3_1 _20087_ (.B(net5286),
    .C(net4882),
    .A(net2525),
    .Y(_03637_));
 sg13g2_o21ai_1 _20088_ (.B1(_03637_),
    .Y(_01570_),
    .A1(_04707_),
    .A2(net4889));
 sg13g2_nand3_1 _20089_ (.B(net5289),
    .C(net4889),
    .A(net1602),
    .Y(_03638_));
 sg13g2_o21ai_1 _20090_ (.B1(_03638_),
    .Y(_01571_),
    .A1(_04708_),
    .A2(net4891));
 sg13g2_nand3_1 _20091_ (.B(net5298),
    .C(net4908),
    .A(net1393),
    .Y(_03639_));
 sg13g2_o21ai_1 _20092_ (.B1(_03639_),
    .Y(_01572_),
    .A1(_04709_),
    .A2(net4908));
 sg13g2_nand3_1 _20093_ (.B(net5298),
    .C(net4909),
    .A(net1916),
    .Y(_03640_));
 sg13g2_o21ai_1 _20094_ (.B1(_03640_),
    .Y(_01573_),
    .A1(_04710_),
    .A2(net4909));
 sg13g2_nand3_1 _20095_ (.B(net5297),
    .C(net4904),
    .A(\TRNG.Word_Out[329] ),
    .Y(_03641_));
 sg13g2_o21ai_1 _20096_ (.B1(_03641_),
    .Y(_01574_),
    .A1(_04711_),
    .A2(net4904));
 sg13g2_nand3_1 _20097_ (.B(net5287),
    .C(net4887),
    .A(net3098),
    .Y(_03642_));
 sg13g2_o21ai_1 _20098_ (.B1(_03642_),
    .Y(_01575_),
    .A1(_04712_),
    .A2(net4872));
 sg13g2_nand3_1 _20099_ (.B(net5278),
    .C(net4869),
    .A(net2556),
    .Y(_03643_));
 sg13g2_o21ai_1 _20100_ (.B1(_03643_),
    .Y(_01576_),
    .A1(_04713_),
    .A2(net4868));
 sg13g2_nand3_1 _20101_ (.B(net5279),
    .C(net4868),
    .A(net1680),
    .Y(_03644_));
 sg13g2_o21ai_1 _20102_ (.B1(_03644_),
    .Y(_01577_),
    .A1(_04714_),
    .A2(net4868));
 sg13g2_nand3_1 _20103_ (.B(net5270),
    .C(net4851),
    .A(net1154),
    .Y(_03645_));
 sg13g2_o21ai_1 _20104_ (.B1(_03645_),
    .Y(_01578_),
    .A1(_04715_),
    .A2(net4851));
 sg13g2_nand3_1 _20105_ (.B(net5270),
    .C(net4850),
    .A(net2101),
    .Y(_03646_));
 sg13g2_o21ai_1 _20106_ (.B1(_03646_),
    .Y(_01579_),
    .A1(_04716_),
    .A2(net4850));
 sg13g2_nand3_1 _20107_ (.B(net5259),
    .C(net4830),
    .A(net3206),
    .Y(_03647_));
 sg13g2_o21ai_1 _20108_ (.B1(_03647_),
    .Y(_01580_),
    .A1(_04717_),
    .A2(net4830));
 sg13g2_nand3_1 _20109_ (.B(net5259),
    .C(net4829),
    .A(net2199),
    .Y(_03648_));
 sg13g2_o21ai_1 _20110_ (.B1(_03648_),
    .Y(_01581_),
    .A1(_04718_),
    .A2(net4837));
 sg13g2_nand3_1 _20111_ (.B(net5263),
    .C(net4837),
    .A(net2638),
    .Y(_03649_));
 sg13g2_o21ai_1 _20112_ (.B1(_03649_),
    .Y(_01582_),
    .A1(_04719_),
    .A2(net4837));
 sg13g2_nand3_1 _20113_ (.B(net5259),
    .C(net4829),
    .A(net2629),
    .Y(_03650_));
 sg13g2_o21ai_1 _20114_ (.B1(_03650_),
    .Y(_01583_),
    .A1(_04720_),
    .A2(net4828));
 sg13g2_nand3_1 _20115_ (.B(net5258),
    .C(net4827),
    .A(net3125),
    .Y(_03651_));
 sg13g2_o21ai_1 _20116_ (.B1(_03651_),
    .Y(_01584_),
    .A1(_04721_),
    .A2(net4802));
 sg13g2_nand3_1 _20117_ (.B(net5243),
    .C(net4801),
    .A(net2770),
    .Y(_03652_));
 sg13g2_o21ai_1 _20118_ (.B1(_03652_),
    .Y(_01585_),
    .A1(_04722_),
    .A2(net4799));
 sg13g2_nand3_1 _20119_ (.B(net5244),
    .C(net4799),
    .A(net2597),
    .Y(_03653_));
 sg13g2_o21ai_1 _20120_ (.B1(_03653_),
    .Y(_01586_),
    .A1(_04723_),
    .A2(net4792));
 sg13g2_nand3_1 _20121_ (.B(net5240),
    .C(net4792),
    .A(net2184),
    .Y(_03654_));
 sg13g2_o21ai_1 _20122_ (.B1(_03654_),
    .Y(_01587_),
    .A1(_04724_),
    .A2(net4791));
 sg13g2_nand3_1 _20123_ (.B(net5239),
    .C(net4793),
    .A(net2776),
    .Y(_03655_));
 sg13g2_o21ai_1 _20124_ (.B1(_03655_),
    .Y(_01588_),
    .A1(_04725_),
    .A2(net4751));
 sg13g2_nand3_1 _20125_ (.B(net5222),
    .C(net4756),
    .A(net2292),
    .Y(_03656_));
 sg13g2_o21ai_1 _20126_ (.B1(_03656_),
    .Y(_01589_),
    .A1(_04726_),
    .A2(net4752));
 sg13g2_nand3_1 _20127_ (.B(net5220),
    .C(net4752),
    .A(net1164),
    .Y(_03657_));
 sg13g2_o21ai_1 _20128_ (.B1(_03657_),
    .Y(_01590_),
    .A1(_04727_),
    .A2(net4752));
 sg13g2_nand3_1 _20129_ (.B(net5225),
    .C(net4761),
    .A(net3381),
    .Y(_03658_));
 sg13g2_o21ai_1 _20130_ (.B1(_03658_),
    .Y(_01591_),
    .A1(_04728_),
    .A2(net4761));
 sg13g2_nand3_1 _20131_ (.B(net5224),
    .C(net4765),
    .A(net2461),
    .Y(_03659_));
 sg13g2_o21ai_1 _20132_ (.B1(_03659_),
    .Y(_01592_),
    .A1(_04729_),
    .A2(net4765));
 sg13g2_nand3_1 _20133_ (.B(net5224),
    .C(net4765),
    .A(net1185),
    .Y(_03660_));
 sg13g2_o21ai_1 _20134_ (.B1(_03660_),
    .Y(_01593_),
    .A1(_04730_),
    .A2(net4772));
 sg13g2_nand3_1 _20135_ (.B(net5275),
    .C(net4772),
    .A(net1381),
    .Y(_03661_));
 sg13g2_o21ai_1 _20136_ (.B1(_03661_),
    .Y(_01594_),
    .A1(_04731_),
    .A2(net4859));
 sg13g2_nand3_1 _20137_ (.B(net5275),
    .C(net4859),
    .A(net2076),
    .Y(_03662_));
 sg13g2_o21ai_1 _20138_ (.B1(_03662_),
    .Y(_01595_),
    .A1(_04732_),
    .A2(net4860));
 sg13g2_nand3_1 _20139_ (.B(net5275),
    .C(net4859),
    .A(net3185),
    .Y(_03663_));
 sg13g2_o21ai_1 _20140_ (.B1(_03663_),
    .Y(_01596_),
    .A1(_04733_),
    .A2(net4863));
 sg13g2_nand3_1 _20141_ (.B(net5277),
    .C(net4863),
    .A(net2087),
    .Y(_03664_));
 sg13g2_o21ai_1 _20142_ (.B1(_03664_),
    .Y(_01597_),
    .A1(_04734_),
    .A2(net4863));
 sg13g2_nand3_1 _20143_ (.B(net5277),
    .C(net4865),
    .A(net2071),
    .Y(_03665_));
 sg13g2_o21ai_1 _20144_ (.B1(_03665_),
    .Y(_01598_),
    .A1(_04735_),
    .A2(net4863));
 sg13g2_nand3_1 _20145_ (.B(net5284),
    .C(net4876),
    .A(net2491),
    .Y(_03666_));
 sg13g2_o21ai_1 _20146_ (.B1(_03666_),
    .Y(_01599_),
    .A1(_04736_),
    .A2(net4876));
 sg13g2_nand3_1 _20147_ (.B(net5285),
    .C(net4880),
    .A(net1187),
    .Y(_03667_));
 sg13g2_o21ai_1 _20148_ (.B1(_03667_),
    .Y(_01600_),
    .A1(_04737_),
    .A2(net4880));
 sg13g2_nand3_1 _20149_ (.B(net5286),
    .C(net4882),
    .A(net2451),
    .Y(_03668_));
 sg13g2_o21ai_1 _20150_ (.B1(_03668_),
    .Y(_01601_),
    .A1(_04738_),
    .A2(net4882));
 sg13g2_nand3_1 _20151_ (.B(net5289),
    .C(net4889),
    .A(net1599),
    .Y(_03669_));
 sg13g2_o21ai_1 _20152_ (.B1(_03669_),
    .Y(_01602_),
    .A1(_04739_),
    .A2(net4889));
 sg13g2_nand3_1 _20153_ (.B(net5290),
    .C(net4891),
    .A(net1991),
    .Y(_03670_));
 sg13g2_o21ai_1 _20154_ (.B1(_03670_),
    .Y(_01603_),
    .A1(_04740_),
    .A2(net4891));
 sg13g2_nand3_1 _20155_ (.B(net5290),
    .C(net4891),
    .A(net1219),
    .Y(_03671_));
 sg13g2_o21ai_1 _20156_ (.B1(_03671_),
    .Y(_01604_),
    .A1(_04741_),
    .A2(net4909));
 sg13g2_nand3_1 _20157_ (.B(net5297),
    .C(net4905),
    .A(net2599),
    .Y(_03672_));
 sg13g2_o21ai_1 _20158_ (.B1(_03672_),
    .Y(_01605_),
    .A1(_04742_),
    .A2(net4905));
 sg13g2_nand3_1 _20159_ (.B(net5297),
    .C(net4904),
    .A(net2588),
    .Y(_03673_));
 sg13g2_o21ai_1 _20160_ (.B1(_03673_),
    .Y(_01606_),
    .A1(_04743_),
    .A2(net4899));
 sg13g2_nand3_1 _20161_ (.B(net5294),
    .C(net4898),
    .A(net3129),
    .Y(_03674_));
 sg13g2_o21ai_1 _20162_ (.B1(_03674_),
    .Y(_01607_),
    .A1(_04744_),
    .A2(net4899));
 sg13g2_nand3_1 _20163_ (.B(net5293),
    .C(net4897),
    .A(net1982),
    .Y(_03675_));
 sg13g2_o21ai_1 _20164_ (.B1(_03675_),
    .Y(_01608_),
    .A1(_04745_),
    .A2(net4895));
 sg13g2_nand3_1 _20165_ (.B(net5293),
    .C(net4895),
    .A(net2610),
    .Y(_03676_));
 sg13g2_o21ai_1 _20166_ (.B1(_03676_),
    .Y(_01609_),
    .A1(_04746_),
    .A2(net4851));
 sg13g2_nand3_1 _20167_ (.B(net5270),
    .C(net4851),
    .A(net2139),
    .Y(_03677_));
 sg13g2_o21ai_1 _20168_ (.B1(_03677_),
    .Y(_01610_),
    .A1(_04747_),
    .A2(net4851));
 sg13g2_nand3_1 _20169_ (.B(net5270),
    .C(net4850),
    .A(net2452),
    .Y(_03678_));
 sg13g2_o21ai_1 _20170_ (.B1(_03678_),
    .Y(_01611_),
    .A1(_04748_),
    .A2(net4847));
 sg13g2_nand3_1 _20171_ (.B(net5265),
    .C(net4841),
    .A(net2561),
    .Y(_03679_));
 sg13g2_o21ai_1 _20172_ (.B1(_03679_),
    .Y(_01612_),
    .A1(_04749_),
    .A2(net4841));
 sg13g2_nand3_1 _20173_ (.B(net5263),
    .C(net4839),
    .A(net2128),
    .Y(_03680_));
 sg13g2_o21ai_1 _20174_ (.B1(_03680_),
    .Y(_01613_),
    .A1(_04750_),
    .A2(net4839));
 sg13g2_nand3_1 _20175_ (.B(net5264),
    .C(net4840),
    .A(net1985),
    .Y(_03681_));
 sg13g2_o21ai_1 _20176_ (.B1(_03681_),
    .Y(_01614_),
    .A1(_04751_),
    .A2(net4840));
 sg13g2_nand3_1 _20177_ (.B(net5264),
    .C(net4840),
    .A(net2843),
    .Y(_03682_));
 sg13g2_o21ai_1 _20178_ (.B1(_03682_),
    .Y(_01615_),
    .A1(_04752_),
    .A2(net4829));
 sg13g2_nand3_1 _20179_ (.B(net5258),
    .C(net4827),
    .A(net2584),
    .Y(_03683_));
 sg13g2_o21ai_1 _20180_ (.B1(_03683_),
    .Y(_01616_),
    .A1(_04753_),
    .A2(net4802));
 sg13g2_nand3_1 _20181_ (.B(net5243),
    .C(net4801),
    .A(net2684),
    .Y(_03684_));
 sg13g2_o21ai_1 _20182_ (.B1(_03684_),
    .Y(_01617_),
    .A1(_04754_),
    .A2(net4801));
 sg13g2_nand3_1 _20183_ (.B(net5244),
    .C(net4799),
    .A(net2414),
    .Y(_03685_));
 sg13g2_o21ai_1 _20184_ (.B1(_03685_),
    .Y(_01618_),
    .A1(_04755_),
    .A2(net4799));
 sg13g2_nand3_1 _20185_ (.B(net5240),
    .C(net4792),
    .A(net2228),
    .Y(_03686_));
 sg13g2_o21ai_1 _20186_ (.B1(_03686_),
    .Y(_01619_),
    .A1(_04756_),
    .A2(net4792));
 sg13g2_nand3_1 _20187_ (.B(net5239),
    .C(net4791),
    .A(net2078),
    .Y(_03687_));
 sg13g2_o21ai_1 _20188_ (.B1(_03687_),
    .Y(_01620_),
    .A1(_04757_),
    .A2(net4793));
 sg13g2_nand3_1 _20189_ (.B(net5241),
    .C(net4794),
    .A(net1178),
    .Y(_03688_));
 sg13g2_o21ai_1 _20190_ (.B1(_03688_),
    .Y(_01621_),
    .A1(_04758_),
    .A2(net4753));
 sg13g2_nand3_1 _20191_ (.B(net5220),
    .C(net4755),
    .A(net3313),
    .Y(_03689_));
 sg13g2_o21ai_1 _20192_ (.B1(_03689_),
    .Y(_01622_),
    .A1(_04759_),
    .A2(net4752));
 sg13g2_nand3_1 _20193_ (.B(net5223),
    .C(net4760),
    .A(net2455),
    .Y(_03690_));
 sg13g2_o21ai_1 _20194_ (.B1(_03690_),
    .Y(_01623_),
    .A1(_04760_),
    .A2(net4762));
 sg13g2_nand3_1 _20195_ (.B(net5225),
    .C(net4762),
    .A(net2594),
    .Y(_03691_));
 sg13g2_o21ai_1 _20196_ (.B1(_03691_),
    .Y(_01624_),
    .A1(_04761_),
    .A2(net4765));
 sg13g2_nand3_1 _20197_ (.B(net5224),
    .C(net4765),
    .A(net2497),
    .Y(_03692_));
 sg13g2_o21ai_1 _20198_ (.B1(_03692_),
    .Y(_01625_),
    .A1(_04762_),
    .A2(net4765));
 sg13g2_nand3_1 _20199_ (.B(net5249),
    .C(net4813),
    .A(net1204),
    .Y(_03693_));
 sg13g2_o21ai_1 _20200_ (.B1(_03693_),
    .Y(_01626_),
    .A1(_04763_),
    .A2(net4859));
 sg13g2_nand3_1 _20201_ (.B(net5275),
    .C(net4859),
    .A(net2896),
    .Y(_03694_));
 sg13g2_o21ai_1 _20202_ (.B1(_03694_),
    .Y(_01627_),
    .A1(_04764_),
    .A2(net4860));
 sg13g2_nand3_1 _20203_ (.B(net5276),
    .C(net4861),
    .A(net2689),
    .Y(_03695_));
 sg13g2_o21ai_1 _20204_ (.B1(_03695_),
    .Y(_01628_),
    .A1(_04765_),
    .A2(net4864));
 sg13g2_nand3_1 _20205_ (.B(net5282),
    .C(net4864),
    .A(net1818),
    .Y(_03696_));
 sg13g2_o21ai_1 _20206_ (.B1(_03696_),
    .Y(_01629_),
    .A1(_04766_),
    .A2(net4864));
 sg13g2_nand3_1 _20207_ (.B(net5277),
    .C(net4865),
    .A(net2157),
    .Y(_03697_));
 sg13g2_o21ai_1 _20208_ (.B1(_03697_),
    .Y(_01630_),
    .A1(_04767_),
    .A2(net4864));
 sg13g2_nand3_1 _20209_ (.B(net5277),
    .C(net4863),
    .A(net2288),
    .Y(_03698_));
 sg13g2_o21ai_1 _20210_ (.B1(_03698_),
    .Y(_01631_),
    .A1(_04768_),
    .A2(net4876));
 sg13g2_nand3_1 _20211_ (.B(net5283),
    .C(net4878),
    .A(net1607),
    .Y(_03699_));
 sg13g2_o21ai_1 _20212_ (.B1(_03699_),
    .Y(_01632_),
    .A1(_04769_),
    .A2(net4878));
 sg13g2_nand3_1 _20213_ (.B(net5283),
    .C(net4878),
    .A(net1425),
    .Y(_03700_));
 sg13g2_o21ai_1 _20214_ (.B1(_03700_),
    .Y(_01633_),
    .A1(_04770_),
    .A2(net4879));
 sg13g2_nand3_1 _20215_ (.B(net5283),
    .C(net4879),
    .A(net1174),
    .Y(_03701_));
 sg13g2_o21ai_1 _20216_ (.B1(_03701_),
    .Y(_01634_),
    .A1(_04771_),
    .A2(net4879));
 sg13g2_nand3_1 _20217_ (.B(net5287),
    .C(net4885),
    .A(net1661),
    .Y(_03702_));
 sg13g2_o21ai_1 _20218_ (.B1(_03702_),
    .Y(_01635_),
    .A1(_04772_),
    .A2(net4885));
 sg13g2_nand3_1 _20219_ (.B(net5287),
    .C(net4885),
    .A(net2449),
    .Y(_03703_));
 sg13g2_o21ai_1 _20220_ (.B1(_03703_),
    .Y(_01636_),
    .A1(_04773_),
    .A2(net4885));
 sg13g2_nand3_1 _20221_ (.B(net5280),
    .C(net4874),
    .A(net3279),
    .Y(_03704_));
 sg13g2_o21ai_1 _20222_ (.B1(_03704_),
    .Y(_01637_),
    .A1(_04774_),
    .A2(net4874));
 sg13g2_nand3_1 _20223_ (.B(net5280),
    .C(net4871),
    .A(net1232),
    .Y(_03705_));
 sg13g2_o21ai_1 _20224_ (.B1(_03705_),
    .Y(_01638_),
    .A1(_04775_),
    .A2(net4871));
 sg13g2_nand3_1 _20225_ (.B(net5278),
    .C(net4867),
    .A(net2587),
    .Y(_03706_));
 sg13g2_o21ai_1 _20226_ (.B1(_03706_),
    .Y(_01639_),
    .A1(_04776_),
    .A2(net4867));
 sg13g2_nand3_1 _20227_ (.B(net5278),
    .C(net4866),
    .A(net1387),
    .Y(_03707_));
 sg13g2_o21ai_1 _20228_ (.B1(_03707_),
    .Y(_01640_),
    .A1(_04777_),
    .A2(net4866));
 sg13g2_nand3_1 _20229_ (.B(net5254),
    .C(net4824),
    .A(net2976),
    .Y(_03708_));
 sg13g2_o21ai_1 _20230_ (.B1(_03708_),
    .Y(_01641_),
    .A1(_04778_),
    .A2(net4821));
 sg13g2_nand3_1 _20231_ (.B(net5254),
    .C(net4821),
    .A(net1227),
    .Y(_03709_));
 sg13g2_o21ai_1 _20232_ (.B1(_03709_),
    .Y(_01642_),
    .A1(_04779_),
    .A2(net4850));
 sg13g2_nand3_1 _20233_ (.B(net5270),
    .C(net4850),
    .A(net2002),
    .Y(_03710_));
 sg13g2_o21ai_1 _20234_ (.B1(_03710_),
    .Y(_01643_),
    .A1(_04780_),
    .A2(net4850));
 sg13g2_nand3_1 _20235_ (.B(net5269),
    .C(net4849),
    .A(net2879),
    .Y(_03711_));
 sg13g2_o21ai_1 _20236_ (.B1(_03711_),
    .Y(_01644_),
    .A1(_04781_),
    .A2(net4842));
 sg13g2_nand3_1 _20237_ (.B(net5265),
    .C(net4841),
    .A(net1471),
    .Y(_03712_));
 sg13g2_o21ai_1 _20238_ (.B1(_03712_),
    .Y(_01645_),
    .A1(_04782_),
    .A2(net4841));
 sg13g2_nand3_1 _20239_ (.B(net5263),
    .C(net4838),
    .A(net2294),
    .Y(_03713_));
 sg13g2_o21ai_1 _20240_ (.B1(_03713_),
    .Y(_01646_),
    .A1(_04783_),
    .A2(net4838));
 sg13g2_nand3_1 _20241_ (.B(net5259),
    .C(net4829),
    .A(net2907),
    .Y(_03714_));
 sg13g2_o21ai_1 _20242_ (.B1(_03714_),
    .Y(_01647_),
    .A1(_04784_),
    .A2(net4829));
 sg13g2_nand3_1 _20243_ (.B(net5243),
    .C(net4801),
    .A(net3263),
    .Y(_03715_));
 sg13g2_o21ai_1 _20244_ (.B1(_03715_),
    .Y(_01648_),
    .A1(_04785_),
    .A2(net4801));
 sg13g2_nand3_1 _20245_ (.B(net5243),
    .C(net4801),
    .A(net2881),
    .Y(_03716_));
 sg13g2_o21ai_1 _20246_ (.B1(_03716_),
    .Y(_01649_),
    .A1(_04786_),
    .A2(net4799));
 sg13g2_nand3_1 _20247_ (.B(net5244),
    .C(net4799),
    .A(net1874),
    .Y(_03717_));
 sg13g2_o21ai_1 _20248_ (.B1(_03717_),
    .Y(_01650_),
    .A1(_04787_),
    .A2(net4799));
 sg13g2_nand3_1 _20249_ (.B(net5239),
    .C(net4791),
    .A(net2534),
    .Y(_03718_));
 sg13g2_o21ai_1 _20250_ (.B1(_03718_),
    .Y(_01651_),
    .A1(_04788_),
    .A2(net4791));
 sg13g2_nand3_1 _20251_ (.B(net5239),
    .C(net4791),
    .A(net2614),
    .Y(_03719_));
 sg13g2_o21ai_1 _20252_ (.B1(_03719_),
    .Y(_01652_),
    .A1(_04789_),
    .A2(net4751));
 sg13g2_nand3_1 _20253_ (.B(net5222),
    .C(net4751),
    .A(net2490),
    .Y(_03720_));
 sg13g2_o21ai_1 _20254_ (.B1(_03720_),
    .Y(_01653_),
    .A1(_04790_),
    .A2(net4756));
 sg13g2_nand3_1 _20255_ (.B(net5221),
    .C(net4753),
    .A(net1168),
    .Y(_03721_));
 sg13g2_o21ai_1 _20256_ (.B1(_03721_),
    .Y(_01654_),
    .A1(_04791_),
    .A2(net4754));
 sg13g2_nand3_1 _20257_ (.B(net5221),
    .C(net4754),
    .A(\TRNG.Word_Out[410] ),
    .Y(_03722_));
 sg13g2_o21ai_1 _20258_ (.B1(_03722_),
    .Y(_01655_),
    .A1(_04792_),
    .A2(net4761));
 sg13g2_nand3_1 _20259_ (.B(net5223),
    .C(net4761),
    .A(net2943),
    .Y(_03723_));
 sg13g2_o21ai_1 _20260_ (.B1(_03723_),
    .Y(_01656_),
    .A1(_04793_),
    .A2(net4765));
 sg13g2_nand3_1 _20261_ (.B(net5250),
    .C(net4815),
    .A(net2641),
    .Y(_03724_));
 sg13g2_o21ai_1 _20262_ (.B1(_03724_),
    .Y(_01657_),
    .A1(_04794_),
    .A2(net4815));
 sg13g2_nand3_1 _20263_ (.B(net5249),
    .C(net4815),
    .A(net1398),
    .Y(_03725_));
 sg13g2_o21ai_1 _20264_ (.B1(_03725_),
    .Y(_01658_),
    .A1(_04795_),
    .A2(net4815));
 sg13g2_nand3_1 _20265_ (.B(net5254),
    .C(net4821),
    .A(net2391),
    .Y(_03726_));
 sg13g2_o21ai_1 _20266_ (.B1(_03726_),
    .Y(_01659_),
    .A1(_04796_),
    .A2(net4855));
 sg13g2_nand3_1 _20267_ (.B(net5272),
    .C(net4855),
    .A(net2030),
    .Y(_03727_));
 sg13g2_o21ai_1 _20268_ (.B1(_03727_),
    .Y(_01660_),
    .A1(_04797_),
    .A2(net4855));
 sg13g2_nand3_1 _20269_ (.B(net5272),
    .C(net4855),
    .A(net2905),
    .Y(_03728_));
 sg13g2_o21ai_1 _20270_ (.B1(_03728_),
    .Y(_01661_),
    .A1(_04798_),
    .A2(net4901));
 sg13g2_nand3_1 _20271_ (.B(net5296),
    .C(net4903),
    .A(net2161),
    .Y(_03729_));
 sg13g2_o21ai_1 _20272_ (.B1(_03729_),
    .Y(_01662_),
    .A1(_04799_),
    .A2(net4901));
 sg13g2_nand3_1 _20273_ (.B(net5296),
    .C(net4903),
    .A(net2370),
    .Y(_03730_));
 sg13g2_o21ai_1 _20274_ (.B1(_03730_),
    .Y(_01663_),
    .A1(_04800_),
    .A2(net4903));
 sg13g2_nand3_1 _20275_ (.B(net5301),
    .C(net4912),
    .A(net2755),
    .Y(_03731_));
 sg13g2_o21ai_1 _20276_ (.B1(_03731_),
    .Y(_01664_),
    .A1(_04801_),
    .A2(net4911));
 sg13g2_nand3_1 _20277_ (.B(net5301),
    .C(net4911),
    .A(net1633),
    .Y(_03732_));
 sg13g2_o21ai_1 _20278_ (.B1(_03732_),
    .Y(_01665_),
    .A1(_04802_),
    .A2(net4911));
 sg13g2_nand3_1 _20279_ (.B(net5301),
    .C(net4911),
    .A(net2421),
    .Y(_03733_));
 sg13g2_o21ai_1 _20280_ (.B1(_03733_),
    .Y(_01666_),
    .A1(_04803_),
    .A2(net4906));
 sg13g2_nand3_1 _20281_ (.B(net5297),
    .C(net4906),
    .A(net2245),
    .Y(_03734_));
 sg13g2_o21ai_1 _20282_ (.B1(_03734_),
    .Y(_01667_),
    .A1(_04804_),
    .A2(net4906));
 sg13g2_nand3_1 _20283_ (.B(net5297),
    .C(net4906),
    .A(net2024),
    .Y(_03735_));
 sg13g2_o21ai_1 _20284_ (.B1(_03735_),
    .Y(_01668_),
    .A1(_04805_),
    .A2(net4906));
 sg13g2_nand3_1 _20285_ (.B(net5296),
    .C(net4901),
    .A(net2231),
    .Y(_03736_));
 sg13g2_o21ai_1 _20286_ (.B1(_03736_),
    .Y(_01669_),
    .A1(_04806_),
    .A2(net4901));
 sg13g2_nand3_1 _20287_ (.B(net5302),
    .C(net4902),
    .A(net2749),
    .Y(_03737_));
 sg13g2_o21ai_1 _20288_ (.B1(_03737_),
    .Y(_01670_),
    .A1(_04807_),
    .A2(net4902));
 sg13g2_nand3_1 _20289_ (.B(net5296),
    .C(net4902),
    .A(net1469),
    .Y(_03738_));
 sg13g2_o21ai_1 _20290_ (.B1(_03738_),
    .Y(_01671_),
    .A1(_04808_),
    .A2(net4902));
 sg13g2_nand3_1 _20291_ (.B(net5272),
    .C(net4856),
    .A(net2273),
    .Y(_03739_));
 sg13g2_o21ai_1 _20292_ (.B1(_03739_),
    .Y(_01672_),
    .A1(_04809_),
    .A2(net4855));
 sg13g2_nand3_1 _20293_ (.B(net5272),
    .C(net4856),
    .A(net1650),
    .Y(_03740_));
 sg13g2_o21ai_1 _20294_ (.B1(_03740_),
    .Y(_01673_),
    .A1(_04810_),
    .A2(net4856));
 sg13g2_nand3_1 _20295_ (.B(net5272),
    .C(net4856),
    .A(net2279),
    .Y(_03741_));
 sg13g2_o21ai_1 _20296_ (.B1(_03741_),
    .Y(_01674_),
    .A1(_04811_),
    .A2(net4855));
 sg13g2_nand3_1 _20297_ (.B(net5273),
    .C(net4856),
    .A(net1795),
    .Y(_03742_));
 sg13g2_o21ai_1 _20298_ (.B1(_03742_),
    .Y(_01675_),
    .A1(_04812_),
    .A2(net4857));
 sg13g2_nand3_1 _20299_ (.B(net5273),
    .C(net4857),
    .A(net2132),
    .Y(_03743_));
 sg13g2_o21ai_1 _20300_ (.B1(_03743_),
    .Y(_01676_),
    .A1(_04813_),
    .A2(net4857));
 sg13g2_nand3_1 _20301_ (.B(net5266),
    .C(net4843),
    .A(net3040),
    .Y(_03744_));
 sg13g2_o21ai_1 _20302_ (.B1(_03744_),
    .Y(_01677_),
    .A1(_04814_),
    .A2(net4844));
 sg13g2_nand3_1 _20303_ (.B(net5266),
    .C(net4844),
    .A(net2298),
    .Y(_03745_));
 sg13g2_o21ai_1 _20304_ (.B1(_03745_),
    .Y(_01678_),
    .A1(_04815_),
    .A2(net4843));
 sg13g2_nand3_1 _20305_ (.B(net5266),
    .C(net4843),
    .A(net1913),
    .Y(_03746_));
 sg13g2_o21ai_1 _20306_ (.B1(_03746_),
    .Y(_01679_),
    .A1(_04816_),
    .A2(net4839));
 sg13g2_nand3_1 _20307_ (.B(net5263),
    .C(net4839),
    .A(net1804),
    .Y(_03747_));
 sg13g2_o21ai_1 _20308_ (.B1(_03747_),
    .Y(_01680_),
    .A1(_04817_),
    .A2(net4839));
 sg13g2_nand3_1 _20309_ (.B(net5266),
    .C(net4843),
    .A(net2346),
    .Y(_03748_));
 sg13g2_o21ai_1 _20310_ (.B1(_03748_),
    .Y(_01681_),
    .A1(_04818_),
    .A2(net4843));
 sg13g2_nand3_1 _20311_ (.B(net5266),
    .C(net4843),
    .A(net2143),
    .Y(_03749_));
 sg13g2_o21ai_1 _20312_ (.B1(_03749_),
    .Y(_01682_),
    .A1(_04819_),
    .A2(net4843));
 sg13g2_nand3_1 _20313_ (.B(net5265),
    .C(net4843),
    .A(net2026),
    .Y(_03750_));
 sg13g2_o21ai_1 _20314_ (.B1(_03750_),
    .Y(_01683_),
    .A1(_04820_),
    .A2(net4854));
 sg13g2_nand3_1 _20315_ (.B(net5272),
    .C(net4857),
    .A(net3034),
    .Y(_03751_));
 sg13g2_o21ai_1 _20316_ (.B1(_03751_),
    .Y(_01684_),
    .A1(_04821_),
    .A2(net4856));
 sg13g2_nand3_1 _20317_ (.B(net5272),
    .C(net4856),
    .A(net2514),
    .Y(_03752_));
 sg13g2_o21ai_1 _20318_ (.B1(_03752_),
    .Y(_01685_),
    .A1(_04822_),
    .A2(net4902));
 sg13g2_nand3_1 _20319_ (.B(net5296),
    .C(net4902),
    .A(net2116),
    .Y(_03753_));
 sg13g2_o21ai_1 _20320_ (.B1(_03753_),
    .Y(_01686_),
    .A1(_04823_),
    .A2(net4902));
 sg13g2_nand3_1 _20321_ (.B(net5296),
    .C(net4901),
    .A(net2572),
    .Y(_03754_));
 sg13g2_o21ai_1 _20322_ (.B1(_03754_),
    .Y(_01687_),
    .A1(_04824_),
    .A2(net4901));
 sg13g2_nand3_1 _20323_ (.B(net5296),
    .C(net4901),
    .A(net2163),
    .Y(_03755_));
 sg13g2_o21ai_1 _20324_ (.B1(_03755_),
    .Y(_01688_),
    .A1(_04825_),
    .A2(net4901));
 sg13g2_nand3_1 _20325_ (.B(net5301),
    .C(net4911),
    .A(net2316),
    .Y(_03756_));
 sg13g2_o21ai_1 _20326_ (.B1(_03756_),
    .Y(_01689_),
    .A1(_04826_),
    .A2(net4911));
 sg13g2_nand3_1 _20327_ (.B(net5301),
    .C(net4911),
    .A(net2217),
    .Y(_03757_));
 sg13g2_o21ai_1 _20328_ (.B1(_03757_),
    .Y(_01690_),
    .A1(_04828_),
    .A2(net4911));
 sg13g2_nor2_1 _20329_ (.A(net5237),
    .B(net5219),
    .Y(_03758_));
 sg13g2_nor2_1 _20330_ (.A(net3449),
    .B(_03758_),
    .Y(_03759_));
 sg13g2_a21oi_1 _20331_ (.A1(_04306_),
    .A2(_03758_),
    .Y(_01691_),
    .B1(_03759_));
 sg13g2_nand2b_1 _20332_ (.Y(_01692_),
    .B(net4681),
    .A_N(net3640));
 sg13g2_nand2_1 _20333_ (.Y(_03760_),
    .A(net1838),
    .B(net4597));
 sg13g2_o21ai_1 _20334_ (.B1(_03760_),
    .Y(_01693_),
    .A1(_04381_),
    .A2(net4597));
 sg13g2_nand2_1 _20335_ (.Y(_03761_),
    .A(net1950),
    .B(net4593));
 sg13g2_o21ai_1 _20336_ (.B1(_03761_),
    .Y(_01694_),
    .A1(_04382_),
    .A2(net4597));
 sg13g2_nand2_1 _20337_ (.Y(_03762_),
    .A(net3589),
    .B(net4681));
 sg13g2_o21ai_1 _20338_ (.B1(_03762_),
    .Y(_01695_),
    .A1(_04383_),
    .A2(net4682));
 sg13g2_nand2_1 _20339_ (.Y(_03763_),
    .A(net1827),
    .B(net4600));
 sg13g2_o21ai_1 _20340_ (.B1(_03763_),
    .Y(_01696_),
    .A1(_04384_),
    .A2(net4600));
 sg13g2_nand2_1 _20341_ (.Y(_03764_),
    .A(net1402),
    .B(net4695));
 sg13g2_o21ai_1 _20342_ (.B1(_03764_),
    .Y(_01697_),
    .A1(_04385_),
    .A2(net4695));
 sg13g2_nand2_1 _20343_ (.Y(_03765_),
    .A(net1757),
    .B(net4698));
 sg13g2_o21ai_1 _20344_ (.B1(_03765_),
    .Y(_01698_),
    .A1(_04386_),
    .A2(net4698));
 sg13g2_nand2_1 _20345_ (.Y(_03766_),
    .A(net1699),
    .B(net4704));
 sg13g2_o21ai_1 _20346_ (.B1(_03766_),
    .Y(_01699_),
    .A1(_04387_),
    .A2(net4704));
 sg13g2_nand2_1 _20347_ (.Y(_03767_),
    .A(net1704),
    .B(net4702));
 sg13g2_o21ai_1 _20348_ (.B1(_03767_),
    .Y(_01700_),
    .A1(_04388_),
    .A2(net4701));
 sg13g2_nand2_1 _20349_ (.Y(_03768_),
    .A(net1553),
    .B(net4701));
 sg13g2_o21ai_1 _20350_ (.B1(_03768_),
    .Y(_01701_),
    .A1(_04389_),
    .A2(net4701));
 sg13g2_nand2_1 _20351_ (.Y(_03769_),
    .A(net1440),
    .B(net4686));
 sg13g2_o21ai_1 _20352_ (.B1(_03769_),
    .Y(_01702_),
    .A1(_04390_),
    .A2(net4687));
 sg13g2_nand2_1 _20353_ (.Y(_03770_),
    .A(net1674),
    .B(net4714));
 sg13g2_o21ai_1 _20354_ (.B1(_03770_),
    .Y(_01703_),
    .A1(_04391_),
    .A2(net4714));
 sg13g2_nand2_1 _20355_ (.Y(_03771_),
    .A(net1952),
    .B(net4685));
 sg13g2_o21ai_1 _20356_ (.B1(_03771_),
    .Y(_01704_),
    .A1(_04392_),
    .A2(net4685));
 sg13g2_nand2_1 _20357_ (.Y(_03772_),
    .A(net1989),
    .B(net4640));
 sg13g2_o21ai_1 _20358_ (.B1(_03772_),
    .Y(_01705_),
    .A1(_04393_),
    .A2(net4640));
 sg13g2_nand2_1 _20359_ (.Y(_03773_),
    .A(net1424),
    .B(net4639));
 sg13g2_o21ai_1 _20360_ (.B1(_03773_),
    .Y(_01706_),
    .A1(_04394_),
    .A2(net4639));
 sg13g2_nand2_1 _20361_ (.Y(_03774_),
    .A(net1259),
    .B(net4636));
 sg13g2_o21ai_1 _20362_ (.B1(_03774_),
    .Y(_01707_),
    .A1(_04395_),
    .A2(net4636));
 sg13g2_nand2_1 _20363_ (.Y(_03775_),
    .A(net1478),
    .B(net4661));
 sg13g2_o21ai_1 _20364_ (.B1(_03775_),
    .Y(_01708_),
    .A1(_04396_),
    .A2(net4661));
 sg13g2_nand2_1 _20365_ (.Y(_03776_),
    .A(net1884),
    .B(net4663));
 sg13g2_o21ai_1 _20366_ (.B1(_03776_),
    .Y(_01709_),
    .A1(_04397_),
    .A2(net4663));
 sg13g2_nand2_1 _20367_ (.Y(_03777_),
    .A(net2174),
    .B(net4647));
 sg13g2_o21ai_1 _20368_ (.B1(_03777_),
    .Y(_01710_),
    .A1(_04398_),
    .A2(net4647));
 sg13g2_nand2_1 _20369_ (.Y(_03778_),
    .A(net1697),
    .B(net4651));
 sg13g2_o21ai_1 _20370_ (.B1(_03778_),
    .Y(_01711_),
    .A1(_04399_),
    .A2(net4648));
 sg13g2_nand2_1 _20371_ (.Y(_03779_),
    .A(net1537),
    .B(net4645));
 sg13g2_o21ai_1 _20372_ (.B1(_03779_),
    .Y(_01712_),
    .A1(_04400_),
    .A2(net4645));
 sg13g2_nand2_1 _20373_ (.Y(_03780_),
    .A(net1539),
    .B(net4620));
 sg13g2_o21ai_1 _20374_ (.B1(_03780_),
    .Y(_01713_),
    .A1(_04401_),
    .A2(net4620));
 sg13g2_nand2_1 _20375_ (.Y(_03781_),
    .A(net1418),
    .B(net4616));
 sg13g2_o21ai_1 _20376_ (.B1(_03781_),
    .Y(_01714_),
    .A1(_04402_),
    .A2(net4616));
 sg13g2_nand2_1 _20377_ (.Y(_03782_),
    .A(net1518),
    .B(net4608));
 sg13g2_o21ai_1 _20378_ (.B1(_03782_),
    .Y(_01715_),
    .A1(_04403_),
    .A2(net4608));
 sg13g2_nand2_1 _20379_ (.Y(_03783_),
    .A(net1292),
    .B(net4608));
 sg13g2_o21ai_1 _20380_ (.B1(_03783_),
    .Y(_01716_),
    .A1(_04404_),
    .A2(net4609));
 sg13g2_nand2_1 _20381_ (.Y(_03784_),
    .A(net2389),
    .B(net4610));
 sg13g2_o21ai_1 _20382_ (.B1(_03784_),
    .Y(_01717_),
    .A1(_04405_),
    .A2(net4610));
 sg13g2_nand2_1 _20383_ (.Y(_03785_),
    .A(net1400),
    .B(net4611));
 sg13g2_o21ai_1 _20384_ (.B1(_03785_),
    .Y(_01718_),
    .A1(_04406_),
    .A2(net4611));
 sg13g2_nand2_1 _20385_ (.Y(_03786_),
    .A(net2066),
    .B(net4573));
 sg13g2_o21ai_1 _20386_ (.B1(_03786_),
    .Y(_01719_),
    .A1(_04407_),
    .A2(net4573));
 sg13g2_nand2_1 _20387_ (.Y(_03787_),
    .A(net2314),
    .B(net4578));
 sg13g2_o21ai_1 _20388_ (.B1(_03787_),
    .Y(_01720_),
    .A1(_04408_),
    .A2(net4578));
 sg13g2_nand2_1 _20389_ (.Y(_03788_),
    .A(net1389),
    .B(net4582));
 sg13g2_o21ai_1 _20390_ (.B1(_03788_),
    .Y(_01721_),
    .A1(_04409_),
    .A2(net4582));
 sg13g2_nand2_1 _20391_ (.Y(_03789_),
    .A(net2390),
    .B(net4583));
 sg13g2_o21ai_1 _20392_ (.B1(_03789_),
    .Y(_01722_),
    .A1(_04410_),
    .A2(net4582));
 sg13g2_nand2_1 _20393_ (.Y(_03790_),
    .A(net1900),
    .B(net4589));
 sg13g2_o21ai_1 _20394_ (.B1(_03790_),
    .Y(_01723_),
    .A1(_04411_),
    .A2(net4589));
 sg13g2_nand2_1 _20395_ (.Y(_03791_),
    .A(net2085),
    .B(net4590));
 sg13g2_o21ai_1 _20396_ (.B1(_03791_),
    .Y(_01724_),
    .A1(_04412_),
    .A2(net4590));
 sg13g2_nand2_1 _20397_ (.Y(_03792_),
    .A(net2186),
    .B(net4593));
 sg13g2_o21ai_1 _20398_ (.B1(_03792_),
    .Y(_01725_),
    .A1(_04413_),
    .A2(net4593));
 sg13g2_nand2_1 _20399_ (.Y(_03793_),
    .A(net2050),
    .B(net4593));
 sg13g2_o21ai_1 _20400_ (.B1(_03793_),
    .Y(_01726_),
    .A1(_04414_),
    .A2(net4593));
 sg13g2_nand2_1 _20401_ (.Y(_03794_),
    .A(net1957),
    .B(net4601));
 sg13g2_o21ai_1 _20402_ (.B1(_03794_),
    .Y(_01727_),
    .A1(_04415_),
    .A2(net4598));
 sg13g2_nand2_1 _20403_ (.Y(_03795_),
    .A(net1845),
    .B(net4603));
 sg13g2_o21ai_1 _20404_ (.B1(_03795_),
    .Y(_01728_),
    .A1(_04416_),
    .A2(net4602));
 sg13g2_nand2_1 _20405_ (.Y(_03796_),
    .A(net2047),
    .B(net4696));
 sg13g2_o21ai_1 _20406_ (.B1(_03796_),
    .Y(_01729_),
    .A1(_04417_),
    .A2(net4604));
 sg13g2_nand2_1 _20407_ (.Y(_03797_),
    .A(net2581),
    .B(net4697));
 sg13g2_o21ai_1 _20408_ (.B1(_03797_),
    .Y(_01730_),
    .A1(_04418_),
    .A2(net4697));
 sg13g2_nand2_1 _20409_ (.Y(_03798_),
    .A(net2107),
    .B(net4705));
 sg13g2_o21ai_1 _20410_ (.B1(_03798_),
    .Y(_01731_),
    .A1(_04419_),
    .A2(net4705));
 sg13g2_nand2_1 _20411_ (.Y(_03799_),
    .A(net2119),
    .B(net4707));
 sg13g2_o21ai_1 _20412_ (.B1(_03799_),
    .Y(_01732_),
    .A1(_04420_),
    .A2(net4706));
 sg13g2_nand2_1 _20413_ (.Y(_03800_),
    .A(net2473),
    .B(net4728));
 sg13g2_o21ai_1 _20414_ (.B1(_03800_),
    .Y(_01733_),
    .A1(_04421_),
    .A2(net4728));
 sg13g2_nand2_1 _20415_ (.Y(_03801_),
    .A(net2149),
    .B(net4727));
 sg13g2_o21ai_1 _20416_ (.B1(_03801_),
    .Y(_01734_),
    .A1(_04422_),
    .A2(net4727));
 sg13g2_nand2_1 _20417_ (.Y(_03802_),
    .A(net1761),
    .B(net4724));
 sg13g2_o21ai_1 _20418_ (.B1(_03802_),
    .Y(_01735_),
    .A1(_04423_),
    .A2(net4724));
 sg13g2_nand2_1 _20419_ (.Y(_03803_),
    .A(net2088),
    .B(net4716));
 sg13g2_o21ai_1 _20420_ (.B1(_03803_),
    .Y(_01736_),
    .A1(_04424_),
    .A2(net4716));
 sg13g2_nand2_1 _20421_ (.Y(_03804_),
    .A(net2182),
    .B(net4712));
 sg13g2_o21ai_1 _20422_ (.B1(_03804_),
    .Y(_01737_),
    .A1(_04425_),
    .A2(net4713));
 sg13g2_nand2_1 _20423_ (.Y(_03805_),
    .A(net2131),
    .B(net4712));
 sg13g2_o21ai_1 _20424_ (.B1(_03805_),
    .Y(_01738_),
    .A1(_04426_),
    .A2(net4712));
 sg13g2_nand2_1 _20425_ (.Y(_03806_),
    .A(net1720),
    .B(net4668));
 sg13g2_o21ai_1 _20426_ (.B1(_03806_),
    .Y(_01739_),
    .A1(_04427_),
    .A2(net4668));
 sg13g2_nand2_1 _20427_ (.Y(_03807_),
    .A(net1861),
    .B(net4667));
 sg13g2_o21ai_1 _20428_ (.B1(_03807_),
    .Y(_01740_),
    .A1(_04428_),
    .A2(net4667));
 sg13g2_nand2_1 _20429_ (.Y(_03808_),
    .A(net1659),
    .B(net4664));
 sg13g2_o21ai_1 _20430_ (.B1(_03808_),
    .Y(_01741_),
    .A1(_04429_),
    .A2(net4664));
 sg13g2_nand2_1 _20431_ (.Y(_03809_),
    .A(net1331),
    .B(net4658));
 sg13g2_o21ai_1 _20432_ (.B1(_03809_),
    .Y(_01742_),
    .A1(_04430_),
    .A2(net4658));
 sg13g2_nand2_1 _20433_ (.Y(_03810_),
    .A(net1830),
    .B(net4650));
 sg13g2_o21ai_1 _20434_ (.B1(_03810_),
    .Y(_01743_),
    .A1(_04431_),
    .A2(net4650));
 sg13g2_nand2_1 _20435_ (.Y(_03811_),
    .A(net1432),
    .B(net4649));
 sg13g2_o21ai_1 _20436_ (.B1(_03811_),
    .Y(_01744_),
    .A1(_04432_),
    .A2(net4649));
 sg13g2_nand2_1 _20437_ (.Y(_03812_),
    .A(net1693),
    .B(net4623));
 sg13g2_o21ai_1 _20438_ (.B1(_03812_),
    .Y(_01745_),
    .A1(_04433_),
    .A2(net4623));
 sg13g2_nand2_1 _20439_ (.Y(_03813_),
    .A(net1949),
    .B(net4622));
 sg13g2_o21ai_1 _20440_ (.B1(_03813_),
    .Y(_01746_),
    .A1(_04434_),
    .A2(net4622));
 sg13g2_nand2_1 _20441_ (.Y(_03814_),
    .A(net1678),
    .B(net4621));
 sg13g2_o21ai_1 _20442_ (.B1(_03814_),
    .Y(_01747_),
    .A1(_04435_),
    .A2(net4621));
 sg13g2_nand2_1 _20443_ (.Y(_03815_),
    .A(net1562),
    .B(net4613));
 sg13g2_o21ai_1 _20444_ (.B1(_03815_),
    .Y(_01748_),
    .A1(_04436_),
    .A2(net4613));
 sg13g2_nand2_1 _20445_ (.Y(_03816_),
    .A(net1448),
    .B(net4610));
 sg13g2_o21ai_1 _20446_ (.B1(_03816_),
    .Y(_01749_),
    .A1(_04437_),
    .A2(net4610));
 sg13g2_nand2_1 _20447_ (.Y(_03817_),
    .A(net1709),
    .B(net4575));
 sg13g2_o21ai_1 _20448_ (.B1(_03817_),
    .Y(_01750_),
    .A1(_04438_),
    .A2(net4575));
 sg13g2_nand2_1 _20449_ (.Y(_03818_),
    .A(net1791),
    .B(net4577));
 sg13g2_o21ai_1 _20450_ (.B1(_03818_),
    .Y(_01751_),
    .A1(_04439_),
    .A2(net4577));
 sg13g2_nand2_1 _20451_ (.Y(_03819_),
    .A(net1933),
    .B(net4582));
 sg13g2_o21ai_1 _20452_ (.B1(_03819_),
    .Y(_01752_),
    .A1(_04440_),
    .A2(net4582));
 sg13g2_nand2_1 _20453_ (.Y(_03820_),
    .A(net2073),
    .B(net4583));
 sg13g2_o21ai_1 _20454_ (.B1(_03820_),
    .Y(_01753_),
    .A1(_04441_),
    .A2(net4583));
 sg13g2_nand2_1 _20455_ (.Y(_03821_),
    .A(net1975),
    .B(net4585));
 sg13g2_o21ai_1 _20456_ (.B1(_03821_),
    .Y(_01754_),
    .A1(_04442_),
    .A2(net4591));
 sg13g2_nand2_1 _20457_ (.Y(_03822_),
    .A(net1772),
    .B(net4591));
 sg13g2_o21ai_1 _20458_ (.B1(_03822_),
    .Y(_01755_),
    .A1(_04443_),
    .A2(net4591));
 sg13g2_nand2_1 _20459_ (.Y(_03823_),
    .A(net1306),
    .B(net4590));
 sg13g2_o21ai_1 _20460_ (.B1(_03823_),
    .Y(_01756_),
    .A1(_04444_),
    .A2(net4590));
 sg13g2_nand2_1 _20461_ (.Y(_03824_),
    .A(net2062),
    .B(net4594));
 sg13g2_o21ai_1 _20462_ (.B1(_03824_),
    .Y(_01757_),
    .A1(_04445_),
    .A2(net4594));
 sg13g2_nand2_1 _20463_ (.Y(_03825_),
    .A(net1786),
    .B(net4598));
 sg13g2_o21ai_1 _20464_ (.B1(_03825_),
    .Y(_01758_),
    .A1(_04446_),
    .A2(net4598));
 sg13g2_nand2_1 _20465_ (.Y(_03826_),
    .A(net1657),
    .B(net4601));
 sg13g2_o21ai_1 _20466_ (.B1(_03826_),
    .Y(_01759_),
    .A1(_04447_),
    .A2(net4602));
 sg13g2_nand2_1 _20467_ (.Y(_03827_),
    .A(net2208),
    .B(net4602));
 sg13g2_o21ai_1 _20468_ (.B1(_03827_),
    .Y(_01760_),
    .A1(_04448_),
    .A2(net4602));
 sg13g2_nand2_1 _20469_ (.Y(_03828_),
    .A(net1583),
    .B(net4602));
 sg13g2_o21ai_1 _20470_ (.B1(_03828_),
    .Y(_01761_),
    .A1(_04449_),
    .A2(net4605));
 sg13g2_nand2_1 _20471_ (.Y(_03829_),
    .A(net2372),
    .B(net4698));
 sg13g2_o21ai_1 _20472_ (.B1(_03829_),
    .Y(_01762_),
    .A1(_04450_),
    .A2(net4697));
 sg13g2_nand2_1 _20473_ (.Y(_03830_),
    .A(net2041),
    .B(net4706));
 sg13g2_o21ai_1 _20474_ (.B1(_03830_),
    .Y(_01763_),
    .A1(_04451_),
    .A2(net4705));
 sg13g2_nand2_1 _20475_ (.Y(_03831_),
    .A(net2420),
    .B(net4706));
 sg13g2_o21ai_1 _20476_ (.B1(_03831_),
    .Y(_01764_),
    .A1(_04452_),
    .A2(net4706));
 sg13g2_nand2_1 _20477_ (.Y(_03832_),
    .A(net2173),
    .B(net4726));
 sg13g2_o21ai_1 _20478_ (.B1(_03832_),
    .Y(_01765_),
    .A1(_04453_),
    .A2(net4726));
 sg13g2_nand2_1 _20479_ (.Y(_03833_),
    .A(net1872),
    .B(net4727));
 sg13g2_o21ai_1 _20480_ (.B1(_03833_),
    .Y(_01766_),
    .A1(_04454_),
    .A2(net4727));
 sg13g2_nand2_1 _20481_ (.Y(_03834_),
    .A(net1685),
    .B(net4717));
 sg13g2_o21ai_1 _20482_ (.B1(_03834_),
    .Y(_01767_),
    .A1(_04455_),
    .A2(net4715));
 sg13g2_nand2_1 _20483_ (.Y(_03835_),
    .A(net1520),
    .B(net4716));
 sg13g2_o21ai_1 _20484_ (.B1(_03835_),
    .Y(_01768_),
    .A1(_04456_),
    .A2(net4716));
 sg13g2_nand2_1 _20485_ (.Y(_03836_),
    .A(net1247),
    .B(net4712));
 sg13g2_o21ai_1 _20486_ (.B1(_03836_),
    .Y(_01769_),
    .A1(_04457_),
    .A2(net4710));
 sg13g2_nand2_1 _20487_ (.Y(_03837_),
    .A(net1375),
    .B(net4639));
 sg13g2_o21ai_1 _20488_ (.B1(_03837_),
    .Y(_01770_),
    .A1(_04458_),
    .A2(net4639));
 sg13g2_nand2_1 _20489_ (.Y(_03838_),
    .A(net1513),
    .B(net4636));
 sg13g2_o21ai_1 _20490_ (.B1(_03838_),
    .Y(_01771_),
    .A1(_04459_),
    .A2(net4637));
 sg13g2_nand2_1 _20491_ (.Y(_03839_),
    .A(net1430),
    .B(net4664));
 sg13g2_o21ai_1 _20492_ (.B1(_03839_),
    .Y(_01772_),
    .A1(_04460_),
    .A2(net4664));
 sg13g2_nand2_1 _20493_ (.Y(_03840_),
    .A(net1234),
    .B(net4663));
 sg13g2_o21ai_1 _20494_ (.B1(_03840_),
    .Y(_01773_),
    .A1(_04461_),
    .A2(net4663));
 sg13g2_nand2_1 _20495_ (.Y(_03841_),
    .A(net1364),
    .B(net4658));
 sg13g2_o21ai_1 _20496_ (.B1(_03841_),
    .Y(_01774_),
    .A1(_04462_),
    .A2(net4670));
 sg13g2_nand2_1 _20497_ (.Y(_03842_),
    .A(net1465),
    .B(net4651));
 sg13g2_o21ai_1 _20498_ (.B1(_03842_),
    .Y(_01775_),
    .A1(_04463_),
    .A2(net4651));
 sg13g2_nand2_1 _20499_ (.Y(_03843_),
    .A(net1780),
    .B(net4649));
 sg13g2_o21ai_1 _20500_ (.B1(_03843_),
    .Y(_01776_),
    .A1(_04464_),
    .A2(net4652));
 sg13g2_nand2_1 _20501_ (.Y(_03844_),
    .A(net1575),
    .B(net4623));
 sg13g2_o21ai_1 _20502_ (.B1(_03844_),
    .Y(_01777_),
    .A1(_04465_),
    .A2(net4623));
 sg13g2_nand2_1 _20503_ (.Y(_03845_),
    .A(net1945),
    .B(net4622));
 sg13g2_o21ai_1 _20504_ (.B1(_03845_),
    .Y(_01778_),
    .A1(_04466_),
    .A2(net4635));
 sg13g2_nand2_1 _20505_ (.Y(_03846_),
    .A(net1734),
    .B(net4622));
 sg13g2_o21ai_1 _20506_ (.B1(_03846_),
    .Y(_01779_),
    .A1(_04467_),
    .A2(net4622));
 sg13g2_nand2_1 _20507_ (.Y(_03847_),
    .A(net1307),
    .B(net4612));
 sg13g2_o21ai_1 _20508_ (.B1(_03847_),
    .Y(_01780_),
    .A1(_04468_),
    .A2(net4612));
 sg13g2_nand2_1 _20509_ (.Y(_03848_),
    .A(net1404),
    .B(net4610));
 sg13g2_o21ai_1 _20510_ (.B1(_03848_),
    .Y(_01781_),
    .A1(_04469_),
    .A2(net4610));
 sg13g2_nand2_1 _20511_ (.Y(_03849_),
    .A(net1373),
    .B(net4611));
 sg13g2_o21ai_1 _20512_ (.B1(_03849_),
    .Y(_01782_),
    .A1(_04470_),
    .A2(net4611));
 sg13g2_nand2_1 _20513_ (.Y(_03850_),
    .A(net1319),
    .B(net4577));
 sg13g2_o21ai_1 _20514_ (.B1(_03850_),
    .Y(_01783_),
    .A1(_04471_),
    .A2(net4577));
 sg13g2_nand2_1 _20515_ (.Y(_03851_),
    .A(net1894),
    .B(net4578));
 sg13g2_o21ai_1 _20516_ (.B1(_03851_),
    .Y(_01784_),
    .A1(_04472_),
    .A2(net4587));
 sg13g2_nand2_1 _20517_ (.Y(_03852_),
    .A(net2056),
    .B(net4582));
 sg13g2_o21ai_1 _20518_ (.B1(_03852_),
    .Y(_01785_),
    .A1(_04473_),
    .A2(net4582));
 sg13g2_nand2_1 _20519_ (.Y(_03853_),
    .A(net2004),
    .B(net4583));
 sg13g2_o21ai_1 _20520_ (.B1(_03853_),
    .Y(_01786_),
    .A1(_04474_),
    .A2(net4583));
 sg13g2_nand2_1 _20521_ (.Y(_03854_),
    .A(net1267),
    .B(net4589));
 sg13g2_o21ai_1 _20522_ (.B1(_03854_),
    .Y(_01787_),
    .A1(_04475_),
    .A2(net4589));
 sg13g2_nand2_1 _20523_ (.Y(_03855_),
    .A(net2568),
    .B(net4592));
 sg13g2_o21ai_1 _20524_ (.B1(_03855_),
    .Y(_01788_),
    .A1(_04476_),
    .A2(net4592));
 sg13g2_nand2_1 _20525_ (.Y(_03856_),
    .A(net1526),
    .B(net4592));
 sg13g2_o21ai_1 _20526_ (.B1(_03856_),
    .Y(_01789_),
    .A1(_04477_),
    .A2(net4591));
 sg13g2_nand2_1 _20527_ (.Y(_03857_),
    .A(net1587),
    .B(net4595));
 sg13g2_o21ai_1 _20528_ (.B1(_03857_),
    .Y(_01790_),
    .A1(_04478_),
    .A2(net4595));
 sg13g2_nand2_1 _20529_ (.Y(_03858_),
    .A(net1603),
    .B(net4599));
 sg13g2_o21ai_1 _20530_ (.B1(_03858_),
    .Y(_01791_),
    .A1(_04479_),
    .A2(net4599));
 sg13g2_nand2_1 _20531_ (.Y(_03859_),
    .A(net1327),
    .B(net4691));
 sg13g2_o21ai_1 _20532_ (.B1(_03859_),
    .Y(_01792_),
    .A1(_04480_),
    .A2(net4691));
 sg13g2_nand2_1 _20533_ (.Y(_03860_),
    .A(net1893),
    .B(net4691));
 sg13g2_o21ai_1 _20534_ (.B1(_03860_),
    .Y(_01793_),
    .A1(_04481_),
    .A2(net4691));
 sg13g2_nand2_1 _20535_ (.Y(_03861_),
    .A(net2012),
    .B(net4693));
 sg13g2_o21ai_1 _20536_ (.B1(_03861_),
    .Y(_01794_),
    .A1(_04482_),
    .A2(net4693));
 sg13g2_nand2_1 _20537_ (.Y(_03862_),
    .A(net1707),
    .B(net4700));
 sg13g2_o21ai_1 _20538_ (.B1(_03862_),
    .Y(_01795_),
    .A1(_04483_),
    .A2(net4700));
 sg13g2_nand2_1 _20539_ (.Y(_03863_),
    .A(net1516),
    .B(net4702));
 sg13g2_o21ai_1 _20540_ (.B1(_03863_),
    .Y(_01796_),
    .A1(_04484_),
    .A2(net4702));
 sg13g2_nand2_1 _20541_ (.Y(_03864_),
    .A(net1610),
    .B(net4722));
 sg13g2_o21ai_1 _20542_ (.B1(_03864_),
    .Y(_01797_),
    .A1(_04485_),
    .A2(net4723));
 sg13g2_nand2_1 _20543_ (.Y(_03865_),
    .A(net1689),
    .B(net4722));
 sg13g2_o21ai_1 _20544_ (.B1(_03865_),
    .Y(_01798_),
    .A1(_04486_),
    .A2(net4722));
 sg13g2_nand2_1 _20545_ (.Y(_03866_),
    .A(net1849),
    .B(net4714));
 sg13g2_o21ai_1 _20546_ (.B1(_03866_),
    .Y(_01799_),
    .A1(_04487_),
    .A2(net4714));
 sg13g2_nand2_1 _20547_ (.Y(_03867_),
    .A(net1422),
    .B(net4684));
 sg13g2_o21ai_1 _20548_ (.B1(_03867_),
    .Y(_01800_),
    .A1(_04488_),
    .A2(net4684));
 sg13g2_nand2_1 _20549_ (.Y(_03868_),
    .A(net1996),
    .B(net4683));
 sg13g2_o21ai_1 _20550_ (.B1(_03868_),
    .Y(_01801_),
    .A1(_04489_),
    .A2(net4683));
 sg13g2_nand2_1 _20551_ (.Y(_03869_),
    .A(net2090),
    .B(net4642));
 sg13g2_o21ai_1 _20552_ (.B1(_03869_),
    .Y(_01802_),
    .A1(_04490_),
    .A2(net4640));
 sg13g2_nand2_1 _20553_ (.Y(_03870_),
    .A(net1712),
    .B(net4636));
 sg13g2_o21ai_1 _20554_ (.B1(_03870_),
    .Y(_01803_),
    .A1(_04491_),
    .A2(net4636));
 sg13g2_nand2_1 _20555_ (.Y(_03871_),
    .A(\TRNG.Padded_Out[176] ),
    .B(net4661));
 sg13g2_o21ai_1 _20556_ (.B1(_03871_),
    .Y(_01804_),
    .A1(_04492_),
    .A2(net4662));
 sg13g2_nand2_1 _20557_ (.Y(_03872_),
    .A(net1238),
    .B(net4663));
 sg13g2_o21ai_1 _20558_ (.B1(_03872_),
    .Y(_01805_),
    .A1(_04493_),
    .A2(net4663));
 sg13g2_nand2_1 _20559_ (.Y(_03873_),
    .A(net2110),
    .B(net4650));
 sg13g2_o21ai_1 _20560_ (.B1(_03873_),
    .Y(_01806_),
    .A1(_04494_),
    .A2(net4650));
 sg13g2_nand2_1 _20561_ (.Y(_03874_),
    .A(net1545),
    .B(net4650));
 sg13g2_o21ai_1 _20562_ (.B1(_03874_),
    .Y(_01807_),
    .A1(_04495_),
    .A2(net4650));
 sg13g2_nand2_1 _20563_ (.Y(_03875_),
    .A(net1261),
    .B(net4649));
 sg13g2_o21ai_1 _20564_ (.B1(_03875_),
    .Y(_01808_),
    .A1(_04496_),
    .A2(net4652));
 sg13g2_nand2_1 _20565_ (.Y(_03876_),
    .A(net1491),
    .B(net4624));
 sg13g2_o21ai_1 _20566_ (.B1(_03876_),
    .Y(_01809_),
    .A1(_04497_),
    .A2(net4624));
 sg13g2_nand2_1 _20567_ (.Y(_03877_),
    .A(net1670),
    .B(net4623));
 sg13g2_o21ai_1 _20568_ (.B1(_03877_),
    .Y(_01810_),
    .A1(_04498_),
    .A2(net4621));
 sg13g2_nand2_1 _20569_ (.Y(_03878_),
    .A(net1808),
    .B(net4607));
 sg13g2_o21ai_1 _20570_ (.B1(_03878_),
    .Y(_01811_),
    .A1(_04499_),
    .A2(net4607));
 sg13g2_nand2_1 _20571_ (.Y(_03879_),
    .A(net1395),
    .B(net4612));
 sg13g2_o21ai_1 _20572_ (.B1(_03879_),
    .Y(_01812_),
    .A1(_04500_),
    .A2(net4612));
 sg13g2_nand2_1 _20573_ (.Y(_03880_),
    .A(net1270),
    .B(net4571));
 sg13g2_o21ai_1 _20574_ (.B1(_03880_),
    .Y(_01813_),
    .A1(_04501_),
    .A2(net4571));
 sg13g2_nand2_1 _20575_ (.Y(_03881_),
    .A(\TRNG.Padded_Out[186] ),
    .B(net4574));
 sg13g2_o21ai_1 _20576_ (.B1(_03881_),
    .Y(_01814_),
    .A1(_04502_),
    .A2(net4574));
 sg13g2_nand2_1 _20577_ (.Y(_03882_),
    .A(net2048),
    .B(net4573));
 sg13g2_o21ai_1 _20578_ (.B1(_03882_),
    .Y(_01815_),
    .A1(_04503_),
    .A2(net4588));
 sg13g2_nand2_1 _20579_ (.Y(_03883_),
    .A(net1870),
    .B(net4578));
 sg13g2_o21ai_1 _20580_ (.B1(_03883_),
    .Y(_01816_),
    .A1(_04504_),
    .A2(net4587));
 sg13g2_nand2_1 _20581_ (.Y(_03884_),
    .A(net1510),
    .B(net4582));
 sg13g2_o21ai_1 _20582_ (.B1(_03884_),
    .Y(_01817_),
    .A1(_04505_),
    .A2(net4587));
 sg13g2_nand2_1 _20583_ (.Y(_03885_),
    .A(net3119),
    .B(net4587));
 sg13g2_o21ai_1 _20584_ (.B1(_03885_),
    .Y(_01818_),
    .A1(_04506_),
    .A2(net4587));
 sg13g2_nand2_1 _20585_ (.Y(_03886_),
    .A(net2079),
    .B(net4589));
 sg13g2_o21ai_1 _20586_ (.B1(_03886_),
    .Y(_01819_),
    .A1(_04507_),
    .A2(net4597));
 sg13g2_nand2_1 _20587_ (.Y(_03887_),
    .A(net1890),
    .B(net4590));
 sg13g2_o21ai_1 _20588_ (.B1(_03887_),
    .Y(_01820_),
    .A1(_04508_),
    .A2(net4590));
 sg13g2_nand2_1 _20589_ (.Y(_03888_),
    .A(net2430),
    .B(net4595));
 sg13g2_o21ai_1 _20590_ (.B1(_03888_),
    .Y(_01821_),
    .A1(_04509_),
    .A2(net4594));
 sg13g2_nand2_1 _20591_ (.Y(_03889_),
    .A(net1793),
    .B(net4595));
 sg13g2_o21ai_1 _20592_ (.B1(_03889_),
    .Y(_01822_),
    .A1(_04510_),
    .A2(net4596));
 sg13g2_nand2_1 _20593_ (.Y(_03890_),
    .A(net1483),
    .B(net4598));
 sg13g2_o21ai_1 _20594_ (.B1(_03890_),
    .Y(_01823_),
    .A1(_04511_),
    .A2(net4598));
 sg13g2_nand2_1 _20595_ (.Y(_03891_),
    .A(net1842),
    .B(net4603));
 sg13g2_o21ai_1 _20596_ (.B1(_03891_),
    .Y(_01824_),
    .A1(_04512_),
    .A2(net4603));
 sg13g2_nand2_1 _20597_ (.Y(_03892_),
    .A(net1414),
    .B(net4603));
 sg13g2_o21ai_1 _20598_ (.B1(_03892_),
    .Y(_01825_),
    .A1(_04513_),
    .A2(net4603));
 sg13g2_nand2_1 _20599_ (.Y(_03893_),
    .A(net1460),
    .B(net4694));
 sg13g2_o21ai_1 _20600_ (.B1(_03893_),
    .Y(_01826_),
    .A1(_04514_),
    .A2(net4693));
 sg13g2_nand2_1 _20601_ (.Y(_03894_),
    .A(net1672),
    .B(net4700));
 sg13g2_o21ai_1 _20602_ (.B1(_03894_),
    .Y(_01827_),
    .A1(_04515_),
    .A2(net4700));
 sg13g2_nand2_1 _20603_ (.Y(_03895_),
    .A(net1475),
    .B(net4702));
 sg13g2_o21ai_1 _20604_ (.B1(_03895_),
    .Y(_01828_),
    .A1(_04516_),
    .A2(net4702));
 sg13g2_nand2_1 _20605_ (.Y(_03896_),
    .A(net1834),
    .B(net4701));
 sg13g2_o21ai_1 _20606_ (.B1(_03896_),
    .Y(_01829_),
    .A1(_04517_),
    .A2(net4701));
 sg13g2_nand2_1 _20607_ (.Y(_03897_),
    .A(net1408),
    .B(net4688));
 sg13g2_o21ai_1 _20608_ (.B1(_03897_),
    .Y(_01830_),
    .A1(_04518_),
    .A2(net4688));
 sg13g2_nand2_1 _20609_ (.Y(_03898_),
    .A(net2040),
    .B(net4714));
 sg13g2_o21ai_1 _20610_ (.B1(_03898_),
    .Y(_01831_),
    .A1(_04519_),
    .A2(net4688));
 sg13g2_nand2_1 _20611_ (.Y(_03899_),
    .A(net1479),
    .B(net4711));
 sg13g2_o21ai_1 _20612_ (.B1(_03899_),
    .Y(_01832_),
    .A1(_04520_),
    .A2(net4714));
 sg13g2_nand2_1 _20613_ (.Y(_03900_),
    .A(net1939),
    .B(net4711));
 sg13g2_o21ai_1 _20614_ (.B1(_03900_),
    .Y(_01833_),
    .A1(_04521_),
    .A2(net4711));
 sg13g2_nand2_1 _20615_ (.Y(_03901_),
    .A(net1826),
    .B(net4710));
 sg13g2_o21ai_1 _20616_ (.B1(_03901_),
    .Y(_01834_),
    .A1(_04522_),
    .A2(net4710));
 sg13g2_nand2_1 _20617_ (.Y(_03902_),
    .A(net1621),
    .B(net4666));
 sg13g2_o21ai_1 _20618_ (.B1(_03902_),
    .Y(_01835_),
    .A1(_04523_),
    .A2(net4666));
 sg13g2_nand2_1 _20619_ (.Y(_03903_),
    .A(net1743),
    .B(net4668));
 sg13g2_o21ai_1 _20620_ (.B1(_03903_),
    .Y(_01836_),
    .A1(_04524_),
    .A2(net4667));
 sg13g2_nand2_1 _20621_ (.Y(_03904_),
    .A(net2052),
    .B(net4670));
 sg13g2_o21ai_1 _20622_ (.B1(_03904_),
    .Y(_01837_),
    .A1(_04525_),
    .A2(net4670));
 sg13g2_nand2_1 _20623_ (.Y(_03905_),
    .A(net1767),
    .B(net4658));
 sg13g2_o21ai_1 _20624_ (.B1(_03905_),
    .Y(_01838_),
    .A1(_04526_),
    .A2(net4658));
 sg13g2_nand2_1 _20625_ (.Y(_03906_),
    .A(net2337),
    .B(net4658));
 sg13g2_o21ai_1 _20626_ (.B1(_03906_),
    .Y(_01839_),
    .A1(_04527_),
    .A2(net4658));
 sg13g2_nand2_1 _20627_ (.Y(_03907_),
    .A(net1755),
    .B(net4649));
 sg13g2_o21ai_1 _20628_ (.B1(_03907_),
    .Y(_01840_),
    .A1(_04528_),
    .A2(net4649));
 sg13g2_nand2_1 _20629_ (.Y(_03908_),
    .A(net1313),
    .B(net4623));
 sg13g2_o21ai_1 _20630_ (.B1(_03908_),
    .Y(_01841_),
    .A1(_04529_),
    .A2(net4623));
 sg13g2_nand2_1 _20631_ (.Y(_03909_),
    .A(net1711),
    .B(net4637));
 sg13g2_o21ai_1 _20632_ (.B1(_03909_),
    .Y(_01842_),
    .A1(_04530_),
    .A2(net4635));
 sg13g2_nand2_1 _20633_ (.Y(_03910_),
    .A(net1965),
    .B(net4635));
 sg13g2_o21ai_1 _20634_ (.B1(_03910_),
    .Y(_01843_),
    .A1(_04531_),
    .A2(net4635));
 sg13g2_nand2_1 _20635_ (.Y(_03911_),
    .A(net2263),
    .B(net4629));
 sg13g2_o21ai_1 _20636_ (.B1(_03911_),
    .Y(_01844_),
    .A1(_04532_),
    .A2(net4629));
 sg13g2_nand2_1 _20637_ (.Y(_03912_),
    .A(net2190),
    .B(net4629));
 sg13g2_o21ai_1 _20638_ (.B1(_03912_),
    .Y(_01845_),
    .A1(_04533_),
    .A2(net4629));
 sg13g2_nand2_1 _20639_ (.Y(_03913_),
    .A(net1765),
    .B(net4627));
 sg13g2_o21ai_1 _20640_ (.B1(_03913_),
    .Y(_01846_),
    .A1(_04534_),
    .A2(net4627));
 sg13g2_nand2_1 _20641_ (.Y(_03914_),
    .A(net1214),
    .B(net4579));
 sg13g2_o21ai_1 _20642_ (.B1(_03914_),
    .Y(_01847_),
    .A1(_04535_),
    .A2(net4579));
 sg13g2_nand2_1 _20643_ (.Y(_03915_),
    .A(net1458),
    .B(net4577));
 sg13g2_o21ai_1 _20644_ (.B1(_03915_),
    .Y(_01848_),
    .A1(_04536_),
    .A2(net4578));
 sg13g2_nand2_1 _20645_ (.Y(_03916_),
    .A(net2007),
    .B(net4583));
 sg13g2_o21ai_1 _20646_ (.B1(_03916_),
    .Y(_01849_),
    .A1(_04537_),
    .A2(net4583));
 sg13g2_nand2_1 _20647_ (.Y(_03917_),
    .A(net2598),
    .B(net4589));
 sg13g2_o21ai_1 _20648_ (.B1(_03917_),
    .Y(_01850_),
    .A1(_04538_),
    .A2(net4589));
 sg13g2_nand2_1 _20649_ (.Y(_03918_),
    .A(net2144),
    .B(net4589));
 sg13g2_o21ai_1 _20650_ (.B1(_03918_),
    .Y(_01851_),
    .A1(_04539_),
    .A2(net4597));
 sg13g2_nand2_1 _20651_ (.Y(_03919_),
    .A(net2092),
    .B(net4590));
 sg13g2_o21ai_1 _20652_ (.B1(_03919_),
    .Y(_01852_),
    .A1(_04540_),
    .A2(net4597));
 sg13g2_nand2_1 _20653_ (.Y(_03920_),
    .A(net1739),
    .B(net4594));
 sg13g2_o21ai_1 _20654_ (.B1(_03920_),
    .Y(_01853_),
    .A1(_04541_),
    .A2(net4594));
 sg13g2_nand2_1 _20655_ (.Y(_03921_),
    .A(net1726),
    .B(net4593));
 sg13g2_o21ai_1 _20656_ (.B1(_03921_),
    .Y(_01854_),
    .A1(_04542_),
    .A2(net4598));
 sg13g2_nand2_1 _20657_ (.Y(_03922_),
    .A(net2180),
    .B(net4598));
 sg13g2_o21ai_1 _20658_ (.B1(_03922_),
    .Y(_01855_),
    .A1(_04543_),
    .A2(net4598));
 sg13g2_nand2_1 _20659_ (.Y(_03923_),
    .A(net2009),
    .B(net4602));
 sg13g2_o21ai_1 _20660_ (.B1(_03923_),
    .Y(_01856_),
    .A1(_04544_),
    .A2(net4602));
 sg13g2_nand2_1 _20661_ (.Y(_03924_),
    .A(net2258),
    .B(net4604));
 sg13g2_o21ai_1 _20662_ (.B1(_03924_),
    .Y(_01857_),
    .A1(_04545_),
    .A2(net4602));
 sg13g2_nand2_1 _20663_ (.Y(_03925_),
    .A(net2028),
    .B(net4697));
 sg13g2_o21ai_1 _20664_ (.B1(_03925_),
    .Y(_01858_),
    .A1(_04546_),
    .A2(net4697));
 sg13g2_nand2_1 _20665_ (.Y(_03926_),
    .A(net1652),
    .B(net4705));
 sg13g2_o21ai_1 _20666_ (.B1(_03926_),
    .Y(_01859_),
    .A1(_04547_),
    .A2(net4705));
 sg13g2_nand2_1 _20667_ (.Y(_03927_),
    .A(net1485),
    .B(net4707));
 sg13g2_o21ai_1 _20668_ (.B1(_03927_),
    .Y(_01860_),
    .A1(_04548_),
    .A2(net4707));
 sg13g2_nand2_1 _20669_ (.Y(_03928_),
    .A(net1454),
    .B(net4701));
 sg13g2_o21ai_1 _20670_ (.B1(_03928_),
    .Y(_01861_),
    .A1(_04549_),
    .A2(net4701));
 sg13g2_nand2_1 _20671_ (.Y(_03929_),
    .A(net1467),
    .B(net4688));
 sg13g2_o21ai_1 _20672_ (.B1(_03929_),
    .Y(_01862_),
    .A1(_04550_),
    .A2(net4688));
 sg13g2_nand2_1 _20673_ (.Y(_03930_),
    .A(net1339),
    .B(net4688));
 sg13g2_o21ai_1 _20674_ (.B1(_03930_),
    .Y(_01863_),
    .A1(_04551_),
    .A2(net4688));
 sg13g2_nand2_1 _20675_ (.Y(_03931_),
    .A(net1655),
    .B(net4684));
 sg13g2_o21ai_1 _20676_ (.B1(_03931_),
    .Y(_01864_),
    .A1(_04552_),
    .A2(net4684));
 sg13g2_nand2_1 _20677_ (.Y(_03932_),
    .A(net1784),
    .B(net4684));
 sg13g2_o21ai_1 _20678_ (.B1(_03932_),
    .Y(_01865_),
    .A1(_04553_),
    .A2(net4684));
 sg13g2_nand2_1 _20679_ (.Y(_03933_),
    .A(net2036),
    .B(net4641));
 sg13g2_o21ai_1 _20680_ (.B1(_03933_),
    .Y(_01866_),
    .A1(_04554_),
    .A2(net4641));
 sg13g2_nand2_1 _20681_ (.Y(_03934_),
    .A(net1437),
    .B(net4666));
 sg13g2_o21ai_1 _20682_ (.B1(_03934_),
    .Y(_01867_),
    .A1(_04555_),
    .A2(net4666));
 sg13g2_nand2_1 _20683_ (.Y(_03935_),
    .A(net2021),
    .B(net4667));
 sg13g2_o21ai_1 _20684_ (.B1(_03935_),
    .Y(_01868_),
    .A1(_04556_),
    .A2(net4667));
 sg13g2_nand2_1 _20685_ (.Y(_03936_),
    .A(net1840),
    .B(net4670));
 sg13g2_o21ai_1 _20686_ (.B1(_03936_),
    .Y(_01869_),
    .A1(_04557_),
    .A2(net4670));
 sg13g2_nand2_1 _20687_ (.Y(_03937_),
    .A(net2257),
    .B(net4653));
 sg13g2_o21ai_1 _20688_ (.B1(_03937_),
    .Y(_01870_),
    .A1(_04558_),
    .A2(net4653));
 sg13g2_nand2_1 _20689_ (.Y(_03938_),
    .A(net1667),
    .B(net4654));
 sg13g2_o21ai_1 _20690_ (.B1(_03938_),
    .Y(_01871_),
    .A1(_04559_),
    .A2(net4654));
 sg13g2_nand2_1 _20691_ (.Y(_03939_),
    .A(net2221),
    .B(net4644));
 sg13g2_o21ai_1 _20692_ (.B1(_03939_),
    .Y(_01872_),
    .A1(_04560_),
    .A2(net4644));
 sg13g2_nand2_1 _20693_ (.Y(_03940_),
    .A(net1446),
    .B(net4619));
 sg13g2_o21ai_1 _20694_ (.B1(_03940_),
    .Y(_01873_),
    .A1(_04561_),
    .A2(net4619));
 sg13g2_nand2_1 _20695_ (.Y(_03941_),
    .A(net1716),
    .B(net4617));
 sg13g2_o21ai_1 _20696_ (.B1(_03941_),
    .Y(_01874_),
    .A1(_04562_),
    .A2(net4617));
 sg13g2_nand2_1 _20697_ (.Y(_03942_),
    .A(net1914),
    .B(net4617));
 sg13g2_o21ai_1 _20698_ (.B1(_03942_),
    .Y(_01875_),
    .A1(_04563_),
    .A2(net4617));
 sg13g2_nand2_1 _20699_ (.Y(_03943_),
    .A(net1284),
    .B(net4612));
 sg13g2_o21ai_1 _20700_ (.B1(_03943_),
    .Y(_01876_),
    .A1(_04564_),
    .A2(net4612));
 sg13g2_nand2_1 _20701_ (.Y(_03944_),
    .A(net1274),
    .B(net4611));
 sg13g2_o21ai_1 _20702_ (.B1(_03944_),
    .Y(_01877_),
    .A1(_04565_),
    .A2(net4611));
 sg13g2_nand2_1 _20703_ (.Y(_03945_),
    .A(net1877),
    .B(net4627));
 sg13g2_o21ai_1 _20704_ (.B1(_03945_),
    .Y(_01878_),
    .A1(_04566_),
    .A2(net4627));
 sg13g2_nand2_1 _20705_ (.Y(_03946_),
    .A(net1802),
    .B(net4627));
 sg13g2_o21ai_1 _20706_ (.B1(_03946_),
    .Y(_01879_),
    .A1(_04567_),
    .A2(net4627));
 sg13g2_nand2_1 _20707_ (.Y(_03947_),
    .A(net1416),
    .B(net4579));
 sg13g2_o21ai_1 _20708_ (.B1(_03947_),
    .Y(_01880_),
    .A1(_04568_),
    .A2(net4579));
 sg13g2_nand2_1 _20709_ (.Y(_03948_),
    .A(net1683),
    .B(net4631));
 sg13g2_o21ai_1 _20710_ (.B1(_03948_),
    .Y(_01881_),
    .A1(_04569_),
    .A2(net4631));
 sg13g2_nand2_1 _20711_ (.Y(_03949_),
    .A(net2023),
    .B(net4632));
 sg13g2_o21ai_1 _20712_ (.B1(_03949_),
    .Y(_01882_),
    .A1(_04570_),
    .A2(net4632));
 sg13g2_nand2_1 _20713_ (.Y(_03950_),
    .A(net2000),
    .B(net4675));
 sg13g2_o21ai_1 _20714_ (.B1(_03950_),
    .Y(_01883_),
    .A1(_04571_),
    .A2(net4675));
 sg13g2_nand2_1 _20715_ (.Y(_03951_),
    .A(net1302),
    .B(net4676));
 sg13g2_o21ai_1 _20716_ (.B1(_03951_),
    .Y(_01884_),
    .A1(_04572_),
    .A2(net4676));
 sg13g2_nand2_1 _20717_ (.Y(_03952_),
    .A(net1495),
    .B(net4679));
 sg13g2_o21ai_1 _20718_ (.B1(_03952_),
    .Y(_01885_),
    .A1(_04573_),
    .A2(net4680));
 sg13g2_nand2_1 _20719_ (.Y(_03953_),
    .A(net1843),
    .B(net4595));
 sg13g2_o21ai_1 _20720_ (.B1(_03953_),
    .Y(_01886_),
    .A1(_04574_),
    .A2(net4596));
 sg13g2_nand2_1 _20721_ (.Y(_03954_),
    .A(net1294),
    .B(net4599));
 sg13g2_o21ai_1 _20722_ (.B1(_03954_),
    .Y(_01887_),
    .A1(_04575_),
    .A2(net4599));
 sg13g2_nand2_1 _20723_ (.Y(_03955_),
    .A(net1701),
    .B(net4603));
 sg13g2_o21ai_1 _20724_ (.B1(_03955_),
    .Y(_01888_),
    .A1(_04576_),
    .A2(net4603));
 sg13g2_nand2_1 _20725_ (.Y(_03956_),
    .A(net1555),
    .B(net4695));
 sg13g2_o21ai_1 _20726_ (.B1(_03956_),
    .Y(_01889_),
    .A1(_04577_),
    .A2(net4603));
 sg13g2_nand2_1 _20727_ (.Y(_03957_),
    .A(net2412),
    .B(net4693));
 sg13g2_o21ai_1 _20728_ (.B1(_03957_),
    .Y(_01890_),
    .A1(_04578_),
    .A2(net4698));
 sg13g2_nand2_1 _20729_ (.Y(_03958_),
    .A(net1278),
    .B(net4705));
 sg13g2_o21ai_1 _20730_ (.B1(_03958_),
    .Y(_01891_),
    .A1(_04579_),
    .A2(net4704));
 sg13g2_nand2_1 _20731_ (.Y(_03959_),
    .A(net1452),
    .B(net4702));
 sg13g2_o21ai_1 _20732_ (.B1(_03959_),
    .Y(_01892_),
    .A1(_04580_),
    .A2(net4701));
 sg13g2_nand2_1 _20733_ (.Y(_03960_),
    .A(net1249),
    .B(net4723));
 sg13g2_o21ai_1 _20734_ (.B1(_03960_),
    .Y(_01893_),
    .A1(_04581_),
    .A2(net4723));
 sg13g2_nand2_1 _20735_ (.Y(_03961_),
    .A(net1969),
    .B(net4725));
 sg13g2_o21ai_1 _20736_ (.B1(_03961_),
    .Y(_01894_),
    .A1(_04582_),
    .A2(net4722));
 sg13g2_nand2_1 _20737_ (.Y(_03962_),
    .A(net1810),
    .B(net4714));
 sg13g2_o21ai_1 _20738_ (.B1(_03962_),
    .Y(_01895_),
    .A1(_04583_),
    .A2(net4714));
 sg13g2_nand2_1 _20739_ (.Y(_03963_),
    .A(net1571),
    .B(net4683));
 sg13g2_o21ai_1 _20740_ (.B1(_03963_),
    .Y(_01896_),
    .A1(_04584_),
    .A2(net4683));
 sg13g2_nand2_1 _20741_ (.Y(_03964_),
    .A(net2155),
    .B(net4640));
 sg13g2_o21ai_1 _20742_ (.B1(_03964_),
    .Y(_01897_),
    .A1(_04585_),
    .A2(net4640));
 sg13g2_nand2_1 _20743_ (.Y(_03965_),
    .A(net1530),
    .B(net4639));
 sg13g2_o21ai_1 _20744_ (.B1(_03965_),
    .Y(_01898_),
    .A1(_04586_),
    .A2(net4639));
 sg13g2_nand2_1 _20745_ (.Y(_03966_),
    .A(net1859),
    .B(net4637));
 sg13g2_o21ai_1 _20746_ (.B1(_03966_),
    .Y(_01899_),
    .A1(_04587_),
    .A2(net4636));
 sg13g2_nand2_1 _20747_ (.Y(_03967_),
    .A(net1618),
    .B(net4661));
 sg13g2_o21ai_1 _20748_ (.B1(_03967_),
    .Y(_01900_),
    .A1(_04588_),
    .A2(net4661));
 sg13g2_nand2_1 _20749_ (.Y(_03968_),
    .A(net1614),
    .B(net4657));
 sg13g2_o21ai_1 _20750_ (.B1(_03968_),
    .Y(_01901_),
    .A1(_04589_),
    .A2(net4651));
 sg13g2_nand2_1 _20751_ (.Y(_03969_),
    .A(net1705),
    .B(net4654));
 sg13g2_o21ai_1 _20752_ (.B1(_03969_),
    .Y(_01902_),
    .A1(_04590_),
    .A2(net4657));
 sg13g2_nand2_1 _20753_ (.Y(_03970_),
    .A(net1263),
    .B(net4650));
 sg13g2_o21ai_1 _20754_ (.B1(_03970_),
    .Y(_01903_),
    .A1(_04591_),
    .A2(net4650));
 sg13g2_nand2_1 _20755_ (.Y(_03971_),
    .A(net1369),
    .B(net4649));
 sg13g2_o21ai_1 _20756_ (.B1(_03971_),
    .Y(_01904_),
    .A1(_04592_),
    .A2(net4649));
 sg13g2_nand2_1 _20757_ (.Y(_03972_),
    .A(net1383),
    .B(net4624));
 sg13g2_o21ai_1 _20758_ (.B1(_03972_),
    .Y(_01905_),
    .A1(_04593_),
    .A2(net4624));
 sg13g2_nand2_1 _20759_ (.Y(_03973_),
    .A(net1377),
    .B(net4635));
 sg13g2_o21ai_1 _20760_ (.B1(_03973_),
    .Y(_01906_),
    .A1(_04594_),
    .A2(net4635));
 sg13g2_nand2_1 _20761_ (.Y(_03974_),
    .A(net1631),
    .B(net4638));
 sg13g2_o21ai_1 _20762_ (.B1(_03974_),
    .Y(_01907_),
    .A1(_04595_),
    .A2(net4638));
 sg13g2_nand2_1 _20763_ (.Y(_03975_),
    .A(net1391),
    .B(net4629));
 sg13g2_o21ai_1 _20764_ (.B1(_03975_),
    .Y(_01908_),
    .A1(_04596_),
    .A2(net4629));
 sg13g2_nand2_1 _20765_ (.Y(_03976_),
    .A(net2341),
    .B(net4629));
 sg13g2_o21ai_1 _20766_ (.B1(_03976_),
    .Y(_01909_),
    .A1(_04597_),
    .A2(net4629));
 sg13g2_nand2_1 _20767_ (.Y(_03977_),
    .A(net1898),
    .B(net4627));
 sg13g2_o21ai_1 _20768_ (.B1(_03977_),
    .Y(_01910_),
    .A1(_04598_),
    .A2(net4628));
 sg13g2_nand2_1 _20769_ (.Y(_03978_),
    .A(net2138),
    .B(net4627));
 sg13g2_o21ai_1 _20770_ (.B1(_03978_),
    .Y(_01911_),
    .A1(_04599_),
    .A2(net4628));
 sg13g2_nand2_1 _20771_ (.Y(_03979_),
    .A(net1737),
    .B(net4584));
 sg13g2_o21ai_1 _20772_ (.B1(_03979_),
    .Y(_01912_),
    .A1(_04600_),
    .A2(net4584));
 sg13g2_nand2_1 _20773_ (.Y(_03980_),
    .A(net1344),
    .B(net4631));
 sg13g2_o21ai_1 _20774_ (.B1(_03980_),
    .Y(_01913_),
    .A1(_04601_),
    .A2(net4631));
 sg13g2_nand2_1 _20775_ (.Y(_03981_),
    .A(net1906),
    .B(net4631));
 sg13g2_o21ai_1 _20776_ (.B1(_03981_),
    .Y(_01914_),
    .A1(_04602_),
    .A2(net4631));
 sg13g2_nand2_1 _20777_ (.Y(_03982_),
    .A(net1498),
    .B(net4677));
 sg13g2_o21ai_1 _20778_ (.B1(_03982_),
    .Y(_01915_),
    .A1(_04603_),
    .A2(net4677));
 sg13g2_nand2_1 _20779_ (.Y(_03983_),
    .A(net2145),
    .B(net4677));
 sg13g2_o21ai_1 _20780_ (.B1(_03983_),
    .Y(_01916_),
    .A1(_04604_),
    .A2(net4678));
 sg13g2_nand2_1 _20781_ (.Y(_03984_),
    .A(net1620),
    .B(net4681));
 sg13g2_o21ai_1 _20782_ (.B1(_03984_),
    .Y(_01917_),
    .A1(_04605_),
    .A2(net4681));
 sg13g2_nand2_1 _20783_ (.Y(_03985_),
    .A(net1728),
    .B(net4595));
 sg13g2_o21ai_1 _20784_ (.B1(_03985_),
    .Y(_01918_),
    .A1(_04606_),
    .A2(net4595));
 sg13g2_nand2_1 _20785_ (.Y(_03986_),
    .A(net1800),
    .B(net4600));
 sg13g2_o21ai_1 _20786_ (.B1(_03986_),
    .Y(_01919_),
    .A1(_04607_),
    .A2(net4600));
 sg13g2_nand2_1 _20787_ (.Y(_03987_),
    .A(net2543),
    .B(net4696));
 sg13g2_o21ai_1 _20788_ (.B1(_03987_),
    .Y(_01920_),
    .A1(_04608_),
    .A2(net4699));
 sg13g2_nand2_1 _20789_ (.Y(_03988_),
    .A(net1876),
    .B(net4696));
 sg13g2_o21ai_1 _20790_ (.B1(_03988_),
    .Y(_01921_),
    .A1(_04609_),
    .A2(net4696));
 sg13g2_nand2_1 _20791_ (.Y(_03989_),
    .A(net1645),
    .B(net4697));
 sg13g2_o21ai_1 _20792_ (.B1(_03989_),
    .Y(_01922_),
    .A1(_04610_),
    .A2(net4698));
 sg13g2_nand2_1 _20793_ (.Y(_03990_),
    .A(net2633),
    .B(net4704));
 sg13g2_o21ai_1 _20794_ (.B1(_03990_),
    .Y(_01923_),
    .A1(_04611_),
    .A2(net4705));
 sg13g2_nand2_1 _20795_ (.Y(_03991_),
    .A(net2264),
    .B(net4726));
 sg13g2_o21ai_1 _20796_ (.B1(_03991_),
    .Y(_01924_),
    .A1(_04612_),
    .A2(net4726));
 sg13g2_nand2_1 _20797_ (.Y(_03992_),
    .A(net2718),
    .B(net4728));
 sg13g2_o21ai_1 _20798_ (.B1(_03992_),
    .Y(_01925_),
    .A1(_04613_),
    .A2(net4728));
 sg13g2_nand2_1 _20799_ (.Y(_03993_),
    .A(net2126),
    .B(net4727));
 sg13g2_o21ai_1 _20800_ (.B1(_03993_),
    .Y(_01926_),
    .A1(_04614_),
    .A2(net4727));
 sg13g2_nand2_1 _20801_ (.Y(_03994_),
    .A(net1691),
    .B(net4724));
 sg13g2_o21ai_1 _20802_ (.B1(_03994_),
    .Y(_01927_),
    .A1(_04615_),
    .A2(net4724));
 sg13g2_nand2_1 _20803_ (.Y(_03995_),
    .A(net1778),
    .B(net4716));
 sg13g2_o21ai_1 _20804_ (.B1(_03995_),
    .Y(_01928_),
    .A1(_04616_),
    .A2(net4716));
 sg13g2_nand2_1 _20805_ (.Y(_03996_),
    .A(net1435),
    .B(net4712));
 sg13g2_o21ai_1 _20806_ (.B1(_03996_),
    .Y(_01929_),
    .A1(_04617_),
    .A2(net4712));
 sg13g2_nand2_1 _20807_ (.Y(_03997_),
    .A(net1855),
    .B(net4712));
 sg13g2_o21ai_1 _20808_ (.B1(_03997_),
    .Y(_01930_),
    .A1(_04618_),
    .A2(net4712));
 sg13g2_nand2_1 _20809_ (.Y(_03998_),
    .A(net2111),
    .B(net4668));
 sg13g2_o21ai_1 _20810_ (.B1(_03998_),
    .Y(_01931_),
    .A1(_04619_),
    .A2(net4668));
 sg13g2_nand2_1 _20811_ (.Y(_03999_),
    .A(net1971),
    .B(net4667));
 sg13g2_o21ai_1 _20812_ (.B1(_03999_),
    .Y(_01932_),
    .A1(_04620_),
    .A2(net4667));
 sg13g2_nand2_1 _20813_ (.Y(_04000_),
    .A(net2044),
    .B(net4657));
 sg13g2_o21ai_1 _20814_ (.B1(_04000_),
    .Y(_01933_),
    .A1(_04621_),
    .A2(net4657));
 sg13g2_nand2_1 _20815_ (.Y(_04001_),
    .A(net2365),
    .B(net4655));
 sg13g2_o21ai_1 _20816_ (.B1(_04001_),
    .Y(_01934_),
    .A1(_04622_),
    .A2(net4656));
 sg13g2_nand2_1 _20817_ (.Y(_04002_),
    .A(net2277),
    .B(net4655));
 sg13g2_o21ai_1 _20818_ (.B1(_04002_),
    .Y(_01935_),
    .A1(_04623_),
    .A2(net4655));
 sg13g2_nand2_1 _20819_ (.Y(_04003_),
    .A(net1438),
    .B(net4645));
 sg13g2_o21ai_1 _20820_ (.B1(_04003_),
    .Y(_01936_),
    .A1(_04624_),
    .A2(net4645));
 sg13g2_nand2_1 _20821_ (.Y(_04004_),
    .A(net1265),
    .B(net4620));
 sg13g2_o21ai_1 _20822_ (.B1(_04004_),
    .Y(_01937_),
    .A1(_04625_),
    .A2(net4623));
 sg13g2_nand2_1 _20823_ (.Y(_04005_),
    .A(net2042),
    .B(net4621));
 sg13g2_o21ai_1 _20824_ (.B1(_04005_),
    .Y(_01938_),
    .A1(_04626_),
    .A2(net4621));
 sg13g2_nand2_1 _20825_ (.Y(_04006_),
    .A(net1966),
    .B(net4635));
 sg13g2_o21ai_1 _20826_ (.B1(_04006_),
    .Y(_01939_),
    .A1(_04627_),
    .A2(net4635));
 sg13g2_nand2_1 _20827_ (.Y(_04007_),
    .A(net1908),
    .B(net4612));
 sg13g2_o21ai_1 _20828_ (.B1(_04007_),
    .Y(_01940_),
    .A1(_04628_),
    .A2(net4613));
 sg13g2_nand2_1 _20829_ (.Y(_04008_),
    .A(net1379),
    .B(net4610));
 sg13g2_o21ai_1 _20830_ (.B1(_04008_),
    .Y(_01941_),
    .A1(_04629_),
    .A2(net4610));
 sg13g2_nand2_1 _20831_ (.Y(_04009_),
    .A(net2167),
    .B(net4575));
 sg13g2_o21ai_1 _20832_ (.B1(_04009_),
    .Y(_01942_),
    .A1(_04630_),
    .A2(net4575));
 sg13g2_nand2_1 _20833_ (.Y(_04010_),
    .A(net1296),
    .B(net4575));
 sg13g2_o21ai_1 _20834_ (.B1(_04010_),
    .Y(_01943_),
    .A1(_04631_),
    .A2(net4576));
 sg13g2_nand2_1 _20835_ (.Y(_04011_),
    .A(net1528),
    .B(net4579));
 sg13g2_o21ai_1 _20836_ (.B1(_04011_),
    .Y(_01944_),
    .A1(_04632_),
    .A2(net4580));
 sg13g2_nand2_1 _20837_ (.Y(_04012_),
    .A(net1641),
    .B(net4633));
 sg13g2_o21ai_1 _20838_ (.B1(_04012_),
    .Y(_01945_),
    .A1(_04633_),
    .A2(net4630));
 sg13g2_nand2_1 _20839_ (.Y(_04013_),
    .A(net2276),
    .B(net4634));
 sg13g2_o21ai_1 _20840_ (.B1(_04013_),
    .Y(_01946_),
    .A1(_04634_),
    .A2(net4634));
 sg13g2_nand2_1 _20841_ (.Y(_04014_),
    .A(net2212),
    .B(net4633));
 sg13g2_o21ai_1 _20842_ (.B1(_04014_),
    .Y(_01947_),
    .A1(_04635_),
    .A2(net4633));
 sg13g2_nand2_1 _20843_ (.Y(_04015_),
    .A(net1847),
    .B(net4677));
 sg13g2_o21ai_1 _20844_ (.B1(_04015_),
    .Y(_01948_),
    .A1(_04636_),
    .A2(net4677));
 sg13g2_nand2_1 _20845_ (.Y(_04016_),
    .A(net1360),
    .B(net4679));
 sg13g2_o21ai_1 _20846_ (.B1(_04016_),
    .Y(_01949_),
    .A1(_04637_),
    .A2(net4679));
 sg13g2_nand2_1 _20847_ (.Y(_04017_),
    .A(net1925),
    .B(net4680));
 sg13g2_o21ai_1 _20848_ (.B1(_04017_),
    .Y(_01950_),
    .A1(_04638_),
    .A2(net4680));
 sg13g2_nand2_1 _20849_ (.Y(_04018_),
    .A(net1321),
    .B(net4691));
 sg13g2_o21ai_1 _20850_ (.B1(_04018_),
    .Y(_01951_),
    .A1(_04639_),
    .A2(net4691));
 sg13g2_nand2_1 _20851_ (.Y(_04019_),
    .A(net1585),
    .B(net4692));
 sg13g2_o21ai_1 _20852_ (.B1(_04019_),
    .Y(_01952_),
    .A1(_04640_),
    .A2(net4692));
 sg13g2_nand2_1 _20853_ (.Y(_04020_),
    .A(net1968),
    .B(net4692));
 sg13g2_o21ai_1 _20854_ (.B1(_04020_),
    .Y(_01953_),
    .A1(_04641_),
    .A2(net4692));
 sg13g2_nand2_1 _20855_ (.Y(_04021_),
    .A(net1798),
    .B(net4693));
 sg13g2_o21ai_1 _20856_ (.B1(_04021_),
    .Y(_01954_),
    .A1(_04642_),
    .A2(net4693));
 sg13g2_nand2_1 _20857_ (.Y(_04022_),
    .A(net1315),
    .B(net4700));
 sg13g2_o21ai_1 _20858_ (.B1(_04022_),
    .Y(_01955_),
    .A1(_04643_),
    .A2(net4681));
 sg13g2_nand2_1 _20859_ (.Y(_04023_),
    .A(net1352),
    .B(net4687));
 sg13g2_o21ai_1 _20860_ (.B1(_04023_),
    .Y(_01956_),
    .A1(_04644_),
    .A2(net4687));
 sg13g2_nand2_1 _20861_ (.Y(_04024_),
    .A(net2328),
    .B(net4686));
 sg13g2_o21ai_1 _20862_ (.B1(_04024_),
    .Y(_01957_),
    .A1(_04645_),
    .A2(net4687));
 sg13g2_nand2_1 _20863_ (.Y(_04025_),
    .A(net2282),
    .B(net4686));
 sg13g2_o21ai_1 _20864_ (.B1(_04025_),
    .Y(_01958_),
    .A1(_04646_),
    .A2(net4686));
 sg13g2_nand2_1 _20865_ (.Y(_04026_),
    .A(net1481),
    .B(net4686));
 sg13g2_o21ai_1 _20866_ (.B1(_04026_),
    .Y(_01959_),
    .A1(_04647_),
    .A2(net4686));
 sg13g2_nand2_1 _20867_ (.Y(_04027_),
    .A(net1329),
    .B(net4685));
 sg13g2_o21ai_1 _20868_ (.B1(_04027_),
    .Y(_01960_),
    .A1(_04648_),
    .A2(net4685));
 sg13g2_nand2_1 _20869_ (.Y(_04028_),
    .A(net1243),
    .B(net4683));
 sg13g2_o21ai_1 _20870_ (.B1(_04028_),
    .Y(_01961_),
    .A1(_04649_),
    .A2(net4683));
 sg13g2_nand2_1 _20871_ (.Y(_04029_),
    .A(net1806),
    .B(net4641));
 sg13g2_o21ai_1 _20872_ (.B1(_04029_),
    .Y(_01962_),
    .A1(_04650_),
    .A2(net4641));
 sg13g2_nand2_1 _20873_ (.Y(_04030_),
    .A(net1514),
    .B(net4636));
 sg13g2_o21ai_1 _20874_ (.B1(_04030_),
    .Y(_01963_),
    .A1(_04651_),
    .A2(net4636));
 sg13g2_nand2_1 _20875_ (.Y(_04031_),
    .A(net1774),
    .B(net4661));
 sg13g2_o21ai_1 _20876_ (.B1(_04031_),
    .Y(_01964_),
    .A1(_04652_),
    .A2(net4661));
 sg13g2_nand2_1 _20877_ (.Y(_04032_),
    .A(net1282),
    .B(net4647));
 sg13g2_o21ai_1 _20878_ (.B1(_04032_),
    .Y(_01965_),
    .A1(_04653_),
    .A2(net4647));
 sg13g2_nand2_1 _20879_ (.Y(_04033_),
    .A(net1770),
    .B(net4653));
 sg13g2_o21ai_1 _20880_ (.B1(_04033_),
    .Y(_01966_),
    .A1(_04654_),
    .A2(net4646));
 sg13g2_nand2_1 _20881_ (.Y(_04034_),
    .A(net2547),
    .B(net4647));
 sg13g2_o21ai_1 _20882_ (.B1(_04034_),
    .Y(_01967_),
    .A1(_04655_),
    .A2(net4646));
 sg13g2_nand2_1 _20883_ (.Y(_04035_),
    .A(net1593),
    .B(net4644));
 sg13g2_o21ai_1 _20884_ (.B1(_04035_),
    .Y(_01968_),
    .A1(_04656_),
    .A2(net4644));
 sg13g2_nand2_1 _20885_ (.Y(_04036_),
    .A(net2068),
    .B(net4644));
 sg13g2_o21ai_1 _20886_ (.B1(_04036_),
    .Y(_01969_),
    .A1(_04657_),
    .A2(net4644));
 sg13g2_nand2_1 _20887_ (.Y(_04037_),
    .A(net2320),
    .B(net4616));
 sg13g2_o21ai_1 _20888_ (.B1(_04037_),
    .Y(_01970_),
    .A1(_04658_),
    .A2(net4616));
 sg13g2_nand2_1 _20889_ (.Y(_04038_),
    .A(net2045),
    .B(net4607));
 sg13g2_o21ai_1 _20890_ (.B1(_04038_),
    .Y(_01971_),
    .A1(_04659_),
    .A2(net4607));
 sg13g2_nand2_1 _20891_ (.Y(_04039_),
    .A(net1745),
    .B(net4607));
 sg13g2_o21ai_1 _20892_ (.B1(_04039_),
    .Y(_01972_),
    .A1(_04660_),
    .A2(net4609));
 sg13g2_nand2_1 _20893_ (.Y(_04040_),
    .A(net2125),
    .B(net4609));
 sg13g2_o21ai_1 _20894_ (.B1(_04040_),
    .Y(_01973_),
    .A1(_04661_),
    .A2(net4572));
 sg13g2_nand2_1 _20895_ (.Y(_04041_),
    .A(net1782),
    .B(net4572));
 sg13g2_o21ai_1 _20896_ (.B1(_04041_),
    .Y(_01974_),
    .A1(_04662_),
    .A2(net4572));
 sg13g2_nand2_1 _20897_ (.Y(_04042_),
    .A(net2246),
    .B(net4573));
 sg13g2_o21ai_1 _20898_ (.B1(_04042_),
    .Y(_01975_),
    .A1(_04663_),
    .A2(net4573));
 sg13g2_nand2_1 _20899_ (.Y(_04043_),
    .A(net1342),
    .B(net4577));
 sg13g2_o21ai_1 _20900_ (.B1(_04043_),
    .Y(_01976_),
    .A1(_04664_),
    .A2(net4577));
 sg13g2_nand2_1 _20901_ (.Y(_04044_),
    .A(net1473),
    .B(net4584));
 sg13g2_o21ai_1 _20902_ (.B1(_04044_),
    .Y(_01977_),
    .A1(_04665_),
    .A2(net4584));
 sg13g2_nand2_1 _20903_ (.Y(_04045_),
    .A(net1630),
    .B(net4585));
 sg13g2_o21ai_1 _20904_ (.B1(_04045_),
    .Y(_01978_),
    .A1(_04666_),
    .A2(net4585));
 sg13g2_nand2_1 _20905_ (.Y(_04046_),
    .A(net1350),
    .B(net4675));
 sg13g2_o21ai_1 _20906_ (.B1(_04046_),
    .Y(_01979_),
    .A1(_04667_),
    .A2(net4675));
 sg13g2_nand2_1 _20907_ (.Y(_04047_),
    .A(net1909),
    .B(net4676));
 sg13g2_o21ai_1 _20908_ (.B1(_04047_),
    .Y(_01980_),
    .A1(_04668_),
    .A2(net4676));
 sg13g2_nand2_1 _20909_ (.Y(_04048_),
    .A(net1923),
    .B(net4594));
 sg13g2_o21ai_1 _20910_ (.B1(_04048_),
    .Y(_01981_),
    .A1(_04669_),
    .A2(net4594));
 sg13g2_nand2_1 _20911_ (.Y(_04049_),
    .A(net1637),
    .B(net4593));
 sg13g2_o21ai_1 _20912_ (.B1(_04049_),
    .Y(_01982_),
    .A1(_04670_),
    .A2(net4593));
 sg13g2_nand2_1 _20913_ (.Y(_04050_),
    .A(net1558),
    .B(net4599));
 sg13g2_o21ai_1 _20914_ (.B1(_04050_),
    .Y(_01983_),
    .A1(_04671_),
    .A2(net4599));
 sg13g2_nand2_1 _20915_ (.Y(_04051_),
    .A(net1647),
    .B(net4604));
 sg13g2_o21ai_1 _20916_ (.B1(_04051_),
    .Y(_01984_),
    .A1(_04672_),
    .A2(net4604));
 sg13g2_nand2_1 _20917_ (.Y(_04052_),
    .A(net2141),
    .B(net4696));
 sg13g2_o21ai_1 _20918_ (.B1(_04052_),
    .Y(_01985_),
    .A1(_04673_),
    .A2(net4696));
 sg13g2_nand2_1 _20919_ (.Y(_04053_),
    .A(net2175),
    .B(net4697));
 sg13g2_o21ai_1 _20920_ (.B1(_04053_),
    .Y(_01986_),
    .A1(_04674_),
    .A2(net4697));
 sg13g2_nand2_1 _20921_ (.Y(_04054_),
    .A(net2460),
    .B(net4706));
 sg13g2_o21ai_1 _20922_ (.B1(_04054_),
    .Y(_01987_),
    .A1(_04675_),
    .A2(net4706));
 sg13g2_nand2_1 _20923_ (.Y(_04055_),
    .A(net2074),
    .B(net4706));
 sg13g2_o21ai_1 _20924_ (.B1(_04055_),
    .Y(_01988_),
    .A1(_04676_),
    .A2(net4706));
 sg13g2_nand2_1 _20925_ (.Y(_04056_),
    .A(net2197),
    .B(net4728));
 sg13g2_o21ai_1 _20926_ (.B1(_04056_),
    .Y(_01989_),
    .A1(_04677_),
    .A2(net4728));
 sg13g2_nand2_1 _20927_ (.Y(_04057_),
    .A(net1476),
    .B(net4688));
 sg13g2_o21ai_1 _20928_ (.B1(_04057_),
    .Y(_01990_),
    .A1(_04678_),
    .A2(net4689));
 sg13g2_nand2_1 _20929_ (.Y(_04058_),
    .A(net1463),
    .B(net4715));
 sg13g2_o21ai_1 _20930_ (.B1(_04058_),
    .Y(_01991_),
    .A1(_04679_),
    .A2(net4715));
 sg13g2_nand2_1 _20931_ (.Y(_04059_),
    .A(net1317),
    .B(net4716));
 sg13g2_o21ai_1 _20932_ (.B1(_04059_),
    .Y(_01992_),
    .A1(_04680_),
    .A2(net4716));
 sg13g2_nand2_1 _20933_ (.Y(_04060_),
    .A(net1789),
    .B(net4710));
 sg13g2_o21ai_1 _20934_ (.B1(_04060_),
    .Y(_01993_),
    .A1(_04681_),
    .A2(net4711));
 sg13g2_nand2_1 _20935_ (.Y(_04061_),
    .A(net1354),
    .B(net4642));
 sg13g2_o21ai_1 _20936_ (.B1(_04061_),
    .Y(_01994_),
    .A1(_04682_),
    .A2(net4642));
 sg13g2_nand2_1 _20937_ (.Y(_04062_),
    .A(net1676),
    .B(net4641));
 sg13g2_o21ai_1 _20938_ (.B1(_04062_),
    .Y(_01995_),
    .A1(_04683_),
    .A2(net4641));
 sg13g2_nand2_1 _20939_ (.Y(_04063_),
    .A(net1797),
    .B(net4662));
 sg13g2_o21ai_1 _20940_ (.B1(_04063_),
    .Y(_01996_),
    .A1(_04684_),
    .A2(net4662));
 sg13g2_nand2_1 _20941_ (.Y(_04064_),
    .A(net2151),
    .B(net4663));
 sg13g2_o21ai_1 _20942_ (.B1(_04064_),
    .Y(_01997_),
    .A1(_04685_),
    .A2(net4663));
 sg13g2_nand2_1 _20943_ (.Y(_04065_),
    .A(net1420),
    .B(net4656));
 sg13g2_o21ai_1 _20944_ (.B1(_04065_),
    .Y(_01998_),
    .A1(_04686_),
    .A2(net4654));
 sg13g2_nand2_1 _20945_ (.Y(_04066_),
    .A(net1543),
    .B(net4653));
 sg13g2_o21ai_1 _20946_ (.B1(_04066_),
    .Y(_01999_),
    .A1(_04687_),
    .A2(net4654));
 sg13g2_nand2_1 _20947_ (.Y(_04067_),
    .A(net1496),
    .B(net4645));
 sg13g2_o21ai_1 _20948_ (.B1(_04067_),
    .Y(_02000_),
    .A1(_04688_),
    .A2(net4645));
 sg13g2_nand2_1 _20949_ (.Y(_04068_),
    .A(net1325),
    .B(net4620));
 sg13g2_o21ai_1 _20950_ (.B1(_04068_),
    .Y(_02001_),
    .A1(_04689_),
    .A2(net4620));
 sg13g2_nand2_1 _20951_ (.Y(_04069_),
    .A(net1776),
    .B(net4617));
 sg13g2_o21ai_1 _20952_ (.B1(_04069_),
    .Y(_02002_),
    .A1(_04690_),
    .A2(net4618));
 sg13g2_nand2_1 _20953_ (.Y(_04070_),
    .A(net1635),
    .B(net4621));
 sg13g2_o21ai_1 _20954_ (.B1(_04070_),
    .Y(_02003_),
    .A1(_04691_),
    .A2(net4621));
 sg13g2_nand2_1 _20955_ (.Y(_04071_),
    .A(net2195),
    .B(net4612));
 sg13g2_o21ai_1 _20956_ (.B1(_04071_),
    .Y(_02004_),
    .A1(_04692_),
    .A2(net4613));
 sg13g2_nand2_1 _20957_ (.Y(_04072_),
    .A(net1517),
    .B(net4571));
 sg13g2_o21ai_1 _20958_ (.B1(_04072_),
    .Y(_02005_),
    .A1(_04693_),
    .A2(net4575));
 sg13g2_nand2_1 _20959_ (.Y(_04073_),
    .A(\TRNG.Padded_Out[378] ),
    .B(net4574));
 sg13g2_o21ai_1 _20960_ (.B1(_04073_),
    .Y(_02006_),
    .A1(_04694_),
    .A2(net4574));
 sg13g2_nand2_1 _20961_ (.Y(_04074_),
    .A(net1346),
    .B(net4573));
 sg13g2_o21ai_1 _20962_ (.B1(_04074_),
    .Y(_02007_),
    .A1(_04695_),
    .A2(net4574));
 sg13g2_nand2_1 _20963_ (.Y(_04075_),
    .A(net1534),
    .B(net4579));
 sg13g2_o21ai_1 _20964_ (.B1(_04075_),
    .Y(_02008_),
    .A1(_04696_),
    .A2(net4577));
 sg13g2_nand2_1 _20965_ (.Y(_04076_),
    .A(net2010),
    .B(net4628));
 sg13g2_o21ai_1 _20966_ (.B1(_04076_),
    .Y(_02009_),
    .A1(_04697_),
    .A2(net4628));
 sg13g2_nand2_1 _20967_ (.Y(_04077_),
    .A(net1323),
    .B(net4631));
 sg13g2_o21ai_1 _20968_ (.B1(_04077_),
    .Y(_02010_),
    .A1(_04698_),
    .A2(net4631));
 sg13g2_nand2_1 _20969_ (.Y(_04078_),
    .A(net1366),
    .B(net4633));
 sg13g2_o21ai_1 _20970_ (.B1(_04078_),
    .Y(_02011_),
    .A1(_04699_),
    .A2(net4634));
 sg13g2_nand2_1 _20971_ (.Y(_04079_),
    .A(net1311),
    .B(net4677));
 sg13g2_o21ai_1 _20972_ (.B1(_04079_),
    .Y(_02012_),
    .A1(_04700_),
    .A2(net4677));
 sg13g2_nand2_1 _20973_ (.Y(_04080_),
    .A(net1987),
    .B(net4591));
 sg13g2_o21ai_1 _20974_ (.B1(_04080_),
    .Y(_02013_),
    .A1(_04701_),
    .A2(net4591));
 sg13g2_nand2_1 _20975_ (.Y(_04081_),
    .A(\TRNG.Padded_Out[386] ),
    .B(net4679));
 sg13g2_o21ai_1 _20976_ (.B1(_04081_),
    .Y(_02014_),
    .A1(_04702_),
    .A2(net4595));
 sg13g2_nand2_1 _20977_ (.Y(_04082_),
    .A(\TRNG.Padded_Out[387] ),
    .B(net4599));
 sg13g2_o21ai_1 _20978_ (.B1(_04082_),
    .Y(_02015_),
    .A1(_04703_),
    .A2(net4599));
 sg13g2_nand2_1 _20979_ (.Y(_04083_),
    .A(net2016),
    .B(net4600));
 sg13g2_o21ai_1 _20980_ (.B1(_04083_),
    .Y(_02016_),
    .A1(_04704_),
    .A2(net4600));
 sg13g2_nand2_1 _20981_ (.Y(_04084_),
    .A(net1629),
    .B(net4695));
 sg13g2_o21ai_1 _20982_ (.B1(_04084_),
    .Y(_02017_),
    .A1(_04705_),
    .A2(net4695));
 sg13g2_nand2_1 _20983_ (.Y(_04085_),
    .A(net1288),
    .B(net4693));
 sg13g2_o21ai_1 _20984_ (.B1(_04085_),
    .Y(_02018_),
    .A1(_04706_),
    .A2(net4693));
 sg13g2_nand2_1 _20985_ (.Y(_04086_),
    .A(net2319),
    .B(net4704));
 sg13g2_o21ai_1 _20986_ (.B1(_04086_),
    .Y(_02019_),
    .A1(_04707_),
    .A2(net4704));
 sg13g2_nand2_1 _20987_ (.Y(_04087_),
    .A(net1337),
    .B(net4707));
 sg13g2_o21ai_1 _20988_ (.B1(_04087_),
    .Y(_02020_),
    .A1(_04708_),
    .A2(net4707));
 sg13g2_nand2_1 _20989_ (.Y(_04088_),
    .A(net1881),
    .B(net4726));
 sg13g2_o21ai_1 _20990_ (.B1(_04088_),
    .Y(_02021_),
    .A1(_04709_),
    .A2(net4726));
 sg13g2_nand2_1 _20991_ (.Y(_04089_),
    .A(net1581),
    .B(net4727));
 sg13g2_o21ai_1 _20992_ (.B1(_04089_),
    .Y(_02022_),
    .A1(_04710_),
    .A2(net4727));
 sg13g2_nand2_1 _20993_ (.Y(_04090_),
    .A(net1304),
    .B(net4722));
 sg13g2_o21ai_1 _20994_ (.B1(_04090_),
    .Y(_02023_),
    .A1(_04711_),
    .A2(net4722));
 sg13g2_nand2_1 _20995_ (.Y(_04091_),
    .A(net1333),
    .B(net4689));
 sg13g2_o21ai_1 _20996_ (.B1(_04091_),
    .Y(_02024_),
    .A1(_04712_),
    .A2(net4689));
 sg13g2_nand2_1 _20997_ (.Y(_04092_),
    .A(net2170),
    .B(net4684));
 sg13g2_o21ai_1 _20998_ (.B1(_04092_),
    .Y(_02025_),
    .A1(_04713_),
    .A2(net4684));
 sg13g2_nand2_1 _20999_ (.Y(_04093_),
    .A(net1769),
    .B(net4710));
 sg13g2_o21ai_1 _21000_ (.B1(_04093_),
    .Y(_02026_),
    .A1(_04714_),
    .A2(net4710));
 sg13g2_nand2_1 _21001_ (.Y(_04094_),
    .A(net1627),
    .B(net4669));
 sg13g2_o21ai_1 _21002_ (.B1(_04094_),
    .Y(_02027_),
    .A1(_04715_),
    .A2(net4666));
 sg13g2_nand2_1 _21003_ (.Y(_04095_),
    .A(net1412),
    .B(net4667));
 sg13g2_o21ai_1 _21004_ (.B1(_04095_),
    .Y(_02028_),
    .A1(_04716_),
    .A2(net4666));
 sg13g2_nand2_1 _21005_ (.Y(_04096_),
    .A(net1300),
    .B(net4647));
 sg13g2_o21ai_1 _21006_ (.B1(_04096_),
    .Y(_02029_),
    .A1(_04717_),
    .A2(net4647));
 sg13g2_nand2_1 _21007_ (.Y(_04097_),
    .A(net1605),
    .B(net4653));
 sg13g2_o21ai_1 _21008_ (.B1(_04097_),
    .Y(_02030_),
    .A1(_04718_),
    .A2(net4653));
 sg13g2_nand2_1 _21009_ (.Y(_04098_),
    .A(net2303),
    .B(net4646));
 sg13g2_o21ai_1 _21010_ (.B1(_04098_),
    .Y(_02031_),
    .A1(_04719_),
    .A2(net4646));
 sg13g2_nand2_1 _21011_ (.Y(_04099_),
    .A(net1358),
    .B(net4644));
 sg13g2_o21ai_1 _21012_ (.B1(_04099_),
    .Y(_02032_),
    .A1(_04720_),
    .A2(net4644));
 sg13g2_nand2_1 _21013_ (.Y(_04100_),
    .A(net1918),
    .B(net4619));
 sg13g2_o21ai_1 _21014_ (.B1(_04100_),
    .Y(_02033_),
    .A1(_04721_),
    .A2(net4619));
 sg13g2_nand2_1 _21015_ (.Y(_04101_),
    .A(net2018),
    .B(net4618));
 sg13g2_o21ai_1 _21016_ (.B1(_04101_),
    .Y(_02034_),
    .A1(_04722_),
    .A2(net4616));
 sg13g2_nand2_1 _21017_ (.Y(_04102_),
    .A(net1902),
    .B(net4607));
 sg13g2_o21ai_1 _21018_ (.B1(_04102_),
    .Y(_02035_),
    .A1(_04723_),
    .A2(net4607));
 sg13g2_nand2_1 _21019_ (.Y(_04103_),
    .A(net2171),
    .B(net4607));
 sg13g2_o21ai_1 _21020_ (.B1(_04103_),
    .Y(_02036_),
    .A1(_04724_),
    .A2(net4609));
 sg13g2_nand2_1 _21021_ (.Y(_04104_),
    .A(net1639),
    .B(net4571));
 sg13g2_o21ai_1 _21022_ (.B1(_04104_),
    .Y(_02037_),
    .A1(_04725_),
    .A2(net4571));
 sg13g2_nand2_1 _21023_ (.Y(_04105_),
    .A(net1269),
    .B(net4572));
 sg13g2_o21ai_1 _21024_ (.B1(_04105_),
    .Y(_02038_),
    .A1(_04726_),
    .A2(net4574));
 sg13g2_nand2_1 _21025_ (.Y(_04106_),
    .A(net1309),
    .B(net4579));
 sg13g2_o21ai_1 _21026_ (.B1(_04106_),
    .Y(_02039_),
    .A1(_04727_),
    .A2(net4579));
 sg13g2_nand2_1 _21027_ (.Y(_04107_),
    .A(net1276),
    .B(net4580));
 sg13g2_o21ai_1 _21028_ (.B1(_04107_),
    .Y(_02040_),
    .A1(_04728_),
    .A2(net4580));
 sg13g2_nand2_1 _21029_ (.Y(_04108_),
    .A(net1255),
    .B(net4585));
 sg13g2_o21ai_1 _21030_ (.B1(_04108_),
    .Y(_02041_),
    .A1(_04729_),
    .A2(net4585));
 sg13g2_nand2_1 _21031_ (.Y(_04109_),
    .A(net1669),
    .B(net4591));
 sg13g2_o21ai_1 _21032_ (.B1(_04109_),
    .Y(_02042_),
    .A1(_04730_),
    .A2(net4591));
 sg13g2_nand2_1 _21033_ (.Y(_04110_),
    .A(net1753),
    .B(net4675));
 sg13g2_o21ai_1 _21034_ (.B1(_04110_),
    .Y(_02043_),
    .A1(_04731_),
    .A2(net4675));
 sg13g2_nand2_1 _21035_ (.Y(_04111_),
    .A(net1502),
    .B(net4676));
 sg13g2_o21ai_1 _21036_ (.B1(_04111_),
    .Y(_02044_),
    .A1(_04732_),
    .A2(net4675));
 sg13g2_nand2_1 _21037_ (.Y(_04112_),
    .A(net1251),
    .B(net4679));
 sg13g2_o21ai_1 _21038_ (.B1(_04112_),
    .Y(_02045_),
    .A1(_04733_),
    .A2(net4679));
 sg13g2_nand2_1 _21039_ (.Y(_04113_),
    .A(net1665),
    .B(net4679));
 sg13g2_o21ai_1 _21040_ (.B1(_04113_),
    .Y(_02046_),
    .A1(_04734_),
    .A2(net4679));
 sg13g2_nand2_1 _21041_ (.Y(_04114_),
    .A(net1335),
    .B(net4680));
 sg13g2_o21ai_1 _21042_ (.B1(_04114_),
    .Y(_02047_),
    .A1(_04735_),
    .A2(net4680));
 sg13g2_nand2_1 _21043_ (.Y(_04115_),
    .A(net1863),
    .B(net4695));
 sg13g2_o21ai_1 _21044_ (.B1(_04115_),
    .Y(_02048_),
    .A1(_04736_),
    .A2(net4695));
 sg13g2_nand2_1 _21045_ (.Y(_04116_),
    .A(net1687),
    .B(net4696));
 sg13g2_o21ai_1 _21046_ (.B1(_04116_),
    .Y(_02049_),
    .A1(_04737_),
    .A2(net4695));
 sg13g2_nand2_1 _21047_ (.Y(_04117_),
    .A(net1500),
    .B(net4698));
 sg13g2_o21ai_1 _21048_ (.B1(_04117_),
    .Y(_02050_),
    .A1(_04738_),
    .A2(net4698));
 sg13g2_nand2_1 _21049_ (.Y(_04118_),
    .A(net1929),
    .B(net4704));
 sg13g2_o21ai_1 _21050_ (.B1(_04118_),
    .Y(_02051_),
    .A1(_04739_),
    .A2(net4704));
 sg13g2_nand2_1 _21051_ (.Y(_04119_),
    .A(net1901),
    .B(net4707));
 sg13g2_o21ai_1 _21052_ (.B1(_04119_),
    .Y(_02052_),
    .A1(_04740_),
    .A2(net4707));
 sg13g2_nand2_1 _21053_ (.Y(_04120_),
    .A(net1868),
    .B(net4726));
 sg13g2_o21ai_1 _21054_ (.B1(_04120_),
    .Y(_02053_),
    .A1(_04741_),
    .A2(net4726));
 sg13g2_nand2_1 _21055_ (.Y(_04121_),
    .A(net1551),
    .B(net4725));
 sg13g2_o21ai_1 _21056_ (.B1(_04121_),
    .Y(_02054_),
    .A1(_04742_),
    .A2(net4723));
 sg13g2_nand2_1 _21057_ (.Y(_04122_),
    .A(net1730),
    .B(net4715));
 sg13g2_o21ai_1 _21058_ (.B1(_04122_),
    .Y(_02055_),
    .A1(_04743_),
    .A2(net4715));
 sg13g2_nand2_1 _21059_ (.Y(_04123_),
    .A(net1648),
    .B(net4711));
 sg13g2_o21ai_1 _21060_ (.B1(_04123_),
    .Y(_02056_),
    .A1(_04744_),
    .A2(net4711));
 sg13g2_nand2_1 _21061_ (.Y(_04124_),
    .A(net1824),
    .B(net4710));
 sg13g2_o21ai_1 _21062_ (.B1(_04124_),
    .Y(_02057_),
    .A1(_04745_),
    .A2(net4710));
 sg13g2_nand2_1 _21063_ (.Y(_04125_),
    .A(net1992),
    .B(net4669));
 sg13g2_o21ai_1 _21064_ (.B1(_04125_),
    .Y(_02058_),
    .A1(_04746_),
    .A2(net4669));
 sg13g2_nand2_1 _21065_ (.Y(_04126_),
    .A(net1524),
    .B(net4641));
 sg13g2_o21ai_1 _21066_ (.B1(_04126_),
    .Y(_02059_),
    .A1(_04747_),
    .A2(net4641));
 sg13g2_nand2_1 _21067_ (.Y(_04127_),
    .A(net1547),
    .B(net4664));
 sg13g2_o21ai_1 _21068_ (.B1(_04127_),
    .Y(_02060_),
    .A1(_04748_),
    .A2(net4661));
 sg13g2_nand2_1 _21069_ (.Y(_04128_),
    .A(net1442),
    .B(net4654));
 sg13g2_o21ai_1 _21070_ (.B1(_04128_),
    .Y(_02061_),
    .A1(_04749_),
    .A2(net4654));
 sg13g2_nand2_1 _21071_ (.Y(_04129_),
    .A(net2201),
    .B(net4656));
 sg13g2_o21ai_1 _21072_ (.B1(_04129_),
    .Y(_02062_),
    .A1(_04750_),
    .A2(net4656));
 sg13g2_nand2_1 _21073_ (.Y(_04130_),
    .A(net2362),
    .B(net4655));
 sg13g2_o21ai_1 _21074_ (.B1(_04130_),
    .Y(_02063_),
    .A1(_04751_),
    .A2(net4655));
 sg13g2_nand2_1 _21075_ (.Y(_04131_),
    .A(net1747),
    .B(net4646));
 sg13g2_o21ai_1 _21076_ (.B1(_04131_),
    .Y(_02064_),
    .A1(_04752_),
    .A2(net4646));
 sg13g2_nand2_1 _21077_ (.Y(_04132_),
    .A(net1489),
    .B(net4620));
 sg13g2_o21ai_1 _21078_ (.B1(_04132_),
    .Y(_02065_),
    .A1(_04753_),
    .A2(net4619));
 sg13g2_nand2_1 _21079_ (.Y(_04133_),
    .A(net1814),
    .B(net4619));
 sg13g2_o21ai_1 _21080_ (.B1(_04133_),
    .Y(_02066_),
    .A1(_04754_),
    .A2(net4616));
 sg13g2_nand2_1 _21081_ (.Y(_04134_),
    .A(net1385),
    .B(net4617));
 sg13g2_o21ai_1 _21082_ (.B1(_04134_),
    .Y(_02067_),
    .A1(_04755_),
    .A2(net4617));
 sg13g2_nand2_1 _21083_ (.Y(_04135_),
    .A(net2256),
    .B(net4608));
 sg13g2_o21ai_1 _21084_ (.B1(_04135_),
    .Y(_02068_),
    .A1(_04756_),
    .A2(net4608));
 sg13g2_nand2_1 _21085_ (.Y(_04136_),
    .A(net1512),
    .B(net4609));
 sg13g2_o21ai_1 _21086_ (.B1(_04136_),
    .Y(_02069_),
    .A1(_04757_),
    .A2(net4609));
 sg13g2_nand2_1 _21087_ (.Y(_04137_),
    .A(net1616),
    .B(net4576));
 sg13g2_o21ai_1 _21088_ (.B1(_04137_),
    .Y(_02070_),
    .A1(_04758_),
    .A2(net4575));
 sg13g2_nand2_1 _21089_ (.Y(_04138_),
    .A(net1426),
    .B(net4573));
 sg13g2_o21ai_1 _21090_ (.B1(_04138_),
    .Y(_02071_),
    .A1(_04759_),
    .A2(net4573));
 sg13g2_nand2_1 _21091_ (.Y(_04139_),
    .A(net1522),
    .B(net4578));
 sg13g2_o21ai_1 _21092_ (.B1(_04139_),
    .Y(_02072_),
    .A1(_04760_),
    .A2(net4578));
 sg13g2_nand2_1 _21093_ (.Y(_04140_),
    .A(net1591),
    .B(net4584));
 sg13g2_o21ai_1 _21094_ (.B1(_04140_),
    .Y(_02073_),
    .A1(_04761_),
    .A2(net4584));
 sg13g2_nand2_1 _21095_ (.Y(_04141_),
    .A(net1397),
    .B(net4632));
 sg13g2_o21ai_1 _21096_ (.B1(_04141_),
    .Y(_02074_),
    .A1(_04762_),
    .A2(net4632));
 sg13g2_nand2_1 _21097_ (.Y(_04142_),
    .A(net1589),
    .B(net4677));
 sg13g2_o21ai_1 _21098_ (.B1(_04142_),
    .Y(_02075_),
    .A1(_04763_),
    .A2(net4675));
 sg13g2_nand2_1 _21099_ (.Y(_04143_),
    .A(net2060),
    .B(net4676));
 sg13g2_o21ai_1 _21100_ (.B1(_04143_),
    .Y(_02076_),
    .A1(_04764_),
    .A2(net4676));
 sg13g2_nand2_1 _21101_ (.Y(_04144_),
    .A(net1487),
    .B(net4681));
 sg13g2_o21ai_1 _21102_ (.B1(_04144_),
    .Y(_02077_),
    .A1(_04765_),
    .A2(net4681));
 sg13g2_nand2_1 _21103_ (.Y(_04145_),
    .A(net2097),
    .B(net4681));
 sg13g2_o21ai_1 _21104_ (.B1(_04145_),
    .Y(_02078_),
    .A1(_04766_),
    .A2(net4682));
 sg13g2_nand2_1 _21105_ (.Y(_04146_),
    .A(net1504),
    .B(net4682));
 sg13g2_o21ai_1 _21106_ (.B1(_04146_),
    .Y(_02079_),
    .A1(_04767_),
    .A2(net4680));
 sg13g2_nand2_1 _21107_ (.Y(_04147_),
    .A(net2020),
    .B(net4691));
 sg13g2_o21ai_1 _21108_ (.B1(_04147_),
    .Y(_02080_),
    .A1(_04768_),
    .A2(net4691));
 sg13g2_nand2_1 _21109_ (.Y(_04148_),
    .A(net1977),
    .B(net4694));
 sg13g2_o21ai_1 _21110_ (.B1(_04148_),
    .Y(_02081_),
    .A1(_04769_),
    .A2(net4694));
 sg13g2_nand2_1 _21111_ (.Y(_04149_),
    .A(net1536),
    .B(net4694));
 sg13g2_o21ai_1 _21112_ (.B1(_04149_),
    .Y(_02082_),
    .A1(_04770_),
    .A2(net4694));
 sg13g2_nand2_1 _21113_ (.Y(_04150_),
    .A(net1829),
    .B(net4703));
 sg13g2_o21ai_1 _21114_ (.B1(_04150_),
    .Y(_02083_),
    .A1(_04771_),
    .A2(net4700));
 sg13g2_nand2_1 _21115_ (.Y(_04151_),
    .A(net1595),
    .B(net4700));
 sg13g2_o21ai_1 _21116_ (.B1(_04151_),
    .Y(_02084_),
    .A1(_04772_),
    .A2(net4700));
 sg13g2_nand2_1 _21117_ (.Y(_04152_),
    .A(net1625),
    .B(net4722));
 sg13g2_o21ai_1 _21118_ (.B1(_04152_),
    .Y(_02085_),
    .A1(_04773_),
    .A2(net4722));
 sg13g2_nand2_1 _21119_ (.Y(_04153_),
    .A(net1256),
    .B(net4687));
 sg13g2_o21ai_1 _21120_ (.B1(_04153_),
    .Y(_02086_),
    .A1(_04774_),
    .A2(net4687));
 sg13g2_nand2_1 _21121_ (.Y(_04154_),
    .A(net1456),
    .B(net4686));
 sg13g2_o21ai_1 _21122_ (.B1(_04154_),
    .Y(_02087_),
    .A1(_04775_),
    .A2(net4686));
 sg13g2_nand2_1 _21123_ (.Y(_04155_),
    .A(net2168),
    .B(net4685));
 sg13g2_o21ai_1 _21124_ (.B1(_04155_),
    .Y(_02088_),
    .A1(_04776_),
    .A2(net4685));
 sg13g2_nand2_1 _21125_ (.Y(_04156_),
    .A(net1714),
    .B(net4683));
 sg13g2_o21ai_1 _21126_ (.B1(_04156_),
    .Y(_02089_),
    .A1(_04777_),
    .A2(net4683));
 sg13g2_nand2_1 _21127_ (.Y(_04157_),
    .A(net1434),
    .B(net4639));
 sg13g2_o21ai_1 _21128_ (.B1(_04157_),
    .Y(_02090_),
    .A1(_04778_),
    .A2(net4639));
 sg13g2_nand2_1 _21129_ (.Y(_04158_),
    .A(net1567),
    .B(net4666));
 sg13g2_o21ai_1 _21130_ (.B1(_04158_),
    .Y(_02091_),
    .A1(_04779_),
    .A2(net4666));
 sg13g2_nand2_1 _21131_ (.Y(_04159_),
    .A(net1450),
    .B(net4662));
 sg13g2_o21ai_1 _21132_ (.B1(_04159_),
    .Y(_02092_),
    .A1(_04780_),
    .A2(net4662));
 sg13g2_nand2_1 _21133_ (.Y(_04160_),
    .A(net1883),
    .B(net4657));
 sg13g2_o21ai_1 _21134_ (.B1(_04160_),
    .Y(_02093_),
    .A1(_04781_),
    .A2(net4657));
 sg13g2_nand2_1 _21135_ (.Y(_04161_),
    .A(net1612),
    .B(net4657));
 sg13g2_o21ai_1 _21136_ (.B1(_04161_),
    .Y(_02094_),
    .A1(_04782_),
    .A2(net4657));
 sg13g2_nand2_1 _21137_ (.Y(_04162_),
    .A(net2223),
    .B(net4653));
 sg13g2_o21ai_1 _21138_ (.B1(_04162_),
    .Y(_02095_),
    .A1(_04783_),
    .A2(net4653));
 sg13g2_nand2_1 _21139_ (.Y(_04163_),
    .A(net2250),
    .B(net4646));
 sg13g2_o21ai_1 _21140_ (.B1(_04163_),
    .Y(_02096_),
    .A1(_04784_),
    .A2(net4646));
 sg13g2_nand2_1 _21141_ (.Y(_04164_),
    .A(net2309),
    .B(net4619));
 sg13g2_o21ai_1 _21142_ (.B1(_04164_),
    .Y(_02097_),
    .A1(_04785_),
    .A2(net4619));
 sg13g2_nand2_1 _21143_ (.Y(_04165_),
    .A(net2096),
    .B(net4616));
 sg13g2_o21ai_1 _21144_ (.B1(_04165_),
    .Y(_02098_),
    .A1(_04786_),
    .A2(net4616));
 sg13g2_nand2_1 _21145_ (.Y(_04166_),
    .A(net1812),
    .B(net4621));
 sg13g2_o21ai_1 _21146_ (.B1(_04166_),
    .Y(_02099_),
    .A1(_04787_),
    .A2(net4617));
 sg13g2_nand2_1 _21147_ (.Y(_04167_),
    .A(net2159),
    .B(net4609));
 sg13g2_o21ai_1 _21148_ (.B1(_04167_),
    .Y(_02100_),
    .A1(_04788_),
    .A2(net4609));
 sg13g2_nand2_1 _21149_ (.Y(_04168_),
    .A(net1695),
    .B(net4571));
 sg13g2_o21ai_1 _21150_ (.B1(_04168_),
    .Y(_02101_),
    .A1(_04789_),
    .A2(net4572));
 sg13g2_nand2_1 _21151_ (.Y(_04169_),
    .A(net1557),
    .B(net4571));
 sg13g2_o21ai_1 _21152_ (.B1(_04169_),
    .Y(_02102_),
    .A1(_04790_),
    .A2(net4571));
 sg13g2_nand2_1 _21153_ (.Y(_04170_),
    .A(net2147),
    .B(net4575));
 sg13g2_o21ai_1 _21154_ (.B1(_04170_),
    .Y(_02103_),
    .A1(_04791_),
    .A2(net4576));
 sg13g2_nand2_1 _21155_ (.Y(_04171_),
    .A(net1444),
    .B(net4580));
 sg13g2_o21ai_1 _21156_ (.B1(_04171_),
    .Y(_02104_),
    .A1(_04792_),
    .A2(net4580));
 sg13g2_nand2_1 _21157_ (.Y(_04172_),
    .A(net1888),
    .B(net4584));
 sg13g2_o21ai_1 _21158_ (.B1(_04172_),
    .Y(_02105_),
    .A1(_04793_),
    .A2(net4584));
 sg13g2_nand2_1 _21159_ (.Y(_04173_),
    .A(net2399),
    .B(net4633));
 sg13g2_o21ai_1 _21160_ (.B1(_04173_),
    .Y(_02106_),
    .A1(_04794_),
    .A2(net4633));
 sg13g2_nand2_1 _21161_ (.Y(_04174_),
    .A(net1597),
    .B(net4633));
 sg13g2_o21ai_1 _21162_ (.B1(_04174_),
    .Y(_02107_),
    .A1(_04795_),
    .A2(net4633));
 sg13g2_nand2_1 _21163_ (.Y(_04175_),
    .A(net2539),
    .B(net4670));
 sg13g2_o21ai_1 _21164_ (.B1(_04175_),
    .Y(_02108_),
    .A1(_04796_),
    .A2(net4672));
 sg13g2_nand2_1 _21165_ (.Y(_04176_),
    .A(net2354),
    .B(net4672));
 sg13g2_o21ai_1 _21166_ (.B1(_04176_),
    .Y(_02109_),
    .A1(_04797_),
    .A2(net4672));
 sg13g2_nand2_1 _21167_ (.Y(_04177_),
    .A(net2213),
    .B(net4719));
 sg13g2_o21ai_1 _21168_ (.B1(_04177_),
    .Y(_02110_),
    .A1(_04798_),
    .A2(net4718));
 sg13g2_nand2_1 _21169_ (.Y(_04178_),
    .A(net1980),
    .B(net4718));
 sg13g2_o21ai_1 _21170_ (.B1(_04178_),
    .Y(_02111_),
    .A1(_04799_),
    .A2(net4718));
 sg13g2_nand2_1 _21171_ (.Y(_04179_),
    .A(net2809),
    .B(net4719));
 sg13g2_o21ai_1 _21172_ (.B1(_04179_),
    .Y(_02112_),
    .A1(_04800_),
    .A2(net4718));
 sg13g2_nand2_1 _21173_ (.Y(_04180_),
    .A(net2860),
    .B(net4730));
 sg13g2_o21ai_1 _21174_ (.B1(_04180_),
    .Y(_02113_),
    .A1(_04801_),
    .A2(net4729));
 sg13g2_nand2_1 _21175_ (.Y(_04181_),
    .A(net1508),
    .B(net4729));
 sg13g2_o21ai_1 _21176_ (.B1(_04181_),
    .Y(_02114_),
    .A1(_04802_),
    .A2(net4729));
 sg13g2_nand2_1 _21177_ (.Y(_04182_),
    .A(net1272),
    .B(net4724));
 sg13g2_o21ai_1 _21178_ (.B1(_04182_),
    .Y(_02115_),
    .A1(_04803_),
    .A2(net4725));
 sg13g2_nand2_1 _21179_ (.Y(_04183_),
    .A(net1663),
    .B(net4724));
 sg13g2_o21ai_1 _21180_ (.B1(_04183_),
    .Y(_02116_),
    .A1(_04804_),
    .A2(net4724));
 sg13g2_nand2_1 _21181_ (.Y(_04184_),
    .A(net2582),
    .B(net4729));
 sg13g2_o21ai_1 _21182_ (.B1(_04184_),
    .Y(_02117_),
    .A1(_04805_),
    .A2(net4724));
 sg13g2_nand2_1 _21183_ (.Y(_04185_),
    .A(net2480),
    .B(net4718));
 sg13g2_o21ai_1 _21184_ (.B1(_04185_),
    .Y(_02118_),
    .A1(_04806_),
    .A2(net4718));
 sg13g2_nand2_1 _21185_ (.Y(_04186_),
    .A(net2442),
    .B(net4720));
 sg13g2_o21ai_1 _21186_ (.B1(_04186_),
    .Y(_02119_),
    .A1(_04807_),
    .A2(net4720));
 sg13g2_nand2_1 _21187_ (.Y(_04187_),
    .A(net2441),
    .B(net4720));
 sg13g2_o21ai_1 _21188_ (.B1(_04187_),
    .Y(_02120_),
    .A1(_04808_),
    .A2(net4720));
 sg13g2_nand2_1 _21189_ (.Y(_04188_),
    .A(net2293),
    .B(net4673));
 sg13g2_o21ai_1 _21190_ (.B1(_04188_),
    .Y(_02121_),
    .A1(_04809_),
    .A2(net4673));
 sg13g2_nand2_1 _21191_ (.Y(_04189_),
    .A(net2472),
    .B(net4672));
 sg13g2_o21ai_1 _21192_ (.B1(_04189_),
    .Y(_02122_),
    .A1(_04810_),
    .A2(net4672));
 sg13g2_nand2_1 _21193_ (.Y(_04190_),
    .A(net2666),
    .B(net4672));
 sg13g2_o21ai_1 _21194_ (.B1(_04190_),
    .Y(_02123_),
    .A1(_04811_),
    .A2(net4672));
 sg13g2_nand2_1 _21195_ (.Y(_04191_),
    .A(net2511),
    .B(net4671));
 sg13g2_o21ai_1 _21196_ (.B1(_04191_),
    .Y(_02124_),
    .A1(_04812_),
    .A2(net4671));
 sg13g2_nand2_1 _21197_ (.Y(_04192_),
    .A(net2733),
    .B(net4670));
 sg13g2_o21ai_1 _21198_ (.B1(_04192_),
    .Y(_02125_),
    .A1(_04813_),
    .A2(net4670));
 sg13g2_nand2_1 _21199_ (.Y(_04193_),
    .A(net2526),
    .B(net4671));
 sg13g2_o21ai_1 _21200_ (.B1(_04193_),
    .Y(_02126_),
    .A1(_04814_),
    .A2(net4671));
 sg13g2_nand2_1 _21201_ (.Y(_04194_),
    .A(net2685),
    .B(net4659));
 sg13g2_o21ai_1 _21202_ (.B1(_04194_),
    .Y(_02127_),
    .A1(_04815_),
    .A2(net4659));
 sg13g2_nand2_1 _21203_ (.Y(_04195_),
    .A(net3356),
    .B(net4655));
 sg13g2_o21ai_1 _21204_ (.B1(_04195_),
    .Y(_02128_),
    .A1(_04816_),
    .A2(net4655));
 sg13g2_nand2_1 _21205_ (.Y(_04196_),
    .A(net2997),
    .B(net4659));
 sg13g2_o21ai_1 _21206_ (.B1(_04196_),
    .Y(_02129_),
    .A1(_04817_),
    .A2(net4655));
 sg13g2_nand2_1 _21207_ (.Y(_04197_),
    .A(net2700),
    .B(net4659));
 sg13g2_o21ai_1 _21208_ (.B1(_04197_),
    .Y(_02130_),
    .A1(_04818_),
    .A2(net4659));
 sg13g2_nand2_1 _21209_ (.Y(_04198_),
    .A(net2464),
    .B(net4659));
 sg13g2_o21ai_1 _21210_ (.B1(_04198_),
    .Y(_02131_),
    .A1(_04819_),
    .A2(net4659));
 sg13g2_nand2_1 _21211_ (.Y(_04199_),
    .A(net2575),
    .B(net4671));
 sg13g2_o21ai_1 _21212_ (.B1(_04199_),
    .Y(_02132_),
    .A1(_04820_),
    .A2(net4671));
 sg13g2_nand2_1 _21213_ (.Y(_04200_),
    .A(net2378),
    .B(net4672));
 sg13g2_o21ai_1 _21214_ (.B1(_04200_),
    .Y(_02133_),
    .A1(_04821_),
    .A2(net4673));
 sg13g2_nand2_1 _21215_ (.Y(_04201_),
    .A(net2580),
    .B(net4720));
 sg13g2_o21ai_1 _21216_ (.B1(_04201_),
    .Y(_02134_),
    .A1(_04822_),
    .A2(net4720));
 sg13g2_nand2_1 _21217_ (.Y(_04202_),
    .A(net1356),
    .B(net4720));
 sg13g2_o21ai_1 _21218_ (.B1(_04202_),
    .Y(_02135_),
    .A1(_04823_),
    .A2(net4720));
 sg13g2_nand2_1 _21219_ (.Y(_04203_),
    .A(net2364),
    .B(net4719));
 sg13g2_o21ai_1 _21220_ (.B1(_04203_),
    .Y(_02136_),
    .A1(_04824_),
    .A2(net4718));
 sg13g2_nand2_1 _21221_ (.Y(_04204_),
    .A(net2357),
    .B(net4718));
 sg13g2_o21ai_1 _21222_ (.B1(_04204_),
    .Y(_02137_),
    .A1(_04825_),
    .A2(net4719));
 sg13g2_nand2_1 _21223_ (.Y(_04205_),
    .A(net1608),
    .B(net4729));
 sg13g2_o21ai_1 _21224_ (.B1(_04205_),
    .Y(_02138_),
    .A1(_04826_),
    .A2(net4729));
 sg13g2_nor2_1 _21225_ (.A(net2501),
    .B(net4729),
    .Y(_04206_));
 sg13g2_a21oi_1 _21226_ (.A1(_04340_),
    .A2(net4729),
    .Y(_02139_),
    .B1(_04206_));
 sg13g2_nor2_1 _21227_ (.A(net3544),
    .B(_03088_),
    .Y(_04207_));
 sg13g2_nor2_2 _21228_ (.A(_04946_),
    .B(_03088_),
    .Y(_04208_));
 sg13g2_a21oi_1 _21229_ (.A1(\TRNG.state[0] ),
    .A2(_04343_),
    .Y(_04209_),
    .B1(_04208_));
 sg13g2_nor2_1 _21230_ (.A(_04207_),
    .B(_04209_),
    .Y(_02140_));
 sg13g2_nor2_1 _21231_ (.A(net5333),
    .B(net5321),
    .Y(_04210_));
 sg13g2_a22oi_1 _21232_ (.Y(_04211_),
    .B1(_04210_),
    .B2(_03088_),
    .A2(_04208_),
    .A1(net3479));
 sg13g2_inv_1 _21233_ (.Y(_02141_),
    .A(_04211_));
 sg13g2_nor2b_1 _21234_ (.A(_00125_),
    .B_N(net5333),
    .Y(_04212_));
 sg13g2_xnor2_1 _21235_ (.Y(_04213_),
    .A(net3443),
    .B(net5333));
 sg13g2_a22oi_1 _21236_ (.Y(_04214_),
    .B1(_04213_),
    .B2(_03088_),
    .A2(_04208_),
    .A1(net5514));
 sg13g2_inv_1 _21237_ (.Y(_02142_),
    .A(net3444));
 sg13g2_xnor2_1 _21238_ (.Y(_04215_),
    .A(net3264),
    .B(_04212_));
 sg13g2_a22oi_1 _21239_ (.Y(_04216_),
    .B1(net3265),
    .B2(_03088_),
    .A2(_04208_),
    .A1(net5509));
 sg13g2_inv_1 _21240_ (.Y(_02143_),
    .A(_04216_));
 sg13g2_nand3_1 _21241_ (.B(net5514),
    .C(net5333),
    .A(net5510),
    .Y(_04217_));
 sg13g2_xor2_1 _21242_ (.B(_04217_),
    .A(net3222),
    .X(_04218_));
 sg13g2_a22oi_1 _21243_ (.Y(_04219_),
    .B1(net3223),
    .B2(_03088_),
    .A2(_04208_),
    .A1(net5508));
 sg13g2_inv_1 _21244_ (.Y(_02144_),
    .A(_04219_));
 sg13g2_buf_1 _21245_ (.A(net2880),
    .X(_01082_));
 sg13g2_dfrbp_1 _21246_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net23),
    .D(net3393),
    .Q_N(_00115_),
    .Q(\TRNG.uart_tx_inst.currentState[4] ));
 sg13g2_dfrbp_1 _21247_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1128),
    .D(net1897),
    .Q_N(_10888_),
    .Q(\TRNG.uart_tx_inst.currentState[3] ));
 sg13g2_dfrbp_1 _21248_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1127),
    .D(net1211),
    .Q_N(_10887_),
    .Q(\TRNG.uart_tx_inst.currentState[2] ));
 sg13g2_dfrbp_1 _21249_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1126),
    .D(_00311_),
    .Q_N(_10886_),
    .Q(\TRNG.uart_tx_inst.currentState[1] ));
 sg13g2_dfrbp_1 _21250_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1125),
    .D(net2681),
    .Q_N(_10885_),
    .Q(\TRNG.uart_tx_inst.currentState[0] ));
 sg13g2_dfrbp_1 _21251_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1124),
    .D(_00313_),
    .Q_N(_10884_),
    .Q(\TRNG.hash[160] ));
 sg13g2_dfrbp_1 _21252_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1123),
    .D(_00314_),
    .Q_N(_10883_),
    .Q(\TRNG.hash[65] ));
 sg13g2_dfrbp_1 _21253_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1122),
    .D(_00315_),
    .Q_N(_10882_),
    .Q(\TRNG.hash[64] ));
 sg13g2_dfrbp_1 _21254_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net24),
    .D(_00316_),
    .Q_N(_10889_),
    .Q(\TRNG.hash[128] ));
 sg13g2_dfrbp_1 _21255_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net25),
    .D(_00064_),
    .Q_N(_10890_),
    .Q(\TRNG.sha256.expand.dout1[0] ));
 sg13g2_dfrbp_1 _21256_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net26),
    .D(net3917),
    .Q_N(_10891_),
    .Q(\TRNG.sha256.expand.dout1[1] ));
 sg13g2_dfrbp_1 _21257_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net27),
    .D(_00086_),
    .Q_N(_10892_),
    .Q(\TRNG.sha256.expand.dout1[2] ));
 sg13g2_dfrbp_1 _21258_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net28),
    .D(_00089_),
    .Q_N(_10893_),
    .Q(\TRNG.sha256.expand.dout1[3] ));
 sg13g2_dfrbp_1 _21259_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net29),
    .D(_00090_),
    .Q_N(_10894_),
    .Q(\TRNG.sha256.expand.dout1[4] ));
 sg13g2_dfrbp_1 _21260_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net30),
    .D(_00091_),
    .Q_N(_10895_),
    .Q(\TRNG.sha256.expand.dout1[5] ));
 sg13g2_dfrbp_1 _21261_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net31),
    .D(net3905),
    .Q_N(_10896_),
    .Q(\TRNG.sha256.expand.dout1[6] ));
 sg13g2_dfrbp_1 _21262_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net32),
    .D(net3908),
    .Q_N(_10897_),
    .Q(\TRNG.sha256.expand.dout1[7] ));
 sg13g2_dfrbp_1 _21263_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net33),
    .D(_00094_),
    .Q_N(_10898_),
    .Q(\TRNG.sha256.expand.dout1[8] ));
 sg13g2_dfrbp_1 _21264_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net34),
    .D(_00095_),
    .Q_N(_10899_),
    .Q(\TRNG.sha256.expand.dout1[9] ));
 sg13g2_dfrbp_1 _21265_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net35),
    .D(_00065_),
    .Q_N(_10900_),
    .Q(\TRNG.sha256.expand.dout1[10] ));
 sg13g2_dfrbp_1 _21266_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net36),
    .D(_00066_),
    .Q_N(_10901_),
    .Q(\TRNG.sha256.expand.dout1[11] ));
 sg13g2_dfrbp_1 _21267_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net37),
    .D(_00067_),
    .Q_N(_10902_),
    .Q(\TRNG.sha256.expand.dout1[12] ));
 sg13g2_dfrbp_1 _21268_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net38),
    .D(_00068_),
    .Q_N(_10903_),
    .Q(\TRNG.sha256.expand.dout1[13] ));
 sg13g2_dfrbp_1 _21269_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net39),
    .D(_00069_),
    .Q_N(_10904_),
    .Q(\TRNG.sha256.expand.dout1[14] ));
 sg13g2_dfrbp_1 _21270_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net40),
    .D(_00070_),
    .Q_N(_10905_),
    .Q(\TRNG.sha256.expand.dout1[15] ));
 sg13g2_dfrbp_1 _21271_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net41),
    .D(_00071_),
    .Q_N(_10906_),
    .Q(\TRNG.sha256.expand.dout1[16] ));
 sg13g2_dfrbp_1 _21272_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net42),
    .D(net3914),
    .Q_N(_10907_),
    .Q(\TRNG.sha256.expand.dout1[17] ));
 sg13g2_dfrbp_1 _21273_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net43),
    .D(net3881),
    .Q_N(_10908_),
    .Q(\TRNG.sha256.expand.dout1[18] ));
 sg13g2_dfrbp_1 _21274_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net44),
    .D(_00074_),
    .Q_N(_10909_),
    .Q(\TRNG.sha256.expand.dout1[19] ));
 sg13g2_dfrbp_1 _21275_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net45),
    .D(_00076_),
    .Q_N(_10910_),
    .Q(\TRNG.sha256.expand.dout1[20] ));
 sg13g2_dfrbp_1 _21276_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net46),
    .D(_00077_),
    .Q_N(_10911_),
    .Q(\TRNG.sha256.expand.dout1[21] ));
 sg13g2_dfrbp_1 _21277_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net47),
    .D(net3930),
    .Q_N(_10912_),
    .Q(\TRNG.sha256.expand.dout1[22] ));
 sg13g2_dfrbp_1 _21278_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net48),
    .D(net3891),
    .Q_N(_10913_),
    .Q(\TRNG.sha256.expand.dout1[23] ));
 sg13g2_dfrbp_1 _21279_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net49),
    .D(_00080_),
    .Q_N(_10914_),
    .Q(\TRNG.sha256.expand.dout1[24] ));
 sg13g2_dfrbp_1 _21280_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net50),
    .D(_00081_),
    .Q_N(_10915_),
    .Q(\TRNG.sha256.expand.dout1[25] ));
 sg13g2_dfrbp_1 _21281_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net51),
    .D(_00082_),
    .Q_N(_10916_),
    .Q(\TRNG.sha256.expand.dout1[26] ));
 sg13g2_dfrbp_1 _21282_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net52),
    .D(_00083_),
    .Q_N(_10917_),
    .Q(\TRNG.sha256.expand.dout1[27] ));
 sg13g2_dfrbp_1 _21283_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net53),
    .D(_00084_),
    .Q_N(_10918_),
    .Q(\TRNG.sha256.expand.dout1[28] ));
 sg13g2_dfrbp_1 _21284_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net54),
    .D(net3927),
    .Q_N(_10919_),
    .Q(\TRNG.sha256.expand.dout1[29] ));
 sg13g2_dfrbp_1 _21285_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net113),
    .D(_00087_),
    .Q_N(_10920_),
    .Q(\TRNG.sha256.expand.dout1[30] ));
 sg13g2_dfrbp_1 _21286_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1121),
    .D(_00088_),
    .Q_N(_10881_),
    .Q(\TRNG.sha256.expand.dout1[31] ));
 sg13g2_dfrbp_1 _21287_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1120),
    .D(_00317_),
    .Q_N(_10880_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][0] ));
 sg13g2_dfrbp_1 _21288_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1119),
    .D(_00318_),
    .Q_N(_10879_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][1] ));
 sg13g2_dfrbp_1 _21289_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1118),
    .D(_00319_),
    .Q_N(_10878_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][2] ));
 sg13g2_dfrbp_1 _21290_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1117),
    .D(_00320_),
    .Q_N(_10877_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][3] ));
 sg13g2_dfrbp_1 _21291_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1116),
    .D(net3205),
    .Q_N(_10876_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][4] ));
 sg13g2_dfrbp_1 _21292_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1115),
    .D(_00322_),
    .Q_N(_10875_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][5] ));
 sg13g2_dfrbp_1 _21293_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1114),
    .D(_00323_),
    .Q_N(_10874_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][6] ));
 sg13g2_dfrbp_1 _21294_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1113),
    .D(_00324_),
    .Q_N(_10873_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][7] ));
 sg13g2_dfrbp_1 _21295_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1112),
    .D(_00325_),
    .Q_N(_10872_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][8] ));
 sg13g2_dfrbp_1 _21296_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1111),
    .D(_00326_),
    .Q_N(_10871_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][9] ));
 sg13g2_dfrbp_1 _21297_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1110),
    .D(_00327_),
    .Q_N(_10870_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][10] ));
 sg13g2_dfrbp_1 _21298_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1109),
    .D(_00328_),
    .Q_N(_10869_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][11] ));
 sg13g2_dfrbp_1 _21299_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1108),
    .D(_00329_),
    .Q_N(_10868_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][12] ));
 sg13g2_dfrbp_1 _21300_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1107),
    .D(_00330_),
    .Q_N(_10867_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][13] ));
 sg13g2_dfrbp_1 _21301_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1106),
    .D(_00331_),
    .Q_N(_10866_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][14] ));
 sg13g2_dfrbp_1 _21302_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1105),
    .D(_00332_),
    .Q_N(_10865_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][15] ));
 sg13g2_dfrbp_1 _21303_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1104),
    .D(_00333_),
    .Q_N(_10864_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][16] ));
 sg13g2_dfrbp_1 _21304_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1103),
    .D(_00334_),
    .Q_N(_10863_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][17] ));
 sg13g2_dfrbp_1 _21305_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1102),
    .D(_00335_),
    .Q_N(_10862_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][18] ));
 sg13g2_dfrbp_1 _21306_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1101),
    .D(_00336_),
    .Q_N(_10861_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][19] ));
 sg13g2_dfrbp_1 _21307_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1100),
    .D(_00337_),
    .Q_N(_10860_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][20] ));
 sg13g2_dfrbp_1 _21308_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1099),
    .D(_00338_),
    .Q_N(_10859_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][21] ));
 sg13g2_dfrbp_1 _21309_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1098),
    .D(_00339_),
    .Q_N(_10858_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][22] ));
 sg13g2_dfrbp_1 _21310_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1097),
    .D(_00340_),
    .Q_N(_10857_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][23] ));
 sg13g2_dfrbp_1 _21311_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1096),
    .D(_00341_),
    .Q_N(_10856_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][24] ));
 sg13g2_dfrbp_1 _21312_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1095),
    .D(_00342_),
    .Q_N(_10855_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][25] ));
 sg13g2_dfrbp_1 _21313_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1094),
    .D(_00343_),
    .Q_N(_10854_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][26] ));
 sg13g2_dfrbp_1 _21314_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1093),
    .D(_00344_),
    .Q_N(_10853_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][27] ));
 sg13g2_dfrbp_1 _21315_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1092),
    .D(_00345_),
    .Q_N(_10852_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][28] ));
 sg13g2_dfrbp_1 _21316_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1091),
    .D(_00346_),
    .Q_N(_10851_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][29] ));
 sg13g2_dfrbp_1 _21317_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1090),
    .D(_00347_),
    .Q_N(_10850_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][30] ));
 sg13g2_dfrbp_1 _21318_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1089),
    .D(_00348_),
    .Q_N(_10849_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[4][31] ));
 sg13g2_dfrbp_1 _21319_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1088),
    .D(_00349_),
    .Q_N(_10848_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][0] ));
 sg13g2_dfrbp_1 _21320_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1087),
    .D(_00350_),
    .Q_N(_10847_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][1] ));
 sg13g2_dfrbp_1 _21321_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1086),
    .D(_00351_),
    .Q_N(_10846_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][2] ));
 sg13g2_dfrbp_1 _21322_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1085),
    .D(_00352_),
    .Q_N(_10845_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][3] ));
 sg13g2_dfrbp_1 _21323_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1084),
    .D(net3112),
    .Q_N(_10844_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][4] ));
 sg13g2_dfrbp_1 _21324_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1083),
    .D(_00354_),
    .Q_N(_10843_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][5] ));
 sg13g2_dfrbp_1 _21325_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1082),
    .D(_00355_),
    .Q_N(_10842_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][6] ));
 sg13g2_dfrbp_1 _21326_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1081),
    .D(_00356_),
    .Q_N(_10841_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][7] ));
 sg13g2_dfrbp_1 _21327_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1080),
    .D(_00357_),
    .Q_N(_10840_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][8] ));
 sg13g2_dfrbp_1 _21328_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1079),
    .D(_00358_),
    .Q_N(_10839_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][9] ));
 sg13g2_dfrbp_1 _21329_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1078),
    .D(_00359_),
    .Q_N(_10838_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][10] ));
 sg13g2_dfrbp_1 _21330_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1077),
    .D(_00360_),
    .Q_N(_10837_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][11] ));
 sg13g2_dfrbp_1 _21331_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1076),
    .D(_00361_),
    .Q_N(_10836_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][12] ));
 sg13g2_dfrbp_1 _21332_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1075),
    .D(_00362_),
    .Q_N(_10835_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][13] ));
 sg13g2_dfrbp_1 _21333_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1074),
    .D(net3377),
    .Q_N(_10834_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][14] ));
 sg13g2_dfrbp_1 _21334_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1073),
    .D(_00364_),
    .Q_N(_10833_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][15] ));
 sg13g2_dfrbp_1 _21335_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1072),
    .D(_00365_),
    .Q_N(_10832_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][16] ));
 sg13g2_dfrbp_1 _21336_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1071),
    .D(_00366_),
    .Q_N(_10831_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][17] ));
 sg13g2_dfrbp_1 _21337_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1070),
    .D(_00367_),
    .Q_N(_10830_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][18] ));
 sg13g2_dfrbp_1 _21338_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1069),
    .D(_00368_),
    .Q_N(_10829_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][19] ));
 sg13g2_dfrbp_1 _21339_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1068),
    .D(_00369_),
    .Q_N(_10828_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][20] ));
 sg13g2_dfrbp_1 _21340_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1067),
    .D(_00370_),
    .Q_N(_10827_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][21] ));
 sg13g2_dfrbp_1 _21341_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1066),
    .D(_00371_),
    .Q_N(_10826_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][22] ));
 sg13g2_dfrbp_1 _21342_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1065),
    .D(_00372_),
    .Q_N(_10825_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][23] ));
 sg13g2_dfrbp_1 _21343_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1064),
    .D(_00373_),
    .Q_N(_10824_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][24] ));
 sg13g2_dfrbp_1 _21344_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1063),
    .D(_00374_),
    .Q_N(_10823_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][25] ));
 sg13g2_dfrbp_1 _21345_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1062),
    .D(_00375_),
    .Q_N(_10822_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][26] ));
 sg13g2_dfrbp_1 _21346_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1061),
    .D(_00376_),
    .Q_N(_10821_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][27] ));
 sg13g2_dfrbp_1 _21347_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1060),
    .D(_00377_),
    .Q_N(_10820_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][28] ));
 sg13g2_dfrbp_1 _21348_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1059),
    .D(_00378_),
    .Q_N(_10819_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][29] ));
 sg13g2_dfrbp_1 _21349_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1058),
    .D(_00379_),
    .Q_N(_10818_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][30] ));
 sg13g2_dfrbp_1 _21350_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1057),
    .D(_00380_),
    .Q_N(_10817_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[3][31] ));
 sg13g2_dfrbp_1 _21351_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1056),
    .D(net3039),
    .Q_N(_10816_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][0] ));
 sg13g2_dfrbp_1 _21352_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1055),
    .D(_00382_),
    .Q_N(_10815_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][1] ));
 sg13g2_dfrbp_1 _21353_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1054),
    .D(_00383_),
    .Q_N(_10814_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][2] ));
 sg13g2_dfrbp_1 _21354_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1053),
    .D(net3213),
    .Q_N(_10813_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][3] ));
 sg13g2_dfrbp_1 _21355_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1052),
    .D(net3143),
    .Q_N(_10812_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][4] ));
 sg13g2_dfrbp_1 _21356_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1051),
    .D(_00386_),
    .Q_N(_10811_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][5] ));
 sg13g2_dfrbp_1 _21357_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1050),
    .D(_00387_),
    .Q_N(_10810_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][6] ));
 sg13g2_dfrbp_1 _21358_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1049),
    .D(_00388_),
    .Q_N(_10809_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][7] ));
 sg13g2_dfrbp_1 _21359_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1048),
    .D(_00389_),
    .Q_N(_10808_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][8] ));
 sg13g2_dfrbp_1 _21360_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1047),
    .D(net3006),
    .Q_N(_10807_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][9] ));
 sg13g2_dfrbp_1 _21361_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1046),
    .D(_00391_),
    .Q_N(_10806_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][10] ));
 sg13g2_dfrbp_1 _21362_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1045),
    .D(net3008),
    .Q_N(_10805_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][11] ));
 sg13g2_dfrbp_1 _21363_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1044),
    .D(_00393_),
    .Q_N(_10804_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][12] ));
 sg13g2_dfrbp_1 _21364_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1043),
    .D(_00394_),
    .Q_N(_10803_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][13] ));
 sg13g2_dfrbp_1 _21365_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1042),
    .D(_00395_),
    .Q_N(_10802_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][14] ));
 sg13g2_dfrbp_1 _21366_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1041),
    .D(_00396_),
    .Q_N(_10801_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][15] ));
 sg13g2_dfrbp_1 _21367_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1040),
    .D(_00397_),
    .Q_N(_10800_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][16] ));
 sg13g2_dfrbp_1 _21368_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1039),
    .D(net2899),
    .Q_N(_10799_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][17] ));
 sg13g2_dfrbp_1 _21369_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1038),
    .D(_00399_),
    .Q_N(_10798_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][18] ));
 sg13g2_dfrbp_1 _21370_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1037),
    .D(net3141),
    .Q_N(_10797_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][19] ));
 sg13g2_dfrbp_1 _21371_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1036),
    .D(_00401_),
    .Q_N(_10796_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][20] ));
 sg13g2_dfrbp_1 _21372_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1035),
    .D(_00402_),
    .Q_N(_10795_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][21] ));
 sg13g2_dfrbp_1 _21373_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1034),
    .D(_00403_),
    .Q_N(_10794_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][22] ));
 sg13g2_dfrbp_1 _21374_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1033),
    .D(_00404_),
    .Q_N(_10793_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][23] ));
 sg13g2_dfrbp_1 _21375_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1032),
    .D(_00405_),
    .Q_N(_10792_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][24] ));
 sg13g2_dfrbp_1 _21376_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1031),
    .D(_00406_),
    .Q_N(_10791_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][25] ));
 sg13g2_dfrbp_1 _21377_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1030),
    .D(_00407_),
    .Q_N(_10790_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][26] ));
 sg13g2_dfrbp_1 _21378_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1029),
    .D(_00408_),
    .Q_N(_10789_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][27] ));
 sg13g2_dfrbp_1 _21379_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1028),
    .D(_00409_),
    .Q_N(_10788_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][28] ));
 sg13g2_dfrbp_1 _21380_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1027),
    .D(_00410_),
    .Q_N(_10787_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][29] ));
 sg13g2_dfrbp_1 _21381_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1026),
    .D(_00411_),
    .Q_N(_10786_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][30] ));
 sg13g2_dfrbp_1 _21382_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1025),
    .D(_00412_),
    .Q_N(_10785_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[15][31] ));
 sg13g2_dfrbp_1 _21383_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1024),
    .D(net2805),
    .Q_N(_10784_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][0] ));
 sg13g2_dfrbp_1 _21384_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1023),
    .D(net2724),
    .Q_N(_10783_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][1] ));
 sg13g2_dfrbp_1 _21385_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1022),
    .D(_00415_),
    .Q_N(_10782_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][2] ));
 sg13g2_dfrbp_1 _21386_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1021),
    .D(_00416_),
    .Q_N(_10781_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][3] ));
 sg13g2_dfrbp_1 _21387_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1020),
    .D(net2688),
    .Q_N(_10780_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][4] ));
 sg13g2_dfrbp_1 _21388_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1019),
    .D(_00418_),
    .Q_N(_10779_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][5] ));
 sg13g2_dfrbp_1 _21389_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1018),
    .D(_00419_),
    .Q_N(_10778_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][6] ));
 sg13g2_dfrbp_1 _21390_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1017),
    .D(_00420_),
    .Q_N(_10777_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][7] ));
 sg13g2_dfrbp_1 _21391_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1016),
    .D(_00421_),
    .Q_N(_10776_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][8] ));
 sg13g2_dfrbp_1 _21392_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1015),
    .D(_00422_),
    .Q_N(_10775_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][9] ));
 sg13g2_dfrbp_1 _21393_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1014),
    .D(_00423_),
    .Q_N(_10774_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][10] ));
 sg13g2_dfrbp_1 _21394_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1013),
    .D(_00424_),
    .Q_N(_10773_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][11] ));
 sg13g2_dfrbp_1 _21395_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1012),
    .D(_00425_),
    .Q_N(_10772_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][12] ));
 sg13g2_dfrbp_1 _21396_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1011),
    .D(_00426_),
    .Q_N(_10771_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][13] ));
 sg13g2_dfrbp_1 _21397_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1010),
    .D(_00427_),
    .Q_N(_10770_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][14] ));
 sg13g2_dfrbp_1 _21398_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1009),
    .D(_00428_),
    .Q_N(_10769_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][15] ));
 sg13g2_dfrbp_1 _21399_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1008),
    .D(_00429_),
    .Q_N(_10768_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][16] ));
 sg13g2_dfrbp_1 _21400_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1007),
    .D(_00430_),
    .Q_N(_10767_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][17] ));
 sg13g2_dfrbp_1 _21401_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1006),
    .D(_00431_),
    .Q_N(_10766_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][18] ));
 sg13g2_dfrbp_1 _21402_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1005),
    .D(_00432_),
    .Q_N(_10765_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][19] ));
 sg13g2_dfrbp_1 _21403_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1004),
    .D(_00433_),
    .Q_N(_10764_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][20] ));
 sg13g2_dfrbp_1 _21404_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1003),
    .D(_00434_),
    .Q_N(_10763_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][21] ));
 sg13g2_dfrbp_1 _21405_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1002),
    .D(_00435_),
    .Q_N(_10762_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][22] ));
 sg13g2_dfrbp_1 _21406_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1001),
    .D(_00436_),
    .Q_N(_10761_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][23] ));
 sg13g2_dfrbp_1 _21407_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1000),
    .D(_00437_),
    .Q_N(_10760_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][24] ));
 sg13g2_dfrbp_1 _21408_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net999),
    .D(_00438_),
    .Q_N(_10759_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][25] ));
 sg13g2_dfrbp_1 _21409_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net998),
    .D(_00439_),
    .Q_N(_10758_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][26] ));
 sg13g2_dfrbp_1 _21410_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net997),
    .D(net2834),
    .Q_N(_10757_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][27] ));
 sg13g2_dfrbp_1 _21411_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net996),
    .D(_00441_),
    .Q_N(_10756_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][28] ));
 sg13g2_dfrbp_1 _21412_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net995),
    .D(_00442_),
    .Q_N(_10755_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][29] ));
 sg13g2_dfrbp_1 _21413_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net994),
    .D(_00443_),
    .Q_N(_10754_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][30] ));
 sg13g2_dfrbp_1 _21414_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net993),
    .D(_00444_),
    .Q_N(_10753_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[2][31] ));
 sg13g2_dfrbp_1 _21415_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net992),
    .D(net2792),
    .Q_N(_10752_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][0] ));
 sg13g2_dfrbp_1 _21416_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net991),
    .D(net2947),
    .Q_N(_10751_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][1] ));
 sg13g2_dfrbp_1 _21417_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net990),
    .D(_00447_),
    .Q_N(_10750_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][2] ));
 sg13g2_dfrbp_1 _21418_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net989),
    .D(_00448_),
    .Q_N(_10749_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][3] ));
 sg13g2_dfrbp_1 _21419_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net988),
    .D(net2706),
    .Q_N(_10748_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][4] ));
 sg13g2_dfrbp_1 _21420_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net987),
    .D(_00450_),
    .Q_N(_10747_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][5] ));
 sg13g2_dfrbp_1 _21421_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net986),
    .D(_00451_),
    .Q_N(_10746_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][6] ));
 sg13g2_dfrbp_1 _21422_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net985),
    .D(_00452_),
    .Q_N(_10745_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][7] ));
 sg13g2_dfrbp_1 _21423_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net984),
    .D(_00453_),
    .Q_N(_10744_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][8] ));
 sg13g2_dfrbp_1 _21424_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net983),
    .D(_00454_),
    .Q_N(_10743_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][9] ));
 sg13g2_dfrbp_1 _21425_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net982),
    .D(_00455_),
    .Q_N(_10742_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][10] ));
 sg13g2_dfrbp_1 _21426_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net981),
    .D(_00456_),
    .Q_N(_10741_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][11] ));
 sg13g2_dfrbp_1 _21427_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net980),
    .D(_00457_),
    .Q_N(_10740_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][12] ));
 sg13g2_dfrbp_1 _21428_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net979),
    .D(_00458_),
    .Q_N(_10739_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][13] ));
 sg13g2_dfrbp_1 _21429_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net978),
    .D(_00459_),
    .Q_N(_10738_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][14] ));
 sg13g2_dfrbp_1 _21430_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net977),
    .D(_00460_),
    .Q_N(_10737_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][15] ));
 sg13g2_dfrbp_1 _21431_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net976),
    .D(_00461_),
    .Q_N(_10736_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][16] ));
 sg13g2_dfrbp_1 _21432_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net975),
    .D(_00462_),
    .Q_N(_10735_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][17] ));
 sg13g2_dfrbp_1 _21433_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net974),
    .D(_00463_),
    .Q_N(_10734_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][18] ));
 sg13g2_dfrbp_1 _21434_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net973),
    .D(_00464_),
    .Q_N(_10733_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][19] ));
 sg13g2_dfrbp_1 _21435_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net972),
    .D(_00465_),
    .Q_N(_10732_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][20] ));
 sg13g2_dfrbp_1 _21436_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net971),
    .D(_00466_),
    .Q_N(_10731_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][21] ));
 sg13g2_dfrbp_1 _21437_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net970),
    .D(_00467_),
    .Q_N(_10730_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][22] ));
 sg13g2_dfrbp_1 _21438_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net969),
    .D(_00468_),
    .Q_N(_10729_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][23] ));
 sg13g2_dfrbp_1 _21439_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net968),
    .D(_00469_),
    .Q_N(_10728_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][24] ));
 sg13g2_dfrbp_1 _21440_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net967),
    .D(_00470_),
    .Q_N(_10727_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][25] ));
 sg13g2_dfrbp_1 _21441_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net966),
    .D(_00471_),
    .Q_N(_10726_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][26] ));
 sg13g2_dfrbp_1 _21442_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net965),
    .D(_00472_),
    .Q_N(_10725_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][27] ));
 sg13g2_dfrbp_1 _21443_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net964),
    .D(_00473_),
    .Q_N(_10724_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][28] ));
 sg13g2_dfrbp_1 _21444_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net963),
    .D(_00474_),
    .Q_N(_10723_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][29] ));
 sg13g2_dfrbp_1 _21445_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net962),
    .D(_00475_),
    .Q_N(_10722_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][30] ));
 sg13g2_dfrbp_1 _21446_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net286),
    .D(_00476_),
    .Q_N(_10921_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[1][31] ));
 sg13g2_dfrbp_1 _21447_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net961),
    .D(net1135),
    .Q_N(_10721_),
    .Q(\TRNG.sha256.compress.hash_gen.temp[0] ));
 sg13g2_dfrbp_1 _21448_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net960),
    .D(net3564),
    .Q_N(_10720_),
    .Q(\TRNG.hash[130] ));
 sg13g2_dfrbp_1 _21449_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net959),
    .D(net3510),
    .Q_N(_00134_),
    .Q(\TRNG.hash[134] ));
 sg13g2_dfrbp_1 _21450_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net958),
    .D(_00479_),
    .Q_N(_10719_),
    .Q(\TRNG.hash[135] ));
 sg13g2_dfrbp_1 _21451_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net957),
    .D(net3498),
    .Q_N(_10718_),
    .Q(\TRNG.hash[137] ));
 sg13g2_dfrbp_1 _21452_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net956),
    .D(net3650),
    .Q_N(_10717_),
    .Q(\TRNG.hash[139] ));
 sg13g2_dfrbp_1 _21453_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net955),
    .D(net3483),
    .Q_N(_00137_),
    .Q(\TRNG.hash[148] ));
 sg13g2_dfrbp_1 _21454_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net954),
    .D(net3618),
    .Q_N(_00139_),
    .Q(\TRNG.hash[149] ));
 sg13g2_dfrbp_1 _21455_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net953),
    .D(_00484_),
    .Q_N(_10716_),
    .Q(\TRNG.hash[151] ));
 sg13g2_dfrbp_1 _21456_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net952),
    .D(_00485_),
    .Q_N(_10715_),
    .Q(\TRNG.hash[153] ));
 sg13g2_dfrbp_1 _21457_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net951),
    .D(net3543),
    .Q_N(_00142_),
    .Q(\TRNG.hash[155] ));
 sg13g2_dfrbp_1 _21458_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net950),
    .D(net2593),
    .Q_N(_10714_),
    .Q(\TRNG.hash[156] ));
 sg13g2_dfrbp_1 _21459_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net949),
    .D(net3507),
    .Q_N(_00144_),
    .Q(\TRNG.hash[158] ));
 sg13g2_dfrbp_1 _21460_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net948),
    .D(net3746),
    .Q_N(_10713_),
    .Q(\TRNG.hash[1] ));
 sg13g2_dfrbp_1 _21461_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net947),
    .D(net3691),
    .Q_N(_00157_),
    .Q(\TRNG.hash[2] ));
 sg13g2_dfrbp_1 _21462_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net946),
    .D(net3548),
    .Q_N(_00149_),
    .Q(\TRNG.hash[5] ));
 sg13g2_dfrbp_1 _21463_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net945),
    .D(net3584),
    .Q_N(_00151_),
    .Q(\TRNG.hash[6] ));
 sg13g2_dfrbp_1 _21464_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net944),
    .D(net3462),
    .Q_N(_10712_),
    .Q(\TRNG.hash[7] ));
 sg13g2_dfrbp_1 _21465_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net943),
    .D(net3621),
    .Q_N(_00152_),
    .Q(\TRNG.hash[9] ));
 sg13g2_dfrbp_1 _21466_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net942),
    .D(net3575),
    .Q_N(_00154_),
    .Q(\TRNG.hash[12] ));
 sg13g2_dfrbp_1 _21467_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net941),
    .D(net3705),
    .Q_N(_10711_),
    .Q(\TRNG.hash[13] ));
 sg13g2_dfrbp_1 _21468_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net940),
    .D(_00497_),
    .Q_N(_10710_),
    .Q(\TRNG.hash[16] ));
 sg13g2_dfrbp_1 _21469_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net939),
    .D(_00498_),
    .Q_N(_10709_),
    .Q(\TRNG.hash[17] ));
 sg13g2_dfrbp_1 _21470_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net938),
    .D(net3578),
    .Q_N(_10708_),
    .Q(\TRNG.hash[18] ));
 sg13g2_dfrbp_1 _21471_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net937),
    .D(_00500_),
    .Q_N(_10707_),
    .Q(\TRNG.hash[19] ));
 sg13g2_dfrbp_1 _21472_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net936),
    .D(_00501_),
    .Q_N(_10706_),
    .Q(\TRNG.hash[20] ));
 sg13g2_dfrbp_1 _21473_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net935),
    .D(_00502_),
    .Q_N(_10705_),
    .Q(\TRNG.hash[26] ));
 sg13g2_dfrbp_1 _21474_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net934),
    .D(net3600),
    .Q_N(_10704_),
    .Q(\TRNG.hash[29] ));
 sg13g2_dfrbp_1 _21475_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net933),
    .D(net3755),
    .Q_N(_10703_),
    .Q(\TRNG.hash[31] ));
 sg13g2_dfrbp_1 _21476_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net932),
    .D(net3518),
    .Q_N(_00160_),
    .Q(\TRNG.hash[34] ));
 sg13g2_dfrbp_1 _21477_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net931),
    .D(net3502),
    .Q_N(_00161_),
    .Q(\TRNG.hash[36] ));
 sg13g2_dfrbp_1 _21478_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net930),
    .D(net3491),
    .Q_N(_00163_),
    .Q(\TRNG.hash[38] ));
 sg13g2_dfrbp_1 _21479_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net929),
    .D(net3562),
    .Q_N(_10702_),
    .Q(\TRNG.hash[41] ));
 sg13g2_dfrbp_1 _21480_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net928),
    .D(net3413),
    .Q_N(_00165_),
    .Q(\TRNG.hash[42] ));
 sg13g2_dfrbp_1 _21481_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net927),
    .D(net3488),
    .Q_N(_00166_),
    .Q(\TRNG.hash[45] ));
 sg13g2_dfrbp_1 _21482_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net926),
    .D(net3481),
    .Q_N(_00168_),
    .Q(\TRNG.hash[50] ));
 sg13g2_dfrbp_1 _21483_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net925),
    .D(_00512_),
    .Q_N(_10701_),
    .Q(\TRNG.hash[51] ));
 sg13g2_dfrbp_1 _21484_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net924),
    .D(net3550),
    .Q_N(_00169_),
    .Q(\TRNG.hash[52] ));
 sg13g2_dfrbp_1 _21485_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net923),
    .D(net3573),
    .Q_N(_00212_),
    .Q(\TRNG.hash[53] ));
 sg13g2_dfrbp_1 _21486_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net922),
    .D(_00515_),
    .Q_N(_00177_),
    .Q(\TRNG.hash[54] ));
 sg13g2_dfrbp_1 _21487_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net921),
    .D(net3471),
    .Q_N(_00170_),
    .Q(\TRNG.hash[61] ));
 sg13g2_dfrbp_1 _21488_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net920),
    .D(_00517_),
    .Q_N(_10700_),
    .Q(\TRNG.hash[62] ));
 sg13g2_dfrbp_1 _21489_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net919),
    .D(_00518_),
    .Q_N(_10699_),
    .Q(\TRNG.hash[63] ));
 sg13g2_dfrbp_1 _21490_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net918),
    .D(net3458),
    .Q_N(_00178_),
    .Q(\TRNG.hash[68] ));
 sg13g2_dfrbp_1 _21491_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net917),
    .D(_00520_),
    .Q_N(_10698_),
    .Q(\TRNG.hash[69] ));
 sg13g2_dfrbp_1 _21492_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net916),
    .D(net3825),
    .Q_N(_00192_),
    .Q(\TRNG.hash[70] ));
 sg13g2_dfrbp_1 _21493_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net915),
    .D(net3494),
    .Q_N(_00179_),
    .Q(\TRNG.hash[72] ));
 sg13g2_dfrbp_1 _21494_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net914),
    .D(net3810),
    .Q_N(_10697_),
    .Q(\TRNG.hash[73] ));
 sg13g2_dfrbp_1 _21495_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net913),
    .D(net3739),
    .Q_N(_00193_),
    .Q(\TRNG.hash[74] ));
 sg13g2_dfrbp_1 _21496_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net912),
    .D(net3420),
    .Q_N(_00181_),
    .Q(\TRNG.hash[76] ));
 sg13g2_dfrbp_1 _21497_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net911),
    .D(net3417),
    .Q_N(_00183_),
    .Q(\TRNG.hash[79] ));
 sg13g2_dfrbp_1 _21498_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net910),
    .D(net3603),
    .Q_N(_10696_),
    .Q(\TRNG.hash[81] ));
 sg13g2_dfrbp_1 _21499_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net909),
    .D(_00528_),
    .Q_N(_10695_),
    .Q(\TRNG.hash[83] ));
 sg13g2_dfrbp_1 _21500_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net908),
    .D(net3383),
    .Q_N(_00186_),
    .Q(\TRNG.hash[84] ));
 sg13g2_dfrbp_1 _21501_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net907),
    .D(_00530_),
    .Q_N(_00213_),
    .Q(\TRNG.hash[85] ));
 sg13g2_dfrbp_1 _21502_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net906),
    .D(net3409),
    .Q_N(_00187_),
    .Q(\TRNG.hash[86] ));
 sg13g2_dfrbp_1 _21503_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net905),
    .D(net3609),
    .Q_N(_00214_),
    .Q(\TRNG.hash[87] ));
 sg13g2_dfrbp_1 _21504_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net904),
    .D(net3473),
    .Q_N(_00188_),
    .Q(\TRNG.hash[90] ));
 sg13g2_dfrbp_1 _21505_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net903),
    .D(net3464),
    .Q_N(_00189_),
    .Q(\TRNG.hash[93] ));
 sg13g2_dfrbp_1 _21506_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net902),
    .D(_00535_),
    .Q_N(_10694_),
    .Q(\TRNG.hash[94] ));
 sg13g2_dfrbp_1 _21507_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net901),
    .D(_00536_),
    .Q_N(_10693_),
    .Q(\TRNG.hash[103] ));
 sg13g2_dfrbp_1 _21508_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net900),
    .D(_00537_),
    .Q_N(_00204_),
    .Q(\TRNG.hash[104] ));
 sg13g2_dfrbp_1 _21509_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net899),
    .D(net3161),
    .Q_N(_00205_),
    .Q(\TRNG.hash[106] ));
 sg13g2_dfrbp_1 _21510_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net898),
    .D(_00539_),
    .Q_N(_10692_),
    .Q(\TRNG.hash[107] ));
 sg13g2_dfrbp_1 _21511_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net897),
    .D(_00540_),
    .Q_N(_10691_),
    .Q(\TRNG.hash[109] ));
 sg13g2_dfrbp_1 _21512_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net896),
    .D(net3135),
    .Q_N(_00209_),
    .Q(\TRNG.hash[111] ));
 sg13g2_dfrbp_1 _21513_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net895),
    .D(_00542_),
    .Q_N(_10690_),
    .Q(\TRNG.hash[112] ));
 sg13g2_dfrbp_1 _21514_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net894),
    .D(net3184),
    .Q_N(_00211_),
    .Q(\TRNG.hash[116] ));
 sg13g2_dfrbp_1 _21515_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net893),
    .D(_00544_),
    .Q_N(_10689_),
    .Q(\TRNG.hash[117] ));
 sg13g2_dfrbp_1 _21516_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net892),
    .D(_00545_),
    .Q_N(_10688_),
    .Q(\TRNG.hash[118] ));
 sg13g2_dfrbp_1 _21517_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net891),
    .D(_00546_),
    .Q_N(_10687_),
    .Q(\TRNG.hash[119] ));
 sg13g2_dfrbp_1 _21518_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net890),
    .D(net3593),
    .Q_N(_00203_),
    .Q(\TRNG.hash[121] ));
 sg13g2_dfrbp_1 _21519_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net889),
    .D(net3660),
    .Q_N(_00202_),
    .Q(\TRNG.hash[122] ));
 sg13g2_dfrbp_1 _21520_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net888),
    .D(_00549_),
    .Q_N(_00201_),
    .Q(\TRNG.hash[123] ));
 sg13g2_dfrbp_1 _21521_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net887),
    .D(_00550_),
    .Q_N(_00199_),
    .Q(\TRNG.hash[125] ));
 sg13g2_dfrbp_1 _21522_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net886),
    .D(_00551_),
    .Q_N(_00198_),
    .Q(\TRNG.hash[127] ));
 sg13g2_dfrbp_1 _21523_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net885),
    .D(net3568),
    .Q_N(_10686_),
    .Q(\TRNG.hash[162] ));
 sg13g2_dfrbp_1 _21524_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net884),
    .D(net3732),
    .Q_N(_10685_),
    .Q(\TRNG.hash[163] ));
 sg13g2_dfrbp_1 _21525_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net883),
    .D(net3514),
    .Q_N(_10684_),
    .Q(\TRNG.hash[167] ));
 sg13g2_dfrbp_1 _21526_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net882),
    .D(net3774),
    .Q_N(_10683_),
    .Q(\TRNG.hash[170] ));
 sg13g2_dfrbp_1 _21527_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net881),
    .D(_00556_),
    .Q_N(_10682_),
    .Q(\TRNG.hash[171] ));
 sg13g2_dfrbp_1 _21528_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net880),
    .D(_00557_),
    .Q_N(_10681_),
    .Q(\TRNG.hash[176] ));
 sg13g2_dfrbp_1 _21529_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net879),
    .D(_00558_),
    .Q_N(_10680_),
    .Q(\TRNG.hash[180] ));
 sg13g2_dfrbp_1 _21530_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net878),
    .D(_00559_),
    .Q_N(_10679_),
    .Q(\TRNG.hash[183] ));
 sg13g2_dfrbp_1 _21531_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net877),
    .D(_00560_),
    .Q_N(_10678_),
    .Q(\TRNG.hash[184] ));
 sg13g2_dfrbp_1 _21532_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net876),
    .D(_00561_),
    .Q_N(_10677_),
    .Q(\TRNG.hash[185] ));
 sg13g2_dfrbp_1 _21533_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net875),
    .D(_00562_),
    .Q_N(_10676_),
    .Q(\TRNG.hash[190] ));
 sg13g2_dfrbp_1 _21534_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net874),
    .D(_00563_),
    .Q_N(_10675_),
    .Q(\TRNG.hash[191] ));
 sg13g2_dfrbp_1 _21535_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net873),
    .D(_00564_),
    .Q_N(_10674_),
    .Q(\TRNG.hash[193] ));
 sg13g2_dfrbp_1 _21536_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net872),
    .D(_00565_),
    .Q_N(_10673_),
    .Q(\TRNG.hash[195] ));
 sg13g2_dfrbp_1 _21537_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net871),
    .D(net3873),
    .Q_N(_10672_),
    .Q(\TRNG.hash[196] ));
 sg13g2_dfrbp_1 _21538_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net870),
    .D(net3864),
    .Q_N(_10671_),
    .Q(\TRNG.hash[197] ));
 sg13g2_dfrbp_1 _21539_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net869),
    .D(_00568_),
    .Q_N(_10670_),
    .Q(\TRNG.hash[198] ));
 sg13g2_dfrbp_1 _21540_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net868),
    .D(net3876),
    .Q_N(_10669_),
    .Q(\TRNG.hash[200] ));
 sg13g2_dfrbp_1 _21541_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net867),
    .D(_00570_),
    .Q_N(_10668_),
    .Q(\TRNG.hash[204] ));
 sg13g2_dfrbp_1 _21542_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net866),
    .D(_00571_),
    .Q_N(_10667_),
    .Q(\TRNG.hash[206] ));
 sg13g2_dfrbp_1 _21543_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net865),
    .D(_00572_),
    .Q_N(_10666_),
    .Q(\TRNG.hash[211] ));
 sg13g2_dfrbp_1 _21544_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net864),
    .D(_00573_),
    .Q_N(_10665_),
    .Q(\TRNG.hash[212] ));
 sg13g2_dfrbp_1 _21545_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net863),
    .D(_00574_),
    .Q_N(_10664_),
    .Q(\TRNG.hash[215] ));
 sg13g2_dfrbp_1 _21546_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net862),
    .D(_00575_),
    .Q_N(_10663_),
    .Q(\TRNG.hash[218] ));
 sg13g2_dfrbp_1 _21547_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net861),
    .D(_00576_),
    .Q_N(_10662_),
    .Q(\TRNG.hash[222] ));
 sg13g2_dfrbp_1 _21548_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net860),
    .D(_00577_),
    .Q_N(_10661_),
    .Q(\TRNG.hash[227] ));
 sg13g2_dfrbp_1 _21549_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net859),
    .D(_00578_),
    .Q_N(_10660_),
    .Q(\TRNG.hash[228] ));
 sg13g2_dfrbp_1 _21550_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net858),
    .D(_00579_),
    .Q_N(_10659_),
    .Q(\TRNG.hash[231] ));
 sg13g2_dfrbp_1 _21551_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net857),
    .D(_00580_),
    .Q_N(_10658_),
    .Q(\TRNG.hash[232] ));
 sg13g2_dfrbp_1 _21552_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net856),
    .D(_00581_),
    .Q_N(_10657_),
    .Q(\TRNG.hash[235] ));
 sg13g2_dfrbp_1 _21553_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net855),
    .D(_00582_),
    .Q_N(_10656_),
    .Q(\TRNG.hash[236] ));
 sg13g2_dfrbp_1 _21554_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net854),
    .D(_00583_),
    .Q_N(_10655_),
    .Q(\TRNG.hash[241] ));
 sg13g2_dfrbp_1 _21555_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net853),
    .D(_00584_),
    .Q_N(_10654_),
    .Q(\TRNG.hash[242] ));
 sg13g2_dfrbp_1 _21556_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net852),
    .D(_00585_),
    .Q_N(_10653_),
    .Q(\TRNG.hash[244] ));
 sg13g2_dfrbp_1 _21557_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net851),
    .D(_00586_),
    .Q_N(_10652_),
    .Q(\TRNG.hash[245] ));
 sg13g2_dfrbp_1 _21558_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net850),
    .D(_00587_),
    .Q_N(_10651_),
    .Q(\TRNG.hash[246] ));
 sg13g2_dfrbp_1 _21559_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net849),
    .D(_00588_),
    .Q_N(_10650_),
    .Q(\TRNG.hash[247] ));
 sg13g2_dfrbp_1 _21560_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net848),
    .D(_00589_),
    .Q_N(_10649_),
    .Q(\TRNG.hash[248] ));
 sg13g2_dfrbp_1 _21561_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net847),
    .D(_00590_),
    .Q_N(_10648_),
    .Q(\TRNG.hash[250] ));
 sg13g2_dfrbp_1 _21562_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net846),
    .D(net3441),
    .Q_N(_10647_),
    .Q(\TRNG.hash[252] ));
 sg13g2_dfrbp_1 _21563_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net845),
    .D(_00592_),
    .Q_N(_10646_),
    .Q(\TRNG.hash[255] ));
 sg13g2_dfrbp_1 _21564_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net844),
    .D(net2551),
    .Q_N(_10645_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][0] ));
 sg13g2_dfrbp_1 _21565_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net843),
    .D(_00594_),
    .Q_N(_10644_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][1] ));
 sg13g2_dfrbp_1 _21566_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net842),
    .D(_00595_),
    .Q_N(_10643_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][2] ));
 sg13g2_dfrbp_1 _21567_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net841),
    .D(_00596_),
    .Q_N(_10642_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][3] ));
 sg13g2_dfrbp_1 _21568_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net840),
    .D(_00597_),
    .Q_N(_10641_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][4] ));
 sg13g2_dfrbp_1 _21569_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net839),
    .D(_00598_),
    .Q_N(_10640_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][5] ));
 sg13g2_dfrbp_1 _21570_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net838),
    .D(_00599_),
    .Q_N(_10639_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][6] ));
 sg13g2_dfrbp_1 _21571_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net837),
    .D(net3020),
    .Q_N(_10638_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][7] ));
 sg13g2_dfrbp_1 _21572_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net836),
    .D(_00601_),
    .Q_N(_10637_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][8] ));
 sg13g2_dfrbp_1 _21573_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net835),
    .D(_00602_),
    .Q_N(_10636_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][9] ));
 sg13g2_dfrbp_1 _21574_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net834),
    .D(_00603_),
    .Q_N(_10635_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][10] ));
 sg13g2_dfrbp_1 _21575_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net833),
    .D(_00604_),
    .Q_N(_10634_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][11] ));
 sg13g2_dfrbp_1 _21576_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net832),
    .D(_00605_),
    .Q_N(_10633_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][12] ));
 sg13g2_dfrbp_1 _21577_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net831),
    .D(_00606_),
    .Q_N(_10632_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][13] ));
 sg13g2_dfrbp_1 _21578_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net830),
    .D(_00607_),
    .Q_N(_10631_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][14] ));
 sg13g2_dfrbp_1 _21579_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net829),
    .D(_00608_),
    .Q_N(_10630_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][15] ));
 sg13g2_dfrbp_1 _21580_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net828),
    .D(_00609_),
    .Q_N(_10629_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][16] ));
 sg13g2_dfrbp_1 _21581_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net827),
    .D(_00610_),
    .Q_N(_10628_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][17] ));
 sg13g2_dfrbp_1 _21582_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net826),
    .D(_00611_),
    .Q_N(_10627_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][18] ));
 sg13g2_dfrbp_1 _21583_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net825),
    .D(_00612_),
    .Q_N(_10626_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][19] ));
 sg13g2_dfrbp_1 _21584_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net824),
    .D(_00613_),
    .Q_N(_10625_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][20] ));
 sg13g2_dfrbp_1 _21585_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net823),
    .D(_00614_),
    .Q_N(_10624_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][21] ));
 sg13g2_dfrbp_1 _21586_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net822),
    .D(_00615_),
    .Q_N(_10623_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][22] ));
 sg13g2_dfrbp_1 _21587_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net821),
    .D(net3308),
    .Q_N(_10622_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][23] ));
 sg13g2_dfrbp_1 _21588_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net820),
    .D(_00617_),
    .Q_N(_10621_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][24] ));
 sg13g2_dfrbp_1 _21589_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net819),
    .D(_00618_),
    .Q_N(_10620_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][25] ));
 sg13g2_dfrbp_1 _21590_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net818),
    .D(_00619_),
    .Q_N(_10619_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][26] ));
 sg13g2_dfrbp_1 _21591_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net817),
    .D(net3278),
    .Q_N(_10618_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][27] ));
 sg13g2_dfrbp_1 _21592_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net816),
    .D(_00621_),
    .Q_N(_10617_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][28] ));
 sg13g2_dfrbp_1 _21593_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net815),
    .D(_00622_),
    .Q_N(_10616_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][29] ));
 sg13g2_dfrbp_1 _21594_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net814),
    .D(_00623_),
    .Q_N(_10615_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][30] ));
 sg13g2_dfrbp_1 _21595_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net813),
    .D(net3103),
    .Q_N(_10614_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[14][31] ));
 sg13g2_dfrbp_1 _21596_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net812),
    .D(_00625_),
    .Q_N(_10613_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][0] ));
 sg13g2_dfrbp_1 _21597_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net811),
    .D(net2856),
    .Q_N(_10612_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][1] ));
 sg13g2_dfrbp_1 _21598_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net810),
    .D(_00627_),
    .Q_N(_10611_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][2] ));
 sg13g2_dfrbp_1 _21599_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net809),
    .D(_00628_),
    .Q_N(_10610_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][3] ));
 sg13g2_dfrbp_1 _21600_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net808),
    .D(net2883),
    .Q_N(_10609_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][4] ));
 sg13g2_dfrbp_1 _21601_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net807),
    .D(_00630_),
    .Q_N(_10608_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][5] ));
 sg13g2_dfrbp_1 _21602_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net806),
    .D(_00631_),
    .Q_N(_10607_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][6] ));
 sg13g2_dfrbp_1 _21603_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net805),
    .D(_00632_),
    .Q_N(_10606_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][7] ));
 sg13g2_dfrbp_1 _21604_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net804),
    .D(_00633_),
    .Q_N(_10605_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][8] ));
 sg13g2_dfrbp_1 _21605_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net803),
    .D(_00634_),
    .Q_N(_10604_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][9] ));
 sg13g2_dfrbp_1 _21606_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net802),
    .D(_00635_),
    .Q_N(_10603_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][10] ));
 sg13g2_dfrbp_1 _21607_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net801),
    .D(_00636_),
    .Q_N(_10602_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][11] ));
 sg13g2_dfrbp_1 _21608_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net800),
    .D(_00637_),
    .Q_N(_10601_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][12] ));
 sg13g2_dfrbp_1 _21609_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net799),
    .D(_00638_),
    .Q_N(_10600_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][13] ));
 sg13g2_dfrbp_1 _21610_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net798),
    .D(_00639_),
    .Q_N(_10599_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][14] ));
 sg13g2_dfrbp_1 _21611_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net797),
    .D(_00640_),
    .Q_N(_10598_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][15] ));
 sg13g2_dfrbp_1 _21612_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net796),
    .D(_00641_),
    .Q_N(_10597_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][16] ));
 sg13g2_dfrbp_1 _21613_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net795),
    .D(_00642_),
    .Q_N(_10596_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][17] ));
 sg13g2_dfrbp_1 _21614_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net794),
    .D(_00643_),
    .Q_N(_10595_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][18] ));
 sg13g2_dfrbp_1 _21615_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net793),
    .D(_00644_),
    .Q_N(_10594_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][19] ));
 sg13g2_dfrbp_1 _21616_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net792),
    .D(_00645_),
    .Q_N(_10593_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][20] ));
 sg13g2_dfrbp_1 _21617_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net791),
    .D(_00646_),
    .Q_N(_10592_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][21] ));
 sg13g2_dfrbp_1 _21618_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net790),
    .D(_00647_),
    .Q_N(_10591_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][22] ));
 sg13g2_dfrbp_1 _21619_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net789),
    .D(_00648_),
    .Q_N(_10590_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][23] ));
 sg13g2_dfrbp_1 _21620_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net788),
    .D(_00649_),
    .Q_N(_10589_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][24] ));
 sg13g2_dfrbp_1 _21621_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net787),
    .D(_00650_),
    .Q_N(_10588_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][25] ));
 sg13g2_dfrbp_1 _21622_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net786),
    .D(_00651_),
    .Q_N(_10587_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][26] ));
 sg13g2_dfrbp_1 _21623_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net785),
    .D(_00652_),
    .Q_N(_10586_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][27] ));
 sg13g2_dfrbp_1 _21624_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net784),
    .D(_00653_),
    .Q_N(_10585_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][28] ));
 sg13g2_dfrbp_1 _21625_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net783),
    .D(_00654_),
    .Q_N(_10584_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][29] ));
 sg13g2_dfrbp_1 _21626_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net782),
    .D(_00655_),
    .Q_N(_10583_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][30] ));
 sg13g2_dfrbp_1 _21627_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net781),
    .D(_00656_),
    .Q_N(_10582_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[5][31] ));
 sg13g2_dfrbp_1 _21628_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net780),
    .D(_00657_),
    .Q_N(_10581_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][0] ));
 sg13g2_dfrbp_1 _21629_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net779),
    .D(_00658_),
    .Q_N(_10580_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][1] ));
 sg13g2_dfrbp_1 _21630_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net778),
    .D(_00659_),
    .Q_N(_10579_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][2] ));
 sg13g2_dfrbp_1 _21631_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net777),
    .D(net2302),
    .Q_N(_10578_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][3] ));
 sg13g2_dfrbp_1 _21632_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net776),
    .D(_00661_),
    .Q_N(_10577_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][4] ));
 sg13g2_dfrbp_1 _21633_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net775),
    .D(_00662_),
    .Q_N(_10576_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][5] ));
 sg13g2_dfrbp_1 _21634_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net774),
    .D(net3349),
    .Q_N(_10575_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][6] ));
 sg13g2_dfrbp_1 _21635_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net773),
    .D(_00664_),
    .Q_N(_10574_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][7] ));
 sg13g2_dfrbp_1 _21636_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net772),
    .D(net3198),
    .Q_N(_10573_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][8] ));
 sg13g2_dfrbp_1 _21637_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net771),
    .D(_00666_),
    .Q_N(_10572_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][9] ));
 sg13g2_dfrbp_1 _21638_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net770),
    .D(_00667_),
    .Q_N(_10571_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][10] ));
 sg13g2_dfrbp_1 _21639_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net769),
    .D(_00668_),
    .Q_N(_10570_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][11] ));
 sg13g2_dfrbp_1 _21640_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net768),
    .D(_00669_),
    .Q_N(_10569_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][12] ));
 sg13g2_dfrbp_1 _21641_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net767),
    .D(_00670_),
    .Q_N(_10568_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][13] ));
 sg13g2_dfrbp_1 _21642_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net766),
    .D(_00671_),
    .Q_N(_10567_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][14] ));
 sg13g2_dfrbp_1 _21643_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net765),
    .D(_00672_),
    .Q_N(_10566_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][15] ));
 sg13g2_dfrbp_1 _21644_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net764),
    .D(_00673_),
    .Q_N(_10565_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][16] ));
 sg13g2_dfrbp_1 _21645_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net762),
    .D(_00674_),
    .Q_N(_10564_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][17] ));
 sg13g2_dfrbp_1 _21646_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net761),
    .D(_00675_),
    .Q_N(_10563_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][18] ));
 sg13g2_dfrbp_1 _21647_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net760),
    .D(net3295),
    .Q_N(_10562_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][19] ));
 sg13g2_dfrbp_1 _21648_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net759),
    .D(_00677_),
    .Q_N(_10561_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][20] ));
 sg13g2_dfrbp_1 _21649_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net758),
    .D(_00678_),
    .Q_N(_10560_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][21] ));
 sg13g2_dfrbp_1 _21650_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net757),
    .D(_00679_),
    .Q_N(_10559_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][22] ));
 sg13g2_dfrbp_1 _21651_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net756),
    .D(_00680_),
    .Q_N(_10558_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][23] ));
 sg13g2_dfrbp_1 _21652_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net755),
    .D(_00681_),
    .Q_N(_10557_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][24] ));
 sg13g2_dfrbp_1 _21653_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net754),
    .D(_00682_),
    .Q_N(_10556_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][25] ));
 sg13g2_dfrbp_1 _21654_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net752),
    .D(_00683_),
    .Q_N(_10555_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][26] ));
 sg13g2_dfrbp_1 _21655_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net751),
    .D(net3346),
    .Q_N(_10554_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][27] ));
 sg13g2_dfrbp_1 _21656_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net750),
    .D(_00685_),
    .Q_N(_10553_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][28] ));
 sg13g2_dfrbp_1 _21657_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net749),
    .D(_00686_),
    .Q_N(_10552_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][29] ));
 sg13g2_dfrbp_1 _21658_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net748),
    .D(net3260),
    .Q_N(_10551_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][30] ));
 sg13g2_dfrbp_1 _21659_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net747),
    .D(_00688_),
    .Q_N(_10550_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[0][31] ));
 sg13g2_dfrbp_1 _21660_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net746),
    .D(net2989),
    .Q_N(_10549_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][0] ));
 sg13g2_dfrbp_1 _21661_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net745),
    .D(net2987),
    .Q_N(_10548_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][1] ));
 sg13g2_dfrbp_1 _21662_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net744),
    .D(_00691_),
    .Q_N(_10547_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][2] ));
 sg13g2_dfrbp_1 _21663_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net743),
    .D(_00692_),
    .Q_N(_10546_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][3] ));
 sg13g2_dfrbp_1 _21664_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net742),
    .D(net3148),
    .Q_N(_10545_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][4] ));
 sg13g2_dfrbp_1 _21665_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net741),
    .D(_00694_),
    .Q_N(_10544_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][5] ));
 sg13g2_dfrbp_1 _21666_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net740),
    .D(_00695_),
    .Q_N(_10543_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][6] ));
 sg13g2_dfrbp_1 _21667_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net739),
    .D(_00696_),
    .Q_N(_10542_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][7] ));
 sg13g2_dfrbp_1 _21668_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net738),
    .D(net2854),
    .Q_N(_10541_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][8] ));
 sg13g2_dfrbp_1 _21669_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net737),
    .D(_00698_),
    .Q_N(_10540_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][9] ));
 sg13g2_dfrbp_1 _21670_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net736),
    .D(net2759),
    .Q_N(_10539_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][10] ));
 sg13g2_dfrbp_1 _21671_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net735),
    .D(_00700_),
    .Q_N(_10538_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][11] ));
 sg13g2_dfrbp_1 _21672_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net734),
    .D(_00701_),
    .Q_N(_10537_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][12] ));
 sg13g2_dfrbp_1 _21673_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net733),
    .D(_00702_),
    .Q_N(_10536_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][13] ));
 sg13g2_dfrbp_1 _21674_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net732),
    .D(_00703_),
    .Q_N(_10535_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][14] ));
 sg13g2_dfrbp_1 _21675_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net731),
    .D(_00704_),
    .Q_N(_10534_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][15] ));
 sg13g2_dfrbp_1 _21676_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net730),
    .D(_00705_),
    .Q_N(_10533_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][16] ));
 sg13g2_dfrbp_1 _21677_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net729),
    .D(_00706_),
    .Q_N(_10532_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][17] ));
 sg13g2_dfrbp_1 _21678_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net728),
    .D(_00707_),
    .Q_N(_10531_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][18] ));
 sg13g2_dfrbp_1 _21679_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net727),
    .D(_00708_),
    .Q_N(_10530_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][19] ));
 sg13g2_dfrbp_1 _21680_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net726),
    .D(_00709_),
    .Q_N(_10529_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][20] ));
 sg13g2_dfrbp_1 _21681_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net725),
    .D(_00710_),
    .Q_N(_10528_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][21] ));
 sg13g2_dfrbp_1 _21682_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net724),
    .D(_00711_),
    .Q_N(_10527_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][22] ));
 sg13g2_dfrbp_1 _21683_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net723),
    .D(_00712_),
    .Q_N(_10526_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][23] ));
 sg13g2_dfrbp_1 _21684_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net722),
    .D(_00713_),
    .Q_N(_10525_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][24] ));
 sg13g2_dfrbp_1 _21685_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net721),
    .D(_00714_),
    .Q_N(_10524_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][25] ));
 sg13g2_dfrbp_1 _21686_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net720),
    .D(_00715_),
    .Q_N(_10523_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][26] ));
 sg13g2_dfrbp_1 _21687_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net719),
    .D(_00716_),
    .Q_N(_10522_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][27] ));
 sg13g2_dfrbp_1 _21688_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net718),
    .D(_00717_),
    .Q_N(_10521_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][28] ));
 sg13g2_dfrbp_1 _21689_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net717),
    .D(_00718_),
    .Q_N(_10520_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][29] ));
 sg13g2_dfrbp_1 _21690_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net716),
    .D(_00719_),
    .Q_N(_10519_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][30] ));
 sg13g2_dfrbp_1 _21691_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net715),
    .D(_00720_),
    .Q_N(_10518_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[7][31] ));
 sg13g2_dfrbp_1 _21692_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net714),
    .D(net3064),
    .Q_N(_10517_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][0] ));
 sg13g2_dfrbp_1 _21693_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net713),
    .D(_00722_),
    .Q_N(_10516_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][1] ));
 sg13g2_dfrbp_1 _21694_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net712),
    .D(_00723_),
    .Q_N(_10515_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][2] ));
 sg13g2_dfrbp_1 _21695_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net711),
    .D(_00724_),
    .Q_N(_10514_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][3] ));
 sg13g2_dfrbp_1 _21696_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net710),
    .D(_00725_),
    .Q_N(_10513_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][4] ));
 sg13g2_dfrbp_1 _21697_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net709),
    .D(_00726_),
    .Q_N(_10512_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][5] ));
 sg13g2_dfrbp_1 _21698_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net708),
    .D(_00727_),
    .Q_N(_10511_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][6] ));
 sg13g2_dfrbp_1 _21699_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net707),
    .D(_00728_),
    .Q_N(_10510_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][7] ));
 sg13g2_dfrbp_1 _21700_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net706),
    .D(_00729_),
    .Q_N(_10509_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][8] ));
 sg13g2_dfrbp_1 _21701_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net705),
    .D(_00730_),
    .Q_N(_10508_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][9] ));
 sg13g2_dfrbp_1 _21702_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net704),
    .D(_00731_),
    .Q_N(_10507_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][10] ));
 sg13g2_dfrbp_1 _21703_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net703),
    .D(_00732_),
    .Q_N(_10506_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][11] ));
 sg13g2_dfrbp_1 _21704_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net702),
    .D(net3334),
    .Q_N(_10505_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][12] ));
 sg13g2_dfrbp_1 _21705_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net701),
    .D(_00734_),
    .Q_N(_10504_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][13] ));
 sg13g2_dfrbp_1 _21706_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net700),
    .D(_00735_),
    .Q_N(_10503_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][14] ));
 sg13g2_dfrbp_1 _21707_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net699),
    .D(net3318),
    .Q_N(_10502_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][15] ));
 sg13g2_dfrbp_1 _21708_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net698),
    .D(_00737_),
    .Q_N(_10501_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][16] ));
 sg13g2_dfrbp_1 _21709_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net697),
    .D(_00738_),
    .Q_N(_10500_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][17] ));
 sg13g2_dfrbp_1 _21710_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net696),
    .D(_00739_),
    .Q_N(_10499_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][18] ));
 sg13g2_dfrbp_1 _21711_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net695),
    .D(_00740_),
    .Q_N(_10498_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][19] ));
 sg13g2_dfrbp_1 _21712_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net694),
    .D(_00741_),
    .Q_N(_10497_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][20] ));
 sg13g2_dfrbp_1 _21713_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net693),
    .D(net3276),
    .Q_N(_10496_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][21] ));
 sg13g2_dfrbp_1 _21714_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net692),
    .D(net3243),
    .Q_N(_10495_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][22] ));
 sg13g2_dfrbp_1 _21715_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net691),
    .D(_00744_),
    .Q_N(_10494_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][23] ));
 sg13g2_dfrbp_1 _21716_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net690),
    .D(_00745_),
    .Q_N(_10493_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][24] ));
 sg13g2_dfrbp_1 _21717_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net689),
    .D(_00746_),
    .Q_N(_10492_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][25] ));
 sg13g2_dfrbp_1 _21718_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net688),
    .D(_00747_),
    .Q_N(_10491_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][26] ));
 sg13g2_dfrbp_1 _21719_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net687),
    .D(net3343),
    .Q_N(_10490_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][27] ));
 sg13g2_dfrbp_1 _21720_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net686),
    .D(net3363),
    .Q_N(_10489_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][28] ));
 sg13g2_dfrbp_1 _21721_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net685),
    .D(_00750_),
    .Q_N(_10488_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][29] ));
 sg13g2_dfrbp_1 _21722_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net684),
    .D(_00751_),
    .Q_N(_10487_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][30] ));
 sg13g2_dfrbp_1 _21723_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net683),
    .D(_00752_),
    .Q_N(_10486_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[8][31] ));
 sg13g2_dfrbp_1 _21724_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net682),
    .D(net2698),
    .Q_N(_10485_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][0] ));
 sg13g2_dfrbp_1 _21725_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net681),
    .D(net2737),
    .Q_N(_10484_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][1] ));
 sg13g2_dfrbp_1 _21726_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net680),
    .D(_00755_),
    .Q_N(_10483_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][2] ));
 sg13g2_dfrbp_1 _21727_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net679),
    .D(_00756_),
    .Q_N(_10482_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][3] ));
 sg13g2_dfrbp_1 _21728_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net678),
    .D(net2971),
    .Q_N(_10481_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][4] ));
 sg13g2_dfrbp_1 _21729_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net677),
    .D(_00758_),
    .Q_N(_10480_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][5] ));
 sg13g2_dfrbp_1 _21730_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net676),
    .D(_00759_),
    .Q_N(_10479_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][6] ));
 sg13g2_dfrbp_1 _21731_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net675),
    .D(_00760_),
    .Q_N(_10478_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][7] ));
 sg13g2_dfrbp_1 _21732_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net674),
    .D(_00761_),
    .Q_N(_10477_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][8] ));
 sg13g2_dfrbp_1 _21733_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net673),
    .D(_00762_),
    .Q_N(_10476_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][9] ));
 sg13g2_dfrbp_1 _21734_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net672),
    .D(_00763_),
    .Q_N(_10475_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][10] ));
 sg13g2_dfrbp_1 _21735_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net671),
    .D(_00764_),
    .Q_N(_10474_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][11] ));
 sg13g2_dfrbp_1 _21736_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net670),
    .D(_00765_),
    .Q_N(_10473_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][12] ));
 sg13g2_dfrbp_1 _21737_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net669),
    .D(_00766_),
    .Q_N(_10472_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][13] ));
 sg13g2_dfrbp_1 _21738_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net668),
    .D(_00767_),
    .Q_N(_10471_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][14] ));
 sg13g2_dfrbp_1 _21739_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net667),
    .D(_00768_),
    .Q_N(_10470_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][15] ));
 sg13g2_dfrbp_1 _21740_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net666),
    .D(net3174),
    .Q_N(_10469_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][16] ));
 sg13g2_dfrbp_1 _21741_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net665),
    .D(_00770_),
    .Q_N(_10468_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][17] ));
 sg13g2_dfrbp_1 _21742_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net664),
    .D(_00771_),
    .Q_N(_10467_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][18] ));
 sg13g2_dfrbp_1 _21743_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net663),
    .D(_00772_),
    .Q_N(_10466_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][19] ));
 sg13g2_dfrbp_1 _21744_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net662),
    .D(_00773_),
    .Q_N(_10465_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][20] ));
 sg13g2_dfrbp_1 _21745_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net661),
    .D(_00774_),
    .Q_N(_10464_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][21] ));
 sg13g2_dfrbp_1 _21746_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net660),
    .D(_00775_),
    .Q_N(_10463_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][22] ));
 sg13g2_dfrbp_1 _21747_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net659),
    .D(_00776_),
    .Q_N(_10462_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][23] ));
 sg13g2_dfrbp_1 _21748_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net658),
    .D(_00777_),
    .Q_N(_10461_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][24] ));
 sg13g2_dfrbp_1 _21749_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net657),
    .D(_00778_),
    .Q_N(_10460_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][25] ));
 sg13g2_dfrbp_1 _21750_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net656),
    .D(_00779_),
    .Q_N(_10459_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][26] ));
 sg13g2_dfrbp_1 _21751_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net655),
    .D(_00780_),
    .Q_N(_10458_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][27] ));
 sg13g2_dfrbp_1 _21752_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net654),
    .D(_00781_),
    .Q_N(_10457_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][28] ));
 sg13g2_dfrbp_1 _21753_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net653),
    .D(_00782_),
    .Q_N(_10456_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][29] ));
 sg13g2_dfrbp_1 _21754_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net652),
    .D(_00783_),
    .Q_N(_10455_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][30] ));
 sg13g2_dfrbp_1 _21755_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net287),
    .D(_00784_),
    .Q_N(_10922_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[6][31] ));
 sg13g2_dfrbp_1 _21756_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net288),
    .D(_00032_),
    .Q_N(_10923_),
    .Q(\TRNG.sha256.expand.dout2[0] ));
 sg13g2_dfrbp_1 _21757_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net289),
    .D(_00043_),
    .Q_N(_10924_),
    .Q(\TRNG.sha256.expand.dout2[1] ));
 sg13g2_dfrbp_1 _21758_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net290),
    .D(_00054_),
    .Q_N(_10925_),
    .Q(\TRNG.sha256.expand.dout2[2] ));
 sg13g2_dfrbp_1 _21759_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net291),
    .D(_00057_),
    .Q_N(_10926_),
    .Q(\TRNG.sha256.expand.dout2[3] ));
 sg13g2_dfrbp_1 _21760_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net292),
    .D(_00058_),
    .Q_N(_10927_),
    .Q(\TRNG.sha256.expand.dout2[4] ));
 sg13g2_dfrbp_1 _21761_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net293),
    .D(_00059_),
    .Q_N(_10928_),
    .Q(\TRNG.sha256.expand.dout2[5] ));
 sg13g2_dfrbp_1 _21762_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net294),
    .D(_00060_),
    .Q_N(_10929_),
    .Q(\TRNG.sha256.expand.dout2[6] ));
 sg13g2_dfrbp_1 _21763_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net295),
    .D(_00061_),
    .Q_N(_10930_),
    .Q(\TRNG.sha256.expand.dout2[7] ));
 sg13g2_dfrbp_1 _21764_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net296),
    .D(_00062_),
    .Q_N(_10931_),
    .Q(\TRNG.sha256.expand.dout2[8] ));
 sg13g2_dfrbp_1 _21765_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net297),
    .D(_00063_),
    .Q_N(_10932_),
    .Q(\TRNG.sha256.expand.dout2[9] ));
 sg13g2_dfrbp_1 _21766_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net298),
    .D(_00033_),
    .Q_N(_10933_),
    .Q(\TRNG.sha256.expand.dout2[10] ));
 sg13g2_dfrbp_1 _21767_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net299),
    .D(_00034_),
    .Q_N(_10934_),
    .Q(\TRNG.sha256.expand.dout2[11] ));
 sg13g2_dfrbp_1 _21768_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net300),
    .D(_00035_),
    .Q_N(_10935_),
    .Q(\TRNG.sha256.expand.dout2[12] ));
 sg13g2_dfrbp_1 _21769_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net301),
    .D(_00036_),
    .Q_N(_10936_),
    .Q(\TRNG.sha256.expand.dout2[13] ));
 sg13g2_dfrbp_1 _21770_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net302),
    .D(_00037_),
    .Q_N(_10937_),
    .Q(\TRNG.sha256.expand.dout2[14] ));
 sg13g2_dfrbp_1 _21771_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net303),
    .D(_00038_),
    .Q_N(_10938_),
    .Q(\TRNG.sha256.expand.dout2[15] ));
 sg13g2_dfrbp_1 _21772_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net304),
    .D(_00039_),
    .Q_N(_10939_),
    .Q(\TRNG.sha256.expand.dout2[16] ));
 sg13g2_dfrbp_1 _21773_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net305),
    .D(_00040_),
    .Q_N(_10940_),
    .Q(\TRNG.sha256.expand.dout2[17] ));
 sg13g2_dfrbp_1 _21774_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net306),
    .D(_00041_),
    .Q_N(_10941_),
    .Q(\TRNG.sha256.expand.dout2[18] ));
 sg13g2_dfrbp_1 _21775_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net307),
    .D(_00042_),
    .Q_N(_10942_),
    .Q(\TRNG.sha256.expand.dout2[19] ));
 sg13g2_dfrbp_1 _21776_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net308),
    .D(_00044_),
    .Q_N(_10943_),
    .Q(\TRNG.sha256.expand.dout2[20] ));
 sg13g2_dfrbp_1 _21777_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net309),
    .D(_00045_),
    .Q_N(_10944_),
    .Q(\TRNG.sha256.expand.dout2[21] ));
 sg13g2_dfrbp_1 _21778_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net310),
    .D(_00046_),
    .Q_N(_10945_),
    .Q(\TRNG.sha256.expand.dout2[22] ));
 sg13g2_dfrbp_1 _21779_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net311),
    .D(_00047_),
    .Q_N(_10946_),
    .Q(\TRNG.sha256.expand.dout2[23] ));
 sg13g2_dfrbp_1 _21780_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net312),
    .D(_00048_),
    .Q_N(_10947_),
    .Q(\TRNG.sha256.expand.dout2[24] ));
 sg13g2_dfrbp_1 _21781_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net313),
    .D(_00049_),
    .Q_N(_10948_),
    .Q(\TRNG.sha256.expand.dout2[25] ));
 sg13g2_dfrbp_1 _21782_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net314),
    .D(_00050_),
    .Q_N(_10949_),
    .Q(\TRNG.sha256.expand.dout2[26] ));
 sg13g2_dfrbp_1 _21783_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net315),
    .D(_00051_),
    .Q_N(_10950_),
    .Q(\TRNG.sha256.expand.dout2[27] ));
 sg13g2_dfrbp_1 _21784_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net316),
    .D(_00052_),
    .Q_N(_10951_),
    .Q(\TRNG.sha256.expand.dout2[28] ));
 sg13g2_dfrbp_1 _21785_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net317),
    .D(_00053_),
    .Q_N(_10952_),
    .Q(\TRNG.sha256.expand.dout2[29] ));
 sg13g2_dfrbp_1 _21786_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net358),
    .D(_00055_),
    .Q_N(_10953_),
    .Q(\TRNG.sha256.expand.dout2[30] ));
 sg13g2_dfrbp_1 _21787_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net651),
    .D(_00056_),
    .Q_N(_10454_),
    .Q(\TRNG.sha256.expand.dout2[31] ));
 sg13g2_dfrbp_1 _21788_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net650),
    .D(_00785_),
    .Q_N(_10453_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][0] ));
 sg13g2_dfrbp_1 _21789_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net649),
    .D(net3030),
    .Q_N(_10452_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][1] ));
 sg13g2_dfrbp_1 _21790_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net648),
    .D(net2524),
    .Q_N(_10451_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][2] ));
 sg13g2_dfrbp_1 _21791_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net647),
    .D(_00788_),
    .Q_N(_10450_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][3] ));
 sg13g2_dfrbp_1 _21792_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net646),
    .D(_00789_),
    .Q_N(_10449_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][4] ));
 sg13g2_dfrbp_1 _21793_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net645),
    .D(_00790_),
    .Q_N(_10448_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][5] ));
 sg13g2_dfrbp_1 _21794_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net644),
    .D(_00791_),
    .Q_N(_10447_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][6] ));
 sg13g2_dfrbp_1 _21795_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net643),
    .D(_00792_),
    .Q_N(_10446_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][7] ));
 sg13g2_dfrbp_1 _21796_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net642),
    .D(_00793_),
    .Q_N(_10445_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][8] ));
 sg13g2_dfrbp_1 _21797_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net641),
    .D(_00794_),
    .Q_N(_10444_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][9] ));
 sg13g2_dfrbp_1 _21798_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net640),
    .D(_00795_),
    .Q_N(_10443_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][10] ));
 sg13g2_dfrbp_1 _21799_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net639),
    .D(_00796_),
    .Q_N(_10442_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][11] ));
 sg13g2_dfrbp_1 _21800_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net638),
    .D(net3036),
    .Q_N(_10441_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][12] ));
 sg13g2_dfrbp_1 _21801_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net637),
    .D(_00798_),
    .Q_N(_10440_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][13] ));
 sg13g2_dfrbp_1 _21802_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net636),
    .D(_00799_),
    .Q_N(_10439_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][14] ));
 sg13g2_dfrbp_1 _21803_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net635),
    .D(net3216),
    .Q_N(_10438_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][15] ));
 sg13g2_dfrbp_1 _21804_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net634),
    .D(_00801_),
    .Q_N(_10437_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][16] ));
 sg13g2_dfrbp_1 _21805_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net633),
    .D(_00802_),
    .Q_N(_10436_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][17] ));
 sg13g2_dfrbp_1 _21806_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net632),
    .D(_00803_),
    .Q_N(_10435_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][18] ));
 sg13g2_dfrbp_1 _21807_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net631),
    .D(_00804_),
    .Q_N(_10434_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][19] ));
 sg13g2_dfrbp_1 _21808_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net630),
    .D(_00805_),
    .Q_N(_10433_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][20] ));
 sg13g2_dfrbp_1 _21809_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net629),
    .D(net2994),
    .Q_N(_10432_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][21] ));
 sg13g2_dfrbp_1 _21810_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net628),
    .D(_00807_),
    .Q_N(_10431_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][22] ));
 sg13g2_dfrbp_1 _21811_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net627),
    .D(_00808_),
    .Q_N(_10430_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][23] ));
 sg13g2_dfrbp_1 _21812_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net626),
    .D(_00809_),
    .Q_N(_10429_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][24] ));
 sg13g2_dfrbp_1 _21813_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net625),
    .D(_00810_),
    .Q_N(_10428_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][25] ));
 sg13g2_dfrbp_1 _21814_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net624),
    .D(_00811_),
    .Q_N(_10427_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][26] ));
 sg13g2_dfrbp_1 _21815_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net623),
    .D(net2747),
    .Q_N(_10426_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][27] ));
 sg13g2_dfrbp_1 _21816_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net622),
    .D(net3060),
    .Q_N(_10425_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][28] ));
 sg13g2_dfrbp_1 _21817_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net621),
    .D(_00814_),
    .Q_N(_10424_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][29] ));
 sg13g2_dfrbp_1 _21818_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net620),
    .D(_00815_),
    .Q_N(_10423_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][30] ));
 sg13g2_dfrbp_1 _21819_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net619),
    .D(_00816_),
    .Q_N(_10422_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[10][31] ));
 sg13g2_dfrbp_1 _21820_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net618),
    .D(net3452),
    .Q_N(_00133_),
    .Q(\TRNG.sha256.control.iteration[6] ));
 sg13g2_dfrbp_1 _21821_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net617),
    .D(net3338),
    .Q_N(_00117_),
    .Q(\TRNG.sha256.control.iteration[8] ));
 sg13g2_dfrbp_1 _21822_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net616),
    .D(net2886),
    .Q_N(_10421_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][0] ));
 sg13g2_dfrbp_1 _21823_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net615),
    .D(net2766),
    .Q_N(_10420_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][1] ));
 sg13g2_dfrbp_1 _21824_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net614),
    .D(_00821_),
    .Q_N(_10419_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][2] ));
 sg13g2_dfrbp_1 _21825_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net613),
    .D(_00822_),
    .Q_N(_10418_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][3] ));
 sg13g2_dfrbp_1 _21826_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net612),
    .D(_00823_),
    .Q_N(_10417_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][4] ));
 sg13g2_dfrbp_1 _21827_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net611),
    .D(_00824_),
    .Q_N(_10416_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][5] ));
 sg13g2_dfrbp_1 _21828_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net610),
    .D(_00825_),
    .Q_N(_10415_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][6] ));
 sg13g2_dfrbp_1 _21829_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net609),
    .D(_00826_),
    .Q_N(_10414_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][7] ));
 sg13g2_dfrbp_1 _21830_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net608),
    .D(_00827_),
    .Q_N(_10413_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][8] ));
 sg13g2_dfrbp_1 _21831_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net607),
    .D(_00828_),
    .Q_N(_10412_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][9] ));
 sg13g2_dfrbp_1 _21832_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net606),
    .D(_00829_),
    .Q_N(_10411_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][10] ));
 sg13g2_dfrbp_1 _21833_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net605),
    .D(_00830_),
    .Q_N(_10410_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][11] ));
 sg13g2_dfrbp_1 _21834_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net604),
    .D(net3018),
    .Q_N(_10409_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][12] ));
 sg13g2_dfrbp_1 _21835_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net603),
    .D(_00832_),
    .Q_N(_10408_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][13] ));
 sg13g2_dfrbp_1 _21836_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net602),
    .D(_00833_),
    .Q_N(_10407_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][14] ));
 sg13g2_dfrbp_1 _21837_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net601),
    .D(net2762),
    .Q_N(_10406_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][15] ));
 sg13g2_dfrbp_1 _21838_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net600),
    .D(_00835_),
    .Q_N(_10405_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][16] ));
 sg13g2_dfrbp_1 _21839_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net599),
    .D(_00836_),
    .Q_N(_10404_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][17] ));
 sg13g2_dfrbp_1 _21840_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net598),
    .D(_00837_),
    .Q_N(_10403_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][18] ));
 sg13g2_dfrbp_1 _21841_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net597),
    .D(_00838_),
    .Q_N(_10402_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][19] ));
 sg13g2_dfrbp_1 _21842_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net596),
    .D(_00839_),
    .Q_N(_10401_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][20] ));
 sg13g2_dfrbp_1 _21843_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net595),
    .D(_00840_),
    .Q_N(_10400_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][21] ));
 sg13g2_dfrbp_1 _21844_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net594),
    .D(_00841_),
    .Q_N(_10399_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][22] ));
 sg13g2_dfrbp_1 _21845_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net593),
    .D(_00842_),
    .Q_N(_10398_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][23] ));
 sg13g2_dfrbp_1 _21846_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net592),
    .D(_00843_),
    .Q_N(_10397_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][24] ));
 sg13g2_dfrbp_1 _21847_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net591),
    .D(_00844_),
    .Q_N(_10396_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][25] ));
 sg13g2_dfrbp_1 _21848_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net590),
    .D(_00845_),
    .Q_N(_10395_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][26] ));
 sg13g2_dfrbp_1 _21849_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net589),
    .D(_00846_),
    .Q_N(_10394_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][27] ));
 sg13g2_dfrbp_1 _21850_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net588),
    .D(_00847_),
    .Q_N(_10393_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][28] ));
 sg13g2_dfrbp_1 _21851_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net587),
    .D(_00848_),
    .Q_N(_10392_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][29] ));
 sg13g2_dfrbp_1 _21852_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net586),
    .D(_00849_),
    .Q_N(_10391_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][30] ));
 sg13g2_dfrbp_1 _21853_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net585),
    .D(_00850_),
    .Q_N(_10390_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[11][31] ));
 sg13g2_dfrbp_1 _21854_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net584),
    .D(_00851_),
    .Q_N(_00118_),
    .Q(\TRNG.sha256.compress.count[4] ));
 sg13g2_dfrbp_1 _21855_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net583),
    .D(_00852_),
    .Q_N(_00275_),
    .Q(\TRNG.sha256.compress.count[0] ));
 sg13g2_dfrbp_1 _21856_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net582),
    .D(_00853_),
    .Q_N(_10389_),
    .Q(\TRNG.sha256.compress.count[1] ));
 sg13g2_dfrbp_1 _21857_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net581),
    .D(_00854_),
    .Q_N(_10388_),
    .Q(\TRNG.sha256.compress.count[2] ));
 sg13g2_dfrbp_1 _21858_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net580),
    .D(_00855_),
    .Q_N(_10387_),
    .Q(\TRNG.sha256.compress.count[3] ));
 sg13g2_dfrbp_1 _21859_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net579),
    .D(net1143),
    .Q_N(_00274_),
    .Q(\TRNG.uart_tx_inst.ticks_counter[0] ));
 sg13g2_dfrbp_1 _21860_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net578),
    .D(net2387),
    .Q_N(_10386_),
    .Q(\TRNG.uart_tx_inst.ticks_counter[1] ));
 sg13g2_dfrbp_1 _21861_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net577),
    .D(net3355),
    .Q_N(_10385_),
    .Q(\TRNG.uart_tx_inst.ticks_counter[2] ));
 sg13g2_dfrbp_1 _21862_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net576),
    .D(_00859_),
    .Q_N(_10384_),
    .Q(\TRNG.uart_tx_inst.ticks_counter[3] ));
 sg13g2_dfrbp_1 _21863_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net575),
    .D(_00860_),
    .Q_N(_10383_),
    .Q(\TRNG.uart_tx_inst.ticks_counter[4] ));
 sg13g2_dfrbp_1 _21864_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net574),
    .D(net3170),
    .Q_N(_10382_),
    .Q(\TRNG.uart_tx_inst.ticks_counter[5] ));
 sg13g2_dfrbp_1 _21865_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net573),
    .D(net2402),
    .Q_N(_10381_),
    .Q(\TRNG.uart_tx_inst.ticks_counter[6] ));
 sg13g2_dfrbp_1 _21866_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net572),
    .D(_00863_),
    .Q_N(_10380_),
    .Q(\TRNG.uart_tx_inst.ticks_counter[7] ));
 sg13g2_dfrbp_1 _21867_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net359),
    .D(_00864_),
    .Q_N(_10954_),
    .Q(\TRNG.uart_tx_inst.ticks_counter[8] ));
 sg13g2_dfrbp_1 _21868_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net360),
    .D(net2484),
    .Q_N(_10955_),
    .Q(\TRNG.uart_tx_inst.tx_reg[0] ));
 sg13g2_dfrbp_1 _21869_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net361),
    .D(net2360),
    .Q_N(_10956_),
    .Q(\TRNG.uart_tx_inst.tx_reg[1] ));
 sg13g2_dfrbp_1 _21870_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net362),
    .D(net2336),
    .Q_N(_10957_),
    .Q(\TRNG.uart_tx_inst.tx_reg[2] ));
 sg13g2_dfrbp_1 _21871_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net363),
    .D(net2327),
    .Q_N(_10958_),
    .Q(\TRNG.uart_tx_inst.tx_reg[3] ));
 sg13g2_dfrbp_1 _21872_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net364),
    .D(net2522),
    .Q_N(_10959_),
    .Q(\TRNG.uart_tx_inst.tx_reg[4] ));
 sg13g2_dfrbp_1 _21873_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net365),
    .D(net2500),
    .Q_N(_10960_),
    .Q(\TRNG.uart_tx_inst.tx_reg[5] ));
 sg13g2_dfrbp_1 _21874_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net366),
    .D(net2260),
    .Q_N(_10961_),
    .Q(\TRNG.uart_tx_inst.tx_reg[6] ));
 sg13g2_dfrbp_1 _21875_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net367),
    .D(net2216),
    .Q_N(_10962_),
    .Q(\TRNG.uart_tx_inst.tx_reg[7] ));
 sg13g2_dfrbp_1 _21876_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net368),
    .D(net1566),
    .Q_N(_00126_),
    .Q(\TRNG.uart_tx_inst.tx_bit_counter[0] ));
 sg13g2_dfrbp_1 _21877_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net369),
    .D(_00103_),
    .Q_N(_00127_),
    .Q(\TRNG.uart_tx_inst.tx_bit_counter[1] ));
 sg13g2_dfrbp_1 _21878_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net452),
    .D(net2194),
    .Q_N(_00128_),
    .Q(\TRNG.uart_tx_inst.tx_bit_counter[2] ));
 sg13g2_dfrbp_1 _21879_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net571),
    .D(net2671),
    .Q_N(_00116_),
    .Q(\TRNG.uart_tx_inst.tx_bit_counter[3] ));
 sg13g2_dfrbp_1 _21880_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net570),
    .D(net2818),
    .Q_N(_10379_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][0] ));
 sg13g2_dfrbp_1 _21881_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net569),
    .D(net2842),
    .Q_N(_10378_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][1] ));
 sg13g2_dfrbp_1 _21882_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net568),
    .D(net2643),
    .Q_N(_10377_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][2] ));
 sg13g2_dfrbp_1 _21883_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net567),
    .D(_00868_),
    .Q_N(_10376_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][3] ));
 sg13g2_dfrbp_1 _21884_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net566),
    .D(_00869_),
    .Q_N(_10375_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][4] ));
 sg13g2_dfrbp_1 _21885_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net565),
    .D(_00870_),
    .Q_N(_10374_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][5] ));
 sg13g2_dfrbp_1 _21886_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net564),
    .D(_00871_),
    .Q_N(_10373_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][6] ));
 sg13g2_dfrbp_1 _21887_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net563),
    .D(_00872_),
    .Q_N(_10372_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][7] ));
 sg13g2_dfrbp_1 _21888_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net562),
    .D(_00873_),
    .Q_N(_10371_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][8] ));
 sg13g2_dfrbp_1 _21889_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net561),
    .D(_00874_),
    .Q_N(_10370_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][9] ));
 sg13g2_dfrbp_1 _21890_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net560),
    .D(_00875_),
    .Q_N(_10369_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][10] ));
 sg13g2_dfrbp_1 _21891_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net559),
    .D(_00876_),
    .Q_N(_10368_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][11] ));
 sg13g2_dfrbp_1 _21892_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net558),
    .D(net2727),
    .Q_N(_10367_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][12] ));
 sg13g2_dfrbp_1 _21893_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net557),
    .D(_00878_),
    .Q_N(_10366_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][13] ));
 sg13g2_dfrbp_1 _21894_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net556),
    .D(_00879_),
    .Q_N(_10365_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][14] ));
 sg13g2_dfrbp_1 _21895_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net555),
    .D(net2673),
    .Q_N(_10364_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][15] ));
 sg13g2_dfrbp_1 _21896_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net554),
    .D(_00881_),
    .Q_N(_10363_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][16] ));
 sg13g2_dfrbp_1 _21897_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net553),
    .D(_00882_),
    .Q_N(_10362_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][17] ));
 sg13g2_dfrbp_1 _21898_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net552),
    .D(_00883_),
    .Q_N(_10361_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][18] ));
 sg13g2_dfrbp_1 _21899_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net551),
    .D(_00884_),
    .Q_N(_10360_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][19] ));
 sg13g2_dfrbp_1 _21900_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net550),
    .D(_00885_),
    .Q_N(_10359_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][20] ));
 sg13g2_dfrbp_1 _21901_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net549),
    .D(_00886_),
    .Q_N(_10358_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][21] ));
 sg13g2_dfrbp_1 _21902_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net548),
    .D(net2602),
    .Q_N(_10357_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][22] ));
 sg13g2_dfrbp_1 _21903_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net451),
    .D(_00888_),
    .Q_N(_10356_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][23] ));
 sg13g2_dfrbp_1 _21904_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net450),
    .D(_00889_),
    .Q_N(_10355_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][24] ));
 sg13g2_dfrbp_1 _21905_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net449),
    .D(_00890_),
    .Q_N(_10354_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][25] ));
 sg13g2_dfrbp_1 _21906_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net448),
    .D(_00891_),
    .Q_N(_10353_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][26] ));
 sg13g2_dfrbp_1 _21907_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net447),
    .D(net2807),
    .Q_N(_10352_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][27] ));
 sg13g2_dfrbp_1 _21908_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net446),
    .D(_00893_),
    .Q_N(_10351_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][28] ));
 sg13g2_dfrbp_1 _21909_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net445),
    .D(_00894_),
    .Q_N(_10350_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][29] ));
 sg13g2_dfrbp_1 _21910_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net444),
    .D(_00895_),
    .Q_N(_10349_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][30] ));
 sg13g2_dfrbp_1 _21911_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net443),
    .D(_00896_),
    .Q_N(_10348_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[9][31] ));
 sg13g2_dfrbp_1 _21912_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net442),
    .D(_00897_),
    .Q_N(_10347_),
    .Q(\TRNG.sha256.W[0] ));
 sg13g2_dfrbp_1 _21913_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net441),
    .D(_00898_),
    .Q_N(_10346_),
    .Q(\TRNG.sha256.W[1] ));
 sg13g2_dfrbp_1 _21914_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net440),
    .D(_00899_),
    .Q_N(_10345_),
    .Q(\TRNG.sha256.W[2] ));
 sg13g2_dfrbp_1 _21915_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net439),
    .D(_00900_),
    .Q_N(_10344_),
    .Q(\TRNG.sha256.W[3] ));
 sg13g2_dfrbp_1 _21916_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net438),
    .D(_00901_),
    .Q_N(_10343_),
    .Q(\TRNG.sha256.W[4] ));
 sg13g2_dfrbp_1 _21917_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net437),
    .D(_00902_),
    .Q_N(_10342_),
    .Q(\TRNG.sha256.W[5] ));
 sg13g2_dfrbp_1 _21918_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net436),
    .D(_00903_),
    .Q_N(_10341_),
    .Q(\TRNG.sha256.W[6] ));
 sg13g2_dfrbp_1 _21919_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net435),
    .D(_00904_),
    .Q_N(_10340_),
    .Q(\TRNG.sha256.W[7] ));
 sg13g2_dfrbp_1 _21920_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net434),
    .D(_00905_),
    .Q_N(_10339_),
    .Q(\TRNG.sha256.W[8] ));
 sg13g2_dfrbp_1 _21921_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net433),
    .D(_00906_),
    .Q_N(_10338_),
    .Q(\TRNG.sha256.W[9] ));
 sg13g2_dfrbp_1 _21922_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net432),
    .D(_00907_),
    .Q_N(_10337_),
    .Q(\TRNG.sha256.W[10] ));
 sg13g2_dfrbp_1 _21923_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net431),
    .D(_00908_),
    .Q_N(_10336_),
    .Q(\TRNG.sha256.W[11] ));
 sg13g2_dfrbp_1 _21924_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net430),
    .D(_00909_),
    .Q_N(_10335_),
    .Q(\TRNG.sha256.W[12] ));
 sg13g2_dfrbp_1 _21925_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net429),
    .D(net3095),
    .Q_N(_10334_),
    .Q(\TRNG.sha256.W[13] ));
 sg13g2_dfrbp_1 _21926_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net428),
    .D(_00911_),
    .Q_N(_10333_),
    .Q(\TRNG.sha256.W[14] ));
 sg13g2_dfrbp_1 _21927_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net427),
    .D(_00912_),
    .Q_N(_10332_),
    .Q(\TRNG.sha256.W[15] ));
 sg13g2_dfrbp_1 _21928_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net426),
    .D(_00913_),
    .Q_N(_10331_),
    .Q(\TRNG.sha256.W[16] ));
 sg13g2_dfrbp_1 _21929_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net425),
    .D(_00914_),
    .Q_N(_10330_),
    .Q(\TRNG.sha256.W[17] ));
 sg13g2_dfrbp_1 _21930_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net424),
    .D(_00915_),
    .Q_N(_10329_),
    .Q(\TRNG.sha256.W[18] ));
 sg13g2_dfrbp_1 _21931_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net423),
    .D(_00916_),
    .Q_N(_10328_),
    .Q(\TRNG.sha256.W[19] ));
 sg13g2_dfrbp_1 _21932_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net422),
    .D(_00917_),
    .Q_N(_10327_),
    .Q(\TRNG.sha256.W[20] ));
 sg13g2_dfrbp_1 _21933_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net421),
    .D(_00918_),
    .Q_N(_10326_),
    .Q(\TRNG.sha256.W[21] ));
 sg13g2_dfrbp_1 _21934_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net420),
    .D(_00919_),
    .Q_N(_10325_),
    .Q(\TRNG.sha256.W[22] ));
 sg13g2_dfrbp_1 _21935_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net419),
    .D(_00920_),
    .Q_N(_10324_),
    .Q(\TRNG.sha256.W[23] ));
 sg13g2_dfrbp_1 _21936_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net418),
    .D(_00921_),
    .Q_N(_10323_),
    .Q(\TRNG.sha256.W[24] ));
 sg13g2_dfrbp_1 _21937_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net417),
    .D(_00922_),
    .Q_N(_10322_),
    .Q(\TRNG.sha256.W[25] ));
 sg13g2_dfrbp_1 _21938_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net416),
    .D(_00923_),
    .Q_N(_10321_),
    .Q(\TRNG.sha256.W[26] ));
 sg13g2_dfrbp_1 _21939_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net415),
    .D(_00924_),
    .Q_N(_10320_),
    .Q(\TRNG.sha256.W[27] ));
 sg13g2_dfrbp_1 _21940_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net414),
    .D(_00925_),
    .Q_N(_10319_),
    .Q(\TRNG.sha256.W[28] ));
 sg13g2_dfrbp_1 _21941_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net413),
    .D(_00926_),
    .Q_N(_10318_),
    .Q(\TRNG.sha256.W[29] ));
 sg13g2_dfrbp_1 _21942_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net412),
    .D(_00927_),
    .Q_N(_10317_),
    .Q(\TRNG.sha256.W[30] ));
 sg13g2_dfrbp_1 _21943_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net411),
    .D(_00928_),
    .Q_N(_10316_),
    .Q(\TRNG.sha256.W[31] ));
 sg13g2_dfrbp_1 _21944_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net410),
    .D(_00929_),
    .Q_N(_10315_),
    .Q(\TRNG.sha256.compress.hash_gen.w_rdy ));
 sg13g2_dfrbp_1 _21945_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net409),
    .D(net3663),
    .Q_N(_10314_),
    .Q(\TRNG.sha256.expand.address1[0] ));
 sg13g2_dfrbp_1 _21946_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net408),
    .D(_00931_),
    .Q_N(_10313_),
    .Q(\TRNG.sha256.expand.address1[1] ));
 sg13g2_dfrbp_1 _21947_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net407),
    .D(net3652),
    .Q_N(_10312_),
    .Q(\TRNG.sha256.expand.address1[2] ));
 sg13g2_dfrbp_1 _21948_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net406),
    .D(net3597),
    .Q_N(_10311_),
    .Q(\TRNG.sha256.expand.address1[3] ));
 sg13g2_dfrbp_1 _21949_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net405),
    .D(_00934_),
    .Q_N(_10310_),
    .Q(\TRNG.sha256.expand.address2[0] ));
 sg13g2_dfrbp_1 _21950_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net404),
    .D(_00935_),
    .Q_N(_10309_),
    .Q(\TRNG.sha256.expand.address2[1] ));
 sg13g2_dfrbp_1 _21951_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net403),
    .D(_00936_),
    .Q_N(_10308_),
    .Q(\TRNG.sha256.expand.address2[2] ));
 sg13g2_dfrbp_1 _21952_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net402),
    .D(_00937_),
    .Q_N(_10307_),
    .Q(\TRNG.sha256.expand.address2[3] ));
 sg13g2_dfrbp_1 _21953_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net401),
    .D(_00938_),
    .Q_N(_10306_),
    .Q(\TRNG.sha256.expand.data1_to_ram[0] ));
 sg13g2_dfrbp_1 _21954_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net400),
    .D(_00939_),
    .Q_N(_10305_),
    .Q(\TRNG.sha256.expand.data1_to_ram[1] ));
 sg13g2_dfrbp_1 _21955_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net399),
    .D(_00940_),
    .Q_N(_10304_),
    .Q(\TRNG.sha256.expand.data1_to_ram[2] ));
 sg13g2_dfrbp_1 _21956_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net398),
    .D(_00941_),
    .Q_N(_10303_),
    .Q(\TRNG.sha256.expand.data1_to_ram[3] ));
 sg13g2_dfrbp_1 _21957_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net397),
    .D(_00942_),
    .Q_N(_10302_),
    .Q(\TRNG.sha256.expand.data1_to_ram[4] ));
 sg13g2_dfrbp_1 _21958_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net396),
    .D(_00943_),
    .Q_N(_10301_),
    .Q(\TRNG.sha256.expand.data1_to_ram[5] ));
 sg13g2_dfrbp_1 _21959_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net395),
    .D(_00944_),
    .Q_N(_10300_),
    .Q(\TRNG.sha256.expand.data1_to_ram[6] ));
 sg13g2_dfrbp_1 _21960_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net394),
    .D(_00945_),
    .Q_N(_10299_),
    .Q(\TRNG.sha256.expand.data1_to_ram[7] ));
 sg13g2_dfrbp_1 _21961_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net393),
    .D(_00946_),
    .Q_N(_10298_),
    .Q(\TRNG.sha256.expand.data1_to_ram[8] ));
 sg13g2_dfrbp_1 _21962_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net392),
    .D(_00947_),
    .Q_N(_10297_),
    .Q(\TRNG.sha256.expand.data1_to_ram[9] ));
 sg13g2_dfrbp_1 _21963_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net391),
    .D(_00948_),
    .Q_N(_10296_),
    .Q(\TRNG.sha256.expand.data1_to_ram[10] ));
 sg13g2_dfrbp_1 _21964_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net390),
    .D(_00949_),
    .Q_N(_10295_),
    .Q(\TRNG.sha256.expand.data1_to_ram[11] ));
 sg13g2_dfrbp_1 _21965_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net389),
    .D(_00950_),
    .Q_N(_10294_),
    .Q(\TRNG.sha256.expand.data1_to_ram[12] ));
 sg13g2_dfrbp_1 _21966_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net388),
    .D(_00951_),
    .Q_N(_10293_),
    .Q(\TRNG.sha256.expand.data1_to_ram[13] ));
 sg13g2_dfrbp_1 _21967_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net387),
    .D(_00952_),
    .Q_N(_10292_),
    .Q(\TRNG.sha256.expand.data1_to_ram[14] ));
 sg13g2_dfrbp_1 _21968_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net386),
    .D(_00953_),
    .Q_N(_10291_),
    .Q(\TRNG.sha256.expand.data1_to_ram[15] ));
 sg13g2_dfrbp_1 _21969_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net385),
    .D(_00954_),
    .Q_N(_10290_),
    .Q(\TRNG.sha256.expand.data1_to_ram[16] ));
 sg13g2_dfrbp_1 _21970_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net384),
    .D(_00955_),
    .Q_N(_10289_),
    .Q(\TRNG.sha256.expand.data1_to_ram[17] ));
 sg13g2_dfrbp_1 _21971_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net383),
    .D(_00956_),
    .Q_N(_10288_),
    .Q(\TRNG.sha256.expand.data1_to_ram[18] ));
 sg13g2_dfrbp_1 _21972_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net382),
    .D(_00957_),
    .Q_N(_10287_),
    .Q(\TRNG.sha256.expand.data1_to_ram[19] ));
 sg13g2_dfrbp_1 _21973_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net381),
    .D(_00958_),
    .Q_N(_10286_),
    .Q(\TRNG.sha256.expand.data1_to_ram[20] ));
 sg13g2_dfrbp_1 _21974_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net380),
    .D(_00959_),
    .Q_N(_10285_),
    .Q(\TRNG.sha256.expand.data1_to_ram[21] ));
 sg13g2_dfrbp_1 _21975_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net379),
    .D(_00960_),
    .Q_N(_10284_),
    .Q(\TRNG.sha256.expand.data1_to_ram[22] ));
 sg13g2_dfrbp_1 _21976_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net378),
    .D(_00961_),
    .Q_N(_10283_),
    .Q(\TRNG.sha256.expand.data1_to_ram[23] ));
 sg13g2_dfrbp_1 _21977_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net377),
    .D(_00962_),
    .Q_N(_10282_),
    .Q(\TRNG.sha256.expand.data1_to_ram[24] ));
 sg13g2_dfrbp_1 _21978_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net376),
    .D(_00963_),
    .Q_N(_10281_),
    .Q(\TRNG.sha256.expand.data1_to_ram[25] ));
 sg13g2_dfrbp_1 _21979_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net375),
    .D(_00964_),
    .Q_N(_10280_),
    .Q(\TRNG.sha256.expand.data1_to_ram[26] ));
 sg13g2_dfrbp_1 _21980_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net374),
    .D(_00965_),
    .Q_N(_10279_),
    .Q(\TRNG.sha256.expand.data1_to_ram[27] ));
 sg13g2_dfrbp_1 _21981_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net373),
    .D(_00966_),
    .Q_N(_10278_),
    .Q(\TRNG.sha256.expand.data1_to_ram[28] ));
 sg13g2_dfrbp_1 _21982_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net372),
    .D(_00967_),
    .Q_N(_10277_),
    .Q(\TRNG.sha256.expand.data1_to_ram[29] ));
 sg13g2_dfrbp_1 _21983_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net371),
    .D(_00968_),
    .Q_N(_10276_),
    .Q(\TRNG.sha256.expand.data1_to_ram[30] ));
 sg13g2_dfrbp_1 _21984_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net370),
    .D(_00969_),
    .Q_N(_10275_),
    .Q(\TRNG.sha256.expand.data1_to_ram[31] ));
 sg13g2_dfrbp_1 _21985_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net357),
    .D(_00970_),
    .Q_N(_10274_),
    .Q(\TRNG.sha256.expand.exp_ctrl.write_en1 ));
 sg13g2_dfrbp_1 _21986_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net356),
    .D(net1137),
    .Q_N(_00273_),
    .Q(\TRNG.sha256.expand.exp_ctrl.j[0] ));
 sg13g2_dfrbp_1 _21987_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net355),
    .D(net2496),
    .Q_N(_10273_),
    .Q(\TRNG.sha256.expand.exp_ctrl.j[1] ));
 sg13g2_dfrbp_1 _21988_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net354),
    .D(_00973_),
    .Q_N(_10272_),
    .Q(\TRNG.sha256.expand.exp_ctrl.j[2] ));
 sg13g2_dfrbp_1 _21989_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net353),
    .D(_00974_),
    .Q_N(_10271_),
    .Q(\TRNG.sha256.expand.exp_ctrl.j[3] ));
 sg13g2_dfrbp_1 _21990_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net352),
    .D(net1181),
    .Q_N(_00272_),
    .Q(\TRNG.sha256.expand.exp_ctrl.j_2[0] ));
 sg13g2_dfrbp_1 _21991_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net351),
    .D(_00976_),
    .Q_N(_10270_),
    .Q(\TRNG.sha256.expand.exp_ctrl.j_2[1] ));
 sg13g2_dfrbp_1 _21992_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net350),
    .D(_00977_),
    .Q_N(_10269_),
    .Q(\TRNG.sha256.expand.exp_ctrl.j_2[2] ));
 sg13g2_dfrbp_1 _21993_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net349),
    .D(net2065),
    .Q_N(_10268_),
    .Q(\TRNG.sha256.expand.exp_ctrl.j_2[3] ));
 sg13g2_dfrbp_1 _21994_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net348),
    .D(net1533),
    .Q_N(_00271_),
    .Q(\TRNG.sha256.expand.exp_ctrl.j_7[0] ));
 sg13g2_dfrbp_1 _21995_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net347),
    .D(_00980_),
    .Q_N(_10267_),
    .Q(\TRNG.sha256.expand.exp_ctrl.j_7[1] ));
 sg13g2_dfrbp_1 _21996_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net346),
    .D(_00981_),
    .Q_N(_10266_),
    .Q(\TRNG.sha256.expand.exp_ctrl.j_7[2] ));
 sg13g2_dfrbp_1 _21997_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net345),
    .D(_00982_),
    .Q_N(_10265_),
    .Q(\TRNG.sha256.expand.exp_ctrl.j_7[3] ));
 sg13g2_dfrbp_1 _21998_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net344),
    .D(net2377),
    .Q_N(_00270_),
    .Q(\TRNG.sha256.expand.exp_ctrl.j_15[0] ));
 sg13g2_dfrbp_1 _21999_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net343),
    .D(net2657),
    .Q_N(_10264_),
    .Q(\TRNG.sha256.expand.exp_ctrl.j_15[1] ));
 sg13g2_dfrbp_1 _22000_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net342),
    .D(_00985_),
    .Q_N(_10263_),
    .Q(\TRNG.sha256.expand.exp_ctrl.j_15[2] ));
 sg13g2_dfrbp_1 _22001_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net341),
    .D(_00986_),
    .Q_N(_10262_),
    .Q(\TRNG.sha256.expand.exp_ctrl.j_15[3] ));
 sg13g2_dfrbp_1 _22002_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net340),
    .D(net2542),
    .Q_N(_10261_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[0] ));
 sg13g2_dfrbp_1 _22003_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net339),
    .D(net2353),
    .Q_N(_10260_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[1] ));
 sg13g2_dfrbp_1 _22004_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net338),
    .D(net2266),
    .Q_N(_10259_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[2] ));
 sg13g2_dfrbp_1 _22005_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net337),
    .D(net2404),
    .Q_N(_10258_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[3] ));
 sg13g2_dfrbp_1 _22006_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net336),
    .D(net2308),
    .Q_N(_10257_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[4] ));
 sg13g2_dfrbp_1 _22007_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net335),
    .D(net2039),
    .Q_N(_10256_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[5] ));
 sg13g2_dfrbp_1 _22008_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net334),
    .D(net2300),
    .Q_N(_10255_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[6] ));
 sg13g2_dfrbp_1 _22009_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net333),
    .D(net2227),
    .Q_N(_10254_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[7] ));
 sg13g2_dfrbp_1 _22010_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net332),
    .D(net2416),
    .Q_N(_10253_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[8] ));
 sg13g2_dfrbp_1 _22011_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net331),
    .D(net2210),
    .Q_N(_10252_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[9] ));
 sg13g2_dfrbp_1 _22012_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net330),
    .D(net2444),
    .Q_N(_10251_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[10] ));
 sg13g2_dfrbp_1 _22013_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net329),
    .D(net2537),
    .Q_N(_10250_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[11] ));
 sg13g2_dfrbp_1 _22014_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net328),
    .D(net2343),
    .Q_N(_10249_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[12] ));
 sg13g2_dfrbp_1 _22015_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net327),
    .D(net2230),
    .Q_N(_10248_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[13] ));
 sg13g2_dfrbp_1 _22016_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net326),
    .D(net2468),
    .Q_N(_10247_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[14] ));
 sg13g2_dfrbp_1 _22017_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net325),
    .D(net2477),
    .Q_N(_10246_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[15] ));
 sg13g2_dfrbp_1 _22018_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net324),
    .D(net2393),
    .Q_N(_10245_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[16] ));
 sg13g2_dfrbp_1 _22019_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net323),
    .D(net2635),
    .Q_N(_10244_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[17] ));
 sg13g2_dfrbp_1 _22020_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net322),
    .D(net2270),
    .Q_N(_10243_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[18] ));
 sg13g2_dfrbp_1 _22021_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net321),
    .D(net2395),
    .Q_N(_10242_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[19] ));
 sg13g2_dfrbp_1 _22022_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net320),
    .D(net1887),
    .Q_N(_10241_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[20] ));
 sg13g2_dfrbp_1 _22023_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net319),
    .D(net2662),
    .Q_N(_10240_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[21] ));
 sg13g2_dfrbp_1 _22024_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net318),
    .D(net1854),
    .Q_N(_10239_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[22] ));
 sg13g2_dfrbp_1 _22025_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net285),
    .D(net2345),
    .Q_N(_10238_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[23] ));
 sg13g2_dfrbp_1 _22026_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net284),
    .D(net2306),
    .Q_N(_10237_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[24] ));
 sg13g2_dfrbp_1 _22027_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net283),
    .D(net2624),
    .Q_N(_10236_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[25] ));
 sg13g2_dfrbp_1 _22028_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net282),
    .D(net2459),
    .Q_N(_10235_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[26] ));
 sg13g2_dfrbp_1 _22029_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net281),
    .D(net2135),
    .Q_N(_10234_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[27] ));
 sg13g2_dfrbp_1 _22030_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net280),
    .D(net2272),
    .Q_N(_10233_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[28] ));
 sg13g2_dfrbp_1 _22031_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net279),
    .D(net1932),
    .Q_N(_10232_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[29] ));
 sg13g2_dfrbp_1 _22032_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net278),
    .D(net2513),
    .Q_N(_10231_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[30] ));
 sg13g2_dfrbp_1 _22033_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net453),
    .D(net2479),
    .Q_N(_10963_),
    .Q(\TRNG.sha256.expand.exp_ctrl.sum[31] ));
 sg13g2_dfrbp_1 _22034_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net454),
    .D(net3485),
    .Q_N(_10964_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[0] ));
 sg13g2_dfrbp_1 _22035_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net455),
    .D(_00277_),
    .Q_N(_10965_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[1] ));
 sg13g2_dfrbp_1 _22036_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net456),
    .D(_00298_),
    .Q_N(_10966_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[2] ));
 sg13g2_dfrbp_1 _22037_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net457),
    .D(_00301_),
    .Q_N(_10967_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[3] ));
 sg13g2_dfrbp_1 _22038_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net458),
    .D(_00302_),
    .Q_N(_10968_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[4] ));
 sg13g2_dfrbp_1 _22039_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net459),
    .D(_00303_),
    .Q_N(_10969_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[5] ));
 sg13g2_dfrbp_1 _22040_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net460),
    .D(_00304_),
    .Q_N(_10970_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[6] ));
 sg13g2_dfrbp_1 _22041_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net461),
    .D(_00305_),
    .Q_N(_10971_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[7] ));
 sg13g2_dfrbp_1 _22042_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net462),
    .D(_00306_),
    .Q_N(_10972_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[8] ));
 sg13g2_dfrbp_1 _22043_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net463),
    .D(_00307_),
    .Q_N(_10973_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[9] ));
 sg13g2_dfrbp_1 _22044_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net464),
    .D(_00278_),
    .Q_N(_10974_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[10] ));
 sg13g2_dfrbp_1 _22045_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net465),
    .D(_00279_),
    .Q_N(_10975_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[11] ));
 sg13g2_dfrbp_1 _22046_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net466),
    .D(_00280_),
    .Q_N(_10976_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[12] ));
 sg13g2_dfrbp_1 _22047_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net467),
    .D(_00281_),
    .Q_N(_10977_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[13] ));
 sg13g2_dfrbp_1 _22048_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net468),
    .D(_00282_),
    .Q_N(_10978_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[14] ));
 sg13g2_dfrbp_1 _22049_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net469),
    .D(_00283_),
    .Q_N(_10979_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[15] ));
 sg13g2_dfrbp_1 _22050_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net470),
    .D(_00284_),
    .Q_N(_10980_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[16] ));
 sg13g2_dfrbp_1 _22051_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net471),
    .D(_00285_),
    .Q_N(_10981_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[17] ));
 sg13g2_dfrbp_1 _22052_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net472),
    .D(_00286_),
    .Q_N(_10982_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[18] ));
 sg13g2_dfrbp_1 _22053_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net473),
    .D(_00287_),
    .Q_N(_10983_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[19] ));
 sg13g2_dfrbp_1 _22054_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net474),
    .D(_00288_),
    .Q_N(_10984_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[20] ));
 sg13g2_dfrbp_1 _22055_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net475),
    .D(_00289_),
    .Q_N(_10985_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[21] ));
 sg13g2_dfrbp_1 _22056_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net476),
    .D(_00290_),
    .Q_N(_10986_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[22] ));
 sg13g2_dfrbp_1 _22057_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net477),
    .D(_00291_),
    .Q_N(_10987_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[23] ));
 sg13g2_dfrbp_1 _22058_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net478),
    .D(_00292_),
    .Q_N(_10988_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[24] ));
 sg13g2_dfrbp_1 _22059_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net479),
    .D(_00293_),
    .Q_N(_10989_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[25] ));
 sg13g2_dfrbp_1 _22060_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net480),
    .D(_00294_),
    .Q_N(_10990_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[26] ));
 sg13g2_dfrbp_1 _22061_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net481),
    .D(_00295_),
    .Q_N(_10991_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[27] ));
 sg13g2_dfrbp_1 _22062_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net482),
    .D(_00296_),
    .Q_N(_10992_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[28] ));
 sg13g2_dfrbp_1 _22063_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net483),
    .D(_00297_),
    .Q_N(_10993_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[29] ));
 sg13g2_dfrbp_1 _22064_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net484),
    .D(_00299_),
    .Q_N(_10994_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[30] ));
 sg13g2_dfrbp_1 _22065_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net485),
    .D(_00300_),
    .Q_N(_10995_),
    .Q(\TRNG.sha256.expand.exp_ctrl.final_sum[31] ));
 sg13g2_dfrbp_1 _22066_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net486),
    .D(_00238_),
    .Q_N(_10996_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[0] ));
 sg13g2_dfrbp_1 _22067_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net487),
    .D(_00249_),
    .Q_N(_10997_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[1] ));
 sg13g2_dfrbp_1 _22068_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net488),
    .D(_00260_),
    .Q_N(_10998_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[2] ));
 sg13g2_dfrbp_1 _22069_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net489),
    .D(_00263_),
    .Q_N(_10999_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[3] ));
 sg13g2_dfrbp_1 _22070_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net490),
    .D(_00264_),
    .Q_N(_11000_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[4] ));
 sg13g2_dfrbp_1 _22071_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net491),
    .D(_00265_),
    .Q_N(_11001_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[5] ));
 sg13g2_dfrbp_1 _22072_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net492),
    .D(_00266_),
    .Q_N(_11002_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[6] ));
 sg13g2_dfrbp_1 _22073_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net493),
    .D(_00267_),
    .Q_N(_11003_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[7] ));
 sg13g2_dfrbp_1 _22074_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net494),
    .D(_00268_),
    .Q_N(_11004_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[8] ));
 sg13g2_dfrbp_1 _22075_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net495),
    .D(_00269_),
    .Q_N(_11005_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[9] ));
 sg13g2_dfrbp_1 _22076_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net496),
    .D(_00239_),
    .Q_N(_11006_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[10] ));
 sg13g2_dfrbp_1 _22077_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net497),
    .D(_00240_),
    .Q_N(_11007_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[11] ));
 sg13g2_dfrbp_1 _22078_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net498),
    .D(_00241_),
    .Q_N(_11008_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[12] ));
 sg13g2_dfrbp_1 _22079_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net499),
    .D(_00242_),
    .Q_N(_11009_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[13] ));
 sg13g2_dfrbp_1 _22080_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net500),
    .D(_00243_),
    .Q_N(_11010_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[14] ));
 sg13g2_dfrbp_1 _22081_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net501),
    .D(_00244_),
    .Q_N(_11011_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[15] ));
 sg13g2_dfrbp_1 _22082_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net502),
    .D(_00245_),
    .Q_N(_11012_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[16] ));
 sg13g2_dfrbp_1 _22083_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net503),
    .D(_00246_),
    .Q_N(_11013_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[17] ));
 sg13g2_dfrbp_1 _22084_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net504),
    .D(_00247_),
    .Q_N(_11014_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[18] ));
 sg13g2_dfrbp_1 _22085_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net505),
    .D(_00248_),
    .Q_N(_11015_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[19] ));
 sg13g2_dfrbp_1 _22086_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net506),
    .D(_00250_),
    .Q_N(_11016_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[20] ));
 sg13g2_dfrbp_1 _22087_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net507),
    .D(_00251_),
    .Q_N(_11017_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[21] ));
 sg13g2_dfrbp_1 _22088_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net508),
    .D(_00252_),
    .Q_N(_11018_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[22] ));
 sg13g2_dfrbp_1 _22089_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net509),
    .D(_00253_),
    .Q_N(_11019_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[23] ));
 sg13g2_dfrbp_1 _22090_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net510),
    .D(_00254_),
    .Q_N(_11020_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[24] ));
 sg13g2_dfrbp_1 _22091_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net511),
    .D(_00255_),
    .Q_N(_11021_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[25] ));
 sg13g2_dfrbp_1 _22092_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net512),
    .D(_00256_),
    .Q_N(_11022_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[26] ));
 sg13g2_dfrbp_1 _22093_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net513),
    .D(_00257_),
    .Q_N(_11023_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[27] ));
 sg13g2_dfrbp_1 _22094_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net514),
    .D(_00258_),
    .Q_N(_11024_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[28] ));
 sg13g2_dfrbp_1 _22095_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net515),
    .D(_00259_),
    .Q_N(_11025_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[29] ));
 sg13g2_dfrbp_1 _22096_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net516),
    .D(_00261_),
    .Q_N(_11026_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[30] ));
 sg13g2_dfrbp_1 _22097_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net517),
    .D(_00262_),
    .Q_N(_11027_),
    .Q(\TRNG.sha256.expand.sm0.sum_0[31] ));
 sg13g2_dfrbp_1 _22098_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net518),
    .D(_00000_),
    .Q_N(_11028_),
    .Q(\TRNG.sha256.K[0] ));
 sg13g2_dfrbp_1 _22099_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net519),
    .D(_00011_),
    .Q_N(_11029_),
    .Q(\TRNG.sha256.K[1] ));
 sg13g2_dfrbp_1 _22100_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net520),
    .D(_00022_),
    .Q_N(_11030_),
    .Q(\TRNG.sha256.K[2] ));
 sg13g2_dfrbp_1 _22101_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net521),
    .D(_00025_),
    .Q_N(_11031_),
    .Q(\TRNG.sha256.K[3] ));
 sg13g2_dfrbp_1 _22102_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net522),
    .D(_00026_),
    .Q_N(_11032_),
    .Q(\TRNG.sha256.K[4] ));
 sg13g2_dfrbp_1 _22103_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net523),
    .D(_00027_),
    .Q_N(_11033_),
    .Q(\TRNG.sha256.K[5] ));
 sg13g2_dfrbp_1 _22104_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net524),
    .D(_00028_),
    .Q_N(_11034_),
    .Q(\TRNG.sha256.K[6] ));
 sg13g2_dfrbp_1 _22105_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net525),
    .D(_00029_),
    .Q_N(_11035_),
    .Q(\TRNG.sha256.K[7] ));
 sg13g2_dfrbp_1 _22106_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net526),
    .D(_00030_),
    .Q_N(_11036_),
    .Q(\TRNG.sha256.K[8] ));
 sg13g2_dfrbp_1 _22107_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net527),
    .D(_00031_),
    .Q_N(_11037_),
    .Q(\TRNG.sha256.K[9] ));
 sg13g2_dfrbp_1 _22108_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net528),
    .D(_00001_),
    .Q_N(_11038_),
    .Q(\TRNG.sha256.K[10] ));
 sg13g2_dfrbp_1 _22109_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net529),
    .D(_00002_),
    .Q_N(_11039_),
    .Q(\TRNG.sha256.K[11] ));
 sg13g2_dfrbp_1 _22110_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net530),
    .D(_00003_),
    .Q_N(_11040_),
    .Q(\TRNG.sha256.K[12] ));
 sg13g2_dfrbp_1 _22111_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net531),
    .D(_00004_),
    .Q_N(_11041_),
    .Q(\TRNG.sha256.K[13] ));
 sg13g2_dfrbp_1 _22112_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net532),
    .D(_00005_),
    .Q_N(_11042_),
    .Q(\TRNG.sha256.K[14] ));
 sg13g2_dfrbp_1 _22113_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net533),
    .D(_00006_),
    .Q_N(_11043_),
    .Q(\TRNG.sha256.K[15] ));
 sg13g2_dfrbp_1 _22114_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net534),
    .D(_00007_),
    .Q_N(_11044_),
    .Q(\TRNG.sha256.K[16] ));
 sg13g2_dfrbp_1 _22115_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net535),
    .D(_00008_),
    .Q_N(_11045_),
    .Q(\TRNG.sha256.K[17] ));
 sg13g2_dfrbp_1 _22116_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net536),
    .D(_00009_),
    .Q_N(_11046_),
    .Q(\TRNG.sha256.K[18] ));
 sg13g2_dfrbp_1 _22117_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net537),
    .D(_00010_),
    .Q_N(_11047_),
    .Q(\TRNG.sha256.K[19] ));
 sg13g2_dfrbp_1 _22118_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net538),
    .D(_00012_),
    .Q_N(_11048_),
    .Q(\TRNG.sha256.K[20] ));
 sg13g2_dfrbp_1 _22119_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net539),
    .D(_00013_),
    .Q_N(_11049_),
    .Q(\TRNG.sha256.K[21] ));
 sg13g2_dfrbp_1 _22120_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net540),
    .D(_00014_),
    .Q_N(_11050_),
    .Q(\TRNG.sha256.K[22] ));
 sg13g2_dfrbp_1 _22121_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net541),
    .D(_00015_),
    .Q_N(_11051_),
    .Q(\TRNG.sha256.K[23] ));
 sg13g2_dfrbp_1 _22122_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net542),
    .D(_00016_),
    .Q_N(_11052_),
    .Q(\TRNG.sha256.K[24] ));
 sg13g2_dfrbp_1 _22123_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net543),
    .D(_00017_),
    .Q_N(_11053_),
    .Q(\TRNG.sha256.K[25] ));
 sg13g2_dfrbp_1 _22124_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net544),
    .D(_00018_),
    .Q_N(_11054_),
    .Q(\TRNG.sha256.K[26] ));
 sg13g2_dfrbp_1 _22125_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net545),
    .D(_00019_),
    .Q_N(_11055_),
    .Q(\TRNG.sha256.K[27] ));
 sg13g2_dfrbp_1 _22126_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net546),
    .D(_00020_),
    .Q_N(_11056_),
    .Q(\TRNG.sha256.K[28] ));
 sg13g2_dfrbp_1 _22127_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net547),
    .D(_00021_),
    .Q_N(_11057_),
    .Q(\TRNG.sha256.K[29] ));
 sg13g2_dfrbp_1 _22128_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net753),
    .D(_00023_),
    .Q_N(_11058_),
    .Q(\TRNG.sha256.K[30] ));
 sg13g2_dfrbp_1 _22129_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net277),
    .D(_00024_),
    .Q_N(_10230_),
    .Q(\TRNG.sha256.K[31] ));
 sg13g2_dfrbp_1 _22130_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net276),
    .D(net2596),
    .Q_N(_10229_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][0] ));
 sg13g2_dfrbp_1 _22131_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net275),
    .D(net2608),
    .Q_N(_10228_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][1] ));
 sg13g2_dfrbp_1 _22132_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net274),
    .D(_01021_),
    .Q_N(_10227_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][2] ));
 sg13g2_dfrbp_1 _22133_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net273),
    .D(net2859),
    .Q_N(_10226_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][3] ));
 sg13g2_dfrbp_1 _22134_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net272),
    .D(_01023_),
    .Q_N(_10225_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][4] ));
 sg13g2_dfrbp_1 _22135_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net271),
    .D(_01024_),
    .Q_N(_10224_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][5] ));
 sg13g2_dfrbp_1 _22136_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net270),
    .D(_01025_),
    .Q_N(_10223_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][6] ));
 sg13g2_dfrbp_1 _22137_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net269),
    .D(_01026_),
    .Q_N(_10222_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][7] ));
 sg13g2_dfrbp_1 _22138_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net268),
    .D(_01027_),
    .Q_N(_10221_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][8] ));
 sg13g2_dfrbp_1 _22139_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net267),
    .D(_01028_),
    .Q_N(_10220_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][9] ));
 sg13g2_dfrbp_1 _22140_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net266),
    .D(_01029_),
    .Q_N(_10219_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][10] ));
 sg13g2_dfrbp_1 _22141_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net265),
    .D(_01030_),
    .Q_N(_10218_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][11] ));
 sg13g2_dfrbp_1 _22142_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net264),
    .D(_01031_),
    .Q_N(_10217_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][12] ));
 sg13g2_dfrbp_1 _22143_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net263),
    .D(_01032_),
    .Q_N(_10216_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][13] ));
 sg13g2_dfrbp_1 _22144_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net262),
    .D(_01033_),
    .Q_N(_10215_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][14] ));
 sg13g2_dfrbp_1 _22145_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net261),
    .D(_01034_),
    .Q_N(_10214_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][15] ));
 sg13g2_dfrbp_1 _22146_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net260),
    .D(_01035_),
    .Q_N(_10213_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][16] ));
 sg13g2_dfrbp_1 _22147_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net259),
    .D(_01036_),
    .Q_N(_10212_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][17] ));
 sg13g2_dfrbp_1 _22148_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net258),
    .D(_01037_),
    .Q_N(_10211_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][18] ));
 sg13g2_dfrbp_1 _22149_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net257),
    .D(_01038_),
    .Q_N(_10210_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][19] ));
 sg13g2_dfrbp_1 _22150_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net256),
    .D(_01039_),
    .Q_N(_10209_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][20] ));
 sg13g2_dfrbp_1 _22151_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net255),
    .D(_01040_),
    .Q_N(_10208_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][21] ));
 sg13g2_dfrbp_1 _22152_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net254),
    .D(_01041_),
    .Q_N(_10207_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][22] ));
 sg13g2_dfrbp_1 _22153_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net253),
    .D(_01042_),
    .Q_N(_10206_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][23] ));
 sg13g2_dfrbp_1 _22154_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net252),
    .D(_01043_),
    .Q_N(_10205_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][24] ));
 sg13g2_dfrbp_1 _22155_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net251),
    .D(_01044_),
    .Q_N(_10204_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][25] ));
 sg13g2_dfrbp_1 _22156_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net250),
    .D(_01045_),
    .Q_N(_10203_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][26] ));
 sg13g2_dfrbp_1 _22157_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net249),
    .D(net2570),
    .Q_N(_10202_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][27] ));
 sg13g2_dfrbp_1 _22158_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net248),
    .D(_01047_),
    .Q_N(_10201_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][28] ));
 sg13g2_dfrbp_1 _22159_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net247),
    .D(_01048_),
    .Q_N(_10200_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][29] ));
 sg13g2_dfrbp_1 _22160_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net246),
    .D(_01049_),
    .Q_N(_10199_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][30] ));
 sg13g2_dfrbp_1 _22161_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net245),
    .D(_01050_),
    .Q_N(_10198_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[12][31] ));
 sg13g2_dfrbp_1 _22162_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net244),
    .D(_01051_),
    .Q_N(_10197_),
    .Q(\TRNG.sha256.compress.done ));
 sg13g2_dfrbp_1 _22163_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net243),
    .D(_01052_),
    .Q_N(_00131_),
    .Q(\TRNG.sha256.connect[0] ));
 sg13g2_dfrbp_1 _22164_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net242),
    .D(_01053_),
    .Q_N(_00132_),
    .Q(\TRNG.sha256.connect[1] ));
 sg13g2_dfrbp_1 _22165_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net241),
    .D(_01054_),
    .Q_N(_00130_),
    .Q(\TRNG.sha256.connect[2] ));
 sg13g2_dfrbp_1 _22166_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net240),
    .D(_01055_),
    .Q_N(_10196_),
    .Q(\TRNG.sha256.connect[3] ));
 sg13g2_dfrbp_1 _22167_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net239),
    .D(_01056_),
    .Q_N(_00129_),
    .Q(\TRNG.sha256.connect[4] ));
 sg13g2_dfrbp_1 _22168_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net238),
    .D(_01057_),
    .Q_N(_10195_),
    .Q(\TRNG.sha256.connect[5] ));
 sg13g2_dfrbp_1 _22169_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net237),
    .D(_01058_),
    .Q_N(_10194_),
    .Q(\TRNG.sha256.control.iteration[7] ));
 sg13g2_dfrbp_1 _22170_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net236),
    .D(_01059_),
    .Q_N(_10193_),
    .Q(\TRNG.sha256.compress.hash_gen.temp[1] ));
 sg13g2_dfrbp_1 _22171_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net235),
    .D(_01060_),
    .Q_N(_10192_),
    .Q(\TRNG.sha256.compress.hash_gen.temp[2] ));
 sg13g2_dfrbp_1 _22172_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net234),
    .D(_01061_),
    .Q_N(_10191_),
    .Q(\TRNG.sha256.compress.hash_gen.temp[3] ));
 sg13g2_dfrbp_1 _22173_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net233),
    .D(_01062_),
    .Q_N(_10190_),
    .Q(\TRNG.sha256.compress.hash_gen.temp[4] ));
 sg13g2_dfrbp_1 _22174_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net232),
    .D(_01063_),
    .Q_N(_00146_),
    .Q(\TRNG.hash[129] ));
 sg13g2_dfrbp_1 _22175_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net231),
    .D(net3631),
    .Q_N(_00147_),
    .Q(\TRNG.hash[131] ));
 sg13g2_dfrbp_1 _22176_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net230),
    .D(net3853),
    .Q_N(_10189_),
    .Q(\TRNG.hash[132] ));
 sg13g2_dfrbp_1 _22177_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net229),
    .D(net3644),
    .Q_N(_00135_),
    .Q(\TRNG.hash[133] ));
 sg13g2_dfrbp_1 _22178_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net228),
    .D(net3516),
    .Q_N(_00148_),
    .Q(\TRNG.hash[136] ));
 sg13g2_dfrbp_1 _22179_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net227),
    .D(net3666),
    .Q_N(_00136_),
    .Q(\TRNG.hash[138] ));
 sg13g2_dfrbp_1 _22180_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net226),
    .D(_01069_),
    .Q_N(_00138_),
    .Q(\TRNG.hash[140] ));
 sg13g2_dfrbp_1 _22181_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net225),
    .D(net3466),
    .Q_N(_00207_),
    .Q(\TRNG.hash[141] ));
 sg13g2_dfrbp_1 _22182_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net224),
    .D(net3843),
    .Q_N(_10188_),
    .Q(\TRNG.hash[142] ));
 sg13g2_dfrbp_1 _22183_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net223),
    .D(_01072_),
    .Q_N(_10187_),
    .Q(\TRNG.hash[143] ));
 sg13g2_dfrbp_1 _22184_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net222),
    .D(_01073_),
    .Q_N(_10186_),
    .Q(\TRNG.hash[144] ));
 sg13g2_dfrbp_1 _22185_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net221),
    .D(net3676),
    .Q_N(_10185_),
    .Q(\TRNG.hash[145] ));
 sg13g2_dfrbp_1 _22186_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net220),
    .D(net3535),
    .Q_N(_10184_),
    .Q(\TRNG.hash[146] ));
 sg13g2_dfrbp_1 _22187_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net219),
    .D(net3656),
    .Q_N(_10183_),
    .Q(\TRNG.hash[147] ));
 sg13g2_dfrbp_1 _22188_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net218),
    .D(net3646),
    .Q_N(_00140_),
    .Q(\TRNG.hash[150] ));
 sg13g2_dfrbp_1 _22189_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net217),
    .D(_01078_),
    .Q_N(_00141_),
    .Q(\TRNG.hash[152] ));
 sg13g2_dfrbp_1 _22190_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net216),
    .D(_01079_),
    .Q_N(_00143_),
    .Q(\TRNG.hash[154] ));
 sg13g2_dfrbp_1 _22191_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net215),
    .D(_01080_),
    .Q_N(_00145_),
    .Q(\TRNG.hash[157] ));
 sg13g2_dfrbp_1 _22192_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net214),
    .D(_01081_),
    .Q_N(_10182_),
    .Q(\TRNG.hash[159] ));
 sg13g2_dfrbp_1 _22193_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net5901),
    .D(_01082_),
    .Q_N(_10181_),
    .Q(\TRNG.Repetition_Count_Test.prev_bit ));
 sg13g2_dfrbp_1 _22194_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net213),
    .D(_01083_),
    .Q_N(_10180_),
    .Q(\TRNG.hash_rdy ));
 sg13g2_dfrbp_1 _22195_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net212),
    .D(_01084_),
    .Q_N(_00228_),
    .Q(\TRNG.hash[224] ));
 sg13g2_dfrbp_1 _22196_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net211),
    .D(_01085_),
    .Q_N(_10179_),
    .Q(\TRNG.hash[225] ));
 sg13g2_dfrbp_1 _22197_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net210),
    .D(_01086_),
    .Q_N(_10178_),
    .Q(\TRNG.hash[226] ));
 sg13g2_dfrbp_1 _22198_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net209),
    .D(_01087_),
    .Q_N(_00231_),
    .Q(\TRNG.hash[229] ));
 sg13g2_dfrbp_1 _22199_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net208),
    .D(_01088_),
    .Q_N(_10177_),
    .Q(\TRNG.hash[230] ));
 sg13g2_dfrbp_1 _22200_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net207),
    .D(_01089_),
    .Q_N(_00232_),
    .Q(\TRNG.hash[233] ));
 sg13g2_dfrbp_1 _22201_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net206),
    .D(_01090_),
    .Q_N(_10176_),
    .Q(\TRNG.hash[234] ));
 sg13g2_dfrbp_1 _22202_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net205),
    .D(_01091_),
    .Q_N(_00237_),
    .Q(\TRNG.hash[237] ));
 sg13g2_dfrbp_1 _22203_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net204),
    .D(_01092_),
    .Q_N(_10175_),
    .Q(\TRNG.hash[238] ));
 sg13g2_dfrbp_1 _22204_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net203),
    .D(_01093_),
    .Q_N(_10174_),
    .Q(\TRNG.hash[239] ));
 sg13g2_dfrbp_1 _22205_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net202),
    .D(_01094_),
    .Q_N(_10173_),
    .Q(\TRNG.hash[240] ));
 sg13g2_dfrbp_1 _22206_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net201),
    .D(net3796),
    .Q_N(_00233_),
    .Q(\TRNG.hash[243] ));
 sg13g2_dfrbp_1 _22207_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net200),
    .D(net3742),
    .Q_N(_00234_),
    .Q(\TRNG.hash[249] ));
 sg13g2_dfrbp_1 _22208_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net199),
    .D(_01097_),
    .Q_N(_00235_),
    .Q(\TRNG.hash[251] ));
 sg13g2_dfrbp_1 _22209_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net198),
    .D(net3789),
    .Q_N(_00236_),
    .Q(\TRNG.hash[253] ));
 sg13g2_dfrbp_1 _22210_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net197),
    .D(_01099_),
    .Q_N(_10172_),
    .Q(\TRNG.hash[254] ));
 sg13g2_dfrbp_1 _22211_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net196),
    .D(_01100_),
    .Q_N(_10171_),
    .Q(\TRNG.hash[192] ));
 sg13g2_dfrbp_1 _22212_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net195),
    .D(_01101_),
    .Q_N(_10170_),
    .Q(\TRNG.hash[194] ));
 sg13g2_dfrbp_1 _22213_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net194),
    .D(_01102_),
    .Q_N(_10169_),
    .Q(\TRNG.hash[199] ));
 sg13g2_dfrbp_1 _22214_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net193),
    .D(net3475),
    .Q_N(_00229_),
    .Q(\TRNG.hash[201] ));
 sg13g2_dfrbp_1 _22215_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net192),
    .D(_01104_),
    .Q_N(_10168_),
    .Q(\TRNG.hash[202] ));
 sg13g2_dfrbp_1 _22216_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net191),
    .D(_01105_),
    .Q_N(_10167_),
    .Q(\TRNG.hash[203] ));
 sg13g2_dfrbp_1 _22217_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net190),
    .D(net3438),
    .Q_N(_00225_),
    .Q(\TRNG.hash[205] ));
 sg13g2_dfrbp_1 _22218_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net189),
    .D(_01107_),
    .Q_N(_10166_),
    .Q(\TRNG.hash[207] ));
 sg13g2_dfrbp_1 _22219_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net188),
    .D(net3637),
    .Q_N(_00230_),
    .Q(\TRNG.hash[208] ));
 sg13g2_dfrbp_1 _22220_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net187),
    .D(_01109_),
    .Q_N(_10165_),
    .Q(\TRNG.hash[209] ));
 sg13g2_dfrbp_1 _22221_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net186),
    .D(_01110_),
    .Q_N(_10164_),
    .Q(\TRNG.hash[210] ));
 sg13g2_dfrbp_1 _22222_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net185),
    .D(net3531),
    .Q_N(_00226_),
    .Q(\TRNG.hash[213] ));
 sg13g2_dfrbp_1 _22223_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net184),
    .D(_01112_),
    .Q_N(_10163_),
    .Q(\TRNG.hash[214] ));
 sg13g2_dfrbp_1 _22224_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net183),
    .D(net3787),
    .Q_N(_10162_),
    .Q(\TRNG.hash[216] ));
 sg13g2_dfrbp_1 _22225_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net182),
    .D(_01114_),
    .Q_N(_10161_),
    .Q(\TRNG.hash[217] ));
 sg13g2_dfrbp_1 _22226_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net181),
    .D(net3477),
    .Q_N(_00227_),
    .Q(\TRNG.hash[219] ));
 sg13g2_dfrbp_1 _22227_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net180),
    .D(_01116_),
    .Q_N(_10160_),
    .Q(\TRNG.hash[220] ));
 sg13g2_dfrbp_1 _22228_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net179),
    .D(_01117_),
    .Q_N(_10159_),
    .Q(\TRNG.hash[221] ));
 sg13g2_dfrbp_1 _22229_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net178),
    .D(_01118_),
    .Q_N(_10158_),
    .Q(\TRNG.hash[223] ));
 sg13g2_dfrbp_1 _22230_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net177),
    .D(_01119_),
    .Q_N(_00222_),
    .Q(\TRNG.hash[161] ));
 sg13g2_dfrbp_1 _22231_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net176),
    .D(net3504),
    .Q_N(_00221_),
    .Q(\TRNG.hash[164] ));
 sg13g2_dfrbp_1 _22232_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net175),
    .D(net3730),
    .Q_N(_10157_),
    .Q(\TRNG.hash[165] ));
 sg13g2_dfrbp_1 _22233_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net174),
    .D(_01122_),
    .Q_N(_10156_),
    .Q(\TRNG.hash[166] ));
 sg13g2_dfrbp_1 _22234_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net173),
    .D(_01123_),
    .Q_N(_10155_),
    .Q(\TRNG.hash[168] ));
 sg13g2_dfrbp_1 _22235_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net172),
    .D(_01124_),
    .Q_N(_10154_),
    .Q(\TRNG.hash[169] ));
 sg13g2_dfrbp_1 _22236_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net171),
    .D(_01125_),
    .Q_N(_10153_),
    .Q(\TRNG.hash[172] ));
 sg13g2_dfrbp_1 _22237_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net170),
    .D(_01126_),
    .Q_N(_10152_),
    .Q(\TRNG.hash[173] ));
 sg13g2_dfrbp_1 _22238_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net169),
    .D(_01127_),
    .Q_N(_10151_),
    .Q(\TRNG.hash[174] ));
 sg13g2_dfrbp_1 _22239_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net168),
    .D(_01128_),
    .Q_N(_10150_),
    .Q(\TRNG.hash[175] ));
 sg13g2_dfrbp_1 _22240_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net167),
    .D(net3685),
    .Q_N(_00223_),
    .Q(\TRNG.hash[177] ));
 sg13g2_dfrbp_1 _22241_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net166),
    .D(_01130_),
    .Q_N(_10149_),
    .Q(\TRNG.hash[178] ));
 sg13g2_dfrbp_1 _22242_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net165),
    .D(_01131_),
    .Q_N(_10148_),
    .Q(\TRNG.hash[179] ));
 sg13g2_dfrbp_1 _22243_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net164),
    .D(_01132_),
    .Q_N(_10147_),
    .Q(\TRNG.hash[181] ));
 sg13g2_dfrbp_1 _22244_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net163),
    .D(net3785),
    .Q_N(_10146_),
    .Q(\TRNG.hash[182] ));
 sg13g2_dfrbp_1 _22245_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net162),
    .D(net3496),
    .Q_N(_00224_),
    .Q(\TRNG.hash[186] ));
 sg13g2_dfrbp_1 _22246_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net161),
    .D(net3869),
    .Q_N(_10145_),
    .Q(\TRNG.hash[187] ));
 sg13g2_dfrbp_1 _22247_ (.CLK(clknet_6_17_0_clk),
    .RESET_B(net160),
    .D(_01136_),
    .Q_N(_10144_),
    .Q(\TRNG.hash[188] ));
 sg13g2_dfrbp_1 _22248_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net159),
    .D(net3831),
    .Q_N(_10143_),
    .Q(\TRNG.hash[189] ));
 sg13g2_dfrbp_1 _22249_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net158),
    .D(_01138_),
    .Q_N(_10142_),
    .Q(\TRNG.hash[96] ));
 sg13g2_dfrbp_1 _22250_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net157),
    .D(_01139_),
    .Q_N(_10141_),
    .Q(\TRNG.hash[97] ));
 sg13g2_dfrbp_1 _22251_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net156),
    .D(_01140_),
    .Q_N(_10140_),
    .Q(\TRNG.hash[98] ));
 sg13g2_dfrbp_1 _22252_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net155),
    .D(_01141_),
    .Q_N(_10139_),
    .Q(\TRNG.hash[99] ));
 sg13g2_dfrbp_1 _22253_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net154),
    .D(_01142_),
    .Q_N(_10138_),
    .Q(\TRNG.hash[100] ));
 sg13g2_dfrbp_1 _22254_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net153),
    .D(_01143_),
    .Q_N(_10137_),
    .Q(\TRNG.hash[101] ));
 sg13g2_dfrbp_1 _22255_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net152),
    .D(_01144_),
    .Q_N(_10136_),
    .Q(\TRNG.hash[102] ));
 sg13g2_dfrbp_1 _22256_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net151),
    .D(net3752),
    .Q_N(_00206_),
    .Q(\TRNG.hash[105] ));
 sg13g2_dfrbp_1 _22257_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net150),
    .D(net3552),
    .Q_N(_00208_),
    .Q(\TRNG.hash[108] ));
 sg13g2_dfrbp_1 _22258_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net149),
    .D(_01147_),
    .Q_N(_10135_),
    .Q(\TRNG.hash[110] ));
 sg13g2_dfrbp_1 _22259_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net148),
    .D(net3715),
    .Q_N(_00220_),
    .Q(\TRNG.hash[113] ));
 sg13g2_dfrbp_1 _22260_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net147),
    .D(_01149_),
    .Q_N(_10134_),
    .Q(\TRNG.hash[114] ));
 sg13g2_dfrbp_1 _22261_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net146),
    .D(_01150_),
    .Q_N(_10133_),
    .Q(\TRNG.hash[115] ));
 sg13g2_dfrbp_1 _22262_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net145),
    .D(_01151_),
    .Q_N(_00215_),
    .Q(\TRNG.hash[120] ));
 sg13g2_dfrbp_1 _22263_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net144),
    .D(_01152_),
    .Q_N(_00200_),
    .Q(\TRNG.hash[124] ));
 sg13g2_dfrbp_1 _22264_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net143),
    .D(_01153_),
    .Q_N(_10132_),
    .Q(\TRNG.hash[126] ));
 sg13g2_dfrbp_1 _22265_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net142),
    .D(_01154_),
    .Q_N(_00191_),
    .Q(\TRNG.hash[66] ));
 sg13g2_dfrbp_1 _22266_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net141),
    .D(net3836),
    .Q_N(_10131_),
    .Q(\TRNG.hash[67] ));
 sg13g2_dfrbp_1 _22267_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net140),
    .D(_01156_),
    .Q_N(_00180_),
    .Q(\TRNG.hash[71] ));
 sg13g2_dfrbp_1 _22268_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net139),
    .D(net3436),
    .Q_N(_00182_),
    .Q(\TRNG.hash[75] ));
 sg13g2_dfrbp_1 _22269_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net138),
    .D(net3448),
    .Q_N(_00194_),
    .Q(\TRNG.hash[77] ));
 sg13g2_dfrbp_1 _22270_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net137),
    .D(net3605),
    .Q_N(_00184_),
    .Q(\TRNG.hash[78] ));
 sg13g2_dfrbp_1 _22271_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net136),
    .D(net3554),
    .Q_N(_00185_),
    .Q(\TRNG.hash[80] ));
 sg13g2_dfrbp_1 _22272_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net135),
    .D(net3456),
    .Q_N(_00195_),
    .Q(\TRNG.hash[82] ));
 sg13g2_dfrbp_1 _22273_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net134),
    .D(net3668),
    .Q_N(_00196_),
    .Q(\TRNG.hash[88] ));
 sg13g2_dfrbp_1 _22274_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net133),
    .D(_01163_),
    .Q_N(_00217_),
    .Q(\TRNG.hash[89] ));
 sg13g2_dfrbp_1 _22275_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net132),
    .D(_01164_),
    .Q_N(_00190_),
    .Q(\TRNG.hash[91] ));
 sg13g2_dfrbp_1 _22276_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net131),
    .D(net3822),
    .Q_N(_10130_),
    .Q(\TRNG.hash[92] ));
 sg13g2_dfrbp_1 _22277_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net130),
    .D(net3389),
    .Q_N(_00197_),
    .Q(\TRNG.hash[95] ));
 sg13g2_dfrbp_1 _22278_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net129),
    .D(net3758),
    .Q_N(_00155_),
    .Q(\TRNG.hash[32] ));
 sg13g2_dfrbp_1 _22279_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net128),
    .D(_01168_),
    .Q_N(_10129_),
    .Q(\TRNG.hash[33] ));
 sg13g2_dfrbp_1 _22280_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net127),
    .D(net3538),
    .Q_N(_00162_),
    .Q(\TRNG.hash[35] ));
 sg13g2_dfrbp_1 _22281_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net126),
    .D(net3771),
    .Q_N(_00164_),
    .Q(\TRNG.hash[37] ));
 sg13g2_dfrbp_1 _22282_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net125),
    .D(_01171_),
    .Q_N(_00173_),
    .Q(\TRNG.hash[39] ));
 sg13g2_dfrbp_1 _22283_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net124),
    .D(_01172_),
    .Q_N(_00174_),
    .Q(\TRNG.hash[40] ));
 sg13g2_dfrbp_1 _22284_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net123),
    .D(net3586),
    .Q_N(_00175_),
    .Q(\TRNG.hash[43] ));
 sg13g2_dfrbp_1 _22285_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net122),
    .D(net3595),
    .Q_N(_00167_),
    .Q(\TRNG.hash[44] ));
 sg13g2_dfrbp_1 _22286_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net121),
    .D(_01175_),
    .Q_N(_10128_),
    .Q(\TRNG.hash[46] ));
 sg13g2_dfrbp_1 _22287_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net120),
    .D(net3607),
    .Q_N(_00210_),
    .Q(\TRNG.hash[47] ));
 sg13g2_dfrbp_1 _22288_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net119),
    .D(net3527),
    .Q_N(_00176_),
    .Q(\TRNG.hash[48] ));
 sg13g2_dfrbp_1 _22289_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net118),
    .D(net3680),
    .Q_N(_10127_),
    .Q(\TRNG.hash[49] ));
 sg13g2_dfrbp_1 _22290_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net117),
    .D(_01179_),
    .Q_N(_00172_),
    .Q(\TRNG.hash[55] ));
 sg13g2_dfrbp_1 _22291_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net116),
    .D(net3804),
    .Q_N(_10126_),
    .Q(\TRNG.hash[56] ));
 sg13g2_dfrbp_1 _22292_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net115),
    .D(_01181_),
    .Q_N(_00216_),
    .Q(\TRNG.hash[57] ));
 sg13g2_dfrbp_1 _22293_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net114),
    .D(_01182_),
    .Q_N(_00218_),
    .Q(\TRNG.hash[58] ));
 sg13g2_dfrbp_1 _22294_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net112),
    .D(_01183_),
    .Q_N(_00219_),
    .Q(\TRNG.hash[59] ));
 sg13g2_dfrbp_1 _22295_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net111),
    .D(net3635),
    .Q_N(_00171_),
    .Q(\TRNG.hash[60] ));
 sg13g2_dfrbp_1 _22296_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net110),
    .D(_01185_),
    .Q_N(_10125_),
    .Q(\TRNG.hash[0] ));
 sg13g2_dfrbp_1 _22297_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net109),
    .D(net3557),
    .Q_N(_00156_),
    .Q(\TRNG.hash[3] ));
 sg13g2_dfrbp_1 _22298_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net108),
    .D(net3540),
    .Q_N(_00150_),
    .Q(\TRNG.hash[4] ));
 sg13g2_dfrbp_1 _22299_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net107),
    .D(net3629),
    .Q_N(_00153_),
    .Q(\TRNG.hash[8] ));
 sg13g2_dfrbp_1 _22300_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net106),
    .D(_01189_),
    .Q_N(_10124_),
    .Q(\TRNG.hash[10] ));
 sg13g2_dfrbp_1 _22301_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net105),
    .D(_01190_),
    .Q_N(_10123_),
    .Q(\TRNG.hash[11] ));
 sg13g2_dfrbp_1 _22302_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net104),
    .D(net3615),
    .Q_N(_00158_),
    .Q(\TRNG.hash[14] ));
 sg13g2_dfrbp_1 _22303_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net103),
    .D(_01192_),
    .Q_N(_10122_),
    .Q(\TRNG.hash[15] ));
 sg13g2_dfrbp_1 _22304_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net102),
    .D(_01193_),
    .Q_N(_00159_),
    .Q(\TRNG.hash[21] ));
 sg13g2_dfrbp_1 _22305_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net101),
    .D(_01194_),
    .Q_N(_10121_),
    .Q(\TRNG.hash[22] ));
 sg13g2_dfrbp_1 _22306_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net100),
    .D(_01195_),
    .Q_N(_10120_),
    .Q(\TRNG.hash[23] ));
 sg13g2_dfrbp_1 _22307_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net99),
    .D(_01196_),
    .Q_N(_10119_),
    .Q(\TRNG.hash[24] ));
 sg13g2_dfrbp_1 _22308_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net98),
    .D(_01197_),
    .Q_N(_10118_),
    .Q(\TRNG.hash[25] ));
 sg13g2_dfrbp_1 _22309_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net97),
    .D(_01198_),
    .Q_N(_10117_),
    .Q(\TRNG.hash[27] ));
 sg13g2_dfrbp_1 _22310_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net96),
    .D(_01199_),
    .Q_N(_10116_),
    .Q(\TRNG.hash[28] ));
 sg13g2_dfrbp_1 _22311_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net95),
    .D(_01200_),
    .Q_N(_10115_),
    .Q(\TRNG.hash[30] ));
 sg13g2_dfrbp_1 _22312_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net94),
    .D(net2838),
    .Q_N(_10114_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][0] ));
 sg13g2_dfrbp_1 _22313_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net93),
    .D(net2775),
    .Q_N(_10113_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][1] ));
 sg13g2_dfrbp_1 _22314_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net92),
    .D(_01203_),
    .Q_N(_10112_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][2] ));
 sg13g2_dfrbp_1 _22315_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net91),
    .D(net2618),
    .Q_N(_10111_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][3] ));
 sg13g2_dfrbp_1 _22316_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net90),
    .D(_01205_),
    .Q_N(_10110_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][4] ));
 sg13g2_dfrbp_1 _22317_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net89),
    .D(_01206_),
    .Q_N(_10109_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][5] ));
 sg13g2_dfrbp_1 _22318_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net88),
    .D(_01207_),
    .Q_N(_10108_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][6] ));
 sg13g2_dfrbp_1 _22319_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net87),
    .D(_01208_),
    .Q_N(_10107_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][7] ));
 sg13g2_dfrbp_1 _22320_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net86),
    .D(_01209_),
    .Q_N(_10106_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][8] ));
 sg13g2_dfrbp_1 _22321_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net85),
    .D(_01210_),
    .Q_N(_10105_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][9] ));
 sg13g2_dfrbp_1 _22322_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net84),
    .D(_01211_),
    .Q_N(_10104_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][10] ));
 sg13g2_dfrbp_1 _22323_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net83),
    .D(_01212_),
    .Q_N(_10103_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][11] ));
 sg13g2_dfrbp_1 _22324_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net82),
    .D(_01213_),
    .Q_N(_10102_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][12] ));
 sg13g2_dfrbp_1 _22325_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net81),
    .D(_01214_),
    .Q_N(_10101_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][13] ));
 sg13g2_dfrbp_1 _22326_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net80),
    .D(_01215_),
    .Q_N(_10100_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][14] ));
 sg13g2_dfrbp_1 _22327_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net79),
    .D(_01216_),
    .Q_N(_10099_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][15] ));
 sg13g2_dfrbp_1 _22328_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net78),
    .D(_01217_),
    .Q_N(_10098_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][16] ));
 sg13g2_dfrbp_1 _22329_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net77),
    .D(_01218_),
    .Q_N(_10097_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][17] ));
 sg13g2_dfrbp_1 _22330_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net76),
    .D(_01219_),
    .Q_N(_10096_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][18] ));
 sg13g2_dfrbp_1 _22331_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net75),
    .D(_01220_),
    .Q_N(_10095_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][19] ));
 sg13g2_dfrbp_1 _22332_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net74),
    .D(_01221_),
    .Q_N(_10094_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][20] ));
 sg13g2_dfrbp_1 _22333_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net73),
    .D(_01222_),
    .Q_N(_10093_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][21] ));
 sg13g2_dfrbp_1 _22334_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net72),
    .D(_01223_),
    .Q_N(_10092_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][22] ));
 sg13g2_dfrbp_1 _22335_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net71),
    .D(_01224_),
    .Q_N(_10091_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][23] ));
 sg13g2_dfrbp_1 _22336_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net70),
    .D(_01225_),
    .Q_N(_10090_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][24] ));
 sg13g2_dfrbp_1 _22337_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net69),
    .D(net2717),
    .Q_N(_10089_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][25] ));
 sg13g2_dfrbp_1 _22338_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net68),
    .D(_01227_),
    .Q_N(_10088_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][26] ));
 sg13g2_dfrbp_1 _22339_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net67),
    .D(net3256),
    .Q_N(_10087_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][27] ));
 sg13g2_dfrbp_1 _22340_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net66),
    .D(_01229_),
    .Q_N(_10086_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][28] ));
 sg13g2_dfrbp_1 _22341_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net65),
    .D(_01230_),
    .Q_N(_10085_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][29] ));
 sg13g2_dfrbp_1 _22342_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net64),
    .D(_01231_),
    .Q_N(_10084_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][30] ));
 sg13g2_dfrbp_1 _22343_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net63),
    .D(_01232_),
    .Q_N(_10083_),
    .Q(\TRNG.sha256.expand.msg_schdl.RAM[13][31] ));
 sg13g2_dfrbp_1 _22344_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net5900),
    .D(net3151),
    .Q_N(_10082_),
    .Q(\TRNG.Repetition_Count_Test.failure ));
 sg13g2_dfrbp_1 _22345_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net5900),
    .D(_01234_),
    .Q_N(_00114_),
    .Q(\TRNG.uart_start ));
 sg13g2_dfrbp_1 _22346_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net5901),
    .D(net1258),
    .Q_N(_11059_),
    .Q(\TRNG.Repetition_Count_Test.count[0] ));
 sg13g2_dfrbp_1 _22347_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net5901),
    .D(net2313),
    .Q_N(_11060_),
    .Q(\TRNG.Repetition_Count_Test.count[1] ));
 sg13g2_dfrbp_1 _22348_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net5901),
    .D(net2369),
    .Q_N(_11061_),
    .Q(\TRNG.Repetition_Count_Test.count[2] ));
 sg13g2_dfrbp_1 _22349_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net5900),
    .D(net1407),
    .Q_N(_11062_),
    .Q(\TRNG.Repetition_Count_Test.count[3] ));
 sg13g2_dfrbp_1 _22350_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net5900),
    .D(_00100_),
    .Q_N(_11063_),
    .Q(\TRNG.Repetition_Count_Test.count[4] ));
 sg13g2_dfrbp_1 _22351_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net5900),
    .D(_00101_),
    .Q_N(_11064_),
    .Q(\TRNG.Repetition_Count_Test.count[5] ));
 sg13g2_dfrbp_1 _22352_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net62),
    .D(\TRNG.NOISE_SOURCE.Noise_Source_Out ),
    .Q_N(_10081_),
    .Q(\TRNG.NOISE_SAMPLER.Sample_Out ));
 sg13g2_dfrbp_1 _22353_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net5904),
    .D(_01235_),
    .Q_N(_10080_),
    .Q(\TRNG.Word_Valid ));
 sg13g2_dfrbp_1 _22354_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net61),
    .D(_01236_),
    .Q_N(_10079_),
    .Q(\TRNG.chunk_reg[0] ));
 sg13g2_dfrbp_1 _22355_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net60),
    .D(_01237_),
    .Q_N(_10078_),
    .Q(\TRNG.chunk_reg[1] ));
 sg13g2_dfrbp_1 _22356_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net59),
    .D(_01238_),
    .Q_N(_10077_),
    .Q(\TRNG.chunk_reg[2] ));
 sg13g2_dfrbp_1 _22357_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net58),
    .D(_01239_),
    .Q_N(_10076_),
    .Q(\TRNG.chunk_reg[3] ));
 sg13g2_dfrbp_1 _22358_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net57),
    .D(_01240_),
    .Q_N(_10075_),
    .Q(\TRNG.chunk_reg[4] ));
 sg13g2_dfrbp_1 _22359_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net56),
    .D(_01241_),
    .Q_N(_10074_),
    .Q(\TRNG.chunk_reg[5] ));
 sg13g2_dfrbp_1 _22360_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net55),
    .D(_01242_),
    .Q_N(_10073_),
    .Q(\TRNG.chunk_reg[6] ));
 sg13g2_dfrbp_1 _22361_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net763),
    .D(_01243_),
    .Q_N(_11065_),
    .Q(\TRNG.chunk_reg[7] ));
 sg13g2_dfrbp_1 _22362_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net5902),
    .D(_02157_),
    .Q_N(_11066_),
    .Q(\TRNG.state[0] ));
 sg13g2_dfrbp_1 _22363_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net5904),
    .D(net3380),
    .Q_N(_11067_),
    .Q(\TRNG.state[1] ));
 sg13g2_dfrbp_1 _22364_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net5903),
    .D(net1147),
    .Q_N(_00119_),
    .Q(\TRNG.state[2] ));
 sg13g2_dfrbp_1 _22365_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net5919),
    .D(_01244_),
    .Q_N(_10072_),
    .Q(\TRNG.Word_Out[0] ));
 sg13g2_dfrbp_1 _22366_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net5920),
    .D(net1865),
    .Q_N(_10071_),
    .Q(\TRNG.Word_Out[1] ));
 sg13g2_dfrbp_1 _22367_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net5926),
    .D(_01246_),
    .Q_N(_10070_),
    .Q(\TRNG.Word_Out[2] ));
 sg13g2_dfrbp_1 _22368_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net5927),
    .D(net2612),
    .Q_N(_10069_),
    .Q(\TRNG.Word_Out[3] ));
 sg13g2_dfrbp_1 _22369_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net5983),
    .D(_01248_),
    .Q_N(_10068_),
    .Q(\TRNG.Word_Out[4] ));
 sg13g2_dfrbp_1 _22370_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net5984),
    .D(net1938),
    .Q_N(_10067_),
    .Q(\TRNG.Word_Out[5] ));
 sg13g2_dfrbp_1 _22371_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net5998),
    .D(_01250_),
    .Q_N(_10066_),
    .Q(\TRNG.Word_Out[6] ));
 sg13g2_dfrbp_1 _22372_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net6002),
    .D(_01251_),
    .Q_N(_10065_),
    .Q(\TRNG.Word_Out[7] ));
 sg13g2_dfrbp_1 _22373_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net6002),
    .D(net1194),
    .Q_N(_10064_),
    .Q(\TRNG.Word_Out[8] ));
 sg13g2_dfrbp_1 _22374_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net5995),
    .D(_01253_),
    .Q_N(_10063_),
    .Q(\TRNG.Word_Out[9] ));
 sg13g2_dfrbp_1 _22375_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net5995),
    .D(net1719),
    .Q_N(_10062_),
    .Q(\TRNG.Word_Out[10] ));
 sg13g2_dfrbp_1 _22376_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net5994),
    .D(net2616),
    .Q_N(_10061_),
    .Q(\TRNG.Word_Out[11] ));
 sg13g2_dfrbp_1 _22377_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net5965),
    .D(net2691),
    .Q_N(_10060_),
    .Q(\TRNG.Word_Out[12] ));
 sg13g2_dfrbp_1 _22378_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net5963),
    .D(_01257_),
    .Q_N(_10059_),
    .Q(\TRNG.Word_Out[13] ));
 sg13g2_dfrbp_1 _22379_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net5964),
    .D(net1230),
    .Q_N(_10058_),
    .Q(\TRNG.Word_Out[14] ));
 sg13g2_dfrbp_1 _22380_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net6018),
    .D(_01259_),
    .Q_N(_10057_),
    .Q(\TRNG.Word_Out[15] ));
 sg13g2_dfrbp_1 _22381_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net6021),
    .D(net1363),
    .Q_N(_10056_),
    .Q(\TRNG.Word_Out[16] ));
 sg13g2_dfrbp_1 _22382_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net6013),
    .D(_01261_),
    .Q_N(_10055_),
    .Q(\TRNG.Word_Out[17] ));
 sg13g2_dfrbp_1 _22383_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net6016),
    .D(net1979),
    .Q_N(_10054_),
    .Q(\TRNG.Word_Out[18] ));
 sg13g2_dfrbp_1 _22384_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net6009),
    .D(net2470),
    .Q_N(_10053_),
    .Q(\TRNG.Word_Out[19] ));
 sg13g2_dfrbp_1 _22385_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net5954),
    .D(_01264_),
    .Q_N(_10052_),
    .Q(\TRNG.Word_Out[20] ));
 sg13g2_dfrbp_1 _22386_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net5950),
    .D(_01265_),
    .Q_N(_10051_),
    .Q(\TRNG.Word_Out[21] ));
 sg13g2_dfrbp_1 _22387_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net5950),
    .D(_01266_),
    .Q_N(_10050_),
    .Q(\TRNG.Word_Out[22] ));
 sg13g2_dfrbp_1 _22388_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net5935),
    .D(net2130),
    .Q_N(_10049_),
    .Q(\TRNG.Word_Out[23] ));
 sg13g2_dfrbp_1 _22389_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net5937),
    .D(_01268_),
    .Q_N(_10048_),
    .Q(\TRNG.Word_Out[24] ));
 sg13g2_dfrbp_1 _22390_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net5933),
    .D(net1151),
    .Q_N(_10047_),
    .Q(\TRNG.Word_Out[25] ));
 sg13g2_dfrbp_1 _22391_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net5911),
    .D(_01270_),
    .Q_N(_10046_),
    .Q(\TRNG.Word_Out[26] ));
 sg13g2_dfrbp_1 _22392_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net5911),
    .D(net2281),
    .Q_N(_10045_),
    .Q(\TRNG.Word_Out[27] ));
 sg13g2_dfrbp_1 _22393_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net5915),
    .D(net2820),
    .Q_N(_10044_),
    .Q(\TRNG.Word_Out[28] ));
 sg13g2_dfrbp_1 _22394_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net5915),
    .D(_01273_),
    .Q_N(_10043_),
    .Q(\TRNG.Word_Out[29] ));
 sg13g2_dfrbp_1 _22395_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net5919),
    .D(_01274_),
    .Q_N(_10042_),
    .Q(\TRNG.Word_Out[30] ));
 sg13g2_dfrbp_1 _22396_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net5919),
    .D(net1192),
    .Q_N(_10041_),
    .Q(\TRNG.Word_Out[31] ));
 sg13g2_dfrbp_1 _22397_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net5920),
    .D(net2487),
    .Q_N(_10040_),
    .Q(\TRNG.Word_Out[32] ));
 sg13g2_dfrbp_1 _22398_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net5926),
    .D(net2574),
    .Q_N(_10039_),
    .Q(\TRNG.Word_Out[33] ));
 sg13g2_dfrbp_1 _22399_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net5926),
    .D(net2710),
    .Q_N(_10038_),
    .Q(\TRNG.Word_Out[34] ));
 sg13g2_dfrbp_1 _22400_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net5928),
    .D(_01279_),
    .Q_N(_10037_),
    .Q(\TRNG.Word_Out[35] ));
 sg13g2_dfrbp_1 _22401_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net5981),
    .D(_01280_),
    .Q_N(_10036_),
    .Q(\TRNG.Word_Out[36] ));
 sg13g2_dfrbp_1 _22402_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net5986),
    .D(net1224),
    .Q_N(_10035_),
    .Q(\TRNG.Word_Out[37] ));
 sg13g2_dfrbp_1 _22403_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net6004),
    .D(_01282_),
    .Q_N(_10034_),
    .Q(\TRNG.Word_Out[38] ));
 sg13g2_dfrbp_1 _22404_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net6005),
    .D(net1240),
    .Q_N(_10033_),
    .Q(\TRNG.Word_Out[39] ));
 sg13g2_dfrbp_1 _22405_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net6057),
    .D(_01284_),
    .Q_N(_10032_),
    .Q(\TRNG.Word_Out[40] ));
 sg13g2_dfrbp_1 _22406_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net6058),
    .D(net1654),
    .Q_N(_10031_),
    .Q(\TRNG.Word_Out[41] ));
 sg13g2_dfrbp_1 _22407_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net6056),
    .D(_01286_),
    .Q_N(_10030_),
    .Q(\TRNG.Word_Out[42] ));
 sg13g2_dfrbp_1 _22408_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net6048),
    .D(_01287_),
    .Q_N(_10029_),
    .Q(\TRNG.Word_Out[43] ));
 sg13g2_dfrbp_1 _22409_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net6045),
    .D(_01288_),
    .Q_N(_10028_),
    .Q(\TRNG.Word_Out[44] ));
 sg13g2_dfrbp_1 _22410_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net6045),
    .D(_01289_),
    .Q_N(_10027_),
    .Q(\TRNG.Word_Out[45] ));
 sg13g2_dfrbp_1 _22411_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net6023),
    .D(_01290_),
    .Q_N(_10026_),
    .Q(\TRNG.Word_Out[46] ));
 sg13g2_dfrbp_1 _22412_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net6024),
    .D(net1822),
    .Q_N(_10025_),
    .Q(\TRNG.Word_Out[47] ));
 sg13g2_dfrbp_1 _22413_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net6035),
    .D(net2463),
    .Q_N(_10024_),
    .Q(\TRNG.Word_Out[48] ));
 sg13g2_dfrbp_1 _22414_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net6028),
    .D(_01293_),
    .Q_N(_10023_),
    .Q(\TRNG.Word_Out[49] ));
 sg13g2_dfrbp_1 _22415_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net6014),
    .D(_01294_),
    .Q_N(_10022_),
    .Q(\TRNG.Word_Out[50] ));
 sg13g2_dfrbp_1 _22416_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net6010),
    .D(net2109),
    .Q_N(_10021_),
    .Q(\TRNG.Word_Out[51] ));
 sg13g2_dfrbp_1 _22417_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net5956),
    .D(_01296_),
    .Q_N(_10020_),
    .Q(\TRNG.Word_Out[52] ));
 sg13g2_dfrbp_1 _22418_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net5955),
    .D(_01297_),
    .Q_N(_10019_),
    .Q(\TRNG.Word_Out[53] ));
 sg13g2_dfrbp_1 _22419_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net5952),
    .D(net1942),
    .Q_N(_10018_),
    .Q(\TRNG.Word_Out[54] ));
 sg13g2_dfrbp_1 _22420_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net5938),
    .D(_01299_),
    .Q_N(_10017_),
    .Q(\TRNG.Word_Out[55] ));
 sg13g2_dfrbp_1 _22421_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net5932),
    .D(net1723),
    .Q_N(_10016_),
    .Q(\TRNG.Word_Out[56] ));
 sg13g2_dfrbp_1 _22422_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net5933),
    .D(net2236),
    .Q_N(_10015_),
    .Q(\TRNG.Word_Out[57] ));
 sg13g2_dfrbp_1 _22423_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net5913),
    .D(_01302_),
    .Q_N(_10014_),
    .Q(\TRNG.Word_Out[58] ));
 sg13g2_dfrbp_1 _22424_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net5915),
    .D(net2579),
    .Q_N(_10013_),
    .Q(\TRNG.Word_Out[59] ));
 sg13g2_dfrbp_1 _22425_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net5916),
    .D(_01304_),
    .Q_N(_10012_),
    .Q(\TRNG.Word_Out[60] ));
 sg13g2_dfrbp_1 _22426_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net5969),
    .D(net1216),
    .Q_N(_10011_),
    .Q(\TRNG.Word_Out[61] ));
 sg13g2_dfrbp_1 _22427_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net5922),
    .D(_01306_),
    .Q_N(_10010_),
    .Q(\TRNG.Word_Out[62] ));
 sg13g2_dfrbp_1 _22428_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net5922),
    .D(_01307_),
    .Q_N(_10009_),
    .Q(\TRNG.Word_Out[63] ));
 sg13g2_dfrbp_1 _22429_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net5924),
    .D(net1171),
    .Q_N(_10008_),
    .Q(\TRNG.Word_Out[64] ));
 sg13g2_dfrbp_1 _22430_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net5930),
    .D(net2891),
    .Q_N(_10007_),
    .Q(\TRNG.Word_Out[65] ));
 sg13g2_dfrbp_1 _22431_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net5929),
    .D(_01310_),
    .Q_N(_10006_),
    .Q(\TRNG.Word_Out[66] ));
 sg13g2_dfrbp_1 _22432_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net5929),
    .D(net1858),
    .Q_N(_10005_),
    .Q(\TRNG.Word_Out[67] ));
 sg13g2_dfrbp_1 _22433_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net5928),
    .D(net2124),
    .Q_N(_10004_),
    .Q(\TRNG.Word_Out[68] ));
 sg13g2_dfrbp_1 _22434_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net6001),
    .D(_01313_),
    .Q_N(_10003_),
    .Q(\TRNG.Word_Out[69] ));
 sg13g2_dfrbp_1 _22435_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net6005),
    .D(_01314_),
    .Q_N(_10002_),
    .Q(\TRNG.Word_Out[70] ));
 sg13g2_dfrbp_1 _22436_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net6052),
    .D(net1207),
    .Q_N(_10001_),
    .Q(\TRNG.Word_Out[71] ));
 sg13g2_dfrbp_1 _22437_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net6053),
    .D(net1578),
    .Q_N(_10000_),
    .Q(\TRNG.Word_Out[72] ));
 sg13g2_dfrbp_1 _22438_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net6057),
    .D(net1725),
    .Q_N(_09999_),
    .Q(\TRNG.Word_Out[73] ));
 sg13g2_dfrbp_1 _22439_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net6047),
    .D(_01318_),
    .Q_N(_09998_),
    .Q(\TRNG.Word_Out[74] ));
 sg13g2_dfrbp_1 _22440_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net6047),
    .D(net2154),
    .Q_N(_09997_),
    .Q(\TRNG.Word_Out[75] ));
 sg13g2_dfrbp_1 _22441_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net6045),
    .D(_01320_),
    .Q_N(_09996_),
    .Q(\TRNG.Word_Out[76] ));
 sg13g2_dfrbp_1 _22442_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net6019),
    .D(_01321_),
    .Q_N(_09995_),
    .Q(\TRNG.Word_Out[77] ));
 sg13g2_dfrbp_1 _22443_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net6018),
    .D(_01322_),
    .Q_N(_09994_),
    .Q(\TRNG.Word_Out[78] ));
 sg13g2_dfrbp_1 _22444_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net6021),
    .D(net1201),
    .Q_N(_09993_),
    .Q(\TRNG.Word_Out[79] ));
 sg13g2_dfrbp_1 _22445_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net6022),
    .D(net1944),
    .Q_N(_09992_),
    .Q(\TRNG.Word_Out[80] ));
 sg13g2_dfrbp_1 _22446_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net6035),
    .D(net2100),
    .Q_N(_09991_),
    .Q(\TRNG.Word_Out[81] ));
 sg13g2_dfrbp_1 _22447_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net6014),
    .D(net2374),
    .Q_N(_09990_),
    .Q(\TRNG.Word_Out[82] ));
 sg13g2_dfrbp_1 _22448_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net6010),
    .D(net2434),
    .Q_N(_09989_),
    .Q(\TRNG.Word_Out[83] ));
 sg13g2_dfrbp_1 _22449_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net5964),
    .D(_01328_),
    .Q_N(_09988_),
    .Q(\TRNG.Word_Out[84] ));
 sg13g2_dfrbp_1 _22450_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net5963),
    .D(net2285),
    .Q_N(_09987_),
    .Q(\TRNG.Word_Out[85] ));
 sg13g2_dfrbp_1 _22451_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net5952),
    .D(_01330_),
    .Q_N(_09986_),
    .Q(\TRNG.Word_Out[86] ));
 sg13g2_dfrbp_1 _22452_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net5951),
    .D(_01331_),
    .Q_N(_09985_),
    .Q(\TRNG.Word_Out[87] ));
 sg13g2_dfrbp_1 _22453_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net5937),
    .D(_01332_),
    .Q_N(_09984_),
    .Q(\TRNG.Word_Out[88] ));
 sg13g2_dfrbp_1 _22454_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net5941),
    .D(net1242),
    .Q_N(_09983_),
    .Q(\TRNG.Word_Out[89] ));
 sg13g2_dfrbp_1 _22455_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net5911),
    .D(_01334_),
    .Q_N(_09982_),
    .Q(\TRNG.Word_Out[90] ));
 sg13g2_dfrbp_1 _22456_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net5911),
    .D(net2203),
    .Q_N(_09981_),
    .Q(\TRNG.Word_Out[91] ));
 sg13g2_dfrbp_1 _22457_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net5912),
    .D(net2702),
    .Q_N(_09980_),
    .Q(\TRNG.Word_Out[92] ));
 sg13g2_dfrbp_1 _22458_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net5915),
    .D(_01337_),
    .Q_N(_09979_),
    .Q(\TRNG.Word_Out[93] ));
 sg13g2_dfrbp_1 _22459_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net5922),
    .D(net1177),
    .Q_N(_09978_),
    .Q(\TRNG.Word_Out[94] ));
 sg13g2_dfrbp_1 _22460_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net5922),
    .D(net1764),
    .Q_N(_09977_),
    .Q(\TRNG.Word_Out[95] ));
 sg13g2_dfrbp_1 _22461_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net5969),
    .D(net2059),
    .Q_N(_09976_),
    .Q(\TRNG.Word_Out[96] ));
 sg13g2_dfrbp_1 _22462_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net5971),
    .D(_01341_),
    .Q_N(_09975_),
    .Q(\TRNG.Word_Out[97] ));
 sg13g2_dfrbp_1 _22463_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net5971),
    .D(_01342_),
    .Q_N(_09974_),
    .Q(\TRNG.Word_Out[98] ));
 sg13g2_dfrbp_1 _22464_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net5979),
    .D(net1817),
    .Q_N(_09973_),
    .Q(\TRNG.Word_Out[99] ));
 sg13g2_dfrbp_1 _22465_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net5983),
    .D(_01344_),
    .Q_N(_09972_),
    .Q(\TRNG.Word_Out[100] ));
 sg13g2_dfrbp_1 _22466_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net5999),
    .D(net1880),
    .Q_N(_09971_),
    .Q(\TRNG.Word_Out[101] ));
 sg13g2_dfrbp_1 _22467_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net5998),
    .D(_01346_),
    .Q_N(_09970_),
    .Q(\TRNG.Word_Out[102] ));
 sg13g2_dfrbp_1 _22468_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net6003),
    .D(_01347_),
    .Q_N(_09969_),
    .Q(\TRNG.Word_Out[103] ));
 sg13g2_dfrbp_1 _22469_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net6050),
    .D(net1183),
    .Q_N(_09968_),
    .Q(\TRNG.Word_Out[104] ));
 sg13g2_dfrbp_1 _22470_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net6051),
    .D(net1644),
    .Q_N(_09967_),
    .Q(\TRNG.Word_Out[105] ));
 sg13g2_dfrbp_1 _22471_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net6043),
    .D(net2033),
    .Q_N(_09966_),
    .Q(\TRNG.Word_Out[106] ));
 sg13g2_dfrbp_1 _22472_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net6042),
    .D(_01351_),
    .Q_N(_09965_),
    .Q(\TRNG.Word_Out[107] ));
 sg13g2_dfrbp_1 _22473_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net5993),
    .D(net1833),
    .Q_N(_09964_),
    .Q(\TRNG.Word_Out[108] ));
 sg13g2_dfrbp_1 _22474_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net5965),
    .D(net2531),
    .Q_N(_09963_),
    .Q(\TRNG.Word_Out[109] ));
 sg13g2_dfrbp_1 _22475_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net5964),
    .D(_01354_),
    .Q_N(_09962_),
    .Q(\TRNG.Word_Out[110] ));
 sg13g2_dfrbp_1 _22476_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net6018),
    .D(_01355_),
    .Q_N(_09961_),
    .Q(\TRNG.Word_Out[111] ));
 sg13g2_dfrbp_1 _22477_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net6021),
    .D(_01356_),
    .Q_N(_09960_),
    .Q(\TRNG.Word_Out[112] ));
 sg13g2_dfrbp_1 _22478_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net6014),
    .D(net1226),
    .Q_N(_09959_),
    .Q(\TRNG.Word_Out[113] ));
 sg13g2_dfrbp_1 _22479_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net6014),
    .D(net1462),
    .Q_N(_09958_),
    .Q(\TRNG.Word_Out[114] ));
 sg13g2_dfrbp_1 _22480_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net6011),
    .D(_01359_),
    .Q_N(_09957_),
    .Q(\TRNG.Word_Out[115] ));
 sg13g2_dfrbp_1 _22481_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net6011),
    .D(_01360_),
    .Q_N(_09956_),
    .Q(\TRNG.Word_Out[116] ));
 sg13g2_dfrbp_1 _22482_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net5955),
    .D(net2241),
    .Q_N(_09955_),
    .Q(\TRNG.Word_Out[117] ));
 sg13g2_dfrbp_1 _22483_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net5951),
    .D(_01362_),
    .Q_N(_09954_),
    .Q(\TRNG.Word_Out[118] ));
 sg13g2_dfrbp_1 _22484_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net5936),
    .D(net2015),
    .Q_N(_09953_),
    .Q(\TRNG.Word_Out[119] ));
 sg13g2_dfrbp_1 _22485_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net5932),
    .D(_01364_),
    .Q_N(_09952_),
    .Q(\TRNG.Word_Out[120] ));
 sg13g2_dfrbp_1 _22486_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net5910),
    .D(net1550),
    .Q_N(_09951_),
    .Q(\TRNG.Word_Out[121] ));
 sg13g2_dfrbp_1 _22487_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net5910),
    .D(_01366_),
    .Q_N(_09950_),
    .Q(\TRNG.Word_Out[122] ));
 sg13g2_dfrbp_1 _22488_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net5911),
    .D(_01367_),
    .Q_N(_09949_),
    .Q(\TRNG.Word_Out[123] ));
 sg13g2_dfrbp_1 _22489_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net5912),
    .D(_01368_),
    .Q_N(_09948_),
    .Q(\TRNG.Word_Out[124] ));
 sg13g2_dfrbp_1 _22490_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net5912),
    .D(_01369_),
    .Q_N(_09947_),
    .Q(\TRNG.Word_Out[125] ));
 sg13g2_dfrbp_1 _22491_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net5919),
    .D(net1218),
    .Q_N(_09946_),
    .Q(\TRNG.Word_Out[126] ));
 sg13g2_dfrbp_1 _22492_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net5921),
    .D(_01371_),
    .Q_N(_09945_),
    .Q(\TRNG.Word_Out[127] ));
 sg13g2_dfrbp_1 _22493_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net5924),
    .D(net1153),
    .Q_N(_09944_),
    .Q(\TRNG.Word_Out[128] ));
 sg13g2_dfrbp_1 _22494_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net5924),
    .D(net1928),
    .Q_N(_09943_),
    .Q(\TRNG.Word_Out[129] ));
 sg13g2_dfrbp_1 _22495_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net5927),
    .D(_01374_),
    .Q_N(_09942_),
    .Q(\TRNG.Word_Out[130] ));
 sg13g2_dfrbp_1 _22496_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net5928),
    .D(_01375_),
    .Q_N(_09941_),
    .Q(\TRNG.Word_Out[131] ));
 sg13g2_dfrbp_1 _22497_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net5981),
    .D(net1368),
    .Q_N(_09940_),
    .Q(\TRNG.Word_Out[132] ));
 sg13g2_dfrbp_1 _22498_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net5984),
    .D(_01377_),
    .Q_N(_09939_),
    .Q(\TRNG.Word_Out[133] ));
 sg13g2_dfrbp_1 _22499_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net6001),
    .D(net1161),
    .Q_N(_09938_),
    .Q(\TRNG.Word_Out[134] ));
 sg13g2_dfrbp_1 _22500_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net6002),
    .D(_01379_),
    .Q_N(_09937_),
    .Q(\TRNG.Word_Out[135] ));
 sg13g2_dfrbp_1 _22501_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net5996),
    .D(net1222),
    .Q_N(_09936_),
    .Q(\TRNG.Word_Out[136] ));
 sg13g2_dfrbp_1 _22502_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net5996),
    .D(_01381_),
    .Q_N(_09935_),
    .Q(\TRNG.Word_Out[137] ));
 sg13g2_dfrbp_1 _22503_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net6044),
    .D(_01382_),
    .Q_N(_09934_),
    .Q(\TRNG.Word_Out[138] ));
 sg13g2_dfrbp_1 _22504_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net6043),
    .D(net1145),
    .Q_N(_09933_),
    .Q(\TRNG.Word_Out[139] ));
 sg13g2_dfrbp_1 _22505_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net6041),
    .D(net2249),
    .Q_N(_09932_),
    .Q(\TRNG.Word_Out[140] ));
 sg13g2_dfrbp_1 _22506_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net6045),
    .D(_01385_),
    .Q_N(_09931_),
    .Q(\TRNG.Word_Out[141] ));
 sg13g2_dfrbp_1 _22507_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net6023),
    .D(net1163),
    .Q_N(_09930_),
    .Q(\TRNG.Word_Out[142] ));
 sg13g2_dfrbp_1 _22508_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net6024),
    .D(net2262),
    .Q_N(_09929_),
    .Q(\TRNG.Word_Out[143] ));
 sg13g2_dfrbp_1 _22509_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net6035),
    .D(net2318),
    .Q_N(_09928_),
    .Q(\TRNG.Word_Out[144] ));
 sg13g2_dfrbp_1 _22510_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net6036),
    .D(net2504),
    .Q_N(_09927_),
    .Q(\TRNG.Word_Out[145] ));
 sg13g2_dfrbp_1 _22511_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net6029),
    .D(net2545),
    .Q_N(_09926_),
    .Q(\TRNG.Word_Out[146] ));
 sg13g2_dfrbp_1 _22512_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net6011),
    .D(_01391_),
    .Q_N(_09925_),
    .Q(\TRNG.Word_Out[147] ));
 sg13g2_dfrbp_1 _22513_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net5956),
    .D(net2397),
    .Q_N(_09924_),
    .Q(\TRNG.Word_Out[148] ));
 sg13g2_dfrbp_1 _22514_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net5963),
    .D(_01393_),
    .Q_N(_09923_),
    .Q(\TRNG.Word_Out[149] ));
 sg13g2_dfrbp_1 _22515_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net5962),
    .D(net1542),
    .Q_N(_09922_),
    .Q(\TRNG.Word_Out[150] ));
 sg13g2_dfrbp_1 _22516_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net5959),
    .D(net1867),
    .Q_N(_09921_),
    .Q(\TRNG.Word_Out[151] ));
 sg13g2_dfrbp_1 _22517_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net5944),
    .D(net1922),
    .Q_N(_09920_),
    .Q(\TRNG.Word_Out[152] ));
 sg13g2_dfrbp_1 _22518_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net5944),
    .D(net2423),
    .Q_N(_09919_),
    .Q(\TRNG.Word_Out[153] ));
 sg13g2_dfrbp_1 _22519_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net5940),
    .D(_01398_),
    .Q_N(_09918_),
    .Q(\TRNG.Word_Out[154] ));
 sg13g2_dfrbp_1 _22520_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net5913),
    .D(net1190),
    .Q_N(_09917_),
    .Q(\TRNG.Word_Out[155] ));
 sg13g2_dfrbp_1 _22521_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net5911),
    .D(_01400_),
    .Q_N(_09916_),
    .Q(\TRNG.Word_Out[156] ));
 sg13g2_dfrbp_1 _22522_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net5919),
    .D(_01401_),
    .Q_N(_09915_),
    .Q(\TRNG.Word_Out[157] ));
 sg13g2_dfrbp_1 _22523_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net5919),
    .D(net1237),
    .Q_N(_09914_),
    .Q(\TRNG.Word_Out[158] ));
 sg13g2_dfrbp_1 _22524_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net5919),
    .D(net1961),
    .Q_N(_09913_),
    .Q(\TRNG.Word_Out[159] ));
 sg13g2_dfrbp_1 _22525_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net5920),
    .D(net2409),
    .Q_N(_09912_),
    .Q(\TRNG.Word_Out[160] ));
 sg13g2_dfrbp_1 _22526_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net5926),
    .D(_01405_),
    .Q_N(_09911_),
    .Q(\TRNG.Word_Out[161] ));
 sg13g2_dfrbp_1 _22527_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net5926),
    .D(net2411),
    .Q_N(_09910_),
    .Q(\TRNG.Word_Out[162] ));
 sg13g2_dfrbp_1 _22528_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net5929),
    .D(_01407_),
    .Q_N(_09909_),
    .Q(\TRNG.Word_Out[163] ));
 sg13g2_dfrbp_1 _22529_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net5929),
    .D(_01408_),
    .Q_N(_09908_),
    .Q(\TRNG.Word_Out[164] ));
 sg13g2_dfrbp_1 _22530_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net5986),
    .D(net1580),
    .Q_N(_09907_),
    .Q(\TRNG.Word_Out[165] ));
 sg13g2_dfrbp_1 _22531_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net6004),
    .D(_01410_),
    .Q_N(_09906_),
    .Q(\TRNG.Word_Out[166] ));
 sg13g2_dfrbp_1 _22532_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net6002),
    .D(net1494),
    .Q_N(_09905_),
    .Q(\TRNG.Word_Out[167] ));
 sg13g2_dfrbp_1 _22533_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net6002),
    .D(net2903),
    .Q_N(_09904_),
    .Q(\TRNG.Word_Out[168] ));
 sg13g2_dfrbp_1 _22534_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net5996),
    .D(_01413_),
    .Q_N(_09903_),
    .Q(\TRNG.Word_Out[169] ));
 sg13g2_dfrbp_1 _22535_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net5996),
    .D(net1570),
    .Q_N(_09902_),
    .Q(\TRNG.Word_Out[170] ));
 sg13g2_dfrbp_1 _22536_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net5994),
    .D(net2406),
    .Q_N(_09901_),
    .Q(\TRNG.Word_Out[171] ));
 sg13g2_dfrbp_1 _22537_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net5994),
    .D(_01416_),
    .Q_N(_09900_),
    .Q(\TRNG.Word_Out[172] ));
 sg13g2_dfrbp_1 _22538_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net5966),
    .D(net2234),
    .Q_N(_09899_),
    .Q(\TRNG.Word_Out[173] ));
 sg13g2_dfrbp_1 _22539_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net6019),
    .D(_01418_),
    .Q_N(_09898_),
    .Q(\TRNG.Word_Out[174] ));
 sg13g2_dfrbp_1 _22540_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net6024),
    .D(net1157),
    .Q_N(_09897_),
    .Q(\TRNG.Word_Out[175] ));
 sg13g2_dfrbp_1 _22541_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net6035),
    .D(net2712),
    .Q_N(_09896_),
    .Q(\TRNG.Word_Out[176] ));
 sg13g2_dfrbp_1 _22542_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net6027),
    .D(_01421_),
    .Q_N(_09895_),
    .Q(\TRNG.Word_Out[177] ));
 sg13g2_dfrbp_1 _22543_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net6027),
    .D(net2104),
    .Q_N(_09894_),
    .Q(\TRNG.Word_Out[178] ));
 sg13g2_dfrbp_1 _22544_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net6009),
    .D(_01423_),
    .Q_N(_09893_),
    .Q(\TRNG.Word_Out[179] ));
 sg13g2_dfrbp_1 _22545_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net6008),
    .D(net2466),
    .Q_N(_09892_),
    .Q(\TRNG.Word_Out[180] ));
 sg13g2_dfrbp_1 _22546_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net5953),
    .D(_01425_),
    .Q_N(_09891_),
    .Q(\TRNG.Word_Out[181] ));
 sg13g2_dfrbp_1 _22547_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net5950),
    .D(net2055),
    .Q_N(_09890_),
    .Q(\TRNG.Word_Out[182] ));
 sg13g2_dfrbp_1 _22548_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net5938),
    .D(_01427_),
    .Q_N(_09889_),
    .Q(\TRNG.Word_Out[183] ));
 sg13g2_dfrbp_1 _22549_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net5938),
    .D(net2220),
    .Q_N(_09888_),
    .Q(\TRNG.Word_Out[184] ));
 sg13g2_dfrbp_1 _22550_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net5945),
    .D(_01429_),
    .Q_N(_09887_),
    .Q(\TRNG.Word_Out[185] ));
 sg13g2_dfrbp_1 _22551_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net5945),
    .D(net1955),
    .Q_N(_09886_),
    .Q(\TRNG.Word_Out[186] ));
 sg13g2_dfrbp_1 _22552_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net5941),
    .D(net2179),
    .Q_N(_09885_),
    .Q(\TRNG.Word_Out[187] ));
 sg13g2_dfrbp_1 _22553_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net5943),
    .D(net2428),
    .Q_N(_09884_),
    .Q(\TRNG.Word_Out[188] ));
 sg13g2_dfrbp_1 _22554_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net5946),
    .D(_01433_),
    .Q_N(_09883_),
    .Q(\TRNG.Word_Out[189] ));
 sg13g2_dfrbp_1 _22555_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net5970),
    .D(net1203),
    .Q_N(_09882_),
    .Q(\TRNG.Word_Out[190] ));
 sg13g2_dfrbp_1 _22556_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net5974),
    .D(net2084),
    .Q_N(_09881_),
    .Q(\TRNG.Word_Out[191] ));
 sg13g2_dfrbp_1 _22557_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net5972),
    .D(_01436_),
    .Q_N(_09880_),
    .Q(\TRNG.Word_Out[192] ));
 sg13g2_dfrbp_1 _22558_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net5971),
    .D(net1134),
    .Q_N(_09879_),
    .Q(\TRNG.Word_Out[193] ));
 sg13g2_dfrbp_1 _22559_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net5980),
    .D(net2876),
    .Q_N(_09878_),
    .Q(\TRNG.Word_Out[194] ));
 sg13g2_dfrbp_1 _22560_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net5981),
    .D(_01439_),
    .Q_N(_09877_),
    .Q(\TRNG.Word_Out[195] ));
 sg13g2_dfrbp_1 _22561_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net5982),
    .D(net1963),
    .Q_N(_09876_),
    .Q(\TRNG.Word_Out[196] ));
 sg13g2_dfrbp_1 _22562_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net6000),
    .D(_01441_),
    .Q_N(_09875_),
    .Q(\TRNG.Word_Out[197] ));
 sg13g2_dfrbp_1 _22563_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net6004),
    .D(net1574),
    .Q_N(_09874_),
    .Q(\TRNG.Word_Out[198] ));
 sg13g2_dfrbp_1 _22564_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net6050),
    .D(net1750),
    .Q_N(_09873_),
    .Q(\TRNG.Word_Out[199] ));
 sg13g2_dfrbp_1 _22565_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net6050),
    .D(_01444_),
    .Q_N(_09872_),
    .Q(\TRNG.Word_Out[200] ));
 sg13g2_dfrbp_1 _22566_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net6051),
    .D(net1281),
    .Q_N(_09871_),
    .Q(\TRNG.Word_Out[201] ));
 sg13g2_dfrbp_1 _22567_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net6044),
    .D(net2985),
    .Q_N(_09870_),
    .Q(\TRNG.Word_Out[202] ));
 sg13g2_dfrbp_1 _22568_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net5990),
    .D(_01447_),
    .Q_N(_09869_),
    .Q(\TRNG.Word_Out[203] ));
 sg13g2_dfrbp_1 _22569_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net5961),
    .D(_01448_),
    .Q_N(_09868_),
    .Q(\TRNG.Word_Out[204] ));
 sg13g2_dfrbp_1 _22570_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net5961),
    .D(_01449_),
    .Q_N(_09867_),
    .Q(\TRNG.Word_Out[205] ));
 sg13g2_dfrbp_1 _22571_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net5964),
    .D(_01450_),
    .Q_N(_09866_),
    .Q(\TRNG.Word_Out[206] ));
 sg13g2_dfrbp_1 _22572_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net6020),
    .D(net2006),
    .Q_N(_09865_),
    .Q(\TRNG.Word_Out[207] ));
 sg13g2_dfrbp_1 _22573_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net6014),
    .D(_01452_),
    .Q_N(_09864_),
    .Q(\TRNG.Word_Out[208] ));
 sg13g2_dfrbp_1 _22574_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net6028),
    .D(net1892),
    .Q_N(_09863_),
    .Q(\TRNG.Word_Out[209] ));
 sg13g2_dfrbp_1 _22575_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net6014),
    .D(net1974),
    .Q_N(_09862_),
    .Q(\TRNG.Word_Out[210] ));
 sg13g2_dfrbp_1 _22576_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net6010),
    .D(net2115),
    .Q_N(_09861_),
    .Q(\TRNG.Word_Out[211] ));
 sg13g2_dfrbp_1 _22577_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net5956),
    .D(_01456_),
    .Q_N(_09860_),
    .Q(\TRNG.Word_Out[212] ));
 sg13g2_dfrbp_1 _22578_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net5963),
    .D(_01457_),
    .Q_N(_09859_),
    .Q(\TRNG.Word_Out[213] ));
 sg13g2_dfrbp_1 _22579_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net5959),
    .D(net2447),
    .Q_N(_09858_),
    .Q(\TRNG.Word_Out[214] ));
 sg13g2_dfrbp_1 _22580_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net5959),
    .D(_01459_),
    .Q_N(_09857_),
    .Q(\TRNG.Word_Out[215] ));
 sg13g2_dfrbp_1 _22581_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net5944),
    .D(net1905),
    .Q_N(_09856_),
    .Q(\TRNG.Word_Out[216] ));
 sg13g2_dfrbp_1 _22582_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net5944),
    .D(_01461_),
    .Q_N(_09855_),
    .Q(\TRNG.Word_Out[217] ));
 sg13g2_dfrbp_1 _22583_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net5941),
    .D(_01462_),
    .Q_N(_09854_),
    .Q(\TRNG.Word_Out[218] ));
 sg13g2_dfrbp_1 _22584_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net5943),
    .D(net1995),
    .Q_N(_09853_),
    .Q(\TRNG.Word_Out[219] ));
 sg13g2_dfrbp_1 _22585_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net5946),
    .D(_01464_),
    .Q_N(_09852_),
    .Q(\TRNG.Word_Out[220] ));
 sg13g2_dfrbp_1 _22586_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net5947),
    .D(net2367),
    .Q_N(_09851_),
    .Q(\TRNG.Word_Out[221] ));
 sg13g2_dfrbp_1 _22587_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net5989),
    .D(_01466_),
    .Q_N(_09850_),
    .Q(\TRNG.Word_Out[222] ));
 sg13g2_dfrbp_1 _22588_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net5989),
    .D(net1948),
    .Q_N(_09849_),
    .Q(\TRNG.Word_Out[223] ));
 sg13g2_dfrbp_1 _22589_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net5991),
    .D(_01468_),
    .Q_N(_09848_),
    .Q(\TRNG.Word_Out[224] ));
 sg13g2_dfrbp_1 _22590_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net5971),
    .D(net1159),
    .Q_N(_09847_),
    .Q(\TRNG.Word_Out[225] ));
 sg13g2_dfrbp_1 _22591_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net5980),
    .D(net3230),
    .Q_N(_09846_),
    .Q(\TRNG.Word_Out[226] ));
 sg13g2_dfrbp_1 _22592_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net5982),
    .D(_01471_),
    .Q_N(_09845_),
    .Q(\TRNG.Word_Out[227] ));
 sg13g2_dfrbp_1 _22593_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net5985),
    .D(_01472_),
    .Q_N(_09844_),
    .Q(\TRNG.Word_Out[228] ));
 sg13g2_dfrbp_1 _22594_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net6000),
    .D(net1209),
    .Q_N(_09843_),
    .Q(\TRNG.Word_Out[229] ));
 sg13g2_dfrbp_1 _22595_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net6000),
    .D(net1742),
    .Q_N(_09842_),
    .Q(\TRNG.Word_Out[230] ));
 sg13g2_dfrbp_1 _22596_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net6053),
    .D(_01475_),
    .Q_N(_09841_),
    .Q(\TRNG.Word_Out[231] ));
 sg13g2_dfrbp_1 _22597_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net6057),
    .D(net1837),
    .Q_N(_09840_),
    .Q(\TRNG.Word_Out[232] ));
 sg13g2_dfrbp_1 _22598_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net6058),
    .D(net2205),
    .Q_N(_09839_),
    .Q(\TRNG.Word_Out[233] ));
 sg13g2_dfrbp_1 _22599_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net6056),
    .D(_01478_),
    .Q_N(_09838_),
    .Q(\TRNG.Word_Out[234] ));
 sg13g2_dfrbp_1 _22600_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net6047),
    .D(net2275),
    .Q_N(_09837_),
    .Q(\TRNG.Word_Out[235] ));
 sg13g2_dfrbp_1 _22601_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net6045),
    .D(net2384),
    .Q_N(_09836_),
    .Q(\TRNG.Word_Out[236] ));
 sg13g2_dfrbp_1 _22602_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net6046),
    .D(_01481_),
    .Q_N(_09835_),
    .Q(\TRNG.Word_Out[237] ));
 sg13g2_dfrbp_1 _22603_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net6024),
    .D(_01482_),
    .Q_N(_09834_),
    .Q(\TRNG.Word_Out[238] ));
 sg13g2_dfrbp_1 _22604_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net6037),
    .D(net2095),
    .Q_N(_09833_),
    .Q(\TRNG.Word_Out[239] ));
 sg13g2_dfrbp_1 _22605_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net6033),
    .D(_01484_),
    .Q_N(_09832_),
    .Q(\TRNG.Word_Out[240] ));
 sg13g2_dfrbp_1 _22606_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net6031),
    .D(net1429),
    .Q_N(_09831_),
    .Q(\TRNG.Word_Out[241] ));
 sg13g2_dfrbp_1 _22607_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net6032),
    .D(net2340),
    .Q_N(_09830_),
    .Q(\TRNG.Word_Out[242] ));
 sg13g2_dfrbp_1 _22608_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net6009),
    .D(_01487_),
    .Q_N(_09829_),
    .Q(\TRNG.Word_Out[243] ));
 sg13g2_dfrbp_1 _22609_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net5956),
    .D(_01488_),
    .Q_N(_09828_),
    .Q(\TRNG.Word_Out[244] ));
 sg13g2_dfrbp_1 _22610_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net5955),
    .D(_01489_),
    .Q_N(_09827_),
    .Q(\TRNG.Word_Out[245] ));
 sg13g2_dfrbp_1 _22611_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net5959),
    .D(net2426),
    .Q_N(_09826_),
    .Q(\TRNG.Word_Out[246] ));
 sg13g2_dfrbp_1 _22612_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net5951),
    .D(_01491_),
    .Q_N(_09825_),
    .Q(\TRNG.Word_Out[247] ));
 sg13g2_dfrbp_1 _22613_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net5937),
    .D(net1561),
    .Q_N(_09824_),
    .Q(\TRNG.Word_Out[248] ));
 sg13g2_dfrbp_1 _22614_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net5932),
    .D(_01493_),
    .Q_N(_09823_),
    .Q(\TRNG.Word_Out[249] ));
 sg13g2_dfrbp_1 _22615_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net5940),
    .D(net1349),
    .Q_N(_09822_),
    .Q(\TRNG.Word_Out[250] ));
 sg13g2_dfrbp_1 _22616_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net5941),
    .D(_01495_),
    .Q_N(_09821_),
    .Q(\TRNG.Word_Out[251] ));
 sg13g2_dfrbp_1 _22617_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net5947),
    .D(net2432),
    .Q_N(_09820_),
    .Q(\TRNG.Word_Out[252] ));
 sg13g2_dfrbp_1 _22618_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net5960),
    .D(_01497_),
    .Q_N(_09819_),
    .Q(\TRNG.Word_Out[253] ));
 sg13g2_dfrbp_1 _22619_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net5960),
    .D(_01498_),
    .Q_N(_09818_),
    .Q(\TRNG.Word_Out[254] ));
 sg13g2_dfrbp_1 _22620_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net5989),
    .D(net1196),
    .Q_N(_09817_),
    .Q(\TRNG.Word_Out[255] ));
 sg13g2_dfrbp_1 _22621_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net5977),
    .D(_01500_),
    .Q_N(_09816_),
    .Q(\TRNG.Word_Out[256] ));
 sg13g2_dfrbp_1 _22622_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net5972),
    .D(net2207),
    .Q_N(_09815_),
    .Q(\TRNG.Word_Out[257] ));
 sg13g2_dfrbp_1 _22623_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net5979),
    .D(_01502_),
    .Q_N(_09814_),
    .Q(\TRNG.Word_Out[258] ));
 sg13g2_dfrbp_1 _22624_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net5979),
    .D(net1852),
    .Q_N(_09813_),
    .Q(\TRNG.Word_Out[259] ));
 sg13g2_dfrbp_1 _22625_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net5983),
    .D(_01504_),
    .Q_N(_09812_),
    .Q(\TRNG.Word_Out[260] ));
 sg13g2_dfrbp_1 _22626_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net5984),
    .D(net1760),
    .Q_N(_09811_),
    .Q(\TRNG.Word_Out[261] ));
 sg13g2_dfrbp_1 _22627_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net5991),
    .D(_01506_),
    .Q_N(_09810_),
    .Q(\TRNG.Word_Out[262] ));
 sg13g2_dfrbp_1 _22628_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net5991),
    .D(_01507_),
    .Q_N(_09809_),
    .Q(\TRNG.Word_Out[263] ));
 sg13g2_dfrbp_1 _22629_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net5991),
    .D(net1372),
    .Q_N(_09808_),
    .Q(\TRNG.Word_Out[264] ));
 sg13g2_dfrbp_1 _22630_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net5991),
    .D(_01509_),
    .Q_N(_09807_),
    .Q(\TRNG.Word_Out[265] ));
 sg13g2_dfrbp_1 _22631_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net5990),
    .D(net1254),
    .Q_N(_09806_),
    .Q(\TRNG.Word_Out[266] ));
 sg13g2_dfrbp_1 _22632_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net5990),
    .D(net1624),
    .Q_N(_09805_),
    .Q(\TRNG.Word_Out[267] ));
 sg13g2_dfrbp_1 _22633_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net5993),
    .D(net1733),
    .Q_N(_09804_),
    .Q(\TRNG.Word_Out[268] ));
 sg13g2_dfrbp_1 _22634_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net5966),
    .D(net3051),
    .Q_N(_09803_),
    .Q(\TRNG.Word_Out[269] ));
 sg13g2_dfrbp_1 _22635_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net5963),
    .D(_01514_),
    .Q_N(_09802_),
    .Q(\TRNG.Word_Out[270] ));
 sg13g2_dfrbp_1 _22636_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net6018),
    .D(net1999),
    .Q_N(_09801_),
    .Q(\TRNG.Word_Out[271] ));
 sg13g2_dfrbp_1 _22637_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net6012),
    .D(_01516_),
    .Q_N(_09800_),
    .Q(\TRNG.Word_Out[272] ));
 sg13g2_dfrbp_1 _22638_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net6013),
    .D(net2082),
    .Q_N(_09799_),
    .Q(\TRNG.Word_Out[273] ));
 sg13g2_dfrbp_1 _22639_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net6013),
    .D(net2297),
    .Q_N(_09798_),
    .Q(\TRNG.Word_Out[274] ));
 sg13g2_dfrbp_1 _22640_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net6009),
    .D(net2437),
    .Q_N(_09797_),
    .Q(\TRNG.Word_Out[275] ));
 sg13g2_dfrbp_1 _22641_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net6008),
    .D(net2640),
    .Q_N(_09796_),
    .Q(\TRNG.Word_Out[276] ));
 sg13g2_dfrbp_1 _22642_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net5953),
    .D(_01521_),
    .Q_N(_09795_),
    .Q(\TRNG.Word_Out[277] ));
 sg13g2_dfrbp_1 _22643_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net5949),
    .D(_01522_),
    .Q_N(_09794_),
    .Q(\TRNG.Word_Out[278] ));
 sg13g2_dfrbp_1 _22644_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net5935),
    .D(net2381),
    .Q_N(_09793_),
    .Q(\TRNG.Word_Out[279] ));
 sg13g2_dfrbp_1 _22645_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net5934),
    .D(_01524_),
    .Q_N(_09792_),
    .Q(\TRNG.Word_Out[280] ));
 sg13g2_dfrbp_1 _22646_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net5909),
    .D(net1139),
    .Q_N(_09791_),
    .Q(\TRNG.Word_Out[281] ));
 sg13g2_dfrbp_1 _22647_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net5907),
    .D(_01526_),
    .Q_N(_09790_),
    .Q(\TRNG.Word_Out[282] ));
 sg13g2_dfrbp_1 _22648_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net5913),
    .D(_01527_),
    .Q_N(_09789_),
    .Q(\TRNG.Word_Out[283] ));
 sg13g2_dfrbp_1 _22649_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net5916),
    .D(net1936),
    .Q_N(_09788_),
    .Q(\TRNG.Word_Out[284] ));
 sg13g2_dfrbp_1 _22650_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net5942),
    .D(_01529_),
    .Q_N(_09787_),
    .Q(\TRNG.Word_Out[285] ));
 sg13g2_dfrbp_1 _22651_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net5970),
    .D(net1411),
    .Q_N(_09786_),
    .Q(\TRNG.Word_Out[286] ));
 sg13g2_dfrbp_1 _22652_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net5970),
    .D(net2166),
    .Q_N(_09785_),
    .Q(\TRNG.Word_Out[287] ));
 sg13g2_dfrbp_1 _22653_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net5923),
    .D(_01532_),
    .Q_N(_09784_),
    .Q(\TRNG.Word_Out[288] ));
 sg13g2_dfrbp_1 _22654_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net5923),
    .D(_01533_),
    .Q_N(_09783_),
    .Q(\TRNG.Word_Out[289] ));
 sg13g2_dfrbp_1 _22655_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net5927),
    .D(net1752),
    .Q_N(_09782_),
    .Q(\TRNG.Word_Out[290] ));
 sg13g2_dfrbp_1 _22656_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net5981),
    .D(_01535_),
    .Q_N(_09781_),
    .Q(\TRNG.Word_Out[291] ));
 sg13g2_dfrbp_1 _22657_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net5981),
    .D(net1213),
    .Q_N(_09780_),
    .Q(\TRNG.Word_Out[292] ));
 sg13g2_dfrbp_1 _22658_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net5985),
    .D(net2291),
    .Q_N(_09779_),
    .Q(\TRNG.Word_Out[293] ));
 sg13g2_dfrbp_1 _22659_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net6005),
    .D(_01538_),
    .Q_N(_09778_),
    .Q(\TRNG.Word_Out[294] ));
 sg13g2_dfrbp_1 _22660_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net6052),
    .D(net1246),
    .Q_N(_09777_),
    .Q(\TRNG.Word_Out[295] ));
 sg13g2_dfrbp_1 _22661_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net6053),
    .D(net1912),
    .Q_N(_09776_),
    .Q(\TRNG.Word_Out[296] ));
 sg13g2_dfrbp_1 _22662_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net6043),
    .D(_01541_),
    .Q_N(_09775_),
    .Q(\TRNG.Word_Out[297] ));
 sg13g2_dfrbp_1 _22663_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net6043),
    .D(net2122),
    .Q_N(_09774_),
    .Q(\TRNG.Word_Out[298] ));
 sg13g2_dfrbp_1 _22664_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net6047),
    .D(net2348),
    .Q_N(_09773_),
    .Q(\TRNG.Word_Out[299] ));
 sg13g2_dfrbp_1 _22665_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net6041),
    .D(net2509),
    .Q_N(_09772_),
    .Q(\TRNG.Word_Out[300] ));
 sg13g2_dfrbp_1 _22666_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net5966),
    .D(_01545_),
    .Q_N(_09771_),
    .Q(\TRNG.Word_Out[301] ));
 sg13g2_dfrbp_1 _22667_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net5966),
    .D(_01546_),
    .Q_N(_09770_),
    .Q(\TRNG.Word_Out[302] ));
 sg13g2_dfrbp_1 _22668_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net6018),
    .D(_01547_),
    .Q_N(_09769_),
    .Q(\TRNG.Word_Out[303] ));
 sg13g2_dfrbp_1 _22669_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net6022),
    .D(net1299),
    .Q_N(_09768_),
    .Q(\TRNG.Word_Out[304] ));
 sg13g2_dfrbp_1 _22670_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net6027),
    .D(_01549_),
    .Q_N(_09767_),
    .Q(\TRNG.Word_Out[305] ));
 sg13g2_dfrbp_1 _22671_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net6027),
    .D(net2350),
    .Q_N(_09766_),
    .Q(\TRNG.Word_Out[306] ));
 sg13g2_dfrbp_1 _22672_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net6008),
    .D(_01551_),
    .Q_N(_09765_),
    .Q(\TRNG.Word_Out[307] ));
 sg13g2_dfrbp_1 _22673_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net5954),
    .D(_01552_),
    .Q_N(_09764_),
    .Q(\TRNG.Word_Out[308] ));
 sg13g2_dfrbp_1 _22674_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net5955),
    .D(_01553_),
    .Q_N(_09763_),
    .Q(\TRNG.Word_Out[309] ));
 sg13g2_dfrbp_1 _22675_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net5952),
    .D(net2035),
    .Q_N(_09762_),
    .Q(\TRNG.Word_Out[310] ));
 sg13g2_dfrbp_1 _22676_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net5938),
    .D(net2137),
    .Q_N(_09761_),
    .Q(\TRNG.Word_Out[311] ));
 sg13g2_dfrbp_1 _22677_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net5932),
    .D(_01556_),
    .Q_N(_09760_),
    .Q(\TRNG.Word_Out[312] ));
 sg13g2_dfrbp_1 _22678_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net5907),
    .D(net1199),
    .Q_N(_09759_),
    .Q(\TRNG.Word_Out[313] ));
 sg13g2_dfrbp_1 _22679_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net5908),
    .D(_01558_),
    .Q_N(_09758_),
    .Q(\TRNG.Word_Out[314] ));
 sg13g2_dfrbp_1 _22680_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net5914),
    .D(_01559_),
    .Q_N(_09757_),
    .Q(\TRNG.Word_Out[315] ));
 sg13g2_dfrbp_1 _22681_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net5945),
    .D(_01560_),
    .Q_N(_09756_),
    .Q(\TRNG.Word_Out[316] ));
 sg13g2_dfrbp_1 _22682_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net5946),
    .D(_01561_),
    .Q_N(_09755_),
    .Q(\TRNG.Word_Out[317] ));
 sg13g2_dfrbp_1 _22683_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net5946),
    .D(_01562_),
    .Q_N(_09754_),
    .Q(\TRNG.Word_Out[318] ));
 sg13g2_dfrbp_1 _22684_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net5975),
    .D(net1291),
    .Q_N(_09753_),
    .Q(\TRNG.Word_Out[319] ));
 sg13g2_dfrbp_1 _22685_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net5970),
    .D(net2555),
    .Q_N(_09752_),
    .Q(\TRNG.Word_Out[320] ));
 sg13g2_dfrbp_1 _22686_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net5972),
    .D(_01565_),
    .Q_N(_09751_),
    .Q(\TRNG.Word_Out[321] ));
 sg13g2_dfrbp_1 _22687_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net5971),
    .D(_01566_),
    .Q_N(_09750_),
    .Q(\TRNG.Word_Out[322] ));
 sg13g2_dfrbp_1 _22688_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net5979),
    .D(_01567_),
    .Q_N(_09749_),
    .Q(\TRNG.Word_Out[323] ));
 sg13g2_dfrbp_1 _22689_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net5983),
    .D(_01568_),
    .Q_N(_09748_),
    .Q(\TRNG.Word_Out[324] ));
 sg13g2_dfrbp_1 _22690_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net5999),
    .D(net1173),
    .Q_N(_09747_),
    .Q(\TRNG.Word_Out[325] ));
 sg13g2_dfrbp_1 _22691_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net6001),
    .D(_01570_),
    .Q_N(_09746_),
    .Q(\TRNG.Word_Out[326] ));
 sg13g2_dfrbp_1 _22692_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net6052),
    .D(_01571_),
    .Q_N(_09745_),
    .Q(\TRNG.Word_Out[327] ));
 sg13g2_dfrbp_1 _22693_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net6053),
    .D(net1394),
    .Q_N(_09744_),
    .Q(\TRNG.Word_Out[328] ));
 sg13g2_dfrbp_1 _22694_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net6057),
    .D(net1917),
    .Q_N(_09743_),
    .Q(\TRNG.Word_Out[329] ));
 sg13g2_dfrbp_1 _22695_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net6050),
    .D(net3099),
    .Q_N(_09742_),
    .Q(\TRNG.Word_Out[330] ));
 sg13g2_dfrbp_1 _22696_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net5997),
    .D(_01575_),
    .Q_N(_09741_),
    .Q(\TRNG.Word_Out[331] ));
 sg13g2_dfrbp_1 _22697_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net6042),
    .D(_01576_),
    .Q_N(_09740_),
    .Q(\TRNG.Word_Out[332] ));
 sg13g2_dfrbp_1 _22698_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net6042),
    .D(_01577_),
    .Q_N(_09739_),
    .Q(\TRNG.Word_Out[333] ));
 sg13g2_dfrbp_1 _22699_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net6020),
    .D(net1155),
    .Q_N(_09738_),
    .Q(\TRNG.Word_Out[334] ));
 sg13g2_dfrbp_1 _22700_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net6023),
    .D(net2102),
    .Q_N(_09737_),
    .Q(\TRNG.Word_Out[335] ));
 sg13g2_dfrbp_1 _22701_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net6013),
    .D(_01580_),
    .Q_N(_09736_),
    .Q(\TRNG.Word_Out[336] ));
 sg13g2_dfrbp_1 _22702_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net6026),
    .D(net2200),
    .Q_N(_09735_),
    .Q(\TRNG.Word_Out[337] ));
 sg13g2_dfrbp_1 _22703_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net6026),
    .D(_01582_),
    .Q_N(_09734_),
    .Q(\TRNG.Word_Out[338] ));
 sg13g2_dfrbp_1 _22704_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net6012),
    .D(net2630),
    .Q_N(_09733_),
    .Q(\TRNG.Word_Out[339] ));
 sg13g2_dfrbp_1 _22705_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net5954),
    .D(_01584_),
    .Q_N(_09732_),
    .Q(\TRNG.Word_Out[340] ));
 sg13g2_dfrbp_1 _22706_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net5950),
    .D(_01585_),
    .Q_N(_09731_),
    .Q(\TRNG.Word_Out[341] ));
 sg13g2_dfrbp_1 _22707_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net5949),
    .D(_01586_),
    .Q_N(_09730_),
    .Q(\TRNG.Word_Out[342] ));
 sg13g2_dfrbp_1 _22708_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net5935),
    .D(net2185),
    .Q_N(_09729_),
    .Q(\TRNG.Word_Out[343] ));
 sg13g2_dfrbp_1 _22709_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net5934),
    .D(_01588_),
    .Q_N(_09728_),
    .Q(\TRNG.Word_Out[344] ));
 sg13g2_dfrbp_1 _22710_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net5908),
    .D(_01589_),
    .Q_N(_09727_),
    .Q(\TRNG.Word_Out[345] ));
 sg13g2_dfrbp_1 _22711_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net5908),
    .D(net1165),
    .Q_N(_09726_),
    .Q(\TRNG.Word_Out[346] ));
 sg13g2_dfrbp_1 _22712_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net5914),
    .D(_01591_),
    .Q_N(_09725_),
    .Q(\TRNG.Word_Out[347] ));
 sg13g2_dfrbp_1 _22713_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net5942),
    .D(_01592_),
    .Q_N(_09724_),
    .Q(\TRNG.Word_Out[348] ));
 sg13g2_dfrbp_1 _22714_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net5969),
    .D(net1186),
    .Q_N(_09723_),
    .Q(\TRNG.Word_Out[349] ));
 sg13g2_dfrbp_1 _22715_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net5974),
    .D(net1382),
    .Q_N(_09722_),
    .Q(\TRNG.Word_Out[350] ));
 sg13g2_dfrbp_1 _22716_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net5974),
    .D(net2077),
    .Q_N(_09721_),
    .Q(\TRNG.Word_Out[351] ));
 sg13g2_dfrbp_1 _22717_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net5977),
    .D(_01596_),
    .Q_N(_09720_),
    .Q(\TRNG.Word_Out[352] ));
 sg13g2_dfrbp_1 _22718_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net5977),
    .D(_01597_),
    .Q_N(_09719_),
    .Q(\TRNG.Word_Out[353] ));
 sg13g2_dfrbp_1 _22719_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net5977),
    .D(net2072),
    .Q_N(_09718_),
    .Q(\TRNG.Word_Out[354] ));
 sg13g2_dfrbp_1 _22720_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net5983),
    .D(_01599_),
    .Q_N(_09717_),
    .Q(\TRNG.Word_Out[355] ));
 sg13g2_dfrbp_1 _22721_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net5986),
    .D(net1188),
    .Q_N(_09716_),
    .Q(\TRNG.Word_Out[356] ));
 sg13g2_dfrbp_1 _22722_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net6000),
    .D(_01601_),
    .Q_N(_09715_),
    .Q(\TRNG.Word_Out[357] ));
 sg13g2_dfrbp_1 _22723_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net6004),
    .D(net1600),
    .Q_N(_09714_),
    .Q(\TRNG.Word_Out[358] ));
 sg13g2_dfrbp_1 _22724_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net6005),
    .D(_01603_),
    .Q_N(_09713_),
    .Q(\TRNG.Word_Out[359] ));
 sg13g2_dfrbp_1 _22725_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net6051),
    .D(net1220),
    .Q_N(_09712_),
    .Q(\TRNG.Word_Out[360] ));
 sg13g2_dfrbp_1 _22726_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net6055),
    .D(_01605_),
    .Q_N(_09711_),
    .Q(\TRNG.Word_Out[361] ));
 sg13g2_dfrbp_1 _22727_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net6043),
    .D(net2589),
    .Q_N(_09710_),
    .Q(\TRNG.Word_Out[362] ));
 sg13g2_dfrbp_1 _22728_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net6042),
    .D(_01607_),
    .Q_N(_09709_),
    .Q(\TRNG.Word_Out[363] ));
 sg13g2_dfrbp_1 _22729_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net6041),
    .D(net1983),
    .Q_N(_09708_),
    .Q(\TRNG.Word_Out[364] ));
 sg13g2_dfrbp_1 _22730_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net6019),
    .D(_01609_),
    .Q_N(_09707_),
    .Q(\TRNG.Word_Out[365] ));
 sg13g2_dfrbp_1 _22731_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net6019),
    .D(net2140),
    .Q_N(_09706_),
    .Q(\TRNG.Word_Out[366] ));
 sg13g2_dfrbp_1 _22732_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net6021),
    .D(net2453),
    .Q_N(_09705_),
    .Q(\TRNG.Word_Out[367] ));
 sg13g2_dfrbp_1 _22733_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net6027),
    .D(_01612_),
    .Q_N(_09704_),
    .Q(\TRNG.Word_Out[368] ));
 sg13g2_dfrbp_1 _22734_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net6031),
    .D(_01613_),
    .Q_N(_09703_),
    .Q(\TRNG.Word_Out[369] ));
 sg13g2_dfrbp_1 _22735_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net6032),
    .D(net1986),
    .Q_N(_09702_),
    .Q(\TRNG.Word_Out[370] ));
 sg13g2_dfrbp_1 _22736_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net6012),
    .D(_01615_),
    .Q_N(_09701_),
    .Q(\TRNG.Word_Out[371] ));
 sg13g2_dfrbp_1 _22737_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net6008),
    .D(net2585),
    .Q_N(_09700_),
    .Q(\TRNG.Word_Out[372] ));
 sg13g2_dfrbp_1 _22738_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net5954),
    .D(_01617_),
    .Q_N(_09699_),
    .Q(\TRNG.Word_Out[373] ));
 sg13g2_dfrbp_1 _22739_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net5949),
    .D(_01618_),
    .Q_N(_09698_),
    .Q(\TRNG.Word_Out[374] ));
 sg13g2_dfrbp_1 _22740_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net5936),
    .D(_01619_),
    .Q_N(_09697_),
    .Q(\TRNG.Word_Out[375] ));
 sg13g2_dfrbp_1 _22741_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net5935),
    .D(_01620_),
    .Q_N(_09696_),
    .Q(\TRNG.Word_Out[376] ));
 sg13g2_dfrbp_1 _22742_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net5932),
    .D(net1179),
    .Q_N(_09695_),
    .Q(\TRNG.Word_Out[377] ));
 sg13g2_dfrbp_1 _22743_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net5908),
    .D(_01622_),
    .Q_N(_09694_),
    .Q(\TRNG.Word_Out[378] ));
 sg13g2_dfrbp_1 _22744_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net5914),
    .D(net2456),
    .Q_N(_09693_),
    .Q(\TRNG.Word_Out[379] ));
 sg13g2_dfrbp_1 _22745_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net5942),
    .D(_01624_),
    .Q_N(_09692_),
    .Q(\TRNG.Word_Out[380] ));
 sg13g2_dfrbp_1 _22746_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net5943),
    .D(_01625_),
    .Q_N(_09691_),
    .Q(\TRNG.Word_Out[381] ));
 sg13g2_dfrbp_1 _22747_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net5974),
    .D(net1205),
    .Q_N(_09690_),
    .Q(\TRNG.Word_Out[382] ));
 sg13g2_dfrbp_1 _22748_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net5975),
    .D(_01627_),
    .Q_N(_09689_),
    .Q(\TRNG.Word_Out[383] ));
 sg13g2_dfrbp_1 _22749_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net5976),
    .D(_01628_),
    .Q_N(_09688_),
    .Q(\TRNG.Word_Out[384] ));
 sg13g2_dfrbp_1 _22750_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net5976),
    .D(net1819),
    .Q_N(_09687_),
    .Q(\TRNG.Word_Out[385] ));
 sg13g2_dfrbp_1 _22751_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net5978),
    .D(net2158),
    .Q_N(_09686_),
    .Q(\TRNG.Word_Out[386] ));
 sg13g2_dfrbp_1 _22752_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net5976),
    .D(_01631_),
    .Q_N(_09685_),
    .Q(\TRNG.Word_Out[387] ));
 sg13g2_dfrbp_1 _22753_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net5976),
    .D(_01632_),
    .Q_N(_09684_),
    .Q(\TRNG.Word_Out[388] ));
 sg13g2_dfrbp_1 _22754_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net5999),
    .D(_01633_),
    .Q_N(_09683_),
    .Q(\TRNG.Word_Out[389] ));
 sg13g2_dfrbp_1 _22755_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net5998),
    .D(net1175),
    .Q_N(_09682_),
    .Q(\TRNG.Word_Out[390] ));
 sg13g2_dfrbp_1 _22756_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net5998),
    .D(net1662),
    .Q_N(_09681_),
    .Q(\TRNG.Word_Out[391] ));
 sg13g2_dfrbp_1 _22757_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net5996),
    .D(net2450),
    .Q_N(_09680_),
    .Q(\TRNG.Word_Out[392] ));
 sg13g2_dfrbp_1 _22758_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net5995),
    .D(_01637_),
    .Q_N(_09679_),
    .Q(\TRNG.Word_Out[393] ));
 sg13g2_dfrbp_1 _22759_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net5995),
    .D(net1233),
    .Q_N(_09678_),
    .Q(\TRNG.Word_Out[394] ));
 sg13g2_dfrbp_1 _22760_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net5990),
    .D(_01639_),
    .Q_N(_09677_),
    .Q(\TRNG.Word_Out[395] ));
 sg13g2_dfrbp_1 _22761_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net5990),
    .D(net1388),
    .Q_N(_09676_),
    .Q(\TRNG.Word_Out[396] ));
 sg13g2_dfrbp_1 _22762_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net5965),
    .D(_01641_),
    .Q_N(_09675_),
    .Q(\TRNG.Word_Out[397] ));
 sg13g2_dfrbp_1 _22763_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net6020),
    .D(net1228),
    .Q_N(_09674_),
    .Q(\TRNG.Word_Out[398] ));
 sg13g2_dfrbp_1 _22764_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net6022),
    .D(net2003),
    .Q_N(_09673_),
    .Q(\TRNG.Word_Out[399] ));
 sg13g2_dfrbp_1 _22765_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net6028),
    .D(_01644_),
    .Q_N(_09672_),
    .Q(\TRNG.Word_Out[400] ));
 sg13g2_dfrbp_1 _22766_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net6029),
    .D(net1472),
    .Q_N(_09671_),
    .Q(\TRNG.Word_Out[401] ));
 sg13g2_dfrbp_1 _22767_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net6027),
    .D(net2295),
    .Q_N(_09670_),
    .Q(\TRNG.Word_Out[402] ));
 sg13g2_dfrbp_1 _22768_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net6012),
    .D(net2908),
    .Q_N(_09669_),
    .Q(\TRNG.Word_Out[403] ));
 sg13g2_dfrbp_1 _22769_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net5954),
    .D(_01648_),
    .Q_N(_09668_),
    .Q(\TRNG.Word_Out[404] ));
 sg13g2_dfrbp_1 _22770_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net5950),
    .D(_01649_),
    .Q_N(_09667_),
    .Q(\TRNG.Word_Out[405] ));
 sg13g2_dfrbp_1 _22771_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net5949),
    .D(net1875),
    .Q_N(_09666_),
    .Q(\TRNG.Word_Out[406] ));
 sg13g2_dfrbp_1 _22772_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net5935),
    .D(net2535),
    .Q_N(_09665_),
    .Q(\TRNG.Word_Out[407] ));
 sg13g2_dfrbp_1 _22773_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net5934),
    .D(_01652_),
    .Q_N(_09664_),
    .Q(\TRNG.Word_Out[408] ));
 sg13g2_dfrbp_1 _22774_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net5909),
    .D(_01653_),
    .Q_N(_09663_),
    .Q(\TRNG.Word_Out[409] ));
 sg13g2_dfrbp_1 _22775_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net5908),
    .D(net1169),
    .Q_N(_09662_),
    .Q(\TRNG.Word_Out[410] ));
 sg13g2_dfrbp_1 _22776_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net5940),
    .D(net2944),
    .Q_N(_09661_),
    .Q(\TRNG.Word_Out[411] ));
 sg13g2_dfrbp_1 _22777_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net5942),
    .D(_01656_),
    .Q_N(_09660_),
    .Q(\TRNG.Word_Out[412] ));
 sg13g2_dfrbp_1 _22778_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net5960),
    .D(_01657_),
    .Q_N(_09659_),
    .Q(\TRNG.Word_Out[413] ));
 sg13g2_dfrbp_1 _22779_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net5961),
    .D(net1399),
    .Q_N(_09658_),
    .Q(\TRNG.Word_Out[414] ));
 sg13g2_dfrbp_1 _22780_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net6037),
    .D(_01659_),
    .Q_N(_09657_),
    .Q(\TRNG.Word_Out[415] ));
 sg13g2_dfrbp_1 _22781_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net6037),
    .D(net2031),
    .Q_N(_09656_),
    .Q(\TRNG.Word_Out[416] ));
 sg13g2_dfrbp_1 _22782_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net6063),
    .D(_01661_),
    .Q_N(_09655_),
    .Q(\TRNG.Word_Out[417] ));
 sg13g2_dfrbp_1 _22783_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net6061),
    .D(net2162),
    .Q_N(_09654_),
    .Q(\TRNG.Word_Out[418] ));
 sg13g2_dfrbp_1 _22784_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net6061),
    .D(net2371),
    .Q_N(_09653_),
    .Q(\TRNG.Word_Out[419] ));
 sg13g2_dfrbp_1 _22785_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net6065),
    .D(_01664_),
    .Q_N(_09652_),
    .Q(\TRNG.Word_Out[420] ));
 sg13g2_dfrbp_1 _22786_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net6064),
    .D(net1634),
    .Q_N(_09651_),
    .Q(\TRNG.Word_Out[421] ));
 sg13g2_dfrbp_1 _22787_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net6055),
    .D(_01666_),
    .Q_N(_09650_),
    .Q(\TRNG.Word_Out[422] ));
 sg13g2_dfrbp_1 _22788_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net6056),
    .D(_01667_),
    .Q_N(_09649_),
    .Q(\TRNG.Word_Out[423] ));
 sg13g2_dfrbp_1 _22789_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net6060),
    .D(net2025),
    .Q_N(_09648_),
    .Q(\TRNG.Word_Out[424] ));
 sg13g2_dfrbp_1 _22790_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net6060),
    .D(net2232),
    .Q_N(_09647_),
    .Q(\TRNG.Word_Out[425] ));
 sg13g2_dfrbp_1 _22791_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net6060),
    .D(_01670_),
    .Q_N(_09646_),
    .Q(\TRNG.Word_Out[426] ));
 sg13g2_dfrbp_1 _22792_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net6060),
    .D(net1470),
    .Q_N(_09645_),
    .Q(\TRNG.Word_Out[427] ));
 sg13g2_dfrbp_1 _22793_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net6037),
    .D(_01672_),
    .Q_N(_09644_),
    .Q(\TRNG.Word_Out[428] ));
 sg13g2_dfrbp_1 _22794_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net6037),
    .D(net1651),
    .Q_N(_09643_),
    .Q(\TRNG.Word_Out[429] ));
 sg13g2_dfrbp_1 _22795_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net6037),
    .D(_01674_),
    .Q_N(_09642_),
    .Q(\TRNG.Word_Out[430] ));
 sg13g2_dfrbp_1 _22796_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net6038),
    .D(net1796),
    .Q_N(_09641_),
    .Q(\TRNG.Word_Out[431] ));
 sg13g2_dfrbp_1 _22797_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net6038),
    .D(net2133),
    .Q_N(_09640_),
    .Q(\TRNG.Word_Out[432] ));
 sg13g2_dfrbp_1 _22798_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net6033),
    .D(_01677_),
    .Q_N(_09639_),
    .Q(\TRNG.Word_Out[433] ));
 sg13g2_dfrbp_1 _22799_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net6033),
    .D(_01678_),
    .Q_N(_09638_),
    .Q(\TRNG.Word_Out[434] ));
 sg13g2_dfrbp_1 _22800_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net6032),
    .D(_01679_),
    .Q_N(_09637_),
    .Q(\TRNG.Word_Out[435] ));
 sg13g2_dfrbp_1 _22801_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net6032),
    .D(net1805),
    .Q_N(_09636_),
    .Q(\TRNG.Word_Out[436] ));
 sg13g2_dfrbp_1 _22802_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net6034),
    .D(_01681_),
    .Q_N(_09635_),
    .Q(\TRNG.Word_Out[437] ));
 sg13g2_dfrbp_1 _22803_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net6033),
    .D(_01682_),
    .Q_N(_09634_),
    .Q(\TRNG.Word_Out[438] ));
 sg13g2_dfrbp_1 _22804_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net6038),
    .D(net2027),
    .Q_N(_09633_),
    .Q(\TRNG.Word_Out[439] ));
 sg13g2_dfrbp_1 _22805_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net6039),
    .D(_01684_),
    .Q_N(_09632_),
    .Q(\TRNG.Word_Out[440] ));
 sg13g2_dfrbp_1 _22806_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net6061),
    .D(_01685_),
    .Q_N(_09631_),
    .Q(\TRNG.Word_Out[441] ));
 sg13g2_dfrbp_1 _22807_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net6061),
    .D(net2117),
    .Q_N(_09630_),
    .Q(\TRNG.Word_Out[442] ));
 sg13g2_dfrbp_1 _22808_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net6062),
    .D(_01687_),
    .Q_N(_09629_),
    .Q(\TRNG.Word_Out[443] ));
 sg13g2_dfrbp_1 _22809_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net6061),
    .D(net2164),
    .Q_N(_09628_),
    .Q(\TRNG.Word_Out[444] ));
 sg13g2_dfrbp_1 _22810_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net6064),
    .D(_01689_),
    .Q_N(_09627_),
    .Q(\TRNG.Word_Out[445] ));
 sg13g2_dfrbp_1 _22811_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net6064),
    .D(net2218),
    .Q_N(_11068_),
    .Q(\TRNG.Word_Out[446] ));
 sg13g2_dfrbp_1 _22812_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net5902),
    .D(_02160_),
    .Q_N(_11069_),
    .Q(\TRNG.raw_byte[0] ));
 sg13g2_dfrbp_1 _22813_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net5905),
    .D(_02161_),
    .Q_N(_11070_),
    .Q(\TRNG.raw_byte[1] ));
 sg13g2_dfrbp_1 _22814_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net5902),
    .D(net2870),
    .Q_N(_11071_),
    .Q(\TRNG.raw_byte[2] ));
 sg13g2_dfrbp_1 _22815_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net5902),
    .D(_02163_),
    .Q_N(_11072_),
    .Q(\TRNG.raw_byte[3] ));
 sg13g2_dfrbp_1 _22816_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net5902),
    .D(_02164_),
    .Q_N(_11073_),
    .Q(\TRNG.raw_byte[4] ));
 sg13g2_dfrbp_1 _22817_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net5902),
    .D(_02165_),
    .Q_N(_11074_),
    .Q(\TRNG.raw_byte[5] ));
 sg13g2_dfrbp_1 _22818_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net5902),
    .D(_02166_),
    .Q_N(_11075_),
    .Q(\TRNG.raw_byte[6] ));
 sg13g2_dfrbp_1 _22819_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net5902),
    .D(net2529),
    .Q_N(_09626_),
    .Q(\TRNG.raw_byte[7] ));
 sg13g2_dfrbp_1 _22820_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net5904),
    .D(_01691_),
    .Q_N(_11076_),
    .Q(\TRNG.discard ));
 sg13g2_dfrbp_1 _22821_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net5900),
    .D(net1),
    .Q_N(_11077_),
    .Q(\TRNG.ctrl_mode_sync[0] ));
 sg13g2_dfrbp_1 _22822_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net5900),
    .D(net1129),
    .Q_N(_00121_),
    .Q(\TRNG.ctrl_mode_sync[1] ));
 sg13g2_dfrbp_1 _22823_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net5992),
    .D(_01692_),
    .Q_N(_09625_),
    .Q(\TRNG.Padded_Out[64] ));
 sg13g2_dfrbp_1 _22824_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net5920),
    .D(net1839),
    .Q_N(_09624_),
    .Q(\TRNG.Padded_Out[65] ));
 sg13g2_dfrbp_1 _22825_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net5920),
    .D(net1951),
    .Q_N(_09623_),
    .Q(\TRNG.Padded_Out[66] ));
 sg13g2_dfrbp_1 _22826_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net5976),
    .D(_01695_),
    .Q_N(_09622_),
    .Q(\TRNG.Padded_Out[67] ));
 sg13g2_dfrbp_1 _22827_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net5927),
    .D(net1828),
    .Q_N(_09621_),
    .Q(\TRNG.Padded_Out[68] ));
 sg13g2_dfrbp_1 _22828_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net5985),
    .D(net1403),
    .Q_N(_09620_),
    .Q(\TRNG.Padded_Out[69] ));
 sg13g2_dfrbp_1 _22829_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net5985),
    .D(net1758),
    .Q_N(_09619_),
    .Q(\TRNG.Padded_Out[70] ));
 sg13g2_dfrbp_1 _22830_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net6002),
    .D(net1700),
    .Q_N(_09618_),
    .Q(\TRNG.Padded_Out[71] ));
 sg13g2_dfrbp_1 _22831_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net6050),
    .D(_01700_),
    .Q_N(_09617_),
    .Q(\TRNG.Padded_Out[72] ));
 sg13g2_dfrbp_1 _22832_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net6003),
    .D(net1554),
    .Q_N(_09616_),
    .Q(\TRNG.Padded_Out[73] ));
 sg13g2_dfrbp_1 _22833_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net5995),
    .D(net1441),
    .Q_N(_09615_),
    .Q(\TRNG.Padded_Out[74] ));
 sg13g2_dfrbp_1 _22834_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net6044),
    .D(net1675),
    .Q_N(_09614_),
    .Q(\TRNG.Padded_Out[75] ));
 sg13g2_dfrbp_1 _22835_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net5994),
    .D(net1953),
    .Q_N(_09613_),
    .Q(\TRNG.Padded_Out[76] ));
 sg13g2_dfrbp_1 _22836_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net5965),
    .D(net1990),
    .Q_N(_09612_),
    .Q(\TRNG.Padded_Out[77] ));
 sg13g2_dfrbp_1 _22837_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net5965),
    .D(_01706_),
    .Q_N(_09611_),
    .Q(\TRNG.Padded_Out[78] ));
 sg13g2_dfrbp_1 _22838_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net5964),
    .D(net1260),
    .Q_N(_09610_),
    .Q(\TRNG.Padded_Out[79] ));
 sg13g2_dfrbp_1 _22839_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net6021),
    .D(_01708_),
    .Q_N(_09609_),
    .Q(\TRNG.Padded_Out[80] ));
 sg13g2_dfrbp_1 _22840_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net6022),
    .D(net1885),
    .Q_N(_09608_),
    .Q(\TRNG.Padded_Out[81] ));
 sg13g2_dfrbp_1 _22841_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net6026),
    .D(_01710_),
    .Q_N(_09607_),
    .Q(\TRNG.Padded_Out[82] ));
 sg13g2_dfrbp_1 _22842_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net6015),
    .D(net1698),
    .Q_N(_09606_),
    .Q(\TRNG.Padded_Out[83] ));
 sg13g2_dfrbp_1 _22843_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net6009),
    .D(net1538),
    .Q_N(_09605_),
    .Q(\TRNG.Padded_Out[84] ));
 sg13g2_dfrbp_1 _22844_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net6008),
    .D(net1540),
    .Q_N(_09604_),
    .Q(\TRNG.Padded_Out[85] ));
 sg13g2_dfrbp_1 _22845_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net5953),
    .D(net1419),
    .Q_N(_09603_),
    .Q(\TRNG.Padded_Out[86] ));
 sg13g2_dfrbp_1 _22846_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net5949),
    .D(net1519),
    .Q_N(_09602_),
    .Q(\TRNG.Padded_Out[87] ));
 sg13g2_dfrbp_1 _22847_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net5935),
    .D(net1293),
    .Q_N(_09601_),
    .Q(\TRNG.Padded_Out[88] ));
 sg13g2_dfrbp_1 _22848_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net5937),
    .D(_01717_),
    .Q_N(_09600_),
    .Q(\TRNG.Padded_Out[89] ));
 sg13g2_dfrbp_1 _22849_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net5937),
    .D(net1401),
    .Q_N(_09599_),
    .Q(\TRNG.Padded_Out[90] ));
 sg13g2_dfrbp_1 _22850_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net5907),
    .D(net2067),
    .Q_N(_09598_),
    .Q(\TRNG.Padded_Out[91] ));
 sg13g2_dfrbp_1 _22851_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net5913),
    .D(net2315),
    .Q_N(_09597_),
    .Q(\TRNG.Padded_Out[92] ));
 sg13g2_dfrbp_1 _22852_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net5916),
    .D(net1390),
    .Q_N(_09596_),
    .Q(\TRNG.Padded_Out[93] ));
 sg13g2_dfrbp_1 _22853_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net5915),
    .D(_01722_),
    .Q_N(_09595_),
    .Q(\TRNG.Padded_Out[94] ));
 sg13g2_dfrbp_1 _22854_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net5921),
    .D(_01723_),
    .Q_N(_09594_),
    .Q(\TRNG.Padded_Out[95] ));
 sg13g2_dfrbp_1 _22855_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net5921),
    .D(net2086),
    .Q_N(_09593_),
    .Q(\TRNG.Padded_Out[96] ));
 sg13g2_dfrbp_1 _22856_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net5924),
    .D(net2187),
    .Q_N(_09592_),
    .Q(\TRNG.Padded_Out[97] ));
 sg13g2_dfrbp_1 _22857_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net5924),
    .D(net2051),
    .Q_N(_09591_),
    .Q(\TRNG.Padded_Out[98] ));
 sg13g2_dfrbp_1 _22858_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net5927),
    .D(net1958),
    .Q_N(_09590_),
    .Q(\TRNG.Padded_Out[99] ));
 sg13g2_dfrbp_1 _22859_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net5928),
    .D(net1846),
    .Q_N(_09589_),
    .Q(\TRNG.Padded_Out[100] ));
 sg13g2_dfrbp_1 _22860_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net5982),
    .D(_01729_),
    .Q_N(_09588_),
    .Q(\TRNG.Padded_Out[101] ));
 sg13g2_dfrbp_1 _22861_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net5985),
    .D(_01730_),
    .Q_N(_09587_),
    .Q(\TRNG.Padded_Out[102] ));
 sg13g2_dfrbp_1 _22862_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net6004),
    .D(_01731_),
    .Q_N(_09586_),
    .Q(\TRNG.Padded_Out[103] ));
 sg13g2_dfrbp_1 _22863_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net6005),
    .D(net2120),
    .Q_N(_09585_),
    .Q(\TRNG.Padded_Out[104] ));
 sg13g2_dfrbp_1 _22864_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net6057),
    .D(_01733_),
    .Q_N(_09584_),
    .Q(\TRNG.Padded_Out[105] ));
 sg13g2_dfrbp_1 _22865_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net6058),
    .D(net2150),
    .Q_N(_09583_),
    .Q(\TRNG.Padded_Out[106] ));
 sg13g2_dfrbp_1 _22866_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net6055),
    .D(net1762),
    .Q_N(_09582_),
    .Q(\TRNG.Padded_Out[107] ));
 sg13g2_dfrbp_1 _22867_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net6048),
    .D(net2089),
    .Q_N(_09581_),
    .Q(\TRNG.Padded_Out[108] ));
 sg13g2_dfrbp_1 _22868_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net6046),
    .D(net2183),
    .Q_N(_09580_),
    .Q(\TRNG.Padded_Out[109] ));
 sg13g2_dfrbp_1 _22869_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net6046),
    .D(_01738_),
    .Q_N(_09579_),
    .Q(\TRNG.Padded_Out[110] ));
 sg13g2_dfrbp_1 _22870_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net6023),
    .D(net1721),
    .Q_N(_09578_),
    .Q(\TRNG.Padded_Out[111] ));
 sg13g2_dfrbp_1 _22871_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net6023),
    .D(net1862),
    .Q_N(_09577_),
    .Q(\TRNG.Padded_Out[112] ));
 sg13g2_dfrbp_1 _22872_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net6036),
    .D(net1660),
    .Q_N(_09576_),
    .Q(\TRNG.Padded_Out[113] ));
 sg13g2_dfrbp_1 _22873_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net6029),
    .D(net1332),
    .Q_N(_09575_),
    .Q(\TRNG.Padded_Out[114] ));
 sg13g2_dfrbp_1 _22874_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net6015),
    .D(net1831),
    .Q_N(_09574_),
    .Q(\TRNG.Padded_Out[115] ));
 sg13g2_dfrbp_1 _22875_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net6010),
    .D(net1433),
    .Q_N(_09573_),
    .Q(\TRNG.Padded_Out[116] ));
 sg13g2_dfrbp_1 _22876_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net5956),
    .D(net1694),
    .Q_N(_09572_),
    .Q(\TRNG.Padded_Out[117] ));
 sg13g2_dfrbp_1 _22877_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net5955),
    .D(_01746_),
    .Q_N(_09571_),
    .Q(\TRNG.Padded_Out[118] ));
 sg13g2_dfrbp_1 _22878_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net5952),
    .D(net1679),
    .Q_N(_09570_),
    .Q(\TRNG.Padded_Out[119] ));
 sg13g2_dfrbp_1 _22879_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net5951),
    .D(net1563),
    .Q_N(_09569_),
    .Q(\TRNG.Padded_Out[120] ));
 sg13g2_dfrbp_1 _22880_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net5933),
    .D(net1449),
    .Q_N(_09568_),
    .Q(\TRNG.Padded_Out[121] ));
 sg13g2_dfrbp_1 _22881_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net5933),
    .D(net1710),
    .Q_N(_09567_),
    .Q(\TRNG.Padded_Out[122] ));
 sg13g2_dfrbp_1 _22882_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net5913),
    .D(net1792),
    .Q_N(_09566_),
    .Q(\TRNG.Padded_Out[123] ));
 sg13g2_dfrbp_1 _22883_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net5916),
    .D(net1934),
    .Q_N(_09565_),
    .Q(\TRNG.Padded_Out[124] ));
 sg13g2_dfrbp_1 _22884_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net5916),
    .D(_01753_),
    .Q_N(_09564_),
    .Q(\TRNG.Padded_Out[125] ));
 sg13g2_dfrbp_1 _22885_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net5943),
    .D(net1976),
    .Q_N(_09563_),
    .Q(\TRNG.Padded_Out[126] ));
 sg13g2_dfrbp_1 _22886_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net5969),
    .D(net1773),
    .Q_N(_09562_),
    .Q(\TRNG.Padded_Out[127] ));
 sg13g2_dfrbp_1 _22887_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net5921),
    .D(_01756_),
    .Q_N(_09561_),
    .Q(\TRNG.Padded_Out[128] ));
 sg13g2_dfrbp_1 _22888_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net5923),
    .D(net2063),
    .Q_N(_09560_),
    .Q(\TRNG.Padded_Out[129] ));
 sg13g2_dfrbp_1 _22889_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net5926),
    .D(net1787),
    .Q_N(_09559_),
    .Q(\TRNG.Padded_Out[130] ));
 sg13g2_dfrbp_1 _22890_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net5926),
    .D(net1658),
    .Q_N(_09558_),
    .Q(\TRNG.Padded_Out[131] ));
 sg13g2_dfrbp_1 _22891_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net5929),
    .D(_01760_),
    .Q_N(_09557_),
    .Q(\TRNG.Padded_Out[132] ));
 sg13g2_dfrbp_1 _22892_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net5928),
    .D(net1584),
    .Q_N(_09556_),
    .Q(\TRNG.Padded_Out[133] ));
 sg13g2_dfrbp_1 _22893_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net6001),
    .D(_01762_),
    .Q_N(_09555_),
    .Q(\TRNG.Padded_Out[134] ));
 sg13g2_dfrbp_1 _22894_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net6005),
    .D(_01763_),
    .Q_N(_09554_),
    .Q(\TRNG.Padded_Out[135] ));
 sg13g2_dfrbp_1 _22895_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net6052),
    .D(_01764_),
    .Q_N(_09553_),
    .Q(\TRNG.Padded_Out[136] ));
 sg13g2_dfrbp_1 _22896_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net6053),
    .D(_01765_),
    .Q_N(_09552_),
    .Q(\TRNG.Padded_Out[137] ));
 sg13g2_dfrbp_1 _22897_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net6056),
    .D(net1873),
    .Q_N(_09551_),
    .Q(\TRNG.Padded_Out[138] ));
 sg13g2_dfrbp_1 _22898_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net6047),
    .D(net1686),
    .Q_N(_09550_),
    .Q(\TRNG.Padded_Out[139] ));
 sg13g2_dfrbp_1 _22899_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net6048),
    .D(net1521),
    .Q_N(_09549_),
    .Q(\TRNG.Padded_Out[140] ));
 sg13g2_dfrbp_1 _22900_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net6045),
    .D(net1248),
    .Q_N(_09548_),
    .Q(\TRNG.Padded_Out[141] ));
 sg13g2_dfrbp_1 _22901_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net5965),
    .D(net1376),
    .Q_N(_09547_),
    .Q(\TRNG.Padded_Out[142] ));
 sg13g2_dfrbp_1 _22902_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net6018),
    .D(_01771_),
    .Q_N(_09546_),
    .Q(\TRNG.Padded_Out[143] ));
 sg13g2_dfrbp_1 _22903_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net6022),
    .D(net1431),
    .Q_N(_09545_),
    .Q(\TRNG.Padded_Out[144] ));
 sg13g2_dfrbp_1 _22904_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net6035),
    .D(net1235),
    .Q_N(_09544_),
    .Q(\TRNG.Padded_Out[145] ));
 sg13g2_dfrbp_1 _22905_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net6035),
    .D(net1365),
    .Q_N(_09543_),
    .Q(\TRNG.Padded_Out[146] ));
 sg13g2_dfrbp_1 _22906_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net6015),
    .D(net1466),
    .Q_N(_09542_),
    .Q(\TRNG.Padded_Out[147] ));
 sg13g2_dfrbp_1 _22907_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net6010),
    .D(net1781),
    .Q_N(_09541_),
    .Q(\TRNG.Padded_Out[148] ));
 sg13g2_dfrbp_1 _22908_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net6011),
    .D(net1576),
    .Q_N(_09540_),
    .Q(\TRNG.Padded_Out[149] ));
 sg13g2_dfrbp_1 _22909_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net5963),
    .D(net1946),
    .Q_N(_09539_),
    .Q(\TRNG.Padded_Out[150] ));
 sg13g2_dfrbp_1 _22910_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net5952),
    .D(net1735),
    .Q_N(_09538_),
    .Q(\TRNG.Padded_Out[151] ));
 sg13g2_dfrbp_1 _22911_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net5951),
    .D(net1308),
    .Q_N(_09537_),
    .Q(\TRNG.Padded_Out[152] ));
 sg13g2_dfrbp_1 _22912_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net5937),
    .D(_01781_),
    .Q_N(_09536_),
    .Q(\TRNG.Padded_Out[153] ));
 sg13g2_dfrbp_1 _22913_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net5945),
    .D(net1374),
    .Q_N(_09535_),
    .Q(\TRNG.Padded_Out[154] ));
 sg13g2_dfrbp_1 _22914_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net5913),
    .D(net1320),
    .Q_N(_09534_),
    .Q(\TRNG.Padded_Out[155] ));
 sg13g2_dfrbp_1 _22915_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net5911),
    .D(net1895),
    .Q_N(_09533_),
    .Q(\TRNG.Padded_Out[156] ));
 sg13g2_dfrbp_1 _22916_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net5915),
    .D(net2057),
    .Q_N(_09532_),
    .Q(\TRNG.Padded_Out[157] ));
 sg13g2_dfrbp_1 _22917_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net5915),
    .D(_01786_),
    .Q_N(_09531_),
    .Q(\TRNG.Padded_Out[158] ));
 sg13g2_dfrbp_1 _22918_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net5922),
    .D(net1268),
    .Q_N(_09530_),
    .Q(\TRNG.Padded_Out[159] ));
 sg13g2_dfrbp_1 _22919_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net5969),
    .D(_01788_),
    .Q_N(_09529_),
    .Q(\TRNG.Padded_Out[160] ));
 sg13g2_dfrbp_1 _22920_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net5969),
    .D(net1527),
    .Q_N(_09528_),
    .Q(\TRNG.Padded_Out[161] ));
 sg13g2_dfrbp_1 _22921_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net5971),
    .D(net1588),
    .Q_N(_09527_),
    .Q(\TRNG.Padded_Out[162] ));
 sg13g2_dfrbp_1 _22922_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net5980),
    .D(net1604),
    .Q_N(_09526_),
    .Q(\TRNG.Padded_Out[163] ));
 sg13g2_dfrbp_1 _22923_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net5979),
    .D(net1328),
    .Q_N(_09525_),
    .Q(\TRNG.Padded_Out[164] ));
 sg13g2_dfrbp_1 _22924_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net5983),
    .D(_01793_),
    .Q_N(_09524_),
    .Q(\TRNG.Padded_Out[165] ));
 sg13g2_dfrbp_1 _22925_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net5999),
    .D(net2013),
    .Q_N(_09523_),
    .Q(\TRNG.Padded_Out[166] ));
 sg13g2_dfrbp_1 _22926_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net5998),
    .D(net1708),
    .Q_N(_09522_),
    .Q(\TRNG.Padded_Out[167] ));
 sg13g2_dfrbp_1 _22927_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net6003),
    .D(_01796_),
    .Q_N(_09521_),
    .Q(\TRNG.Padded_Out[168] ));
 sg13g2_dfrbp_1 _22928_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net6050),
    .D(net1611),
    .Q_N(_09520_),
    .Q(\TRNG.Padded_Out[169] ));
 sg13g2_dfrbp_1 _22929_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net6055),
    .D(net1690),
    .Q_N(_09519_),
    .Q(\TRNG.Padded_Out[170] ));
 sg13g2_dfrbp_1 _22930_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net6043),
    .D(net1850),
    .Q_N(_09518_),
    .Q(\TRNG.Padded_Out[171] ));
 sg13g2_dfrbp_1 _22931_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net6042),
    .D(net1423),
    .Q_N(_09517_),
    .Q(\TRNG.Padded_Out[172] ));
 sg13g2_dfrbp_1 _22932_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net5993),
    .D(net1997),
    .Q_N(_09516_),
    .Q(\TRNG.Padded_Out[173] ));
 sg13g2_dfrbp_1 _22933_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net5966),
    .D(net2091),
    .Q_N(_09515_),
    .Q(\TRNG.Padded_Out[174] ));
 sg13g2_dfrbp_1 _22934_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net5964),
    .D(net1713),
    .Q_N(_09514_),
    .Q(\TRNG.Padded_Out[175] ));
 sg13g2_dfrbp_1 _22935_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net6018),
    .D(net1507),
    .Q_N(_09513_),
    .Q(\TRNG.Padded_Out[176] ));
 sg13g2_dfrbp_1 _22936_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net6022),
    .D(_01805_),
    .Q_N(_09512_),
    .Q(\TRNG.Padded_Out[177] ));
 sg13g2_dfrbp_1 _22937_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net6028),
    .D(_01806_),
    .Q_N(_09511_),
    .Q(\TRNG.Padded_Out[178] ));
 sg13g2_dfrbp_1 _22938_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net6014),
    .D(net1546),
    .Q_N(_09510_),
    .Q(\TRNG.Padded_Out[179] ));
 sg13g2_dfrbp_1 _22939_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net6010),
    .D(net1262),
    .Q_N(_09509_),
    .Q(\TRNG.Padded_Out[180] ));
 sg13g2_dfrbp_1 _22940_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net6011),
    .D(net1492),
    .Q_N(_09508_),
    .Q(\TRNG.Padded_Out[181] ));
 sg13g2_dfrbp_1 _22941_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net5955),
    .D(net1671),
    .Q_N(_09507_),
    .Q(\TRNG.Padded_Out[182] ));
 sg13g2_dfrbp_1 _22942_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net5949),
    .D(net1809),
    .Q_N(_09506_),
    .Q(\TRNG.Padded_Out[183] ));
 sg13g2_dfrbp_1 _22943_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net5951),
    .D(net1396),
    .Q_N(_09505_),
    .Q(\TRNG.Padded_Out[184] ));
 sg13g2_dfrbp_1 _22944_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net5934),
    .D(net1271),
    .Q_N(_09504_),
    .Q(\TRNG.Padded_Out[185] ));
 sg13g2_dfrbp_1 _22945_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net5907),
    .D(net1682),
    .Q_N(_09503_),
    .Q(\TRNG.Padded_Out[186] ));
 sg13g2_dfrbp_1 _22946_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net5910),
    .D(net2049),
    .Q_N(_09502_),
    .Q(\TRNG.Padded_Out[187] ));
 sg13g2_dfrbp_1 _22947_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net5911),
    .D(net1871),
    .Q_N(_09501_),
    .Q(\TRNG.Padded_Out[188] ));
 sg13g2_dfrbp_1 _22948_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net5912),
    .D(net1511),
    .Q_N(_09500_),
    .Q(\TRNG.Padded_Out[189] ));
 sg13g2_dfrbp_1 _22949_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net5912),
    .D(_01818_),
    .Q_N(_09499_),
    .Q(\TRNG.Padded_Out[190] ));
 sg13g2_dfrbp_1 _22950_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net5921),
    .D(net2080),
    .Q_N(_09498_),
    .Q(\TRNG.Padded_Out[191] ));
 sg13g2_dfrbp_1 _22951_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net5921),
    .D(_01820_),
    .Q_N(_09497_),
    .Q(\TRNG.Padded_Out[192] ));
 sg13g2_dfrbp_1 _22952_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net5923),
    .D(_01821_),
    .Q_N(_09496_),
    .Q(\TRNG.Padded_Out[193] ));
 sg13g2_dfrbp_1 _22953_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net5924),
    .D(net1794),
    .Q_N(_09495_),
    .Q(\TRNG.Padded_Out[194] ));
 sg13g2_dfrbp_1 _22954_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net5926),
    .D(net1484),
    .Q_N(_09494_),
    .Q(\TRNG.Padded_Out[195] ));
 sg13g2_dfrbp_1 _22955_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net5928),
    .D(_01824_),
    .Q_N(_09493_),
    .Q(\TRNG.Padded_Out[196] ));
 sg13g2_dfrbp_1 _22956_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net5982),
    .D(net1415),
    .Q_N(_09492_),
    .Q(\TRNG.Padded_Out[197] ));
 sg13g2_dfrbp_1 _22957_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net5999),
    .D(_01826_),
    .Q_N(_09491_),
    .Q(\TRNG.Padded_Out[198] ));
 sg13g2_dfrbp_1 _22958_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net5998),
    .D(net1673),
    .Q_N(_09490_),
    .Q(\TRNG.Padded_Out[199] ));
 sg13g2_dfrbp_1 _22959_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net6003),
    .D(_01828_),
    .Q_N(_09489_),
    .Q(\TRNG.Padded_Out[200] ));
 sg13g2_dfrbp_1 _22960_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net6050),
    .D(net1835),
    .Q_N(_09488_),
    .Q(\TRNG.Padded_Out[201] ));
 sg13g2_dfrbp_1 _22961_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net5996),
    .D(net1409),
    .Q_N(_09487_),
    .Q(\TRNG.Padded_Out[202] ));
 sg13g2_dfrbp_1 _22962_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net6044),
    .D(_01831_),
    .Q_N(_09486_),
    .Q(\TRNG.Padded_Out[203] ));
 sg13g2_dfrbp_1 _22963_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net6041),
    .D(net1480),
    .Q_N(_09485_),
    .Q(\TRNG.Padded_Out[204] ));
 sg13g2_dfrbp_1 _22964_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net6045),
    .D(net1940),
    .Q_N(_09484_),
    .Q(\TRNG.Padded_Out[205] ));
 sg13g2_dfrbp_1 _22965_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net6041),
    .D(_01834_),
    .Q_N(_09483_),
    .Q(\TRNG.Padded_Out[206] ));
 sg13g2_dfrbp_1 _22966_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net6023),
    .D(net1622),
    .Q_N(_09482_),
    .Q(\TRNG.Padded_Out[207] ));
 sg13g2_dfrbp_1 _22967_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net6024),
    .D(net1744),
    .Q_N(_09481_),
    .Q(\TRNG.Padded_Out[208] ));
 sg13g2_dfrbp_1 _22968_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net6035),
    .D(net2053),
    .Q_N(_09480_),
    .Q(\TRNG.Padded_Out[209] ));
 sg13g2_dfrbp_1 _22969_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net6028),
    .D(net1768),
    .Q_N(_09479_),
    .Q(\TRNG.Padded_Out[210] ));
 sg13g2_dfrbp_1 _22970_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net6029),
    .D(net2338),
    .Q_N(_09478_),
    .Q(\TRNG.Padded_Out[211] ));
 sg13g2_dfrbp_1 _22971_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net6010),
    .D(net1756),
    .Q_N(_09477_),
    .Q(\TRNG.Padded_Out[212] ));
 sg13g2_dfrbp_1 _22972_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net6011),
    .D(net1314),
    .Q_N(_09476_),
    .Q(\TRNG.Padded_Out[213] ));
 sg13g2_dfrbp_1 _22973_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net5963),
    .D(_01842_),
    .Q_N(_09475_),
    .Q(\TRNG.Padded_Out[214] ));
 sg13g2_dfrbp_1 _22974_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net5962),
    .D(_01843_),
    .Q_N(_09474_),
    .Q(\TRNG.Padded_Out[215] ));
 sg13g2_dfrbp_1 _22975_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net5959),
    .D(_01844_),
    .Q_N(_09473_),
    .Q(\TRNG.Padded_Out[216] ));
 sg13g2_dfrbp_1 _22976_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net5944),
    .D(net2191),
    .Q_N(_09472_),
    .Q(\TRNG.Padded_Out[217] ));
 sg13g2_dfrbp_1 _22977_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net5944),
    .D(net1766),
    .Q_N(_09471_),
    .Q(\TRNG.Padded_Out[218] ));
 sg13g2_dfrbp_1 _22978_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net5940),
    .D(_01847_),
    .Q_N(_09470_),
    .Q(\TRNG.Padded_Out[219] ));
 sg13g2_dfrbp_1 _22979_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net5914),
    .D(net1459),
    .Q_N(_09469_),
    .Q(\TRNG.Padded_Out[220] ));
 sg13g2_dfrbp_1 _22980_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net5915),
    .D(net2008),
    .Q_N(_09468_),
    .Q(\TRNG.Padded_Out[221] ));
 sg13g2_dfrbp_1 _22981_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net5921),
    .D(_01850_),
    .Q_N(_09467_),
    .Q(\TRNG.Padded_Out[222] ));
 sg13g2_dfrbp_1 _22982_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net5921),
    .D(_01851_),
    .Q_N(_09466_),
    .Q(\TRNG.Padded_Out[223] ));
 sg13g2_dfrbp_1 _22983_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net5919),
    .D(net2093),
    .Q_N(_09465_),
    .Q(\TRNG.Padded_Out[224] ));
 sg13g2_dfrbp_1 _22984_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net5924),
    .D(net1740),
    .Q_N(_09464_),
    .Q(\TRNG.Padded_Out[225] ));
 sg13g2_dfrbp_1 _22985_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net5923),
    .D(net1727),
    .Q_N(_09463_),
    .Q(\TRNG.Padded_Out[226] ));
 sg13g2_dfrbp_1 _22986_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net5927),
    .D(net2181),
    .Q_N(_09462_),
    .Q(\TRNG.Padded_Out[227] ));
 sg13g2_dfrbp_1 _22987_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net5928),
    .D(_01856_),
    .Q_N(_09461_),
    .Q(\TRNG.Padded_Out[228] ));
 sg13g2_dfrbp_1 _22988_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net5928),
    .D(_01857_),
    .Q_N(_09460_),
    .Q(\TRNG.Padded_Out[229] ));
 sg13g2_dfrbp_1 _22989_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net5986),
    .D(net2029),
    .Q_N(_09459_),
    .Q(\TRNG.Padded_Out[230] ));
 sg13g2_dfrbp_1 _22990_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net6004),
    .D(_01859_),
    .Q_N(_09458_),
    .Q(\TRNG.Padded_Out[231] ));
 sg13g2_dfrbp_1 _22991_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net6003),
    .D(net1486),
    .Q_N(_09457_),
    .Q(\TRNG.Padded_Out[232] ));
 sg13g2_dfrbp_1 _22992_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net6002),
    .D(net1455),
    .Q_N(_09456_),
    .Q(\TRNG.Padded_Out[233] ));
 sg13g2_dfrbp_1 _22993_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net5996),
    .D(net1468),
    .Q_N(_09455_),
    .Q(\TRNG.Padded_Out[234] ));
 sg13g2_dfrbp_1 _22994_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net6044),
    .D(net1340),
    .Q_N(_09454_),
    .Q(\TRNG.Padded_Out[235] ));
 sg13g2_dfrbp_1 _22995_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net6042),
    .D(net1656),
    .Q_N(_09453_),
    .Q(\TRNG.Padded_Out[236] ));
 sg13g2_dfrbp_1 _22996_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net5994),
    .D(net1785),
    .Q_N(_09452_),
    .Q(\TRNG.Padded_Out[237] ));
 sg13g2_dfrbp_1 _22997_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net5966),
    .D(net2037),
    .Q_N(_09451_),
    .Q(\TRNG.Padded_Out[238] ));
 sg13g2_dfrbp_1 _22998_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net6019),
    .D(_01867_),
    .Q_N(_09450_),
    .Q(\TRNG.Padded_Out[239] ));
 sg13g2_dfrbp_1 _22999_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net6024),
    .D(net2022),
    .Q_N(_09449_),
    .Q(\TRNG.Padded_Out[240] ));
 sg13g2_dfrbp_1 _23000_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net6035),
    .D(net1841),
    .Q_N(_09448_),
    .Q(\TRNG.Padded_Out[241] ));
 sg13g2_dfrbp_1 _23001_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net6027),
    .D(_01870_),
    .Q_N(_09447_),
    .Q(\TRNG.Padded_Out[242] ));
 sg13g2_dfrbp_1 _23002_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net6031),
    .D(net1668),
    .Q_N(_09446_),
    .Q(\TRNG.Padded_Out[243] ));
 sg13g2_dfrbp_1 _23003_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net6009),
    .D(net2222),
    .Q_N(_09445_),
    .Q(\TRNG.Padded_Out[244] ));
 sg13g2_dfrbp_1 _23004_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net6008),
    .D(net1447),
    .Q_N(_09444_),
    .Q(\TRNG.Padded_Out[245] ));
 sg13g2_dfrbp_1 _23005_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net5953),
    .D(net1717),
    .Q_N(_09443_),
    .Q(\TRNG.Padded_Out[246] ));
 sg13g2_dfrbp_1 _23006_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net5952),
    .D(net1915),
    .Q_N(_09442_),
    .Q(\TRNG.Padded_Out[247] ));
 sg13g2_dfrbp_1 _23007_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net5938),
    .D(net1285),
    .Q_N(_09441_),
    .Q(\TRNG.Padded_Out[248] ));
 sg13g2_dfrbp_1 _23008_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net5937),
    .D(net1275),
    .Q_N(_09440_),
    .Q(\TRNG.Padded_Out[249] ));
 sg13g2_dfrbp_1 _23009_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net5945),
    .D(net1878),
    .Q_N(_09439_),
    .Q(\TRNG.Padded_Out[250] ));
 sg13g2_dfrbp_1 _23010_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net5941),
    .D(net1803),
    .Q_N(_09438_),
    .Q(\TRNG.Padded_Out[251] ));
 sg13g2_dfrbp_1 _23011_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net5941),
    .D(net1417),
    .Q_N(_09437_),
    .Q(\TRNG.Padded_Out[252] ));
 sg13g2_dfrbp_1 _23012_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net5946),
    .D(net1684),
    .Q_N(_09436_),
    .Q(\TRNG.Padded_Out[253] ));
 sg13g2_dfrbp_1 _23013_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net5946),
    .D(_01882_),
    .Q_N(_09435_),
    .Q(\TRNG.Padded_Out[254] ));
 sg13g2_dfrbp_1 _23014_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net5970),
    .D(net2001),
    .Q_N(_09434_),
    .Q(\TRNG.Padded_Out[255] ));
 sg13g2_dfrbp_1 _23015_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net5974),
    .D(net1303),
    .Q_N(_09433_),
    .Q(\TRNG.Padded_Out[256] ));
 sg13g2_dfrbp_1 _23016_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net5974),
    .D(_01885_),
    .Q_N(_09432_),
    .Q(\TRNG.Padded_Out[257] ));
 sg13g2_dfrbp_1 _23017_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net5923),
    .D(net1844),
    .Q_N(_09431_),
    .Q(\TRNG.Padded_Out[258] ));
 sg13g2_dfrbp_1 _23018_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net5980),
    .D(net1295),
    .Q_N(_09430_),
    .Q(\TRNG.Padded_Out[259] ));
 sg13g2_dfrbp_1 _23019_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net5981),
    .D(net1702),
    .Q_N(_09429_),
    .Q(\TRNG.Padded_Out[260] ));
 sg13g2_dfrbp_1 _23020_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net5982),
    .D(net1556),
    .Q_N(_09428_),
    .Q(\TRNG.Padded_Out[261] ));
 sg13g2_dfrbp_1 _23021_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net5999),
    .D(_01890_),
    .Q_N(_09427_),
    .Q(\TRNG.Padded_Out[262] ));
 sg13g2_dfrbp_1 _23022_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net6004),
    .D(net1279),
    .Q_N(_09426_),
    .Q(\TRNG.Padded_Out[263] ));
 sg13g2_dfrbp_1 _23023_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net6050),
    .D(net1453),
    .Q_N(_09425_),
    .Q(\TRNG.Padded_Out[264] ));
 sg13g2_dfrbp_1 _23024_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net6051),
    .D(net1250),
    .Q_N(_09424_),
    .Q(\TRNG.Padded_Out[265] ));
 sg13g2_dfrbp_1 _23025_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net6055),
    .D(net1970),
    .Q_N(_09423_),
    .Q(\TRNG.Padded_Out[266] ));
 sg13g2_dfrbp_1 _23026_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net6043),
    .D(net1811),
    .Q_N(_09422_),
    .Q(\TRNG.Padded_Out[267] ));
 sg13g2_dfrbp_1 _23027_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net5993),
    .D(net1572),
    .Q_N(_09421_),
    .Q(\TRNG.Padded_Out[268] ));
 sg13g2_dfrbp_1 _23028_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net5961),
    .D(net2156),
    .Q_N(_09420_),
    .Q(\TRNG.Padded_Out[269] ));
 sg13g2_dfrbp_1 _23029_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net5960),
    .D(net1531),
    .Q_N(_09419_),
    .Q(\TRNG.Padded_Out[270] ));
 sg13g2_dfrbp_1 _23030_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net6018),
    .D(net1860),
    .Q_N(_09418_),
    .Q(\TRNG.Padded_Out[271] ));
 sg13g2_dfrbp_1 _23031_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net6021),
    .D(net1619),
    .Q_N(_09417_),
    .Q(\TRNG.Padded_Out[272] ));
 sg13g2_dfrbp_1 _23032_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net6028),
    .D(net1615),
    .Q_N(_09416_),
    .Q(\TRNG.Padded_Out[273] ));
 sg13g2_dfrbp_1 _23033_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net6028),
    .D(net1706),
    .Q_N(_09415_),
    .Q(\TRNG.Padded_Out[274] ));
 sg13g2_dfrbp_1 _23034_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net6015),
    .D(net1264),
    .Q_N(_09414_),
    .Q(\TRNG.Padded_Out[275] ));
 sg13g2_dfrbp_1 _23035_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net6014),
    .D(net1370),
    .Q_N(_09413_),
    .Q(\TRNG.Padded_Out[276] ));
 sg13g2_dfrbp_1 _23036_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net5956),
    .D(net1384),
    .Q_N(_09412_),
    .Q(\TRNG.Padded_Out[277] ));
 sg13g2_dfrbp_1 _23037_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net5963),
    .D(net1378),
    .Q_N(_09411_),
    .Q(\TRNG.Padded_Out[278] ));
 sg13g2_dfrbp_1 _23038_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net5959),
    .D(net1632),
    .Q_N(_09410_),
    .Q(\TRNG.Padded_Out[279] ));
 sg13g2_dfrbp_1 _23039_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net5959),
    .D(net1392),
    .Q_N(_09409_),
    .Q(\TRNG.Padded_Out[280] ));
 sg13g2_dfrbp_1 _23040_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net5944),
    .D(_01909_),
    .Q_N(_09408_),
    .Q(\TRNG.Padded_Out[281] ));
 sg13g2_dfrbp_1 _23041_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net5944),
    .D(net1899),
    .Q_N(_09407_),
    .Q(\TRNG.Padded_Out[282] ));
 sg13g2_dfrbp_1 _23042_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net5941),
    .D(_01911_),
    .Q_N(_09406_),
    .Q(\TRNG.Padded_Out[283] ));
 sg13g2_dfrbp_1 _23043_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net5942),
    .D(net1738),
    .Q_N(_09405_),
    .Q(\TRNG.Padded_Out[284] ));
 sg13g2_dfrbp_1 _23044_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net5946),
    .D(net1345),
    .Q_N(_09404_),
    .Q(\TRNG.Padded_Out[285] ));
 sg13g2_dfrbp_1 _23045_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net5947),
    .D(net1907),
    .Q_N(_09403_),
    .Q(\TRNG.Padded_Out[286] ));
 sg13g2_dfrbp_1 _23046_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net5989),
    .D(net1499),
    .Q_N(_09402_),
    .Q(\TRNG.Padded_Out[287] ));
 sg13g2_dfrbp_1 _23047_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net5989),
    .D(net2146),
    .Q_N(_09401_),
    .Q(\TRNG.Padded_Out[288] ));
 sg13g2_dfrbp_1 _23048_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net5989),
    .D(_01917_),
    .Q_N(_09400_),
    .Q(\TRNG.Padded_Out[289] ));
 sg13g2_dfrbp_1 _23049_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net5971),
    .D(net1729),
    .Q_N(_09399_),
    .Q(\TRNG.Padded_Out[290] ));
 sg13g2_dfrbp_1 _23050_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net5980),
    .D(net1801),
    .Q_N(_09398_),
    .Q(\TRNG.Padded_Out[291] ));
 sg13g2_dfrbp_1 _23051_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net5981),
    .D(_01920_),
    .Q_N(_09397_),
    .Q(\TRNG.Padded_Out[292] ));
 sg13g2_dfrbp_1 _23052_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net5985),
    .D(_01921_),
    .Q_N(_09396_),
    .Q(\TRNG.Padded_Out[293] ));
 sg13g2_dfrbp_1 _23053_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net6000),
    .D(net1646),
    .Q_N(_09395_),
    .Q(\TRNG.Padded_Out[294] ));
 sg13g2_dfrbp_1 _23054_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net6000),
    .D(_01923_),
    .Q_N(_09394_),
    .Q(\TRNG.Padded_Out[295] ));
 sg13g2_dfrbp_1 _23055_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net6052),
    .D(_01924_),
    .Q_N(_09393_),
    .Q(\TRNG.Padded_Out[296] ));
 sg13g2_dfrbp_1 _23056_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net6057),
    .D(_01925_),
    .Q_N(_09392_),
    .Q(\TRNG.Padded_Out[297] ));
 sg13g2_dfrbp_1 _23057_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net6057),
    .D(net2127),
    .Q_N(_09391_),
    .Q(\TRNG.Padded_Out[298] ));
 sg13g2_dfrbp_1 _23058_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net6047),
    .D(net1692),
    .Q_N(_09390_),
    .Q(\TRNG.Padded_Out[299] ));
 sg13g2_dfrbp_1 _23059_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net6048),
    .D(net1779),
    .Q_N(_09389_),
    .Q(\TRNG.Padded_Out[300] ));
 sg13g2_dfrbp_1 _23060_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net6045),
    .D(net1436),
    .Q_N(_09388_),
    .Q(\TRNG.Padded_Out[301] ));
 sg13g2_dfrbp_1 _23061_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net6046),
    .D(net1856),
    .Q_N(_09387_),
    .Q(\TRNG.Padded_Out[302] ));
 sg13g2_dfrbp_1 _23062_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net6024),
    .D(_01931_),
    .Q_N(_09386_),
    .Q(\TRNG.Padded_Out[303] ));
 sg13g2_dfrbp_1 _23063_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net6037),
    .D(net1972),
    .Q_N(_09385_),
    .Q(\TRNG.Padded_Out[304] ));
 sg13g2_dfrbp_1 _23064_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net6033),
    .D(_01933_),
    .Q_N(_09384_),
    .Q(\TRNG.Padded_Out[305] ));
 sg13g2_dfrbp_1 _23065_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net6031),
    .D(_01934_),
    .Q_N(_09383_),
    .Q(\TRNG.Padded_Out[306] ));
 sg13g2_dfrbp_1 _23066_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net6031),
    .D(net2278),
    .Q_N(_09382_),
    .Q(\TRNG.Padded_Out[307] ));
 sg13g2_dfrbp_1 _23067_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net6013),
    .D(net1439),
    .Q_N(_09381_),
    .Q(\TRNG.Padded_Out[308] ));
 sg13g2_dfrbp_1 _23068_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net6011),
    .D(net1266),
    .Q_N(_09380_),
    .Q(\TRNG.Padded_Out[309] ));
 sg13g2_dfrbp_1 _23069_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net5955),
    .D(net2043),
    .Q_N(_09379_),
    .Q(\TRNG.Padded_Out[310] ));
 sg13g2_dfrbp_1 _23070_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net5959),
    .D(net1967),
    .Q_N(_09378_),
    .Q(\TRNG.Padded_Out[311] ));
 sg13g2_dfrbp_1 _23071_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net5951),
    .D(_01940_),
    .Q_N(_09377_),
    .Q(\TRNG.Padded_Out[312] ));
 sg13g2_dfrbp_1 _23072_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net5937),
    .D(net1380),
    .Q_N(_09376_),
    .Q(\TRNG.Padded_Out[313] ));
 sg13g2_dfrbp_1 _23073_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net5907),
    .D(_01942_),
    .Q_N(_09375_),
    .Q(\TRNG.Padded_Out[314] ));
 sg13g2_dfrbp_1 _23074_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net5932),
    .D(net1297),
    .Q_N(_09374_),
    .Q(\TRNG.Padded_Out[315] ));
 sg13g2_dfrbp_1 _23075_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net5940),
    .D(net1529),
    .Q_N(_09373_),
    .Q(\TRNG.Padded_Out[316] ));
 sg13g2_dfrbp_1 _23076_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net5947),
    .D(net1642),
    .Q_N(_09372_),
    .Q(\TRNG.Padded_Out[317] ));
 sg13g2_dfrbp_1 _23077_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net5960),
    .D(_01946_),
    .Q_N(_09371_),
    .Q(\TRNG.Padded_Out[318] ));
 sg13g2_dfrbp_1 _23078_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net5960),
    .D(_01947_),
    .Q_N(_09370_),
    .Q(\TRNG.Padded_Out[319] ));
 sg13g2_dfrbp_1 _23079_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net5989),
    .D(net1848),
    .Q_N(_09369_),
    .Q(\TRNG.Padded_Out[320] ));
 sg13g2_dfrbp_1 _23080_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net5977),
    .D(net1361),
    .Q_N(_09368_),
    .Q(\TRNG.Padded_Out[321] ));
 sg13g2_dfrbp_1 _23081_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net5972),
    .D(net1926),
    .Q_N(_09367_),
    .Q(\TRNG.Padded_Out[322] ));
 sg13g2_dfrbp_1 _23082_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net5979),
    .D(net1322),
    .Q_N(_09366_),
    .Q(\TRNG.Padded_Out[323] ));
 sg13g2_dfrbp_1 _23083_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net5979),
    .D(net1586),
    .Q_N(_09365_),
    .Q(\TRNG.Padded_Out[324] ));
 sg13g2_dfrbp_1 _23084_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net5983),
    .D(_01953_),
    .Q_N(_09364_),
    .Q(\TRNG.Padded_Out[325] ));
 sg13g2_dfrbp_1 _23085_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net5984),
    .D(net1799),
    .Q_N(_09363_),
    .Q(\TRNG.Padded_Out[326] ));
 sg13g2_dfrbp_1 _23086_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net5991),
    .D(net1316),
    .Q_N(_09362_),
    .Q(\TRNG.Padded_Out[327] ));
 sg13g2_dfrbp_1 _23087_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net5991),
    .D(net1353),
    .Q_N(_09361_),
    .Q(\TRNG.Padded_Out[328] ));
 sg13g2_dfrbp_1 _23088_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net5991),
    .D(_01957_),
    .Q_N(_09360_),
    .Q(\TRNG.Padded_Out[329] ));
 sg13g2_dfrbp_1 _23089_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net5995),
    .D(_01958_),
    .Q_N(_09359_),
    .Q(\TRNG.Padded_Out[330] ));
 sg13g2_dfrbp_1 _23090_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net5993),
    .D(net1482),
    .Q_N(_09358_),
    .Q(\TRNG.Padded_Out[331] ));
 sg13g2_dfrbp_1 _23091_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net5993),
    .D(net1330),
    .Q_N(_09357_),
    .Q(\TRNG.Padded_Out[332] ));
 sg13g2_dfrbp_1 _23092_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net5993),
    .D(net1244),
    .Q_N(_09356_),
    .Q(\TRNG.Padded_Out[333] ));
 sg13g2_dfrbp_1 _23093_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net6019),
    .D(net1807),
    .Q_N(_09355_),
    .Q(\TRNG.Padded_Out[334] ));
 sg13g2_dfrbp_1 _23094_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net5964),
    .D(net1515),
    .Q_N(_09354_),
    .Q(\TRNG.Padded_Out[335] ));
 sg13g2_dfrbp_1 _23095_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net6020),
    .D(net1775),
    .Q_N(_09353_),
    .Q(\TRNG.Padded_Out[336] ));
 sg13g2_dfrbp_1 _23096_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net6013),
    .D(net1283),
    .Q_N(_09352_),
    .Q(\TRNG.Padded_Out[337] ));
 sg13g2_dfrbp_1 _23097_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net6026),
    .D(net1771),
    .Q_N(_09351_),
    .Q(\TRNG.Padded_Out[338] ));
 sg13g2_dfrbp_1 _23098_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net6013),
    .D(_01967_),
    .Q_N(_09350_),
    .Q(\TRNG.Padded_Out[339] ));
 sg13g2_dfrbp_1 _23099_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net6012),
    .D(net1594),
    .Q_N(_09349_),
    .Q(\TRNG.Padded_Out[340] ));
 sg13g2_dfrbp_1 _23100_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net6008),
    .D(net2069),
    .Q_N(_09348_),
    .Q(\TRNG.Padded_Out[341] ));
 sg13g2_dfrbp_1 _23101_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net5953),
    .D(net2321),
    .Q_N(_09347_),
    .Q(\TRNG.Padded_Out[342] ));
 sg13g2_dfrbp_1 _23102_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net5949),
    .D(net2046),
    .Q_N(_09346_),
    .Q(\TRNG.Padded_Out[343] ));
 sg13g2_dfrbp_1 _23103_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net5936),
    .D(net1746),
    .Q_N(_09345_),
    .Q(\TRNG.Padded_Out[344] ));
 sg13g2_dfrbp_1 _23104_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net5934),
    .D(_01973_),
    .Q_N(_09344_),
    .Q(\TRNG.Padded_Out[345] ));
 sg13g2_dfrbp_1 _23105_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net5909),
    .D(net1783),
    .Q_N(_09343_),
    .Q(\TRNG.Padded_Out[346] ));
 sg13g2_dfrbp_1 _23106_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net5907),
    .D(net2247),
    .Q_N(_09342_),
    .Q(\TRNG.Padded_Out[347] ));
 sg13g2_dfrbp_1 _23107_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net5913),
    .D(net1343),
    .Q_N(_09341_),
    .Q(\TRNG.Padded_Out[348] ));
 sg13g2_dfrbp_1 _23108_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net5942),
    .D(net1474),
    .Q_N(_09340_),
    .Q(\TRNG.Padded_Out[349] ));
 sg13g2_dfrbp_1 _23109_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net5943),
    .D(_01978_),
    .Q_N(_09339_),
    .Q(\TRNG.Padded_Out[350] ));
 sg13g2_dfrbp_1 _23110_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net5975),
    .D(net1351),
    .Q_N(_09338_),
    .Q(\TRNG.Padded_Out[351] ));
 sg13g2_dfrbp_1 _23111_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net5970),
    .D(net1910),
    .Q_N(_09337_),
    .Q(\TRNG.Padded_Out[352] ));
 sg13g2_dfrbp_1 _23112_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net5923),
    .D(net1924),
    .Q_N(_09336_),
    .Q(\TRNG.Padded_Out[353] ));
 sg13g2_dfrbp_1 _23113_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net5923),
    .D(net1638),
    .Q_N(_09335_),
    .Q(\TRNG.Padded_Out[354] ));
 sg13g2_dfrbp_1 _23114_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net5980),
    .D(net1559),
    .Q_N(_09334_),
    .Q(\TRNG.Padded_Out[355] ));
 sg13g2_dfrbp_1 _23115_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net5981),
    .D(_01984_),
    .Q_N(_09333_),
    .Q(\TRNG.Padded_Out[356] ));
 sg13g2_dfrbp_1 _23116_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net5985),
    .D(net2142),
    .Q_N(_09332_),
    .Q(\TRNG.Padded_Out[357] ));
 sg13g2_dfrbp_1 _23117_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net6000),
    .D(net2176),
    .Q_N(_09331_),
    .Q(\TRNG.Padded_Out[358] ));
 sg13g2_dfrbp_1 _23118_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net6005),
    .D(_01987_),
    .Q_N(_09330_),
    .Q(\TRNG.Padded_Out[359] ));
 sg13g2_dfrbp_1 _23119_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net6052),
    .D(_01988_),
    .Q_N(_09329_),
    .Q(\TRNG.Padded_Out[360] ));
 sg13g2_dfrbp_1 _23120_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net6053),
    .D(net2198),
    .Q_N(_09328_),
    .Q(\TRNG.Padded_Out[361] ));
 sg13g2_dfrbp_1 _23121_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net6044),
    .D(net1477),
    .Q_N(_09327_),
    .Q(\TRNG.Padded_Out[362] ));
 sg13g2_dfrbp_1 _23122_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net6043),
    .D(net1464),
    .Q_N(_09326_),
    .Q(\TRNG.Padded_Out[363] ));
 sg13g2_dfrbp_1 _23123_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net6047),
    .D(net1318),
    .Q_N(_09325_),
    .Q(\TRNG.Padded_Out[364] ));
 sg13g2_dfrbp_1 _23124_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net6041),
    .D(net1790),
    .Q_N(_09324_),
    .Q(\TRNG.Padded_Out[365] ));
 sg13g2_dfrbp_1 _23125_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net5966),
    .D(net1355),
    .Q_N(_09323_),
    .Q(\TRNG.Padded_Out[366] ));
 sg13g2_dfrbp_1 _23126_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net5965),
    .D(net1677),
    .Q_N(_09322_),
    .Q(\TRNG.Padded_Out[367] ));
 sg13g2_dfrbp_1 _23127_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net6020),
    .D(_01996_),
    .Q_N(_09321_),
    .Q(\TRNG.Padded_Out[368] ));
 sg13g2_dfrbp_1 _23128_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net6022),
    .D(net2152),
    .Q_N(_09320_),
    .Q(\TRNG.Padded_Out[369] ));
 sg13g2_dfrbp_1 _23129_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net6026),
    .D(net1421),
    .Q_N(_09319_),
    .Q(\TRNG.Padded_Out[370] ));
 sg13g2_dfrbp_1 _23130_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net6031),
    .D(net1544),
    .Q_N(_09318_),
    .Q(\TRNG.Padded_Out[371] ));
 sg13g2_dfrbp_1 _23131_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net6010),
    .D(net1497),
    .Q_N(_09317_),
    .Q(\TRNG.Padded_Out[372] ));
 sg13g2_dfrbp_1 _23132_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net5954),
    .D(net1326),
    .Q_N(_09316_),
    .Q(\TRNG.Padded_Out[373] ));
 sg13g2_dfrbp_1 _23133_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net5955),
    .D(net1777),
    .Q_N(_09315_),
    .Q(\TRNG.Padded_Out[374] ));
 sg13g2_dfrbp_1 _23134_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net5952),
    .D(net1636),
    .Q_N(_09314_),
    .Q(\TRNG.Padded_Out[375] ));
 sg13g2_dfrbp_1 _23135_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net5951),
    .D(net2196),
    .Q_N(_09313_),
    .Q(\TRNG.Padded_Out[376] ));
 sg13g2_dfrbp_1 _23136_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net5932),
    .D(_02005_),
    .Q_N(_09312_),
    .Q(\TRNG.Padded_Out[377] ));
 sg13g2_dfrbp_1 _23137_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net5907),
    .D(net1287),
    .Q_N(_09311_),
    .Q(\TRNG.Padded_Out[378] ));
 sg13g2_dfrbp_1 _23138_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net5907),
    .D(net1347),
    .Q_N(_09310_),
    .Q(\TRNG.Padded_Out[379] ));
 sg13g2_dfrbp_1 _23139_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net5914),
    .D(net1535),
    .Q_N(_09309_),
    .Q(\TRNG.Padded_Out[380] ));
 sg13g2_dfrbp_1 _23140_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net5945),
    .D(net2011),
    .Q_N(_09308_),
    .Q(\TRNG.Padded_Out[381] ));
 sg13g2_dfrbp_1 _23141_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net5947),
    .D(net1324),
    .Q_N(_09307_),
    .Q(\TRNG.Padded_Out[382] ));
 sg13g2_dfrbp_1 _23142_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net5960),
    .D(_02011_),
    .Q_N(_09306_),
    .Q(\TRNG.Padded_Out[383] ));
 sg13g2_dfrbp_1 _23143_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net5989),
    .D(net1312),
    .Q_N(_09305_),
    .Q(\TRNG.Padded_Out[384] ));
 sg13g2_dfrbp_1 _23144_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net5969),
    .D(net1988),
    .Q_N(_09304_),
    .Q(\TRNG.Padded_Out[385] ));
 sg13g2_dfrbp_1 _23145_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net5971),
    .D(net1141),
    .Q_N(_09303_),
    .Q(\TRNG.Padded_Out[386] ));
 sg13g2_dfrbp_1 _23146_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net5972),
    .D(net1167),
    .Q_N(_09302_),
    .Q(\TRNG.Padded_Out[387] ));
 sg13g2_dfrbp_1 _23147_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net5980),
    .D(_02016_),
    .Q_N(_09301_),
    .Q(\TRNG.Padded_Out[388] ));
 sg13g2_dfrbp_1 _23148_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net5985),
    .D(_02017_),
    .Q_N(_09300_),
    .Q(\TRNG.Padded_Out[389] ));
 sg13g2_dfrbp_1 _23149_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net5999),
    .D(net1289),
    .Q_N(_09299_),
    .Q(\TRNG.Padded_Out[390] ));
 sg13g2_dfrbp_1 _23150_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net5998),
    .D(_02019_),
    .Q_N(_09298_),
    .Q(\TRNG.Padded_Out[391] ));
 sg13g2_dfrbp_1 _23151_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net6052),
    .D(net1338),
    .Q_N(_09297_),
    .Q(\TRNG.Padded_Out[392] ));
 sg13g2_dfrbp_1 _23152_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net6053),
    .D(net1882),
    .Q_N(_09296_),
    .Q(\TRNG.Padded_Out[393] ));
 sg13g2_dfrbp_1 _23153_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net6057),
    .D(net1582),
    .Q_N(_09295_),
    .Q(\TRNG.Padded_Out[394] ));
 sg13g2_dfrbp_1 _23154_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net6055),
    .D(net1305),
    .Q_N(_09294_),
    .Q(\TRNG.Padded_Out[395] ));
 sg13g2_dfrbp_1 _23155_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net5994),
    .D(net1334),
    .Q_N(_09293_),
    .Q(\TRNG.Padded_Out[396] ));
 sg13g2_dfrbp_1 _23156_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net5994),
    .D(_02025_),
    .Q_N(_09292_),
    .Q(\TRNG.Padded_Out[397] ));
 sg13g2_dfrbp_1 _23157_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net6041),
    .D(_02026_),
    .Q_N(_09291_),
    .Q(\TRNG.Padded_Out[398] ));
 sg13g2_dfrbp_1 _23158_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net6019),
    .D(net1628),
    .Q_N(_09290_),
    .Q(\TRNG.Padded_Out[399] ));
 sg13g2_dfrbp_1 _23159_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net6023),
    .D(net1413),
    .Q_N(_09289_),
    .Q(\TRNG.Padded_Out[400] ));
 sg13g2_dfrbp_1 _23160_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net6026),
    .D(net1301),
    .Q_N(_09288_),
    .Q(\TRNG.Padded_Out[401] ));
 sg13g2_dfrbp_1 _23161_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net6026),
    .D(net1606),
    .Q_N(_09287_),
    .Q(\TRNG.Padded_Out[402] ));
 sg13g2_dfrbp_1 _23162_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net6026),
    .D(net2304),
    .Q_N(_09286_),
    .Q(\TRNG.Padded_Out[403] ));
 sg13g2_dfrbp_1 _23163_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net6012),
    .D(net1359),
    .Q_N(_09285_),
    .Q(\TRNG.Padded_Out[404] ));
 sg13g2_dfrbp_1 _23164_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net5954),
    .D(net1919),
    .Q_N(_09284_),
    .Q(\TRNG.Padded_Out[405] ));
 sg13g2_dfrbp_1 _23165_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net5953),
    .D(net2019),
    .Q_N(_09283_),
    .Q(\TRNG.Padded_Out[406] ));
 sg13g2_dfrbp_1 _23166_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net5949),
    .D(net1903),
    .Q_N(_09282_),
    .Q(\TRNG.Padded_Out[407] ));
 sg13g2_dfrbp_1 _23167_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net5936),
    .D(net2172),
    .Q_N(_09281_),
    .Q(\TRNG.Padded_Out[408] ));
 sg13g2_dfrbp_1 _23168_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net5933),
    .D(net1640),
    .Q_N(_09280_),
    .Q(\TRNG.Padded_Out[409] ));
 sg13g2_dfrbp_1 _23169_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net5908),
    .D(_02038_),
    .Q_N(_09279_),
    .Q(\TRNG.Padded_Out[410] ));
 sg13g2_dfrbp_1 _23170_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net5940),
    .D(net1310),
    .Q_N(_09278_),
    .Q(\TRNG.Padded_Out[411] ));
 sg13g2_dfrbp_1 _23171_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net5940),
    .D(net1277),
    .Q_N(_09277_),
    .Q(\TRNG.Padded_Out[412] ));
 sg13g2_dfrbp_1 _23172_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net5943),
    .D(_02041_),
    .Q_N(_09276_),
    .Q(\TRNG.Padded_Out[413] ));
 sg13g2_dfrbp_1 _23173_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net5969),
    .D(_02042_),
    .Q_N(_09275_),
    .Q(\TRNG.Padded_Out[414] ));
 sg13g2_dfrbp_1 _23174_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net5974),
    .D(net1754),
    .Q_N(_09274_),
    .Q(\TRNG.Padded_Out[415] ));
 sg13g2_dfrbp_1 _23175_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net5974),
    .D(net1503),
    .Q_N(_09273_),
    .Q(\TRNG.Padded_Out[416] ));
 sg13g2_dfrbp_1 _23176_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net5976),
    .D(net1252),
    .Q_N(_09272_),
    .Q(\TRNG.Padded_Out[417] ));
 sg13g2_dfrbp_1 _23177_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net5977),
    .D(net1666),
    .Q_N(_09271_),
    .Q(\TRNG.Padded_Out[418] ));
 sg13g2_dfrbp_1 _23178_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net5977),
    .D(net1336),
    .Q_N(_09270_),
    .Q(\TRNG.Padded_Out[419] ));
 sg13g2_dfrbp_1 _23179_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net5979),
    .D(_02048_),
    .Q_N(_09269_),
    .Q(\TRNG.Padded_Out[420] ));
 sg13g2_dfrbp_1 _23180_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net5986),
    .D(net1688),
    .Q_N(_09268_),
    .Q(\TRNG.Padded_Out[421] ));
 sg13g2_dfrbp_1 _23181_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net6000),
    .D(net1501),
    .Q_N(_09267_),
    .Q(\TRNG.Padded_Out[422] ));
 sg13g2_dfrbp_1 _23182_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net6004),
    .D(net1930),
    .Q_N(_09266_),
    .Q(\TRNG.Padded_Out[423] ));
 sg13g2_dfrbp_1 _23183_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net6052),
    .D(_02052_),
    .Q_N(_09265_),
    .Q(\TRNG.Padded_Out[424] ));
 sg13g2_dfrbp_1 _23184_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net6051),
    .D(net1869),
    .Q_N(_09264_),
    .Q(\TRNG.Padded_Out[425] ));
 sg13g2_dfrbp_1 _23185_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net6055),
    .D(net1552),
    .Q_N(_09263_),
    .Q(\TRNG.Padded_Out[426] ));
 sg13g2_dfrbp_1 _23186_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net6047),
    .D(net1731),
    .Q_N(_09262_),
    .Q(\TRNG.Padded_Out[427] ));
 sg13g2_dfrbp_1 _23187_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net6042),
    .D(net1649),
    .Q_N(_09261_),
    .Q(\TRNG.Padded_Out[428] ));
 sg13g2_dfrbp_1 _23188_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net6041),
    .D(net1825),
    .Q_N(_09260_),
    .Q(\TRNG.Padded_Out[429] ));
 sg13g2_dfrbp_1 _23189_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net6020),
    .D(net1993),
    .Q_N(_09259_),
    .Q(\TRNG.Padded_Out[430] ));
 sg13g2_dfrbp_1 _23190_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net6019),
    .D(net1525),
    .Q_N(_09258_),
    .Q(\TRNG.Padded_Out[431] ));
 sg13g2_dfrbp_1 _23191_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net6021),
    .D(net1548),
    .Q_N(_09257_),
    .Q(\TRNG.Padded_Out[432] ));
 sg13g2_dfrbp_1 _23192_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net6029),
    .D(net1443),
    .Q_N(_09256_),
    .Q(\TRNG.Padded_Out[433] ));
 sg13g2_dfrbp_1 _23193_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net6031),
    .D(_02062_),
    .Q_N(_09255_),
    .Q(\TRNG.Padded_Out[434] ));
 sg13g2_dfrbp_1 _23194_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net6032),
    .D(net2363),
    .Q_N(_09254_),
    .Q(\TRNG.Padded_Out[435] ));
 sg13g2_dfrbp_1 _23195_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net6012),
    .D(net1748),
    .Q_N(_09253_),
    .Q(\TRNG.Padded_Out[436] ));
 sg13g2_dfrbp_1 _23196_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net6008),
    .D(net1490),
    .Q_N(_09252_),
    .Q(\TRNG.Padded_Out[437] ));
 sg13g2_dfrbp_1 _23197_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net5953),
    .D(net1815),
    .Q_N(_09251_),
    .Q(\TRNG.Padded_Out[438] ));
 sg13g2_dfrbp_1 _23198_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net5950),
    .D(net1386),
    .Q_N(_09250_),
    .Q(\TRNG.Padded_Out[439] ));
 sg13g2_dfrbp_1 _23199_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net5950),
    .D(_02068_),
    .Q_N(_09249_),
    .Q(\TRNG.Padded_Out[440] ));
 sg13g2_dfrbp_1 _23200_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net5935),
    .D(_02069_),
    .Q_N(_09248_),
    .Q(\TRNG.Padded_Out[441] ));
 sg13g2_dfrbp_1 _23201_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net5933),
    .D(net1617),
    .Q_N(_09247_),
    .Q(\TRNG.Padded_Out[442] ));
 sg13g2_dfrbp_1 _23202_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net5913),
    .D(net1427),
    .Q_N(_09246_),
    .Q(\TRNG.Padded_Out[443] ));
 sg13g2_dfrbp_1 _23203_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net5914),
    .D(net1523),
    .Q_N(_09245_),
    .Q(\TRNG.Padded_Out[444] ));
 sg13g2_dfrbp_1 _23204_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net5942),
    .D(net1592),
    .Q_N(_09244_),
    .Q(\TRNG.Padded_Out[445] ));
 sg13g2_dfrbp_1 _23205_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net5943),
    .D(_02074_),
    .Q_N(_09243_),
    .Q(\TRNG.Padded_Out[446] ));
 sg13g2_dfrbp_1 _23206_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net5975),
    .D(net1590),
    .Q_N(_09242_),
    .Q(\TRNG.Padded_Out[447] ));
 sg13g2_dfrbp_1 _23207_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net5975),
    .D(net2061),
    .Q_N(_09241_),
    .Q(\TRNG.Padded_Out[448] ));
 sg13g2_dfrbp_1 _23208_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net5976),
    .D(net1488),
    .Q_N(_09240_),
    .Q(\TRNG.Padded_Out[449] ));
 sg13g2_dfrbp_1 _23209_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net5976),
    .D(net2098),
    .Q_N(_09239_),
    .Q(\TRNG.Padded_Out[450] ));
 sg13g2_dfrbp_1 _23210_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net5978),
    .D(net1505),
    .Q_N(_09238_),
    .Q(\TRNG.Padded_Out[451] ));
 sg13g2_dfrbp_1 _23211_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net5983),
    .D(_02080_),
    .Q_N(_09237_),
    .Q(\TRNG.Padded_Out[452] ));
 sg13g2_dfrbp_1 _23212_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net5984),
    .D(_02081_),
    .Q_N(_09236_),
    .Q(\TRNG.Padded_Out[453] ));
 sg13g2_dfrbp_1 _23213_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net5999),
    .D(_02082_),
    .Q_N(_09235_),
    .Q(\TRNG.Padded_Out[454] ));
 sg13g2_dfrbp_1 _23214_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net5998),
    .D(_02083_),
    .Q_N(_09234_),
    .Q(\TRNG.Padded_Out[455] ));
 sg13g2_dfrbp_1 _23215_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net6002),
    .D(net1596),
    .Q_N(_09233_),
    .Q(\TRNG.Padded_Out[456] ));
 sg13g2_dfrbp_1 _23216_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net6051),
    .D(net1626),
    .Q_N(_09232_),
    .Q(\TRNG.Padded_Out[457] ));
 sg13g2_dfrbp_1 _23217_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net5995),
    .D(_02086_),
    .Q_N(_09231_),
    .Q(\TRNG.Padded_Out[458] ));
 sg13g2_dfrbp_1 _23218_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net5995),
    .D(net1457),
    .Q_N(_09230_),
    .Q(\TRNG.Padded_Out[459] ));
 sg13g2_dfrbp_1 _23219_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net5993),
    .D(_02088_),
    .Q_N(_09229_),
    .Q(\TRNG.Padded_Out[460] ));
 sg13g2_dfrbp_1 _23220_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net5990),
    .D(net1715),
    .Q_N(_09228_),
    .Q(\TRNG.Padded_Out[461] ));
 sg13g2_dfrbp_1 _23221_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net5965),
    .D(_02090_),
    .Q_N(_09227_),
    .Q(\TRNG.Padded_Out[462] ));
 sg13g2_dfrbp_1 _23222_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net6023),
    .D(net1568),
    .Q_N(_09226_),
    .Q(\TRNG.Padded_Out[463] ));
 sg13g2_dfrbp_1 _23223_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net6021),
    .D(net1451),
    .Q_N(_09225_),
    .Q(\TRNG.Padded_Out[464] ));
 sg13g2_dfrbp_1 _23224_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net6028),
    .D(_02093_),
    .Q_N(_09224_),
    .Q(\TRNG.Padded_Out[465] ));
 sg13g2_dfrbp_1 _23225_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net6029),
    .D(net1613),
    .Q_N(_09223_),
    .Q(\TRNG.Padded_Out[466] ));
 sg13g2_dfrbp_1 _23226_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net6031),
    .D(net2224),
    .Q_N(_09222_),
    .Q(\TRNG.Padded_Out[467] ));
 sg13g2_dfrbp_1 _23227_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net6012),
    .D(net2251),
    .Q_N(_09221_),
    .Q(\TRNG.Padded_Out[468] ));
 sg13g2_dfrbp_1 _23228_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net5954),
    .D(net2310),
    .Q_N(_09220_),
    .Q(\TRNG.Padded_Out[469] ));
 sg13g2_dfrbp_1 _23229_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net5953),
    .D(_02098_),
    .Q_N(_09219_),
    .Q(\TRNG.Padded_Out[470] ));
 sg13g2_dfrbp_1 _23230_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net5952),
    .D(net1813),
    .Q_N(_09218_),
    .Q(\TRNG.Padded_Out[471] ));
 sg13g2_dfrbp_1 _23231_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net5935),
    .D(net2160),
    .Q_N(_09217_),
    .Q(\TRNG.Padded_Out[472] ));
 sg13g2_dfrbp_1 _23232_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net5934),
    .D(net1696),
    .Q_N(_09216_),
    .Q(\TRNG.Padded_Out[473] ));
 sg13g2_dfrbp_1 _23233_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net5909),
    .D(_02102_),
    .Q_N(_09215_),
    .Q(\TRNG.Padded_Out[474] ));
 sg13g2_dfrbp_1 _23234_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net5932),
    .D(net2148),
    .Q_N(_09214_),
    .Q(\TRNG.Padded_Out[475] ));
 sg13g2_dfrbp_1 _23235_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net5940),
    .D(net1445),
    .Q_N(_09213_),
    .Q(\TRNG.Padded_Out[476] ));
 sg13g2_dfrbp_1 _23236_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net5942),
    .D(net1889),
    .Q_N(_09212_),
    .Q(\TRNG.Padded_Out[477] ));
 sg13g2_dfrbp_1 _23237_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net5946),
    .D(_02106_),
    .Q_N(_09211_),
    .Q(\TRNG.Padded_Out[478] ));
 sg13g2_dfrbp_1 _23238_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net5960),
    .D(net1598),
    .Q_N(_09210_),
    .Q(\TRNG.Padded_Out[479] ));
 sg13g2_dfrbp_1 _23239_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net6039),
    .D(_02108_),
    .Q_N(_09209_),
    .Q(\TRNG.Padded_Out[480] ));
 sg13g2_dfrbp_1 _23240_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net6038),
    .D(net2355),
    .Q_N(_09208_),
    .Q(\TRNG.Padded_Out[481] ));
 sg13g2_dfrbp_1 _23241_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net6062),
    .D(_02110_),
    .Q_N(_09207_),
    .Q(\TRNG.Padded_Out[482] ));
 sg13g2_dfrbp_1 _23242_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net6063),
    .D(net1981),
    .Q_N(_09206_),
    .Q(\TRNG.Padded_Out[483] ));
 sg13g2_dfrbp_1 _23243_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net6061),
    .D(_02112_),
    .Q_N(_09205_),
    .Q(\TRNG.Padded_Out[484] ));
 sg13g2_dfrbp_1 _23244_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net6064),
    .D(_02113_),
    .Q_N(_09204_),
    .Q(\TRNG.Padded_Out[485] ));
 sg13g2_dfrbp_1 _23245_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net6064),
    .D(net1509),
    .Q_N(_09203_),
    .Q(\TRNG.Padded_Out[486] ));
 sg13g2_dfrbp_1 _23246_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net6064),
    .D(net1273),
    .Q_N(_09202_),
    .Q(\TRNG.Padded_Out[487] ));
 sg13g2_dfrbp_1 _23247_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net6055),
    .D(net1664),
    .Q_N(_09201_),
    .Q(\TRNG.Padded_Out[488] ));
 sg13g2_dfrbp_1 _23248_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net6060),
    .D(_02117_),
    .Q_N(_09200_),
    .Q(\TRNG.Padded_Out[489] ));
 sg13g2_dfrbp_1 _23249_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net6060),
    .D(net2481),
    .Q_N(_09199_),
    .Q(\TRNG.Padded_Out[490] ));
 sg13g2_dfrbp_1 _23250_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net6060),
    .D(_02119_),
    .Q_N(_09198_),
    .Q(\TRNG.Padded_Out[491] ));
 sg13g2_dfrbp_1 _23251_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net6060),
    .D(_02120_),
    .Q_N(_09197_),
    .Q(\TRNG.Padded_Out[492] ));
 sg13g2_dfrbp_1 _23252_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net6039),
    .D(_02121_),
    .Q_N(_09196_),
    .Q(\TRNG.Padded_Out[493] ));
 sg13g2_dfrbp_1 _23253_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net6038),
    .D(_02122_),
    .Q_N(_09195_),
    .Q(\TRNG.Padded_Out[494] ));
 sg13g2_dfrbp_1 _23254_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net6037),
    .D(_02123_),
    .Q_N(_09194_),
    .Q(\TRNG.Padded_Out[495] ));
 sg13g2_dfrbp_1 _23255_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net6038),
    .D(_02124_),
    .Q_N(_09193_),
    .Q(\TRNG.Padded_Out[496] ));
 sg13g2_dfrbp_1 _23256_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net6036),
    .D(net2734),
    .Q_N(_09192_),
    .Q(\TRNG.Padded_Out[497] ));
 sg13g2_dfrbp_1 _23257_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net6038),
    .D(_02126_),
    .Q_N(_09191_),
    .Q(\TRNG.Padded_Out[498] ));
 sg13g2_dfrbp_1 _23258_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net6034),
    .D(_02127_),
    .Q_N(_09190_),
    .Q(\TRNG.Padded_Out[499] ));
 sg13g2_dfrbp_1 _23259_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net6032),
    .D(_02128_),
    .Q_N(_09189_),
    .Q(\TRNG.Padded_Out[500] ));
 sg13g2_dfrbp_1 _23260_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net6033),
    .D(_02129_),
    .Q_N(_09188_),
    .Q(\TRNG.Padded_Out[501] ));
 sg13g2_dfrbp_1 _23261_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net6033),
    .D(_02130_),
    .Q_N(_09187_),
    .Q(\TRNG.Padded_Out[502] ));
 sg13g2_dfrbp_1 _23262_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net6033),
    .D(_02131_),
    .Q_N(_09186_),
    .Q(\TRNG.Padded_Out[503] ));
 sg13g2_dfrbp_1 _23263_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net6038),
    .D(net2576),
    .Q_N(_09185_),
    .Q(\TRNG.Padded_Out[504] ));
 sg13g2_dfrbp_1 _23264_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net6039),
    .D(net2379),
    .Q_N(_09184_),
    .Q(\TRNG.Padded_Out[505] ));
 sg13g2_dfrbp_1 _23265_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net6061),
    .D(_02134_),
    .Q_N(_09183_),
    .Q(\TRNG.Padded_Out[506] ));
 sg13g2_dfrbp_1 _23266_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net6061),
    .D(net1357),
    .Q_N(_09182_),
    .Q(\TRNG.Padded_Out[507] ));
 sg13g2_dfrbp_1 _23267_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net6062),
    .D(_02136_),
    .Q_N(_09181_),
    .Q(\TRNG.Padded_Out[508] ));
 sg13g2_dfrbp_1 _23268_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net6062),
    .D(_02137_),
    .Q_N(_09180_),
    .Q(\TRNG.Padded_Out[509] ));
 sg13g2_dfrbp_1 _23269_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net6064),
    .D(net1609),
    .Q_N(_09179_),
    .Q(\TRNG.Padded_Out[510] ));
 sg13g2_dfrbp_1 _23270_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net6064),
    .D(net2502),
    .Q_N(_11078_),
    .Q(\TRNG.Padded_Out[511] ));
 sg13g2_dfrbp_1 _23271_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net5906),
    .D(_02145_),
    .Q_N(_11079_),
    .Q(\TRNG.raw_bit_counter[0] ));
 sg13g2_dfrbp_1 _23272_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net5906),
    .D(net3402),
    .Q_N(_11080_),
    .Q(\TRNG.raw_bit_counter[1] ));
 sg13g2_dfrbp_1 _23273_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net5906),
    .D(net3315),
    .Q_N(_09178_),
    .Q(\TRNG.raw_bit_counter[2] ));
 sg13g2_dfrbp_1 _23274_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net5899),
    .D(net3545),
    .Q_N(_09177_),
    .Q(\TRNG.chunk_index[0] ));
 sg13g2_dfrbp_1 _23275_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net5899),
    .D(_02141_),
    .Q_N(_09176_),
    .Q(\TRNG.chunk_index[1] ));
 sg13g2_dfrbp_1 _23276_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net5898),
    .D(_02142_),
    .Q_N(_00125_),
    .Q(\TRNG.chunk_index[2] ));
 sg13g2_dfrbp_1 _23277_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net5898),
    .D(_02143_),
    .Q_N(_00124_),
    .Q(\TRNG.chunk_index[3] ));
 sg13g2_dfrbp_1 _23278_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net5898),
    .D(_02144_),
    .Q_N(_00123_),
    .Q(\TRNG.chunk_index[4] ));
 sg13g2_dfrbp_1 _23279_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net5903),
    .D(_02148_),
    .Q_N(_00122_),
    .Q(\TRNG.bit_counter[0] ));
 sg13g2_dfrbp_1 _23280_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net5903),
    .D(net2333),
    .Q_N(_11081_),
    .Q(\TRNG.bit_counter[1] ));
 sg13g2_dfrbp_1 _23281_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net5903),
    .D(_02150_),
    .Q_N(_11082_),
    .Q(\TRNG.bit_counter[2] ));
 sg13g2_dfrbp_1 _23282_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net5903),
    .D(_02151_),
    .Q_N(_11083_),
    .Q(\TRNG.bit_counter[3] ));
 sg13g2_dfrbp_1 _23283_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net5903),
    .D(net2330),
    .Q_N(_11084_),
    .Q(\TRNG.bit_counter[4] ));
 sg13g2_dfrbp_1 _23284_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net5904),
    .D(_02153_),
    .Q_N(_11085_),
    .Q(\TRNG.bit_counter[5] ));
 sg13g2_dfrbp_1 _23285_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net5906),
    .D(_02154_),
    .Q_N(_11086_),
    .Q(\TRNG.bit_counter[6] ));
 sg13g2_dfrbp_1 _23286_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net5903),
    .D(_02155_),
    .Q_N(_11087_),
    .Q(\TRNG.bit_counter[7] ));
 sg13g2_dfrbp_1 _23287_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net5903),
    .D(net2653),
    .Q_N(_00120_),
    .Q(\TRNG.bit_counter[8] ));
 sg13g2_dfrbp_1 _23288_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net5900),
    .D(net5517),
    .Q_N(_09175_),
    .Q(\TRNG.prev_ctrl_mode ));
 sg13g2_tiehi _21254__24 (.L_HI(net24));
 sg13g2_tiehi _21255__25 (.L_HI(net25));
 sg13g2_tiehi _21256__26 (.L_HI(net26));
 sg13g2_tiehi _21257__27 (.L_HI(net27));
 sg13g2_tiehi _21258__28 (.L_HI(net28));
 sg13g2_tiehi _21259__29 (.L_HI(net29));
 sg13g2_tiehi _21260__30 (.L_HI(net30));
 sg13g2_tiehi _21261__31 (.L_HI(net31));
 sg13g2_tiehi _21262__32 (.L_HI(net32));
 sg13g2_tiehi _21263__33 (.L_HI(net33));
 sg13g2_tiehi _21264__34 (.L_HI(net34));
 sg13g2_tiehi _21265__35 (.L_HI(net35));
 sg13g2_tiehi _21266__36 (.L_HI(net36));
 sg13g2_tiehi _21267__37 (.L_HI(net37));
 sg13g2_tiehi _21268__38 (.L_HI(net38));
 sg13g2_tiehi _21269__39 (.L_HI(net39));
 sg13g2_tiehi _21270__40 (.L_HI(net40));
 sg13g2_tiehi _21271__41 (.L_HI(net41));
 sg13g2_tiehi _21272__42 (.L_HI(net42));
 sg13g2_tiehi _21273__43 (.L_HI(net43));
 sg13g2_tiehi _21274__44 (.L_HI(net44));
 sg13g2_tiehi _21275__45 (.L_HI(net45));
 sg13g2_tiehi _21276__46 (.L_HI(net46));
 sg13g2_tiehi _21277__47 (.L_HI(net47));
 sg13g2_tiehi _21278__48 (.L_HI(net48));
 sg13g2_tiehi _21279__49 (.L_HI(net49));
 sg13g2_tiehi _21280__50 (.L_HI(net50));
 sg13g2_tiehi _21281__51 (.L_HI(net51));
 sg13g2_tiehi _21282__52 (.L_HI(net52));
 sg13g2_tiehi _21283__53 (.L_HI(net53));
 sg13g2_tiehi _21284__54 (.L_HI(net54));
 sg13g2_tiehi _22360__55 (.L_HI(net55));
 sg13g2_tiehi _22359__56 (.L_HI(net56));
 sg13g2_tiehi _22358__57 (.L_HI(net57));
 sg13g2_tiehi _22357__58 (.L_HI(net58));
 sg13g2_tiehi _22356__59 (.L_HI(net59));
 sg13g2_tiehi _22355__60 (.L_HI(net60));
 sg13g2_tiehi _22354__61 (.L_HI(net61));
 sg13g2_tiehi _22352__62 (.L_HI(net62));
 sg13g2_tiehi _22343__63 (.L_HI(net63));
 sg13g2_tiehi _22342__64 (.L_HI(net64));
 sg13g2_tiehi _22341__65 (.L_HI(net65));
 sg13g2_tiehi _22340__66 (.L_HI(net66));
 sg13g2_tiehi _22339__67 (.L_HI(net67));
 sg13g2_tiehi _22338__68 (.L_HI(net68));
 sg13g2_tiehi _22337__69 (.L_HI(net69));
 sg13g2_tiehi _22336__70 (.L_HI(net70));
 sg13g2_tiehi _22335__71 (.L_HI(net71));
 sg13g2_tiehi _22334__72 (.L_HI(net72));
 sg13g2_tiehi _22333__73 (.L_HI(net73));
 sg13g2_tiehi _22332__74 (.L_HI(net74));
 sg13g2_tiehi _22331__75 (.L_HI(net75));
 sg13g2_tiehi _22330__76 (.L_HI(net76));
 sg13g2_tiehi _22329__77 (.L_HI(net77));
 sg13g2_tiehi _22328__78 (.L_HI(net78));
 sg13g2_tiehi _22327__79 (.L_HI(net79));
 sg13g2_tiehi _22326__80 (.L_HI(net80));
 sg13g2_tiehi _22325__81 (.L_HI(net81));
 sg13g2_tiehi _22324__82 (.L_HI(net82));
 sg13g2_tiehi _22323__83 (.L_HI(net83));
 sg13g2_tiehi _22322__84 (.L_HI(net84));
 sg13g2_tiehi _22321__85 (.L_HI(net85));
 sg13g2_tiehi _22320__86 (.L_HI(net86));
 sg13g2_tiehi _22319__87 (.L_HI(net87));
 sg13g2_tiehi _22318__88 (.L_HI(net88));
 sg13g2_tiehi _22317__89 (.L_HI(net89));
 sg13g2_tiehi _22316__90 (.L_HI(net90));
 sg13g2_tiehi _22315__91 (.L_HI(net91));
 sg13g2_tiehi _22314__92 (.L_HI(net92));
 sg13g2_tiehi _22313__93 (.L_HI(net93));
 sg13g2_tiehi _22312__94 (.L_HI(net94));
 sg13g2_tiehi _22311__95 (.L_HI(net95));
 sg13g2_tiehi _22310__96 (.L_HI(net96));
 sg13g2_tiehi _22309__97 (.L_HI(net97));
 sg13g2_tiehi _22308__98 (.L_HI(net98));
 sg13g2_tiehi _22307__99 (.L_HI(net99));
 sg13g2_tiehi _22306__100 (.L_HI(net100));
 sg13g2_tiehi _22305__101 (.L_HI(net101));
 sg13g2_tiehi _22304__102 (.L_HI(net102));
 sg13g2_tiehi _22303__103 (.L_HI(net103));
 sg13g2_tiehi _22302__104 (.L_HI(net104));
 sg13g2_tiehi _22301__105 (.L_HI(net105));
 sg13g2_tiehi _22300__106 (.L_HI(net106));
 sg13g2_tiehi _22299__107 (.L_HI(net107));
 sg13g2_tiehi _22298__108 (.L_HI(net108));
 sg13g2_tiehi _22297__109 (.L_HI(net109));
 sg13g2_tiehi _22296__110 (.L_HI(net110));
 sg13g2_tiehi _22295__111 (.L_HI(net111));
 sg13g2_tiehi _22294__112 (.L_HI(net112));
 sg13g2_tiehi _21285__113 (.L_HI(net113));
 sg13g2_tiehi _22293__114 (.L_HI(net114));
 sg13g2_tiehi _22292__115 (.L_HI(net115));
 sg13g2_tiehi _22291__116 (.L_HI(net116));
 sg13g2_tiehi _22290__117 (.L_HI(net117));
 sg13g2_tiehi _22289__118 (.L_HI(net118));
 sg13g2_tiehi _22288__119 (.L_HI(net119));
 sg13g2_tiehi _22287__120 (.L_HI(net120));
 sg13g2_tiehi _22286__121 (.L_HI(net121));
 sg13g2_tiehi _22285__122 (.L_HI(net122));
 sg13g2_tiehi _22284__123 (.L_HI(net123));
 sg13g2_tiehi _22283__124 (.L_HI(net124));
 sg13g2_tiehi _22282__125 (.L_HI(net125));
 sg13g2_tiehi _22281__126 (.L_HI(net126));
 sg13g2_tiehi _22280__127 (.L_HI(net127));
 sg13g2_tiehi _22279__128 (.L_HI(net128));
 sg13g2_tiehi _22278__129 (.L_HI(net129));
 sg13g2_tiehi _22277__130 (.L_HI(net130));
 sg13g2_tiehi _22276__131 (.L_HI(net131));
 sg13g2_tiehi _22275__132 (.L_HI(net132));
 sg13g2_tiehi _22274__133 (.L_HI(net133));
 sg13g2_tiehi _22273__134 (.L_HI(net134));
 sg13g2_tiehi _22272__135 (.L_HI(net135));
 sg13g2_tiehi _22271__136 (.L_HI(net136));
 sg13g2_tiehi _22270__137 (.L_HI(net137));
 sg13g2_tiehi _22269__138 (.L_HI(net138));
 sg13g2_tiehi _22268__139 (.L_HI(net139));
 sg13g2_tiehi _22267__140 (.L_HI(net140));
 sg13g2_tiehi _22266__141 (.L_HI(net141));
 sg13g2_tiehi _22265__142 (.L_HI(net142));
 sg13g2_tiehi _22264__143 (.L_HI(net143));
 sg13g2_tiehi _22263__144 (.L_HI(net144));
 sg13g2_tiehi _22262__145 (.L_HI(net145));
 sg13g2_tiehi _22261__146 (.L_HI(net146));
 sg13g2_tiehi _22260__147 (.L_HI(net147));
 sg13g2_tiehi _22259__148 (.L_HI(net148));
 sg13g2_tiehi _22258__149 (.L_HI(net149));
 sg13g2_tiehi _22257__150 (.L_HI(net150));
 sg13g2_tiehi _22256__151 (.L_HI(net151));
 sg13g2_tiehi _22255__152 (.L_HI(net152));
 sg13g2_tiehi _22254__153 (.L_HI(net153));
 sg13g2_tiehi _22253__154 (.L_HI(net154));
 sg13g2_tiehi _22252__155 (.L_HI(net155));
 sg13g2_tiehi _22251__156 (.L_HI(net156));
 sg13g2_tiehi _22250__157 (.L_HI(net157));
 sg13g2_tiehi _22249__158 (.L_HI(net158));
 sg13g2_tiehi _22248__159 (.L_HI(net159));
 sg13g2_tiehi _22247__160 (.L_HI(net160));
 sg13g2_tiehi _22246__161 (.L_HI(net161));
 sg13g2_tiehi _22245__162 (.L_HI(net162));
 sg13g2_tiehi _22244__163 (.L_HI(net163));
 sg13g2_tiehi _22243__164 (.L_HI(net164));
 sg13g2_tiehi _22242__165 (.L_HI(net165));
 sg13g2_tiehi _22241__166 (.L_HI(net166));
 sg13g2_tiehi _22240__167 (.L_HI(net167));
 sg13g2_tiehi _22239__168 (.L_HI(net168));
 sg13g2_tiehi _22238__169 (.L_HI(net169));
 sg13g2_tiehi _22237__170 (.L_HI(net170));
 sg13g2_tiehi _22236__171 (.L_HI(net171));
 sg13g2_tiehi _22235__172 (.L_HI(net172));
 sg13g2_tiehi _22234__173 (.L_HI(net173));
 sg13g2_tiehi _22233__174 (.L_HI(net174));
 sg13g2_tiehi _22232__175 (.L_HI(net175));
 sg13g2_tiehi _22231__176 (.L_HI(net176));
 sg13g2_tiehi _22230__177 (.L_HI(net177));
 sg13g2_tiehi _22229__178 (.L_HI(net178));
 sg13g2_tiehi _22228__179 (.L_HI(net179));
 sg13g2_tiehi _22227__180 (.L_HI(net180));
 sg13g2_tiehi _22226__181 (.L_HI(net181));
 sg13g2_tiehi _22225__182 (.L_HI(net182));
 sg13g2_tiehi _22224__183 (.L_HI(net183));
 sg13g2_tiehi _22223__184 (.L_HI(net184));
 sg13g2_tiehi _22222__185 (.L_HI(net185));
 sg13g2_tiehi _22221__186 (.L_HI(net186));
 sg13g2_tiehi _22220__187 (.L_HI(net187));
 sg13g2_tiehi _22219__188 (.L_HI(net188));
 sg13g2_tiehi _22218__189 (.L_HI(net189));
 sg13g2_tiehi _22217__190 (.L_HI(net190));
 sg13g2_tiehi _22216__191 (.L_HI(net191));
 sg13g2_tiehi _22215__192 (.L_HI(net192));
 sg13g2_tiehi _22214__193 (.L_HI(net193));
 sg13g2_tiehi _22213__194 (.L_HI(net194));
 sg13g2_tiehi _22212__195 (.L_HI(net195));
 sg13g2_tiehi _22211__196 (.L_HI(net196));
 sg13g2_tiehi _22210__197 (.L_HI(net197));
 sg13g2_tiehi _22209__198 (.L_HI(net198));
 sg13g2_tiehi _22208__199 (.L_HI(net199));
 sg13g2_tiehi _22207__200 (.L_HI(net200));
 sg13g2_tiehi _22206__201 (.L_HI(net201));
 sg13g2_tiehi _22205__202 (.L_HI(net202));
 sg13g2_tiehi _22204__203 (.L_HI(net203));
 sg13g2_tiehi _22203__204 (.L_HI(net204));
 sg13g2_tiehi _22202__205 (.L_HI(net205));
 sg13g2_tiehi _22201__206 (.L_HI(net206));
 sg13g2_tiehi _22200__207 (.L_HI(net207));
 sg13g2_tiehi _22199__208 (.L_HI(net208));
 sg13g2_tiehi _22198__209 (.L_HI(net209));
 sg13g2_tiehi _22197__210 (.L_HI(net210));
 sg13g2_tiehi _22196__211 (.L_HI(net211));
 sg13g2_tiehi _22195__212 (.L_HI(net212));
 sg13g2_tiehi _22194__213 (.L_HI(net213));
 sg13g2_tiehi _22192__214 (.L_HI(net214));
 sg13g2_tiehi _22191__215 (.L_HI(net215));
 sg13g2_tiehi _22190__216 (.L_HI(net216));
 sg13g2_tiehi _22189__217 (.L_HI(net217));
 sg13g2_tiehi _22188__218 (.L_HI(net218));
 sg13g2_tiehi _22187__219 (.L_HI(net219));
 sg13g2_tiehi _22186__220 (.L_HI(net220));
 sg13g2_tiehi _22185__221 (.L_HI(net221));
 sg13g2_tiehi _22184__222 (.L_HI(net222));
 sg13g2_tiehi _22183__223 (.L_HI(net223));
 sg13g2_tiehi _22182__224 (.L_HI(net224));
 sg13g2_tiehi _22181__225 (.L_HI(net225));
 sg13g2_tiehi _22180__226 (.L_HI(net226));
 sg13g2_tiehi _22179__227 (.L_HI(net227));
 sg13g2_tiehi _22178__228 (.L_HI(net228));
 sg13g2_tiehi _22177__229 (.L_HI(net229));
 sg13g2_tiehi _22176__230 (.L_HI(net230));
 sg13g2_tiehi _22175__231 (.L_HI(net231));
 sg13g2_tiehi _22174__232 (.L_HI(net232));
 sg13g2_tiehi _22173__233 (.L_HI(net233));
 sg13g2_tiehi _22172__234 (.L_HI(net234));
 sg13g2_tiehi _22171__235 (.L_HI(net235));
 sg13g2_tiehi _22170__236 (.L_HI(net236));
 sg13g2_tiehi _22169__237 (.L_HI(net237));
 sg13g2_tiehi _22168__238 (.L_HI(net238));
 sg13g2_tiehi _22167__239 (.L_HI(net239));
 sg13g2_tiehi _22166__240 (.L_HI(net240));
 sg13g2_tiehi _22165__241 (.L_HI(net241));
 sg13g2_tiehi _22164__242 (.L_HI(net242));
 sg13g2_tiehi _22163__243 (.L_HI(net243));
 sg13g2_tiehi _22162__244 (.L_HI(net244));
 sg13g2_tiehi _22161__245 (.L_HI(net245));
 sg13g2_tiehi _22160__246 (.L_HI(net246));
 sg13g2_tiehi _22159__247 (.L_HI(net247));
 sg13g2_tiehi _22158__248 (.L_HI(net248));
 sg13g2_tiehi _22157__249 (.L_HI(net249));
 sg13g2_tiehi _22156__250 (.L_HI(net250));
 sg13g2_tiehi _22155__251 (.L_HI(net251));
 sg13g2_tiehi _22154__252 (.L_HI(net252));
 sg13g2_tiehi _22153__253 (.L_HI(net253));
 sg13g2_tiehi _22152__254 (.L_HI(net254));
 sg13g2_tiehi _22151__255 (.L_HI(net255));
 sg13g2_tiehi _22150__256 (.L_HI(net256));
 sg13g2_tiehi _22149__257 (.L_HI(net257));
 sg13g2_tiehi _22148__258 (.L_HI(net258));
 sg13g2_tiehi _22147__259 (.L_HI(net259));
 sg13g2_tiehi _22146__260 (.L_HI(net260));
 sg13g2_tiehi _22145__261 (.L_HI(net261));
 sg13g2_tiehi _22144__262 (.L_HI(net262));
 sg13g2_tiehi _22143__263 (.L_HI(net263));
 sg13g2_tiehi _22142__264 (.L_HI(net264));
 sg13g2_tiehi _22141__265 (.L_HI(net265));
 sg13g2_tiehi _22140__266 (.L_HI(net266));
 sg13g2_tiehi _22139__267 (.L_HI(net267));
 sg13g2_tiehi _22138__268 (.L_HI(net268));
 sg13g2_tiehi _22137__269 (.L_HI(net269));
 sg13g2_tiehi _22136__270 (.L_HI(net270));
 sg13g2_tiehi _22135__271 (.L_HI(net271));
 sg13g2_tiehi _22134__272 (.L_HI(net272));
 sg13g2_tiehi _22133__273 (.L_HI(net273));
 sg13g2_tiehi _22132__274 (.L_HI(net274));
 sg13g2_tiehi _22131__275 (.L_HI(net275));
 sg13g2_tiehi _22130__276 (.L_HI(net276));
 sg13g2_tiehi _22129__277 (.L_HI(net277));
 sg13g2_tiehi _22032__278 (.L_HI(net278));
 sg13g2_tiehi _22031__279 (.L_HI(net279));
 sg13g2_tiehi _22030__280 (.L_HI(net280));
 sg13g2_tiehi _22029__281 (.L_HI(net281));
 sg13g2_tiehi _22028__282 (.L_HI(net282));
 sg13g2_tiehi _22027__283 (.L_HI(net283));
 sg13g2_tiehi _22026__284 (.L_HI(net284));
 sg13g2_tiehi _22025__285 (.L_HI(net285));
 sg13g2_tiehi _21446__286 (.L_HI(net286));
 sg13g2_tiehi _21755__287 (.L_HI(net287));
 sg13g2_tiehi _21756__288 (.L_HI(net288));
 sg13g2_tiehi _21757__289 (.L_HI(net289));
 sg13g2_tiehi _21758__290 (.L_HI(net290));
 sg13g2_tiehi _21759__291 (.L_HI(net291));
 sg13g2_tiehi _21760__292 (.L_HI(net292));
 sg13g2_tiehi _21761__293 (.L_HI(net293));
 sg13g2_tiehi _21762__294 (.L_HI(net294));
 sg13g2_tiehi _21763__295 (.L_HI(net295));
 sg13g2_tiehi _21764__296 (.L_HI(net296));
 sg13g2_tiehi _21765__297 (.L_HI(net297));
 sg13g2_tiehi _21766__298 (.L_HI(net298));
 sg13g2_tiehi _21767__299 (.L_HI(net299));
 sg13g2_tiehi _21768__300 (.L_HI(net300));
 sg13g2_tiehi _21769__301 (.L_HI(net301));
 sg13g2_tiehi _21770__302 (.L_HI(net302));
 sg13g2_tiehi _21771__303 (.L_HI(net303));
 sg13g2_tiehi _21772__304 (.L_HI(net304));
 sg13g2_tiehi _21773__305 (.L_HI(net305));
 sg13g2_tiehi _21774__306 (.L_HI(net306));
 sg13g2_tiehi _21775__307 (.L_HI(net307));
 sg13g2_tiehi _21776__308 (.L_HI(net308));
 sg13g2_tiehi _21777__309 (.L_HI(net309));
 sg13g2_tiehi _21778__310 (.L_HI(net310));
 sg13g2_tiehi _21779__311 (.L_HI(net311));
 sg13g2_tiehi _21780__312 (.L_HI(net312));
 sg13g2_tiehi _21781__313 (.L_HI(net313));
 sg13g2_tiehi _21782__314 (.L_HI(net314));
 sg13g2_tiehi _21783__315 (.L_HI(net315));
 sg13g2_tiehi _21784__316 (.L_HI(net316));
 sg13g2_tiehi _21785__317 (.L_HI(net317));
 sg13g2_tiehi _22024__318 (.L_HI(net318));
 sg13g2_tiehi _22023__319 (.L_HI(net319));
 sg13g2_tiehi _22022__320 (.L_HI(net320));
 sg13g2_tiehi _22021__321 (.L_HI(net321));
 sg13g2_tiehi _22020__322 (.L_HI(net322));
 sg13g2_tiehi _22019__323 (.L_HI(net323));
 sg13g2_tiehi _22018__324 (.L_HI(net324));
 sg13g2_tiehi _22017__325 (.L_HI(net325));
 sg13g2_tiehi _22016__326 (.L_HI(net326));
 sg13g2_tiehi _22015__327 (.L_HI(net327));
 sg13g2_tiehi _22014__328 (.L_HI(net328));
 sg13g2_tiehi _22013__329 (.L_HI(net329));
 sg13g2_tiehi _22012__330 (.L_HI(net330));
 sg13g2_tiehi _22011__331 (.L_HI(net331));
 sg13g2_tiehi _22010__332 (.L_HI(net332));
 sg13g2_tiehi _22009__333 (.L_HI(net333));
 sg13g2_tiehi _22008__334 (.L_HI(net334));
 sg13g2_tiehi _22007__335 (.L_HI(net335));
 sg13g2_tiehi _22006__336 (.L_HI(net336));
 sg13g2_tiehi _22005__337 (.L_HI(net337));
 sg13g2_tiehi _22004__338 (.L_HI(net338));
 sg13g2_tiehi _22003__339 (.L_HI(net339));
 sg13g2_tiehi _22002__340 (.L_HI(net340));
 sg13g2_tiehi _22001__341 (.L_HI(net341));
 sg13g2_tiehi _22000__342 (.L_HI(net342));
 sg13g2_tiehi _21999__343 (.L_HI(net343));
 sg13g2_tiehi _21998__344 (.L_HI(net344));
 sg13g2_tiehi _21997__345 (.L_HI(net345));
 sg13g2_tiehi _21996__346 (.L_HI(net346));
 sg13g2_tiehi _21995__347 (.L_HI(net347));
 sg13g2_tiehi _21994__348 (.L_HI(net348));
 sg13g2_tiehi _21993__349 (.L_HI(net349));
 sg13g2_tiehi _21992__350 (.L_HI(net350));
 sg13g2_tiehi _21991__351 (.L_HI(net351));
 sg13g2_tiehi _21990__352 (.L_HI(net352));
 sg13g2_tiehi _21989__353 (.L_HI(net353));
 sg13g2_tiehi _21988__354 (.L_HI(net354));
 sg13g2_tiehi _21987__355 (.L_HI(net355));
 sg13g2_tiehi _21986__356 (.L_HI(net356));
 sg13g2_tiehi _21985__357 (.L_HI(net357));
 sg13g2_tiehi _21786__358 (.L_HI(net358));
 sg13g2_tiehi _21867__359 (.L_HI(net359));
 sg13g2_tiehi _21868__360 (.L_HI(net360));
 sg13g2_tiehi _21869__361 (.L_HI(net361));
 sg13g2_tiehi _21870__362 (.L_HI(net362));
 sg13g2_tiehi _21871__363 (.L_HI(net363));
 sg13g2_tiehi _21872__364 (.L_HI(net364));
 sg13g2_tiehi _21873__365 (.L_HI(net365));
 sg13g2_tiehi _21874__366 (.L_HI(net366));
 sg13g2_tiehi _21875__367 (.L_HI(net367));
 sg13g2_tiehi _21876__368 (.L_HI(net368));
 sg13g2_tiehi _21877__369 (.L_HI(net369));
 sg13g2_tiehi _21984__370 (.L_HI(net370));
 sg13g2_tiehi _21983__371 (.L_HI(net371));
 sg13g2_tiehi _21982__372 (.L_HI(net372));
 sg13g2_tiehi _21981__373 (.L_HI(net373));
 sg13g2_tiehi _21980__374 (.L_HI(net374));
 sg13g2_tiehi _21979__375 (.L_HI(net375));
 sg13g2_tiehi _21978__376 (.L_HI(net376));
 sg13g2_tiehi _21977__377 (.L_HI(net377));
 sg13g2_tiehi _21976__378 (.L_HI(net378));
 sg13g2_tiehi _21975__379 (.L_HI(net379));
 sg13g2_tiehi _21974__380 (.L_HI(net380));
 sg13g2_tiehi _21973__381 (.L_HI(net381));
 sg13g2_tiehi _21972__382 (.L_HI(net382));
 sg13g2_tiehi _21971__383 (.L_HI(net383));
 sg13g2_tiehi _21970__384 (.L_HI(net384));
 sg13g2_tiehi _21969__385 (.L_HI(net385));
 sg13g2_tiehi _21968__386 (.L_HI(net386));
 sg13g2_tiehi _21967__387 (.L_HI(net387));
 sg13g2_tiehi _21966__388 (.L_HI(net388));
 sg13g2_tiehi _21965__389 (.L_HI(net389));
 sg13g2_tiehi _21964__390 (.L_HI(net390));
 sg13g2_tiehi _21963__391 (.L_HI(net391));
 sg13g2_tiehi _21962__392 (.L_HI(net392));
 sg13g2_tiehi _21961__393 (.L_HI(net393));
 sg13g2_tiehi _21960__394 (.L_HI(net394));
 sg13g2_tiehi _21959__395 (.L_HI(net395));
 sg13g2_tiehi _21958__396 (.L_HI(net396));
 sg13g2_tiehi _21957__397 (.L_HI(net397));
 sg13g2_tiehi _21956__398 (.L_HI(net398));
 sg13g2_tiehi _21955__399 (.L_HI(net399));
 sg13g2_tiehi _21954__400 (.L_HI(net400));
 sg13g2_tiehi _21953__401 (.L_HI(net401));
 sg13g2_tiehi _21952__402 (.L_HI(net402));
 sg13g2_tiehi _21951__403 (.L_HI(net403));
 sg13g2_tiehi _21950__404 (.L_HI(net404));
 sg13g2_tiehi _21949__405 (.L_HI(net405));
 sg13g2_tiehi _21948__406 (.L_HI(net406));
 sg13g2_tiehi _21947__407 (.L_HI(net407));
 sg13g2_tiehi _21946__408 (.L_HI(net408));
 sg13g2_tiehi _21945__409 (.L_HI(net409));
 sg13g2_tiehi _21944__410 (.L_HI(net410));
 sg13g2_tiehi _21943__411 (.L_HI(net411));
 sg13g2_tiehi _21942__412 (.L_HI(net412));
 sg13g2_tiehi _21941__413 (.L_HI(net413));
 sg13g2_tiehi _21940__414 (.L_HI(net414));
 sg13g2_tiehi _21939__415 (.L_HI(net415));
 sg13g2_tiehi _21938__416 (.L_HI(net416));
 sg13g2_tiehi _21937__417 (.L_HI(net417));
 sg13g2_tiehi _21936__418 (.L_HI(net418));
 sg13g2_tiehi _21935__419 (.L_HI(net419));
 sg13g2_tiehi _21934__420 (.L_HI(net420));
 sg13g2_tiehi _21933__421 (.L_HI(net421));
 sg13g2_tiehi _21932__422 (.L_HI(net422));
 sg13g2_tiehi _21931__423 (.L_HI(net423));
 sg13g2_tiehi _21930__424 (.L_HI(net424));
 sg13g2_tiehi _21929__425 (.L_HI(net425));
 sg13g2_tiehi _21928__426 (.L_HI(net426));
 sg13g2_tiehi _21927__427 (.L_HI(net427));
 sg13g2_tiehi _21926__428 (.L_HI(net428));
 sg13g2_tiehi _21925__429 (.L_HI(net429));
 sg13g2_tiehi _21924__430 (.L_HI(net430));
 sg13g2_tiehi _21923__431 (.L_HI(net431));
 sg13g2_tiehi _21922__432 (.L_HI(net432));
 sg13g2_tiehi _21921__433 (.L_HI(net433));
 sg13g2_tiehi _21920__434 (.L_HI(net434));
 sg13g2_tiehi _21919__435 (.L_HI(net435));
 sg13g2_tiehi _21918__436 (.L_HI(net436));
 sg13g2_tiehi _21917__437 (.L_HI(net437));
 sg13g2_tiehi _21916__438 (.L_HI(net438));
 sg13g2_tiehi _21915__439 (.L_HI(net439));
 sg13g2_tiehi _21914__440 (.L_HI(net440));
 sg13g2_tiehi _21913__441 (.L_HI(net441));
 sg13g2_tiehi _21912__442 (.L_HI(net442));
 sg13g2_tiehi _21911__443 (.L_HI(net443));
 sg13g2_tiehi _21910__444 (.L_HI(net444));
 sg13g2_tiehi _21909__445 (.L_HI(net445));
 sg13g2_tiehi _21908__446 (.L_HI(net446));
 sg13g2_tiehi _21907__447 (.L_HI(net447));
 sg13g2_tiehi _21906__448 (.L_HI(net448));
 sg13g2_tiehi _21905__449 (.L_HI(net449));
 sg13g2_tiehi _21904__450 (.L_HI(net450));
 sg13g2_tiehi _21903__451 (.L_HI(net451));
 sg13g2_tiehi _21878__452 (.L_HI(net452));
 sg13g2_tiehi _22033__453 (.L_HI(net453));
 sg13g2_tiehi _22034__454 (.L_HI(net454));
 sg13g2_tiehi _22035__455 (.L_HI(net455));
 sg13g2_tiehi _22036__456 (.L_HI(net456));
 sg13g2_tiehi _22037__457 (.L_HI(net457));
 sg13g2_tiehi _22038__458 (.L_HI(net458));
 sg13g2_tiehi _22039__459 (.L_HI(net459));
 sg13g2_tiehi _22040__460 (.L_HI(net460));
 sg13g2_tiehi _22041__461 (.L_HI(net461));
 sg13g2_tiehi _22042__462 (.L_HI(net462));
 sg13g2_tiehi _22043__463 (.L_HI(net463));
 sg13g2_tiehi _22044__464 (.L_HI(net464));
 sg13g2_tiehi _22045__465 (.L_HI(net465));
 sg13g2_tiehi _22046__466 (.L_HI(net466));
 sg13g2_tiehi _22047__467 (.L_HI(net467));
 sg13g2_tiehi _22048__468 (.L_HI(net468));
 sg13g2_tiehi _22049__469 (.L_HI(net469));
 sg13g2_tiehi _22050__470 (.L_HI(net470));
 sg13g2_tiehi _22051__471 (.L_HI(net471));
 sg13g2_tiehi _22052__472 (.L_HI(net472));
 sg13g2_tiehi _22053__473 (.L_HI(net473));
 sg13g2_tiehi _22054__474 (.L_HI(net474));
 sg13g2_tiehi _22055__475 (.L_HI(net475));
 sg13g2_tiehi _22056__476 (.L_HI(net476));
 sg13g2_tiehi _22057__477 (.L_HI(net477));
 sg13g2_tiehi _22058__478 (.L_HI(net478));
 sg13g2_tiehi _22059__479 (.L_HI(net479));
 sg13g2_tiehi _22060__480 (.L_HI(net480));
 sg13g2_tiehi _22061__481 (.L_HI(net481));
 sg13g2_tiehi _22062__482 (.L_HI(net482));
 sg13g2_tiehi _22063__483 (.L_HI(net483));
 sg13g2_tiehi _22064__484 (.L_HI(net484));
 sg13g2_tiehi _22065__485 (.L_HI(net485));
 sg13g2_tiehi _22066__486 (.L_HI(net486));
 sg13g2_tiehi _22067__487 (.L_HI(net487));
 sg13g2_tiehi _22068__488 (.L_HI(net488));
 sg13g2_tiehi _22069__489 (.L_HI(net489));
 sg13g2_tiehi _22070__490 (.L_HI(net490));
 sg13g2_tiehi _22071__491 (.L_HI(net491));
 sg13g2_tiehi _22072__492 (.L_HI(net492));
 sg13g2_tiehi _22073__493 (.L_HI(net493));
 sg13g2_tiehi _22074__494 (.L_HI(net494));
 sg13g2_tiehi _22075__495 (.L_HI(net495));
 sg13g2_tiehi _22076__496 (.L_HI(net496));
 sg13g2_tiehi _22077__497 (.L_HI(net497));
 sg13g2_tiehi _22078__498 (.L_HI(net498));
 sg13g2_tiehi _22079__499 (.L_HI(net499));
 sg13g2_tiehi _22080__500 (.L_HI(net500));
 sg13g2_tiehi _22081__501 (.L_HI(net501));
 sg13g2_tiehi _22082__502 (.L_HI(net502));
 sg13g2_tiehi _22083__503 (.L_HI(net503));
 sg13g2_tiehi _22084__504 (.L_HI(net504));
 sg13g2_tiehi _22085__505 (.L_HI(net505));
 sg13g2_tiehi _22086__506 (.L_HI(net506));
 sg13g2_tiehi _22087__507 (.L_HI(net507));
 sg13g2_tiehi _22088__508 (.L_HI(net508));
 sg13g2_tiehi _22089__509 (.L_HI(net509));
 sg13g2_tiehi _22090__510 (.L_HI(net510));
 sg13g2_tiehi _22091__511 (.L_HI(net511));
 sg13g2_tiehi _22092__512 (.L_HI(net512));
 sg13g2_tiehi _22093__513 (.L_HI(net513));
 sg13g2_tiehi _22094__514 (.L_HI(net514));
 sg13g2_tiehi _22095__515 (.L_HI(net515));
 sg13g2_tiehi _22096__516 (.L_HI(net516));
 sg13g2_tiehi _22097__517 (.L_HI(net517));
 sg13g2_tiehi _22098__518 (.L_HI(net518));
 sg13g2_tiehi _22099__519 (.L_HI(net519));
 sg13g2_tiehi _22100__520 (.L_HI(net520));
 sg13g2_tiehi _22101__521 (.L_HI(net521));
 sg13g2_tiehi _22102__522 (.L_HI(net522));
 sg13g2_tiehi _22103__523 (.L_HI(net523));
 sg13g2_tiehi _22104__524 (.L_HI(net524));
 sg13g2_tiehi _22105__525 (.L_HI(net525));
 sg13g2_tiehi _22106__526 (.L_HI(net526));
 sg13g2_tiehi _22107__527 (.L_HI(net527));
 sg13g2_tiehi _22108__528 (.L_HI(net528));
 sg13g2_tiehi _22109__529 (.L_HI(net529));
 sg13g2_tiehi _22110__530 (.L_HI(net530));
 sg13g2_tiehi _22111__531 (.L_HI(net531));
 sg13g2_tiehi _22112__532 (.L_HI(net532));
 sg13g2_tiehi _22113__533 (.L_HI(net533));
 sg13g2_tiehi _22114__534 (.L_HI(net534));
 sg13g2_tiehi _22115__535 (.L_HI(net535));
 sg13g2_tiehi _22116__536 (.L_HI(net536));
 sg13g2_tiehi _22117__537 (.L_HI(net537));
 sg13g2_tiehi _22118__538 (.L_HI(net538));
 sg13g2_tiehi _22119__539 (.L_HI(net539));
 sg13g2_tiehi _22120__540 (.L_HI(net540));
 sg13g2_tiehi _22121__541 (.L_HI(net541));
 sg13g2_tiehi _22122__542 (.L_HI(net542));
 sg13g2_tiehi _22123__543 (.L_HI(net543));
 sg13g2_tiehi _22124__544 (.L_HI(net544));
 sg13g2_tiehi _22125__545 (.L_HI(net545));
 sg13g2_tiehi _22126__546 (.L_HI(net546));
 sg13g2_tiehi _22127__547 (.L_HI(net547));
 sg13g2_tiehi _21902__548 (.L_HI(net548));
 sg13g2_tiehi _21901__549 (.L_HI(net549));
 sg13g2_tiehi _21900__550 (.L_HI(net550));
 sg13g2_tiehi _21899__551 (.L_HI(net551));
 sg13g2_tiehi _21898__552 (.L_HI(net552));
 sg13g2_tiehi _21897__553 (.L_HI(net553));
 sg13g2_tiehi _21896__554 (.L_HI(net554));
 sg13g2_tiehi _21895__555 (.L_HI(net555));
 sg13g2_tiehi _21894__556 (.L_HI(net556));
 sg13g2_tiehi _21893__557 (.L_HI(net557));
 sg13g2_tiehi _21892__558 (.L_HI(net558));
 sg13g2_tiehi _21891__559 (.L_HI(net559));
 sg13g2_tiehi _21890__560 (.L_HI(net560));
 sg13g2_tiehi _21889__561 (.L_HI(net561));
 sg13g2_tiehi _21888__562 (.L_HI(net562));
 sg13g2_tiehi _21887__563 (.L_HI(net563));
 sg13g2_tiehi _21886__564 (.L_HI(net564));
 sg13g2_tiehi _21885__565 (.L_HI(net565));
 sg13g2_tiehi _21884__566 (.L_HI(net566));
 sg13g2_tiehi _21883__567 (.L_HI(net567));
 sg13g2_tiehi _21882__568 (.L_HI(net568));
 sg13g2_tiehi _21881__569 (.L_HI(net569));
 sg13g2_tiehi _21880__570 (.L_HI(net570));
 sg13g2_tiehi _21879__571 (.L_HI(net571));
 sg13g2_tiehi _21866__572 (.L_HI(net572));
 sg13g2_tiehi _21865__573 (.L_HI(net573));
 sg13g2_tiehi _21864__574 (.L_HI(net574));
 sg13g2_tiehi _21863__575 (.L_HI(net575));
 sg13g2_tiehi _21862__576 (.L_HI(net576));
 sg13g2_tiehi _21861__577 (.L_HI(net577));
 sg13g2_tiehi _21860__578 (.L_HI(net578));
 sg13g2_tiehi _21859__579 (.L_HI(net579));
 sg13g2_tiehi _21858__580 (.L_HI(net580));
 sg13g2_tiehi _21857__581 (.L_HI(net581));
 sg13g2_tiehi _21856__582 (.L_HI(net582));
 sg13g2_tiehi _21855__583 (.L_HI(net583));
 sg13g2_tiehi _21854__584 (.L_HI(net584));
 sg13g2_tiehi _21853__585 (.L_HI(net585));
 sg13g2_tiehi _21852__586 (.L_HI(net586));
 sg13g2_tiehi _21851__587 (.L_HI(net587));
 sg13g2_tiehi _21850__588 (.L_HI(net588));
 sg13g2_tiehi _21849__589 (.L_HI(net589));
 sg13g2_tiehi _21848__590 (.L_HI(net590));
 sg13g2_tiehi _21847__591 (.L_HI(net591));
 sg13g2_tiehi _21846__592 (.L_HI(net592));
 sg13g2_tiehi _21845__593 (.L_HI(net593));
 sg13g2_tiehi _21844__594 (.L_HI(net594));
 sg13g2_tiehi _21843__595 (.L_HI(net595));
 sg13g2_tiehi _21842__596 (.L_HI(net596));
 sg13g2_tiehi _21841__597 (.L_HI(net597));
 sg13g2_tiehi _21840__598 (.L_HI(net598));
 sg13g2_tiehi _21839__599 (.L_HI(net599));
 sg13g2_tiehi _21838__600 (.L_HI(net600));
 sg13g2_tiehi _21837__601 (.L_HI(net601));
 sg13g2_tiehi _21836__602 (.L_HI(net602));
 sg13g2_tiehi _21835__603 (.L_HI(net603));
 sg13g2_tiehi _21834__604 (.L_HI(net604));
 sg13g2_tiehi _21833__605 (.L_HI(net605));
 sg13g2_tiehi _21832__606 (.L_HI(net606));
 sg13g2_tiehi _21831__607 (.L_HI(net607));
 sg13g2_tiehi _21830__608 (.L_HI(net608));
 sg13g2_tiehi _21829__609 (.L_HI(net609));
 sg13g2_tiehi _21828__610 (.L_HI(net610));
 sg13g2_tiehi _21827__611 (.L_HI(net611));
 sg13g2_tiehi _21826__612 (.L_HI(net612));
 sg13g2_tiehi _21825__613 (.L_HI(net613));
 sg13g2_tiehi _21824__614 (.L_HI(net614));
 sg13g2_tiehi _21823__615 (.L_HI(net615));
 sg13g2_tiehi _21822__616 (.L_HI(net616));
 sg13g2_tiehi _21821__617 (.L_HI(net617));
 sg13g2_tiehi _21820__618 (.L_HI(net618));
 sg13g2_tiehi _21819__619 (.L_HI(net619));
 sg13g2_tiehi _21818__620 (.L_HI(net620));
 sg13g2_tiehi _21817__621 (.L_HI(net621));
 sg13g2_tiehi _21816__622 (.L_HI(net622));
 sg13g2_tiehi _21815__623 (.L_HI(net623));
 sg13g2_tiehi _21814__624 (.L_HI(net624));
 sg13g2_tiehi _21813__625 (.L_HI(net625));
 sg13g2_tiehi _21812__626 (.L_HI(net626));
 sg13g2_tiehi _21811__627 (.L_HI(net627));
 sg13g2_tiehi _21810__628 (.L_HI(net628));
 sg13g2_tiehi _21809__629 (.L_HI(net629));
 sg13g2_tiehi _21808__630 (.L_HI(net630));
 sg13g2_tiehi _21807__631 (.L_HI(net631));
 sg13g2_tiehi _21806__632 (.L_HI(net632));
 sg13g2_tiehi _21805__633 (.L_HI(net633));
 sg13g2_tiehi _21804__634 (.L_HI(net634));
 sg13g2_tiehi _21803__635 (.L_HI(net635));
 sg13g2_tiehi _21802__636 (.L_HI(net636));
 sg13g2_tiehi _21801__637 (.L_HI(net637));
 sg13g2_tiehi _21800__638 (.L_HI(net638));
 sg13g2_tiehi _21799__639 (.L_HI(net639));
 sg13g2_tiehi _21798__640 (.L_HI(net640));
 sg13g2_tiehi _21797__641 (.L_HI(net641));
 sg13g2_tiehi _21796__642 (.L_HI(net642));
 sg13g2_tiehi _21795__643 (.L_HI(net643));
 sg13g2_tiehi _21794__644 (.L_HI(net644));
 sg13g2_tiehi _21793__645 (.L_HI(net645));
 sg13g2_tiehi _21792__646 (.L_HI(net646));
 sg13g2_tiehi _21791__647 (.L_HI(net647));
 sg13g2_tiehi _21790__648 (.L_HI(net648));
 sg13g2_tiehi _21789__649 (.L_HI(net649));
 sg13g2_tiehi _21788__650 (.L_HI(net650));
 sg13g2_tiehi _21787__651 (.L_HI(net651));
 sg13g2_tiehi _21754__652 (.L_HI(net652));
 sg13g2_tiehi _21753__653 (.L_HI(net653));
 sg13g2_tiehi _21752__654 (.L_HI(net654));
 sg13g2_tiehi _21751__655 (.L_HI(net655));
 sg13g2_tiehi _21750__656 (.L_HI(net656));
 sg13g2_tiehi _21749__657 (.L_HI(net657));
 sg13g2_tiehi _21748__658 (.L_HI(net658));
 sg13g2_tiehi _21747__659 (.L_HI(net659));
 sg13g2_tiehi _21746__660 (.L_HI(net660));
 sg13g2_tiehi _21745__661 (.L_HI(net661));
 sg13g2_tiehi _21744__662 (.L_HI(net662));
 sg13g2_tiehi _21743__663 (.L_HI(net663));
 sg13g2_tiehi _21742__664 (.L_HI(net664));
 sg13g2_tiehi _21741__665 (.L_HI(net665));
 sg13g2_tiehi _21740__666 (.L_HI(net666));
 sg13g2_tiehi _21739__667 (.L_HI(net667));
 sg13g2_tiehi _21738__668 (.L_HI(net668));
 sg13g2_tiehi _21737__669 (.L_HI(net669));
 sg13g2_tiehi _21736__670 (.L_HI(net670));
 sg13g2_tiehi _21735__671 (.L_HI(net671));
 sg13g2_tiehi _21734__672 (.L_HI(net672));
 sg13g2_tiehi _21733__673 (.L_HI(net673));
 sg13g2_tiehi _21732__674 (.L_HI(net674));
 sg13g2_tiehi _21731__675 (.L_HI(net675));
 sg13g2_tiehi _21730__676 (.L_HI(net676));
 sg13g2_tiehi _21729__677 (.L_HI(net677));
 sg13g2_tiehi _21728__678 (.L_HI(net678));
 sg13g2_tiehi _21727__679 (.L_HI(net679));
 sg13g2_tiehi _21726__680 (.L_HI(net680));
 sg13g2_tiehi _21725__681 (.L_HI(net681));
 sg13g2_tiehi _21724__682 (.L_HI(net682));
 sg13g2_tiehi _21723__683 (.L_HI(net683));
 sg13g2_tiehi _21722__684 (.L_HI(net684));
 sg13g2_tiehi _21721__685 (.L_HI(net685));
 sg13g2_tiehi _21720__686 (.L_HI(net686));
 sg13g2_tiehi _21719__687 (.L_HI(net687));
 sg13g2_tiehi _21718__688 (.L_HI(net688));
 sg13g2_tiehi _21717__689 (.L_HI(net689));
 sg13g2_tiehi _21716__690 (.L_HI(net690));
 sg13g2_tiehi _21715__691 (.L_HI(net691));
 sg13g2_tiehi _21714__692 (.L_HI(net692));
 sg13g2_tiehi _21713__693 (.L_HI(net693));
 sg13g2_tiehi _21712__694 (.L_HI(net694));
 sg13g2_tiehi _21711__695 (.L_HI(net695));
 sg13g2_tiehi _21710__696 (.L_HI(net696));
 sg13g2_tiehi _21709__697 (.L_HI(net697));
 sg13g2_tiehi _21708__698 (.L_HI(net698));
 sg13g2_tiehi _21707__699 (.L_HI(net699));
 sg13g2_tiehi _21706__700 (.L_HI(net700));
 sg13g2_tiehi _21705__701 (.L_HI(net701));
 sg13g2_tiehi _21704__702 (.L_HI(net702));
 sg13g2_tiehi _21703__703 (.L_HI(net703));
 sg13g2_tiehi _21702__704 (.L_HI(net704));
 sg13g2_tiehi _21701__705 (.L_HI(net705));
 sg13g2_tiehi _21700__706 (.L_HI(net706));
 sg13g2_tiehi _21699__707 (.L_HI(net707));
 sg13g2_tiehi _21698__708 (.L_HI(net708));
 sg13g2_tiehi _21697__709 (.L_HI(net709));
 sg13g2_tiehi _21696__710 (.L_HI(net710));
 sg13g2_tiehi _21695__711 (.L_HI(net711));
 sg13g2_tiehi _21694__712 (.L_HI(net712));
 sg13g2_tiehi _21693__713 (.L_HI(net713));
 sg13g2_tiehi _21692__714 (.L_HI(net714));
 sg13g2_tiehi _21691__715 (.L_HI(net715));
 sg13g2_tiehi _21690__716 (.L_HI(net716));
 sg13g2_tiehi _21689__717 (.L_HI(net717));
 sg13g2_tiehi _21688__718 (.L_HI(net718));
 sg13g2_tiehi _21687__719 (.L_HI(net719));
 sg13g2_tiehi _21686__720 (.L_HI(net720));
 sg13g2_tiehi _21685__721 (.L_HI(net721));
 sg13g2_tiehi _21684__722 (.L_HI(net722));
 sg13g2_tiehi _21683__723 (.L_HI(net723));
 sg13g2_tiehi _21682__724 (.L_HI(net724));
 sg13g2_tiehi _21681__725 (.L_HI(net725));
 sg13g2_tiehi _21680__726 (.L_HI(net726));
 sg13g2_tiehi _21679__727 (.L_HI(net727));
 sg13g2_tiehi _21678__728 (.L_HI(net728));
 sg13g2_tiehi _21677__729 (.L_HI(net729));
 sg13g2_tiehi _21676__730 (.L_HI(net730));
 sg13g2_tiehi _21675__731 (.L_HI(net731));
 sg13g2_tiehi _21674__732 (.L_HI(net732));
 sg13g2_tiehi _21673__733 (.L_HI(net733));
 sg13g2_tiehi _21672__734 (.L_HI(net734));
 sg13g2_tiehi _21671__735 (.L_HI(net735));
 sg13g2_tiehi _21670__736 (.L_HI(net736));
 sg13g2_tiehi _21669__737 (.L_HI(net737));
 sg13g2_tiehi _21668__738 (.L_HI(net738));
 sg13g2_tiehi _21667__739 (.L_HI(net739));
 sg13g2_tiehi _21666__740 (.L_HI(net740));
 sg13g2_tiehi _21665__741 (.L_HI(net741));
 sg13g2_tiehi _21664__742 (.L_HI(net742));
 sg13g2_tiehi _21663__743 (.L_HI(net743));
 sg13g2_tiehi _21662__744 (.L_HI(net744));
 sg13g2_tiehi _21661__745 (.L_HI(net745));
 sg13g2_tiehi _21660__746 (.L_HI(net746));
 sg13g2_tiehi _21659__747 (.L_HI(net747));
 sg13g2_tiehi _21658__748 (.L_HI(net748));
 sg13g2_tiehi _21657__749 (.L_HI(net749));
 sg13g2_tiehi _21656__750 (.L_HI(net750));
 sg13g2_tiehi _21655__751 (.L_HI(net751));
 sg13g2_tiehi _21654__752 (.L_HI(net752));
 sg13g2_tiehi _22128__753 (.L_HI(net753));
 sg13g2_tiehi _21653__754 (.L_HI(net754));
 sg13g2_tiehi _21652__755 (.L_HI(net755));
 sg13g2_tiehi _21651__756 (.L_HI(net756));
 sg13g2_tiehi _21650__757 (.L_HI(net757));
 sg13g2_tiehi _21649__758 (.L_HI(net758));
 sg13g2_tiehi _21648__759 (.L_HI(net759));
 sg13g2_tiehi _21647__760 (.L_HI(net760));
 sg13g2_tiehi _21646__761 (.L_HI(net761));
 sg13g2_tiehi _21645__762 (.L_HI(net762));
 sg13g2_tiehi _22361__763 (.L_HI(net763));
 sg13g2_tiehi _21644__764 (.L_HI(net764));
 sg13g2_tiehi _21643__765 (.L_HI(net765));
 sg13g2_tiehi _21642__766 (.L_HI(net766));
 sg13g2_tiehi _21641__767 (.L_HI(net767));
 sg13g2_tiehi _21640__768 (.L_HI(net768));
 sg13g2_tiehi _21639__769 (.L_HI(net769));
 sg13g2_tiehi _21638__770 (.L_HI(net770));
 sg13g2_tiehi _21637__771 (.L_HI(net771));
 sg13g2_tiehi _21636__772 (.L_HI(net772));
 sg13g2_tiehi _21635__773 (.L_HI(net773));
 sg13g2_tiehi _21634__774 (.L_HI(net774));
 sg13g2_tiehi _21633__775 (.L_HI(net775));
 sg13g2_tiehi _21632__776 (.L_HI(net776));
 sg13g2_tiehi _21631__777 (.L_HI(net777));
 sg13g2_tiehi _21630__778 (.L_HI(net778));
 sg13g2_tiehi _21629__779 (.L_HI(net779));
 sg13g2_tiehi _21628__780 (.L_HI(net780));
 sg13g2_tiehi _21627__781 (.L_HI(net781));
 sg13g2_tiehi _21626__782 (.L_HI(net782));
 sg13g2_tiehi _21625__783 (.L_HI(net783));
 sg13g2_tiehi _21624__784 (.L_HI(net784));
 sg13g2_tiehi _21623__785 (.L_HI(net785));
 sg13g2_tiehi _21622__786 (.L_HI(net786));
 sg13g2_tiehi _21621__787 (.L_HI(net787));
 sg13g2_tiehi _21620__788 (.L_HI(net788));
 sg13g2_tiehi _21619__789 (.L_HI(net789));
 sg13g2_tiehi _21618__790 (.L_HI(net790));
 sg13g2_tiehi _21617__791 (.L_HI(net791));
 sg13g2_tiehi _21616__792 (.L_HI(net792));
 sg13g2_tiehi _21615__793 (.L_HI(net793));
 sg13g2_tiehi _21614__794 (.L_HI(net794));
 sg13g2_tiehi _21613__795 (.L_HI(net795));
 sg13g2_tiehi _21612__796 (.L_HI(net796));
 sg13g2_tiehi _21611__797 (.L_HI(net797));
 sg13g2_tiehi _21610__798 (.L_HI(net798));
 sg13g2_tiehi _21609__799 (.L_HI(net799));
 sg13g2_tiehi _21608__800 (.L_HI(net800));
 sg13g2_tiehi _21607__801 (.L_HI(net801));
 sg13g2_tiehi _21606__802 (.L_HI(net802));
 sg13g2_tiehi _21605__803 (.L_HI(net803));
 sg13g2_tiehi _21604__804 (.L_HI(net804));
 sg13g2_tiehi _21603__805 (.L_HI(net805));
 sg13g2_tiehi _21602__806 (.L_HI(net806));
 sg13g2_tiehi _21601__807 (.L_HI(net807));
 sg13g2_tiehi _21600__808 (.L_HI(net808));
 sg13g2_tiehi _21599__809 (.L_HI(net809));
 sg13g2_tiehi _21598__810 (.L_HI(net810));
 sg13g2_tiehi _21597__811 (.L_HI(net811));
 sg13g2_tiehi _21596__812 (.L_HI(net812));
 sg13g2_tiehi _21595__813 (.L_HI(net813));
 sg13g2_tiehi _21594__814 (.L_HI(net814));
 sg13g2_tiehi _21593__815 (.L_HI(net815));
 sg13g2_tiehi _21592__816 (.L_HI(net816));
 sg13g2_tiehi _21591__817 (.L_HI(net817));
 sg13g2_tiehi _21590__818 (.L_HI(net818));
 sg13g2_tiehi _21589__819 (.L_HI(net819));
 sg13g2_tiehi _21588__820 (.L_HI(net820));
 sg13g2_tiehi _21587__821 (.L_HI(net821));
 sg13g2_tiehi _21586__822 (.L_HI(net822));
 sg13g2_tiehi _21585__823 (.L_HI(net823));
 sg13g2_tiehi _21584__824 (.L_HI(net824));
 sg13g2_tiehi _21583__825 (.L_HI(net825));
 sg13g2_tiehi _21582__826 (.L_HI(net826));
 sg13g2_tiehi _21581__827 (.L_HI(net827));
 sg13g2_tiehi _21580__828 (.L_HI(net828));
 sg13g2_tiehi _21579__829 (.L_HI(net829));
 sg13g2_tiehi _21578__830 (.L_HI(net830));
 sg13g2_tiehi _21577__831 (.L_HI(net831));
 sg13g2_tiehi _21576__832 (.L_HI(net832));
 sg13g2_tiehi _21575__833 (.L_HI(net833));
 sg13g2_tiehi _21574__834 (.L_HI(net834));
 sg13g2_tiehi _21573__835 (.L_HI(net835));
 sg13g2_tiehi _21572__836 (.L_HI(net836));
 sg13g2_tiehi _21571__837 (.L_HI(net837));
 sg13g2_tiehi _21570__838 (.L_HI(net838));
 sg13g2_tiehi _21569__839 (.L_HI(net839));
 sg13g2_tiehi _21568__840 (.L_HI(net840));
 sg13g2_tiehi _21567__841 (.L_HI(net841));
 sg13g2_tiehi _21566__842 (.L_HI(net842));
 sg13g2_tiehi _21565__843 (.L_HI(net843));
 sg13g2_tiehi _21564__844 (.L_HI(net844));
 sg13g2_tiehi _21563__845 (.L_HI(net845));
 sg13g2_tiehi _21562__846 (.L_HI(net846));
 sg13g2_tiehi _21561__847 (.L_HI(net847));
 sg13g2_tiehi _21560__848 (.L_HI(net848));
 sg13g2_tiehi _21559__849 (.L_HI(net849));
 sg13g2_tiehi _21558__850 (.L_HI(net850));
 sg13g2_tiehi _21557__851 (.L_HI(net851));
 sg13g2_tiehi _21556__852 (.L_HI(net852));
 sg13g2_tiehi _21555__853 (.L_HI(net853));
 sg13g2_tiehi _21554__854 (.L_HI(net854));
 sg13g2_tiehi _21553__855 (.L_HI(net855));
 sg13g2_tiehi _21552__856 (.L_HI(net856));
 sg13g2_tiehi _21551__857 (.L_HI(net857));
 sg13g2_tiehi _21550__858 (.L_HI(net858));
 sg13g2_tiehi _21549__859 (.L_HI(net859));
 sg13g2_tiehi _21548__860 (.L_HI(net860));
 sg13g2_tiehi _21547__861 (.L_HI(net861));
 sg13g2_tiehi _21546__862 (.L_HI(net862));
 sg13g2_tiehi _21545__863 (.L_HI(net863));
 sg13g2_tiehi _21544__864 (.L_HI(net864));
 sg13g2_tiehi _21543__865 (.L_HI(net865));
 sg13g2_tiehi _21542__866 (.L_HI(net866));
 sg13g2_tiehi _21541__867 (.L_HI(net867));
 sg13g2_tiehi _21540__868 (.L_HI(net868));
 sg13g2_tiehi _21539__869 (.L_HI(net869));
 sg13g2_tiehi _21538__870 (.L_HI(net870));
 sg13g2_tiehi _21537__871 (.L_HI(net871));
 sg13g2_tiehi _21536__872 (.L_HI(net872));
 sg13g2_tiehi _21535__873 (.L_HI(net873));
 sg13g2_tiehi _21534__874 (.L_HI(net874));
 sg13g2_tiehi _21533__875 (.L_HI(net875));
 sg13g2_tiehi _21532__876 (.L_HI(net876));
 sg13g2_tiehi _21531__877 (.L_HI(net877));
 sg13g2_tiehi _21530__878 (.L_HI(net878));
 sg13g2_tiehi _21529__879 (.L_HI(net879));
 sg13g2_tiehi _21528__880 (.L_HI(net880));
 sg13g2_tiehi _21527__881 (.L_HI(net881));
 sg13g2_tiehi _21526__882 (.L_HI(net882));
 sg13g2_tiehi _21525__883 (.L_HI(net883));
 sg13g2_tiehi _21524__884 (.L_HI(net884));
 sg13g2_tiehi _21523__885 (.L_HI(net885));
 sg13g2_tiehi _21522__886 (.L_HI(net886));
 sg13g2_tiehi _21521__887 (.L_HI(net887));
 sg13g2_tiehi _21520__888 (.L_HI(net888));
 sg13g2_tiehi _21519__889 (.L_HI(net889));
 sg13g2_tiehi _21518__890 (.L_HI(net890));
 sg13g2_tiehi _21517__891 (.L_HI(net891));
 sg13g2_tiehi _21516__892 (.L_HI(net892));
 sg13g2_tiehi _21515__893 (.L_HI(net893));
 sg13g2_tiehi _21514__894 (.L_HI(net894));
 sg13g2_tiehi _21513__895 (.L_HI(net895));
 sg13g2_tiehi _21512__896 (.L_HI(net896));
 sg13g2_tiehi _21511__897 (.L_HI(net897));
 sg13g2_tiehi _21510__898 (.L_HI(net898));
 sg13g2_tiehi _21509__899 (.L_HI(net899));
 sg13g2_tiehi _21508__900 (.L_HI(net900));
 sg13g2_tiehi _21507__901 (.L_HI(net901));
 sg13g2_tiehi _21506__902 (.L_HI(net902));
 sg13g2_tiehi _21505__903 (.L_HI(net903));
 sg13g2_tiehi _21504__904 (.L_HI(net904));
 sg13g2_tiehi _21503__905 (.L_HI(net905));
 sg13g2_tiehi _21502__906 (.L_HI(net906));
 sg13g2_tiehi _21501__907 (.L_HI(net907));
 sg13g2_tiehi _21500__908 (.L_HI(net908));
 sg13g2_tiehi _21499__909 (.L_HI(net909));
 sg13g2_tiehi _21498__910 (.L_HI(net910));
 sg13g2_tiehi _21497__911 (.L_HI(net911));
 sg13g2_tiehi _21496__912 (.L_HI(net912));
 sg13g2_tiehi _21495__913 (.L_HI(net913));
 sg13g2_tiehi _21494__914 (.L_HI(net914));
 sg13g2_tiehi _21493__915 (.L_HI(net915));
 sg13g2_tiehi _21492__916 (.L_HI(net916));
 sg13g2_tiehi _21491__917 (.L_HI(net917));
 sg13g2_tiehi _21490__918 (.L_HI(net918));
 sg13g2_tiehi _21489__919 (.L_HI(net919));
 sg13g2_tiehi _21488__920 (.L_HI(net920));
 sg13g2_tiehi _21487__921 (.L_HI(net921));
 sg13g2_tiehi _21486__922 (.L_HI(net922));
 sg13g2_tiehi _21485__923 (.L_HI(net923));
 sg13g2_tiehi _21484__924 (.L_HI(net924));
 sg13g2_tiehi _21483__925 (.L_HI(net925));
 sg13g2_tiehi _21482__926 (.L_HI(net926));
 sg13g2_tiehi _21481__927 (.L_HI(net927));
 sg13g2_tiehi _21480__928 (.L_HI(net928));
 sg13g2_tiehi _21479__929 (.L_HI(net929));
 sg13g2_tiehi _21478__930 (.L_HI(net930));
 sg13g2_tiehi _21477__931 (.L_HI(net931));
 sg13g2_tiehi _21476__932 (.L_HI(net932));
 sg13g2_tiehi _21475__933 (.L_HI(net933));
 sg13g2_tiehi _21474__934 (.L_HI(net934));
 sg13g2_tiehi _21473__935 (.L_HI(net935));
 sg13g2_tiehi _21472__936 (.L_HI(net936));
 sg13g2_tiehi _21471__937 (.L_HI(net937));
 sg13g2_tiehi _21470__938 (.L_HI(net938));
 sg13g2_tiehi _21469__939 (.L_HI(net939));
 sg13g2_tiehi _21468__940 (.L_HI(net940));
 sg13g2_tiehi _21467__941 (.L_HI(net941));
 sg13g2_tiehi _21466__942 (.L_HI(net942));
 sg13g2_tiehi _21465__943 (.L_HI(net943));
 sg13g2_tiehi _21464__944 (.L_HI(net944));
 sg13g2_tiehi _21463__945 (.L_HI(net945));
 sg13g2_tiehi _21462__946 (.L_HI(net946));
 sg13g2_tiehi _21461__947 (.L_HI(net947));
 sg13g2_tiehi _21460__948 (.L_HI(net948));
 sg13g2_tiehi _21459__949 (.L_HI(net949));
 sg13g2_tiehi _21458__950 (.L_HI(net950));
 sg13g2_tiehi _21457__951 (.L_HI(net951));
 sg13g2_tiehi _21456__952 (.L_HI(net952));
 sg13g2_tiehi _21455__953 (.L_HI(net953));
 sg13g2_tiehi _21454__954 (.L_HI(net954));
 sg13g2_tiehi _21453__955 (.L_HI(net955));
 sg13g2_tiehi _21452__956 (.L_HI(net956));
 sg13g2_tiehi _21451__957 (.L_HI(net957));
 sg13g2_tiehi _21450__958 (.L_HI(net958));
 sg13g2_tiehi _21449__959 (.L_HI(net959));
 sg13g2_tiehi _21448__960 (.L_HI(net960));
 sg13g2_tiehi _21447__961 (.L_HI(net961));
 sg13g2_tiehi _21445__962 (.L_HI(net962));
 sg13g2_tiehi _21444__963 (.L_HI(net963));
 sg13g2_tiehi _21443__964 (.L_HI(net964));
 sg13g2_tiehi _21442__965 (.L_HI(net965));
 sg13g2_tiehi _21441__966 (.L_HI(net966));
 sg13g2_tiehi _21440__967 (.L_HI(net967));
 sg13g2_tiehi _21439__968 (.L_HI(net968));
 sg13g2_tiehi _21438__969 (.L_HI(net969));
 sg13g2_tiehi _21437__970 (.L_HI(net970));
 sg13g2_tiehi _21436__971 (.L_HI(net971));
 sg13g2_tiehi _21435__972 (.L_HI(net972));
 sg13g2_tiehi _21434__973 (.L_HI(net973));
 sg13g2_tiehi _21433__974 (.L_HI(net974));
 sg13g2_tiehi _21432__975 (.L_HI(net975));
 sg13g2_tiehi _21431__976 (.L_HI(net976));
 sg13g2_tiehi _21430__977 (.L_HI(net977));
 sg13g2_tiehi _21429__978 (.L_HI(net978));
 sg13g2_tiehi _21428__979 (.L_HI(net979));
 sg13g2_tiehi _21427__980 (.L_HI(net980));
 sg13g2_tiehi _21426__981 (.L_HI(net981));
 sg13g2_tiehi _21425__982 (.L_HI(net982));
 sg13g2_tiehi _21424__983 (.L_HI(net983));
 sg13g2_tiehi _21423__984 (.L_HI(net984));
 sg13g2_tiehi _21422__985 (.L_HI(net985));
 sg13g2_tiehi _21421__986 (.L_HI(net986));
 sg13g2_tiehi _21420__987 (.L_HI(net987));
 sg13g2_tiehi _21419__988 (.L_HI(net988));
 sg13g2_tiehi _21418__989 (.L_HI(net989));
 sg13g2_tiehi _21417__990 (.L_HI(net990));
 sg13g2_tiehi _21416__991 (.L_HI(net991));
 sg13g2_tiehi _21415__992 (.L_HI(net992));
 sg13g2_tiehi _21414__993 (.L_HI(net993));
 sg13g2_tiehi _21413__994 (.L_HI(net994));
 sg13g2_tiehi _21412__995 (.L_HI(net995));
 sg13g2_tiehi _21411__996 (.L_HI(net996));
 sg13g2_tiehi _21410__997 (.L_HI(net997));
 sg13g2_tiehi _21409__998 (.L_HI(net998));
 sg13g2_tiehi _21408__999 (.L_HI(net999));
 sg13g2_tiehi _21407__1000 (.L_HI(net1000));
 sg13g2_tiehi _21406__1001 (.L_HI(net1001));
 sg13g2_tiehi _21405__1002 (.L_HI(net1002));
 sg13g2_tiehi _21404__1003 (.L_HI(net1003));
 sg13g2_tiehi _21403__1004 (.L_HI(net1004));
 sg13g2_tiehi _21402__1005 (.L_HI(net1005));
 sg13g2_tiehi _21401__1006 (.L_HI(net1006));
 sg13g2_tiehi _21400__1007 (.L_HI(net1007));
 sg13g2_tiehi _21399__1008 (.L_HI(net1008));
 sg13g2_tiehi _21398__1009 (.L_HI(net1009));
 sg13g2_tiehi _21397__1010 (.L_HI(net1010));
 sg13g2_tiehi _21396__1011 (.L_HI(net1011));
 sg13g2_tiehi _21395__1012 (.L_HI(net1012));
 sg13g2_tiehi _21394__1013 (.L_HI(net1013));
 sg13g2_tiehi _21393__1014 (.L_HI(net1014));
 sg13g2_tiehi _21392__1015 (.L_HI(net1015));
 sg13g2_tiehi _21391__1016 (.L_HI(net1016));
 sg13g2_tiehi _21390__1017 (.L_HI(net1017));
 sg13g2_tiehi _21389__1018 (.L_HI(net1018));
 sg13g2_tiehi _21388__1019 (.L_HI(net1019));
 sg13g2_tiehi _21387__1020 (.L_HI(net1020));
 sg13g2_tiehi _21386__1021 (.L_HI(net1021));
 sg13g2_tiehi _21385__1022 (.L_HI(net1022));
 sg13g2_tiehi _21384__1023 (.L_HI(net1023));
 sg13g2_tiehi _21383__1024 (.L_HI(net1024));
 sg13g2_tiehi _21382__1025 (.L_HI(net1025));
 sg13g2_tiehi _21381__1026 (.L_HI(net1026));
 sg13g2_tiehi _21380__1027 (.L_HI(net1027));
 sg13g2_tiehi _21379__1028 (.L_HI(net1028));
 sg13g2_tiehi _21378__1029 (.L_HI(net1029));
 sg13g2_tiehi _21377__1030 (.L_HI(net1030));
 sg13g2_tiehi _21376__1031 (.L_HI(net1031));
 sg13g2_tiehi _21375__1032 (.L_HI(net1032));
 sg13g2_tiehi _21374__1033 (.L_HI(net1033));
 sg13g2_tiehi _21373__1034 (.L_HI(net1034));
 sg13g2_tiehi _21372__1035 (.L_HI(net1035));
 sg13g2_tiehi _21371__1036 (.L_HI(net1036));
 sg13g2_tiehi _21370__1037 (.L_HI(net1037));
 sg13g2_tiehi _21369__1038 (.L_HI(net1038));
 sg13g2_tiehi _21368__1039 (.L_HI(net1039));
 sg13g2_tiehi _21367__1040 (.L_HI(net1040));
 sg13g2_tiehi _21366__1041 (.L_HI(net1041));
 sg13g2_tiehi _21365__1042 (.L_HI(net1042));
 sg13g2_tiehi _21364__1043 (.L_HI(net1043));
 sg13g2_tiehi _21363__1044 (.L_HI(net1044));
 sg13g2_tiehi _21362__1045 (.L_HI(net1045));
 sg13g2_tiehi _21361__1046 (.L_HI(net1046));
 sg13g2_tiehi _21360__1047 (.L_HI(net1047));
 sg13g2_tiehi _21359__1048 (.L_HI(net1048));
 sg13g2_tiehi _21358__1049 (.L_HI(net1049));
 sg13g2_tiehi _21357__1050 (.L_HI(net1050));
 sg13g2_tiehi _21356__1051 (.L_HI(net1051));
 sg13g2_tiehi _21355__1052 (.L_HI(net1052));
 sg13g2_tiehi _21354__1053 (.L_HI(net1053));
 sg13g2_tiehi _21353__1054 (.L_HI(net1054));
 sg13g2_tiehi _21352__1055 (.L_HI(net1055));
 sg13g2_tiehi _21351__1056 (.L_HI(net1056));
 sg13g2_tiehi _21350__1057 (.L_HI(net1057));
 sg13g2_tiehi _21349__1058 (.L_HI(net1058));
 sg13g2_tiehi _21348__1059 (.L_HI(net1059));
 sg13g2_tiehi _21347__1060 (.L_HI(net1060));
 sg13g2_tiehi _21346__1061 (.L_HI(net1061));
 sg13g2_tiehi _21345__1062 (.L_HI(net1062));
 sg13g2_tiehi _21344__1063 (.L_HI(net1063));
 sg13g2_tiehi _21343__1064 (.L_HI(net1064));
 sg13g2_tiehi _21342__1065 (.L_HI(net1065));
 sg13g2_tiehi _21341__1066 (.L_HI(net1066));
 sg13g2_tiehi _21340__1067 (.L_HI(net1067));
 sg13g2_tiehi _21339__1068 (.L_HI(net1068));
 sg13g2_tiehi _21338__1069 (.L_HI(net1069));
 sg13g2_tiehi _21337__1070 (.L_HI(net1070));
 sg13g2_tiehi _21336__1071 (.L_HI(net1071));
 sg13g2_tiehi _21335__1072 (.L_HI(net1072));
 sg13g2_tiehi _21334__1073 (.L_HI(net1073));
 sg13g2_tiehi _21333__1074 (.L_HI(net1074));
 sg13g2_tiehi _21332__1075 (.L_HI(net1075));
 sg13g2_tiehi _21331__1076 (.L_HI(net1076));
 sg13g2_tiehi _21330__1077 (.L_HI(net1077));
 sg13g2_tiehi _21329__1078 (.L_HI(net1078));
 sg13g2_tiehi _21328__1079 (.L_HI(net1079));
 sg13g2_tiehi _21327__1080 (.L_HI(net1080));
 sg13g2_tiehi _21326__1081 (.L_HI(net1081));
 sg13g2_tiehi _21325__1082 (.L_HI(net1082));
 sg13g2_tiehi _21324__1083 (.L_HI(net1083));
 sg13g2_tiehi _21323__1084 (.L_HI(net1084));
 sg13g2_tiehi _21322__1085 (.L_HI(net1085));
 sg13g2_tiehi _21321__1086 (.L_HI(net1086));
 sg13g2_tiehi _21320__1087 (.L_HI(net1087));
 sg13g2_tiehi _21319__1088 (.L_HI(net1088));
 sg13g2_tiehi _21318__1089 (.L_HI(net1089));
 sg13g2_tiehi _21317__1090 (.L_HI(net1090));
 sg13g2_tiehi _21316__1091 (.L_HI(net1091));
 sg13g2_tiehi _21315__1092 (.L_HI(net1092));
 sg13g2_tiehi _21314__1093 (.L_HI(net1093));
 sg13g2_tiehi _21313__1094 (.L_HI(net1094));
 sg13g2_tiehi _21312__1095 (.L_HI(net1095));
 sg13g2_tiehi _21311__1096 (.L_HI(net1096));
 sg13g2_tiehi _21310__1097 (.L_HI(net1097));
 sg13g2_tiehi _21309__1098 (.L_HI(net1098));
 sg13g2_tiehi _21308__1099 (.L_HI(net1099));
 sg13g2_tiehi _21307__1100 (.L_HI(net1100));
 sg13g2_tiehi _21306__1101 (.L_HI(net1101));
 sg13g2_tiehi _21305__1102 (.L_HI(net1102));
 sg13g2_tiehi _21304__1103 (.L_HI(net1103));
 sg13g2_tiehi _21303__1104 (.L_HI(net1104));
 sg13g2_tiehi _21302__1105 (.L_HI(net1105));
 sg13g2_tiehi _21301__1106 (.L_HI(net1106));
 sg13g2_tiehi _21300__1107 (.L_HI(net1107));
 sg13g2_tiehi _21299__1108 (.L_HI(net1108));
 sg13g2_tiehi _21298__1109 (.L_HI(net1109));
 sg13g2_tiehi _21297__1110 (.L_HI(net1110));
 sg13g2_tiehi _21296__1111 (.L_HI(net1111));
 sg13g2_tiehi _21295__1112 (.L_HI(net1112));
 sg13g2_tiehi _21294__1113 (.L_HI(net1113));
 sg13g2_tiehi _21293__1114 (.L_HI(net1114));
 sg13g2_tiehi _21292__1115 (.L_HI(net1115));
 sg13g2_tiehi _21291__1116 (.L_HI(net1116));
 sg13g2_tiehi _21290__1117 (.L_HI(net1117));
 sg13g2_tiehi _21289__1118 (.L_HI(net1118));
 sg13g2_tiehi _21288__1119 (.L_HI(net1119));
 sg13g2_tiehi _21287__1120 (.L_HI(net1120));
 sg13g2_tiehi _21286__1121 (.L_HI(net1121));
 sg13g2_tiehi _21253__1122 (.L_HI(net1122));
 sg13g2_tiehi _21252__1123 (.L_HI(net1123));
 sg13g2_tiehi _21251__1124 (.L_HI(net1124));
 sg13g2_tiehi _21250__1125 (.L_HI(net1125));
 sg13g2_tiehi _21249__1126 (.L_HI(net1126));
 sg13g2_tiehi _21248__1127 (.L_HI(net1127));
 sg13g2_tiehi _21247__1128 (.L_HI(net1128));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_6_3_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_bilal_trng_3 (.L_LO(net3));
 sg13g2_tielo tt_um_bilal_trng_4 (.L_LO(net4));
 sg13g2_tielo tt_um_bilal_trng_5 (.L_LO(net5));
 sg13g2_tielo tt_um_bilal_trng_6 (.L_LO(net6));
 sg13g2_tielo tt_um_bilal_trng_7 (.L_LO(net7));
 sg13g2_tielo tt_um_bilal_trng_8 (.L_LO(net8));
 sg13g2_tielo tt_um_bilal_trng_9 (.L_LO(net9));
 sg13g2_tielo tt_um_bilal_trng_10 (.L_LO(net10));
 sg13g2_tielo tt_um_bilal_trng_11 (.L_LO(net11));
 sg13g2_tielo tt_um_bilal_trng_12 (.L_LO(net12));
 sg13g2_tielo tt_um_bilal_trng_13 (.L_LO(net13));
 sg13g2_tielo tt_um_bilal_trng_14 (.L_LO(net14));
 sg13g2_tielo tt_um_bilal_trng_15 (.L_LO(net15));
 sg13g2_tielo tt_um_bilal_trng_16 (.L_LO(net16));
 sg13g2_tielo tt_um_bilal_trng_17 (.L_LO(net17));
 sg13g2_tielo tt_um_bilal_trng_18 (.L_LO(net18));
 sg13g2_tielo tt_um_bilal_trng_19 (.L_LO(net19));
 sg13g2_tielo tt_um_bilal_trng_20 (.L_LO(net20));
 sg13g2_tielo tt_um_bilal_trng_21 (.L_LO(net21));
 sg13g2_tielo tt_um_bilal_trng_22 (.L_LO(net22));
 sg13g2_tiehi _21246__23 (.L_HI(net23));
 sg13g2_buf_2 _24416_ (.A(\TRNG.Repetition_Count_Test.failure ),
    .X(uo_out[0]));
 sg13g2_buf_2 _24417_ (.A(\TRNG.hash_rdy ),
    .X(uo_out[1]));
 sg13g2_buf_2 _24418_ (.A(\TRNG.UART_Tx ),
    .X(uo_out[2]));
 sg13g2_buf_4 fanout4555 (.X(net4555),
    .A(net4556));
 sg13g2_buf_4 fanout4556 (.X(net4556),
    .A(_03091_));
 sg13g2_buf_2 fanout4557 (.A(net4558),
    .X(net4557));
 sg13g2_buf_2 fanout4558 (.A(net4559),
    .X(net4558));
 sg13g2_buf_1 fanout4559 (.A(_02255_),
    .X(net4559));
 sg13g2_buf_2 fanout4560 (.A(net4561),
    .X(net4560));
 sg13g2_buf_2 fanout4561 (.A(_02255_),
    .X(net4561));
 sg13g2_buf_2 fanout4562 (.A(net4566),
    .X(net4562));
 sg13g2_buf_2 fanout4563 (.A(net4566),
    .X(net4563));
 sg13g2_buf_2 fanout4564 (.A(net4566),
    .X(net4564));
 sg13g2_buf_2 fanout4565 (.A(net4566),
    .X(net4565));
 sg13g2_buf_2 fanout4566 (.A(_02255_),
    .X(net4566));
 sg13g2_buf_2 fanout4567 (.A(net4570),
    .X(net4567));
 sg13g2_buf_2 fanout4568 (.A(net4570),
    .X(net4568));
 sg13g2_buf_4 fanout4569 (.X(net4569),
    .A(net4570));
 sg13g2_buf_2 fanout4570 (.A(_08890_),
    .X(net4570));
 sg13g2_buf_2 fanout4571 (.A(net4572),
    .X(net4571));
 sg13g2_buf_2 fanout4572 (.A(net4588),
    .X(net4572));
 sg13g2_buf_2 fanout4573 (.A(net4574),
    .X(net4573));
 sg13g2_buf_2 fanout4574 (.A(net4576),
    .X(net4574));
 sg13g2_buf_2 fanout4575 (.A(net4576),
    .X(net4575));
 sg13g2_buf_2 fanout4576 (.A(net4588),
    .X(net4576));
 sg13g2_buf_2 fanout4577 (.A(net4581),
    .X(net4577));
 sg13g2_buf_2 fanout4578 (.A(net4581),
    .X(net4578));
 sg13g2_buf_2 fanout4579 (.A(net4581),
    .X(net4579));
 sg13g2_buf_1 fanout4580 (.A(net4581),
    .X(net4580));
 sg13g2_buf_1 fanout4581 (.A(net4587),
    .X(net4581));
 sg13g2_buf_2 fanout4582 (.A(net4586),
    .X(net4582));
 sg13g2_buf_2 fanout4583 (.A(net4586),
    .X(net4583));
 sg13g2_buf_2 fanout4584 (.A(net4586),
    .X(net4584));
 sg13g2_buf_1 fanout4585 (.A(net4586),
    .X(net4585));
 sg13g2_buf_1 fanout4586 (.A(net4587),
    .X(net4586));
 sg13g2_buf_2 fanout4587 (.A(net4588),
    .X(net4587));
 sg13g2_buf_2 fanout4588 (.A(_04949_),
    .X(net4588));
 sg13g2_buf_2 fanout4589 (.A(net4592),
    .X(net4589));
 sg13g2_buf_2 fanout4590 (.A(net4592),
    .X(net4590));
 sg13g2_buf_2 fanout4591 (.A(net4592),
    .X(net4591));
 sg13g2_buf_2 fanout4592 (.A(net4597),
    .X(net4592));
 sg13g2_buf_2 fanout4593 (.A(net4594),
    .X(net4593));
 sg13g2_buf_2 fanout4594 (.A(net4596),
    .X(net4594));
 sg13g2_buf_2 fanout4595 (.A(net4596),
    .X(net4595));
 sg13g2_buf_1 fanout4596 (.A(net4597),
    .X(net4596));
 sg13g2_buf_4 fanout4597 (.X(net4597),
    .A(net4606));
 sg13g2_buf_2 fanout4598 (.A(net4601),
    .X(net4598));
 sg13g2_buf_2 fanout4599 (.A(net4601),
    .X(net4599));
 sg13g2_buf_2 fanout4600 (.A(net4601),
    .X(net4600));
 sg13g2_buf_2 fanout4601 (.A(net4606),
    .X(net4601));
 sg13g2_buf_2 fanout4602 (.A(net4605),
    .X(net4602));
 sg13g2_buf_2 fanout4603 (.A(net4605),
    .X(net4603));
 sg13g2_buf_1 fanout4604 (.A(net4605),
    .X(net4604));
 sg13g2_buf_1 fanout4605 (.A(net4606),
    .X(net4605));
 sg13g2_buf_4 fanout4606 (.X(net4606),
    .A(_04949_));
 sg13g2_buf_2 fanout4607 (.A(net4615),
    .X(net4607));
 sg13g2_buf_1 fanout4608 (.A(net4615),
    .X(net4608));
 sg13g2_buf_2 fanout4609 (.A(net4615),
    .X(net4609));
 sg13g2_buf_2 fanout4610 (.A(net4614),
    .X(net4610));
 sg13g2_buf_2 fanout4611 (.A(net4614),
    .X(net4611));
 sg13g2_buf_2 fanout4612 (.A(net4614),
    .X(net4612));
 sg13g2_buf_1 fanout4613 (.A(net4614),
    .X(net4613));
 sg13g2_buf_2 fanout4614 (.A(net4615),
    .X(net4614));
 sg13g2_buf_2 fanout4615 (.A(net4626),
    .X(net4615));
 sg13g2_buf_2 fanout4616 (.A(net4618),
    .X(net4616));
 sg13g2_buf_2 fanout4617 (.A(net4618),
    .X(net4617));
 sg13g2_buf_1 fanout4618 (.A(net4626),
    .X(net4618));
 sg13g2_buf_2 fanout4619 (.A(net4620),
    .X(net4619));
 sg13g2_buf_2 fanout4620 (.A(net4626),
    .X(net4620));
 sg13g2_buf_2 fanout4621 (.A(net4625),
    .X(net4621));
 sg13g2_buf_2 fanout4622 (.A(net4625),
    .X(net4622));
 sg13g2_buf_2 fanout4623 (.A(net4625),
    .X(net4623));
 sg13g2_buf_1 fanout4624 (.A(net4625),
    .X(net4624));
 sg13g2_buf_1 fanout4625 (.A(net4626),
    .X(net4625));
 sg13g2_buf_2 fanout4626 (.A(net4731),
    .X(net4626));
 sg13g2_buf_2 fanout4627 (.A(net4630),
    .X(net4627));
 sg13g2_buf_1 fanout4628 (.A(net4630),
    .X(net4628));
 sg13g2_buf_2 fanout4629 (.A(net4630),
    .X(net4629));
 sg13g2_buf_1 fanout4630 (.A(net4643),
    .X(net4630));
 sg13g2_buf_2 fanout4631 (.A(net4634),
    .X(net4631));
 sg13g2_buf_1 fanout4632 (.A(net4634),
    .X(net4632));
 sg13g2_buf_2 fanout4633 (.A(net4634),
    .X(net4633));
 sg13g2_buf_2 fanout4634 (.A(net4643),
    .X(net4634));
 sg13g2_buf_2 fanout4635 (.A(net4638),
    .X(net4635));
 sg13g2_buf_2 fanout4636 (.A(net4637),
    .X(net4636));
 sg13g2_buf_2 fanout4637 (.A(net4638),
    .X(net4637));
 sg13g2_buf_1 fanout4638 (.A(net4643),
    .X(net4638));
 sg13g2_buf_2 fanout4639 (.A(net4642),
    .X(net4639));
 sg13g2_buf_2 fanout4640 (.A(net4642),
    .X(net4640));
 sg13g2_buf_2 fanout4641 (.A(net4642),
    .X(net4641));
 sg13g2_buf_2 fanout4642 (.A(net4643),
    .X(net4642));
 sg13g2_buf_2 fanout4643 (.A(net4731),
    .X(net4643));
 sg13g2_buf_2 fanout4644 (.A(net4648),
    .X(net4644));
 sg13g2_buf_2 fanout4645 (.A(net4648),
    .X(net4645));
 sg13g2_buf_2 fanout4646 (.A(net4647),
    .X(net4646));
 sg13g2_buf_2 fanout4647 (.A(net4648),
    .X(net4647));
 sg13g2_buf_2 fanout4648 (.A(net4660),
    .X(net4648));
 sg13g2_buf_2 fanout4649 (.A(net4652),
    .X(net4649));
 sg13g2_buf_2 fanout4650 (.A(net4651),
    .X(net4650));
 sg13g2_buf_2 fanout4651 (.A(net4652),
    .X(net4651));
 sg13g2_buf_1 fanout4652 (.A(net4660),
    .X(net4652));
 sg13g2_buf_2 fanout4653 (.A(net4654),
    .X(net4653));
 sg13g2_buf_2 fanout4654 (.A(net4656),
    .X(net4654));
 sg13g2_buf_2 fanout4655 (.A(net4656),
    .X(net4655));
 sg13g2_buf_2 fanout4656 (.A(net4660),
    .X(net4656));
 sg13g2_buf_2 fanout4657 (.A(net4658),
    .X(net4657));
 sg13g2_buf_2 fanout4658 (.A(net4659),
    .X(net4658));
 sg13g2_buf_2 fanout4659 (.A(net4660),
    .X(net4659));
 sg13g2_buf_2 fanout4660 (.A(net4674),
    .X(net4660));
 sg13g2_buf_2 fanout4661 (.A(net4665),
    .X(net4661));
 sg13g2_buf_2 fanout4662 (.A(net4665),
    .X(net4662));
 sg13g2_buf_2 fanout4663 (.A(net4665),
    .X(net4663));
 sg13g2_buf_1 fanout4664 (.A(net4665),
    .X(net4664));
 sg13g2_buf_1 fanout4665 (.A(net4674),
    .X(net4665));
 sg13g2_buf_2 fanout4666 (.A(net4669),
    .X(net4666));
 sg13g2_buf_2 fanout4667 (.A(net4668),
    .X(net4667));
 sg13g2_buf_2 fanout4668 (.A(net4669),
    .X(net4668));
 sg13g2_buf_1 fanout4669 (.A(net4674),
    .X(net4669));
 sg13g2_buf_2 fanout4670 (.A(net4673),
    .X(net4670));
 sg13g2_buf_2 fanout4671 (.A(net4673),
    .X(net4671));
 sg13g2_buf_2 fanout4672 (.A(net4673),
    .X(net4672));
 sg13g2_buf_2 fanout4673 (.A(net4674),
    .X(net4673));
 sg13g2_buf_2 fanout4674 (.A(net4731),
    .X(net4674));
 sg13g2_buf_2 fanout4675 (.A(net4678),
    .X(net4675));
 sg13g2_buf_2 fanout4676 (.A(net4678),
    .X(net4676));
 sg13g2_buf_2 fanout4677 (.A(net4678),
    .X(net4677));
 sg13g2_buf_1 fanout4678 (.A(net4709),
    .X(net4678));
 sg13g2_buf_2 fanout4679 (.A(net4680),
    .X(net4679));
 sg13g2_buf_2 fanout4680 (.A(net4682),
    .X(net4680));
 sg13g2_buf_2 fanout4681 (.A(net4682),
    .X(net4681));
 sg13g2_buf_2 fanout4682 (.A(net4709),
    .X(net4682));
 sg13g2_buf_2 fanout4683 (.A(net4685),
    .X(net4683));
 sg13g2_buf_2 fanout4684 (.A(net4685),
    .X(net4684));
 sg13g2_buf_2 fanout4685 (.A(net4690),
    .X(net4685));
 sg13g2_buf_2 fanout4686 (.A(net4690),
    .X(net4686));
 sg13g2_buf_2 fanout4687 (.A(net4690),
    .X(net4687));
 sg13g2_buf_2 fanout4688 (.A(net4689),
    .X(net4688));
 sg13g2_buf_2 fanout4689 (.A(net4690),
    .X(net4689));
 sg13g2_buf_1 fanout4690 (.A(net4709),
    .X(net4690));
 sg13g2_buf_2 fanout4691 (.A(net4699),
    .X(net4691));
 sg13g2_buf_1 fanout4692 (.A(net4699),
    .X(net4692));
 sg13g2_buf_2 fanout4693 (.A(net4694),
    .X(net4693));
 sg13g2_buf_2 fanout4694 (.A(net4699),
    .X(net4694));
 sg13g2_buf_2 fanout4695 (.A(net4696),
    .X(net4695));
 sg13g2_buf_2 fanout4696 (.A(net4699),
    .X(net4696));
 sg13g2_buf_2 fanout4697 (.A(net4698),
    .X(net4697));
 sg13g2_buf_2 fanout4698 (.A(net4699),
    .X(net4698));
 sg13g2_buf_2 fanout4699 (.A(net4708),
    .X(net4699));
 sg13g2_buf_2 fanout4700 (.A(net4703),
    .X(net4700));
 sg13g2_buf_2 fanout4701 (.A(net4703),
    .X(net4701));
 sg13g2_buf_2 fanout4702 (.A(net4703),
    .X(net4702));
 sg13g2_buf_1 fanout4703 (.A(net4708),
    .X(net4703));
 sg13g2_buf_2 fanout4704 (.A(net4705),
    .X(net4704));
 sg13g2_buf_2 fanout4705 (.A(net4708),
    .X(net4705));
 sg13g2_buf_2 fanout4706 (.A(net4707),
    .X(net4706));
 sg13g2_buf_2 fanout4707 (.A(net4708),
    .X(net4707));
 sg13g2_buf_2 fanout4708 (.A(net4709),
    .X(net4708));
 sg13g2_buf_2 fanout4709 (.A(net4731),
    .X(net4709));
 sg13g2_buf_2 fanout4710 (.A(net4713),
    .X(net4710));
 sg13g2_buf_2 fanout4711 (.A(net4713),
    .X(net4711));
 sg13g2_buf_2 fanout4712 (.A(net4713),
    .X(net4712));
 sg13g2_buf_2 fanout4713 (.A(net4721),
    .X(net4713));
 sg13g2_buf_2 fanout4714 (.A(net4717),
    .X(net4714));
 sg13g2_buf_1 fanout4715 (.A(net4717),
    .X(net4715));
 sg13g2_buf_2 fanout4716 (.A(net4717),
    .X(net4716));
 sg13g2_buf_1 fanout4717 (.A(net4721),
    .X(net4717));
 sg13g2_buf_2 fanout4718 (.A(net4721),
    .X(net4718));
 sg13g2_buf_2 fanout4719 (.A(net4721),
    .X(net4719));
 sg13g2_buf_2 fanout4720 (.A(net4721),
    .X(net4720));
 sg13g2_buf_2 fanout4721 (.A(net4731),
    .X(net4721));
 sg13g2_buf_2 fanout4722 (.A(net4725),
    .X(net4722));
 sg13g2_buf_1 fanout4723 (.A(net4725),
    .X(net4723));
 sg13g2_buf_2 fanout4724 (.A(net4725),
    .X(net4724));
 sg13g2_buf_2 fanout4725 (.A(net4730),
    .X(net4725));
 sg13g2_buf_2 fanout4726 (.A(net4728),
    .X(net4726));
 sg13g2_buf_2 fanout4727 (.A(net4728),
    .X(net4727));
 sg13g2_buf_2 fanout4728 (.A(net4730),
    .X(net4728));
 sg13g2_buf_2 fanout4729 (.A(net4730),
    .X(net4729));
 sg13g2_buf_2 fanout4730 (.A(net4731),
    .X(net4730));
 sg13g2_buf_8 fanout4731 (.A(_04949_),
    .X(net4731));
 sg13g2_buf_2 fanout4732 (.A(net4733),
    .X(net4732));
 sg13g2_buf_2 fanout4733 (.A(net4734),
    .X(net4733));
 sg13g2_buf_1 fanout4734 (.A(net4742),
    .X(net4734));
 sg13g2_buf_2 fanout4735 (.A(net4742),
    .X(net4735));
 sg13g2_buf_1 fanout4736 (.A(net4742),
    .X(net4736));
 sg13g2_buf_2 fanout4737 (.A(net4738),
    .X(net4737));
 sg13g2_buf_2 fanout4738 (.A(net4741),
    .X(net4738));
 sg13g2_buf_2 fanout4739 (.A(net4741),
    .X(net4739));
 sg13g2_buf_2 fanout4740 (.A(net4741),
    .X(net4740));
 sg13g2_buf_2 fanout4741 (.A(net4742),
    .X(net4741));
 sg13g2_buf_2 fanout4742 (.A(_02288_),
    .X(net4742));
 sg13g2_buf_4 fanout4743 (.X(net4743),
    .A(net4745));
 sg13g2_buf_2 fanout4744 (.A(net4745),
    .X(net4744));
 sg13g2_buf_4 fanout4745 (.X(net4745),
    .A(_06878_));
 sg13g2_buf_4 fanout4746 (.X(net4746),
    .A(net4747));
 sg13g2_buf_2 fanout4747 (.A(net4748),
    .X(net4747));
 sg13g2_buf_2 fanout4748 (.A(_06877_),
    .X(net4748));
 sg13g2_buf_2 fanout4749 (.A(_05906_),
    .X(net4749));
 sg13g2_buf_1 fanout4750 (.A(_05906_),
    .X(net4750));
 sg13g2_buf_2 fanout4751 (.A(net4756),
    .X(net4751));
 sg13g2_buf_2 fanout4752 (.A(net4755),
    .X(net4752));
 sg13g2_buf_2 fanout4753 (.A(net4755),
    .X(net4753));
 sg13g2_buf_2 fanout4754 (.A(net4755),
    .X(net4754));
 sg13g2_buf_2 fanout4755 (.A(net4756),
    .X(net4755));
 sg13g2_buf_2 fanout4756 (.A(net4757),
    .X(net4756));
 sg13g2_buf_1 fanout4757 (.A(net4914),
    .X(net4757));
 sg13g2_buf_2 fanout4758 (.A(net4767),
    .X(net4758));
 sg13g2_buf_2 fanout4759 (.A(net4767),
    .X(net4759));
 sg13g2_buf_2 fanout4760 (.A(net4762),
    .X(net4760));
 sg13g2_buf_2 fanout4761 (.A(net4762),
    .X(net4761));
 sg13g2_buf_2 fanout4762 (.A(net4767),
    .X(net4762));
 sg13g2_buf_2 fanout4763 (.A(net4766),
    .X(net4763));
 sg13g2_buf_1 fanout4764 (.A(net4766),
    .X(net4764));
 sg13g2_buf_2 fanout4765 (.A(net4766),
    .X(net4765));
 sg13g2_buf_1 fanout4766 (.A(net4767),
    .X(net4766));
 sg13g2_buf_1 fanout4767 (.A(net4914),
    .X(net4767));
 sg13g2_buf_2 fanout4768 (.A(net4769),
    .X(net4768));
 sg13g2_buf_1 fanout4769 (.A(net4770),
    .X(net4769));
 sg13g2_buf_2 fanout4770 (.A(net4790),
    .X(net4770));
 sg13g2_buf_2 fanout4771 (.A(net4774),
    .X(net4771));
 sg13g2_buf_2 fanout4772 (.A(net4774),
    .X(net4772));
 sg13g2_buf_2 fanout4773 (.A(net4774),
    .X(net4773));
 sg13g2_buf_2 fanout4774 (.A(net4779),
    .X(net4774));
 sg13g2_buf_2 fanout4775 (.A(net4779),
    .X(net4775));
 sg13g2_buf_1 fanout4776 (.A(net4779),
    .X(net4776));
 sg13g2_buf_2 fanout4777 (.A(net4778),
    .X(net4777));
 sg13g2_buf_2 fanout4778 (.A(net4779),
    .X(net4778));
 sg13g2_buf_1 fanout4779 (.A(net4790),
    .X(net4779));
 sg13g2_buf_2 fanout4780 (.A(net4783),
    .X(net4780));
 sg13g2_buf_1 fanout4781 (.A(net4783),
    .X(net4781));
 sg13g2_buf_2 fanout4782 (.A(net4783),
    .X(net4782));
 sg13g2_buf_2 fanout4783 (.A(net4789),
    .X(net4783));
 sg13g2_buf_2 fanout4784 (.A(net4788),
    .X(net4784));
 sg13g2_buf_1 fanout4785 (.A(net4788),
    .X(net4785));
 sg13g2_buf_2 fanout4786 (.A(net4788),
    .X(net4786));
 sg13g2_buf_2 fanout4787 (.A(net4788),
    .X(net4787));
 sg13g2_buf_2 fanout4788 (.A(net4789),
    .X(net4788));
 sg13g2_buf_1 fanout4789 (.A(net4790),
    .X(net4789));
 sg13g2_buf_2 fanout4790 (.A(net4914),
    .X(net4790));
 sg13g2_buf_2 fanout4791 (.A(net4793),
    .X(net4791));
 sg13g2_buf_2 fanout4792 (.A(net4793),
    .X(net4792));
 sg13g2_buf_2 fanout4793 (.A(net4826),
    .X(net4793));
 sg13g2_buf_2 fanout4794 (.A(net4798),
    .X(net4794));
 sg13g2_buf_1 fanout4795 (.A(net4798),
    .X(net4795));
 sg13g2_buf_2 fanout4796 (.A(net4798),
    .X(net4796));
 sg13g2_buf_2 fanout4797 (.A(net4798),
    .X(net4797));
 sg13g2_buf_1 fanout4798 (.A(net4826),
    .X(net4798));
 sg13g2_buf_2 fanout4799 (.A(net4800),
    .X(net4799));
 sg13g2_buf_2 fanout4800 (.A(net4807),
    .X(net4800));
 sg13g2_buf_2 fanout4801 (.A(net4802),
    .X(net4801));
 sg13g2_buf_2 fanout4802 (.A(net4807),
    .X(net4802));
 sg13g2_buf_2 fanout4803 (.A(net4806),
    .X(net4803));
 sg13g2_buf_1 fanout4804 (.A(net4806),
    .X(net4804));
 sg13g2_buf_2 fanout4805 (.A(net4806),
    .X(net4805));
 sg13g2_buf_2 fanout4806 (.A(net4807),
    .X(net4806));
 sg13g2_buf_2 fanout4807 (.A(net4826),
    .X(net4807));
 sg13g2_buf_2 fanout4808 (.A(net4809),
    .X(net4808));
 sg13g2_buf_2 fanout4809 (.A(net4812),
    .X(net4809));
 sg13g2_buf_2 fanout4810 (.A(net4812),
    .X(net4810));
 sg13g2_buf_1 fanout4811 (.A(net4812),
    .X(net4811));
 sg13g2_buf_1 fanout4812 (.A(net4825),
    .X(net4812));
 sg13g2_buf_2 fanout4813 (.A(net4817),
    .X(net4813));
 sg13g2_buf_1 fanout4814 (.A(net4817),
    .X(net4814));
 sg13g2_buf_2 fanout4815 (.A(net4817),
    .X(net4815));
 sg13g2_buf_1 fanout4816 (.A(net4817),
    .X(net4816));
 sg13g2_buf_1 fanout4817 (.A(net4825),
    .X(net4817));
 sg13g2_buf_2 fanout4818 (.A(net4820),
    .X(net4818));
 sg13g2_buf_2 fanout4819 (.A(net4820),
    .X(net4819));
 sg13g2_buf_2 fanout4820 (.A(net4825),
    .X(net4820));
 sg13g2_buf_2 fanout4821 (.A(net4824),
    .X(net4821));
 sg13g2_buf_2 fanout4822 (.A(net4824),
    .X(net4822));
 sg13g2_buf_2 fanout4823 (.A(net4824),
    .X(net4823));
 sg13g2_buf_2 fanout4824 (.A(net4825),
    .X(net4824));
 sg13g2_buf_2 fanout4825 (.A(net4826),
    .X(net4825));
 sg13g2_buf_2 fanout4826 (.A(net4914),
    .X(net4826));
 sg13g2_buf_2 fanout4827 (.A(net4828),
    .X(net4827));
 sg13g2_buf_2 fanout4828 (.A(net4831),
    .X(net4828));
 sg13g2_buf_2 fanout4829 (.A(net4830),
    .X(net4829));
 sg13g2_buf_2 fanout4830 (.A(net4831),
    .X(net4830));
 sg13g2_buf_1 fanout4831 (.A(net4845),
    .X(net4831));
 sg13g2_buf_2 fanout4832 (.A(net4836),
    .X(net4832));
 sg13g2_buf_1 fanout4833 (.A(net4836),
    .X(net4833));
 sg13g2_buf_2 fanout4834 (.A(net4836),
    .X(net4834));
 sg13g2_buf_1 fanout4835 (.A(net4836),
    .X(net4835));
 sg13g2_buf_1 fanout4836 (.A(net4845),
    .X(net4836));
 sg13g2_buf_2 fanout4837 (.A(net4838),
    .X(net4837));
 sg13g2_buf_2 fanout4838 (.A(net4845),
    .X(net4838));
 sg13g2_buf_2 fanout4839 (.A(net4840),
    .X(net4839));
 sg13g2_buf_2 fanout4840 (.A(net4845),
    .X(net4840));
 sg13g2_buf_2 fanout4841 (.A(net4844),
    .X(net4841));
 sg13g2_buf_2 fanout4842 (.A(net4844),
    .X(net4842));
 sg13g2_buf_2 fanout4843 (.A(net4844),
    .X(net4843));
 sg13g2_buf_2 fanout4844 (.A(net4845),
    .X(net4844));
 sg13g2_buf_2 fanout4845 (.A(net4858),
    .X(net4845));
 sg13g2_buf_2 fanout4846 (.A(net4849),
    .X(net4846));
 sg13g2_buf_1 fanout4847 (.A(net4849),
    .X(net4847));
 sg13g2_buf_2 fanout4848 (.A(net4849),
    .X(net4848));
 sg13g2_buf_2 fanout4849 (.A(net4858),
    .X(net4849));
 sg13g2_buf_2 fanout4850 (.A(net4853),
    .X(net4850));
 sg13g2_buf_2 fanout4851 (.A(net4853),
    .X(net4851));
 sg13g2_buf_2 fanout4852 (.A(net4853),
    .X(net4852));
 sg13g2_buf_2 fanout4853 (.A(net4858),
    .X(net4853));
 sg13g2_buf_2 fanout4854 (.A(net4857),
    .X(net4854));
 sg13g2_buf_2 fanout4855 (.A(net4856),
    .X(net4855));
 sg13g2_buf_2 fanout4856 (.A(net4857),
    .X(net4856));
 sg13g2_buf_2 fanout4857 (.A(net4858),
    .X(net4857));
 sg13g2_buf_2 fanout4858 (.A(net4914),
    .X(net4858));
 sg13g2_buf_2 fanout4859 (.A(net4862),
    .X(net4859));
 sg13g2_buf_2 fanout4860 (.A(net4862),
    .X(net4860));
 sg13g2_buf_2 fanout4861 (.A(net4862),
    .X(net4861));
 sg13g2_buf_1 fanout4862 (.A(net4875),
    .X(net4862));
 sg13g2_buf_2 fanout4863 (.A(net4865),
    .X(net4863));
 sg13g2_buf_2 fanout4864 (.A(net4865),
    .X(net4864));
 sg13g2_buf_2 fanout4865 (.A(net4875),
    .X(net4865));
 sg13g2_buf_2 fanout4866 (.A(net4870),
    .X(net4866));
 sg13g2_buf_1 fanout4867 (.A(net4870),
    .X(net4867));
 sg13g2_buf_2 fanout4868 (.A(net4870),
    .X(net4868));
 sg13g2_buf_1 fanout4869 (.A(net4870),
    .X(net4869));
 sg13g2_buf_1 fanout4870 (.A(net4875),
    .X(net4870));
 sg13g2_buf_2 fanout4871 (.A(net4874),
    .X(net4871));
 sg13g2_buf_2 fanout4872 (.A(net4874),
    .X(net4872));
 sg13g2_buf_1 fanout4873 (.A(net4874),
    .X(net4873));
 sg13g2_buf_1 fanout4874 (.A(net4875),
    .X(net4874));
 sg13g2_buf_2 fanout4875 (.A(net4913),
    .X(net4875));
 sg13g2_buf_2 fanout4876 (.A(net4884),
    .X(net4876));
 sg13g2_buf_1 fanout4877 (.A(net4884),
    .X(net4877));
 sg13g2_buf_2 fanout4878 (.A(net4879),
    .X(net4878));
 sg13g2_buf_2 fanout4879 (.A(net4884),
    .X(net4879));
 sg13g2_buf_2 fanout4880 (.A(net4883),
    .X(net4880));
 sg13g2_buf_2 fanout4881 (.A(net4883),
    .X(net4881));
 sg13g2_buf_2 fanout4882 (.A(net4883),
    .X(net4882));
 sg13g2_buf_2 fanout4883 (.A(net4884),
    .X(net4883));
 sg13g2_buf_1 fanout4884 (.A(net4913),
    .X(net4884));
 sg13g2_buf_2 fanout4885 (.A(net4894),
    .X(net4885));
 sg13g2_buf_1 fanout4886 (.A(net4894),
    .X(net4886));
 sg13g2_buf_2 fanout4887 (.A(net4888),
    .X(net4887));
 sg13g2_buf_2 fanout4888 (.A(net4894),
    .X(net4888));
 sg13g2_buf_2 fanout4889 (.A(net4893),
    .X(net4889));
 sg13g2_buf_2 fanout4890 (.A(net4893),
    .X(net4890));
 sg13g2_buf_2 fanout4891 (.A(net4893),
    .X(net4891));
 sg13g2_buf_1 fanout4892 (.A(net4893),
    .X(net4892));
 sg13g2_buf_2 fanout4893 (.A(net4894),
    .X(net4893));
 sg13g2_buf_1 fanout4894 (.A(net4913),
    .X(net4894));
 sg13g2_buf_2 fanout4895 (.A(net4897),
    .X(net4895));
 sg13g2_buf_2 fanout4896 (.A(net4897),
    .X(net4896));
 sg13g2_buf_2 fanout4897 (.A(net4903),
    .X(net4897));
 sg13g2_buf_2 fanout4898 (.A(net4899),
    .X(net4898));
 sg13g2_buf_2 fanout4899 (.A(net4900),
    .X(net4899));
 sg13g2_buf_2 fanout4900 (.A(net4903),
    .X(net4900));
 sg13g2_buf_2 fanout4901 (.A(net4902),
    .X(net4901));
 sg13g2_buf_2 fanout4902 (.A(net4903),
    .X(net4902));
 sg13g2_buf_2 fanout4903 (.A(net4913),
    .X(net4903));
 sg13g2_buf_2 fanout4904 (.A(net4907),
    .X(net4904));
 sg13g2_buf_1 fanout4905 (.A(net4907),
    .X(net4905));
 sg13g2_buf_2 fanout4906 (.A(net4907),
    .X(net4906));
 sg13g2_buf_1 fanout4907 (.A(net4912),
    .X(net4907));
 sg13g2_buf_2 fanout4908 (.A(net4909),
    .X(net4908));
 sg13g2_buf_2 fanout4909 (.A(net4910),
    .X(net4909));
 sg13g2_buf_2 fanout4910 (.A(net4912),
    .X(net4910));
 sg13g2_buf_2 fanout4911 (.A(net4912),
    .X(net4911));
 sg13g2_buf_2 fanout4912 (.A(net4913),
    .X(net4912));
 sg13g2_buf_4 fanout4913 (.X(net4913),
    .A(net4914));
 sg13g2_buf_8 fanout4914 (.A(_03310_),
    .X(net4914));
 sg13g2_buf_2 fanout4915 (.A(net4916),
    .X(net4915));
 sg13g2_buf_2 fanout4916 (.A(net4924),
    .X(net4916));
 sg13g2_buf_4 fanout4917 (.X(net4917),
    .A(net4918));
 sg13g2_buf_1 fanout4918 (.A(net4924),
    .X(net4918));
 sg13g2_buf_4 fanout4919 (.X(net4919),
    .A(net4920));
 sg13g2_buf_4 fanout4920 (.X(net4920),
    .A(net4924));
 sg13g2_buf_4 fanout4921 (.X(net4921),
    .A(net4922));
 sg13g2_buf_2 fanout4922 (.A(net4923),
    .X(net4922));
 sg13g2_buf_4 fanout4923 (.X(net4923),
    .A(net4924));
 sg13g2_buf_4 fanout4924 (.X(net4924),
    .A(_02493_));
 sg13g2_buf_4 fanout4925 (.X(net4925),
    .A(net4933));
 sg13g2_buf_2 fanout4926 (.A(net4933),
    .X(net4926));
 sg13g2_buf_4 fanout4927 (.X(net4927),
    .A(net4928));
 sg13g2_buf_2 fanout4928 (.A(net4933),
    .X(net4928));
 sg13g2_buf_4 fanout4929 (.X(net4929),
    .A(net4930));
 sg13g2_buf_4 fanout4930 (.X(net4930),
    .A(net4933));
 sg13g2_buf_4 fanout4931 (.X(net4931),
    .A(net4933));
 sg13g2_buf_2 fanout4932 (.A(net4933),
    .X(net4932));
 sg13g2_buf_4 fanout4933 (.X(net4933),
    .A(_02493_));
 sg13g2_buf_8 fanout4934 (.A(_02492_),
    .X(net4934));
 sg13g2_buf_2 fanout4935 (.A(_02492_),
    .X(net4935));
 sg13g2_buf_2 fanout4936 (.A(net4938),
    .X(net4936));
 sg13g2_buf_2 fanout4937 (.A(net4938),
    .X(net4937));
 sg13g2_buf_4 fanout4938 (.X(net4938),
    .A(net4944));
 sg13g2_buf_2 fanout4939 (.A(net4944),
    .X(net4939));
 sg13g2_buf_1 fanout4940 (.A(net4944),
    .X(net4940));
 sg13g2_buf_2 fanout4941 (.A(net4943),
    .X(net4941));
 sg13g2_buf_2 fanout4942 (.A(net4943),
    .X(net4942));
 sg13g2_buf_2 fanout4943 (.A(net4944),
    .X(net4943));
 sg13g2_buf_2 fanout4944 (.A(net4952),
    .X(net4944));
 sg13g2_buf_2 fanout4945 (.A(net4946),
    .X(net4945));
 sg13g2_buf_2 fanout4946 (.A(net4947),
    .X(net4946));
 sg13g2_buf_2 fanout4947 (.A(net4952),
    .X(net4947));
 sg13g2_buf_2 fanout4948 (.A(net4949),
    .X(net4948));
 sg13g2_buf_2 fanout4949 (.A(net4952),
    .X(net4949));
 sg13g2_buf_2 fanout4950 (.A(net4951),
    .X(net4950));
 sg13g2_buf_4 fanout4951 (.X(net4951),
    .A(net4952));
 sg13g2_buf_4 fanout4952 (.X(net4952),
    .A(_02487_));
 sg13g2_buf_4 fanout4953 (.X(net4953),
    .A(_02486_));
 sg13g2_buf_2 fanout4954 (.A(_02486_),
    .X(net4954));
 sg13g2_buf_4 fanout4955 (.X(net4955),
    .A(net4956));
 sg13g2_buf_4 fanout4956 (.X(net4956),
    .A(net4957));
 sg13g2_buf_4 fanout4957 (.X(net4957),
    .A(_02486_));
 sg13g2_buf_2 fanout4958 (.A(_08888_),
    .X(net4958));
 sg13g2_buf_2 fanout4959 (.A(_08886_),
    .X(net4959));
 sg13g2_buf_4 fanout4960 (.X(net4960),
    .A(net4964));
 sg13g2_buf_2 fanout4961 (.A(net4964),
    .X(net4961));
 sg13g2_buf_4 fanout4962 (.X(net4962),
    .A(net4964));
 sg13g2_buf_2 fanout4963 (.A(net4964),
    .X(net4963));
 sg13g2_buf_2 fanout4964 (.A(_06875_),
    .X(net4964));
 sg13g2_buf_4 fanout4965 (.X(net4965),
    .A(net4967));
 sg13g2_buf_2 fanout4966 (.A(net4967),
    .X(net4966));
 sg13g2_buf_4 fanout4967 (.X(net4967),
    .A(_06875_));
 sg13g2_buf_4 fanout4968 (.X(net4968),
    .A(net4972));
 sg13g2_buf_2 fanout4969 (.A(net4972),
    .X(net4969));
 sg13g2_buf_2 fanout4970 (.A(net4972),
    .X(net4970));
 sg13g2_buf_2 fanout4971 (.A(net4972),
    .X(net4971));
 sg13g2_buf_2 fanout4972 (.A(_06875_),
    .X(net4972));
 sg13g2_buf_4 fanout4973 (.X(net4973),
    .A(net4974));
 sg13g2_buf_4 fanout4974 (.X(net4974),
    .A(_06874_));
 sg13g2_buf_4 fanout4975 (.X(net4975),
    .A(net4976));
 sg13g2_buf_2 fanout4976 (.A(net4977),
    .X(net4976));
 sg13g2_buf_2 fanout4977 (.A(_06874_),
    .X(net4977));
 sg13g2_buf_2 fanout4978 (.A(net4979),
    .X(net4978));
 sg13g2_buf_2 fanout4979 (.A(_05916_),
    .X(net4979));
 sg13g2_buf_8 fanout4980 (.A(net4981),
    .X(net4980));
 sg13g2_buf_8 fanout4981 (.A(_03085_),
    .X(net4981));
 sg13g2_buf_8 fanout4982 (.A(net4984),
    .X(net4982));
 sg13g2_buf_8 fanout4983 (.A(net4984),
    .X(net4983));
 sg13g2_buf_8 fanout4984 (.A(_03085_),
    .X(net4984));
 sg13g2_buf_2 fanout4985 (.A(_02263_),
    .X(net4985));
 sg13g2_buf_2 fanout4986 (.A(_02263_),
    .X(net4986));
 sg13g2_buf_4 fanout4987 (.X(net4987),
    .A(_02259_));
 sg13g2_buf_2 fanout4988 (.A(net4989),
    .X(net4988));
 sg13g2_buf_2 fanout4989 (.A(net4990),
    .X(net4989));
 sg13g2_buf_2 fanout4990 (.A(net4992),
    .X(net4990));
 sg13g2_buf_2 fanout4991 (.A(net4992),
    .X(net4991));
 sg13g2_buf_2 fanout4992 (.A(_02254_),
    .X(net4992));
 sg13g2_buf_2 fanout4993 (.A(net4997),
    .X(net4993));
 sg13g2_buf_2 fanout4994 (.A(net4997),
    .X(net4994));
 sg13g2_buf_2 fanout4995 (.A(net4996),
    .X(net4995));
 sg13g2_buf_2 fanout4996 (.A(net4997),
    .X(net4996));
 sg13g2_buf_2 fanout4997 (.A(_02254_),
    .X(net4997));
 sg13g2_buf_8 fanout4998 (.A(net5002),
    .X(net4998));
 sg13g2_buf_8 fanout4999 (.A(net5002),
    .X(net4999));
 sg13g2_buf_8 fanout5000 (.A(net5001),
    .X(net5000));
 sg13g2_buf_8 fanout5001 (.A(net5002),
    .X(net5001));
 sg13g2_buf_4 fanout5002 (.X(net5002),
    .A(_08873_));
 sg13g2_buf_8 fanout5003 (.A(net5007),
    .X(net5003));
 sg13g2_buf_4 fanout5004 (.X(net5004),
    .A(net5007));
 sg13g2_buf_4 fanout5005 (.X(net5005),
    .A(net5006));
 sg13g2_buf_8 fanout5006 (.A(net5007),
    .X(net5006));
 sg13g2_buf_4 fanout5007 (.X(net5007),
    .A(_08867_));
 sg13g2_buf_8 fanout5008 (.A(net5012),
    .X(net5008));
 sg13g2_buf_4 fanout5009 (.X(net5009),
    .A(net5012));
 sg13g2_buf_4 fanout5010 (.X(net5010),
    .A(net5011));
 sg13g2_buf_8 fanout5011 (.A(net5012),
    .X(net5011));
 sg13g2_buf_8 fanout5012 (.A(_08864_),
    .X(net5012));
 sg13g2_buf_4 fanout5013 (.X(net5013),
    .A(net5017));
 sg13g2_buf_4 fanout5014 (.X(net5014),
    .A(net5017));
 sg13g2_buf_4 fanout5015 (.X(net5015),
    .A(net5016));
 sg13g2_buf_4 fanout5016 (.X(net5016),
    .A(net5017));
 sg13g2_buf_4 fanout5017 (.X(net5017),
    .A(_08863_));
 sg13g2_buf_4 fanout5018 (.X(net5018),
    .A(net5019));
 sg13g2_buf_8 fanout5019 (.A(net5022),
    .X(net5019));
 sg13g2_buf_4 fanout5020 (.X(net5020),
    .A(net5022));
 sg13g2_buf_4 fanout5021 (.X(net5021),
    .A(net5022));
 sg13g2_buf_8 fanout5022 (.A(_08859_),
    .X(net5022));
 sg13g2_buf_4 fanout5023 (.X(net5023),
    .A(net5024));
 sg13g2_buf_8 fanout5024 (.A(net5027),
    .X(net5024));
 sg13g2_buf_4 fanout5025 (.X(net5025),
    .A(net5026));
 sg13g2_buf_4 fanout5026 (.X(net5026),
    .A(net5027));
 sg13g2_buf_4 fanout5027 (.X(net5027),
    .A(_08857_));
 sg13g2_buf_8 fanout5028 (.A(_08854_),
    .X(net5028));
 sg13g2_buf_4 fanout5029 (.X(net5029),
    .A(_08854_));
 sg13g2_buf_4 fanout5030 (.X(net5030),
    .A(net5032));
 sg13g2_buf_4 fanout5031 (.X(net5031),
    .A(net5032));
 sg13g2_buf_8 fanout5032 (.A(_08854_),
    .X(net5032));
 sg13g2_buf_8 fanout5033 (.A(_08830_),
    .X(net5033));
 sg13g2_buf_4 fanout5034 (.X(net5034),
    .A(_08830_));
 sg13g2_buf_4 fanout5035 (.X(net5035),
    .A(net5037));
 sg13g2_buf_8 fanout5036 (.A(net5037),
    .X(net5036));
 sg13g2_buf_8 fanout5037 (.A(_08830_),
    .X(net5037));
 sg13g2_buf_8 fanout5038 (.A(_08789_),
    .X(net5038));
 sg13g2_buf_4 fanout5039 (.X(net5039),
    .A(_08789_));
 sg13g2_buf_4 fanout5040 (.X(net5040),
    .A(net5042));
 sg13g2_buf_4 fanout5041 (.X(net5041),
    .A(net5042));
 sg13g2_buf_8 fanout5042 (.A(_08789_),
    .X(net5042));
 sg13g2_buf_4 fanout5043 (.X(net5043),
    .A(net5044));
 sg13g2_buf_8 fanout5044 (.A(net5047),
    .X(net5044));
 sg13g2_buf_8 fanout5045 (.A(net5047),
    .X(net5045));
 sg13g2_buf_4 fanout5046 (.X(net5046),
    .A(net5047));
 sg13g2_buf_8 fanout5047 (.A(_08787_),
    .X(net5047));
 sg13g2_buf_8 fanout5048 (.A(_08773_),
    .X(net5048));
 sg13g2_buf_2 fanout5049 (.A(net5050),
    .X(net5049));
 sg13g2_buf_8 fanout5050 (.A(_08773_),
    .X(net5050));
 sg13g2_buf_4 fanout5051 (.X(net5051),
    .A(net5054));
 sg13g2_buf_4 fanout5052 (.X(net5052),
    .A(net5054));
 sg13g2_buf_2 fanout5053 (.A(net5054),
    .X(net5053));
 sg13g2_buf_2 fanout5054 (.A(_08773_),
    .X(net5054));
 sg13g2_buf_4 fanout5055 (.X(net5055),
    .A(net5056));
 sg13g2_buf_8 fanout5056 (.A(net5059),
    .X(net5056));
 sg13g2_buf_8 fanout5057 (.A(net5059),
    .X(net5057));
 sg13g2_buf_4 fanout5058 (.X(net5058),
    .A(net5059));
 sg13g2_buf_8 fanout5059 (.A(_08769_),
    .X(net5059));
 sg13g2_buf_8 fanout5060 (.A(net5061),
    .X(net5060));
 sg13g2_buf_8 fanout5061 (.A(_08767_),
    .X(net5061));
 sg13g2_buf_8 fanout5062 (.A(net5064),
    .X(net5062));
 sg13g2_buf_8 fanout5063 (.A(net5064),
    .X(net5063));
 sg13g2_buf_8 fanout5064 (.A(_08767_),
    .X(net5064));
 sg13g2_buf_8 fanout5065 (.A(net5069),
    .X(net5065));
 sg13g2_buf_4 fanout5066 (.X(net5066),
    .A(net5069));
 sg13g2_buf_8 fanout5067 (.A(net5068),
    .X(net5067));
 sg13g2_buf_8 fanout5068 (.A(net5069),
    .X(net5068));
 sg13g2_buf_8 fanout5069 (.A(_06914_),
    .X(net5069));
 sg13g2_buf_8 fanout5070 (.A(net5074),
    .X(net5070));
 sg13g2_buf_8 fanout5071 (.A(net5074),
    .X(net5071));
 sg13g2_buf_8 fanout5072 (.A(net5073),
    .X(net5072));
 sg13g2_buf_8 fanout5073 (.A(net5074),
    .X(net5073));
 sg13g2_buf_8 fanout5074 (.A(_06911_),
    .X(net5074));
 sg13g2_buf_4 fanout5075 (.X(net5075),
    .A(net5076));
 sg13g2_buf_4 fanout5076 (.X(net5076),
    .A(net5078));
 sg13g2_buf_4 fanout5077 (.X(net5077),
    .A(net5078));
 sg13g2_buf_4 fanout5078 (.X(net5078),
    .A(net5083));
 sg13g2_buf_4 fanout5079 (.X(net5079),
    .A(net5083));
 sg13g2_buf_4 fanout5080 (.X(net5080),
    .A(net5083));
 sg13g2_buf_4 fanout5081 (.X(net5081),
    .A(net5082));
 sg13g2_buf_4 fanout5082 (.X(net5082),
    .A(net5083));
 sg13g2_buf_4 fanout5083 (.X(net5083),
    .A(_06888_));
 sg13g2_buf_8 fanout5084 (.A(net5088),
    .X(net5084));
 sg13g2_buf_4 fanout5085 (.X(net5085),
    .A(net5088));
 sg13g2_buf_8 fanout5086 (.A(net5087),
    .X(net5086));
 sg13g2_buf_8 fanout5087 (.A(net5088),
    .X(net5087));
 sg13g2_buf_8 fanout5088 (.A(_06886_),
    .X(net5088));
 sg13g2_buf_4 fanout5089 (.X(net5089),
    .A(net5090));
 sg13g2_buf_8 fanout5090 (.A(_06873_),
    .X(net5090));
 sg13g2_buf_2 fanout5091 (.A(net5092),
    .X(net5091));
 sg13g2_buf_2 fanout5092 (.A(net5096),
    .X(net5092));
 sg13g2_buf_2 fanout5093 (.A(net5096),
    .X(net5093));
 sg13g2_buf_2 fanout5094 (.A(net5096),
    .X(net5094));
 sg13g2_buf_2 fanout5095 (.A(net5096),
    .X(net5095));
 sg13g2_buf_2 fanout5096 (.A(net5097),
    .X(net5096));
 sg13g2_buf_8 fanout5097 (.A(_06872_),
    .X(net5097));
 sg13g2_buf_4 fanout5098 (.X(net5098),
    .A(_05985_));
 sg13g2_buf_2 fanout5099 (.A(_05985_),
    .X(net5099));
 sg13g2_buf_2 fanout5100 (.A(_04854_),
    .X(net5100));
 sg13g2_buf_2 fanout5101 (.A(_03105_),
    .X(net5101));
 sg13g2_buf_2 fanout5102 (.A(_03105_),
    .X(net5102));
 sg13g2_buf_2 fanout5103 (.A(net5105),
    .X(net5103));
 sg13g2_buf_1 fanout5104 (.A(net5105),
    .X(net5104));
 sg13g2_buf_1 fanout5105 (.A(net5106),
    .X(net5105));
 sg13g2_buf_2 fanout5106 (.A(net5107),
    .X(net5106));
 sg13g2_buf_2 fanout5107 (.A(net5108),
    .X(net5107));
 sg13g2_buf_2 fanout5108 (.A(_03093_),
    .X(net5108));
 sg13g2_buf_2 fanout5109 (.A(net5113),
    .X(net5109));
 sg13g2_buf_1 fanout5110 (.A(net5113),
    .X(net5110));
 sg13g2_buf_2 fanout5111 (.A(net5113),
    .X(net5111));
 sg13g2_buf_2 fanout5112 (.A(net5113),
    .X(net5112));
 sg13g2_buf_2 fanout5113 (.A(net5114),
    .X(net5113));
 sg13g2_buf_4 fanout5114 (.X(net5114),
    .A(_03093_));
 sg13g2_buf_8 fanout5115 (.A(_02461_),
    .X(net5115));
 sg13g2_buf_4 fanout5116 (.X(net5116),
    .A(_02461_));
 sg13g2_buf_8 fanout5117 (.A(net5119),
    .X(net5117));
 sg13g2_buf_8 fanout5118 (.A(net5119),
    .X(net5118));
 sg13g2_buf_8 fanout5119 (.A(_02461_),
    .X(net5119));
 sg13g2_buf_8 fanout5120 (.A(net5122),
    .X(net5120));
 sg13g2_buf_4 fanout5121 (.X(net5121),
    .A(net5122));
 sg13g2_buf_8 fanout5122 (.A(net5124),
    .X(net5122));
 sg13g2_buf_8 fanout5123 (.A(net5124),
    .X(net5123));
 sg13g2_buf_4 fanout5124 (.X(net5124),
    .A(_08871_));
 sg13g2_buf_8 fanout5125 (.A(net5127),
    .X(net5125));
 sg13g2_buf_4 fanout5126 (.X(net5126),
    .A(net5127));
 sg13g2_buf_4 fanout5127 (.X(net5127),
    .A(_08869_));
 sg13g2_buf_8 fanout5128 (.A(_08869_),
    .X(net5128));
 sg13g2_buf_4 fanout5129 (.X(net5129),
    .A(_08869_));
 sg13g2_buf_4 fanout5130 (.X(net5130),
    .A(net5134));
 sg13g2_buf_4 fanout5131 (.X(net5131),
    .A(net5134));
 sg13g2_buf_4 fanout5132 (.X(net5132),
    .A(net5133));
 sg13g2_buf_4 fanout5133 (.X(net5133),
    .A(net5134));
 sg13g2_buf_4 fanout5134 (.X(net5134),
    .A(_08868_));
 sg13g2_buf_4 fanout5135 (.X(net5135),
    .A(net5139));
 sg13g2_buf_8 fanout5136 (.A(net5139),
    .X(net5136));
 sg13g2_buf_4 fanout5137 (.X(net5137),
    .A(net5139));
 sg13g2_buf_4 fanout5138 (.X(net5138),
    .A(net5139));
 sg13g2_buf_4 fanout5139 (.X(net5139),
    .A(_08866_));
 sg13g2_buf_4 fanout5140 (.X(net5140),
    .A(net5141));
 sg13g2_buf_8 fanout5141 (.A(net5144),
    .X(net5141));
 sg13g2_buf_4 fanout5142 (.X(net5142),
    .A(net5143));
 sg13g2_buf_8 fanout5143 (.A(net5144),
    .X(net5143));
 sg13g2_buf_4 fanout5144 (.X(net5144),
    .A(_08862_));
 sg13g2_buf_4 fanout5145 (.X(net5145),
    .A(_08861_));
 sg13g2_buf_4 fanout5146 (.X(net5146),
    .A(_08861_));
 sg13g2_buf_4 fanout5147 (.X(net5147),
    .A(net5149));
 sg13g2_buf_8 fanout5148 (.A(net5149),
    .X(net5148));
 sg13g2_buf_4 fanout5149 (.X(net5149),
    .A(_08861_));
 sg13g2_buf_4 fanout5150 (.X(net5150),
    .A(net5154));
 sg13g2_buf_8 fanout5151 (.A(net5154),
    .X(net5151));
 sg13g2_buf_4 fanout5152 (.X(net5152),
    .A(net5154));
 sg13g2_buf_4 fanout5153 (.X(net5153),
    .A(net5154));
 sg13g2_buf_8 fanout5154 (.A(_08858_),
    .X(net5154));
 sg13g2_buf_2 fanout5155 (.A(net5158),
    .X(net5155));
 sg13g2_buf_2 fanout5156 (.A(net5158),
    .X(net5156));
 sg13g2_buf_2 fanout5157 (.A(net5158),
    .X(net5157));
 sg13g2_buf_2 fanout5158 (.A(_08835_),
    .X(net5158));
 sg13g2_buf_2 fanout5159 (.A(net5160),
    .X(net5159));
 sg13g2_buf_2 fanout5160 (.A(net5163),
    .X(net5160));
 sg13g2_buf_4 fanout5161 (.X(net5161),
    .A(net5162));
 sg13g2_buf_2 fanout5162 (.A(net5163),
    .X(net5162));
 sg13g2_buf_2 fanout5163 (.A(_08833_),
    .X(net5163));
 sg13g2_buf_8 fanout5164 (.A(_08785_),
    .X(net5164));
 sg13g2_buf_4 fanout5165 (.X(net5165),
    .A(_08785_));
 sg13g2_buf_4 fanout5166 (.X(net5166),
    .A(net5168));
 sg13g2_buf_4 fanout5167 (.X(net5167),
    .A(net5168));
 sg13g2_buf_8 fanout5168 (.A(_08785_),
    .X(net5168));
 sg13g2_buf_8 fanout5169 (.A(net5173),
    .X(net5169));
 sg13g2_buf_4 fanout5170 (.X(net5170),
    .A(net5173));
 sg13g2_buf_8 fanout5171 (.A(net5172),
    .X(net5171));
 sg13g2_buf_8 fanout5172 (.A(net5173),
    .X(net5172));
 sg13g2_buf_8 fanout5173 (.A(_08771_),
    .X(net5173));
 sg13g2_buf_4 fanout5174 (.X(net5174),
    .A(net5175));
 sg13g2_buf_4 fanout5175 (.X(net5175),
    .A(net5178));
 sg13g2_buf_4 fanout5176 (.X(net5176),
    .A(net5178));
 sg13g2_buf_4 fanout5177 (.X(net5177),
    .A(net5178));
 sg13g2_buf_2 fanout5178 (.A(_06927_),
    .X(net5178));
 sg13g2_buf_4 fanout5179 (.X(net5179),
    .A(net5180));
 sg13g2_buf_4 fanout5180 (.X(net5180),
    .A(_06920_));
 sg13g2_buf_4 fanout5181 (.X(net5181),
    .A(_06920_));
 sg13g2_buf_4 fanout5182 (.X(net5182),
    .A(net5183));
 sg13g2_buf_4 fanout5183 (.X(net5183),
    .A(_06919_));
 sg13g2_buf_4 fanout5184 (.X(net5184),
    .A(net5185));
 sg13g2_buf_4 fanout5185 (.X(net5185),
    .A(_06919_));
 sg13g2_buf_4 fanout5186 (.X(net5186),
    .A(net5188));
 sg13g2_buf_4 fanout5187 (.X(net5187),
    .A(net5188));
 sg13g2_buf_4 fanout5188 (.X(net5188),
    .A(net5192));
 sg13g2_buf_4 fanout5189 (.X(net5189),
    .A(net5191));
 sg13g2_buf_4 fanout5190 (.X(net5190),
    .A(net5191));
 sg13g2_buf_4 fanout5191 (.X(net5191),
    .A(net5192));
 sg13g2_buf_4 fanout5192 (.X(net5192),
    .A(_06919_));
 sg13g2_buf_8 fanout5193 (.A(net5194),
    .X(net5193));
 sg13g2_buf_8 fanout5194 (.A(net5197),
    .X(net5194));
 sg13g2_buf_8 fanout5195 (.A(net5196),
    .X(net5195));
 sg13g2_buf_8 fanout5196 (.A(net5197),
    .X(net5196));
 sg13g2_buf_4 fanout5197 (.X(net5197),
    .A(_06883_));
 sg13g2_buf_4 fanout5198 (.X(net5198),
    .A(_06049_));
 sg13g2_buf_4 fanout5199 (.X(net5199),
    .A(_06039_));
 sg13g2_buf_2 fanout5200 (.A(_06039_),
    .X(net5200));
 sg13g2_buf_4 fanout5201 (.X(net5201),
    .A(_05962_));
 sg13g2_buf_4 fanout5202 (.X(net5202),
    .A(net5206));
 sg13g2_buf_8 fanout5203 (.A(net5206),
    .X(net5203));
 sg13g2_buf_4 fanout5204 (.X(net5204),
    .A(net5205));
 sg13g2_buf_8 fanout5205 (.A(net5206),
    .X(net5205));
 sg13g2_buf_8 fanout5206 (.A(_04966_),
    .X(net5206));
 sg13g2_buf_4 fanout5207 (.X(net5207),
    .A(net5208));
 sg13g2_buf_4 fanout5208 (.X(net5208),
    .A(net5212));
 sg13g2_buf_4 fanout5209 (.X(net5209),
    .A(net5211));
 sg13g2_buf_4 fanout5210 (.X(net5210),
    .A(net5211));
 sg13g2_buf_8 fanout5211 (.A(net5212),
    .X(net5211));
 sg13g2_buf_4 fanout5212 (.X(net5212),
    .A(_04962_));
 sg13g2_buf_4 fanout5213 (.X(net5213),
    .A(net5214));
 sg13g2_buf_8 fanout5214 (.A(net5217),
    .X(net5214));
 sg13g2_buf_4 fanout5215 (.X(net5215),
    .A(net5216));
 sg13g2_buf_8 fanout5216 (.A(net5217),
    .X(net5216));
 sg13g2_buf_8 fanout5217 (.A(_04954_),
    .X(net5217));
 sg13g2_buf_2 fanout5218 (.A(net5219),
    .X(net5218));
 sg13g2_buf_1 fanout5219 (.A(_04896_),
    .X(net5219));
 sg13g2_buf_2 fanout5220 (.A(net5222),
    .X(net5220));
 sg13g2_buf_2 fanout5221 (.A(net5222),
    .X(net5221));
 sg13g2_buf_2 fanout5222 (.A(net5238),
    .X(net5222));
 sg13g2_buf_2 fanout5223 (.A(net5225),
    .X(net5223));
 sg13g2_buf_2 fanout5224 (.A(net5225),
    .X(net5224));
 sg13g2_buf_2 fanout5225 (.A(net5226),
    .X(net5225));
 sg13g2_buf_2 fanout5226 (.A(net5238),
    .X(net5226));
 sg13g2_buf_2 fanout5227 (.A(net5231),
    .X(net5227));
 sg13g2_buf_1 fanout5228 (.A(net5231),
    .X(net5228));
 sg13g2_buf_2 fanout5229 (.A(net5231),
    .X(net5229));
 sg13g2_buf_2 fanout5230 (.A(net5231),
    .X(net5230));
 sg13g2_buf_2 fanout5231 (.A(net5232),
    .X(net5231));
 sg13g2_buf_2 fanout5232 (.A(net5237),
    .X(net5232));
 sg13g2_buf_2 fanout5233 (.A(net5236),
    .X(net5233));
 sg13g2_buf_2 fanout5234 (.A(net5236),
    .X(net5234));
 sg13g2_buf_2 fanout5235 (.A(net5236),
    .X(net5235));
 sg13g2_buf_2 fanout5236 (.A(net5237),
    .X(net5236));
 sg13g2_buf_4 fanout5237 (.X(net5237),
    .A(net5238));
 sg13g2_buf_2 fanout5238 (.A(_04845_),
    .X(net5238));
 sg13g2_buf_2 fanout5239 (.A(net5242),
    .X(net5239));
 sg13g2_buf_1 fanout5240 (.A(net5242),
    .X(net5240));
 sg13g2_buf_2 fanout5241 (.A(net5242),
    .X(net5241));
 sg13g2_buf_2 fanout5242 (.A(net5257),
    .X(net5242));
 sg13g2_buf_2 fanout5243 (.A(net5244),
    .X(net5243));
 sg13g2_buf_2 fanout5244 (.A(net5246),
    .X(net5244));
 sg13g2_buf_2 fanout5245 (.A(net5246),
    .X(net5245));
 sg13g2_buf_2 fanout5246 (.A(net5257),
    .X(net5246));
 sg13g2_buf_2 fanout5247 (.A(net5248),
    .X(net5247));
 sg13g2_buf_2 fanout5248 (.A(net5251),
    .X(net5248));
 sg13g2_buf_4 fanout5249 (.X(net5249),
    .A(net5251));
 sg13g2_buf_2 fanout5250 (.A(net5251),
    .X(net5250));
 sg13g2_buf_2 fanout5251 (.A(net5257),
    .X(net5251));
 sg13g2_buf_2 fanout5252 (.A(net5256),
    .X(net5252));
 sg13g2_buf_1 fanout5253 (.A(net5256),
    .X(net5253));
 sg13g2_buf_2 fanout5254 (.A(net5256),
    .X(net5254));
 sg13g2_buf_2 fanout5255 (.A(net5256),
    .X(net5255));
 sg13g2_buf_2 fanout5256 (.A(net5257),
    .X(net5256));
 sg13g2_buf_2 fanout5257 (.A(net5274),
    .X(net5257));
 sg13g2_buf_2 fanout5258 (.A(net5260),
    .X(net5258));
 sg13g2_buf_2 fanout5259 (.A(net5260),
    .X(net5259));
 sg13g2_buf_1 fanout5260 (.A(net5268),
    .X(net5260));
 sg13g2_buf_2 fanout5261 (.A(net5268),
    .X(net5261));
 sg13g2_buf_2 fanout5262 (.A(net5268),
    .X(net5262));
 sg13g2_buf_2 fanout5263 (.A(net5267),
    .X(net5263));
 sg13g2_buf_1 fanout5264 (.A(net5267),
    .X(net5264));
 sg13g2_buf_2 fanout5265 (.A(net5267),
    .X(net5265));
 sg13g2_buf_2 fanout5266 (.A(net5267),
    .X(net5266));
 sg13g2_buf_1 fanout5267 (.A(net5268),
    .X(net5267));
 sg13g2_buf_2 fanout5268 (.A(net5274),
    .X(net5268));
 sg13g2_buf_2 fanout5269 (.A(net5271),
    .X(net5269));
 sg13g2_buf_2 fanout5270 (.A(net5271),
    .X(net5270));
 sg13g2_buf_2 fanout5271 (.A(net5274),
    .X(net5271));
 sg13g2_buf_2 fanout5272 (.A(net5273),
    .X(net5272));
 sg13g2_buf_2 fanout5273 (.A(net5274),
    .X(net5273));
 sg13g2_buf_4 fanout5274 (.X(net5274),
    .A(_04845_));
 sg13g2_buf_2 fanout5275 (.A(net5277),
    .X(net5275));
 sg13g2_buf_2 fanout5276 (.A(net5277),
    .X(net5276));
 sg13g2_buf_4 fanout5277 (.X(net5277),
    .A(net5282));
 sg13g2_buf_2 fanout5278 (.A(net5281),
    .X(net5278));
 sg13g2_buf_1 fanout5279 (.A(net5281),
    .X(net5279));
 sg13g2_buf_2 fanout5280 (.A(net5281),
    .X(net5280));
 sg13g2_buf_2 fanout5281 (.A(net5282),
    .X(net5281));
 sg13g2_buf_2 fanout5282 (.A(net5302),
    .X(net5282));
 sg13g2_buf_2 fanout5283 (.A(net5284),
    .X(net5283));
 sg13g2_buf_2 fanout5284 (.A(net5292),
    .X(net5284));
 sg13g2_buf_2 fanout5285 (.A(net5292),
    .X(net5285));
 sg13g2_buf_1 fanout5286 (.A(net5292),
    .X(net5286));
 sg13g2_buf_2 fanout5287 (.A(net5291),
    .X(net5287));
 sg13g2_buf_2 fanout5288 (.A(net5291),
    .X(net5288));
 sg13g2_buf_2 fanout5289 (.A(net5291),
    .X(net5289));
 sg13g2_buf_2 fanout5290 (.A(net5291),
    .X(net5290));
 sg13g2_buf_1 fanout5291 (.A(net5292),
    .X(net5291));
 sg13g2_buf_2 fanout5292 (.A(net5302),
    .X(net5292));
 sg13g2_buf_2 fanout5293 (.A(net5295),
    .X(net5293));
 sg13g2_buf_2 fanout5294 (.A(net5295),
    .X(net5294));
 sg13g2_buf_2 fanout5295 (.A(net5296),
    .X(net5295));
 sg13g2_buf_2 fanout5296 (.A(net5302),
    .X(net5296));
 sg13g2_buf_2 fanout5297 (.A(net5300),
    .X(net5297));
 sg13g2_buf_2 fanout5298 (.A(net5300),
    .X(net5298));
 sg13g2_buf_1 fanout5299 (.A(net5300),
    .X(net5299));
 sg13g2_buf_2 fanout5300 (.A(net5301),
    .X(net5300));
 sg13g2_buf_2 fanout5301 (.A(net5302),
    .X(net5301));
 sg13g2_buf_4 fanout5302 (.X(net5302),
    .A(_04845_));
 sg13g2_buf_2 fanout5303 (.A(_03101_),
    .X(net5303));
 sg13g2_buf_2 fanout5304 (.A(_03101_),
    .X(net5304));
 sg13g2_buf_2 fanout5305 (.A(net5306),
    .X(net5305));
 sg13g2_buf_2 fanout5306 (.A(net5307),
    .X(net5306));
 sg13g2_buf_2 fanout5307 (.A(net5308),
    .X(net5307));
 sg13g2_buf_2 fanout5308 (.A(net5309),
    .X(net5308));
 sg13g2_buf_2 fanout5309 (.A(net5315),
    .X(net5309));
 sg13g2_buf_4 fanout5310 (.X(net5310),
    .A(net5315));
 sg13g2_buf_2 fanout5311 (.A(net5315),
    .X(net5311));
 sg13g2_buf_2 fanout5312 (.A(net5313),
    .X(net5312));
 sg13g2_buf_2 fanout5313 (.A(net5314),
    .X(net5313));
 sg13g2_buf_2 fanout5314 (.A(net5315),
    .X(net5314));
 sg13g2_buf_4 fanout5315 (.X(net5315),
    .A(_03096_));
 sg13g2_buf_4 fanout5316 (.X(net5316),
    .A(net5319));
 sg13g2_buf_2 fanout5317 (.A(net5319),
    .X(net5317));
 sg13g2_buf_1 fanout5318 (.A(net5319),
    .X(net5318));
 sg13g2_buf_2 fanout5319 (.A(net5320),
    .X(net5319));
 sg13g2_buf_2 fanout5320 (.A(net5321),
    .X(net5320));
 sg13g2_buf_4 fanout5321 (.X(net5321),
    .A(_03094_));
 sg13g2_buf_2 fanout5322 (.A(net5326),
    .X(net5322));
 sg13g2_buf_1 fanout5323 (.A(net5326),
    .X(net5323));
 sg13g2_buf_4 fanout5324 (.X(net5324),
    .A(net5326));
 sg13g2_buf_1 fanout5325 (.A(net5326),
    .X(net5325));
 sg13g2_buf_2 fanout5326 (.A(_03094_),
    .X(net5326));
 sg13g2_buf_4 fanout5327 (.X(net5327),
    .A(_03094_));
 sg13g2_buf_2 fanout5328 (.A(net5329),
    .X(net5328));
 sg13g2_buf_2 fanout5329 (.A(net5330),
    .X(net5329));
 sg13g2_buf_2 fanout5330 (.A(net5331),
    .X(net5330));
 sg13g2_buf_1 fanout5331 (.A(net5340),
    .X(net5331));
 sg13g2_buf_2 fanout5332 (.A(net5333),
    .X(net5332));
 sg13g2_buf_4 fanout5333 (.X(net5333),
    .A(net5340));
 sg13g2_buf_2 fanout5334 (.A(net5340),
    .X(net5334));
 sg13g2_buf_1 fanout5335 (.A(net5340),
    .X(net5335));
 sg13g2_buf_2 fanout5336 (.A(net5338),
    .X(net5336));
 sg13g2_buf_1 fanout5337 (.A(net5338),
    .X(net5337));
 sg13g2_buf_2 fanout5338 (.A(net5339),
    .X(net5338));
 sg13g2_buf_2 fanout5339 (.A(net5340),
    .X(net5339));
 sg13g2_buf_4 fanout5340 (.X(net5340),
    .A(_03092_));
 sg13g2_buf_2 fanout5341 (.A(net5342),
    .X(net5341));
 sg13g2_buf_4 fanout5342 (.X(net5342),
    .A(_08834_));
 sg13g2_buf_2 fanout5343 (.A(net5344),
    .X(net5343));
 sg13g2_buf_4 fanout5344 (.X(net5344),
    .A(_08814_));
 sg13g2_buf_4 fanout5345 (.X(net5345),
    .A(net5349));
 sg13g2_buf_2 fanout5346 (.A(net5349),
    .X(net5346));
 sg13g2_buf_4 fanout5347 (.X(net5347),
    .A(net5349));
 sg13g2_buf_2 fanout5348 (.A(net5349),
    .X(net5348));
 sg13g2_buf_2 fanout5349 (.A(_06926_),
    .X(net5349));
 sg13g2_buf_4 fanout5350 (.X(net5350),
    .A(net5357));
 sg13g2_buf_4 fanout5351 (.X(net5351),
    .A(net5357));
 sg13g2_buf_4 fanout5352 (.X(net5352),
    .A(net5357));
 sg13g2_buf_4 fanout5353 (.X(net5353),
    .A(net5357));
 sg13g2_buf_2 fanout5354 (.A(net5357),
    .X(net5354));
 sg13g2_buf_4 fanout5355 (.X(net5355),
    .A(net5356));
 sg13g2_buf_4 fanout5356 (.X(net5356),
    .A(net5357));
 sg13g2_buf_4 fanout5357 (.X(net5357),
    .A(_06926_));
 sg13g2_buf_4 fanout5358 (.X(net5358),
    .A(_06050_));
 sg13g2_buf_4 fanout5359 (.X(net5359),
    .A(_05954_));
 sg13g2_buf_4 fanout5360 (.X(net5360),
    .A(net5364));
 sg13g2_buf_4 fanout5361 (.X(net5361),
    .A(net5364));
 sg13g2_buf_4 fanout5362 (.X(net5362),
    .A(net5364));
 sg13g2_buf_4 fanout5363 (.X(net5363),
    .A(net5364));
 sg13g2_buf_8 fanout5364 (.A(_04970_),
    .X(net5364));
 sg13g2_buf_4 fanout5365 (.X(net5365),
    .A(net5367));
 sg13g2_buf_2 fanout5366 (.A(net5367),
    .X(net5366));
 sg13g2_buf_4 fanout5367 (.X(net5367),
    .A(net5387));
 sg13g2_buf_4 fanout5368 (.X(net5368),
    .A(net5369));
 sg13g2_buf_2 fanout5369 (.A(net5387),
    .X(net5369));
 sg13g2_buf_4 fanout5370 (.X(net5370),
    .A(net5374));
 sg13g2_buf_4 fanout5371 (.X(net5371),
    .A(net5374));
 sg13g2_buf_4 fanout5372 (.X(net5372),
    .A(net5373));
 sg13g2_buf_2 fanout5373 (.A(net5374),
    .X(net5373));
 sg13g2_buf_4 fanout5374 (.X(net5374),
    .A(net5387));
 sg13g2_buf_4 fanout5375 (.X(net5375),
    .A(net5376));
 sg13g2_buf_4 fanout5376 (.X(net5376),
    .A(net5386));
 sg13g2_buf_4 fanout5377 (.X(net5377),
    .A(net5379));
 sg13g2_buf_4 fanout5378 (.X(net5378),
    .A(net5379));
 sg13g2_buf_4 fanout5379 (.X(net5379),
    .A(net5386));
 sg13g2_buf_4 fanout5380 (.X(net5380),
    .A(net5386));
 sg13g2_buf_2 fanout5381 (.A(net5386),
    .X(net5381));
 sg13g2_buf_4 fanout5382 (.X(net5382),
    .A(net5385));
 sg13g2_buf_4 fanout5383 (.X(net5383),
    .A(net5385));
 sg13g2_buf_2 fanout5384 (.A(net5385),
    .X(net5384));
 sg13g2_buf_2 fanout5385 (.A(net5386),
    .X(net5385));
 sg13g2_buf_4 fanout5386 (.X(net5386),
    .A(net5387));
 sg13g2_buf_4 fanout5387 (.X(net5387),
    .A(_04959_));
 sg13g2_buf_2 fanout5388 (.A(net5390),
    .X(net5388));
 sg13g2_buf_2 fanout5389 (.A(net5390),
    .X(net5389));
 sg13g2_buf_4 fanout5390 (.X(net5390),
    .A(net5392));
 sg13g2_buf_4 fanout5391 (.X(net5391),
    .A(net5392));
 sg13g2_buf_2 fanout5392 (.A(_04958_),
    .X(net5392));
 sg13g2_buf_4 fanout5393 (.X(net5393),
    .A(net5398));
 sg13g2_buf_2 fanout5394 (.A(net5398),
    .X(net5394));
 sg13g2_buf_2 fanout5395 (.A(net5398),
    .X(net5395));
 sg13g2_buf_4 fanout5396 (.X(net5396),
    .A(net5398));
 sg13g2_buf_2 fanout5397 (.A(net5398),
    .X(net5397));
 sg13g2_buf_2 fanout5398 (.A(_04958_),
    .X(net5398));
 sg13g2_buf_4 fanout5399 (.X(net5399),
    .A(net5400));
 sg13g2_buf_4 fanout5400 (.X(net5400),
    .A(net5411));
 sg13g2_buf_4 fanout5401 (.X(net5401),
    .A(net5404));
 sg13g2_buf_2 fanout5402 (.A(net5404),
    .X(net5402));
 sg13g2_buf_4 fanout5403 (.X(net5403),
    .A(net5404));
 sg13g2_buf_2 fanout5404 (.A(net5411),
    .X(net5404));
 sg13g2_buf_4 fanout5405 (.X(net5405),
    .A(net5411));
 sg13g2_buf_2 fanout5406 (.A(net5411),
    .X(net5406));
 sg13g2_buf_4 fanout5407 (.X(net5407),
    .A(net5410));
 sg13g2_buf_4 fanout5408 (.X(net5408),
    .A(net5410));
 sg13g2_buf_1 fanout5409 (.A(net5410),
    .X(net5409));
 sg13g2_buf_2 fanout5410 (.A(net5411),
    .X(net5410));
 sg13g2_buf_4 fanout5411 (.X(net5411),
    .A(_04958_));
 sg13g2_buf_4 fanout5412 (.X(net5412),
    .A(net5414));
 sg13g2_buf_2 fanout5413 (.A(net5414),
    .X(net5413));
 sg13g2_buf_4 fanout5414 (.X(net5414),
    .A(net5433));
 sg13g2_buf_4 fanout5415 (.X(net5415),
    .A(net5416));
 sg13g2_buf_2 fanout5416 (.A(net5433),
    .X(net5416));
 sg13g2_buf_4 fanout5417 (.X(net5417),
    .A(net5421));
 sg13g2_buf_4 fanout5418 (.X(net5418),
    .A(net5421));
 sg13g2_buf_4 fanout5419 (.X(net5419),
    .A(net5420));
 sg13g2_buf_2 fanout5420 (.A(net5421),
    .X(net5420));
 sg13g2_buf_4 fanout5421 (.X(net5421),
    .A(net5433));
 sg13g2_buf_4 fanout5422 (.X(net5422),
    .A(net5423));
 sg13g2_buf_4 fanout5423 (.X(net5423),
    .A(net5432));
 sg13g2_buf_4 fanout5424 (.X(net5424),
    .A(net5426));
 sg13g2_buf_4 fanout5425 (.X(net5425),
    .A(net5426));
 sg13g2_buf_4 fanout5426 (.X(net5426),
    .A(net5432));
 sg13g2_buf_4 fanout5427 (.X(net5427),
    .A(net5428));
 sg13g2_buf_4 fanout5428 (.X(net5428),
    .A(net5432));
 sg13g2_buf_4 fanout5429 (.X(net5429),
    .A(net5431));
 sg13g2_buf_4 fanout5430 (.X(net5430),
    .A(net5431));
 sg13g2_buf_4 fanout5431 (.X(net5431),
    .A(net5432));
 sg13g2_buf_2 fanout5432 (.A(net5433),
    .X(net5432));
 sg13g2_buf_4 fanout5433 (.X(net5433),
    .A(_04956_));
 sg13g2_buf_2 fanout5434 (.A(net5436),
    .X(net5434));
 sg13g2_buf_2 fanout5435 (.A(net5436),
    .X(net5435));
 sg13g2_buf_2 fanout5436 (.A(net5455),
    .X(net5436));
 sg13g2_buf_4 fanout5437 (.X(net5437),
    .A(net5438));
 sg13g2_buf_2 fanout5438 (.A(net5455),
    .X(net5438));
 sg13g2_buf_4 fanout5439 (.X(net5439),
    .A(net5443));
 sg13g2_buf_2 fanout5440 (.A(net5443),
    .X(net5440));
 sg13g2_buf_4 fanout5441 (.X(net5441),
    .A(net5442));
 sg13g2_buf_2 fanout5442 (.A(net5443),
    .X(net5442));
 sg13g2_buf_4 fanout5443 (.X(net5443),
    .A(net5455));
 sg13g2_buf_2 fanout5444 (.A(net5445),
    .X(net5444));
 sg13g2_buf_2 fanout5445 (.A(net5454),
    .X(net5445));
 sg13g2_buf_4 fanout5446 (.X(net5446),
    .A(net5448));
 sg13g2_buf_4 fanout5447 (.X(net5447),
    .A(net5448));
 sg13g2_buf_4 fanout5448 (.X(net5448),
    .A(net5454));
 sg13g2_buf_4 fanout5449 (.X(net5449),
    .A(net5450));
 sg13g2_buf_2 fanout5450 (.A(net5454),
    .X(net5450));
 sg13g2_buf_4 fanout5451 (.X(net5451),
    .A(net5453));
 sg13g2_buf_2 fanout5452 (.A(net5453),
    .X(net5452));
 sg13g2_buf_2 fanout5453 (.A(net5454),
    .X(net5453));
 sg13g2_buf_2 fanout5454 (.A(net5455),
    .X(net5454));
 sg13g2_buf_4 fanout5455 (.X(net5455),
    .A(_04955_));
 sg13g2_buf_2 fanout5456 (.A(_04852_),
    .X(net5456));
 sg13g2_buf_2 fanout5457 (.A(_04848_),
    .X(net5457));
 sg13g2_buf_2 fanout5458 (.A(_04848_),
    .X(net5458));
 sg13g2_buf_2 fanout5459 (.A(net5460),
    .X(net5459));
 sg13g2_buf_4 fanout5460 (.X(net5460),
    .A(_04342_));
 sg13g2_buf_2 fanout5461 (.A(net5463),
    .X(net5461));
 sg13g2_buf_2 fanout5462 (.A(net5463),
    .X(net5462));
 sg13g2_buf_4 fanout5463 (.X(net5463),
    .A(net5468));
 sg13g2_buf_4 fanout5464 (.X(net5464),
    .A(net5465));
 sg13g2_buf_4 fanout5465 (.X(net5465),
    .A(net5468));
 sg13g2_buf_4 fanout5466 (.X(net5466),
    .A(net5468));
 sg13g2_buf_2 fanout5467 (.A(net5468),
    .X(net5467));
 sg13g2_buf_4 fanout5468 (.X(net5468),
    .A(_04304_));
 sg13g2_buf_4 fanout5469 (.X(net5469),
    .A(net5471));
 sg13g2_buf_4 fanout5470 (.X(net5470),
    .A(net5471));
 sg13g2_buf_2 fanout5471 (.A(net5472),
    .X(net5471));
 sg13g2_buf_2 fanout5472 (.A(net5474),
    .X(net5472));
 sg13g2_buf_4 fanout5473 (.X(net5473),
    .A(net5474));
 sg13g2_buf_2 fanout5474 (.A(_04304_),
    .X(net5474));
 sg13g2_buf_2 fanout5475 (.A(net5476),
    .X(net5475));
 sg13g2_buf_2 fanout5476 (.A(net5482),
    .X(net5476));
 sg13g2_buf_2 fanout5477 (.A(net5481),
    .X(net5477));
 sg13g2_buf_4 fanout5478 (.X(net5478),
    .A(net5479));
 sg13g2_buf_2 fanout5479 (.A(net5480),
    .X(net5479));
 sg13g2_buf_2 fanout5480 (.A(net5481),
    .X(net5480));
 sg13g2_buf_2 fanout5481 (.A(net5482),
    .X(net5481));
 sg13g2_buf_2 fanout5482 (.A(_04304_),
    .X(net5482));
 sg13g2_buf_4 fanout5483 (.X(net5483),
    .A(net5485));
 sg13g2_buf_4 fanout5484 (.X(net5484),
    .A(net5485));
 sg13g2_buf_2 fanout5485 (.A(net5489),
    .X(net5485));
 sg13g2_buf_4 fanout5486 (.X(net5486),
    .A(net5488));
 sg13g2_buf_1 fanout5487 (.A(net5488),
    .X(net5487));
 sg13g2_buf_4 fanout5488 (.X(net5488),
    .A(net5489));
 sg13g2_buf_4 fanout5489 (.X(net5489),
    .A(_04279_));
 sg13g2_buf_4 fanout5490 (.X(net5490),
    .A(net5493));
 sg13g2_buf_4 fanout5491 (.X(net5491),
    .A(net5493));
 sg13g2_buf_4 fanout5492 (.X(net5492),
    .A(net5493));
 sg13g2_buf_2 fanout5493 (.A(_04279_),
    .X(net5493));
 sg13g2_buf_4 fanout5494 (.X(net5494),
    .A(net5496));
 sg13g2_buf_1 fanout5495 (.A(net5496),
    .X(net5495));
 sg13g2_buf_2 fanout5496 (.A(_04276_),
    .X(net5496));
 sg13g2_buf_4 fanout5497 (.X(net5497),
    .A(_04239_));
 sg13g2_buf_4 fanout5498 (.X(net5498),
    .A(_04238_));
 sg13g2_buf_2 fanout5499 (.A(net5500),
    .X(net5499));
 sg13g2_buf_4 fanout5500 (.X(net5500),
    .A(net5502));
 sg13g2_buf_2 fanout5501 (.A(net5502),
    .X(net5501));
 sg13g2_buf_2 fanout5502 (.A(_04237_),
    .X(net5502));
 sg13g2_buf_4 fanout5503 (.X(net5503),
    .A(net5504));
 sg13g2_buf_4 fanout5504 (.X(net5504),
    .A(_04236_));
 sg13g2_buf_2 fanout5505 (.A(net5507),
    .X(net5505));
 sg13g2_buf_1 fanout5506 (.A(net5507),
    .X(net5506));
 sg13g2_buf_2 fanout5507 (.A(_04235_),
    .X(net5507));
 sg13g2_buf_4 fanout5508 (.X(net5508),
    .A(\TRNG.chunk_index[4] ));
 sg13g2_buf_4 fanout5509 (.X(net5509),
    .A(net5511));
 sg13g2_buf_2 fanout5510 (.A(net5511),
    .X(net5510));
 sg13g2_buf_4 fanout5511 (.X(net5511),
    .A(\TRNG.chunk_index[3] ));
 sg13g2_buf_2 fanout5512 (.A(net5514),
    .X(net5512));
 sg13g2_buf_2 fanout5513 (.A(net5514),
    .X(net5513));
 sg13g2_buf_4 fanout5514 (.X(net5514),
    .A(\TRNG.chunk_index[2] ));
 sg13g2_buf_2 fanout5515 (.A(net5516),
    .X(net5515));
 sg13g2_buf_2 fanout5516 (.A(net5517),
    .X(net5516));
 sg13g2_buf_2 fanout5517 (.A(net2375),
    .X(net5517));
 sg13g2_buf_4 fanout5518 (.X(net5518),
    .A(net5522));
 sg13g2_buf_1 fanout5519 (.A(net5522),
    .X(net5519));
 sg13g2_buf_4 fanout5520 (.X(net5520),
    .A(net5521));
 sg13g2_buf_4 fanout5521 (.X(net5521),
    .A(net5522));
 sg13g2_buf_2 fanout5522 (.A(net5528),
    .X(net5522));
 sg13g2_buf_4 fanout5523 (.X(net5523),
    .A(net5528));
 sg13g2_buf_4 fanout5524 (.X(net5524),
    .A(net5528));
 sg13g2_buf_4 fanout5525 (.X(net5525),
    .A(net5526));
 sg13g2_buf_4 fanout5526 (.X(net5526),
    .A(net5528));
 sg13g2_buf_4 fanout5527 (.X(net5527),
    .A(net5528));
 sg13g2_buf_4 fanout5528 (.X(net5528),
    .A(\TRNG.Word_Valid ));
 sg13g2_buf_2 fanout5529 (.A(net5530),
    .X(net5529));
 sg13g2_buf_2 fanout5530 (.A(net5533),
    .X(net5530));
 sg13g2_buf_2 fanout5531 (.A(net5533),
    .X(net5531));
 sg13g2_buf_2 fanout5532 (.A(net5533),
    .X(net5532));
 sg13g2_buf_2 fanout5533 (.A(\TRNG.Word_Valid ),
    .X(net5533));
 sg13g2_buf_2 fanout5534 (.A(net5535),
    .X(net5534));
 sg13g2_buf_4 fanout5535 (.X(net5535),
    .A(net5542));
 sg13g2_buf_2 fanout5536 (.A(net5537),
    .X(net5536));
 sg13g2_buf_2 fanout5537 (.A(net5541),
    .X(net5537));
 sg13g2_buf_2 fanout5538 (.A(net5539),
    .X(net5538));
 sg13g2_buf_4 fanout5539 (.X(net5539),
    .A(net5540));
 sg13g2_buf_2 fanout5540 (.A(net5541),
    .X(net5540));
 sg13g2_buf_2 fanout5541 (.A(net5542),
    .X(net5541));
 sg13g2_buf_2 fanout5542 (.A(net5543),
    .X(net5542));
 sg13g2_buf_2 fanout5543 (.A(\TRNG.Word_Valid ),
    .X(net5543));
 sg13g2_buf_4 fanout5544 (.X(net5544),
    .A(\TRNG.hash[115] ));
 sg13g2_buf_4 fanout5545 (.X(net5545),
    .A(\TRNG.hash[114] ));
 sg13g2_buf_4 fanout5546 (.X(net5546),
    .A(\TRNG.hash[113] ));
 sg13g2_buf_4 fanout5547 (.X(net5547),
    .A(net3867));
 sg13g2_buf_4 fanout5548 (.X(net5548),
    .A(\TRNG.hash[108] ));
 sg13g2_buf_4 fanout5549 (.X(net5549),
    .A(\TRNG.hash[102] ));
 sg13g2_buf_4 fanout5550 (.X(net5550),
    .A(\TRNG.hash[101] ));
 sg13g2_buf_4 fanout5551 (.X(net5551),
    .A(\TRNG.hash[100] ));
 sg13g2_buf_4 fanout5552 (.X(net5552),
    .A(\TRNG.hash[99] ));
 sg13g2_buf_4 fanout5553 (.X(net5553),
    .A(\TRNG.hash[98] ));
 sg13g2_buf_4 fanout5554 (.X(net5554),
    .A(\TRNG.hash[97] ));
 sg13g2_buf_4 fanout5555 (.X(net5555),
    .A(\TRNG.hash[96] ));
 sg13g2_buf_4 fanout5556 (.X(net5556),
    .A(net3427));
 sg13g2_buf_4 fanout5557 (.X(net5557),
    .A(\TRNG.hash[253] ));
 sg13g2_buf_4 fanout5558 (.X(net5558),
    .A(\TRNG.hash[251] ));
 sg13g2_buf_4 fanout5559 (.X(net5559),
    .A(\TRNG.hash[249] ));
 sg13g2_buf_4 fanout5560 (.X(net5560),
    .A(\TRNG.hash[243] ));
 sg13g2_buf_4 fanout5561 (.X(net5561),
    .A(net3921));
 sg13g2_buf_4 fanout5562 (.X(net5562),
    .A(\TRNG.hash[238] ));
 sg13g2_buf_4 fanout5563 (.X(net5563),
    .A(\TRNG.hash[237] ));
 sg13g2_buf_4 fanout5564 (.X(net5564),
    .A(\TRNG.hash[234] ));
 sg13g2_buf_4 fanout5565 (.X(net5565),
    .A(\TRNG.hash[233] ));
 sg13g2_buf_4 fanout5566 (.X(net5566),
    .A(\TRNG.hash[230] ));
 sg13g2_buf_4 fanout5567 (.X(net5567),
    .A(\TRNG.hash[229] ));
 sg13g2_buf_4 fanout5568 (.X(net5568),
    .A(\TRNG.hash[226] ));
 sg13g2_buf_4 fanout5569 (.X(net5569),
    .A(\TRNG.hash[225] ));
 sg13g2_buf_4 fanout5570 (.X(net5570),
    .A(\TRNG.hash[224] ));
 sg13g2_buf_4 fanout5571 (.X(net5571),
    .A(net5572));
 sg13g2_buf_4 fanout5572 (.X(net5572),
    .A(net5574));
 sg13g2_buf_4 fanout5573 (.X(net5573),
    .A(net5574));
 sg13g2_buf_2 fanout5574 (.A(net3756),
    .X(net5574));
 sg13g2_buf_2 fanout5575 (.A(net3826),
    .X(net5575));
 sg13g2_buf_2 fanout5576 (.A(net5578),
    .X(net5576));
 sg13g2_buf_2 fanout5577 (.A(net5578),
    .X(net5577));
 sg13g2_buf_4 fanout5578 (.X(net5578),
    .A(net3283));
 sg13g2_buf_4 fanout5579 (.X(net5579),
    .A(net3283));
 sg13g2_buf_2 fanout5580 (.A(net5583),
    .X(net5580));
 sg13g2_buf_2 fanout5581 (.A(net5583),
    .X(net5581));
 sg13g2_buf_1 fanout5582 (.A(net5583),
    .X(net5582));
 sg13g2_buf_2 fanout5583 (.A(\TRNG.sha256.connect[4] ),
    .X(net5583));
 sg13g2_buf_2 fanout5584 (.A(net5587),
    .X(net5584));
 sg13g2_buf_2 fanout5585 (.A(net5587),
    .X(net5585));
 sg13g2_buf_1 fanout5586 (.A(net5587),
    .X(net5586));
 sg13g2_buf_1 fanout5587 (.A(\TRNG.sha256.connect[4] ),
    .X(net5587));
 sg13g2_buf_2 fanout5588 (.A(net5591),
    .X(net5588));
 sg13g2_buf_2 fanout5589 (.A(net5591),
    .X(net5589));
 sg13g2_buf_2 fanout5590 (.A(net5591),
    .X(net5590));
 sg13g2_buf_1 fanout5591 (.A(net5602),
    .X(net5591));
 sg13g2_buf_2 fanout5592 (.A(net5593),
    .X(net5592));
 sg13g2_buf_2 fanout5593 (.A(net5595),
    .X(net5593));
 sg13g2_buf_2 fanout5594 (.A(net5595),
    .X(net5594));
 sg13g2_buf_1 fanout5595 (.A(net5602),
    .X(net5595));
 sg13g2_buf_2 fanout5596 (.A(net5598),
    .X(net5596));
 sg13g2_buf_1 fanout5597 (.A(net5598),
    .X(net5597));
 sg13g2_buf_2 fanout5598 (.A(net5602),
    .X(net5598));
 sg13g2_buf_2 fanout5599 (.A(net5600),
    .X(net5599));
 sg13g2_buf_2 fanout5600 (.A(net5601),
    .X(net5600));
 sg13g2_buf_1 fanout5601 (.A(net5602),
    .X(net5601));
 sg13g2_buf_2 fanout5602 (.A(\TRNG.sha256.connect[3] ),
    .X(net5602));
 sg13g2_buf_2 fanout5603 (.A(_00130_),
    .X(net5603));
 sg13g2_buf_2 fanout5604 (.A(net5609),
    .X(net5604));
 sg13g2_buf_1 fanout5605 (.A(net5606),
    .X(net5605));
 sg13g2_buf_4 fanout5606 (.X(net5606),
    .A(net5609));
 sg13g2_buf_2 fanout5607 (.A(net5608),
    .X(net5607));
 sg13g2_buf_4 fanout5608 (.X(net5608),
    .A(net5609));
 sg13g2_buf_2 fanout5609 (.A(\TRNG.sha256.connect[2] ),
    .X(net5609));
 sg13g2_buf_4 fanout5610 (.X(net5610),
    .A(\TRNG.sha256.connect[1] ));
 sg13g2_buf_2 fanout5611 (.A(net5612),
    .X(net5611));
 sg13g2_buf_4 fanout5612 (.X(net5612),
    .A(\TRNG.sha256.connect[1] ));
 sg13g2_buf_4 fanout5613 (.X(net5613),
    .A(net5615));
 sg13g2_buf_4 fanout5614 (.X(net5614),
    .A(net5615));
 sg13g2_buf_2 fanout5615 (.A(\TRNG.sha256.connect[0] ),
    .X(net5615));
 sg13g2_buf_2 fanout5616 (.A(net5617),
    .X(net5616));
 sg13g2_buf_2 fanout5617 (.A(net3934),
    .X(net5617));
 sg13g2_buf_2 fanout5618 (.A(net5620),
    .X(net5618));
 sg13g2_buf_2 fanout5619 (.A(net5620),
    .X(net5619));
 sg13g2_buf_2 fanout5620 (.A(net3687),
    .X(net5620));
 sg13g2_buf_4 fanout5621 (.X(net5621),
    .A(net5623));
 sg13g2_buf_1 fanout5622 (.A(net5623),
    .X(net5622));
 sg13g2_buf_4 fanout5623 (.X(net5623),
    .A(net2492));
 sg13g2_buf_4 fanout5624 (.X(net5624),
    .A(net5626));
 sg13g2_buf_2 fanout5625 (.A(net5626),
    .X(net5625));
 sg13g2_buf_1 fanout5626 (.A(\TRNG.sha256.expand.data1_to_ram[28] ),
    .X(net5626));
 sg13g2_buf_2 fanout5627 (.A(net5628),
    .X(net5627));
 sg13g2_buf_2 fanout5628 (.A(net3345),
    .X(net5628));
 sg13g2_buf_2 fanout5629 (.A(\TRNG.sha256.expand.data1_to_ram[26] ),
    .X(net5629));
 sg13g2_buf_2 fanout5630 (.A(\TRNG.sha256.expand.data1_to_ram[26] ),
    .X(net5630));
 sg13g2_buf_2 fanout5631 (.A(net5632),
    .X(net5631));
 sg13g2_buf_2 fanout5632 (.A(\TRNG.sha256.expand.data1_to_ram[25] ),
    .X(net5632));
 sg13g2_buf_2 fanout5633 (.A(\TRNG.sha256.expand.data1_to_ram[24] ),
    .X(net5633));
 sg13g2_buf_2 fanout5634 (.A(\TRNG.sha256.expand.data1_to_ram[24] ),
    .X(net5634));
 sg13g2_buf_2 fanout5635 (.A(net5636),
    .X(net5635));
 sg13g2_buf_2 fanout5636 (.A(\TRNG.sha256.expand.data1_to_ram[23] ),
    .X(net5636));
 sg13g2_buf_2 fanout5637 (.A(net5638),
    .X(net5637));
 sg13g2_buf_2 fanout5638 (.A(net5639),
    .X(net5638));
 sg13g2_buf_4 fanout5639 (.X(net5639),
    .A(net3632));
 sg13g2_buf_2 fanout5640 (.A(net5641),
    .X(net5640));
 sg13g2_buf_2 fanout5641 (.A(net5642),
    .X(net5641));
 sg13g2_buf_2 fanout5642 (.A(net3720),
    .X(net5642));
 sg13g2_buf_2 fanout5643 (.A(net5645),
    .X(net5643));
 sg13g2_buf_2 fanout5644 (.A(net5645),
    .X(net5644));
 sg13g2_buf_4 fanout5645 (.X(net5645),
    .A(net2631));
 sg13g2_buf_2 fanout5646 (.A(\TRNG.sha256.expand.data1_to_ram[19] ),
    .X(net5646));
 sg13g2_buf_2 fanout5647 (.A(\TRNG.sha256.expand.data1_to_ram[19] ),
    .X(net5647));
 sg13g2_buf_2 fanout5648 (.A(net5650),
    .X(net5648));
 sg13g2_buf_1 fanout5649 (.A(net5650),
    .X(net5649));
 sg13g2_buf_2 fanout5650 (.A(net2418),
    .X(net5650));
 sg13g2_buf_2 fanout5651 (.A(net5652),
    .X(net5651));
 sg13g2_buf_2 fanout5652 (.A(\TRNG.sha256.expand.data1_to_ram[17] ),
    .X(net5652));
 sg13g2_buf_2 fanout5653 (.A(net5654),
    .X(net5653));
 sg13g2_buf_2 fanout5654 (.A(\TRNG.sha256.expand.data1_to_ram[16] ),
    .X(net5654));
 sg13g2_buf_2 fanout5655 (.A(net5657),
    .X(net5655));
 sg13g2_buf_1 fanout5656 (.A(net5657),
    .X(net5656));
 sg13g2_buf_4 fanout5657 (.X(net5657),
    .A(\TRNG.sha256.expand.data1_to_ram[15] ));
 sg13g2_buf_2 fanout5658 (.A(net5659),
    .X(net5658));
 sg13g2_buf_2 fanout5659 (.A(\TRNG.sha256.expand.data1_to_ram[14] ),
    .X(net5659));
 sg13g2_buf_2 fanout5660 (.A(\TRNG.sha256.expand.data1_to_ram[13] ),
    .X(net5660));
 sg13g2_buf_2 fanout5661 (.A(\TRNG.sha256.expand.data1_to_ram[13] ),
    .X(net5661));
 sg13g2_buf_2 fanout5662 (.A(net5664),
    .X(net5662));
 sg13g2_buf_1 fanout5663 (.A(net5664),
    .X(net5663));
 sg13g2_buf_2 fanout5664 (.A(\TRNG.sha256.expand.data1_to_ram[12] ),
    .X(net5664));
 sg13g2_buf_2 fanout5665 (.A(\TRNG.sha256.expand.data1_to_ram[11] ),
    .X(net5665));
 sg13g2_buf_2 fanout5666 (.A(\TRNG.sha256.expand.data1_to_ram[11] ),
    .X(net5666));
 sg13g2_buf_2 fanout5667 (.A(net5668),
    .X(net5667));
 sg13g2_buf_2 fanout5668 (.A(\TRNG.sha256.expand.data1_to_ram[10] ),
    .X(net5668));
 sg13g2_buf_2 fanout5669 (.A(\TRNG.sha256.expand.data1_to_ram[9] ),
    .X(net5669));
 sg13g2_buf_2 fanout5670 (.A(\TRNG.sha256.expand.data1_to_ram[9] ),
    .X(net5670));
 sg13g2_buf_4 fanout5671 (.X(net5671),
    .A(net5673));
 sg13g2_buf_2 fanout5672 (.A(net5673),
    .X(net5672));
 sg13g2_buf_4 fanout5673 (.X(net5673),
    .A(net3657));
 sg13g2_buf_2 fanout5674 (.A(net5675),
    .X(net5674));
 sg13g2_buf_2 fanout5675 (.A(\TRNG.sha256.expand.data1_to_ram[7] ),
    .X(net5675));
 sg13g2_buf_2 fanout5676 (.A(net5678),
    .X(net5676));
 sg13g2_buf_2 fanout5677 (.A(net5678),
    .X(net5677));
 sg13g2_buf_2 fanout5678 (.A(net3701),
    .X(net5678));
 sg13g2_buf_2 fanout5679 (.A(net5681),
    .X(net5679));
 sg13g2_buf_1 fanout5680 (.A(net5681),
    .X(net5680));
 sg13g2_buf_2 fanout5681 (.A(net2439),
    .X(net5681));
 sg13g2_buf_2 fanout5682 (.A(net5683),
    .X(net5682));
 sg13g2_buf_2 fanout5683 (.A(net3204),
    .X(net5683));
 sg13g2_buf_2 fanout5684 (.A(net5686),
    .X(net5684));
 sg13g2_buf_1 fanout5685 (.A(net5686),
    .X(net5685));
 sg13g2_buf_2 fanout5686 (.A(net3079),
    .X(net5686));
 sg13g2_buf_2 fanout5687 (.A(net3068),
    .X(net5687));
 sg13g2_buf_2 fanout5688 (.A(net3068),
    .X(net5688));
 sg13g2_buf_4 fanout5689 (.X(net5689),
    .A(net3063));
 sg13g2_buf_2 fanout5690 (.A(net3063),
    .X(net5690));
 sg13g2_buf_4 fanout5691 (.X(net5691),
    .A(net5692));
 sg13g2_buf_4 fanout5692 (.X(net5692),
    .A(net5701));
 sg13g2_buf_4 fanout5693 (.X(net5693),
    .A(net5694));
 sg13g2_buf_4 fanout5694 (.X(net5694),
    .A(net5701));
 sg13g2_buf_4 fanout5695 (.X(net5695),
    .A(net5701));
 sg13g2_buf_2 fanout5696 (.A(net5697),
    .X(net5696));
 sg13g2_buf_4 fanout5697 (.X(net5697),
    .A(net5701));
 sg13g2_buf_4 fanout5698 (.X(net5698),
    .A(net5700));
 sg13g2_buf_2 fanout5699 (.A(net5700),
    .X(net5699));
 sg13g2_buf_2 fanout5700 (.A(net5701),
    .X(net5700));
 sg13g2_buf_8 fanout5701 (.A(\TRNG.sha256.expand.address2[3] ),
    .X(net5701));
 sg13g2_buf_2 fanout5702 (.A(net5704),
    .X(net5702));
 sg13g2_buf_2 fanout5703 (.A(net5704),
    .X(net5703));
 sg13g2_buf_4 fanout5704 (.X(net5704),
    .A(net5711));
 sg13g2_buf_2 fanout5705 (.A(net5711),
    .X(net5705));
 sg13g2_buf_4 fanout5706 (.X(net5706),
    .A(net5710));
 sg13g2_buf_2 fanout5707 (.A(net5710),
    .X(net5707));
 sg13g2_buf_2 fanout5708 (.A(net5710),
    .X(net5708));
 sg13g2_buf_2 fanout5709 (.A(net5710),
    .X(net5709));
 sg13g2_buf_2 fanout5710 (.A(net5711),
    .X(net5710));
 sg13g2_buf_4 fanout5711 (.X(net5711),
    .A(\TRNG.sha256.expand.address2[2] ));
 sg13g2_buf_2 fanout5712 (.A(net5713),
    .X(net5712));
 sg13g2_buf_4 fanout5713 (.X(net5713),
    .A(net5725));
 sg13g2_buf_4 fanout5714 (.X(net5714),
    .A(net5717));
 sg13g2_buf_2 fanout5715 (.A(net5717),
    .X(net5715));
 sg13g2_buf_2 fanout5716 (.A(net5717),
    .X(net5716));
 sg13g2_buf_2 fanout5717 (.A(net5725),
    .X(net5717));
 sg13g2_buf_2 fanout5718 (.A(net5724),
    .X(net5718));
 sg13g2_buf_2 fanout5719 (.A(net5723),
    .X(net5719));
 sg13g2_buf_1 fanout5720 (.A(net5723),
    .X(net5720));
 sg13g2_buf_4 fanout5721 (.X(net5721),
    .A(net5723));
 sg13g2_buf_2 fanout5722 (.A(net5723),
    .X(net5722));
 sg13g2_buf_2 fanout5723 (.A(net5724),
    .X(net5723));
 sg13g2_buf_2 fanout5724 (.A(net5725),
    .X(net5724));
 sg13g2_buf_4 fanout5725 (.X(net5725),
    .A(\TRNG.sha256.expand.address2[2] ));
 sg13g2_buf_2 fanout5726 (.A(net5728),
    .X(net5726));
 sg13g2_buf_2 fanout5727 (.A(net5728),
    .X(net5727));
 sg13g2_buf_4 fanout5728 (.X(net5728),
    .A(net5729));
 sg13g2_buf_4 fanout5729 (.X(net5729),
    .A(net5733));
 sg13g2_buf_2 fanout5730 (.A(net5732),
    .X(net5730));
 sg13g2_buf_2 fanout5731 (.A(net5732),
    .X(net5731));
 sg13g2_buf_2 fanout5732 (.A(net5733),
    .X(net5732));
 sg13g2_buf_4 fanout5733 (.X(net5733),
    .A(\TRNG.sha256.expand.address2[1] ));
 sg13g2_buf_2 fanout5734 (.A(net5741),
    .X(net5734));
 sg13g2_buf_2 fanout5735 (.A(net5741),
    .X(net5735));
 sg13g2_buf_2 fanout5736 (.A(net5737),
    .X(net5736));
 sg13g2_buf_4 fanout5737 (.X(net5737),
    .A(net5741));
 sg13g2_buf_4 fanout5738 (.X(net5738),
    .A(net5740));
 sg13g2_buf_2 fanout5739 (.A(net5740),
    .X(net5739));
 sg13g2_buf_2 fanout5740 (.A(net5741),
    .X(net5740));
 sg13g2_buf_2 fanout5741 (.A(\TRNG.sha256.expand.address2[1] ),
    .X(net5741));
 sg13g2_buf_2 fanout5742 (.A(net5743),
    .X(net5742));
 sg13g2_buf_4 fanout5743 (.X(net5743),
    .A(net5744));
 sg13g2_buf_4 fanout5744 (.X(net5744),
    .A(net5751));
 sg13g2_buf_4 fanout5745 (.X(net5745),
    .A(net5750));
 sg13g2_buf_2 fanout5746 (.A(net5747),
    .X(net5746));
 sg13g2_buf_4 fanout5747 (.X(net5747),
    .A(net5750));
 sg13g2_buf_2 fanout5748 (.A(net5749),
    .X(net5748));
 sg13g2_buf_2 fanout5749 (.A(net5750),
    .X(net5749));
 sg13g2_buf_2 fanout5750 (.A(net5751),
    .X(net5750));
 sg13g2_buf_2 fanout5751 (.A(net5760),
    .X(net5751));
 sg13g2_buf_4 fanout5752 (.X(net5752),
    .A(net5753));
 sg13g2_buf_4 fanout5753 (.X(net5753),
    .A(net5760));
 sg13g2_buf_2 fanout5754 (.A(net5759),
    .X(net5754));
 sg13g2_buf_2 fanout5755 (.A(net5759),
    .X(net5755));
 sg13g2_buf_2 fanout5756 (.A(net5759),
    .X(net5756));
 sg13g2_buf_1 fanout5757 (.A(net5759),
    .X(net5757));
 sg13g2_buf_2 fanout5758 (.A(net5759),
    .X(net5758));
 sg13g2_buf_4 fanout5759 (.X(net5759),
    .A(net5760));
 sg13g2_buf_4 fanout5760 (.X(net5760),
    .A(\TRNG.sha256.expand.address2[1] ));
 sg13g2_buf_4 fanout5761 (.X(net5761),
    .A(net5762));
 sg13g2_buf_4 fanout5762 (.X(net5762),
    .A(net5765));
 sg13g2_buf_4 fanout5763 (.X(net5763),
    .A(net5765));
 sg13g2_buf_2 fanout5764 (.A(net5765),
    .X(net5764));
 sg13g2_buf_2 fanout5765 (.A(net5767),
    .X(net5765));
 sg13g2_buf_4 fanout5766 (.X(net5766),
    .A(net5767));
 sg13g2_buf_2 fanout5767 (.A(net5815),
    .X(net5767));
 sg13g2_buf_4 fanout5768 (.X(net5768),
    .A(net5771));
 sg13g2_buf_4 fanout5769 (.X(net5769),
    .A(net5771));
 sg13g2_buf_2 fanout5770 (.A(net5771),
    .X(net5770));
 sg13g2_buf_2 fanout5771 (.A(net5772),
    .X(net5771));
 sg13g2_buf_2 fanout5772 (.A(net5815),
    .X(net5772));
 sg13g2_buf_2 fanout5773 (.A(net5774),
    .X(net5773));
 sg13g2_buf_2 fanout5774 (.A(net5784),
    .X(net5774));
 sg13g2_buf_2 fanout5775 (.A(net5776),
    .X(net5775));
 sg13g2_buf_2 fanout5776 (.A(net5784),
    .X(net5776));
 sg13g2_buf_2 fanout5777 (.A(net5779),
    .X(net5777));
 sg13g2_buf_2 fanout5778 (.A(net5779),
    .X(net5778));
 sg13g2_buf_4 fanout5779 (.X(net5779),
    .A(net5784));
 sg13g2_buf_4 fanout5780 (.X(net5780),
    .A(net5781));
 sg13g2_buf_4 fanout5781 (.X(net5781),
    .A(net5784));
 sg13g2_buf_4 fanout5782 (.X(net5782),
    .A(net5783));
 sg13g2_buf_2 fanout5783 (.A(net5784),
    .X(net5783));
 sg13g2_buf_2 fanout5784 (.A(net5815),
    .X(net5784));
 sg13g2_buf_2 fanout5785 (.A(net5787),
    .X(net5785));
 sg13g2_buf_2 fanout5786 (.A(net5787),
    .X(net5786));
 sg13g2_buf_4 fanout5787 (.X(net5787),
    .A(net5790));
 sg13g2_buf_2 fanout5788 (.A(net5790),
    .X(net5788));
 sg13g2_buf_2 fanout5789 (.A(net5790),
    .X(net5789));
 sg13g2_buf_4 fanout5790 (.X(net5790),
    .A(net5800));
 sg13g2_buf_2 fanout5791 (.A(net5795),
    .X(net5791));
 sg13g2_buf_4 fanout5792 (.X(net5792),
    .A(net5794));
 sg13g2_buf_2 fanout5793 (.A(net5794),
    .X(net5793));
 sg13g2_buf_2 fanout5794 (.A(net5795),
    .X(net5794));
 sg13g2_buf_2 fanout5795 (.A(net5800),
    .X(net5795));
 sg13g2_buf_2 fanout5796 (.A(net5797),
    .X(net5796));
 sg13g2_buf_2 fanout5797 (.A(net5800),
    .X(net5797));
 sg13g2_buf_4 fanout5798 (.X(net5798),
    .A(net5799));
 sg13g2_buf_4 fanout5799 (.X(net5799),
    .A(net5800));
 sg13g2_buf_2 fanout5800 (.A(net5814),
    .X(net5800));
 sg13g2_buf_4 fanout5801 (.X(net5801),
    .A(net5804));
 sg13g2_buf_4 fanout5802 (.X(net5802),
    .A(net5803));
 sg13g2_buf_4 fanout5803 (.X(net5803),
    .A(net5804));
 sg13g2_buf_2 fanout5804 (.A(net5814),
    .X(net5804));
 sg13g2_buf_2 fanout5805 (.A(net5808),
    .X(net5805));
 sg13g2_buf_4 fanout5806 (.X(net5806),
    .A(net5808));
 sg13g2_buf_2 fanout5807 (.A(net5808),
    .X(net5807));
 sg13g2_buf_2 fanout5808 (.A(net5814),
    .X(net5808));
 sg13g2_buf_2 fanout5809 (.A(net5810),
    .X(net5809));
 sg13g2_buf_2 fanout5810 (.A(net5813),
    .X(net5810));
 sg13g2_buf_2 fanout5811 (.A(net5812),
    .X(net5811));
 sg13g2_buf_2 fanout5812 (.A(net5813),
    .X(net5812));
 sg13g2_buf_2 fanout5813 (.A(net5814),
    .X(net5813));
 sg13g2_buf_4 fanout5814 (.X(net5814),
    .A(net5815));
 sg13g2_buf_4 fanout5815 (.X(net5815),
    .A(\TRNG.sha256.expand.address2[0] ));
 sg13g2_buf_2 fanout5816 (.A(net5819),
    .X(net5816));
 sg13g2_buf_2 fanout5817 (.A(net5819),
    .X(net5817));
 sg13g2_buf_1 fanout5818 (.A(net5819),
    .X(net5818));
 sg13g2_buf_1 fanout5819 (.A(net5821),
    .X(net5819));
 sg13g2_buf_2 fanout5820 (.A(net5821),
    .X(net5820));
 sg13g2_buf_2 fanout5821 (.A(net5826),
    .X(net5821));
 sg13g2_buf_2 fanout5822 (.A(net5823),
    .X(net5822));
 sg13g2_buf_2 fanout5823 (.A(net5826),
    .X(net5823));
 sg13g2_buf_2 fanout5824 (.A(net5825),
    .X(net5824));
 sg13g2_buf_1 fanout5825 (.A(net5826),
    .X(net5825));
 sg13g2_buf_2 fanout5826 (.A(net5872),
    .X(net5826));
 sg13g2_buf_2 fanout5827 (.A(net5829),
    .X(net5827));
 sg13g2_buf_1 fanout5828 (.A(net5829),
    .X(net5828));
 sg13g2_buf_2 fanout5829 (.A(net5836),
    .X(net5829));
 sg13g2_buf_2 fanout5830 (.A(net5831),
    .X(net5830));
 sg13g2_buf_2 fanout5831 (.A(net5836),
    .X(net5831));
 sg13g2_buf_2 fanout5832 (.A(net5835),
    .X(net5832));
 sg13g2_buf_2 fanout5833 (.A(net5835),
    .X(net5833));
 sg13g2_buf_2 fanout5834 (.A(net5835),
    .X(net5834));
 sg13g2_buf_2 fanout5835 (.A(net5836),
    .X(net5835));
 sg13g2_buf_2 fanout5836 (.A(net5872),
    .X(net5836));
 sg13g2_buf_2 fanout5837 (.A(net5838),
    .X(net5837));
 sg13g2_buf_2 fanout5838 (.A(net5840),
    .X(net5838));
 sg13g2_buf_4 fanout5839 (.X(net5839),
    .A(net5840));
 sg13g2_buf_2 fanout5840 (.A(net5844),
    .X(net5840));
 sg13g2_buf_2 fanout5841 (.A(net5842),
    .X(net5841));
 sg13g2_buf_2 fanout5842 (.A(net5843),
    .X(net5842));
 sg13g2_buf_2 fanout5843 (.A(net5844),
    .X(net5843));
 sg13g2_buf_2 fanout5844 (.A(net5872),
    .X(net5844));
 sg13g2_buf_2 fanout5845 (.A(net5846),
    .X(net5845));
 sg13g2_buf_2 fanout5846 (.A(net5849),
    .X(net5846));
 sg13g2_buf_2 fanout5847 (.A(net5849),
    .X(net5847));
 sg13g2_buf_2 fanout5848 (.A(net5849),
    .X(net5848));
 sg13g2_buf_2 fanout5849 (.A(net5858),
    .X(net5849));
 sg13g2_buf_2 fanout5850 (.A(net5853),
    .X(net5850));
 sg13g2_buf_2 fanout5851 (.A(net5852),
    .X(net5851));
 sg13g2_buf_2 fanout5852 (.A(net5853),
    .X(net5852));
 sg13g2_buf_2 fanout5853 (.A(net5858),
    .X(net5853));
 sg13g2_buf_2 fanout5854 (.A(net5855),
    .X(net5854));
 sg13g2_buf_2 fanout5855 (.A(net5856),
    .X(net5855));
 sg13g2_buf_2 fanout5856 (.A(net5858),
    .X(net5856));
 sg13g2_buf_4 fanout5857 (.X(net5857),
    .A(net5858));
 sg13g2_buf_2 fanout5858 (.A(net5871),
    .X(net5858));
 sg13g2_buf_2 fanout5859 (.A(net5860),
    .X(net5859));
 sg13g2_buf_4 fanout5860 (.X(net5860),
    .A(net5866));
 sg13g2_buf_2 fanout5861 (.A(net5865),
    .X(net5861));
 sg13g2_buf_1 fanout5862 (.A(net5865),
    .X(net5862));
 sg13g2_buf_2 fanout5863 (.A(net5865),
    .X(net5863));
 sg13g2_buf_1 fanout5864 (.A(net5865),
    .X(net5864));
 sg13g2_buf_2 fanout5865 (.A(net5866),
    .X(net5865));
 sg13g2_buf_2 fanout5866 (.A(net5871),
    .X(net5866));
 sg13g2_buf_2 fanout5867 (.A(net5868),
    .X(net5867));
 sg13g2_buf_2 fanout5868 (.A(net5869),
    .X(net5868));
 sg13g2_buf_2 fanout5869 (.A(net5870),
    .X(net5869));
 sg13g2_buf_2 fanout5870 (.A(net5871),
    .X(net5870));
 sg13g2_buf_2 fanout5871 (.A(net5872),
    .X(net5871));
 sg13g2_buf_4 fanout5872 (.X(net5872),
    .A(\TRNG.sha256.compress.hash_gen.w_rdy ));
 sg13g2_buf_2 fanout5873 (.A(net3596),
    .X(net5873));
 sg13g2_buf_4 fanout5874 (.X(net5874),
    .A(net3651));
 sg13g2_buf_2 fanout5875 (.A(net5876),
    .X(net5875));
 sg13g2_buf_2 fanout5876 (.A(net3889),
    .X(net5876));
 sg13g2_buf_4 fanout5877 (.X(net5877),
    .A(net3440));
 sg13g2_buf_4 fanout5878 (.X(net5878),
    .A(net3569));
 sg13g2_buf_4 fanout5879 (.X(net5879),
    .A(net3882));
 sg13g2_buf_4 fanout5880 (.X(net5880),
    .A(net3395));
 sg13g2_buf_4 fanout5881 (.X(net5881),
    .A(\TRNG.hash[245] ));
 sg13g2_buf_4 fanout5882 (.X(net5882),
    .A(net3432));
 sg13g2_buf_4 fanout5883 (.X(net5883),
    .A(net3865));
 sg13g2_buf_4 fanout5884 (.X(net5884),
    .A(net3906));
 sg13g2_buf_4 fanout5885 (.X(net5885),
    .A(net3918));
 sg13g2_buf_4 fanout5886 (.X(net5886),
    .A(net3875));
 sg13g2_buf_4 fanout5887 (.X(net5887),
    .A(\TRNG.hash[228] ));
 sg13g2_buf_4 fanout5888 (.X(net5888),
    .A(net3736));
 sg13g2_buf_4 fanout5889 (.X(net5889),
    .A(net3892));
 sg13g2_buf_4 fanout5890 (.X(net5890),
    .A(\TRNG.hash[116] ));
 sg13g2_buf_4 fanout5891 (.X(net5891),
    .A(net3871));
 sg13g2_buf_4 fanout5892 (.X(net5892),
    .A(\TRNG.hash[111] ));
 sg13g2_buf_4 fanout5893 (.X(net5893),
    .A(net3895));
 sg13g2_buf_4 fanout5894 (.X(net5894),
    .A(net3434));
 sg13g2_buf_4 fanout5895 (.X(net5895),
    .A(\TRNG.hash[106] ));
 sg13g2_buf_4 fanout5896 (.X(net5896),
    .A(net3877));
 sg13g2_buf_4 fanout5897 (.X(net5897),
    .A(\TRNG.hash[103] ));
 sg13g2_buf_4 fanout5898 (.X(net5898),
    .A(net5899));
 sg13g2_buf_2 fanout5899 (.A(net5906),
    .X(net5899));
 sg13g2_buf_4 fanout5900 (.X(net5900),
    .A(net5905));
 sg13g2_buf_2 fanout5901 (.A(net5905),
    .X(net5901));
 sg13g2_buf_4 fanout5902 (.X(net5902),
    .A(net5904));
 sg13g2_buf_4 fanout5903 (.X(net5903),
    .A(net5904));
 sg13g2_buf_4 fanout5904 (.X(net5904),
    .A(net5905));
 sg13g2_buf_2 fanout5905 (.A(net5906),
    .X(net5905));
 sg13g2_buf_4 fanout5906 (.X(net5906),
    .A(net5931));
 sg13g2_buf_4 fanout5907 (.X(net5907),
    .A(net5909));
 sg13g2_buf_4 fanout5908 (.X(net5908),
    .A(net5909));
 sg13g2_buf_4 fanout5909 (.X(net5909),
    .A(net5910));
 sg13g2_buf_2 fanout5910 (.A(net5918),
    .X(net5910));
 sg13g2_buf_4 fanout5911 (.X(net5911),
    .A(net5918));
 sg13g2_buf_2 fanout5912 (.A(net5918),
    .X(net5912));
 sg13g2_buf_4 fanout5913 (.X(net5913),
    .A(net5917));
 sg13g2_buf_4 fanout5914 (.X(net5914),
    .A(net5917));
 sg13g2_buf_4 fanout5915 (.X(net5915),
    .A(net5917));
 sg13g2_buf_2 fanout5916 (.A(net5917),
    .X(net5916));
 sg13g2_buf_2 fanout5917 (.A(net5918),
    .X(net5917));
 sg13g2_buf_2 fanout5918 (.A(net5931),
    .X(net5918));
 sg13g2_buf_4 fanout5919 (.X(net5919),
    .A(net5925));
 sg13g2_buf_2 fanout5920 (.A(net5925),
    .X(net5920));
 sg13g2_buf_4 fanout5921 (.X(net5921),
    .A(net5922));
 sg13g2_buf_4 fanout5922 (.X(net5922),
    .A(net5925));
 sg13g2_buf_4 fanout5923 (.X(net5923),
    .A(net5924));
 sg13g2_buf_4 fanout5924 (.X(net5924),
    .A(net5925));
 sg13g2_buf_2 fanout5925 (.A(net5931),
    .X(net5925));
 sg13g2_buf_4 fanout5926 (.X(net5926),
    .A(net5930));
 sg13g2_buf_4 fanout5927 (.X(net5927),
    .A(net5930));
 sg13g2_buf_4 fanout5928 (.X(net5928),
    .A(net5929));
 sg13g2_buf_4 fanout5929 (.X(net5929),
    .A(net5930));
 sg13g2_buf_2 fanout5930 (.A(net5931),
    .X(net5930));
 sg13g2_buf_2 fanout5931 (.A(ui_in[0]),
    .X(net5931));
 sg13g2_buf_4 fanout5932 (.X(net5932),
    .A(net5934));
 sg13g2_buf_4 fanout5933 (.X(net5933),
    .A(net5934));
 sg13g2_buf_4 fanout5934 (.X(net5934),
    .A(net5968));
 sg13g2_buf_4 fanout5935 (.X(net5935),
    .A(net5939));
 sg13g2_buf_2 fanout5936 (.A(net5939),
    .X(net5936));
 sg13g2_buf_4 fanout5937 (.X(net5937),
    .A(net5939));
 sg13g2_buf_2 fanout5938 (.A(net5939),
    .X(net5938));
 sg13g2_buf_2 fanout5939 (.A(net5968),
    .X(net5939));
 sg13g2_buf_4 fanout5940 (.X(net5940),
    .A(net5948));
 sg13g2_buf_4 fanout5941 (.X(net5941),
    .A(net5948));
 sg13g2_buf_4 fanout5942 (.X(net5942),
    .A(net5943));
 sg13g2_buf_4 fanout5943 (.X(net5943),
    .A(net5948));
 sg13g2_buf_4 fanout5944 (.X(net5944),
    .A(net5945));
 sg13g2_buf_4 fanout5945 (.X(net5945),
    .A(net5948));
 sg13g2_buf_4 fanout5946 (.X(net5946),
    .A(net5948));
 sg13g2_buf_4 fanout5947 (.X(net5947),
    .A(net5948));
 sg13g2_buf_2 fanout5948 (.A(net5968),
    .X(net5948));
 sg13g2_buf_4 fanout5949 (.X(net5949),
    .A(net5950));
 sg13g2_buf_4 fanout5950 (.X(net5950),
    .A(net5958));
 sg13g2_buf_4 fanout5951 (.X(net5951),
    .A(net5958));
 sg13g2_buf_4 fanout5952 (.X(net5952),
    .A(net5958));
 sg13g2_buf_4 fanout5953 (.X(net5953),
    .A(net5957));
 sg13g2_buf_4 fanout5954 (.X(net5954),
    .A(net5957));
 sg13g2_buf_4 fanout5955 (.X(net5955),
    .A(net5957));
 sg13g2_buf_4 fanout5956 (.X(net5956),
    .A(net5957));
 sg13g2_buf_2 fanout5957 (.A(net5958),
    .X(net5957));
 sg13g2_buf_2 fanout5958 (.A(net5968),
    .X(net5958));
 sg13g2_buf_4 fanout5959 (.X(net5959),
    .A(net5962));
 sg13g2_buf_4 fanout5960 (.X(net5960),
    .A(net5962));
 sg13g2_buf_2 fanout5961 (.A(net5962),
    .X(net5961));
 sg13g2_buf_2 fanout5962 (.A(net5968),
    .X(net5962));
 sg13g2_buf_4 fanout5963 (.X(net5963),
    .A(net5967));
 sg13g2_buf_4 fanout5964 (.X(net5964),
    .A(net5967));
 sg13g2_buf_4 fanout5965 (.X(net5965),
    .A(net5967));
 sg13g2_buf_4 fanout5966 (.X(net5966),
    .A(net5967));
 sg13g2_buf_2 fanout5967 (.A(net5968),
    .X(net5967));
 sg13g2_buf_4 fanout5968 (.X(net5968),
    .A(net6066));
 sg13g2_buf_4 fanout5969 (.X(net5969),
    .A(net5973));
 sg13g2_buf_4 fanout5970 (.X(net5970),
    .A(net5973));
 sg13g2_buf_4 fanout5971 (.X(net5971),
    .A(net5973));
 sg13g2_buf_4 fanout5972 (.X(net5972),
    .A(net5973));
 sg13g2_buf_2 fanout5973 (.A(net6007),
    .X(net5973));
 sg13g2_buf_4 fanout5974 (.X(net5974),
    .A(net5978));
 sg13g2_buf_2 fanout5975 (.A(net5978),
    .X(net5975));
 sg13g2_buf_4 fanout5976 (.X(net5976),
    .A(net5977));
 sg13g2_buf_4 fanout5977 (.X(net5977),
    .A(net5978));
 sg13g2_buf_2 fanout5978 (.A(net6007),
    .X(net5978));
 sg13g2_buf_4 fanout5979 (.X(net5979),
    .A(net5980));
 sg13g2_buf_4 fanout5980 (.X(net5980),
    .A(net5988));
 sg13g2_buf_4 fanout5981 (.X(net5981),
    .A(net5988));
 sg13g2_buf_2 fanout5982 (.A(net5988),
    .X(net5982));
 sg13g2_buf_4 fanout5983 (.X(net5983),
    .A(net5987));
 sg13g2_buf_2 fanout5984 (.A(net5987),
    .X(net5984));
 sg13g2_buf_4 fanout5985 (.X(net5985),
    .A(net5987));
 sg13g2_buf_2 fanout5986 (.A(net5987),
    .X(net5986));
 sg13g2_buf_2 fanout5987 (.A(net5988),
    .X(net5987));
 sg13g2_buf_2 fanout5988 (.A(net6007),
    .X(net5988));
 sg13g2_buf_4 fanout5989 (.X(net5989),
    .A(net5992));
 sg13g2_buf_4 fanout5990 (.X(net5990),
    .A(net5992));
 sg13g2_buf_4 fanout5991 (.X(net5991),
    .A(net5992));
 sg13g2_buf_2 fanout5992 (.A(net5997),
    .X(net5992));
 sg13g2_buf_4 fanout5993 (.X(net5993),
    .A(net5994));
 sg13g2_buf_4 fanout5994 (.X(net5994),
    .A(net5997));
 sg13g2_buf_4 fanout5995 (.X(net5995),
    .A(net5996));
 sg13g2_buf_4 fanout5996 (.X(net5996),
    .A(net5997));
 sg13g2_buf_2 fanout5997 (.A(net6007),
    .X(net5997));
 sg13g2_buf_4 fanout5998 (.X(net5998),
    .A(net6001));
 sg13g2_buf_4 fanout5999 (.X(net5999),
    .A(net6001));
 sg13g2_buf_4 fanout6000 (.X(net6000),
    .A(net6001));
 sg13g2_buf_4 fanout6001 (.X(net6001),
    .A(net6007));
 sg13g2_buf_4 fanout6002 (.X(net6002),
    .A(net6006));
 sg13g2_buf_4 fanout6003 (.X(net6003),
    .A(net6006));
 sg13g2_buf_4 fanout6004 (.X(net6004),
    .A(net6006));
 sg13g2_buf_4 fanout6005 (.X(net6005),
    .A(net6006));
 sg13g2_buf_2 fanout6006 (.A(net6007),
    .X(net6006));
 sg13g2_buf_4 fanout6007 (.X(net6007),
    .A(net6066));
 sg13g2_buf_4 fanout6008 (.X(net6008),
    .A(net6017));
 sg13g2_buf_4 fanout6009 (.X(net6009),
    .A(net6017));
 sg13g2_buf_4 fanout6010 (.X(net6010),
    .A(net6011));
 sg13g2_buf_4 fanout6011 (.X(net6011),
    .A(net6017));
 sg13g2_buf_4 fanout6012 (.X(net6012),
    .A(net6013));
 sg13g2_buf_4 fanout6013 (.X(net6013),
    .A(net6016));
 sg13g2_buf_4 fanout6014 (.X(net6014),
    .A(net6016));
 sg13g2_buf_2 fanout6015 (.A(net6016),
    .X(net6015));
 sg13g2_buf_2 fanout6016 (.A(net6017),
    .X(net6016));
 sg13g2_buf_2 fanout6017 (.A(net6040),
    .X(net6017));
 sg13g2_buf_4 fanout6018 (.X(net6018),
    .A(net6020));
 sg13g2_buf_4 fanout6019 (.X(net6019),
    .A(net6020));
 sg13g2_buf_4 fanout6020 (.X(net6020),
    .A(net6025));
 sg13g2_buf_4 fanout6021 (.X(net6021),
    .A(net6022));
 sg13g2_buf_4 fanout6022 (.X(net6022),
    .A(net6025));
 sg13g2_buf_4 fanout6023 (.X(net6023),
    .A(net6025));
 sg13g2_buf_4 fanout6024 (.X(net6024),
    .A(net6025));
 sg13g2_buf_2 fanout6025 (.A(net6040),
    .X(net6025));
 sg13g2_buf_4 fanout6026 (.X(net6026),
    .A(net6030));
 sg13g2_buf_4 fanout6027 (.X(net6027),
    .A(net6030));
 sg13g2_buf_4 fanout6028 (.X(net6028),
    .A(net6030));
 sg13g2_buf_4 fanout6029 (.X(net6029),
    .A(net6030));
 sg13g2_buf_2 fanout6030 (.A(net6040),
    .X(net6030));
 sg13g2_buf_4 fanout6031 (.X(net6031),
    .A(net6034));
 sg13g2_buf_4 fanout6032 (.X(net6032),
    .A(net6034));
 sg13g2_buf_4 fanout6033 (.X(net6033),
    .A(net6034));
 sg13g2_buf_2 fanout6034 (.A(net6040),
    .X(net6034));
 sg13g2_buf_4 fanout6035 (.X(net6035),
    .A(net6036));
 sg13g2_buf_2 fanout6036 (.A(net6039),
    .X(net6036));
 sg13g2_buf_4 fanout6037 (.X(net6037),
    .A(net6039));
 sg13g2_buf_4 fanout6038 (.X(net6038),
    .A(net6039));
 sg13g2_buf_4 fanout6039 (.X(net6039),
    .A(net6040));
 sg13g2_buf_4 fanout6040 (.X(net6040),
    .A(net6066));
 sg13g2_buf_4 fanout6041 (.X(net6041),
    .A(net6042));
 sg13g2_buf_4 fanout6042 (.X(net6042),
    .A(net6059));
 sg13g2_buf_4 fanout6043 (.X(net6043),
    .A(net6044));
 sg13g2_buf_4 fanout6044 (.X(net6044),
    .A(net6059));
 sg13g2_buf_4 fanout6045 (.X(net6045),
    .A(net6049));
 sg13g2_buf_2 fanout6046 (.A(net6049),
    .X(net6046));
 sg13g2_buf_4 fanout6047 (.X(net6047),
    .A(net6049));
 sg13g2_buf_2 fanout6048 (.A(net6049),
    .X(net6048));
 sg13g2_buf_2 fanout6049 (.A(net6059),
    .X(net6049));
 sg13g2_buf_4 fanout6050 (.X(net6050),
    .A(net6054));
 sg13g2_buf_4 fanout6051 (.X(net6051),
    .A(net6054));
 sg13g2_buf_4 fanout6052 (.X(net6052),
    .A(net6054));
 sg13g2_buf_4 fanout6053 (.X(net6053),
    .A(net6054));
 sg13g2_buf_2 fanout6054 (.A(net6059),
    .X(net6054));
 sg13g2_buf_4 fanout6055 (.X(net6055),
    .A(net6058));
 sg13g2_buf_2 fanout6056 (.A(net6058),
    .X(net6056));
 sg13g2_buf_4 fanout6057 (.X(net6057),
    .A(net6058));
 sg13g2_buf_2 fanout6058 (.A(net6059),
    .X(net6058));
 sg13g2_buf_4 fanout6059 (.X(net6059),
    .A(net6065));
 sg13g2_buf_4 fanout6060 (.X(net6060),
    .A(net6063));
 sg13g2_buf_4 fanout6061 (.X(net6061),
    .A(net6063));
 sg13g2_buf_2 fanout6062 (.A(net6063),
    .X(net6062));
 sg13g2_buf_2 fanout6063 (.A(net6065),
    .X(net6063));
 sg13g2_buf_4 fanout6064 (.X(net6064),
    .A(net6065));
 sg13g2_buf_2 fanout6065 (.A(net6066),
    .X(net6065));
 sg13g2_buf_8 fanout6066 (.A(ui_in[0]),
    .X(net6066));
 sg13g2_buf_1 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_tielo tt_um_bilal_trng_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_6_3_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_6_3_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_6_0_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_6_2_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_6_0_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_6_0_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_6_0_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_6_1_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_6_0_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_6_1_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_6_1_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_6_1_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_6_6_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_6_6_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_6_7_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_6_7_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_6_7_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_6_14_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_6_14_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_6_13_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_6_24_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_6_25_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_6_25_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_6_22_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_6_7_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_6_20_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_6_22_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_6_20_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_6_16_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_6_16_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_6_16_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_6_16_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_6_17_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_6_16_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_6_17_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_6_17_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_6_18_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_6_18_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_6_21_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_6_18_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_6_18_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_6_19_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_6_19_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_6_21_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_6_19_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_6_19_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_6_21_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_6_21_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_6_20_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_6_28_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_6_28_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_6_28_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_6_29_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_6_29_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_6_28_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_6_25_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_6_31_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_6_31_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_6_31_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_6_23_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_6_23_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_6_23_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_6_20_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_6_22_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_6_22_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_6_23_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_6_27_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_6_27_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_6_27_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_6_25_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_72_clk (.A(clknet_6_24_0_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_6_26_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_74_clk (.A(clknet_6_24_0_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_2 clkbuf_leaf_75_clk (.A(clknet_6_26_0_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_2 clkbuf_leaf_76_clk (.A(clknet_6_26_0_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_2 clkbuf_leaf_77_clk (.A(clknet_6_48_0_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_2 clkbuf_leaf_78_clk (.A(clknet_6_26_0_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_2 clkbuf_leaf_79_clk (.A(clknet_6_27_0_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_2 clkbuf_leaf_80_clk (.A(clknet_6_30_0_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_2 clkbuf_leaf_81_clk (.A(clknet_6_49_0_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_2 clkbuf_leaf_82_clk (.A(clknet_6_48_0_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_2 clkbuf_leaf_83_clk (.A(clknet_6_49_0_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_2 clkbuf_leaf_84_clk (.A(clknet_6_49_0_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_2 clkbuf_leaf_85_clk (.A(clknet_6_49_0_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_2 clkbuf_leaf_86_clk (.A(clknet_6_54_0_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_2 clkbuf_leaf_87_clk (.A(clknet_6_52_0_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_2 clkbuf_leaf_88_clk (.A(clknet_6_52_0_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_2 clkbuf_leaf_89_clk (.A(clknet_6_52_0_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_2 clkbuf_leaf_90_clk (.A(clknet_6_30_0_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_2 clkbuf_leaf_91_clk (.A(clknet_6_31_0_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_2 clkbuf_leaf_92_clk (.A(clknet_6_29_0_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_2 clkbuf_leaf_93_clk (.A(clknet_6_53_0_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_2 clkbuf_leaf_94_clk (.A(clknet_6_30_0_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_2 clkbuf_leaf_95_clk (.A(clknet_6_30_0_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_2 clkbuf_leaf_96_clk (.A(clknet_6_29_0_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_2 clkbuf_leaf_97_clk (.A(clknet_6_53_0_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_2 clkbuf_leaf_98_clk (.A(clknet_6_53_0_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_2 clkbuf_leaf_99_clk (.A(clknet_6_52_0_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_2 clkbuf_leaf_100_clk (.A(clknet_6_53_0_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_2 clkbuf_leaf_101_clk (.A(clknet_6_55_0_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_2 clkbuf_leaf_102_clk (.A(clknet_6_55_0_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_2 clkbuf_leaf_103_clk (.A(clknet_6_55_0_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_2 clkbuf_leaf_104_clk (.A(clknet_6_55_0_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_2 clkbuf_leaf_105_clk (.A(clknet_6_54_0_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_2 clkbuf_leaf_106_clk (.A(clknet_6_54_0_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_2 clkbuf_leaf_107_clk (.A(clknet_6_54_0_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_2 clkbuf_leaf_108_clk (.A(clknet_6_60_0_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_2 clkbuf_leaf_109_clk (.A(clknet_6_61_0_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_2 clkbuf_leaf_110_clk (.A(clknet_6_61_0_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_2 clkbuf_leaf_111_clk (.A(clknet_6_61_0_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_2 clkbuf_leaf_112_clk (.A(clknet_6_61_0_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_2 clkbuf_leaf_113_clk (.A(clknet_6_63_0_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_2 clkbuf_leaf_114_clk (.A(clknet_6_63_0_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_2 clkbuf_leaf_115_clk (.A(clknet_6_63_0_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_2 clkbuf_leaf_116_clk (.A(clknet_6_63_0_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_2 clkbuf_leaf_117_clk (.A(clknet_6_62_0_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_2 clkbuf_leaf_118_clk (.A(clknet_6_62_0_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_2 clkbuf_leaf_119_clk (.A(clknet_6_62_0_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_2 clkbuf_leaf_120_clk (.A(clknet_6_62_0_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_2 clkbuf_leaf_121_clk (.A(clknet_6_60_0_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_2 clkbuf_leaf_122_clk (.A(clknet_6_60_0_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_2 clkbuf_leaf_123_clk (.A(clknet_6_60_0_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_2 clkbuf_leaf_124_clk (.A(clknet_6_57_0_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_2 clkbuf_leaf_125_clk (.A(clknet_6_57_0_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_2 clkbuf_leaf_126_clk (.A(clknet_6_59_0_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_2 clkbuf_leaf_127_clk (.A(clknet_6_59_0_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_2 clkbuf_leaf_128_clk (.A(clknet_6_59_0_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_2 clkbuf_leaf_129_clk (.A(clknet_6_59_0_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_2 clkbuf_leaf_130_clk (.A(clknet_6_58_0_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_2 clkbuf_leaf_131_clk (.A(clknet_6_58_0_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_2 clkbuf_leaf_132_clk (.A(clknet_6_56_0_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_2 clkbuf_leaf_133_clk (.A(clknet_6_56_0_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_2 clkbuf_leaf_134_clk (.A(clknet_6_57_0_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_2 clkbuf_leaf_135_clk (.A(clknet_6_50_0_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_2 clkbuf_leaf_136_clk (.A(clknet_6_57_0_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_2 clkbuf_leaf_137_clk (.A(clknet_6_51_0_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_2 clkbuf_leaf_138_clk (.A(clknet_6_51_0_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_2 clkbuf_leaf_139_clk (.A(clknet_6_51_0_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_2 clkbuf_leaf_140_clk (.A(clknet_6_50_0_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_2 clkbuf_leaf_141_clk (.A(clknet_6_51_0_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_2 clkbuf_leaf_142_clk (.A(clknet_6_50_0_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_2 clkbuf_leaf_143_clk (.A(clknet_6_50_0_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_2 clkbuf_leaf_144_clk (.A(clknet_6_48_0_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_2 clkbuf_leaf_145_clk (.A(clknet_6_48_0_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_2 clkbuf_leaf_146_clk (.A(clknet_6_48_0_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_2 clkbuf_leaf_147_clk (.A(clknet_6_24_0_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_2 clkbuf_leaf_148_clk (.A(clknet_6_15_0_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_2 clkbuf_leaf_149_clk (.A(clknet_6_15_0_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_2 clkbuf_leaf_150_clk (.A(clknet_6_37_0_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_2 clkbuf_leaf_151_clk (.A(clknet_6_37_0_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_2 clkbuf_leaf_152_clk (.A(clknet_6_37_0_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_2 clkbuf_leaf_153_clk (.A(clknet_6_37_0_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_2 clkbuf_leaf_154_clk (.A(clknet_6_39_0_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_2 clkbuf_leaf_155_clk (.A(clknet_6_39_0_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_2 clkbuf_leaf_156_clk (.A(clknet_6_39_0_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_2 clkbuf_leaf_157_clk (.A(clknet_6_39_0_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_2 clkbuf_leaf_158_clk (.A(clknet_6_38_0_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_2 clkbuf_leaf_159_clk (.A(clknet_6_38_0_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_2 clkbuf_leaf_160_clk (.A(clknet_6_44_0_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_2 clkbuf_leaf_161_clk (.A(clknet_6_45_0_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_2 clkbuf_leaf_162_clk (.A(clknet_6_44_0_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_2 clkbuf_leaf_163_clk (.A(clknet_6_45_0_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_2 clkbuf_leaf_164_clk (.A(clknet_6_56_0_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_2 clkbuf_leaf_165_clk (.A(clknet_6_45_0_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_2 clkbuf_leaf_166_clk (.A(clknet_6_56_0_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_2 clkbuf_leaf_167_clk (.A(clknet_6_58_0_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_2 clkbuf_leaf_168_clk (.A(clknet_6_58_0_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_2 clkbuf_leaf_169_clk (.A(clknet_6_47_0_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_2 clkbuf_leaf_170_clk (.A(clknet_6_45_0_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_2 clkbuf_leaf_171_clk (.A(clknet_6_47_0_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_2 clkbuf_leaf_172_clk (.A(clknet_6_47_0_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_2 clkbuf_leaf_173_clk (.A(clknet_6_47_0_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_2 clkbuf_leaf_174_clk (.A(clknet_6_44_0_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_2 clkbuf_leaf_175_clk (.A(clknet_6_44_0_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_2 clkbuf_leaf_176_clk (.A(clknet_6_41_0_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_2 clkbuf_leaf_177_clk (.A(clknet_6_41_0_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_2 clkbuf_leaf_178_clk (.A(clknet_6_43_0_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_2 clkbuf_leaf_179_clk (.A(clknet_6_46_0_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_2 clkbuf_leaf_180_clk (.A(clknet_6_46_0_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_2 clkbuf_leaf_181_clk (.A(clknet_6_46_0_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_2 clkbuf_leaf_182_clk (.A(clknet_6_46_0_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_2 clkbuf_leaf_183_clk (.A(clknet_6_42_0_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_2 clkbuf_leaf_184_clk (.A(clknet_6_42_0_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_2 clkbuf_leaf_185_clk (.A(clknet_6_42_0_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_2 clkbuf_leaf_186_clk (.A(clknet_6_42_0_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_2 clkbuf_leaf_187_clk (.A(clknet_6_43_0_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_2 clkbuf_leaf_188_clk (.A(clknet_6_43_0_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_2 clkbuf_leaf_189_clk (.A(clknet_6_40_0_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_2 clkbuf_leaf_190_clk (.A(clknet_6_40_0_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_2 clkbuf_leaf_191_clk (.A(clknet_6_40_0_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_2 clkbuf_leaf_192_clk (.A(clknet_6_43_0_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_2 clkbuf_leaf_193_clk (.A(clknet_6_41_0_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_2 clkbuf_leaf_194_clk (.A(clknet_6_41_0_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_2 clkbuf_leaf_195_clk (.A(clknet_6_35_0_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_2 clkbuf_leaf_196_clk (.A(clknet_6_35_0_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_2 clkbuf_leaf_197_clk (.A(clknet_6_34_0_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_2 clkbuf_leaf_198_clk (.A(clknet_6_40_0_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_2 clkbuf_leaf_199_clk (.A(clknet_6_34_0_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_2 clkbuf_leaf_200_clk (.A(clknet_6_34_0_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_2 clkbuf_leaf_201_clk (.A(clknet_6_34_0_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_2 clkbuf_leaf_202_clk (.A(clknet_6_32_0_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_2 clkbuf_leaf_203_clk (.A(clknet_6_32_0_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_2 clkbuf_leaf_204_clk (.A(clknet_6_32_0_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_2 clkbuf_leaf_205_clk (.A(clknet_6_10_0_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_2 clkbuf_leaf_206_clk (.A(clknet_6_8_0_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_2 clkbuf_leaf_207_clk (.A(clknet_6_32_0_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_2 clkbuf_leaf_208_clk (.A(clknet_6_32_0_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_2 clkbuf_leaf_209_clk (.A(clknet_6_10_0_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_2 clkbuf_leaf_210_clk (.A(clknet_6_11_0_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_2 clkbuf_leaf_211_clk (.A(clknet_6_10_0_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_2 clkbuf_leaf_212_clk (.A(clknet_6_33_0_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_2 clkbuf_leaf_213_clk (.A(clknet_6_33_0_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_2 clkbuf_leaf_214_clk (.A(clknet_6_33_0_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_2 clkbuf_leaf_215_clk (.A(clknet_6_35_0_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_2 clkbuf_leaf_216_clk (.A(clknet_6_35_0_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_2 clkbuf_leaf_217_clk (.A(clknet_6_38_0_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_2 clkbuf_leaf_218_clk (.A(clknet_6_38_0_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_2 clkbuf_leaf_219_clk (.A(clknet_6_36_0_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_2 clkbuf_leaf_220_clk (.A(clknet_6_36_0_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_2 clkbuf_leaf_221_clk (.A(clknet_6_33_0_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_2 clkbuf_leaf_222_clk (.A(clknet_6_11_0_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_2 clkbuf_leaf_223_clk (.A(clknet_6_11_0_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_2 clkbuf_leaf_224_clk (.A(clknet_6_13_0_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_2 clkbuf_leaf_225_clk (.A(clknet_6_36_0_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_2 clkbuf_leaf_226_clk (.A(clknet_6_36_0_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_2 clkbuf_leaf_227_clk (.A(clknet_6_15_0_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_2 clkbuf_leaf_228_clk (.A(clknet_6_15_0_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_2 clkbuf_leaf_229_clk (.A(clknet_6_14_0_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_2 clkbuf_leaf_230_clk (.A(clknet_6_13_0_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_2 clkbuf_leaf_231_clk (.A(clknet_6_14_0_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_2 clkbuf_leaf_232_clk (.A(clknet_6_12_0_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_2 clkbuf_leaf_233_clk (.A(clknet_6_13_0_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_2 clkbuf_leaf_234_clk (.A(clknet_6_12_0_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_2 clkbuf_leaf_235_clk (.A(clknet_6_12_0_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_2 clkbuf_leaf_236_clk (.A(clknet_6_5_0_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_2 clkbuf_leaf_237_clk (.A(clknet_6_6_0_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_2 clkbuf_leaf_238_clk (.A(clknet_6_5_0_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_2 clkbuf_leaf_239_clk (.A(clknet_6_6_0_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_2 clkbuf_leaf_240_clk (.A(clknet_6_5_0_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_2 clkbuf_leaf_241_clk (.A(clknet_6_5_0_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_2 clkbuf_leaf_242_clk (.A(clknet_6_4_0_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_2 clkbuf_leaf_243_clk (.A(clknet_6_4_0_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_2 clkbuf_leaf_244_clk (.A(clknet_6_11_0_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_2 clkbuf_leaf_245_clk (.A(clknet_6_10_0_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_2 clkbuf_leaf_246_clk (.A(clknet_6_8_0_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_2 clkbuf_leaf_247_clk (.A(clknet_6_12_0_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_2 clkbuf_leaf_248_clk (.A(clknet_6_8_0_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_2 clkbuf_leaf_249_clk (.A(clknet_6_9_0_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_2 clkbuf_leaf_250_clk (.A(clknet_6_9_0_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_2 clkbuf_leaf_251_clk (.A(clknet_6_8_0_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_2 clkbuf_leaf_252_clk (.A(clknet_6_9_0_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_2 clkbuf_leaf_253_clk (.A(clknet_6_9_0_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_2 clkbuf_leaf_254_clk (.A(clknet_6_4_0_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_2 clkbuf_leaf_255_clk (.A(clknet_6_4_0_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_2 clkbuf_leaf_256_clk (.A(clknet_6_2_0_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_2 clkbuf_leaf_257_clk (.A(clknet_6_2_0_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_2 clkbuf_leaf_258_clk (.A(clknet_6_2_0_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_2 clkbuf_leaf_259_clk (.A(clknet_6_3_0_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_2 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_2 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_2 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_2 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_2 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_2 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_2 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_2 clkbuf_6_0_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_0_0_clk));
 sg13g2_buf_2 clkbuf_6_1_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_1_0_clk));
 sg13g2_buf_2 clkbuf_6_2_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_2_0_clk));
 sg13g2_buf_2 clkbuf_6_3_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_3_0_clk));
 sg13g2_buf_2 clkbuf_6_4_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_4_0_clk));
 sg13g2_buf_2 clkbuf_6_5_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_5_0_clk));
 sg13g2_buf_2 clkbuf_6_6_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_6_0_clk));
 sg13g2_buf_2 clkbuf_6_7_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_7_0_clk));
 sg13g2_buf_2 clkbuf_6_8_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_8_0_clk));
 sg13g2_buf_2 clkbuf_6_9_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_9_0_clk));
 sg13g2_buf_2 clkbuf_6_10_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_10_0_clk));
 sg13g2_buf_2 clkbuf_6_11_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_11_0_clk));
 sg13g2_buf_2 clkbuf_6_12_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_12_0_clk));
 sg13g2_buf_2 clkbuf_6_13_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_13_0_clk));
 sg13g2_buf_2 clkbuf_6_14_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_14_0_clk));
 sg13g2_buf_2 clkbuf_6_15_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_15_0_clk));
 sg13g2_buf_2 clkbuf_6_16_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_16_0_clk));
 sg13g2_buf_2 clkbuf_6_17_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_17_0_clk));
 sg13g2_buf_2 clkbuf_6_18_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_18_0_clk));
 sg13g2_buf_2 clkbuf_6_19_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_19_0_clk));
 sg13g2_buf_2 clkbuf_6_20_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_20_0_clk));
 sg13g2_buf_2 clkbuf_6_21_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_21_0_clk));
 sg13g2_buf_2 clkbuf_6_22_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_22_0_clk));
 sg13g2_buf_2 clkbuf_6_23_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_23_0_clk));
 sg13g2_buf_2 clkbuf_6_24_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_24_0_clk));
 sg13g2_buf_2 clkbuf_6_25_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_25_0_clk));
 sg13g2_buf_2 clkbuf_6_26_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_26_0_clk));
 sg13g2_buf_2 clkbuf_6_27_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_27_0_clk));
 sg13g2_buf_2 clkbuf_6_28_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_28_0_clk));
 sg13g2_buf_2 clkbuf_6_29_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_29_0_clk));
 sg13g2_buf_2 clkbuf_6_30_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_30_0_clk));
 sg13g2_buf_2 clkbuf_6_31_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_31_0_clk));
 sg13g2_buf_2 clkbuf_6_32_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_32_0_clk));
 sg13g2_buf_2 clkbuf_6_33_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_33_0_clk));
 sg13g2_buf_2 clkbuf_6_34_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_34_0_clk));
 sg13g2_buf_2 clkbuf_6_35_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_35_0_clk));
 sg13g2_buf_2 clkbuf_6_36_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_36_0_clk));
 sg13g2_buf_2 clkbuf_6_37_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_37_0_clk));
 sg13g2_buf_2 clkbuf_6_38_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_38_0_clk));
 sg13g2_buf_2 clkbuf_6_39_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_39_0_clk));
 sg13g2_buf_2 clkbuf_6_40_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_40_0_clk));
 sg13g2_buf_2 clkbuf_6_41_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_41_0_clk));
 sg13g2_buf_2 clkbuf_6_42_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_42_0_clk));
 sg13g2_buf_2 clkbuf_6_43_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_43_0_clk));
 sg13g2_buf_2 clkbuf_6_44_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_44_0_clk));
 sg13g2_buf_2 clkbuf_6_45_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_45_0_clk));
 sg13g2_buf_2 clkbuf_6_46_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_46_0_clk));
 sg13g2_buf_2 clkbuf_6_47_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_47_0_clk));
 sg13g2_buf_2 clkbuf_6_48_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_48_0_clk));
 sg13g2_buf_2 clkbuf_6_49_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_49_0_clk));
 sg13g2_buf_2 clkbuf_6_50_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_50_0_clk));
 sg13g2_buf_2 clkbuf_6_51_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_51_0_clk));
 sg13g2_buf_2 clkbuf_6_52_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_52_0_clk));
 sg13g2_buf_2 clkbuf_6_53_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_53_0_clk));
 sg13g2_buf_2 clkbuf_6_54_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_54_0_clk));
 sg13g2_buf_2 clkbuf_6_55_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_55_0_clk));
 sg13g2_buf_2 clkbuf_6_56_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_56_0_clk));
 sg13g2_buf_2 clkbuf_6_57_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_57_0_clk));
 sg13g2_buf_2 clkbuf_6_58_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_58_0_clk));
 sg13g2_buf_2 clkbuf_6_59_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_59_0_clk));
 sg13g2_buf_2 clkbuf_6_60_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_60_0_clk));
 sg13g2_buf_2 clkbuf_6_61_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_61_0_clk));
 sg13g2_buf_2 clkbuf_6_62_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_62_0_clk));
 sg13g2_buf_2 clkbuf_6_63_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_63_0_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_6_1_0_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_6_2_0_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_6_3_0_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_6_4_0_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_6_5_0_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_6_6_0_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_6_7_0_clk));
 sg13g2_buf_1 clkload7 (.A(clknet_6_17_0_clk));
 sg13g2_buf_2 clkload8 (.A(clknet_6_18_0_clk));
 sg13g2_buf_2 clkload9 (.A(clknet_6_19_0_clk));
 sg13g2_buf_2 clkload10 (.A(clknet_6_20_0_clk));
 sg13g2_buf_2 clkload11 (.A(clknet_6_21_0_clk));
 sg13g2_buf_2 clkload12 (.A(clknet_6_22_0_clk));
 sg13g2_buf_2 clkload13 (.A(clknet_6_23_0_clk));
 sg13g2_buf_2 clkload14 (.A(clknet_6_33_0_clk));
 sg13g2_buf_2 clkload15 (.A(clknet_6_34_0_clk));
 sg13g2_buf_2 clkload16 (.A(clknet_6_35_0_clk));
 sg13g2_buf_2 clkload17 (.A(clknet_6_36_0_clk));
 sg13g2_buf_2 clkload18 (.A(clknet_6_37_0_clk));
 sg13g2_buf_2 clkload19 (.A(clknet_6_38_0_clk));
 sg13g2_buf_2 clkload20 (.A(clknet_6_39_0_clk));
 sg13g2_buf_2 clkload21 (.A(clknet_6_49_0_clk));
 sg13g2_buf_2 clkload22 (.A(clknet_6_50_0_clk));
 sg13g2_buf_2 clkload23 (.A(clknet_6_51_0_clk));
 sg13g2_buf_2 clkload24 (.A(clknet_6_52_0_clk));
 sg13g2_buf_2 clkload25 (.A(clknet_6_53_0_clk));
 sg13g2_buf_2 clkload26 (.A(clknet_6_54_0_clk));
 sg13g2_buf_2 clkload27 (.A(clknet_6_55_0_clk));
 sg13g2_inv_1 clkload28 (.A(clknet_leaf_9_clk));
 sg13g2_inv_1 clkload29 (.A(clknet_leaf_11_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_258_clk));
 sg13g2_inv_2 clkload31 (.A(clknet_leaf_254_clk));
 sg13g2_inv_1 clkload32 (.A(clknet_leaf_14_clk));
 sg13g2_inv_1 clkload33 (.A(clknet_leaf_29_clk));
 sg13g2_inv_1 clkload34 (.A(clknet_leaf_31_clk));
 sg13g2_inv_1 clkload35 (.A(clknet_leaf_33_clk));
 sg13g2_inv_4 clkload36 (.A(clknet_leaf_41_clk));
 sg13g2_inv_4 clkload37 (.A(clknet_leaf_28_clk));
 sg13g2_inv_4 clkload38 (.A(clknet_leaf_64_clk));
 sg13g2_inv_4 clkload39 (.A(clknet_leaf_63_clk));
 sg13g2_inv_8 clkload40 (.A(clknet_leaf_164_clk));
 sg13g2_inv_1 clkload41 (.A(clknet_leaf_134_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\TRNG.ctrl_mode_sync[0] ),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold2 (.A(_00275_),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold3 (.A(_00122_),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold4 (.A(_04855_),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold5 (.A(\TRNG.Word_Out[192] ),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold6 (.A(_01437_),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold7 (.A(\TRNG.sha256.compress.done ),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold8 (.A(_00273_),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold9 (.A(_00971_),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold10 (.A(\TRNG.Word_Out[280] ),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold11 (.A(_01525_),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold12 (.A(\TRNG.Word_Out[321] ),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold13 (.A(_02014_),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold14 (.A(_00274_),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold15 (.A(_00856_),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold16 (.A(\TRNG.Word_Out[138] ),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold17 (.A(_01383_),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold18 (.A(_00121_),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold19 (.A(_02159_),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold20 (.A(\TRNG.sha256.compress.hash_gen.temp[2] ),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold21 (.A(\TRNG.sha256.compress.hash_gen.temp[1] ),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold22 (.A(\TRNG.Word_Out[24] ),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold23 (.A(_01269_),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold24 (.A(\TRNG.Word_Out[127] ),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold25 (.A(_01372_),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold26 (.A(\TRNG.Word_Out[333] ),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold27 (.A(_01578_),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold28 (.A(\TRNG.Word_Out[174] ),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold29 (.A(_01419_),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold30 (.A(\TRNG.Word_Out[224] ),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold31 (.A(_01469_),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold32 (.A(\TRNG.Word_Out[133] ),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold33 (.A(_01378_),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold34 (.A(\TRNG.Word_Out[141] ),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold35 (.A(_01386_),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold36 (.A(\TRNG.Word_Out[345] ),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold37 (.A(_01590_),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold38 (.A(\TRNG.Word_Out[322] ),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold39 (.A(_02015_),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold40 (.A(\TRNG.Word_Out[409] ),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold41 (.A(_01654_),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold42 (.A(\TRNG.Word_Out[63] ),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold43 (.A(_01308_),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold44 (.A(\TRNG.Word_Out[324] ),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold45 (.A(_01569_),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold46 (.A(\TRNG.Word_Out[389] ),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold47 (.A(_01634_),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold48 (.A(\TRNG.Word_Out[93] ),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold49 (.A(_01338_),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold50 (.A(\TRNG.Word_Out[376] ),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold51 (.A(_01621_),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold52 (.A(_00272_),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold53 (.A(_00975_),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold54 (.A(\TRNG.Word_Out[103] ),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold55 (.A(_01348_),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold56 (.A(\TRNG.sha256.compress.hash_gen.temp[0] ),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold57 (.A(\TRNG.Word_Out[348] ),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold58 (.A(_01593_),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold59 (.A(\TRNG.Word_Out[355] ),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold60 (.A(_01600_),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold61 (.A(\TRNG.Word_Out[154] ),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold62 (.A(_01399_),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold63 (.A(\TRNG.Word_Out[30] ),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold64 (.A(_01275_),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold65 (.A(\TRNG.Word_Out[7] ),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold66 (.A(_01252_),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold67 (.A(\TRNG.Word_Out[254] ),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold68 (.A(_01499_),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold69 (.A(\TRNG.Word_Out[323] ),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold70 (.A(\TRNG.Word_Out[312] ),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold71 (.A(_01557_),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold72 (.A(\TRNG.Word_Out[78] ),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold73 (.A(_01323_),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold74 (.A(\TRNG.Word_Out[189] ),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold75 (.A(_01434_),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold76 (.A(\TRNG.Word_Out[381] ),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold77 (.A(_01626_),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold78 (.A(\TRNG.Word_Out[70] ),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold79 (.A(_01315_),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold80 (.A(\TRNG.Word_Out[228] ),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold81 (.A(_01473_),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold82 (.A(_00116_),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold83 (.A(_00310_),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold84 (.A(\TRNG.Word_Out[291] ),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold85 (.A(_01536_),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold86 (.A(\TRNG.Padded_Out[219] ),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold87 (.A(\TRNG.Word_Out[60] ),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold88 (.A(_01305_),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold89 (.A(\TRNG.Word_Out[125] ),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold90 (.A(_01370_),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold91 (.A(\TRNG.Word_Out[359] ),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold92 (.A(_01604_),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold93 (.A(\TRNG.Word_Out[135] ),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold94 (.A(_01380_),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold95 (.A(\TRNG.Word_Out[36] ),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold96 (.A(_01281_),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold97 (.A(\TRNG.Word_Out[112] ),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold98 (.A(_01357_),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold99 (.A(\TRNG.Word_Out[397] ),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold100 (.A(_01642_),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold101 (.A(\TRNG.Word_Out[13] ),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold102 (.A(_01258_),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold103 (.A(\TRNG.Word_Out[29] ),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold104 (.A(\TRNG.Word_Out[393] ),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold105 (.A(_01638_),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold106 (.A(\TRNG.Padded_Out[145] ),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold107 (.A(_01773_),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold108 (.A(\TRNG.Word_Out[157] ),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold109 (.A(_01402_),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold110 (.A(\TRNG.Padded_Out[177] ),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold111 (.A(\TRNG.Word_Out[38] ),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold112 (.A(_01283_),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold113 (.A(\TRNG.Word_Out[88] ),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold114 (.A(_01333_),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold115 (.A(\TRNG.Padded_Out[333] ),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold116 (.A(_01961_),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold117 (.A(\TRNG.Word_Out[294] ),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold118 (.A(_01539_),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold119 (.A(\TRNG.Padded_Out[141] ),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold120 (.A(_01769_),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold121 (.A(\TRNG.Padded_Out[265] ),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold122 (.A(_01893_),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold123 (.A(\TRNG.Padded_Out[417] ),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold124 (.A(_02045_),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold125 (.A(\TRNG.Word_Out[265] ),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold126 (.A(_01510_),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold127 (.A(\TRNG.Padded_Out[413] ),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold128 (.A(\TRNG.Padded_Out[458] ),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold129 (.A(\TRNG.Repetition_Count_Test.count[0] ),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold130 (.A(_00096_),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold131 (.A(\TRNG.Padded_Out[79] ),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold132 (.A(_01707_),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold133 (.A(\TRNG.Padded_Out[180] ),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold134 (.A(_01808_),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold135 (.A(\TRNG.Padded_Out[275] ),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold136 (.A(_01903_),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold137 (.A(\TRNG.Padded_Out[309] ),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold138 (.A(_01937_),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold139 (.A(\TRNG.Padded_Out[159] ),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold140 (.A(_01787_),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold141 (.A(\TRNG.Padded_Out[410] ),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold142 (.A(\TRNG.Padded_Out[185] ),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold143 (.A(_01813_),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold144 (.A(\TRNG.Padded_Out[487] ),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold145 (.A(_02115_),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold146 (.A(\TRNG.Padded_Out[249] ),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold147 (.A(_01877_),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold148 (.A(\TRNG.Padded_Out[412] ),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold149 (.A(_02040_),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold150 (.A(\TRNG.Padded_Out[263] ),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold151 (.A(_01891_),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold152 (.A(\TRNG.Word_Out[200] ),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold153 (.A(_01445_),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold154 (.A(\TRNG.Padded_Out[337] ),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold155 (.A(_01965_),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold156 (.A(\TRNG.Padded_Out[248] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold157 (.A(_01876_),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold158 (.A(\TRNG.Word_Out[313] ),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold159 (.A(_02006_),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold160 (.A(\TRNG.Padded_Out[390] ),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold161 (.A(_02018_),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold162 (.A(\TRNG.Word_Out[318] ),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold163 (.A(_01563_),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold164 (.A(\TRNG.Padded_Out[88] ),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold165 (.A(_01716_),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold166 (.A(\TRNG.Padded_Out[259] ),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold167 (.A(_01887_),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold168 (.A(\TRNG.Padded_Out[315] ),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold169 (.A(_01943_),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold170 (.A(\TRNG.Word_Out[303] ),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold171 (.A(_01548_),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold172 (.A(\TRNG.Padded_Out[401] ),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold173 (.A(_02029_),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold174 (.A(\TRNG.Padded_Out[256] ),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold175 (.A(_01884_),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold176 (.A(\TRNG.Padded_Out[395] ),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold177 (.A(_02023_),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold178 (.A(\TRNG.Padded_Out[128] ),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold179 (.A(\TRNG.Padded_Out[152] ),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold180 (.A(_01780_),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold181 (.A(\TRNG.Padded_Out[411] ),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold182 (.A(_02039_),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold183 (.A(\TRNG.Padded_Out[384] ),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold184 (.A(_02012_),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold185 (.A(\TRNG.Padded_Out[213] ),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold186 (.A(_01841_),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold187 (.A(\TRNG.Padded_Out[327] ),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold188 (.A(_01955_),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold189 (.A(\TRNG.Padded_Out[364] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold190 (.A(_01992_),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold191 (.A(\TRNG.Padded_Out[155] ),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold192 (.A(_01783_),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold193 (.A(\TRNG.Padded_Out[323] ),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold194 (.A(_01951_),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold195 (.A(\TRNG.Padded_Out[382] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold196 (.A(_02010_),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold197 (.A(\TRNG.Padded_Out[373] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold198 (.A(_02001_),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold199 (.A(\TRNG.Padded_Out[164] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold200 (.A(_01792_),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold201 (.A(\TRNG.Padded_Out[332] ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold202 (.A(_01960_),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold203 (.A(\TRNG.Padded_Out[114] ),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold204 (.A(_01742_),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold205 (.A(\TRNG.Padded_Out[396] ),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold206 (.A(_02024_),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold207 (.A(\TRNG.Padded_Out[419] ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold208 (.A(_02047_),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold209 (.A(\TRNG.Padded_Out[392] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold210 (.A(_02020_),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold211 (.A(\TRNG.Padded_Out[235] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold212 (.A(_01863_),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold213 (.A(\TRNG.Word_Out[87] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold214 (.A(\TRNG.Padded_Out[348] ),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold215 (.A(_01976_),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold216 (.A(\TRNG.Padded_Out[285] ),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold217 (.A(_01913_),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold218 (.A(\TRNG.Padded_Out[379] ),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold219 (.A(_02007_),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold220 (.A(\TRNG.Word_Out[249] ),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold221 (.A(_01494_),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold222 (.A(\TRNG.Padded_Out[351] ),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold223 (.A(_01979_),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold224 (.A(\TRNG.Padded_Out[328] ),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold225 (.A(_01956_),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold226 (.A(\TRNG.Padded_Out[366] ),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold227 (.A(_01994_),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold228 (.A(\TRNG.Padded_Out[507] ),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold229 (.A(_02135_),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold230 (.A(\TRNG.Padded_Out[404] ),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold231 (.A(_02032_),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold232 (.A(\TRNG.Padded_Out[321] ),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold233 (.A(_01949_),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold234 (.A(\TRNG.Word_Out[15] ),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold235 (.A(_01260_),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold236 (.A(\TRNG.Padded_Out[146] ),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold237 (.A(_01774_),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold238 (.A(\TRNG.Padded_Out[383] ),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold239 (.A(\TRNG.Word_Out[131] ),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold240 (.A(_01376_),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold241 (.A(\TRNG.Padded_Out[276] ),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold242 (.A(_01904_),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold243 (.A(\TRNG.Word_Out[263] ),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold244 (.A(_01508_),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold245 (.A(\TRNG.Padded_Out[154] ),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold246 (.A(_01782_),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold247 (.A(\TRNG.Padded_Out[142] ),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold248 (.A(_01770_),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold249 (.A(\TRNG.Padded_Out[278] ),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold250 (.A(_01906_),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold251 (.A(\TRNG.Padded_Out[313] ),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold252 (.A(_01941_),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold253 (.A(\TRNG.Word_Out[349] ),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold254 (.A(_01594_),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold255 (.A(\TRNG.Padded_Out[277] ),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold256 (.A(_01905_),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold257 (.A(\TRNG.Padded_Out[439] ),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold258 (.A(_02067_),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold259 (.A(\TRNG.Word_Out[395] ),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold260 (.A(_01640_),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold261 (.A(\TRNG.Padded_Out[93] ),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold262 (.A(_01721_),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold263 (.A(\TRNG.Padded_Out[280] ),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold264 (.A(_01908_),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold265 (.A(\TRNG.Word_Out[327] ),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold266 (.A(_01572_),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold267 (.A(\TRNG.Padded_Out[184] ),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold268 (.A(_01812_),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold269 (.A(\TRNG.Padded_Out[446] ),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold270 (.A(\TRNG.Word_Out[413] ),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold271 (.A(_01658_),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold272 (.A(\TRNG.Padded_Out[90] ),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold273 (.A(_01718_),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold274 (.A(\TRNG.Padded_Out[69] ),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold275 (.A(_01697_),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold276 (.A(\TRNG.Padded_Out[153] ),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold277 (.A(\TRNG.Repetition_Count_Test.count[3] ),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold278 (.A(_06333_),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold279 (.A(_00099_),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold280 (.A(\TRNG.Padded_Out[202] ),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold281 (.A(_01830_),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold282 (.A(\TRNG.Word_Out[285] ),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold283 (.A(_01530_),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold284 (.A(\TRNG.Padded_Out[400] ),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold285 (.A(_02028_),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold286 (.A(\TRNG.Padded_Out[197] ),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold287 (.A(_01825_),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold288 (.A(\TRNG.Padded_Out[252] ),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold289 (.A(_01880_),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold290 (.A(\TRNG.Padded_Out[86] ),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold291 (.A(_01714_),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold292 (.A(\TRNG.Padded_Out[370] ),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold293 (.A(_01998_),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold294 (.A(\TRNG.Padded_Out[172] ),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold295 (.A(_01800_),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold296 (.A(\TRNG.Padded_Out[78] ),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold297 (.A(\TRNG.Word_Out[388] ),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold298 (.A(\TRNG.Padded_Out[443] ),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold299 (.A(_02071_),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold300 (.A(\TRNG.Word_Out[240] ),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold301 (.A(_01485_),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold302 (.A(\TRNG.Padded_Out[144] ),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold303 (.A(_01772_),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold304 (.A(\TRNG.Padded_Out[116] ),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold305 (.A(_01744_),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold306 (.A(\TRNG.Padded_Out[462] ),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold307 (.A(\TRNG.Padded_Out[301] ),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold308 (.A(_01929_),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold309 (.A(\TRNG.Padded_Out[239] ),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold310 (.A(\TRNG.Padded_Out[308] ),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold311 (.A(_01936_),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold312 (.A(\TRNG.Padded_Out[74] ),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold313 (.A(_01702_),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold314 (.A(\TRNG.Padded_Out[433] ),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold315 (.A(_02061_),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold316 (.A(\TRNG.Padded_Out[476] ),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold317 (.A(_02104_),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold318 (.A(\TRNG.Padded_Out[245] ),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold319 (.A(_01873_),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold320 (.A(\TRNG.Padded_Out[121] ),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold321 (.A(_01749_),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold322 (.A(\TRNG.Padded_Out[464] ),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold323 (.A(_02092_),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold324 (.A(\TRNG.Padded_Out[264] ),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold325 (.A(_01892_),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold326 (.A(\TRNG.Padded_Out[233] ),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold327 (.A(_01861_),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold328 (.A(\TRNG.Padded_Out[459] ),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold329 (.A(_02087_),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold330 (.A(\TRNG.Padded_Out[220] ),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold331 (.A(_01848_),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold332 (.A(\TRNG.Padded_Out[198] ),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold333 (.A(\TRNG.Word_Out[113] ),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold334 (.A(_01358_),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold335 (.A(\TRNG.Padded_Out[363] ),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold336 (.A(_01991_),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold337 (.A(\TRNG.Padded_Out[147] ),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold338 (.A(_01775_),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold339 (.A(\TRNG.Padded_Out[234] ),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold340 (.A(_01862_),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold341 (.A(\TRNG.Word_Out[426] ),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold342 (.A(_01671_),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold343 (.A(\TRNG.Word_Out[400] ),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold344 (.A(_01645_),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold345 (.A(\TRNG.Padded_Out[349] ),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold346 (.A(_01977_),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold347 (.A(\TRNG.Padded_Out[200] ),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold348 (.A(\TRNG.Padded_Out[362] ),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold349 (.A(_01990_),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold350 (.A(\TRNG.Padded_Out[80] ),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold351 (.A(\TRNG.Padded_Out[204] ),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold352 (.A(_01832_),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold353 (.A(\TRNG.Padded_Out[331] ),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold354 (.A(_01959_),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold355 (.A(\TRNG.Padded_Out[195] ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold356 (.A(_01823_),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold357 (.A(\TRNG.Padded_Out[232] ),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold358 (.A(_01860_),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold359 (.A(\TRNG.Padded_Out[449] ),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold360 (.A(_02077_),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold361 (.A(\TRNG.Padded_Out[437] ),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold362 (.A(_02065_),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold363 (.A(\TRNG.Padded_Out[181] ),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold364 (.A(_01809_),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold365 (.A(\TRNG.Word_Out[166] ),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold366 (.A(_01411_),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold367 (.A(\TRNG.Padded_Out[257] ),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold368 (.A(\TRNG.Padded_Out[372] ),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold369 (.A(_02000_),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold370 (.A(\TRNG.Padded_Out[287] ),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold371 (.A(_01915_),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold372 (.A(\TRNG.Padded_Out[422] ),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold373 (.A(_02050_),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold374 (.A(\TRNG.Padded_Out[416] ),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold375 (.A(_02044_),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold376 (.A(\TRNG.Padded_Out[451] ),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold377 (.A(_02079_),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold378 (.A(\TRNG.Word_Out[111] ),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold379 (.A(_01804_),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold380 (.A(\TRNG.Padded_Out[486] ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold381 (.A(_02114_),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold382 (.A(\TRNG.Padded_Out[189] ),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold383 (.A(_01817_),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold384 (.A(\TRNG.Padded_Out[441] ),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold385 (.A(\TRNG.Padded_Out[143] ),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold386 (.A(\TRNG.Padded_Out[335] ),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold387 (.A(_01963_),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold388 (.A(\TRNG.Padded_Out[168] ),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold389 (.A(\TRNG.Padded_Out[377] ),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold390 (.A(\TRNG.Padded_Out[87] ),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold391 (.A(_01715_),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold392 (.A(\TRNG.Padded_Out[140] ),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold393 (.A(_01768_),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold394 (.A(\TRNG.Padded_Out[444] ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold395 (.A(_02072_),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold396 (.A(\TRNG.Padded_Out[431] ),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold397 (.A(_02059_),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold398 (.A(\TRNG.Padded_Out[161] ),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold399 (.A(_01789_),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold400 (.A(\TRNG.Padded_Out[316] ),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold401 (.A(_01944_),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold402 (.A(\TRNG.Padded_Out[270] ),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold403 (.A(_01898_),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold404 (.A(_00271_),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold405 (.A(_00979_),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold406 (.A(\TRNG.Padded_Out[380] ),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold407 (.A(_02008_),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold408 (.A(\TRNG.Padded_Out[454] ),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold409 (.A(\TRNG.Padded_Out[84] ),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold410 (.A(_01712_),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold411 (.A(\TRNG.Padded_Out[85] ),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold412 (.A(_01713_),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold413 (.A(\TRNG.Word_Out[149] ),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold414 (.A(_01394_),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold415 (.A(\TRNG.Padded_Out[371] ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold416 (.A(_01999_),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold417 (.A(\TRNG.Padded_Out[179] ),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold418 (.A(_01807_),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold419 (.A(\TRNG.Padded_Out[432] ),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold420 (.A(_02060_),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold421 (.A(\TRNG.Word_Out[120] ),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold422 (.A(_01365_),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold423 (.A(\TRNG.Padded_Out[426] ),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold424 (.A(_02054_),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold425 (.A(\TRNG.Padded_Out[73] ),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold426 (.A(_01701_),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold427 (.A(\TRNG.Padded_Out[261] ),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold428 (.A(_01889_),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold429 (.A(\TRNG.Padded_Out[474] ),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold430 (.A(\TRNG.Padded_Out[355] ),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold431 (.A(_01983_),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold432 (.A(\TRNG.Word_Out[247] ),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold433 (.A(_01492_),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold434 (.A(\TRNG.Padded_Out[120] ),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold435 (.A(_01748_),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold436 (.A(_00126_),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold437 (.A(_05905_),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold438 (.A(_00102_),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold439 (.A(\TRNG.Padded_Out[463] ),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold440 (.A(_02091_),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold441 (.A(\TRNG.Word_Out[169] ),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold442 (.A(_01414_),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold443 (.A(\TRNG.Padded_Out[268] ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold444 (.A(_01896_),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold445 (.A(\TRNG.Word_Out[197] ),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold446 (.A(_01442_),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold447 (.A(\TRNG.Padded_Out[149] ),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold448 (.A(_01777_),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold449 (.A(\TRNG.Word_Out[71] ),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold450 (.A(_01316_),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold451 (.A(\TRNG.Word_Out[164] ),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold452 (.A(_01409_),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold453 (.A(\TRNG.Padded_Out[394] ),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold454 (.A(_02022_),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold455 (.A(\TRNG.Padded_Out[133] ),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold456 (.A(_01761_),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold457 (.A(\TRNG.Padded_Out[324] ),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold458 (.A(_01952_),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold459 (.A(\TRNG.Padded_Out[162] ),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold460 (.A(_01790_),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold461 (.A(\TRNG.Padded_Out[447] ),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold462 (.A(_02075_),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold463 (.A(\TRNG.Padded_Out[445] ),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold464 (.A(_02073_),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold465 (.A(\TRNG.Padded_Out[340] ),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold466 (.A(_01968_),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold467 (.A(\TRNG.Padded_Out[456] ),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold468 (.A(_02084_),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold469 (.A(\TRNG.Padded_Out[479] ),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold470 (.A(_02107_),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold471 (.A(\TRNG.Word_Out[357] ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold472 (.A(_01602_),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold473 (.A(\TRNG.Word_Out[14] ),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold474 (.A(\TRNG.Word_Out[326] ),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold475 (.A(\TRNG.Padded_Out[163] ),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold476 (.A(_01791_),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold477 (.A(\TRNG.Padded_Out[402] ),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold478 (.A(_02030_),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold479 (.A(\TRNG.Word_Out[387] ),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold480 (.A(\TRNG.Padded_Out[510] ),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold481 (.A(_02138_),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold482 (.A(\TRNG.Padded_Out[169] ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold483 (.A(_01797_),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold484 (.A(\TRNG.Padded_Out[466] ),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold485 (.A(_02094_),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold486 (.A(\TRNG.Padded_Out[273] ),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold487 (.A(_01901_),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold488 (.A(\TRNG.Padded_Out[442] ),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold489 (.A(_02070_),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold490 (.A(\TRNG.Padded_Out[272] ),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold491 (.A(_01900_),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold492 (.A(\TRNG.Padded_Out[289] ),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold493 (.A(\TRNG.Padded_Out[207] ),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold494 (.A(_01835_),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold495 (.A(\TRNG.Word_Out[266] ),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold496 (.A(_01511_),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold497 (.A(\TRNG.Padded_Out[457] ),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold498 (.A(_02085_),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold499 (.A(\TRNG.Padded_Out[399] ),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold500 (.A(_02027_),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold501 (.A(\TRNG.Padded_Out[389] ),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold502 (.A(\TRNG.Padded_Out[350] ),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold503 (.A(\TRNG.Padded_Out[279] ),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold504 (.A(_01907_),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold505 (.A(\TRNG.Word_Out[420] ),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold506 (.A(_01665_),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold507 (.A(\TRNG.Padded_Out[375] ),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold508 (.A(_02003_),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold509 (.A(\TRNG.Padded_Out[354] ),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold510 (.A(_01982_),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold511 (.A(\TRNG.Padded_Out[409] ),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold512 (.A(_02037_),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold513 (.A(\TRNG.Padded_Out[317] ),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold514 (.A(_01945_),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold515 (.A(\TRNG.Word_Out[104] ),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold516 (.A(_01349_),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold517 (.A(\TRNG.Padded_Out[294] ),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold518 (.A(_01922_),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold519 (.A(\TRNG.Padded_Out[356] ),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold520 (.A(\TRNG.Padded_Out[428] ),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold521 (.A(_02056_),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold522 (.A(\TRNG.Word_Out[428] ),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold523 (.A(_01673_),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold524 (.A(\TRNG.Padded_Out[231] ),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold525 (.A(\TRNG.Word_Out[40] ),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold526 (.A(_01285_),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold527 (.A(\TRNG.Padded_Out[236] ),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold528 (.A(_01864_),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold529 (.A(\TRNG.Padded_Out[131] ),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold530 (.A(_01759_),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold531 (.A(\TRNG.Padded_Out[113] ),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold532 (.A(_01741_),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold533 (.A(\TRNG.Word_Out[390] ),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold534 (.A(_01635_),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold535 (.A(\TRNG.Padded_Out[488] ),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold536 (.A(_02116_),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold537 (.A(\TRNG.Padded_Out[418] ),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold538 (.A(_02046_),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold539 (.A(\TRNG.Padded_Out[243] ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold540 (.A(_01871_),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold541 (.A(\TRNG.Padded_Out[414] ),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold542 (.A(\TRNG.Padded_Out[182] ),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold543 (.A(_01810_),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold544 (.A(\TRNG.Padded_Out[199] ),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold545 (.A(_01827_),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold546 (.A(\TRNG.Padded_Out[75] ),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold547 (.A(_01703_),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold548 (.A(\TRNG.Padded_Out[367] ),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold549 (.A(_01995_),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold550 (.A(\TRNG.Padded_Out[119] ),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold551 (.A(_01747_),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold552 (.A(\TRNG.Word_Out[332] ),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold553 (.A(\TRNG.Word_Out[121] ),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold554 (.A(_01814_),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold555 (.A(\TRNG.Padded_Out[253] ),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold556 (.A(_01881_),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold557 (.A(\TRNG.Padded_Out[139] ),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold558 (.A(_01767_),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold559 (.A(\TRNG.Padded_Out[421] ),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold560 (.A(_02049_),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold561 (.A(\TRNG.Padded_Out[170] ),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold562 (.A(_01798_),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold563 (.A(\TRNG.Padded_Out[299] ),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold564 (.A(_01927_),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold565 (.A(\TRNG.Padded_Out[117] ),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold566 (.A(_01745_),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold567 (.A(\TRNG.Padded_Out[473] ),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold568 (.A(_02101_),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold569 (.A(\TRNG.Padded_Out[83] ),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold570 (.A(_01711_),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold571 (.A(\TRNG.Padded_Out[71] ),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold572 (.A(_01699_),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold573 (.A(\TRNG.Padded_Out[260] ),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold574 (.A(_01888_),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold575 (.A(\TRNG.sha256.compress.hash_gen.temp[3] ),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold576 (.A(\TRNG.Padded_Out[72] ),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold577 (.A(\TRNG.Padded_Out[274] ),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold578 (.A(_01902_),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold579 (.A(\TRNG.Padded_Out[167] ),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold580 (.A(_01795_),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold581 (.A(\TRNG.Padded_Out[122] ),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold582 (.A(_01750_),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold583 (.A(\TRNG.Padded_Out[214] ),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold584 (.A(\TRNG.Padded_Out[175] ),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold585 (.A(_01803_),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold586 (.A(\TRNG.Padded_Out[461] ),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold587 (.A(_02089_),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold588 (.A(\TRNG.Padded_Out[246] ),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold589 (.A(_01874_),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold590 (.A(\TRNG.Word_Out[9] ),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold591 (.A(_01254_),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold592 (.A(\TRNG.Padded_Out[111] ),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold593 (.A(_01739_),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold594 (.A(\TRNG.Word_Out[55] ),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold595 (.A(_01300_),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold596 (.A(\TRNG.Word_Out[72] ),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold597 (.A(_01317_),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold598 (.A(\TRNG.Padded_Out[226] ),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold599 (.A(_01854_),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold600 (.A(\TRNG.Padded_Out[290] ),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold601 (.A(_01918_),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold602 (.A(\TRNG.Padded_Out[427] ),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold603 (.A(_02055_),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold604 (.A(\TRNG.Word_Out[267] ),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold605 (.A(_01512_),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold606 (.A(\TRNG.Padded_Out[151] ),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold607 (.A(_01779_),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold608 (.A(\TRNG.Word_Out[102] ),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold609 (.A(\TRNG.Padded_Out[284] ),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold610 (.A(_01912_),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold611 (.A(\TRNG.Padded_Out[225] ),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold612 (.A(_01853_),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold613 (.A(\TRNG.Word_Out[229] ),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold614 (.A(_01474_),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold615 (.A(\TRNG.Padded_Out[208] ),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold616 (.A(_01836_),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold617 (.A(\TRNG.Padded_Out[344] ),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold618 (.A(_01972_),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold619 (.A(\TRNG.Padded_Out[436] ),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold620 (.A(_02064_),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold621 (.A(\TRNG.Word_Out[198] ),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold622 (.A(_01443_),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold623 (.A(\TRNG.Word_Out[289] ),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold624 (.A(_01534_),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold625 (.A(\TRNG.Padded_Out[415] ),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold626 (.A(_02043_),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold627 (.A(\TRNG.Padded_Out[212] ),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold628 (.A(_01840_),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold629 (.A(\TRNG.Padded_Out[70] ),
    .X(net1757));
 sg13g2_dlygate4sd3_1 hold630 (.A(_01698_),
    .X(net1758));
 sg13g2_dlygate4sd3_1 hold631 (.A(\TRNG.Word_Out[260] ),
    .X(net1759));
 sg13g2_dlygate4sd3_1 hold632 (.A(_01505_),
    .X(net1760));
 sg13g2_dlygate4sd3_1 hold633 (.A(\TRNG.Padded_Out[107] ),
    .X(net1761));
 sg13g2_dlygate4sd3_1 hold634 (.A(_01735_),
    .X(net1762));
 sg13g2_dlygate4sd3_1 hold635 (.A(\TRNG.Word_Out[94] ),
    .X(net1763));
 sg13g2_dlygate4sd3_1 hold636 (.A(_01339_),
    .X(net1764));
 sg13g2_dlygate4sd3_1 hold637 (.A(\TRNG.Padded_Out[218] ),
    .X(net1765));
 sg13g2_dlygate4sd3_1 hold638 (.A(_01846_),
    .X(net1766));
 sg13g2_dlygate4sd3_1 hold639 (.A(\TRNG.Padded_Out[210] ),
    .X(net1767));
 sg13g2_dlygate4sd3_1 hold640 (.A(_01838_),
    .X(net1768));
 sg13g2_dlygate4sd3_1 hold641 (.A(\TRNG.Padded_Out[398] ),
    .X(net1769));
 sg13g2_dlygate4sd3_1 hold642 (.A(\TRNG.Padded_Out[338] ),
    .X(net1770));
 sg13g2_dlygate4sd3_1 hold643 (.A(_01966_),
    .X(net1771));
 sg13g2_dlygate4sd3_1 hold644 (.A(\TRNG.Padded_Out[127] ),
    .X(net1772));
 sg13g2_dlygate4sd3_1 hold645 (.A(_01755_),
    .X(net1773));
 sg13g2_dlygate4sd3_1 hold646 (.A(\TRNG.Padded_Out[336] ),
    .X(net1774));
 sg13g2_dlygate4sd3_1 hold647 (.A(_01964_),
    .X(net1775));
 sg13g2_dlygate4sd3_1 hold648 (.A(\TRNG.Padded_Out[374] ),
    .X(net1776));
 sg13g2_dlygate4sd3_1 hold649 (.A(_02002_),
    .X(net1777));
 sg13g2_dlygate4sd3_1 hold650 (.A(\TRNG.Padded_Out[300] ),
    .X(net1778));
 sg13g2_dlygate4sd3_1 hold651 (.A(_01928_),
    .X(net1779));
 sg13g2_dlygate4sd3_1 hold652 (.A(\TRNG.Padded_Out[148] ),
    .X(net1780));
 sg13g2_dlygate4sd3_1 hold653 (.A(_01776_),
    .X(net1781));
 sg13g2_dlygate4sd3_1 hold654 (.A(\TRNG.Padded_Out[346] ),
    .X(net1782));
 sg13g2_dlygate4sd3_1 hold655 (.A(_01974_),
    .X(net1783));
 sg13g2_dlygate4sd3_1 hold656 (.A(\TRNG.Padded_Out[237] ),
    .X(net1784));
 sg13g2_dlygate4sd3_1 hold657 (.A(_01865_),
    .X(net1785));
 sg13g2_dlygate4sd3_1 hold658 (.A(\TRNG.Padded_Out[130] ),
    .X(net1786));
 sg13g2_dlygate4sd3_1 hold659 (.A(_01758_),
    .X(net1787));
 sg13g2_dlygate4sd3_1 hold660 (.A(\TRNG.Word_Out[262] ),
    .X(net1788));
 sg13g2_dlygate4sd3_1 hold661 (.A(\TRNG.Padded_Out[365] ),
    .X(net1789));
 sg13g2_dlygate4sd3_1 hold662 (.A(_01993_),
    .X(net1790));
 sg13g2_dlygate4sd3_1 hold663 (.A(\TRNG.Padded_Out[123] ),
    .X(net1791));
 sg13g2_dlygate4sd3_1 hold664 (.A(_01751_),
    .X(net1792));
 sg13g2_dlygate4sd3_1 hold665 (.A(\TRNG.Padded_Out[194] ),
    .X(net1793));
 sg13g2_dlygate4sd3_1 hold666 (.A(_01822_),
    .X(net1794));
 sg13g2_dlygate4sd3_1 hold667 (.A(\TRNG.Word_Out[430] ),
    .X(net1795));
 sg13g2_dlygate4sd3_1 hold668 (.A(_01675_),
    .X(net1796));
 sg13g2_dlygate4sd3_1 hold669 (.A(\TRNG.Padded_Out[368] ),
    .X(net1797));
 sg13g2_dlygate4sd3_1 hold670 (.A(\TRNG.Padded_Out[326] ),
    .X(net1798));
 sg13g2_dlygate4sd3_1 hold671 (.A(_01954_),
    .X(net1799));
 sg13g2_dlygate4sd3_1 hold672 (.A(\TRNG.Padded_Out[291] ),
    .X(net1800));
 sg13g2_dlygate4sd3_1 hold673 (.A(_01919_),
    .X(net1801));
 sg13g2_dlygate4sd3_1 hold674 (.A(\TRNG.Padded_Out[251] ),
    .X(net1802));
 sg13g2_dlygate4sd3_1 hold675 (.A(_01879_),
    .X(net1803));
 sg13g2_dlygate4sd3_1 hold676 (.A(\TRNG.Word_Out[435] ),
    .X(net1804));
 sg13g2_dlygate4sd3_1 hold677 (.A(_01680_),
    .X(net1805));
 sg13g2_dlygate4sd3_1 hold678 (.A(\TRNG.Padded_Out[334] ),
    .X(net1806));
 sg13g2_dlygate4sd3_1 hold679 (.A(_01962_),
    .X(net1807));
 sg13g2_dlygate4sd3_1 hold680 (.A(\TRNG.Padded_Out[183] ),
    .X(net1808));
 sg13g2_dlygate4sd3_1 hold681 (.A(_01811_),
    .X(net1809));
 sg13g2_dlygate4sd3_1 hold682 (.A(\TRNG.Padded_Out[267] ),
    .X(net1810));
 sg13g2_dlygate4sd3_1 hold683 (.A(_01895_),
    .X(net1811));
 sg13g2_dlygate4sd3_1 hold684 (.A(\TRNG.Padded_Out[471] ),
    .X(net1812));
 sg13g2_dlygate4sd3_1 hold685 (.A(_02099_),
    .X(net1813));
 sg13g2_dlygate4sd3_1 hold686 (.A(\TRNG.Padded_Out[438] ),
    .X(net1814));
 sg13g2_dlygate4sd3_1 hold687 (.A(_02066_),
    .X(net1815));
 sg13g2_dlygate4sd3_1 hold688 (.A(\TRNG.Word_Out[98] ),
    .X(net1816));
 sg13g2_dlygate4sd3_1 hold689 (.A(_01343_),
    .X(net1817));
 sg13g2_dlygate4sd3_1 hold690 (.A(\TRNG.Word_Out[384] ),
    .X(net1818));
 sg13g2_dlygate4sd3_1 hold691 (.A(_01629_),
    .X(net1819));
 sg13g2_dlygate4sd3_1 hold692 (.A(\TRNG.Word_Out[6] ),
    .X(net1820));
 sg13g2_dlygate4sd3_1 hold693 (.A(\TRNG.Word_Out[46] ),
    .X(net1821));
 sg13g2_dlygate4sd3_1 hold694 (.A(_01291_),
    .X(net1822));
 sg13g2_dlygate4sd3_1 hold695 (.A(\TRNG.Word_Out[163] ),
    .X(net1823));
 sg13g2_dlygate4sd3_1 hold696 (.A(\TRNG.Padded_Out[429] ),
    .X(net1824));
 sg13g2_dlygate4sd3_1 hold697 (.A(_02057_),
    .X(net1825));
 sg13g2_dlygate4sd3_1 hold698 (.A(\TRNG.Padded_Out[206] ),
    .X(net1826));
 sg13g2_dlygate4sd3_1 hold699 (.A(\TRNG.Padded_Out[68] ),
    .X(net1827));
 sg13g2_dlygate4sd3_1 hold700 (.A(_01696_),
    .X(net1828));
 sg13g2_dlygate4sd3_1 hold701 (.A(\TRNG.Padded_Out[455] ),
    .X(net1829));
 sg13g2_dlygate4sd3_1 hold702 (.A(\TRNG.Padded_Out[115] ),
    .X(net1830));
 sg13g2_dlygate4sd3_1 hold703 (.A(_01743_),
    .X(net1831));
 sg13g2_dlygate4sd3_1 hold704 (.A(\TRNG.Word_Out[107] ),
    .X(net1832));
 sg13g2_dlygate4sd3_1 hold705 (.A(_01352_),
    .X(net1833));
 sg13g2_dlygate4sd3_1 hold706 (.A(\TRNG.Padded_Out[201] ),
    .X(net1834));
 sg13g2_dlygate4sd3_1 hold707 (.A(_01829_),
    .X(net1835));
 sg13g2_dlygate4sd3_1 hold708 (.A(\TRNG.Word_Out[231] ),
    .X(net1836));
 sg13g2_dlygate4sd3_1 hold709 (.A(_01476_),
    .X(net1837));
 sg13g2_dlygate4sd3_1 hold710 (.A(\TRNG.Padded_Out[65] ),
    .X(net1838));
 sg13g2_dlygate4sd3_1 hold711 (.A(_01693_),
    .X(net1839));
 sg13g2_dlygate4sd3_1 hold712 (.A(\TRNG.Padded_Out[241] ),
    .X(net1840));
 sg13g2_dlygate4sd3_1 hold713 (.A(_01869_),
    .X(net1841));
 sg13g2_dlygate4sd3_1 hold714 (.A(\TRNG.Padded_Out[196] ),
    .X(net1842));
 sg13g2_dlygate4sd3_1 hold715 (.A(\TRNG.Padded_Out[258] ),
    .X(net1843));
 sg13g2_dlygate4sd3_1 hold716 (.A(_01886_),
    .X(net1844));
 sg13g2_dlygate4sd3_1 hold717 (.A(\TRNG.Padded_Out[100] ),
    .X(net1845));
 sg13g2_dlygate4sd3_1 hold718 (.A(_01728_),
    .X(net1846));
 sg13g2_dlygate4sd3_1 hold719 (.A(\TRNG.Padded_Out[320] ),
    .X(net1847));
 sg13g2_dlygate4sd3_1 hold720 (.A(_01948_),
    .X(net1848));
 sg13g2_dlygate4sd3_1 hold721 (.A(\TRNG.Padded_Out[171] ),
    .X(net1849));
 sg13g2_dlygate4sd3_1 hold722 (.A(_01799_),
    .X(net1850));
 sg13g2_dlygate4sd3_1 hold723 (.A(\TRNG.Word_Out[258] ),
    .X(net1851));
 sg13g2_dlygate4sd3_1 hold724 (.A(_01503_),
    .X(net1852));
 sg13g2_dlygate4sd3_1 hold725 (.A(\TRNG.sha256.expand.exp_ctrl.sum[22] ),
    .X(net1853));
 sg13g2_dlygate4sd3_1 hold726 (.A(_01009_),
    .X(net1854));
 sg13g2_dlygate4sd3_1 hold727 (.A(\TRNG.Padded_Out[302] ),
    .X(net1855));
 sg13g2_dlygate4sd3_1 hold728 (.A(_01930_),
    .X(net1856));
 sg13g2_dlygate4sd3_1 hold729 (.A(\TRNG.Word_Out[66] ),
    .X(net1857));
 sg13g2_dlygate4sd3_1 hold730 (.A(_01311_),
    .X(net1858));
 sg13g2_dlygate4sd3_1 hold731 (.A(\TRNG.Padded_Out[271] ),
    .X(net1859));
 sg13g2_dlygate4sd3_1 hold732 (.A(_01899_),
    .X(net1860));
 sg13g2_dlygate4sd3_1 hold733 (.A(\TRNG.Padded_Out[112] ),
    .X(net1861));
 sg13g2_dlygate4sd3_1 hold734 (.A(_01740_),
    .X(net1862));
 sg13g2_dlygate4sd3_1 hold735 (.A(\TRNG.Padded_Out[420] ),
    .X(net1863));
 sg13g2_dlygate4sd3_1 hold736 (.A(\TRNG.Word_Out[0] ),
    .X(net1864));
 sg13g2_dlygate4sd3_1 hold737 (.A(_01245_),
    .X(net1865));
 sg13g2_dlygate4sd3_1 hold738 (.A(\TRNG.Word_Out[150] ),
    .X(net1866));
 sg13g2_dlygate4sd3_1 hold739 (.A(_01395_),
    .X(net1867));
 sg13g2_dlygate4sd3_1 hold740 (.A(\TRNG.Padded_Out[425] ),
    .X(net1868));
 sg13g2_dlygate4sd3_1 hold741 (.A(_02053_),
    .X(net1869));
 sg13g2_dlygate4sd3_1 hold742 (.A(\TRNG.Padded_Out[188] ),
    .X(net1870));
 sg13g2_dlygate4sd3_1 hold743 (.A(_01816_),
    .X(net1871));
 sg13g2_dlygate4sd3_1 hold744 (.A(\TRNG.Padded_Out[138] ),
    .X(net1872));
 sg13g2_dlygate4sd3_1 hold745 (.A(_01766_),
    .X(net1873));
 sg13g2_dlygate4sd3_1 hold746 (.A(\TRNG.Word_Out[405] ),
    .X(net1874));
 sg13g2_dlygate4sd3_1 hold747 (.A(_01650_),
    .X(net1875));
 sg13g2_dlygate4sd3_1 hold748 (.A(\TRNG.Padded_Out[293] ),
    .X(net1876));
 sg13g2_dlygate4sd3_1 hold749 (.A(\TRNG.Padded_Out[250] ),
    .X(net1877));
 sg13g2_dlygate4sd3_1 hold750 (.A(_01878_),
    .X(net1878));
 sg13g2_dlygate4sd3_1 hold751 (.A(\TRNG.Word_Out[100] ),
    .X(net1879));
 sg13g2_dlygate4sd3_1 hold752 (.A(_01345_),
    .X(net1880));
 sg13g2_dlygate4sd3_1 hold753 (.A(\TRNG.Padded_Out[393] ),
    .X(net1881));
 sg13g2_dlygate4sd3_1 hold754 (.A(_02021_),
    .X(net1882));
 sg13g2_dlygate4sd3_1 hold755 (.A(\TRNG.Padded_Out[465] ),
    .X(net1883));
 sg13g2_dlygate4sd3_1 hold756 (.A(\TRNG.Padded_Out[81] ),
    .X(net1884));
 sg13g2_dlygate4sd3_1 hold757 (.A(_01709_),
    .X(net1885));
 sg13g2_dlygate4sd3_1 hold758 (.A(\TRNG.sha256.expand.exp_ctrl.sum[20] ),
    .X(net1886));
 sg13g2_dlygate4sd3_1 hold759 (.A(_01007_),
    .X(net1887));
 sg13g2_dlygate4sd3_1 hold760 (.A(\TRNG.Padded_Out[477] ),
    .X(net1888));
 sg13g2_dlygate4sd3_1 hold761 (.A(_02105_),
    .X(net1889));
 sg13g2_dlygate4sd3_1 hold762 (.A(\TRNG.Padded_Out[192] ),
    .X(net1890));
 sg13g2_dlygate4sd3_1 hold763 (.A(\TRNG.Word_Out[208] ),
    .X(net1891));
 sg13g2_dlygate4sd3_1 hold764 (.A(_01453_),
    .X(net1892));
 sg13g2_dlygate4sd3_1 hold765 (.A(\TRNG.Padded_Out[165] ),
    .X(net1893));
 sg13g2_dlygate4sd3_1 hold766 (.A(\TRNG.Padded_Out[156] ),
    .X(net1894));
 sg13g2_dlygate4sd3_1 hold767 (.A(_01784_),
    .X(net1895));
 sg13g2_dlygate4sd3_1 hold768 (.A(\TRNG.uart_tx_inst.tx_bit_counter[3] ),
    .X(net1896));
 sg13g2_dlygate4sd3_1 hold769 (.A(_00309_),
    .X(net1897));
 sg13g2_dlygate4sd3_1 hold770 (.A(\TRNG.Padded_Out[282] ),
    .X(net1898));
 sg13g2_dlygate4sd3_1 hold771 (.A(_01910_),
    .X(net1899));
 sg13g2_dlygate4sd3_1 hold772 (.A(\TRNG.Padded_Out[95] ),
    .X(net1900));
 sg13g2_dlygate4sd3_1 hold773 (.A(\TRNG.Padded_Out[424] ),
    .X(net1901));
 sg13g2_dlygate4sd3_1 hold774 (.A(\TRNG.Padded_Out[407] ),
    .X(net1902));
 sg13g2_dlygate4sd3_1 hold775 (.A(_02035_),
    .X(net1903));
 sg13g2_dlygate4sd3_1 hold776 (.A(\TRNG.Word_Out[215] ),
    .X(net1904));
 sg13g2_dlygate4sd3_1 hold777 (.A(_01460_),
    .X(net1905));
 sg13g2_dlygate4sd3_1 hold778 (.A(\TRNG.Padded_Out[286] ),
    .X(net1906));
 sg13g2_dlygate4sd3_1 hold779 (.A(_01914_),
    .X(net1907));
 sg13g2_dlygate4sd3_1 hold780 (.A(\TRNG.Padded_Out[312] ),
    .X(net1908));
 sg13g2_dlygate4sd3_1 hold781 (.A(\TRNG.Padded_Out[352] ),
    .X(net1909));
 sg13g2_dlygate4sd3_1 hold782 (.A(_01980_),
    .X(net1910));
 sg13g2_dlygate4sd3_1 hold783 (.A(\TRNG.Word_Out[295] ),
    .X(net1911));
 sg13g2_dlygate4sd3_1 hold784 (.A(_01540_),
    .X(net1912));
 sg13g2_dlygate4sd3_1 hold785 (.A(\TRNG.Word_Out[434] ),
    .X(net1913));
 sg13g2_dlygate4sd3_1 hold786 (.A(\TRNG.Padded_Out[247] ),
    .X(net1914));
 sg13g2_dlygate4sd3_1 hold787 (.A(_01875_),
    .X(net1915));
 sg13g2_dlygate4sd3_1 hold788 (.A(\TRNG.Word_Out[328] ),
    .X(net1916));
 sg13g2_dlygate4sd3_1 hold789 (.A(_01573_),
    .X(net1917));
 sg13g2_dlygate4sd3_1 hold790 (.A(\TRNG.Padded_Out[405] ),
    .X(net1918));
 sg13g2_dlygate4sd3_1 hold791 (.A(_02033_),
    .X(net1919));
 sg13g2_dlygate4sd3_1 hold792 (.A(\TRNG.Word_Out[259] ),
    .X(net1920));
 sg13g2_dlygate4sd3_1 hold793 (.A(\TRNG.Word_Out[151] ),
    .X(net1921));
 sg13g2_dlygate4sd3_1 hold794 (.A(_01396_),
    .X(net1922));
 sg13g2_dlygate4sd3_1 hold795 (.A(\TRNG.Padded_Out[353] ),
    .X(net1923));
 sg13g2_dlygate4sd3_1 hold796 (.A(_01981_),
    .X(net1924));
 sg13g2_dlygate4sd3_1 hold797 (.A(\TRNG.Padded_Out[322] ),
    .X(net1925));
 sg13g2_dlygate4sd3_1 hold798 (.A(_01950_),
    .X(net1926));
 sg13g2_dlygate4sd3_1 hold799 (.A(\TRNG.Word_Out[128] ),
    .X(net1927));
 sg13g2_dlygate4sd3_1 hold800 (.A(_01373_),
    .X(net1928));
 sg13g2_dlygate4sd3_1 hold801 (.A(\TRNG.Padded_Out[423] ),
    .X(net1929));
 sg13g2_dlygate4sd3_1 hold802 (.A(_02051_),
    .X(net1930));
 sg13g2_dlygate4sd3_1 hold803 (.A(\TRNG.sha256.expand.exp_ctrl.sum[29] ),
    .X(net1931));
 sg13g2_dlygate4sd3_1 hold804 (.A(_01016_),
    .X(net1932));
 sg13g2_dlygate4sd3_1 hold805 (.A(\TRNG.Padded_Out[124] ),
    .X(net1933));
 sg13g2_dlygate4sd3_1 hold806 (.A(_01752_),
    .X(net1934));
 sg13g2_dlygate4sd3_1 hold807 (.A(\TRNG.Word_Out[283] ),
    .X(net1935));
 sg13g2_dlygate4sd3_1 hold808 (.A(_01528_),
    .X(net1936));
 sg13g2_dlygate4sd3_1 hold809 (.A(\TRNG.Word_Out[4] ),
    .X(net1937));
 sg13g2_dlygate4sd3_1 hold810 (.A(_01249_),
    .X(net1938));
 sg13g2_dlygate4sd3_1 hold811 (.A(\TRNG.Padded_Out[205] ),
    .X(net1939));
 sg13g2_dlygate4sd3_1 hold812 (.A(_01833_),
    .X(net1940));
 sg13g2_dlygate4sd3_1 hold813 (.A(\TRNG.Word_Out[53] ),
    .X(net1941));
 sg13g2_dlygate4sd3_1 hold814 (.A(_01298_),
    .X(net1942));
 sg13g2_dlygate4sd3_1 hold815 (.A(\TRNG.Word_Out[79] ),
    .X(net1943));
 sg13g2_dlygate4sd3_1 hold816 (.A(_01324_),
    .X(net1944));
 sg13g2_dlygate4sd3_1 hold817 (.A(\TRNG.Padded_Out[150] ),
    .X(net1945));
 sg13g2_dlygate4sd3_1 hold818 (.A(_01778_),
    .X(net1946));
 sg13g2_dlygate4sd3_1 hold819 (.A(\TRNG.Word_Out[222] ),
    .X(net1947));
 sg13g2_dlygate4sd3_1 hold820 (.A(_01467_),
    .X(net1948));
 sg13g2_dlygate4sd3_1 hold821 (.A(\TRNG.Padded_Out[118] ),
    .X(net1949));
 sg13g2_dlygate4sd3_1 hold822 (.A(\TRNG.Padded_Out[66] ),
    .X(net1950));
 sg13g2_dlygate4sd3_1 hold823 (.A(_01694_),
    .X(net1951));
 sg13g2_dlygate4sd3_1 hold824 (.A(\TRNG.Padded_Out[76] ),
    .X(net1952));
 sg13g2_dlygate4sd3_1 hold825 (.A(_01704_),
    .X(net1953));
 sg13g2_dlygate4sd3_1 hold826 (.A(\TRNG.Word_Out[185] ),
    .X(net1954));
 sg13g2_dlygate4sd3_1 hold827 (.A(_01430_),
    .X(net1955));
 sg13g2_dlygate4sd3_1 hold828 (.A(\TRNG.Word_Out[227] ),
    .X(net1956));
 sg13g2_dlygate4sd3_1 hold829 (.A(\TRNG.Padded_Out[99] ),
    .X(net1957));
 sg13g2_dlygate4sd3_1 hold830 (.A(_01727_),
    .X(net1958));
 sg13g2_dlygate4sd3_1 hold831 (.A(\TRNG.Word_Out[317] ),
    .X(net1959));
 sg13g2_dlygate4sd3_1 hold832 (.A(\TRNG.Word_Out[158] ),
    .X(net1960));
 sg13g2_dlygate4sd3_1 hold833 (.A(_01403_),
    .X(net1961));
 sg13g2_dlygate4sd3_1 hold834 (.A(\TRNG.Word_Out[195] ),
    .X(net1962));
 sg13g2_dlygate4sd3_1 hold835 (.A(_01440_),
    .X(net1963));
 sg13g2_dlygate4sd3_1 hold836 (.A(\TRNG.Word_Out[110] ),
    .X(net1964));
 sg13g2_dlygate4sd3_1 hold837 (.A(\TRNG.Padded_Out[215] ),
    .X(net1965));
 sg13g2_dlygate4sd3_1 hold838 (.A(\TRNG.Padded_Out[311] ),
    .X(net1966));
 sg13g2_dlygate4sd3_1 hold839 (.A(_01939_),
    .X(net1967));
 sg13g2_dlygate4sd3_1 hold840 (.A(\TRNG.Padded_Out[325] ),
    .X(net1968));
 sg13g2_dlygate4sd3_1 hold841 (.A(\TRNG.Padded_Out[266] ),
    .X(net1969));
 sg13g2_dlygate4sd3_1 hold842 (.A(_01894_),
    .X(net1970));
 sg13g2_dlygate4sd3_1 hold843 (.A(\TRNG.Padded_Out[304] ),
    .X(net1971));
 sg13g2_dlygate4sd3_1 hold844 (.A(_01932_),
    .X(net1972));
 sg13g2_dlygate4sd3_1 hold845 (.A(\TRNG.Word_Out[209] ),
    .X(net1973));
 sg13g2_dlygate4sd3_1 hold846 (.A(_01454_),
    .X(net1974));
 sg13g2_dlygate4sd3_1 hold847 (.A(\TRNG.Padded_Out[126] ),
    .X(net1975));
 sg13g2_dlygate4sd3_1 hold848 (.A(_01754_),
    .X(net1976));
 sg13g2_dlygate4sd3_1 hold849 (.A(\TRNG.Padded_Out[453] ),
    .X(net1977));
 sg13g2_dlygate4sd3_1 hold850 (.A(\TRNG.Word_Out[17] ),
    .X(net1978));
 sg13g2_dlygate4sd3_1 hold851 (.A(_01262_),
    .X(net1979));
 sg13g2_dlygate4sd3_1 hold852 (.A(\TRNG.Padded_Out[483] ),
    .X(net1980));
 sg13g2_dlygate4sd3_1 hold853 (.A(_02111_),
    .X(net1981));
 sg13g2_dlygate4sd3_1 hold854 (.A(\TRNG.Word_Out[363] ),
    .X(net1982));
 sg13g2_dlygate4sd3_1 hold855 (.A(_01608_),
    .X(net1983));
 sg13g2_dlygate4sd3_1 hold856 (.A(\TRNG.Word_Out[16] ),
    .X(net1984));
 sg13g2_dlygate4sd3_1 hold857 (.A(\TRNG.Word_Out[369] ),
    .X(net1985));
 sg13g2_dlygate4sd3_1 hold858 (.A(_01614_),
    .X(net1986));
 sg13g2_dlygate4sd3_1 hold859 (.A(\TRNG.Padded_Out[385] ),
    .X(net1987));
 sg13g2_dlygate4sd3_1 hold860 (.A(_02013_),
    .X(net1988));
 sg13g2_dlygate4sd3_1 hold861 (.A(\TRNG.Padded_Out[77] ),
    .X(net1989));
 sg13g2_dlygate4sd3_1 hold862 (.A(_01705_),
    .X(net1990));
 sg13g2_dlygate4sd3_1 hold863 (.A(\TRNG.Word_Out[358] ),
    .X(net1991));
 sg13g2_dlygate4sd3_1 hold864 (.A(\TRNG.Padded_Out[430] ),
    .X(net1992));
 sg13g2_dlygate4sd3_1 hold865 (.A(_02058_),
    .X(net1993));
 sg13g2_dlygate4sd3_1 hold866 (.A(\TRNG.Word_Out[218] ),
    .X(net1994));
 sg13g2_dlygate4sd3_1 hold867 (.A(_01463_),
    .X(net1995));
 sg13g2_dlygate4sd3_1 hold868 (.A(\TRNG.Padded_Out[173] ),
    .X(net1996));
 sg13g2_dlygate4sd3_1 hold869 (.A(_01801_),
    .X(net1997));
 sg13g2_dlygate4sd3_1 hold870 (.A(\TRNG.Word_Out[270] ),
    .X(net1998));
 sg13g2_dlygate4sd3_1 hold871 (.A(_01515_),
    .X(net1999));
 sg13g2_dlygate4sd3_1 hold872 (.A(\TRNG.Padded_Out[255] ),
    .X(net2000));
 sg13g2_dlygate4sd3_1 hold873 (.A(_01883_),
    .X(net2001));
 sg13g2_dlygate4sd3_1 hold874 (.A(\TRNG.Word_Out[398] ),
    .X(net2002));
 sg13g2_dlygate4sd3_1 hold875 (.A(_01643_),
    .X(net2003));
 sg13g2_dlygate4sd3_1 hold876 (.A(\TRNG.Padded_Out[158] ),
    .X(net2004));
 sg13g2_dlygate4sd3_1 hold877 (.A(\TRNG.Word_Out[206] ),
    .X(net2005));
 sg13g2_dlygate4sd3_1 hold878 (.A(_01451_),
    .X(net2006));
 sg13g2_dlygate4sd3_1 hold879 (.A(\TRNG.Padded_Out[221] ),
    .X(net2007));
 sg13g2_dlygate4sd3_1 hold880 (.A(_01849_),
    .X(net2008));
 sg13g2_dlygate4sd3_1 hold881 (.A(\TRNG.Padded_Out[228] ),
    .X(net2009));
 sg13g2_dlygate4sd3_1 hold882 (.A(\TRNG.Padded_Out[381] ),
    .X(net2010));
 sg13g2_dlygate4sd3_1 hold883 (.A(_02009_),
    .X(net2011));
 sg13g2_dlygate4sd3_1 hold884 (.A(\TRNG.Padded_Out[166] ),
    .X(net2012));
 sg13g2_dlygate4sd3_1 hold885 (.A(_01794_),
    .X(net2013));
 sg13g2_dlygate4sd3_1 hold886 (.A(\TRNG.Word_Out[118] ),
    .X(net2014));
 sg13g2_dlygate4sd3_1 hold887 (.A(_01363_),
    .X(net2015));
 sg13g2_dlygate4sd3_1 hold888 (.A(\TRNG.Padded_Out[388] ),
    .X(net2016));
 sg13g2_dlygate4sd3_1 hold889 (.A(\TRNG.Word_Out[217] ),
    .X(net2017));
 sg13g2_dlygate4sd3_1 hold890 (.A(\TRNG.Padded_Out[406] ),
    .X(net2018));
 sg13g2_dlygate4sd3_1 hold891 (.A(_02034_),
    .X(net2019));
 sg13g2_dlygate4sd3_1 hold892 (.A(\TRNG.Padded_Out[452] ),
    .X(net2020));
 sg13g2_dlygate4sd3_1 hold893 (.A(\TRNG.Padded_Out[240] ),
    .X(net2021));
 sg13g2_dlygate4sd3_1 hold894 (.A(_01868_),
    .X(net2022));
 sg13g2_dlygate4sd3_1 hold895 (.A(\TRNG.Padded_Out[254] ),
    .X(net2023));
 sg13g2_dlygate4sd3_1 hold896 (.A(\TRNG.Word_Out[423] ),
    .X(net2024));
 sg13g2_dlygate4sd3_1 hold897 (.A(_01668_),
    .X(net2025));
 sg13g2_dlygate4sd3_1 hold898 (.A(\TRNG.Word_Out[438] ),
    .X(net2026));
 sg13g2_dlygate4sd3_1 hold899 (.A(_01683_),
    .X(net2027));
 sg13g2_dlygate4sd3_1 hold900 (.A(\TRNG.Padded_Out[230] ),
    .X(net2028));
 sg13g2_dlygate4sd3_1 hold901 (.A(_01858_),
    .X(net2029));
 sg13g2_dlygate4sd3_1 hold902 (.A(\TRNG.Word_Out[415] ),
    .X(net2030));
 sg13g2_dlygate4sd3_1 hold903 (.A(_01660_),
    .X(net2031));
 sg13g2_dlygate4sd3_1 hold904 (.A(\TRNG.Word_Out[105] ),
    .X(net2032));
 sg13g2_dlygate4sd3_1 hold905 (.A(_01350_),
    .X(net2033));
 sg13g2_dlygate4sd3_1 hold906 (.A(\TRNG.Word_Out[309] ),
    .X(net2034));
 sg13g2_dlygate4sd3_1 hold907 (.A(_01554_),
    .X(net2035));
 sg13g2_dlygate4sd3_1 hold908 (.A(\TRNG.Padded_Out[238] ),
    .X(net2036));
 sg13g2_dlygate4sd3_1 hold909 (.A(_01866_),
    .X(net2037));
 sg13g2_dlygate4sd3_1 hold910 (.A(\TRNG.sha256.expand.exp_ctrl.sum[5] ),
    .X(net2038));
 sg13g2_dlygate4sd3_1 hold911 (.A(_00992_),
    .X(net2039));
 sg13g2_dlygate4sd3_1 hold912 (.A(\TRNG.Padded_Out[203] ),
    .X(net2040));
 sg13g2_dlygate4sd3_1 hold913 (.A(\TRNG.Padded_Out[135] ),
    .X(net2041));
 sg13g2_dlygate4sd3_1 hold914 (.A(\TRNG.Padded_Out[310] ),
    .X(net2042));
 sg13g2_dlygate4sd3_1 hold915 (.A(_01938_),
    .X(net2043));
 sg13g2_dlygate4sd3_1 hold916 (.A(\TRNG.Padded_Out[305] ),
    .X(net2044));
 sg13g2_dlygate4sd3_1 hold917 (.A(\TRNG.Padded_Out[343] ),
    .X(net2045));
 sg13g2_dlygate4sd3_1 hold918 (.A(_01971_),
    .X(net2046));
 sg13g2_dlygate4sd3_1 hold919 (.A(\TRNG.Padded_Out[101] ),
    .X(net2047));
 sg13g2_dlygate4sd3_1 hold920 (.A(\TRNG.Padded_Out[187] ),
    .X(net2048));
 sg13g2_dlygate4sd3_1 hold921 (.A(_01815_),
    .X(net2049));
 sg13g2_dlygate4sd3_1 hold922 (.A(\TRNG.Padded_Out[98] ),
    .X(net2050));
 sg13g2_dlygate4sd3_1 hold923 (.A(_01726_),
    .X(net2051));
 sg13g2_dlygate4sd3_1 hold924 (.A(\TRNG.Padded_Out[209] ),
    .X(net2052));
 sg13g2_dlygate4sd3_1 hold925 (.A(_01837_),
    .X(net2053));
 sg13g2_dlygate4sd3_1 hold926 (.A(\TRNG.Word_Out[181] ),
    .X(net2054));
 sg13g2_dlygate4sd3_1 hold927 (.A(_01426_),
    .X(net2055));
 sg13g2_dlygate4sd3_1 hold928 (.A(\TRNG.Padded_Out[157] ),
    .X(net2056));
 sg13g2_dlygate4sd3_1 hold929 (.A(_01785_),
    .X(net2057));
 sg13g2_dlygate4sd3_1 hold930 (.A(\TRNG.Word_Out[95] ),
    .X(net2058));
 sg13g2_dlygate4sd3_1 hold931 (.A(_01340_),
    .X(net2059));
 sg13g2_dlygate4sd3_1 hold932 (.A(\TRNG.Padded_Out[448] ),
    .X(net2060));
 sg13g2_dlygate4sd3_1 hold933 (.A(_02076_),
    .X(net2061));
 sg13g2_dlygate4sd3_1 hold934 (.A(\TRNG.Padded_Out[129] ),
    .X(net2062));
 sg13g2_dlygate4sd3_1 hold935 (.A(_01757_),
    .X(net2063));
 sg13g2_dlygate4sd3_1 hold936 (.A(\TRNG.sha256.expand.exp_ctrl.j_2[3] ),
    .X(net2064));
 sg13g2_dlygate4sd3_1 hold937 (.A(_00978_),
    .X(net2065));
 sg13g2_dlygate4sd3_1 hold938 (.A(\TRNG.Padded_Out[91] ),
    .X(net2066));
 sg13g2_dlygate4sd3_1 hold939 (.A(_01719_),
    .X(net2067));
 sg13g2_dlygate4sd3_1 hold940 (.A(\TRNG.Padded_Out[341] ),
    .X(net2068));
 sg13g2_dlygate4sd3_1 hold941 (.A(_01969_),
    .X(net2069));
 sg13g2_dlygate4sd3_1 hold942 (.A(\TRNG.Word_Out[122] ),
    .X(net2070));
 sg13g2_dlygate4sd3_1 hold943 (.A(\TRNG.Word_Out[353] ),
    .X(net2071));
 sg13g2_dlygate4sd3_1 hold944 (.A(_01598_),
    .X(net2072));
 sg13g2_dlygate4sd3_1 hold945 (.A(\TRNG.Padded_Out[125] ),
    .X(net2073));
 sg13g2_dlygate4sd3_1 hold946 (.A(\TRNG.Padded_Out[360] ),
    .X(net2074));
 sg13g2_dlygate4sd3_1 hold947 (.A(\TRNG.Word_Out[97] ),
    .X(net2075));
 sg13g2_dlygate4sd3_1 hold948 (.A(\TRNG.Word_Out[350] ),
    .X(net2076));
 sg13g2_dlygate4sd3_1 hold949 (.A(_01595_),
    .X(net2077));
 sg13g2_dlygate4sd3_1 hold950 (.A(\TRNG.Word_Out[375] ),
    .X(net2078));
 sg13g2_dlygate4sd3_1 hold951 (.A(\TRNG.Padded_Out[191] ),
    .X(net2079));
 sg13g2_dlygate4sd3_1 hold952 (.A(_01819_),
    .X(net2080));
 sg13g2_dlygate4sd3_1 hold953 (.A(\TRNG.Word_Out[272] ),
    .X(net2081));
 sg13g2_dlygate4sd3_1 hold954 (.A(_01517_),
    .X(net2082));
 sg13g2_dlygate4sd3_1 hold955 (.A(\TRNG.Word_Out[190] ),
    .X(net2083));
 sg13g2_dlygate4sd3_1 hold956 (.A(_01435_),
    .X(net2084));
 sg13g2_dlygate4sd3_1 hold957 (.A(\TRNG.Padded_Out[96] ),
    .X(net2085));
 sg13g2_dlygate4sd3_1 hold958 (.A(_01724_),
    .X(net2086));
 sg13g2_dlygate4sd3_1 hold959 (.A(\TRNG.Word_Out[352] ),
    .X(net2087));
 sg13g2_dlygate4sd3_1 hold960 (.A(\TRNG.Padded_Out[108] ),
    .X(net2088));
 sg13g2_dlygate4sd3_1 hold961 (.A(_01736_),
    .X(net2089));
 sg13g2_dlygate4sd3_1 hold962 (.A(\TRNG.Padded_Out[174] ),
    .X(net2090));
 sg13g2_dlygate4sd3_1 hold963 (.A(_01802_),
    .X(net2091));
 sg13g2_dlygate4sd3_1 hold964 (.A(\TRNG.Padded_Out[224] ),
    .X(net2092));
 sg13g2_dlygate4sd3_1 hold965 (.A(_01852_),
    .X(net2093));
 sg13g2_dlygate4sd3_1 hold966 (.A(\TRNG.Word_Out[238] ),
    .X(net2094));
 sg13g2_dlygate4sd3_1 hold967 (.A(_01483_),
    .X(net2095));
 sg13g2_dlygate4sd3_1 hold968 (.A(\TRNG.Padded_Out[470] ),
    .X(net2096));
 sg13g2_dlygate4sd3_1 hold969 (.A(\TRNG.Padded_Out[450] ),
    .X(net2097));
 sg13g2_dlygate4sd3_1 hold970 (.A(_02078_),
    .X(net2098));
 sg13g2_dlygate4sd3_1 hold971 (.A(\TRNG.Word_Out[80] ),
    .X(net2099));
 sg13g2_dlygate4sd3_1 hold972 (.A(_01325_),
    .X(net2100));
 sg13g2_dlygate4sd3_1 hold973 (.A(\TRNG.Word_Out[334] ),
    .X(net2101));
 sg13g2_dlygate4sd3_1 hold974 (.A(_01579_),
    .X(net2102));
 sg13g2_dlygate4sd3_1 hold975 (.A(\TRNG.Word_Out[177] ),
    .X(net2103));
 sg13g2_dlygate4sd3_1 hold976 (.A(_01422_),
    .X(net2104));
 sg13g2_dlygate4sd3_1 hold977 (.A(\TRNG.Word_Out[205] ),
    .X(net2105));
 sg13g2_dlygate4sd3_1 hold978 (.A(\TRNG.Word_Out[62] ),
    .X(net2106));
 sg13g2_dlygate4sd3_1 hold979 (.A(\TRNG.Padded_Out[103] ),
    .X(net2107));
 sg13g2_dlygate4sd3_1 hold980 (.A(\TRNG.Word_Out[50] ),
    .X(net2108));
 sg13g2_dlygate4sd3_1 hold981 (.A(_01295_),
    .X(net2109));
 sg13g2_dlygate4sd3_1 hold982 (.A(\TRNG.Padded_Out[178] ),
    .X(net2110));
 sg13g2_dlygate4sd3_1 hold983 (.A(\TRNG.Padded_Out[303] ),
    .X(net2111));
 sg13g2_dlygate4sd3_1 hold984 (.A(\TRNG.Word_Out[45] ),
    .X(net2112));
 sg13g2_dlygate4sd3_1 hold985 (.A(\TRNG.Word_Out[35] ),
    .X(net2113));
 sg13g2_dlygate4sd3_1 hold986 (.A(\TRNG.Word_Out[210] ),
    .X(net2114));
 sg13g2_dlygate4sd3_1 hold987 (.A(_01455_),
    .X(net2115));
 sg13g2_dlygate4sd3_1 hold988 (.A(\TRNG.Word_Out[441] ),
    .X(net2116));
 sg13g2_dlygate4sd3_1 hold989 (.A(_01686_),
    .X(net2117));
 sg13g2_dlygate4sd3_1 hold990 (.A(\TRNG.Word_Out[137] ),
    .X(net2118));
 sg13g2_dlygate4sd3_1 hold991 (.A(\TRNG.Padded_Out[104] ),
    .X(net2119));
 sg13g2_dlygate4sd3_1 hold992 (.A(_01732_),
    .X(net2120));
 sg13g2_dlygate4sd3_1 hold993 (.A(\TRNG.Word_Out[297] ),
    .X(net2121));
 sg13g2_dlygate4sd3_1 hold994 (.A(_01542_),
    .X(net2122));
 sg13g2_dlygate4sd3_1 hold995 (.A(\TRNG.Word_Out[67] ),
    .X(net2123));
 sg13g2_dlygate4sd3_1 hold996 (.A(_01312_),
    .X(net2124));
 sg13g2_dlygate4sd3_1 hold997 (.A(\TRNG.Padded_Out[345] ),
    .X(net2125));
 sg13g2_dlygate4sd3_1 hold998 (.A(\TRNG.Padded_Out[298] ),
    .X(net2126));
 sg13g2_dlygate4sd3_1 hold999 (.A(_01926_),
    .X(net2127));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\TRNG.Word_Out[368] ),
    .X(net2128));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\TRNG.Word_Out[22] ),
    .X(net2129));
 sg13g2_dlygate4sd3_1 hold1002 (.A(_01267_),
    .X(net2130));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\TRNG.Padded_Out[110] ),
    .X(net2131));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\TRNG.Word_Out[431] ),
    .X(net2132));
 sg13g2_dlygate4sd3_1 hold1005 (.A(_01676_),
    .X(net2133));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\TRNG.sha256.expand.exp_ctrl.sum[27] ),
    .X(net2134));
 sg13g2_dlygate4sd3_1 hold1007 (.A(_01014_),
    .X(net2135));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\TRNG.Word_Out[310] ),
    .X(net2136));
 sg13g2_dlygate4sd3_1 hold1009 (.A(_01555_),
    .X(net2137));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\TRNG.Padded_Out[283] ),
    .X(net2138));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\TRNG.Word_Out[365] ),
    .X(net2139));
 sg13g2_dlygate4sd3_1 hold1012 (.A(_01610_),
    .X(net2140));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\TRNG.Padded_Out[357] ),
    .X(net2141));
 sg13g2_dlygate4sd3_1 hold1014 (.A(_01985_),
    .X(net2142));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\TRNG.Word_Out[437] ),
    .X(net2143));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\TRNG.Padded_Out[223] ),
    .X(net2144));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\TRNG.Padded_Out[288] ),
    .X(net2145));
 sg13g2_dlygate4sd3_1 hold1018 (.A(_01916_),
    .X(net2146));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\TRNG.Padded_Out[475] ),
    .X(net2147));
 sg13g2_dlygate4sd3_1 hold1020 (.A(_02103_),
    .X(net2148));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\TRNG.Padded_Out[106] ),
    .X(net2149));
 sg13g2_dlygate4sd3_1 hold1022 (.A(_01734_),
    .X(net2150));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\TRNG.Padded_Out[369] ),
    .X(net2151));
 sg13g2_dlygate4sd3_1 hold1024 (.A(_01997_),
    .X(net2152));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\TRNG.Word_Out[74] ),
    .X(net2153));
 sg13g2_dlygate4sd3_1 hold1026 (.A(_01319_),
    .X(net2154));
 sg13g2_dlygate4sd3_1 hold1027 (.A(\TRNG.Padded_Out[269] ),
    .X(net2155));
 sg13g2_dlygate4sd3_1 hold1028 (.A(_01897_),
    .X(net2156));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\TRNG.Word_Out[385] ),
    .X(net2157));
 sg13g2_dlygate4sd3_1 hold1030 (.A(_01630_),
    .X(net2158));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\TRNG.Padded_Out[472] ),
    .X(net2159));
 sg13g2_dlygate4sd3_1 hold1032 (.A(_02100_),
    .X(net2160));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\TRNG.Word_Out[417] ),
    .X(net2161));
 sg13g2_dlygate4sd3_1 hold1034 (.A(_01662_),
    .X(net2162));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\TRNG.Word_Out[443] ),
    .X(net2163));
 sg13g2_dlygate4sd3_1 hold1036 (.A(_01688_),
    .X(net2164));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\TRNG.Word_Out[286] ),
    .X(net2165));
 sg13g2_dlygate4sd3_1 hold1038 (.A(_01531_),
    .X(net2166));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\TRNG.Padded_Out[314] ),
    .X(net2167));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\TRNG.Padded_Out[460] ),
    .X(net2168));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\TRNG.Word_Out[96] ),
    .X(net2169));
 sg13g2_dlygate4sd3_1 hold1042 (.A(\TRNG.Padded_Out[397] ),
    .X(net2170));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\TRNG.Padded_Out[408] ),
    .X(net2171));
 sg13g2_dlygate4sd3_1 hold1044 (.A(_02036_),
    .X(net2172));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\TRNG.Padded_Out[137] ),
    .X(net2173));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\TRNG.Padded_Out[82] ),
    .X(net2174));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\TRNG.Padded_Out[358] ),
    .X(net2175));
 sg13g2_dlygate4sd3_1 hold1048 (.A(_01986_),
    .X(net2176));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\TRNG.Word_Out[271] ),
    .X(net2177));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\TRNG.Word_Out[186] ),
    .X(net2178));
 sg13g2_dlygate4sd3_1 hold1051 (.A(_01431_),
    .X(net2179));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\TRNG.Padded_Out[227] ),
    .X(net2180));
 sg13g2_dlygate4sd3_1 hold1053 (.A(_01855_),
    .X(net2181));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\TRNG.Padded_Out[109] ),
    .X(net2182));
 sg13g2_dlygate4sd3_1 hold1055 (.A(_01737_),
    .X(net2183));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\TRNG.Word_Out[342] ),
    .X(net2184));
 sg13g2_dlygate4sd3_1 hold1057 (.A(_01587_),
    .X(net2185));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\TRNG.Padded_Out[97] ),
    .X(net2186));
 sg13g2_dlygate4sd3_1 hold1059 (.A(_01725_),
    .X(net2187));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\TRNG.Word_Out[264] ),
    .X(net2188));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\TRNG.Word_Out[69] ),
    .X(net2189));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\TRNG.Padded_Out[217] ),
    .X(net2190));
 sg13g2_dlygate4sd3_1 hold1063 (.A(_01845_),
    .X(net2191));
 sg13g2_dlygate4sd3_1 hold1064 (.A(_00128_),
    .X(net2192));
 sg13g2_dlygate4sd3_1 hold1065 (.A(_05912_),
    .X(net2193));
 sg13g2_dlygate4sd3_1 hold1066 (.A(_00104_),
    .X(net2194));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\TRNG.Padded_Out[376] ),
    .X(net2195));
 sg13g2_dlygate4sd3_1 hold1068 (.A(_02004_),
    .X(net2196));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\TRNG.Padded_Out[361] ),
    .X(net2197));
 sg13g2_dlygate4sd3_1 hold1070 (.A(_01989_),
    .X(net2198));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\TRNG.Word_Out[336] ),
    .X(net2199));
 sg13g2_dlygate4sd3_1 hold1072 (.A(_01581_),
    .X(net2200));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\TRNG.Padded_Out[434] ),
    .X(net2201));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\TRNG.Word_Out[90] ),
    .X(net2202));
 sg13g2_dlygate4sd3_1 hold1075 (.A(_01335_),
    .X(net2203));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\TRNG.Word_Out[232] ),
    .X(net2204));
 sg13g2_dlygate4sd3_1 hold1077 (.A(_01477_),
    .X(net2205));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\TRNG.Word_Out[256] ),
    .X(net2206));
 sg13g2_dlygate4sd3_1 hold1079 (.A(_01501_),
    .X(net2207));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\TRNG.Padded_Out[132] ),
    .X(net2208));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\TRNG.sha256.expand.exp_ctrl.sum[9] ),
    .X(net2209));
 sg13g2_dlygate4sd3_1 hold1082 (.A(_00996_),
    .X(net2210));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\TRNG.Word_Out[86] ),
    .X(net2211));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\TRNG.Padded_Out[319] ),
    .X(net2212));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\TRNG.Padded_Out[482] ),
    .X(net2213));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\TRNG.uart_tx_inst.tx_reg[7] ),
    .X(net2214));
 sg13g2_dlygate4sd3_1 hold1087 (.A(_05946_),
    .X(net2215));
 sg13g2_dlygate4sd3_1 hold1088 (.A(_00113_),
    .X(net2216));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\TRNG.Word_Out[445] ),
    .X(net2217));
 sg13g2_dlygate4sd3_1 hold1090 (.A(_01690_),
    .X(net2218));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\TRNG.Word_Out[183] ),
    .X(net2219));
 sg13g2_dlygate4sd3_1 hold1092 (.A(_01428_),
    .X(net2220));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\TRNG.Padded_Out[244] ),
    .X(net2221));
 sg13g2_dlygate4sd3_1 hold1094 (.A(_01872_),
    .X(net2222));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\TRNG.Padded_Out[467] ),
    .X(net2223));
 sg13g2_dlygate4sd3_1 hold1096 (.A(_02095_),
    .X(net2224));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\TRNG.Word_Out[216] ),
    .X(net2225));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\TRNG.sha256.expand.exp_ctrl.sum[7] ),
    .X(net2226));
 sg13g2_dlygate4sd3_1 hold1099 (.A(_00994_),
    .X(net2227));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\TRNG.Word_Out[374] ),
    .X(net2228));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\TRNG.sha256.expand.exp_ctrl.sum[13] ),
    .X(net2229));
 sg13g2_dlygate4sd3_1 hold1102 (.A(_01000_),
    .X(net2230));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\TRNG.Word_Out[424] ),
    .X(net2231));
 sg13g2_dlygate4sd3_1 hold1104 (.A(_01669_),
    .X(net2232));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\TRNG.Word_Out[172] ),
    .X(net2233));
 sg13g2_dlygate4sd3_1 hold1106 (.A(_01417_),
    .X(net2234));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\TRNG.Word_Out[56] ),
    .X(net2235));
 sg13g2_dlygate4sd3_1 hold1108 (.A(_01301_),
    .X(net2236));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\TRNG.Word_Out[302] ),
    .X(net2237));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\TRNG.Word_Out[207] ),
    .X(net2238));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\TRNG.Word_Out[173] ),
    .X(net2239));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\TRNG.Word_Out[116] ),
    .X(net2240));
 sg13g2_dlygate4sd3_1 hold1113 (.A(_01361_),
    .X(net2241));
 sg13g2_dlygate4sd3_1 hold1114 (.A(\TRNG.Word_Out[124] ),
    .X(net2242));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\TRNG.Word_Out[237] ),
    .X(net2243));
 sg13g2_dlygate4sd3_1 hold1116 (.A(\TRNG.Word_Out[52] ),
    .X(net2244));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\TRNG.Word_Out[422] ),
    .X(net2245));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\TRNG.Padded_Out[347] ),
    .X(net2246));
 sg13g2_dlygate4sd3_1 hold1119 (.A(_01975_),
    .X(net2247));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\TRNG.Word_Out[139] ),
    .X(net2248));
 sg13g2_dlygate4sd3_1 hold1121 (.A(_01384_),
    .X(net2249));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\TRNG.Padded_Out[468] ),
    .X(net2250));
 sg13g2_dlygate4sd3_1 hold1123 (.A(_02096_),
    .X(net2251));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\TRNG.Word_Out[199] ),
    .X(net2252));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\TRNG.Word_Out[101] ),
    .X(net2253));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\TRNG.Word_Out[253] ),
    .X(net2254));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\TRNG.Word_Out[314] ),
    .X(net2255));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\TRNG.Padded_Out[440] ),
    .X(net2256));
 sg13g2_dlygate4sd3_1 hold1129 (.A(\TRNG.Padded_Out[242] ),
    .X(net2257));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\TRNG.Padded_Out[229] ),
    .X(net2258));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\TRNG.uart_tx_inst.tx_reg[6] ),
    .X(net2259));
 sg13g2_dlygate4sd3_1 hold1132 (.A(_00112_),
    .X(net2260));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\TRNG.Word_Out[142] ),
    .X(net2261));
 sg13g2_dlygate4sd3_1 hold1134 (.A(_01387_),
    .X(net2262));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\TRNG.Padded_Out[216] ),
    .X(net2263));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\TRNG.Padded_Out[296] ),
    .X(net2264));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\TRNG.sha256.expand.exp_ctrl.sum[2] ),
    .X(net2265));
 sg13g2_dlygate4sd3_1 hold1138 (.A(_00989_),
    .X(net2266));
 sg13g2_dlygate4sd3_1 hold1139 (.A(\TRNG.Word_Out[115] ),
    .X(net2267));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\TRNG.Word_Out[44] ),
    .X(net2268));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\TRNG.sha256.expand.exp_ctrl.sum[18] ),
    .X(net2269));
 sg13g2_dlygate4sd3_1 hold1142 (.A(_01005_),
    .X(net2270));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\TRNG.sha256.expand.exp_ctrl.sum[28] ),
    .X(net2271));
 sg13g2_dlygate4sd3_1 hold1144 (.A(_01015_),
    .X(net2272));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\TRNG.Word_Out[427] ),
    .X(net2273));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\TRNG.Word_Out[234] ),
    .X(net2274));
 sg13g2_dlygate4sd3_1 hold1147 (.A(_01479_),
    .X(net2275));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\TRNG.Padded_Out[318] ),
    .X(net2276));
 sg13g2_dlygate4sd3_1 hold1149 (.A(\TRNG.Padded_Out[307] ),
    .X(net2277));
 sg13g2_dlygate4sd3_1 hold1150 (.A(_01935_),
    .X(net2278));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\TRNG.Word_Out[429] ),
    .X(net2279));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\TRNG.Word_Out[26] ),
    .X(net2280));
 sg13g2_dlygate4sd3_1 hold1153 (.A(_01271_),
    .X(net2281));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\TRNG.Padded_Out[330] ),
    .X(net2282));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\TRNG.Word_Out[230] ),
    .X(net2283));
 sg13g2_dlygate4sd3_1 hold1156 (.A(\TRNG.Word_Out[84] ),
    .X(net2284));
 sg13g2_dlygate4sd3_1 hold1157 (.A(_01329_),
    .X(net2285));
 sg13g2_dlygate4sd3_1 hold1158 (.A(\TRNG.Word_Out[288] ),
    .X(net2286));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\TRNG.Word_Out[123] ),
    .X(net2287));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\TRNG.Word_Out[386] ),
    .X(net2288));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\TRNG.sha256.expand.exp_ctrl.j_7[3] ),
    .X(net2289));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\TRNG.Word_Out[292] ),
    .X(net2290));
 sg13g2_dlygate4sd3_1 hold1163 (.A(_01537_),
    .X(net2291));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\TRNG.Word_Out[344] ),
    .X(net2292));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\TRNG.Padded_Out[493] ),
    .X(net2293));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\TRNG.Word_Out[401] ),
    .X(net2294));
 sg13g2_dlygate4sd3_1 hold1167 (.A(_01646_),
    .X(net2295));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\TRNG.Word_Out[273] ),
    .X(net2296));
 sg13g2_dlygate4sd3_1 hold1169 (.A(_01518_),
    .X(net2297));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\TRNG.Word_Out[433] ),
    .X(net2298));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\TRNG.sha256.expand.exp_ctrl.sum[6] ),
    .X(net2299));
 sg13g2_dlygate4sd3_1 hold1172 (.A(_00993_),
    .X(net2300));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][3] ),
    .X(net2301));
 sg13g2_dlygate4sd3_1 hold1174 (.A(_00660_),
    .X(net2302));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\TRNG.Padded_Out[403] ),
    .X(net2303));
 sg13g2_dlygate4sd3_1 hold1176 (.A(_02031_),
    .X(net2304));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\TRNG.sha256.expand.exp_ctrl.sum[24] ),
    .X(net2305));
 sg13g2_dlygate4sd3_1 hold1178 (.A(_01011_),
    .X(net2306));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\TRNG.sha256.expand.exp_ctrl.sum[4] ),
    .X(net2307));
 sg13g2_dlygate4sd3_1 hold1180 (.A(_00991_),
    .X(net2308));
 sg13g2_dlygate4sd3_1 hold1181 (.A(\TRNG.Padded_Out[469] ),
    .X(net2309));
 sg13g2_dlygate4sd3_1 hold1182 (.A(_02097_),
    .X(net2310));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\TRNG.sha256.expand.exp_ctrl.j_7[0] ),
    .X(net2311));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\TRNG.Repetition_Count_Test.count[1] ),
    .X(net2312));
 sg13g2_dlygate4sd3_1 hold1185 (.A(_00097_),
    .X(net2313));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\TRNG.Padded_Out[92] ),
    .X(net2314));
 sg13g2_dlygate4sd3_1 hold1187 (.A(_01720_),
    .X(net2315));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\TRNG.Word_Out[444] ),
    .X(net2316));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\TRNG.Word_Out[143] ),
    .X(net2317));
 sg13g2_dlygate4sd3_1 hold1190 (.A(_01388_),
    .X(net2318));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\TRNG.Padded_Out[391] ),
    .X(net2319));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\TRNG.Padded_Out[342] ),
    .X(net2320));
 sg13g2_dlygate4sd3_1 hold1193 (.A(_01970_),
    .X(net2321));
 sg13g2_dlygate4sd3_1 hold1194 (.A(_00127_),
    .X(net2322));
 sg13g2_dlygate4sd3_1 hold1195 (.A(_05908_),
    .X(net2323));
 sg13g2_dlygate4sd3_1 hold1196 (.A(_05911_),
    .X(net2324));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\TRNG.uart_tx_inst.tx_reg[4] ),
    .X(net2325));
 sg13g2_dlygate4sd3_1 hold1198 (.A(_05932_),
    .X(net2326));
 sg13g2_dlygate4sd3_1 hold1199 (.A(_00109_),
    .X(net2327));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\TRNG.Padded_Out[329] ),
    .X(net2328));
 sg13g2_dlygate4sd3_1 hold1201 (.A(\TRNG.bit_counter[4] ),
    .X(net2329));
 sg13g2_dlygate4sd3_1 hold1202 (.A(_02152_),
    .X(net2330));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\TRNG.bit_counter[1] ),
    .X(net2331));
 sg13g2_dlygate4sd3_1 hold1204 (.A(_04856_),
    .X(net2332));
 sg13g2_dlygate4sd3_1 hold1205 (.A(_02149_),
    .X(net2333));
 sg13g2_dlygate4sd3_1 hold1206 (.A(\TRNG.uart_tx_inst.tx_reg[3] ),
    .X(net2334));
 sg13g2_dlygate4sd3_1 hold1207 (.A(_05928_),
    .X(net2335));
 sg13g2_dlygate4sd3_1 hold1208 (.A(_00108_),
    .X(net2336));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\TRNG.Padded_Out[211] ),
    .X(net2337));
 sg13g2_dlygate4sd3_1 hold1210 (.A(_01839_),
    .X(net2338));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\TRNG.Word_Out[241] ),
    .X(net2339));
 sg13g2_dlygate4sd3_1 hold1212 (.A(_01486_),
    .X(net2340));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\TRNG.Padded_Out[281] ),
    .X(net2341));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\TRNG.sha256.expand.exp_ctrl.sum[12] ),
    .X(net2342));
 sg13g2_dlygate4sd3_1 hold1215 (.A(_00999_),
    .X(net2343));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\TRNG.sha256.expand.exp_ctrl.sum[23] ),
    .X(net2344));
 sg13g2_dlygate4sd3_1 hold1217 (.A(_01010_),
    .X(net2345));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\TRNG.Word_Out[436] ),
    .X(net2346));
 sg13g2_dlygate4sd3_1 hold1219 (.A(\TRNG.Word_Out[298] ),
    .X(net2347));
 sg13g2_dlygate4sd3_1 hold1220 (.A(_01543_),
    .X(net2348));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\TRNG.Word_Out[305] ),
    .X(net2349));
 sg13g2_dlygate4sd3_1 hold1222 (.A(_01550_),
    .X(net2350));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\TRNG.Word_Out[49] ),
    .X(net2351));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\TRNG.sha256.expand.exp_ctrl.sum[1] ),
    .X(net2352));
 sg13g2_dlygate4sd3_1 hold1225 (.A(_00988_),
    .X(net2353));
 sg13g2_dlygate4sd3_1 hold1226 (.A(\TRNG.Padded_Out[481] ),
    .X(net2354));
 sg13g2_dlygate4sd3_1 hold1227 (.A(_02109_),
    .X(net2355));
 sg13g2_dlygate4sd3_1 hold1228 (.A(\TRNG.Word_Out[315] ),
    .X(net2356));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\TRNG.Padded_Out[509] ),
    .X(net2357));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\TRNG.uart_tx_inst.tx_reg[2] ),
    .X(net2358));
 sg13g2_dlygate4sd3_1 hold1231 (.A(_05924_),
    .X(net2359));
 sg13g2_dlygate4sd3_1 hold1232 (.A(_00107_),
    .X(net2360));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\TRNG.bit_counter[5] ),
    .X(net2361));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\TRNG.Padded_Out[435] ),
    .X(net2362));
 sg13g2_dlygate4sd3_1 hold1235 (.A(_02063_),
    .X(net2363));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\TRNG.Padded_Out[508] ),
    .X(net2364));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\TRNG.Padded_Out[306] ),
    .X(net2365));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\TRNG.Word_Out[220] ),
    .X(net2366));
 sg13g2_dlygate4sd3_1 hold1239 (.A(_01465_),
    .X(net2367));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\TRNG.Repetition_Count_Test.count[2] ),
    .X(net2368));
 sg13g2_dlygate4sd3_1 hold1241 (.A(_00098_),
    .X(net2369));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\TRNG.Word_Out[418] ),
    .X(net2370));
 sg13g2_dlygate4sd3_1 hold1243 (.A(_01663_),
    .X(net2371));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\TRNG.Padded_Out[134] ),
    .X(net2372));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\TRNG.Word_Out[81] ),
    .X(net2373));
 sg13g2_dlygate4sd3_1 hold1246 (.A(_01326_),
    .X(net2374));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\TRNG.ctrl_mode_sync[1] ),
    .X(net2375));
 sg13g2_dlygate4sd3_1 hold1248 (.A(_00270_),
    .X(net2376));
 sg13g2_dlygate4sd3_1 hold1249 (.A(_00983_),
    .X(net2377));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\TRNG.Padded_Out[505] ),
    .X(net2378));
 sg13g2_dlygate4sd3_1 hold1251 (.A(_02133_),
    .X(net2379));
 sg13g2_dlygate4sd3_1 hold1252 (.A(\TRNG.Word_Out[278] ),
    .X(net2380));
 sg13g2_dlygate4sd3_1 hold1253 (.A(_01523_),
    .X(net2381));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\TRNG.Word_Out[287] ),
    .X(net2382));
 sg13g2_dlygate4sd3_1 hold1255 (.A(\TRNG.Word_Out[235] ),
    .X(net2383));
 sg13g2_dlygate4sd3_1 hold1256 (.A(_01480_),
    .X(net2384));
 sg13g2_dlygate4sd3_1 hold1257 (.A(\TRNG.uart_tx_inst.ticks_counter[1] ),
    .X(net2385));
 sg13g2_dlygate4sd3_1 hold1258 (.A(_08841_),
    .X(net2386));
 sg13g2_dlygate4sd3_1 hold1259 (.A(_00857_),
    .X(net2387));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\TRNG.sha256.expand.exp_ctrl.j_7[1] ),
    .X(net2388));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\TRNG.Padded_Out[89] ),
    .X(net2389));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\TRNG.Padded_Out[94] ),
    .X(net2390));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\TRNG.Word_Out[414] ),
    .X(net2391));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\TRNG.sha256.expand.exp_ctrl.sum[16] ),
    .X(net2392));
 sg13g2_dlygate4sd3_1 hold1265 (.A(_01003_),
    .X(net2393));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\TRNG.sha256.expand.exp_ctrl.sum[19] ),
    .X(net2394));
 sg13g2_dlygate4sd3_1 hold1267 (.A(_01006_),
    .X(net2395));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\TRNG.Word_Out[147] ),
    .X(net2396));
 sg13g2_dlygate4sd3_1 hold1269 (.A(_01392_),
    .X(net2397));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\TRNG.Word_Out[257] ),
    .X(net2398));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\TRNG.Padded_Out[478] ),
    .X(net2399));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\TRNG.uart_tx_inst.ticks_counter[6] ),
    .X(net2400));
 sg13g2_dlygate4sd3_1 hold1273 (.A(_08850_),
    .X(net2401));
 sg13g2_dlygate4sd3_1 hold1274 (.A(_00862_),
    .X(net2402));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\TRNG.sha256.expand.exp_ctrl.sum[3] ),
    .X(net2403));
 sg13g2_dlygate4sd3_1 hold1276 (.A(_00990_),
    .X(net2404));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\TRNG.Word_Out[170] ),
    .X(net2405));
 sg13g2_dlygate4sd3_1 hold1278 (.A(_01415_),
    .X(net2406));
 sg13g2_dlygate4sd3_1 hold1279 (.A(\TRNG.Word_Out[219] ),
    .X(net2407));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\TRNG.Word_Out[159] ),
    .X(net2408));
 sg13g2_dlygate4sd3_1 hold1281 (.A(_01404_),
    .X(net2409));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\TRNG.Word_Out[161] ),
    .X(net2410));
 sg13g2_dlygate4sd3_1 hold1283 (.A(_01406_),
    .X(net2411));
 sg13g2_dlygate4sd3_1 hold1284 (.A(\TRNG.Padded_Out[262] ),
    .X(net2412));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][3] ),
    .X(net2413));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\TRNG.Word_Out[373] ),
    .X(net2414));
 sg13g2_dlygate4sd3_1 hold1287 (.A(\TRNG.sha256.expand.exp_ctrl.sum[8] ),
    .X(net2415));
 sg13g2_dlygate4sd3_1 hold1288 (.A(_00995_),
    .X(net2416));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\TRNG.Word_Out[196] ),
    .X(net2417));
 sg13g2_dlygate4sd3_1 hold1290 (.A(\TRNG.sha256.expand.data1_to_ram[18] ),
    .X(net2418));
 sg13g2_dlygate4sd3_1 hold1291 (.A(_02356_),
    .X(net2419));
 sg13g2_dlygate4sd3_1 hold1292 (.A(\TRNG.Padded_Out[136] ),
    .X(net2420));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\TRNG.Word_Out[421] ),
    .X(net2421));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\TRNG.Word_Out[152] ),
    .X(net2422));
 sg13g2_dlygate4sd3_1 hold1295 (.A(_01397_),
    .X(net2423));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\TRNG.Word_Out[279] ),
    .X(net2424));
 sg13g2_dlygate4sd3_1 hold1297 (.A(\TRNG.Word_Out[245] ),
    .X(net2425));
 sg13g2_dlygate4sd3_1 hold1298 (.A(_01490_),
    .X(net2426));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\TRNG.Word_Out[187] ),
    .X(net2427));
 sg13g2_dlygate4sd3_1 hold1300 (.A(_01432_),
    .X(net2428));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\TRNG.Word_Out[171] ),
    .X(net2429));
 sg13g2_dlygate4sd3_1 hold1302 (.A(\TRNG.Padded_Out[193] ),
    .X(net2430));
 sg13g2_dlygate4sd3_1 hold1303 (.A(\TRNG.Word_Out[251] ),
    .X(net2431));
 sg13g2_dlygate4sd3_1 hold1304 (.A(_01496_),
    .X(net2432));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\TRNG.Word_Out[82] ),
    .X(net2433));
 sg13g2_dlygate4sd3_1 hold1306 (.A(_01327_),
    .X(net2434));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\TRNG.Word_Out[311] ),
    .X(net2435));
 sg13g2_dlygate4sd3_1 hold1308 (.A(\TRNG.Word_Out[274] ),
    .X(net2436));
 sg13g2_dlygate4sd3_1 hold1309 (.A(_01519_),
    .X(net2437));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\TRNG.Word_Out[184] ),
    .X(net2438));
 sg13g2_dlygate4sd3_1 hold1311 (.A(\TRNG.sha256.expand.data1_to_ram[5] ),
    .X(net2439));
 sg13g2_dlygate4sd3_1 hold1312 (.A(_02309_),
    .X(net2440));
 sg13g2_dlygate4sd3_1 hold1313 (.A(\TRNG.Padded_Out[492] ),
    .X(net2441));
 sg13g2_dlygate4sd3_1 hold1314 (.A(\TRNG.Padded_Out[491] ),
    .X(net2442));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\TRNG.sha256.expand.exp_ctrl.sum[10] ),
    .X(net2443));
 sg13g2_dlygate4sd3_1 hold1316 (.A(_00997_),
    .X(net2444));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\TRNG.Word_Out[221] ),
    .X(net2445));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\TRNG.Word_Out[213] ),
    .X(net2446));
 sg13g2_dlygate4sd3_1 hold1319 (.A(_01458_),
    .X(net2447));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\TRNG.Word_Out[188] ),
    .X(net2448));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\TRNG.Word_Out[391] ),
    .X(net2449));
 sg13g2_dlygate4sd3_1 hold1322 (.A(_01636_),
    .X(net2450));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\TRNG.Word_Out[356] ),
    .X(net2451));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\TRNG.Word_Out[366] ),
    .X(net2452));
 sg13g2_dlygate4sd3_1 hold1325 (.A(_01611_),
    .X(net2453));
 sg13g2_dlygate4sd3_1 hold1326 (.A(\TRNG.Word_Out[156] ),
    .X(net2454));
 sg13g2_dlygate4sd3_1 hold1327 (.A(\TRNG.Word_Out[378] ),
    .X(net2455));
 sg13g2_dlygate4sd3_1 hold1328 (.A(_01623_),
    .X(net2456));
 sg13g2_dlygate4sd3_1 hold1329 (.A(\TRNG.Word_Out[61] ),
    .X(net2457));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\TRNG.sha256.expand.exp_ctrl.sum[26] ),
    .X(net2458));
 sg13g2_dlygate4sd3_1 hold1331 (.A(_01013_),
    .X(net2459));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\TRNG.Padded_Out[359] ),
    .X(net2460));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\TRNG.Word_Out[347] ),
    .X(net2461));
 sg13g2_dlygate4sd3_1 hold1334 (.A(\TRNG.Word_Out[47] ),
    .X(net2462));
 sg13g2_dlygate4sd3_1 hold1335 (.A(_01292_),
    .X(net2463));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\TRNG.Padded_Out[503] ),
    .X(net2464));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\TRNG.Word_Out[179] ),
    .X(net2465));
 sg13g2_dlygate4sd3_1 hold1338 (.A(_01424_),
    .X(net2466));
 sg13g2_dlygate4sd3_1 hold1339 (.A(\TRNG.sha256.expand.exp_ctrl.sum[14] ),
    .X(net2467));
 sg13g2_dlygate4sd3_1 hold1340 (.A(_01001_),
    .X(net2468));
 sg13g2_dlygate4sd3_1 hold1341 (.A(\TRNG.Word_Out[18] ),
    .X(net2469));
 sg13g2_dlygate4sd3_1 hold1342 (.A(_01263_),
    .X(net2470));
 sg13g2_dlygate4sd3_1 hold1343 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][5] ),
    .X(net2471));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\TRNG.Padded_Out[494] ),
    .X(net2472));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\TRNG.Padded_Out[105] ),
    .X(net2473));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\TRNG.Word_Out[77] ),
    .X(net2474));
 sg13g2_dlygate4sd3_1 hold1347 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][4] ),
    .X(net2475));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\TRNG.sha256.expand.exp_ctrl.sum[15] ),
    .X(net2476));
 sg13g2_dlygate4sd3_1 hold1349 (.A(_01002_),
    .X(net2477));
 sg13g2_dlygate4sd3_1 hold1350 (.A(\TRNG.sha256.expand.exp_ctrl.sum[31] ),
    .X(net2478));
 sg13g2_dlygate4sd3_1 hold1351 (.A(_01018_),
    .X(net2479));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\TRNG.Padded_Out[490] ),
    .X(net2480));
 sg13g2_dlygate4sd3_1 hold1353 (.A(_02118_),
    .X(net2481));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\TRNG.uart_tx_inst.tx_reg[1] ),
    .X(net2482));
 sg13g2_dlygate4sd3_1 hold1355 (.A(_05920_),
    .X(net2483));
 sg13g2_dlygate4sd3_1 hold1356 (.A(_00106_),
    .X(net2484));
 sg13g2_dlygate4sd3_1 hold1357 (.A(\TRNG.Word_Out[246] ),
    .X(net2485));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\TRNG.Word_Out[31] ),
    .X(net2486));
 sg13g2_dlygate4sd3_1 hold1359 (.A(_01276_),
    .X(net2487));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\TRNG.Word_Out[244] ),
    .X(net2488));
 sg13g2_dlygate4sd3_1 hold1361 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][14] ),
    .X(net2489));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\TRNG.Word_Out[408] ),
    .X(net2490));
 sg13g2_dlygate4sd3_1 hold1363 (.A(\TRNG.Word_Out[354] ),
    .X(net2491));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\TRNG.sha256.expand.data1_to_ram[29] ),
    .X(net2492));
 sg13g2_dlygate4sd3_1 hold1365 (.A(_02393_),
    .X(net2493));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\TRNG.sha256.expand.exp_ctrl.j[1] ),
    .X(net2494));
 sg13g2_dlygate4sd3_1 hold1367 (.A(_02404_),
    .X(net2495));
 sg13g2_dlygate4sd3_1 hold1368 (.A(_00972_),
    .X(net2496));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\TRNG.Word_Out[380] ),
    .X(net2497));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][17] ),
    .X(net2498));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\TRNG.uart_tx_inst.tx_reg[5] ),
    .X(net2499));
 sg13g2_dlygate4sd3_1 hold1372 (.A(_00111_),
    .X(net2500));
 sg13g2_dlygate4sd3_1 hold1373 (.A(\TRNG.Word_Out[446] ),
    .X(net2501));
 sg13g2_dlygate4sd3_1 hold1374 (.A(_02139_),
    .X(net2502));
 sg13g2_dlygate4sd3_1 hold1375 (.A(\TRNG.Word_Out[144] ),
    .X(net2503));
 sg13g2_dlygate4sd3_1 hold1376 (.A(_01389_),
    .X(net2504));
 sg13g2_dlygate4sd3_1 hold1377 (.A(\TRNG.Word_Out[119] ),
    .X(net2505));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\TRNG.Word_Out[54] ),
    .X(net2506));
 sg13g2_dlygate4sd3_1 hold1379 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][10] ),
    .X(net2507));
 sg13g2_dlygate4sd3_1 hold1380 (.A(\TRNG.Word_Out[299] ),
    .X(net2508));
 sg13g2_dlygate4sd3_1 hold1381 (.A(_01544_),
    .X(net2509));
 sg13g2_dlygate4sd3_1 hold1382 (.A(\TRNG.Word_Out[39] ),
    .X(net2510));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\TRNG.Padded_Out[496] ),
    .X(net2511));
 sg13g2_dlygate4sd3_1 hold1384 (.A(\TRNG.sha256.expand.exp_ctrl.sum[30] ),
    .X(net2512));
 sg13g2_dlygate4sd3_1 hold1385 (.A(_01017_),
    .X(net2513));
 sg13g2_dlygate4sd3_1 hold1386 (.A(\TRNG.Word_Out[440] ),
    .X(net2514));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][28] ),
    .X(net2515));
 sg13g2_dlygate4sd3_1 hold1388 (.A(\TRNG.Word_Out[182] ),
    .X(net2516));
 sg13g2_dlygate4sd3_1 hold1389 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][9] ),
    .X(net2517));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][30] ),
    .X(net2518));
 sg13g2_dlygate4sd3_1 hold1391 (.A(\TRNG.Word_Out[293] ),
    .X(net2519));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\TRNG.raw_byte[4] ),
    .X(net2520));
 sg13g2_dlygate4sd3_1 hold1393 (.A(_05935_),
    .X(net2521));
 sg13g2_dlygate4sd3_1 hold1394 (.A(_00110_),
    .X(net2522));
 sg13g2_dlygate4sd3_1 hold1395 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][2] ),
    .X(net2523));
 sg13g2_dlygate4sd3_1 hold1396 (.A(_00787_),
    .X(net2524));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\TRNG.Word_Out[325] ),
    .X(net2525));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\TRNG.Padded_Out[498] ),
    .X(net2526));
 sg13g2_dlygate4sd3_1 hold1399 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][14] ),
    .X(net2527));
 sg13g2_dlygate4sd3_1 hold1400 (.A(\TRNG.raw_byte[7] ),
    .X(net2528));
 sg13g2_dlygate4sd3_1 hold1401 (.A(_02167_),
    .X(net2529));
 sg13g2_dlygate4sd3_1 hold1402 (.A(\TRNG.Word_Out[108] ),
    .X(net2530));
 sg13g2_dlygate4sd3_1 hold1403 (.A(_01353_),
    .X(net2531));
 sg13g2_dlygate4sd3_1 hold1404 (.A(\TRNG.sha256.expand.exp_ctrl.j_7[2] ),
    .X(net2532));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\TRNG.Word_Out[304] ),
    .X(net2533));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\TRNG.Word_Out[406] ),
    .X(net2534));
 sg13g2_dlygate4sd3_1 hold1407 (.A(_01651_),
    .X(net2535));
 sg13g2_dlygate4sd3_1 hold1408 (.A(\TRNG.sha256.expand.exp_ctrl.sum[11] ),
    .X(net2536));
 sg13g2_dlygate4sd3_1 hold1409 (.A(_00998_),
    .X(net2537));
 sg13g2_dlygate4sd3_1 hold1410 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][22] ),
    .X(net2538));
 sg13g2_dlygate4sd3_1 hold1411 (.A(\TRNG.Padded_Out[480] ),
    .X(net2539));
 sg13g2_dlygate4sd3_1 hold1412 (.A(\TRNG.Word_Out[214] ),
    .X(net2540));
 sg13g2_dlygate4sd3_1 hold1413 (.A(\TRNG.sha256.expand.exp_ctrl.sum[0] ),
    .X(net2541));
 sg13g2_dlygate4sd3_1 hold1414 (.A(_00987_),
    .X(net2542));
 sg13g2_dlygate4sd3_1 hold1415 (.A(\TRNG.Padded_Out[292] ),
    .X(net2543));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\TRNG.Word_Out[145] ),
    .X(net2544));
 sg13g2_dlygate4sd3_1 hold1417 (.A(_01390_),
    .X(net2545));
 sg13g2_dlygate4sd3_1 hold1418 (.A(\TRNG.Word_Out[261] ),
    .X(net2546));
 sg13g2_dlygate4sd3_1 hold1419 (.A(\TRNG.Padded_Out[339] ),
    .X(net2547));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\TRNG.Word_Out[21] ),
    .X(net2548));
 sg13g2_dlygate4sd3_1 hold1421 (.A(\TRNG.Word_Out[37] ),
    .X(net2549));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][0] ),
    .X(net2550));
 sg13g2_dlygate4sd3_1 hold1423 (.A(_00593_),
    .X(net2551));
 sg13g2_dlygate4sd3_1 hold1424 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][22] ),
    .X(net2552));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][13] ),
    .X(net2553));
 sg13g2_dlygate4sd3_1 hold1426 (.A(\TRNG.Word_Out[319] ),
    .X(net2554));
 sg13g2_dlygate4sd3_1 hold1427 (.A(_01564_),
    .X(net2555));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\TRNG.Word_Out[331] ),
    .X(net2556));
 sg13g2_dlygate4sd3_1 hold1429 (.A(\TRNG.bit_counter[7] ),
    .X(net2557));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\TRNG.Word_Out[85] ),
    .X(net2558));
 sg13g2_dlygate4sd3_1 hold1431 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][11] ),
    .X(net2559));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\TRNG.chunk_reg[6] ),
    .X(net2560));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\TRNG.Word_Out[367] ),
    .X(net2561));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][26] ),
    .X(net2562));
 sg13g2_dlygate4sd3_1 hold1435 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][29] ),
    .X(net2563));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\TRNG.Word_Out[212] ),
    .X(net2564));
 sg13g2_dlygate4sd3_1 hold1437 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][2] ),
    .X(net2565));
 sg13g2_dlygate4sd3_1 hold1438 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][19] ),
    .X(net2566));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][6] ),
    .X(net2567));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\TRNG.Padded_Out[160] ),
    .X(net2568));
 sg13g2_dlygate4sd3_1 hold1441 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][27] ),
    .X(net2569));
 sg13g2_dlygate4sd3_1 hold1442 (.A(_01046_),
    .X(net2570));
 sg13g2_dlygate4sd3_1 hold1443 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][2] ),
    .X(net2571));
 sg13g2_dlygate4sd3_1 hold1444 (.A(\TRNG.Word_Out[442] ),
    .X(net2572));
 sg13g2_dlygate4sd3_1 hold1445 (.A(\TRNG.Word_Out[32] ),
    .X(net2573));
 sg13g2_dlygate4sd3_1 hold1446 (.A(_01277_),
    .X(net2574));
 sg13g2_dlygate4sd3_1 hold1447 (.A(\TRNG.Padded_Out[504] ),
    .X(net2575));
 sg13g2_dlygate4sd3_1 hold1448 (.A(_02132_),
    .X(net2576));
 sg13g2_dlygate4sd3_1 hold1449 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][29] ),
    .X(net2577));
 sg13g2_dlygate4sd3_1 hold1450 (.A(\TRNG.Word_Out[58] ),
    .X(net2578));
 sg13g2_dlygate4sd3_1 hold1451 (.A(_01303_),
    .X(net2579));
 sg13g2_dlygate4sd3_1 hold1452 (.A(\TRNG.Padded_Out[506] ),
    .X(net2580));
 sg13g2_dlygate4sd3_1 hold1453 (.A(\TRNG.Padded_Out[102] ),
    .X(net2581));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\TRNG.Padded_Out[489] ),
    .X(net2582));
 sg13g2_dlygate4sd3_1 hold1455 (.A(\TRNG.Word_Out[248] ),
    .X(net2583));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\TRNG.Word_Out[371] ),
    .X(net2584));
 sg13g2_dlygate4sd3_1 hold1457 (.A(_01616_),
    .X(net2585));
 sg13g2_dlygate4sd3_1 hold1458 (.A(\TRNG.Word_Out[43] ),
    .X(net2586));
 sg13g2_dlygate4sd3_1 hold1459 (.A(\TRNG.Word_Out[394] ),
    .X(net2587));
 sg13g2_dlygate4sd3_1 hold1460 (.A(\TRNG.Word_Out[361] ),
    .X(net2588));
 sg13g2_dlygate4sd3_1 hold1461 (.A(_01606_),
    .X(net2589));
 sg13g2_dlygate4sd3_1 hold1462 (.A(\TRNG.Word_Out[178] ),
    .X(net2590));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\TRNG.hash[188] ),
    .X(net2591));
 sg13g2_dlygate4sd3_1 hold1464 (.A(_06981_),
    .X(net2592));
 sg13g2_dlygate4sd3_1 hold1465 (.A(_00487_),
    .X(net2593));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\TRNG.Word_Out[379] ),
    .X(net2594));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][0] ),
    .X(net2595));
 sg13g2_dlygate4sd3_1 hold1468 (.A(_01019_),
    .X(net2596));
 sg13g2_dlygate4sd3_1 hold1469 (.A(\TRNG.Word_Out[341] ),
    .X(net2597));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\TRNG.Padded_Out[222] ),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold1471 (.A(\TRNG.Word_Out[360] ),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][19] ),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold1473 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][22] ),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold1474 (.A(_00887_),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\TRNG.Word_Out[153] ),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold1476 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][18] ),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold1477 (.A(\TRNG.Word_Out[252] ),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold1478 (.A(\TRNG.Word_Out[5] ),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold1479 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][1] ),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold1480 (.A(_01020_),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold1481 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][28] ),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\TRNG.Word_Out[364] ),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold1483 (.A(\TRNG.Word_Out[2] ),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold1484 (.A(_01247_),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][31] ),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold1486 (.A(\TRNG.Word_Out[407] ),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\TRNG.Word_Out[10] ),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold1488 (.A(_01255_),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][3] ),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold1490 (.A(_01204_),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold1491 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][7] ),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold1492 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][20] ),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][14] ),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold1494 (.A(\TRNG.Word_Out[23] ),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\TRNG.sha256.expand.exp_ctrl.sum[25] ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold1496 (.A(_01012_),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold1497 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][15] ),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][3] ),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold1499 (.A(\TRNG.Word_Out[316] ),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][27] ),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold1501 (.A(\TRNG.Word_Out[338] ),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold1502 (.A(_01583_),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\TRNG.sha256.expand.data1_to_ram[20] ),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold1504 (.A(_02362_),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\TRNG.Padded_Out[295] ),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold1506 (.A(\TRNG.sha256.expand.exp_ctrl.sum[17] ),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold1507 (.A(_01004_),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\TRNG.sha256.W[14] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold1509 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][30] ),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\TRNG.Word_Out[337] ),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold1511 (.A(\TRNG.Word_Out[275] ),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold1512 (.A(_01520_),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\TRNG.Word_Out[412] ),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold1514 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][2] ),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold1515 (.A(_00867_),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][20] ),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold1517 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][7] ),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][16] ),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold1519 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][19] ),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\TRNG.Word_Out[204] ),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][5] ),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold1522 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][25] ),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold1523 (.A(\TRNG.Word_Out[160] ),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold1524 (.A(\TRNG.bit_counter[8] ),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold1525 (.A(_02156_),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold1526 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][27] ),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold1527 (.A(\TRNG.sha256.expand.exp_ctrl.j_15[1] ),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold1528 (.A(_02423_),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold1529 (.A(_00984_),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\TRNG.chunk_reg[4] ),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold1531 (.A(\TRNG.Word_Out[236] ),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold1532 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][22] ),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold1533 (.A(\TRNG.sha256.expand.exp_ctrl.sum[21] ),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold1534 (.A(_01008_),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][4] ),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][4] ),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold1537 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][23] ),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold1538 (.A(\TRNG.Padded_Out[495] ),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][24] ),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold1540 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][5] ),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\TRNG.Word_Out[282] ),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold1542 (.A(_00114_),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold1543 (.A(_00105_),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold1544 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][15] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold1545 (.A(_00880_),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold1546 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][3] ),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold1547 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][11] ),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold1548 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][3] ),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold1549 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][5] ),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold1550 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][29] ),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\TRNG.uart_tx_inst.currentState[4] ),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold1552 (.A(_05903_),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold1553 (.A(_00312_),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold1554 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][3] ),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\TRNG.Word_Out[308] ),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\TRNG.Word_Out[372] ),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold1557 (.A(\TRNG.Padded_Out[499] ),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold1558 (.A(\TRNG.Word_Out[155] ),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][4] ),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold1560 (.A(_00417_),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold1561 (.A(\TRNG.Word_Out[383] ),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold1562 (.A(\TRNG.Word_Out[11] ),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold1563 (.A(_01256_),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold1564 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][3] ),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold1565 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][28] ),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold1566 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][11] ),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold1567 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][23] ),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][20] ),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold1569 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][0] ),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold1570 (.A(_00753_),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold1571 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][23] ),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold1572 (.A(\TRNG.Padded_Out[502] ),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\TRNG.Word_Out[91] ),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold1574 (.A(_01336_),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][24] ),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold1576 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][12] ),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][4] ),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold1578 (.A(_00449_),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold1579 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][16] ),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold1580 (.A(\TRNG.Word_Out[117] ),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold1581 (.A(\TRNG.Word_Out[33] ),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold1582 (.A(_01278_),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold1583 (.A(\TRNG.Word_Out[175] ),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold1584 (.A(_01420_),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold1585 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][31] ),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][31] ),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold1587 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][5] ),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold1588 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][25] ),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold1589 (.A(_01226_),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold1590 (.A(\TRNG.Padded_Out[297] ),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold1591 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][10] ),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold1592 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][28] ),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold1593 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][23] ),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold1594 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][20] ),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][1] ),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold1596 (.A(_00414_),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\TRNG.raw_byte[5] ),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold1598 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][12] ),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold1599 (.A(_00877_),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][28] ),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold1601 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][23] ),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\TRNG.Word_Out[301] ),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold1603 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][9] ),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold1604 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][23] ),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold1605 (.A(\TRNG.Padded_Out[497] ),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold1606 (.A(_02125_),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold1607 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][15] ),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold1608 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][1] ),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold1609 (.A(_00754_),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][17] ),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold1611 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][20] ),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold1612 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][9] ),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold1613 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][6] ),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold1614 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][7] ),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][29] ),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold1616 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][20] ),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][10] ),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold1618 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][27] ),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold1619 (.A(_00812_),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold1620 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][5] ),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold1621 (.A(\TRNG.Word_Out[425] ),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold1622 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][24] ),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold1623 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][6] ),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold1624 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][13] ),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold1625 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][3] ),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\TRNG.bit_counter[6] ),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\TRNG.Word_Out[419] ),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][18] ),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold1629 (.A(\TRNG.Word_Out[20] ),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold1630 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][10] ),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold1631 (.A(_00699_),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold1632 (.A(\TRNG.chunk_reg[5] ),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold1633 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][15] ),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold1634 (.A(_00834_),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold1635 (.A(\TRNG.chunk_reg[2] ),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold1636 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][13] ),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold1637 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][1] ),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold1638 (.A(_00820_),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold1639 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][22] ),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold1640 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][20] ),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold1641 (.A(\TRNG.Word_Out[223] ),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold1642 (.A(\TRNG.Word_Out[340] ),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold1643 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][18] ),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold1644 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][12] ),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold1645 (.A(\TRNG.Word_Out[68] ),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold1646 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][1] ),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold1647 (.A(_01202_),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold1648 (.A(\TRNG.Word_Out[343] ),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold1649 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][11] ),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold1650 (.A(\TRNG.sha256.W[29] ),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold1651 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][13] ),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][10] ),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold1653 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][25] ),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][28] ),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold1655 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][24] ),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold1656 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][14] ),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold1657 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][9] ),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\TRNG.Word_Out[130] ),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold1659 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][27] ),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold1660 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][21] ),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold1661 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][8] ),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold1662 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][2] ),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold1663 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][0] ),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold1664 (.A(_00445_),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold1665 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][2] ),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold1666 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][26] ),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold1667 (.A(\TRNG.raw_byte[3] ),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold1668 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][9] ),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold1669 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][30] ),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold1670 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][6] ),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold1671 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][17] ),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold1672 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][10] ),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold1673 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][26] ),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold1674 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][18] ),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold1675 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][6] ),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold1676 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][0] ),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold1677 (.A(_00413_),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold1678 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][27] ),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold1679 (.A(_00892_),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold1680 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][7] ),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold1681 (.A(\TRNG.Padded_Out[484] ),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold1682 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][26] ),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold1683 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][15] ),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold1684 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][25] ),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold1685 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][30] ),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold1686 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][22] ),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold1687 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][17] ),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold1688 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][15] ),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold1689 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][0] ),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold1690 (.A(_00865_),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold1691 (.A(\TRNG.Word_Out[27] ),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold1692 (.A(_01272_),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold1693 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][14] ),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold1694 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][10] ),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold1695 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][9] ),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold1696 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][13] ),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold1697 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][17] ),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold1698 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][21] ),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold1699 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][26] ),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold1700 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][9] ),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold1701 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][11] ),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold1702 (.A(\TRNG.chunk_reg[7] ),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\TRNG.Word_Out[165] ),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold1704 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][20] ),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold1705 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][27] ),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold1706 (.A(_00440_),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold1707 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][16] ),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold1708 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][26] ),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold1709 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][0] ),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold1710 (.A(_01201_),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold1711 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][30] ),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][8] ),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][1] ),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold1714 (.A(_00866_),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold1715 (.A(\TRNG.Word_Out[370] ),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold1716 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][2] ),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold1717 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][11] ),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][26] ),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold1719 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][4] ),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold1720 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][25] ),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold1721 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][18] ),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold1722 (.A(\TRNG.Word_Out[42] ),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold1723 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][15] ),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold1724 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][13] ),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold1725 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][8] ),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold1726 (.A(_00697_),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold1727 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][1] ),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold1728 (.A(_00626_),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold1729 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][18] ),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold1730 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][3] ),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold1731 (.A(_01022_),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold1732 (.A(\TRNG.Padded_Out[485] ),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold1733 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][22] ),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold1734 (.A(\TRNG.chunk_reg[1] ),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold1735 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][4] ),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold1736 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][23] ),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold1737 (.A(\TRNG.Word_Out[277] ),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold1738 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][9] ),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold1739 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][14] ),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold1740 (.A(\TRNG.Word_Out[126] ),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold1741 (.A(\TRNG.raw_byte[2] ),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold1742 (.A(_02162_),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold1743 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][31] ),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold1744 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][22] ),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold1745 (.A(\TRNG.hash_rdy ),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold1746 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][3] ),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\TRNG.Word_Out[194] ),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold1748 (.A(_01438_),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][24] ),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold1750 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][26] ),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\TRNG.Word_Out[399] ),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold1752 (.A(\TRNG.NOISE_SAMPLER.Sample_Out ),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold1753 (.A(\TRNG.Word_Out[404] ),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold1754 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][4] ),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold1755 (.A(_00629_),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold1756 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][23] ),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold1757 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][0] ),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold1758 (.A(_00819_),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold1759 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][6] ),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold1760 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][16] ),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold1761 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][21] ),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold1762 (.A(\TRNG.Word_Out[64] ),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold1763 (.A(_01309_),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold1764 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][19] ),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold1765 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][21] ),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold1766 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][29] ),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold1767 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][28] ),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold1768 (.A(\TRNG.Word_Out[382] ),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold1769 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][10] ),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold1770 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][17] ),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold1771 (.A(_00398_),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold1772 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][21] ),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold1773 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][10] ),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold1774 (.A(\TRNG.Word_Out[167] ),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold1775 (.A(_01412_),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold1776 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][22] ),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold1777 (.A(\TRNG.Word_Out[416] ),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold1778 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][23] ),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold1779 (.A(\TRNG.Word_Out[402] ),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold1780 (.A(_01647_),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold1781 (.A(\TRNG.Word_Out[8] ),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold1782 (.A(\TRNG.Word_Out[132] ),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold1783 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][20] ),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold1784 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][12] ),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold1785 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][31] ),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold1786 (.A(\TRNG.Word_Out[134] ),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold1787 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][22] ),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold1788 (.A(\TRNG.Word_Out[307] ),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold1789 (.A(\TRNG.Word_Out[109] ),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold1790 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][30] ),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold1791 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][10] ),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold1792 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][17] ),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold1793 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][29] ),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold1794 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][14] ),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold1795 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][16] ),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold1796 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][31] ),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold1797 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][7] ),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold1798 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][31] ),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold1799 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][4] ),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold1800 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][24] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold1801 (.A(\TRNG.sha256.expand.msg_schdl.RAM[9][8] ),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold1802 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][3] ),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold1803 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][12] ),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold1804 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][20] ),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold1805 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][9] ),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold1806 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][25] ),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold1807 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][29] ),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold1808 (.A(\TRNG.discard ),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold1809 (.A(_04851_),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold1810 (.A(\TRNG.Word_Out[57] ),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold1811 (.A(\TRNG.Word_Out[48] ),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold1812 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][11] ),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold1813 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][11] ),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold1814 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][18] ),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold1815 (.A(\TRNG.Word_Out[411] ),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold1816 (.A(_01655_),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold1817 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][8] ),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold1818 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][1] ),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold1819 (.A(_00446_),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold1820 (.A(\TRNG.chunk_reg[3] ),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold1821 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][26] ),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold1822 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][7] ),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold1823 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][12] ),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold1824 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][15] ),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold1825 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][29] ),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold1826 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][5] ),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold1827 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][29] ),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold1828 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][18] ),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold1829 (.A(\TRNG.Word_Out[148] ),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold1830 (.A(\TRNG.Word_Out[73] ),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold1831 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][20] ),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold1832 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][21] ),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold1833 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][16] ),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold1834 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][16] ),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold1835 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][19] ),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold1836 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][14] ),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold1837 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][10] ),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold1838 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][17] ),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold1839 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][28] ),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold1840 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][8] ),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold1841 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][13] ),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold1842 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][4] ),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold1843 (.A(_00757_),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold1844 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][25] ),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold1845 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][6] ),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold1846 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][3] ),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold1847 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][26] ),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold1848 (.A(\TRNG.Word_Out[396] ),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold1849 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][28] ),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold1850 (.A(\TRNG.Word_Out[92] ),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold1851 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][7] ),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold1852 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][31] ),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold1853 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][16] ),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold1854 (.A(\TRNG.Word_Out[106] ),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold1855 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][18] ),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold1856 (.A(\TRNG.Word_Out[201] ),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold1857 (.A(_01446_),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold1858 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][1] ),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold1859 (.A(_00690_),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold1860 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][0] ),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold1861 (.A(_00689_),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold1862 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][6] ),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold1863 (.A(\TRNG.Word_Out[306] ),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold1864 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][7] ),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold1865 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][21] ),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold1866 (.A(_00806_),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold1867 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][19] ),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold1868 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][17] ),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold1869 (.A(\TRNG.Padded_Out[501] ),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold1870 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][5] ),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold1871 (.A(\TRNG.uart_start ),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold1872 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][31] ),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold1873 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][23] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold1874 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][3] ),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold1875 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][29] ),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold1876 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][19] ),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold1877 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][9] ),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold1878 (.A(_00390_),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold1879 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][11] ),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold1880 (.A(_00392_),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold1881 (.A(\TRNG.bit_counter[2] ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold1882 (.A(_04861_),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold1883 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][11] ),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold1884 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][24] ),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold1885 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][26] ),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold1886 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][15] ),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold1887 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][18] ),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold1888 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][17] ),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold1889 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][12] ),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold1890 (.A(_00831_),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold1891 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][7] ),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold1892 (.A(_00600_),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold1893 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][17] ),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold1894 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][30] ),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold1895 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][29] ),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold1896 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][20] ),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold1897 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][20] ),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold1898 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][25] ),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold1899 (.A(\TRNG.Word_Out[320] ),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold1900 (.A(\TRNG.Word_Out[136] ),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold1901 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][1] ),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold1902 (.A(_00786_),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold1903 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][7] ),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold1904 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][13] ),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold1905 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][29] ),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold1906 (.A(\TRNG.Word_Out[439] ),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold1907 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][12] ),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold1908 (.A(_00797_),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold1909 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][29] ),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold1910 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][0] ),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold1911 (.A(_00381_),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold1912 (.A(\TRNG.Word_Out[432] ),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold1913 (.A(\TRNG.raw_byte[0] ),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold1914 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][5] ),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold1915 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][24] ),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold1916 (.A(\TRNG.Word_Out[203] ),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold1917 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][28] ),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold1918 (.A(\TRNG.Word_Out[255] ),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold1919 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][14] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold1920 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][12] ),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold1921 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][30] ),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold1922 (.A(\TRNG.Word_Out[268] ),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold1923 (.A(_01513_),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold1924 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][17] ),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold1925 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][16] ),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold1926 (.A(\TRNG.Word_Out[99] ),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold1927 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][9] ),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold1928 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][18] ),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold1929 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][26] ),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold1930 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][27] ),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold1931 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][28] ),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold1932 (.A(_00813_),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold1933 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][27] ),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold1934 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][15] ),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold1935 (.A(\TRNG.sha256.expand.data1_to_ram[0] ),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold1936 (.A(_00721_),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold1937 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][17] ),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold1938 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][30] ),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold1939 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][28] ),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold1940 (.A(\TRNG.sha256.expand.data1_to_ram[1] ),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold1941 (.A(_02295_),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold1942 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][24] ),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold1943 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][5] ),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold1944 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][8] ),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold1945 (.A(\TRNG.bit_counter[3] ),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold1946 (.A(_04864_),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold1947 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][12] ),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold1948 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][15] ),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold1949 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][14] ),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold1950 (.A(\TRNG.Word_Out[290] ),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold1951 (.A(\TRNG.sha256.expand.data1_to_ram[2] ),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold1952 (.A(_02299_),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold1953 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][0] ),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold1954 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][6] ),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold1955 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][24] ),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold1956 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][10] ),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold1957 (.A(\TRNG.Word_Out[1] ),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold1958 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][14] ),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold1959 (.A(\TRNG.Word_Out[12] ),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold1960 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][13] ),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold1961 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][13] ),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold1962 (.A(\TRNG.Word_Out[168] ),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold1963 (.A(\TRNG.Word_Out[269] ),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold1964 (.A(\TRNG.Word_Out[180] ),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold1965 (.A(\TRNG.Word_Out[51] ),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold1966 (.A(\TRNG.sha256.W[13] ),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold1967 (.A(_00910_),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold1968 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][21] ),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold1969 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][8] ),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold1970 (.A(\TRNG.Word_Out[330] ),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold1971 (.A(_01574_),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold1972 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][15] ),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold1973 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][1] ),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold1974 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][31] ),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold1975 (.A(_00624_),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold1976 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][9] ),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold1977 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][2] ),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold1978 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][27] ),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold1979 (.A(\TRNG.Word_Out[176] ),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold1980 (.A(\TRNG.chunk_reg[0] ),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold1981 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][23] ),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold1982 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][18] ),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold1983 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][4] ),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold1984 (.A(_00353_),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold1985 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][21] ),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold1986 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][2] ),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold1987 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][12] ),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold1988 (.A(\TRNG.Word_Out[19] ),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold1989 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][12] ),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold1990 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][6] ),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold1991 (.A(\TRNG.Padded_Out[190] ),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold1992 (.A(\TRNG.Word_Out[41] ),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold1993 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][11] ),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold1994 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][8] ),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold1995 (.A(\TRNG.raw_byte[6] ),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold1996 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][1] ),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold1997 (.A(\TRNG.Word_Out[339] ),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold1998 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][25] ),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold1999 (.A(\TRNG.Word_Out[243] ),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold2000 (.A(\TRNG.Word_Out[162] ),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold2001 (.A(\TRNG.Word_Out[362] ),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold2002 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][30] ),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold2003 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][19] ),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold2004 (.A(\TRNG.raw_byte[1] ),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold2005 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][5] ),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold2006 (.A(_00209_),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold2007 (.A(_00541_),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold2008 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][6] ),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold2009 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][1] ),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold2010 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][9] ),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold2011 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][30] ),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold2012 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][19] ),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold2013 (.A(_00400_),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold2014 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][4] ),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold2015 (.A(_00385_),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold2016 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][30] ),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold2017 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][25] ),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold2018 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][22] ),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold2019 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][4] ),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold2020 (.A(_00693_),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold2021 (.A(\TRNG.Repetition_Count_Test.count[5] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold2022 (.A(_03087_),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold2023 (.A(_01233_),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold2024 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][25] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold2025 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][0] ),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold2026 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][25] ),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold2027 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][5] ),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold2028 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][25] ),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold2029 (.A(\TRNG.Word_Out[114] ),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold2030 (.A(\TRNG.Word_Out[83] ),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold2031 (.A(_00205_),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold2032 (.A(_07494_),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold2033 (.A(_00538_),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold2034 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][22] ),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold2035 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][31] ),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold2036 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][31] ),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold2037 (.A(\TRNG.Word_Out[65] ),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold2038 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][29] ),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold2039 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][11] ),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold2040 (.A(\TRNG.sha256.expand.msg_schdl.RAM[12][14] ),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold2041 (.A(\TRNG.uart_tx_inst.ticks_counter[5] ),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold2042 (.A(_00861_),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold2043 (.A(\TRNG.Word_Out[202] ),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold2044 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][5] ),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold2045 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][16] ),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold2046 (.A(_00769_),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold2047 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][6] ),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold2048 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][13] ),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold2049 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][24] ),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold2050 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][8] ),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold2051 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][28] ),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold2052 (.A(\TRNG.Word_Out[276] ),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold2053 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][26] ),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold2054 (.A(\TRNG.Word_Out[25] ),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold2055 (.A(_00211_),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold2056 (.A(_00543_),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold2057 (.A(\TRNG.Word_Out[351] ),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold2058 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][1] ),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold2059 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][31] ),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold2060 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][8] ),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold2061 (.A(\TRNG.Word_Out[28] ),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold2062 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][25] ),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold2063 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][22] ),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold2064 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][16] ),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold2065 (.A(\TRNG.Word_Out[76] ),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold2066 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][6] ),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold2067 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][13] ),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold2068 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][24] ),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold2069 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][8] ),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold2070 (.A(_00665_),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold2071 (.A(\TRNG.Word_Out[34] ),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold2072 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][18] ),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold2073 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][7] ),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold2074 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][29] ),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold2075 (.A(\TRNG.Word_Out[242] ),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold2076 (.A(\TRNG.sha256.expand.data1_to_ram[4] ),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold2077 (.A(_00321_),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold2078 (.A(\TRNG.Word_Out[335] ),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold2079 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][2] ),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold2080 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][27] ),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold2081 (.A(\TRNG.Word_Out[3] ),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold2082 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][22] ),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold2083 (.A(\TRNG.Word_Out[191] ),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold2084 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][3] ),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold2085 (.A(_00384_),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold2086 (.A(\TRNG.Word_Out[75] ),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold2087 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][15] ),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold2088 (.A(_00800_),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold2089 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][24] ),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold2090 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][5] ),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold2091 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][12] ),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold2092 (.A(\TRNG.Word_Out[239] ),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold2093 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][17] ),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold2094 (.A(_00123_),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold2095 (.A(_04218_),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold2096 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][17] ),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold2097 (.A(\TRNG.Word_Out[284] ),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold2098 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][23] ),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold2099 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][16] ),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold2100 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][18] ),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold2101 (.A(\TRNG.Word_Out[226] ),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold2102 (.A(_01470_),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold2103 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][10] ),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold2104 (.A(\TRNG.sha256.expand.data1_to_ram[3] ),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold2105 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][7] ),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold2106 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][2] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold2107 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][14] ),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold2108 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][2] ),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold2109 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][23] ),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold2110 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][19] ),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold2111 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][19] ),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold2112 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][21] ),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold2113 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][21] ),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold2114 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][22] ),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold2115 (.A(_00743_),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold2116 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][1] ),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold2117 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][8] ),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold2118 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][28] ),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold2119 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][23] ),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold2120 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][2] ),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold2121 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][19] ),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold2122 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][21] ),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold2123 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][7] ),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold2124 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][0] ),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold2125 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][10] ),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold2126 (.A(\TRNG.Word_Out[146] ),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold2127 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][27] ),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold2128 (.A(_01228_),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold2129 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][13] ),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold2130 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][23] ),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold2131 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][30] ),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold2132 (.A(_00687_),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold2133 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][26] ),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold2134 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][16] ),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold2135 (.A(\TRNG.Word_Out[403] ),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold2136 (.A(_00124_),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold2137 (.A(_04215_),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold2138 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][11] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold2139 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][9] ),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold2140 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][20] ),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold2141 (.A(\TRNG.uart_tx_inst.ticks_counter[8] ),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold2142 (.A(_08853_),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold2143 (.A(\TRNG.Word_Out[140] ),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold2144 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][10] ),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold2145 (.A(\TRNG.Word_Out[129] ),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold2146 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][11] ),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold2147 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][21] ),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold2148 (.A(_00742_),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold2149 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][27] ),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold2150 (.A(_00620_),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold2151 (.A(\TRNG.Word_Out[392] ),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold2152 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][27] ),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold2153 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][0] ),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold2154 (.A(\TRNG.Word_Out[296] ),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold2155 (.A(\TRNG.sha256.connect[5] ),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold2156 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][29] ),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold2157 (.A(\TRNG.sha256.expand.exp_ctrl.j_2[2] ),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold2158 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][31] ),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold2159 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][17] ),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold2160 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][2] ),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold2161 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][26] ),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold2162 (.A(\TRNG.Word_Out[250] ),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold2163 (.A(_00115_),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold2164 (.A(_04834_),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold2165 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][5] ),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold2166 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][19] ),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold2167 (.A(_00676_),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold2168 (.A(\TRNG.Word_Out[211] ),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold2169 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][19] ),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold2170 (.A(\TRNG.Word_Out[59] ),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold2171 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][3] ),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold2172 (.A(\TRNG.sha256.W[12] ),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold2173 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][20] ),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold2174 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][7] ),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold2175 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][8] ),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold2176 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][26] ),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold2177 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][15] ),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold2178 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][24] ),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold2179 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][23] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold2180 (.A(_00616_),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold2181 (.A(\TRNG.Padded_Out[511] ),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold2182 (.A(_02253_),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold2183 (.A(\TRNG.Word_Out[233] ),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold2184 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][24] ),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold2185 (.A(\TRNG.Word_Out[377] ),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold2186 (.A(\TRNG.raw_bit_counter[2] ),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold2187 (.A(_02147_),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold2188 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][2] ),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold2189 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][15] ),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold2190 (.A(_00736_),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold2191 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][16] ),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold2192 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][0] ),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold2193 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][18] ),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold2194 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][6] ),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold2195 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][13] ),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold2196 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][10] ),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold2197 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][2] ),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold2198 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][21] ),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold2199 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][13] ),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold2200 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][14] ),
    .X(net3328));
 sg13g2_dlygate4sd3_1 hold2201 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][28] ),
    .X(net3329));
 sg13g2_dlygate4sd3_1 hold2202 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][12] ),
    .X(net3330));
 sg13g2_dlygate4sd3_1 hold2203 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][5] ),
    .X(net3331));
 sg13g2_dlygate4sd3_1 hold2204 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][30] ),
    .X(net3332));
 sg13g2_dlygate4sd3_1 hold2205 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][12] ),
    .X(net3333));
 sg13g2_dlygate4sd3_1 hold2206 (.A(_00733_),
    .X(net3334));
 sg13g2_dlygate4sd3_1 hold2207 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][18] ),
    .X(net3335));
 sg13g2_dlygate4sd3_1 hold2208 (.A(\TRNG.sha256.control.iteration[8] ),
    .X(net3336));
 sg13g2_dlygate4sd3_1 hold2209 (.A(_08829_),
    .X(net3337));
 sg13g2_dlygate4sd3_1 hold2210 (.A(_00818_),
    .X(net3338));
 sg13g2_dlygate4sd3_1 hold2211 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][1] ),
    .X(net3339));
 sg13g2_dlygate4sd3_1 hold2212 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][31] ),
    .X(net3340));
 sg13g2_dlygate4sd3_1 hold2213 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][24] ),
    .X(net3341));
 sg13g2_dlygate4sd3_1 hold2214 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][27] ),
    .X(net3342));
 sg13g2_dlygate4sd3_1 hold2215 (.A(_00748_),
    .X(net3343));
 sg13g2_dlygate4sd3_1 hold2216 (.A(\TRNG.Word_Out[89] ),
    .X(net3344));
 sg13g2_dlygate4sd3_1 hold2217 (.A(\TRNG.sha256.expand.data1_to_ram[27] ),
    .X(net3345));
 sg13g2_dlygate4sd3_1 hold2218 (.A(_00684_),
    .X(net3346));
 sg13g2_dlygate4sd3_1 hold2219 (.A(\TRNG.sha256.W[18] ),
    .X(net3347));
 sg13g2_dlygate4sd3_1 hold2220 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][6] ),
    .X(net3348));
 sg13g2_dlygate4sd3_1 hold2221 (.A(_00663_),
    .X(net3349));
 sg13g2_dlygate4sd3_1 hold2222 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][9] ),
    .X(net3350));
 sg13g2_dlygate4sd3_1 hold2223 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][7] ),
    .X(net3351));
 sg13g2_dlygate4sd3_1 hold2224 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][4] ),
    .X(net3352));
 sg13g2_dlygate4sd3_1 hold2225 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][6] ),
    .X(net3353));
 sg13g2_dlygate4sd3_1 hold2226 (.A(\TRNG.uart_tx_inst.ticks_counter[2] ),
    .X(net3354));
 sg13g2_dlygate4sd3_1 hold2227 (.A(_00858_),
    .X(net3355));
 sg13g2_dlygate4sd3_1 hold2228 (.A(\TRNG.Padded_Out[500] ),
    .X(net3356));
 sg13g2_dlygate4sd3_1 hold2229 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][11] ),
    .X(net3357));
 sg13g2_dlygate4sd3_1 hold2230 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][30] ),
    .X(net3358));
 sg13g2_dlygate4sd3_1 hold2231 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][8] ),
    .X(net3359));
 sg13g2_dlygate4sd3_1 hold2232 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][14] ),
    .X(net3360));
 sg13g2_dlygate4sd3_1 hold2233 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][8] ),
    .X(net3361));
 sg13g2_dlygate4sd3_1 hold2234 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][28] ),
    .X(net3362));
 sg13g2_dlygate4sd3_1 hold2235 (.A(_00749_),
    .X(net3363));
 sg13g2_dlygate4sd3_1 hold2236 (.A(\TRNG.sha256.expand.msg_schdl.RAM[5][19] ),
    .X(net3364));
 sg13g2_dlygate4sd3_1 hold2237 (.A(\TRNG.Word_Out[300] ),
    .X(net3365));
 sg13g2_dlygate4sd3_1 hold2238 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][9] ),
    .X(net3366));
 sg13g2_dlygate4sd3_1 hold2239 (.A(\TRNG.sha256.expand.msg_schdl.RAM[8][30] ),
    .X(net3367));
 sg13g2_dlygate4sd3_1 hold2240 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][22] ),
    .X(net3368));
 sg13g2_dlygate4sd3_1 hold2241 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][4] ),
    .X(net3369));
 sg13g2_dlygate4sd3_1 hold2242 (.A(\TRNG.Repetition_Count_Test.count[4] ),
    .X(net3370));
 sg13g2_dlygate4sd3_1 hold2243 (.A(\TRNG.sha256.W[1] ),
    .X(net3371));
 sg13g2_dlygate4sd3_1 hold2244 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][16] ),
    .X(net3372));
 sg13g2_dlygate4sd3_1 hold2245 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][15] ),
    .X(net3373));
 sg13g2_dlygate4sd3_1 hold2246 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][20] ),
    .X(net3374));
 sg13g2_dlygate4sd3_1 hold2247 (.A(\TRNG.sha256.W[5] ),
    .X(net3375));
 sg13g2_dlygate4sd3_1 hold2248 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][14] ),
    .X(net3376));
 sg13g2_dlygate4sd3_1 hold2249 (.A(_00363_),
    .X(net3377));
 sg13g2_dlygate4sd3_1 hold2250 (.A(_00119_),
    .X(net3378));
 sg13g2_dlygate4sd3_1 hold2251 (.A(_04945_),
    .X(net3379));
 sg13g2_dlygate4sd3_1 hold2252 (.A(_02158_),
    .X(net3380));
 sg13g2_dlygate4sd3_1 hold2253 (.A(\TRNG.Word_Out[346] ),
    .X(net3381));
 sg13g2_dlygate4sd3_1 hold2254 (.A(_00186_),
    .X(net3382));
 sg13g2_dlygate4sd3_1 hold2255 (.A(_00529_),
    .X(net3383));
 sg13g2_dlygate4sd3_1 hold2256 (.A(_00129_),
    .X(net3384));
 sg13g2_dlygate4sd3_1 hold2257 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][25] ),
    .X(net3385));
 sg13g2_dlygate4sd3_1 hold2258 (.A(\TRNG.sha256.expand.exp_ctrl.j_2[1] ),
    .X(net3386));
 sg13g2_dlygate4sd3_1 hold2259 (.A(\TRNG.sha256.expand.msg_schdl.RAM[3][19] ),
    .X(net3387));
 sg13g2_dlygate4sd3_1 hold2260 (.A(_00197_),
    .X(net3388));
 sg13g2_dlygate4sd3_1 hold2261 (.A(_01166_),
    .X(net3389));
 sg13g2_dlygate4sd3_1 hold2262 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][31] ),
    .X(net3390));
 sg13g2_dlygate4sd3_1 hold2263 (.A(\TRNG.uart_tx_inst.currentState[3] ),
    .X(net3391));
 sg13g2_dlygate4sd3_1 hold2264 (.A(_04884_),
    .X(net3392));
 sg13g2_dlygate4sd3_1 hold2265 (.A(_00308_),
    .X(net3393));
 sg13g2_dlygate4sd3_1 hold2266 (.A(\TRNG.Repetition_Count_Test.prev_bit ),
    .X(net3394));
 sg13g2_dlygate4sd3_1 hold2267 (.A(\TRNG.hash[247] ),
    .X(net3395));
 sg13g2_dlygate4sd3_1 hold2268 (.A(_08236_),
    .X(net3396));
 sg13g2_dlygate4sd3_1 hold2269 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][25] ),
    .X(net3397));
 sg13g2_dlygate4sd3_1 hold2270 (.A(\TRNG.sha256.expand.exp_ctrl.j[3] ),
    .X(net3398));
 sg13g2_dlygate4sd3_1 hold2271 (.A(_02409_),
    .X(net3399));
 sg13g2_dlygate4sd3_1 hold2272 (.A(\TRNG.raw_bit_counter[1] ),
    .X(net3400));
 sg13g2_dlygate4sd3_1 hold2273 (.A(_04900_),
    .X(net3401));
 sg13g2_dlygate4sd3_1 hold2274 (.A(_02146_),
    .X(net3402));
 sg13g2_dlygate4sd3_1 hold2275 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][16] ),
    .X(net3403));
 sg13g2_dlygate4sd3_1 hold2276 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][13] ),
    .X(net3404));
 sg13g2_dlygate4sd3_1 hold2277 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][11] ),
    .X(net3405));
 sg13g2_dlygate4sd3_1 hold2278 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][7] ),
    .X(net3406));
 sg13g2_dlygate4sd3_1 hold2279 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][12] ),
    .X(net3407));
 sg13g2_dlygate4sd3_1 hold2280 (.A(_00187_),
    .X(net3408));
 sg13g2_dlygate4sd3_1 hold2281 (.A(_00531_),
    .X(net3409));
 sg13g2_dlygate4sd3_1 hold2282 (.A(\TRNG.hash[160] ),
    .X(net3410));
 sg13g2_dlygate4sd3_1 hold2283 (.A(_06882_),
    .X(net3411));
 sg13g2_dlygate4sd3_1 hold2284 (.A(_00165_),
    .X(net3412));
 sg13g2_dlygate4sd3_1 hold2285 (.A(_00509_),
    .X(net3413));
 sg13g2_dlygate4sd3_1 hold2286 (.A(\TRNG.sha256.expand.msg_schdl.RAM[4][21] ),
    .X(net3414));
 sg13g2_dlygate4sd3_1 hold2287 (.A(_00184_),
    .X(net3415));
 sg13g2_dlygate4sd3_1 hold2288 (.A(_07164_),
    .X(net3416));
 sg13g2_dlygate4sd3_1 hold2289 (.A(_00526_),
    .X(net3417));
 sg13g2_dlygate4sd3_1 hold2290 (.A(\TRNG.uart_tx_inst.ticks_counter[7] ),
    .X(net3418));
 sg13g2_dlygate4sd3_1 hold2291 (.A(_00181_),
    .X(net3419));
 sg13g2_dlygate4sd3_1 hold2292 (.A(_00525_),
    .X(net3420));
 sg13g2_dlygate4sd3_1 hold2293 (.A(\TRNG.sha256.expand.data1_to_ram[15] ),
    .X(net3421));
 sg13g2_dlygate4sd3_1 hold2294 (.A(_02346_),
    .X(net3422));
 sg13g2_dlygate4sd3_1 hold2295 (.A(_00222_),
    .X(net3423));
 sg13g2_dlygate4sd3_1 hold2296 (.A(_02726_),
    .X(net3424));
 sg13g2_dlygate4sd3_1 hold2297 (.A(\TRNG.Word_Out[281] ),
    .X(net3425));
 sg13g2_dlygate4sd3_1 hold2298 (.A(\TRNG.sha256.W[25] ),
    .X(net3426));
 sg13g2_dlygate4sd3_1 hold2299 (.A(\TRNG.hash[254] ),
    .X(net3427));
 sg13g2_dlygate4sd3_1 hold2300 (.A(_08250_),
    .X(net3428));
 sg13g2_dlygate4sd3_1 hold2301 (.A(\TRNG.sha256.expand.msg_schdl.RAM[0][21] ),
    .X(net3429));
 sg13g2_dlygate4sd3_1 hold2302 (.A(\TRNG.sha256.expand.exp_ctrl.j_15[2] ),
    .X(net3430));
 sg13g2_dlygate4sd3_1 hold2303 (.A(_02426_),
    .X(net3431));
 sg13g2_dlygate4sd3_1 hold2304 (.A(\TRNG.hash[244] ),
    .X(net3432));
 sg13g2_dlygate4sd3_1 hold2305 (.A(_08231_),
    .X(net3433));
 sg13g2_dlygate4sd3_1 hold2306 (.A(\TRNG.hash[107] ),
    .X(net3434));
 sg13g2_dlygate4sd3_1 hold2307 (.A(_02904_),
    .X(net3435));
 sg13g2_dlygate4sd3_1 hold2308 (.A(_01157_),
    .X(net3436));
 sg13g2_dlygate4sd3_1 hold2309 (.A(_00225_),
    .X(net3437));
 sg13g2_dlygate4sd3_1 hold2310 (.A(_01106_),
    .X(net3438));
 sg13g2_dlygate4sd3_1 hold2311 (.A(_00228_),
    .X(net3439));
 sg13g2_dlygate4sd3_1 hold2312 (.A(\TRNG.hash[252] ),
    .X(net3440));
 sg13g2_dlygate4sd3_1 hold2313 (.A(_00591_),
    .X(net3441));
 sg13g2_dlygate4sd3_1 hold2314 (.A(\TRNG.sha256.W[15] ),
    .X(net3442));
 sg13g2_dlygate4sd3_1 hold2315 (.A(_00125_),
    .X(net3443));
 sg13g2_dlygate4sd3_1 hold2316 (.A(_04214_),
    .X(net3444));
 sg13g2_dlygate4sd3_1 hold2317 (.A(_00191_),
    .X(net3445));
 sg13g2_dlygate4sd3_1 hold2318 (.A(_02891_),
    .X(net3446));
 sg13g2_dlygate4sd3_1 hold2319 (.A(\TRNG.hash[77] ),
    .X(net3447));
 sg13g2_dlygate4sd3_1 hold2320 (.A(_01158_),
    .X(net3448));
 sg13g2_dlygate4sd3_1 hold2321 (.A(\TRNG.Repetition_Count_Test.failure ),
    .X(net3449));
 sg13g2_dlygate4sd3_1 hold2322 (.A(\TRNG.sha256.expand.exp_ctrl.j_15[3] ),
    .X(net3450));
 sg13g2_dlygate4sd3_1 hold2323 (.A(\TRNG.sha256.control.iteration[6] ),
    .X(net3451));
 sg13g2_dlygate4sd3_1 hold2324 (.A(_00817_),
    .X(net3452));
 sg13g2_dlygate4sd3_1 hold2325 (.A(\TRNG.sha256.expand.data1_to_ram[19] ),
    .X(net3453));
 sg13g2_dlygate4sd3_1 hold2326 (.A(_02359_),
    .X(net3454));
 sg13g2_dlygate4sd3_1 hold2327 (.A(_00195_),
    .X(net3455));
 sg13g2_dlygate4sd3_1 hold2328 (.A(_01161_),
    .X(net3456));
 sg13g2_dlygate4sd3_1 hold2329 (.A(_00178_),
    .X(net3457));
 sg13g2_dlygate4sd3_1 hold2330 (.A(_00519_),
    .X(net3458));
 sg13g2_dlygate4sd3_1 hold2331 (.A(\TRNG.sha256.expand.exp_ctrl.j[2] ),
    .X(net3459));
 sg13g2_dlygate4sd3_1 hold2332 (.A(_02407_),
    .X(net3460));
 sg13g2_dlygate4sd3_1 hold2333 (.A(\TRNG.hash[39] ),
    .X(net3461));
 sg13g2_dlygate4sd3_1 hold2334 (.A(_00493_),
    .X(net3462));
 sg13g2_dlygate4sd3_1 hold2335 (.A(_00189_),
    .X(net3463));
 sg13g2_dlygate4sd3_1 hold2336 (.A(_00534_),
    .X(net3464));
 sg13g2_dlygate4sd3_1 hold2337 (.A(\TRNG.hash[141] ),
    .X(net3465));
 sg13g2_dlygate4sd3_1 hold2338 (.A(_01070_),
    .X(net3466));
 sg13g2_dlygate4sd3_1 hold2339 (.A(\TRNG.sha256.expand.data1_to_ram[28] ),
    .X(net3467));
 sg13g2_dlygate4sd3_1 hold2340 (.A(_02389_),
    .X(net3468));
 sg13g2_dlygate4sd3_1 hold2341 (.A(_00170_),
    .X(net3469));
 sg13g2_dlygate4sd3_1 hold2342 (.A(_07119_),
    .X(net3470));
 sg13g2_dlygate4sd3_1 hold2343 (.A(_00516_),
    .X(net3471));
 sg13g2_dlygate4sd3_1 hold2344 (.A(_00188_),
    .X(net3472));
 sg13g2_dlygate4sd3_1 hold2345 (.A(_00533_),
    .X(net3473));
 sg13g2_dlygate4sd3_1 hold2346 (.A(_00229_),
    .X(net3474));
 sg13g2_dlygate4sd3_1 hold2347 (.A(_01103_),
    .X(net3475));
 sg13g2_dlygate4sd3_1 hold2348 (.A(_00227_),
    .X(net3476));
 sg13g2_dlygate4sd3_1 hold2349 (.A(_01115_),
    .X(net3477));
 sg13g2_dlygate4sd3_1 hold2350 (.A(\TRNG.sha256.W[4] ),
    .X(net3478));
 sg13g2_dlygate4sd3_1 hold2351 (.A(\TRNG.chunk_index[1] ),
    .X(net3479));
 sg13g2_dlygate4sd3_1 hold2352 (.A(_00168_),
    .X(net3480));
 sg13g2_dlygate4sd3_1 hold2353 (.A(_00511_),
    .X(net3481));
 sg13g2_dlygate4sd3_1 hold2354 (.A(_00137_),
    .X(net3482));
 sg13g2_dlygate4sd3_1 hold2355 (.A(_00482_),
    .X(net3483));
 sg13g2_dlygate4sd3_1 hold2356 (.A(\TRNG.sha256.expand.dout2[0] ),
    .X(net3484));
 sg13g2_dlygate4sd3_1 hold2357 (.A(_00276_),
    .X(net3485));
 sg13g2_dlygate4sd3_1 hold2358 (.A(_00166_),
    .X(net3486));
 sg13g2_dlygate4sd3_1 hold2359 (.A(_07089_),
    .X(net3487));
 sg13g2_dlygate4sd3_1 hold2360 (.A(_00510_),
    .X(net3488));
 sg13g2_dlygate4sd3_1 hold2361 (.A(_00163_),
    .X(net3489));
 sg13g2_dlygate4sd3_1 hold2362 (.A(_07073_),
    .X(net3490));
 sg13g2_dlygate4sd3_1 hold2363 (.A(_00507_),
    .X(net3491));
 sg13g2_dlygate4sd3_1 hold2364 (.A(_00179_),
    .X(net3492));
 sg13g2_dlygate4sd3_1 hold2365 (.A(_07143_),
    .X(net3493));
 sg13g2_dlygate4sd3_1 hold2366 (.A(_00522_),
    .X(net3494));
 sg13g2_dlygate4sd3_1 hold2367 (.A(_00224_),
    .X(net3495));
 sg13g2_dlygate4sd3_1 hold2368 (.A(_01134_),
    .X(net3496));
 sg13g2_dlygate4sd3_1 hold2369 (.A(\TRNG.hash[169] ),
    .X(net3497));
 sg13g2_dlygate4sd3_1 hold2370 (.A(_00480_),
    .X(net3498));
 sg13g2_dlygate4sd3_1 hold2371 (.A(\TRNG.hash[245] ),
    .X(net3499));
 sg13g2_dlygate4sd3_1 hold2372 (.A(_00161_),
    .X(net3500));
 sg13g2_dlygate4sd3_1 hold2373 (.A(_07068_),
    .X(net3501));
 sg13g2_dlygate4sd3_1 hold2374 (.A(_00506_),
    .X(net3502));
 sg13g2_dlygate4sd3_1 hold2375 (.A(_00221_),
    .X(net3503));
 sg13g2_dlygate4sd3_1 hold2376 (.A(_01120_),
    .X(net3504));
 sg13g2_dlygate4sd3_1 hold2377 (.A(_00144_),
    .X(net3505));
 sg13g2_dlygate4sd3_1 hold2378 (.A(_06985_),
    .X(net3506));
 sg13g2_dlygate4sd3_1 hold2379 (.A(_00488_),
    .X(net3507));
 sg13g2_dlygate4sd3_1 hold2380 (.A(_00134_),
    .X(net3508));
 sg13g2_dlygate4sd3_1 hold2381 (.A(_06924_),
    .X(net3509));
 sg13g2_dlygate4sd3_1 hold2382 (.A(_00478_),
    .X(net3510));
 sg13g2_dlygate4sd3_1 hold2383 (.A(\TRNG.sha256.expand.data1_to_ram[17] ),
    .X(net3511));
 sg13g2_dlygate4sd3_1 hold2384 (.A(_02352_),
    .X(net3512));
 sg13g2_dlygate4sd3_1 hold2385 (.A(\TRNG.hash[199] ),
    .X(net3513));
 sg13g2_dlygate4sd3_1 hold2386 (.A(_00554_),
    .X(net3514));
 sg13g2_dlygate4sd3_1 hold2387 (.A(\TRNG.hash[136] ),
    .X(net3515));
 sg13g2_dlygate4sd3_1 hold2388 (.A(_01067_),
    .X(net3516));
 sg13g2_dlygate4sd3_1 hold2389 (.A(_00160_),
    .X(net3517));
 sg13g2_dlygate4sd3_1 hold2390 (.A(_00505_),
    .X(net3518));
 sg13g2_dlygate4sd3_1 hold2391 (.A(\TRNG.sha256.expand.data1_to_ram[13] ),
    .X(net3519));
 sg13g2_dlygate4sd3_1 hold2392 (.A(_02338_),
    .X(net3520));
 sg13g2_dlygate4sd3_1 hold2393 (.A(\TRNG.hash[192] ),
    .X(net3521));
 sg13g2_dlygate4sd3_1 hold2394 (.A(_00173_),
    .X(net3522));
 sg13g2_dlygate4sd3_1 hold2395 (.A(_02961_),
    .X(net3523));
 sg13g2_dlygate4sd3_1 hold2396 (.A(\TRNG.sha256.W[30] ),
    .X(net3524));
 sg13g2_dlygate4sd3_1 hold2397 (.A(\TRNG.raw_bit_counter[0] ),
    .X(net3525));
 sg13g2_dlygate4sd3_1 hold2398 (.A(\TRNG.hash[48] ),
    .X(net3526));
 sg13g2_dlygate4sd3_1 hold2399 (.A(_01177_),
    .X(net3527));
 sg13g2_dlygate4sd3_1 hold2400 (.A(\TRNG.sha256.expand.data1_to_ram[11] ),
    .X(net3528));
 sg13g2_dlygate4sd3_1 hold2401 (.A(\TRNG.sha256.expand.data1_to_ram[25] ),
    .X(net3529));
 sg13g2_dlygate4sd3_1 hold2402 (.A(_00226_),
    .X(net3530));
 sg13g2_dlygate4sd3_1 hold2403 (.A(_01111_),
    .X(net3531));
 sg13g2_dlygate4sd3_1 hold2404 (.A(\TRNG.sha256.expand.data1_to_ram[12] ),
    .X(net3532));
 sg13g2_dlygate4sd3_1 hold2405 (.A(_02334_),
    .X(net3533));
 sg13g2_dlygate4sd3_1 hold2406 (.A(\TRNG.hash[146] ),
    .X(net3534));
 sg13g2_dlygate4sd3_1 hold2407 (.A(_01075_),
    .X(net3535));
 sg13g2_dlygate4sd3_1 hold2408 (.A(\TRNG.hash[16] ),
    .X(net3536));
 sg13g2_dlygate4sd3_1 hold2409 (.A(_00162_),
    .X(net3537));
 sg13g2_dlygate4sd3_1 hold2410 (.A(_01169_),
    .X(net3538));
 sg13g2_dlygate4sd3_1 hold2411 (.A(\TRNG.hash[4] ),
    .X(net3539));
 sg13g2_dlygate4sd3_1 hold2412 (.A(_01187_),
    .X(net3540));
 sg13g2_dlygate4sd3_1 hold2413 (.A(_00142_),
    .X(net3541));
 sg13g2_dlygate4sd3_1 hold2414 (.A(_06974_),
    .X(net3542));
 sg13g2_dlygate4sd3_1 hold2415 (.A(_00486_),
    .X(net3543));
 sg13g2_dlygate4sd3_1 hold2416 (.A(\TRNG.chunk_index[0] ),
    .X(net3544));
 sg13g2_dlygate4sd3_1 hold2417 (.A(_02140_),
    .X(net3545));
 sg13g2_dlygate4sd3_1 hold2418 (.A(_00149_),
    .X(net3546));
 sg13g2_dlygate4sd3_1 hold2419 (.A(_06997_),
    .X(net3547));
 sg13g2_dlygate4sd3_1 hold2420 (.A(_00491_),
    .X(net3548));
 sg13g2_dlygate4sd3_1 hold2421 (.A(_00169_),
    .X(net3549));
 sg13g2_dlygate4sd3_1 hold2422 (.A(_00513_),
    .X(net3550));
 sg13g2_dlygate4sd3_1 hold2423 (.A(_00208_),
    .X(net3551));
 sg13g2_dlygate4sd3_1 hold2424 (.A(_01146_),
    .X(net3552));
 sg13g2_dlygate4sd3_1 hold2425 (.A(\TRNG.hash[80] ),
    .X(net3553));
 sg13g2_dlygate4sd3_1 hold2426 (.A(_01160_),
    .X(net3554));
 sg13g2_dlygate4sd3_1 hold2427 (.A(_00156_),
    .X(net3555));
 sg13g2_dlygate4sd3_1 hold2428 (.A(_03021_),
    .X(net3556));
 sg13g2_dlygate4sd3_1 hold2429 (.A(_01186_),
    .X(net3557));
 sg13g2_dlygate4sd3_1 hold2430 (.A(\TRNG.hash[54] ),
    .X(net3558));
 sg13g2_dlygate4sd3_1 hold2431 (.A(_07113_),
    .X(net3559));
 sg13g2_dlygate4sd3_1 hold2432 (.A(\TRNG.hash[41] ),
    .X(net3560));
 sg13g2_dlygate4sd3_1 hold2433 (.A(_07081_),
    .X(net3561));
 sg13g2_dlygate4sd3_1 hold2434 (.A(_00508_),
    .X(net3562));
 sg13g2_dlygate4sd3_1 hold2435 (.A(\TRNG.hash[162] ),
    .X(net3563));
 sg13g2_dlygate4sd3_1 hold2436 (.A(_00477_),
    .X(net3564));
 sg13g2_dlygate4sd3_1 hold2437 (.A(\TRNG.hash[65] ),
    .X(net3565));
 sg13g2_dlygate4sd3_1 hold2438 (.A(_06880_),
    .X(net3566));
 sg13g2_dlygate4sd3_1 hold2439 (.A(\TRNG.hash[194] ),
    .X(net3567));
 sg13g2_dlygate4sd3_1 hold2440 (.A(_00552_),
    .X(net3568));
 sg13g2_dlygate4sd3_1 hold2441 (.A(\TRNG.hash[250] ),
    .X(net3569));
 sg13g2_dlygate4sd3_1 hold2442 (.A(_08243_),
    .X(net3570));
 sg13g2_dlygate4sd3_1 hold2443 (.A(\TRNG.hash[53] ),
    .X(net3571));
 sg13g2_dlygate4sd3_1 hold2444 (.A(_07109_),
    .X(net3572));
 sg13g2_dlygate4sd3_1 hold2445 (.A(_00514_),
    .X(net3573));
 sg13g2_dlygate4sd3_1 hold2446 (.A(_00154_),
    .X(net3574));
 sg13g2_dlygate4sd3_1 hold2447 (.A(_00495_),
    .X(net3575));
 sg13g2_dlygate4sd3_1 hold2448 (.A(\TRNG.hash[50] ),
    .X(net3576));
 sg13g2_dlygate4sd3_1 hold2449 (.A(_07036_),
    .X(net3577));
 sg13g2_dlygate4sd3_1 hold2450 (.A(_00499_),
    .X(net3578));
 sg13g2_dlygate4sd3_1 hold2451 (.A(\TRNG.hash[180] ),
    .X(net3579));
 sg13g2_dlygate4sd3_1 hold2452 (.A(_08160_),
    .X(net3580));
 sg13g2_dlygate4sd3_1 hold2453 (.A(\TRNG.hash[85] ),
    .X(net3581));
 sg13g2_dlygate4sd3_1 hold2454 (.A(_07186_),
    .X(net3582));
 sg13g2_dlygate4sd3_1 hold2455 (.A(_00151_),
    .X(net3583));
 sg13g2_dlygate4sd3_1 hold2456 (.A(_00492_),
    .X(net3584));
 sg13g2_dlygate4sd3_1 hold2457 (.A(\TRNG.hash[43] ),
    .X(net3585));
 sg13g2_dlygate4sd3_1 hold2458 (.A(_01173_),
    .X(net3586));
 sg13g2_dlygate4sd3_1 hold2459 (.A(\TRNG.hash[51] ),
    .X(net3587));
 sg13g2_dlygate4sd3_1 hold2460 (.A(_07102_),
    .X(net3588));
 sg13g2_dlygate4sd3_1 hold2461 (.A(\TRNG.Padded_Out[67] ),
    .X(net3589));
 sg13g2_dlygate4sd3_1 hold2462 (.A(\TRNG.sha256.W[27] ),
    .X(net3590));
 sg13g2_dlygate4sd3_1 hold2463 (.A(_00203_),
    .X(net3591));
 sg13g2_dlygate4sd3_1 hold2464 (.A(_07957_),
    .X(net3592));
 sg13g2_dlygate4sd3_1 hold2465 (.A(_00547_),
    .X(net3593));
 sg13g2_dlygate4sd3_1 hold2466 (.A(\TRNG.hash[44] ),
    .X(net3594));
 sg13g2_dlygate4sd3_1 hold2467 (.A(_01174_),
    .X(net3595));
 sg13g2_dlygate4sd3_1 hold2468 (.A(\TRNG.sha256.compress.count[3] ),
    .X(net3596));
 sg13g2_dlygate4sd3_1 hold2469 (.A(_00933_),
    .X(net3597));
 sg13g2_dlygate4sd3_1 hold2470 (.A(\TRNG.hash[61] ),
    .X(net3598));
 sg13g2_dlygate4sd3_1 hold2471 (.A(_07057_),
    .X(net3599));
 sg13g2_dlygate4sd3_1 hold2472 (.A(_00503_),
    .X(net3600));
 sg13g2_dlygate4sd3_1 hold2473 (.A(_00185_),
    .X(net3601));
 sg13g2_dlygate4sd3_1 hold2474 (.A(_07170_),
    .X(net3602));
 sg13g2_dlygate4sd3_1 hold2475 (.A(_00527_),
    .X(net3603));
 sg13g2_dlygate4sd3_1 hold2476 (.A(\TRNG.hash[78] ),
    .X(net3604));
 sg13g2_dlygate4sd3_1 hold2477 (.A(_01159_),
    .X(net3605));
 sg13g2_dlygate4sd3_1 hold2478 (.A(\TRNG.hash[79] ),
    .X(net3606));
 sg13g2_dlygate4sd3_1 hold2479 (.A(_01176_),
    .X(net3607));
 sg13g2_dlygate4sd3_1 hold2480 (.A(\TRNG.hash[87] ),
    .X(net3608));
 sg13g2_dlygate4sd3_1 hold2481 (.A(_00532_),
    .X(net3609));
 sg13g2_dlygate4sd3_1 hold2482 (.A(\TRNG.hash[64] ),
    .X(net3610));
 sg13g2_dlygate4sd3_1 hold2483 (.A(_06881_),
    .X(net3611));
 sg13g2_dlygate4sd3_1 hold2484 (.A(\TRNG.hash[20] ),
    .X(net3612));
 sg13g2_dlygate4sd3_1 hold2485 (.A(_07045_),
    .X(net3613));
 sg13g2_dlygate4sd3_1 hold2486 (.A(\TRNG.hash[46] ),
    .X(net3614));
 sg13g2_dlygate4sd3_1 hold2487 (.A(_01191_),
    .X(net3615));
 sg13g2_dlygate4sd3_1 hold2488 (.A(\TRNG.hash[149] ),
    .X(net3616));
 sg13g2_dlygate4sd3_1 hold2489 (.A(_06958_),
    .X(net3617));
 sg13g2_dlygate4sd3_1 hold2490 (.A(_00483_),
    .X(net3618));
 sg13g2_dlygate4sd3_1 hold2491 (.A(_00198_),
    .X(net3619));
 sg13g2_dlygate4sd3_1 hold2492 (.A(\TRNG.hash[9] ),
    .X(net3620));
 sg13g2_dlygate4sd3_1 hold2493 (.A(_00494_),
    .X(net3621));
 sg13g2_dlygate4sd3_1 hold2494 (.A(\TRNG.sha256.expand.data1_to_ram[7] ),
    .X(net3622));
 sg13g2_dlygate4sd3_1 hold2495 (.A(_02317_),
    .X(net3623));
 sg13g2_dlygate4sd3_1 hold2496 (.A(\TRNG.hash[140] ),
    .X(net3624));
 sg13g2_dlygate4sd3_1 hold2497 (.A(_02513_),
    .X(net3625));
 sg13g2_dlygate4sd3_1 hold2498 (.A(\TRNG.sha256.expand.data1_to_ram[9] ),
    .X(net3626));
 sg13g2_dlygate4sd3_1 hold2499 (.A(_02324_),
    .X(net3627));
 sg13g2_dlygate4sd3_1 hold2500 (.A(_00153_),
    .X(net3628));
 sg13g2_dlygate4sd3_1 hold2501 (.A(_01188_),
    .X(net3629));
 sg13g2_dlygate4sd3_1 hold2502 (.A(\TRNG.hash[131] ),
    .X(net3630));
 sg13g2_dlygate4sd3_1 hold2503 (.A(_01064_),
    .X(net3631));
 sg13g2_dlygate4sd3_1 hold2504 (.A(\TRNG.sha256.expand.data1_to_ram[22] ),
    .X(net3632));
 sg13g2_dlygate4sd3_1 hold2505 (.A(_02369_),
    .X(net3633));
 sg13g2_dlygate4sd3_1 hold2506 (.A(\TRNG.hash[60] ),
    .X(net3634));
 sg13g2_dlygate4sd3_1 hold2507 (.A(_01184_),
    .X(net3635));
 sg13g2_dlygate4sd3_1 hold2508 (.A(\TRNG.hash[208] ),
    .X(net3636));
 sg13g2_dlygate4sd3_1 hold2509 (.A(_01108_),
    .X(net3637));
 sg13g2_dlygate4sd3_1 hold2510 (.A(\TRNG.sha256.expand.data1_to_ram[31] ),
    .X(net3638));
 sg13g2_dlygate4sd3_1 hold2511 (.A(_02401_),
    .X(net3639));
 sg13g2_dlygate4sd3_1 hold2512 (.A(\TRNG.Padded_Out[64] ),
    .X(net3640));
 sg13g2_dlygate4sd3_1 hold2513 (.A(\TRNG.sha256.expand.data1_to_ram[10] ),
    .X(net3641));
 sg13g2_dlygate4sd3_1 hold2514 (.A(_02327_),
    .X(net3642));
 sg13g2_dlygate4sd3_1 hold2515 (.A(_00135_),
    .X(net3643));
 sg13g2_dlygate4sd3_1 hold2516 (.A(_01066_),
    .X(net3644));
 sg13g2_dlygate4sd3_1 hold2517 (.A(_00140_),
    .X(net3645));
 sg13g2_dlygate4sd3_1 hold2518 (.A(_01077_),
    .X(net3646));
 sg13g2_dlygate4sd3_1 hold2519 (.A(\TRNG.hash[176] ),
    .X(net3647));
 sg13g2_dlygate4sd3_1 hold2520 (.A(\TRNG.hash[139] ),
    .X(net3648));
 sg13g2_dlygate4sd3_1 hold2521 (.A(_06944_),
    .X(net3649));
 sg13g2_dlygate4sd3_1 hold2522 (.A(_00481_),
    .X(net3650));
 sg13g2_dlygate4sd3_1 hold2523 (.A(\TRNG.sha256.compress.count[2] ),
    .X(net3651));
 sg13g2_dlygate4sd3_1 hold2524 (.A(_00932_),
    .X(net3652));
 sg13g2_dlygate4sd3_1 hold2525 (.A(\TRNG.sha256.expand.address1[1] ),
    .X(net3653));
 sg13g2_dlygate4sd3_1 hold2526 (.A(_00155_),
    .X(net3654));
 sg13g2_dlygate4sd3_1 hold2527 (.A(\TRNG.hash[147] ),
    .X(net3655));
 sg13g2_dlygate4sd3_1 hold2528 (.A(_01076_),
    .X(net3656));
 sg13g2_dlygate4sd3_1 hold2529 (.A(\TRNG.sha256.expand.data1_to_ram[8] ),
    .X(net3657));
 sg13g2_dlygate4sd3_1 hold2530 (.A(_02321_),
    .X(net3658));
 sg13g2_dlygate4sd3_1 hold2531 (.A(_00202_),
    .X(net3659));
 sg13g2_dlygate4sd3_1 hold2532 (.A(_00548_),
    .X(net3660));
 sg13g2_dlygate4sd3_1 hold2533 (.A(\TRNG.sha256.expand.exp_ctrl.j[0] ),
    .X(net3661));
 sg13g2_dlygate4sd3_1 hold2534 (.A(_02268_),
    .X(net3662));
 sg13g2_dlygate4sd3_1 hold2535 (.A(_00930_),
    .X(net3663));
 sg13g2_dlygate4sd3_1 hold2536 (.A(\TRNG.Padded_Out[151] ),
    .X(net3664));
 sg13g2_dlygate4sd3_1 hold2537 (.A(\TRNG.hash[138] ),
    .X(net3665));
 sg13g2_dlygate4sd3_1 hold2538 (.A(_01068_),
    .X(net3666));
 sg13g2_dlygate4sd3_1 hold2539 (.A(_00196_),
    .X(net3667));
 sg13g2_dlygate4sd3_1 hold2540 (.A(_01162_),
    .X(net3668));
 sg13g2_dlygate4sd3_1 hold2541 (.A(\TRNG.hash[40] ),
    .X(net3669));
 sg13g2_dlygate4sd3_1 hold2542 (.A(_02966_),
    .X(net3670));
 sg13g2_dlygate4sd3_1 hold2543 (.A(\TRNG.sha256.expand.data1_to_ram[23] ),
    .X(net3671));
 sg13g2_dlygate4sd3_1 hold2544 (.A(_02372_),
    .X(net3672));
 sg13g2_dlygate4sd3_1 hold2545 (.A(\TRNG.sha256.expand.data1_to_ram[26] ),
    .X(net3673));
 sg13g2_dlygate4sd3_1 hold2546 (.A(_02381_),
    .X(net3674));
 sg13g2_dlygate4sd3_1 hold2547 (.A(\TRNG.hash[145] ),
    .X(net3675));
 sg13g2_dlygate4sd3_1 hold2548 (.A(_01074_),
    .X(net3676));
 sg13g2_dlygate4sd3_1 hold2549 (.A(_00159_),
    .X(net3677));
 sg13g2_dlygate4sd3_1 hold2550 (.A(_03053_),
    .X(net3678));
 sg13g2_dlygate4sd3_1 hold2551 (.A(\TRNG.hash[49] ),
    .X(net3679));
 sg13g2_dlygate4sd3_1 hold2552 (.A(_01178_),
    .X(net3680));
 sg13g2_dlygate4sd3_1 hold2553 (.A(\TRNG.hash[157] ),
    .X(net3681));
 sg13g2_dlygate4sd3_1 hold2554 (.A(_02553_),
    .X(net3682));
 sg13g2_dlygate4sd3_1 hold2555 (.A(\TRNG.hash[45] ),
    .X(net3683));
 sg13g2_dlygate4sd3_1 hold2556 (.A(\TRNG.hash[177] ),
    .X(net3684));
 sg13g2_dlygate4sd3_1 hold2557 (.A(_01129_),
    .X(net3685));
 sg13g2_dlygate4sd3_1 hold2558 (.A(\TRNG.hash[167] ),
    .X(net3686));
 sg13g2_dlygate4sd3_1 hold2559 (.A(\TRNG.sha256.expand.data1_to_ram[30] ),
    .X(net3687));
 sg13g2_dlygate4sd3_1 hold2560 (.A(_02397_),
    .X(net3688));
 sg13g2_dlygate4sd3_1 hold2561 (.A(\TRNG.hash[34] ),
    .X(net3689));
 sg13g2_dlygate4sd3_1 hold2562 (.A(_06994_),
    .X(net3690));
 sg13g2_dlygate4sd3_1 hold2563 (.A(_00490_),
    .X(net3691));
 sg13g2_dlygate4sd3_1 hold2564 (.A(\TRNG.hash[181] ),
    .X(net3692));
 sg13g2_dlygate4sd3_1 hold2565 (.A(_02781_),
    .X(net3693));
 sg13g2_dlygate4sd3_1 hold2566 (.A(\TRNG.hash[55] ),
    .X(net3694));
 sg13g2_dlygate4sd3_1 hold2567 (.A(_02996_),
    .X(net3695));
 sg13g2_dlygate4sd3_1 hold2568 (.A(\TRNG.uart_tx_inst.ticks_counter[3] ),
    .X(net3696));
 sg13g2_dlygate4sd3_1 hold2569 (.A(\TRNG.Padded_Out[203] ),
    .X(net3697));
 sg13g2_dlygate4sd3_1 hold2570 (.A(\TRNG.sha256.expand.data1_to_ram[16] ),
    .X(net3698));
 sg13g2_dlygate4sd3_1 hold2571 (.A(\TRNG.hash[152] ),
    .X(net3699));
 sg13g2_dlygate4sd3_1 hold2572 (.A(_02545_),
    .X(net3700));
 sg13g2_dlygate4sd3_1 hold2573 (.A(\TRNG.sha256.expand.data1_to_ram[6] ),
    .X(net3701));
 sg13g2_dlygate4sd3_1 hold2574 (.A(_02313_),
    .X(net3702));
 sg13g2_dlygate4sd3_1 hold2575 (.A(\TRNG.hash[194] ),
    .X(net3703));
 sg13g2_dlygate4sd3_1 hold2576 (.A(\TRNG.hash[13] ),
    .X(net3704));
 sg13g2_dlygate4sd3_1 hold2577 (.A(_00496_),
    .X(net3705));
 sg13g2_dlygate4sd3_1 hold2578 (.A(\TRNG.sha256.expand.data1_to_ram[24] ),
    .X(net3706));
 sg13g2_dlygate4sd3_1 hold2579 (.A(_02375_),
    .X(net3707));
 sg13g2_dlygate4sd3_1 hold2580 (.A(\TRNG.Padded_Out[201] ),
    .X(net3708));
 sg13g2_dlygate4sd3_1 hold2581 (.A(_09001_),
    .X(net3709));
 sg13g2_dlygate4sd3_1 hold2582 (.A(_00199_),
    .X(net3710));
 sg13g2_dlygate4sd3_1 hold2583 (.A(_08073_),
    .X(net3711));
 sg13g2_dlygate4sd3_1 hold2584 (.A(\TRNG.hash[154] ),
    .X(net3712));
 sg13g2_dlygate4sd3_1 hold2585 (.A(_02549_),
    .X(net3713));
 sg13g2_dlygate4sd3_1 hold2586 (.A(_00220_),
    .X(net3714));
 sg13g2_dlygate4sd3_1 hold2587 (.A(_01148_),
    .X(net3715));
 sg13g2_dlygate4sd3_1 hold2588 (.A(_00232_),
    .X(net3716));
 sg13g2_dlygate4sd3_1 hold2589 (.A(\TRNG.hash[83] ),
    .X(net3717));
 sg13g2_dlygate4sd3_1 hold2590 (.A(\TRNG.hash[144] ),
    .X(net3718));
 sg13g2_dlygate4sd3_1 hold2591 (.A(_02528_),
    .X(net3719));
 sg13g2_dlygate4sd3_1 hold2592 (.A(\TRNG.sha256.expand.data1_to_ram[21] ),
    .X(net3720));
 sg13g2_dlygate4sd3_1 hold2593 (.A(_02365_),
    .X(net3721));
 sg13g2_dlygate4sd3_1 hold2594 (.A(\TRNG.hash[62] ),
    .X(net3722));
 sg13g2_dlygate4sd3_1 hold2595 (.A(_07127_),
    .X(net3723));
 sg13g2_dlygate4sd3_1 hold2596 (.A(\TRNG.hash[95] ),
    .X(net3724));
 sg13g2_dlygate4sd3_1 hold2597 (.A(_07130_),
    .X(net3725));
 sg13g2_dlygate4sd3_1 hold2598 (.A(\TRNG.Padded_Out[152] ),
    .X(net3726));
 sg13g2_dlygate4sd3_1 hold2599 (.A(\TRNG.uart_tx_inst.ticks_counter[4] ),
    .X(net3727));
 sg13g2_dlygate4sd3_1 hold2600 (.A(\TRNG.hash[22] ),
    .X(net3728));
 sg13g2_dlygate4sd3_1 hold2601 (.A(\TRNG.hash[165] ),
    .X(net3729));
 sg13g2_dlygate4sd3_1 hold2602 (.A(_01121_),
    .X(net3730));
 sg13g2_dlygate4sd3_1 hold2603 (.A(\TRNG.hash[195] ),
    .X(net3731));
 sg13g2_dlygate4sd3_1 hold2604 (.A(_00553_),
    .X(net3732));
 sg13g2_dlygate4sd3_1 hold2605 (.A(\TRNG.hash[71] ),
    .X(net3733));
 sg13g2_dlygate4sd3_1 hold2606 (.A(_02900_),
    .X(net3734));
 sg13g2_dlygate4sd3_1 hold2607 (.A(\TRNG.hash[28] ),
    .X(net3735));
 sg13g2_dlygate4sd3_1 hold2608 (.A(\TRNG.hash[227] ),
    .X(net3736));
 sg13g2_dlygate4sd3_1 hold2609 (.A(\TRNG.Padded_Out[288] ),
    .X(net3737));
 sg13g2_dlygate4sd3_1 hold2610 (.A(\TRNG.hash[74] ),
    .X(net3738));
 sg13g2_dlygate4sd3_1 hold2611 (.A(_00524_),
    .X(net3739));
 sg13g2_dlygate4sd3_1 hold2612 (.A(_00215_),
    .X(net3740));
 sg13g2_dlygate4sd3_1 hold2613 (.A(_00234_),
    .X(net3741));
 sg13g2_dlygate4sd3_1 hold2614 (.A(_01096_),
    .X(net3742));
 sg13g2_dlygate4sd3_1 hold2615 (.A(\TRNG.sha256.expand.data1_to_ram[14] ),
    .X(net3743));
 sg13g2_dlygate4sd3_1 hold2616 (.A(_02342_),
    .X(net3744));
 sg13g2_dlygate4sd3_1 hold2617 (.A(\TRNG.hash[33] ),
    .X(net3745));
 sg13g2_dlygate4sd3_1 hold2618 (.A(_00489_),
    .X(net3746));
 sg13g2_dlygate4sd3_1 hold2619 (.A(\TRNG.hash[10] ),
    .X(net3747));
 sg13g2_dlygate4sd3_1 hold2620 (.A(_03036_),
    .X(net3748));
 sg13g2_dlygate4sd3_1 hold2621 (.A(\TRNG.sha256.expand.exp_ctrl.j_2[0] ),
    .X(net3749));
 sg13g2_dlygate4sd3_1 hold2622 (.A(_00206_),
    .X(net3750));
 sg13g2_dlygate4sd3_1 hold2623 (.A(_02841_),
    .X(net3751));
 sg13g2_dlygate4sd3_1 hold2624 (.A(_01145_),
    .X(net3752));
 sg13g2_dlygate4sd3_1 hold2625 (.A(\TRNG.hash[31] ),
    .X(net3753));
 sg13g2_dlygate4sd3_1 hold2626 (.A(_07061_),
    .X(net3754));
 sg13g2_dlygate4sd3_1 hold2627 (.A(_00504_),
    .X(net3755));
 sg13g2_dlygate4sd3_1 hold2628 (.A(\TRNG.sha256.compress.hash_gen.temp[4] ),
    .X(net3756));
 sg13g2_dlygate4sd3_1 hold2629 (.A(_00118_),
    .X(net3757));
 sg13g2_dlygate4sd3_1 hold2630 (.A(_01167_),
    .X(net3758));
 sg13g2_dlygate4sd3_1 hold2631 (.A(\TRNG.hash[143] ),
    .X(net3759));
 sg13g2_dlygate4sd3_1 hold2632 (.A(\TRNG.hash[202] ),
    .X(net3760));
 sg13g2_dlygate4sd3_1 hold2633 (.A(\TRNG.hash[26] ),
    .X(net3761));
 sg13g2_dlygate4sd3_1 hold2634 (.A(_07052_),
    .X(net3762));
 sg13g2_dlygate4sd3_1 hold2635 (.A(\TRNG.hash[58] ),
    .X(net3763));
 sg13g2_dlygate4sd3_1 hold2636 (.A(_03009_),
    .X(net3764));
 sg13g2_dlygate4sd3_1 hold2637 (.A(_00146_),
    .X(net3765));
 sg13g2_dlygate4sd3_1 hold2638 (.A(_02485_),
    .X(net3766));
 sg13g2_dlygate4sd3_1 hold2639 (.A(_00231_),
    .X(net3767));
 sg13g2_dlygate4sd3_1 hold2640 (.A(\TRNG.hash[11] ),
    .X(net3768));
 sg13g2_dlygate4sd3_1 hold2641 (.A(_00164_),
    .X(net3769));
 sg13g2_dlygate4sd3_1 hold2642 (.A(_02956_),
    .X(net3770));
 sg13g2_dlygate4sd3_1 hold2643 (.A(_01170_),
    .X(net3771));
 sg13g2_dlygate4sd3_1 hold2644 (.A(\TRNG.hash[159] ),
    .X(net3772));
 sg13g2_dlygate4sd3_1 hold2645 (.A(\TRNG.hash[170] ),
    .X(net3773));
 sg13g2_dlygate4sd3_1 hold2646 (.A(_00555_),
    .X(net3774));
 sg13g2_dlygate4sd3_1 hold2647 (.A(\TRNG.hash[59] ),
    .X(net3775));
 sg13g2_dlygate4sd3_1 hold2648 (.A(_03013_),
    .X(net3776));
 sg13g2_dlygate4sd3_1 hold2649 (.A(\TRNG.hash[179] ),
    .X(net3777));
 sg13g2_dlygate4sd3_1 hold2650 (.A(\TRNG.hash[222] ),
    .X(net3778));
 sg13g2_dlygate4sd3_1 hold2651 (.A(_08181_),
    .X(net3779));
 sg13g2_dlygate4sd3_1 hold2652 (.A(\TRNG.Padded_Out[480] ),
    .X(net3780));
 sg13g2_dlygate4sd3_1 hold2653 (.A(\TRNG.hash[91] ),
    .X(net3781));
 sg13g2_dlygate4sd3_1 hold2654 (.A(_02935_),
    .X(net3782));
 sg13g2_dlygate4sd3_1 hold2655 (.A(_00235_),
    .X(net3783));
 sg13g2_dlygate4sd3_1 hold2656 (.A(\TRNG.hash[214] ),
    .X(net3784));
 sg13g2_dlygate4sd3_1 hold2657 (.A(_01133_),
    .X(net3785));
 sg13g2_dlygate4sd3_1 hold2658 (.A(\TRNG.hash[216] ),
    .X(net3786));
 sg13g2_dlygate4sd3_1 hold2659 (.A(_01113_),
    .X(net3787));
 sg13g2_dlygate4sd3_1 hold2660 (.A(_00236_),
    .X(net3788));
 sg13g2_dlygate4sd3_1 hold2661 (.A(_01098_),
    .X(net3789));
 sg13g2_dlygate4sd3_1 hold2662 (.A(\TRNG.sha256.expand.sm0.sum_0[0] ),
    .X(net3790));
 sg13g2_dlygate4sd3_1 hold2663 (.A(_06597_),
    .X(net3791));
 sg13g2_dlygate4sd3_1 hold2664 (.A(\TRNG.hash[210] ),
    .X(net3792));
 sg13g2_dlygate4sd3_1 hold2665 (.A(\TRNG.hash[153] ),
    .X(net3793));
 sg13g2_dlygate4sd3_1 hold2666 (.A(_06972_),
    .X(net3794));
 sg13g2_dlygate4sd3_1 hold2667 (.A(_00233_),
    .X(net3795));
 sg13g2_dlygate4sd3_1 hold2668 (.A(_01095_),
    .X(net3796));
 sg13g2_dlygate4sd3_1 hold2669 (.A(\TRNG.Padded_Out[209] ),
    .X(net3797));
 sg13g2_dlygate4sd3_1 hold2670 (.A(\TRNG.hash[173] ),
    .X(net3798));
 sg13g2_dlygate4sd3_1 hold2671 (.A(\TRNG.hash[211] ),
    .X(net3799));
 sg13g2_dlygate4sd3_1 hold2672 (.A(_08227_),
    .X(net3800));
 sg13g2_dlygate4sd3_1 hold2673 (.A(\TRNG.hash[191] ),
    .X(net3801));
 sg13g2_dlygate4sd3_1 hold2674 (.A(_08184_),
    .X(net3802));
 sg13g2_dlygate4sd3_1 hold2675 (.A(\TRNG.hash[88] ),
    .X(net3803));
 sg13g2_dlygate4sd3_1 hold2676 (.A(_01180_),
    .X(net3804));
 sg13g2_dlygate4sd3_1 hold2677 (.A(\TRNG.hash[183] ),
    .X(net3805));
 sg13g2_dlygate4sd3_1 hold2678 (.A(_08166_),
    .X(net3806));
 sg13g2_dlygate4sd3_1 hold2679 (.A(\TRNG.sha256.compress.hash_gen.w_rdy ),
    .X(net3807));
 sg13g2_dlygate4sd3_1 hold2680 (.A(\TRNG.hash[206] ),
    .X(net3808));
 sg13g2_dlygate4sd3_1 hold2681 (.A(\TRNG.hash[73] ),
    .X(net3809));
 sg13g2_dlygate4sd3_1 hold2682 (.A(_00523_),
    .X(net3810));
 sg13g2_dlygate4sd3_1 hold2683 (.A(\TRNG.Padded_Out[181] ),
    .X(net3811));
 sg13g2_dlygate4sd3_1 hold2684 (.A(_09137_),
    .X(net3812));
 sg13g2_dlygate4sd3_1 hold2685 (.A(\TRNG.hash[23] ),
    .X(net3813));
 sg13g2_dlygate4sd3_1 hold2686 (.A(\TRNG.hash[217] ),
    .X(net3814));
 sg13g2_dlygate4sd3_1 hold2687 (.A(\TRNG.hash[89] ),
    .X(net3815));
 sg13g2_dlygate4sd3_1 hold2688 (.A(\TRNG.sha256.expand.exp_ctrl.final_sum[27] ),
    .X(net3816));
 sg13g2_dlygate4sd3_1 hold2689 (.A(\TRNG.sha256.compress.count[1] ),
    .X(net3817));
 sg13g2_dlygate4sd3_1 hold2690 (.A(\TRNG.hash[168] ),
    .X(net3818));
 sg13g2_dlygate4sd3_1 hold2691 (.A(\TRNG.sha256.W[20] ),
    .X(net3819));
 sg13g2_dlygate4sd3_1 hold2692 (.A(\TRNG.hash[27] ),
    .X(net3820));
 sg13g2_dlygate4sd3_1 hold2693 (.A(\TRNG.hash[92] ),
    .X(net3821));
 sg13g2_dlygate4sd3_1 hold2694 (.A(_01165_),
    .X(net3822));
 sg13g2_dlygate4sd3_1 hold2695 (.A(\TRNG.hash[184] ),
    .X(net3823));
 sg13g2_dlygate4sd3_1 hold2696 (.A(\TRNG.hash[70] ),
    .X(net3824));
 sg13g2_dlygate4sd3_1 hold2697 (.A(_00521_),
    .X(net3825));
 sg13g2_dlygate4sd3_1 hold2698 (.A(\TRNG.sha256.control.iteration[7] ),
    .X(net3826));
 sg13g2_dlygate4sd3_1 hold2699 (.A(_02483_),
    .X(net3827));
 sg13g2_dlygate4sd3_1 hold2700 (.A(\TRNG.hash[214] ),
    .X(net3828));
 sg13g2_dlygate4sd3_1 hold2701 (.A(\TRNG.hash[24] ),
    .X(net3829));
 sg13g2_dlygate4sd3_1 hold2702 (.A(\TRNG.hash[189] ),
    .X(net3830));
 sg13g2_dlygate4sd3_1 hold2703 (.A(_01137_),
    .X(net3831));
 sg13g2_dlygate4sd3_1 hold2704 (.A(\TRNG.hash[207] ),
    .X(net3832));
 sg13g2_dlygate4sd3_1 hold2705 (.A(_00237_),
    .X(net3833));
 sg13g2_dlygate4sd3_1 hold2706 (.A(\TRNG.hash[25] ),
    .X(net3834));
 sg13g2_dlygate4sd3_1 hold2707 (.A(\TRNG.hash[67] ),
    .X(net3835));
 sg13g2_dlygate4sd3_1 hold2708 (.A(_01155_),
    .X(net3836));
 sg13g2_dlygate4sd3_1 hold2709 (.A(\TRNG.hash[94] ),
    .X(net3837));
 sg13g2_dlygate4sd3_1 hold2710 (.A(\TRNG.hash[204] ),
    .X(net3838));
 sg13g2_dlygate4sd3_1 hold2711 (.A(_08214_),
    .X(net3839));
 sg13g2_dlygate4sd3_1 hold2712 (.A(\TRNG.hash[175] ),
    .X(net3840));
 sg13g2_dlygate4sd3_1 hold2713 (.A(\TRNG.hash[69] ),
    .X(net3841));
 sg13g2_dlygate4sd3_1 hold2714 (.A(\TRNG.hash[142] ),
    .X(net3842));
 sg13g2_dlygate4sd3_1 hold2715 (.A(_01071_),
    .X(net3843));
 sg13g2_dlygate4sd3_1 hold2716 (.A(\TRNG.hash[209] ),
    .X(net3844));
 sg13g2_dlygate4sd3_1 hold2717 (.A(\TRNG.hash[203] ),
    .X(net3845));
 sg13g2_dlygate4sd3_1 hold2718 (.A(\TRNG.hash[223] ),
    .X(net3846));
 sg13g2_dlygate4sd3_1 hold2719 (.A(\TRNG.sha256.expand.exp_ctrl.final_sum[4] ),
    .X(net3847));
 sg13g2_dlygate4sd3_1 hold2720 (.A(\TRNG.hash[166] ),
    .X(net3848));
 sg13g2_dlygate4sd3_1 hold2721 (.A(\TRNG.hash[172] ),
    .X(net3849));
 sg13g2_dlygate4sd3_1 hold2722 (.A(\TRNG.hash[57] ),
    .X(net3850));
 sg13g2_dlygate4sd3_1 hold2723 (.A(_03005_),
    .X(net3851));
 sg13g2_dlygate4sd3_1 hold2724 (.A(\TRNG.hash[132] ),
    .X(net3852));
 sg13g2_dlygate4sd3_1 hold2725 (.A(_01065_),
    .X(net3853));
 sg13g2_dlygate4sd3_1 hold2726 (.A(\TRNG.hash[151] ),
    .X(net3854));
 sg13g2_dlygate4sd3_1 hold2727 (.A(_00131_),
    .X(net3855));
 sg13g2_dlygate4sd3_1 hold2728 (.A(\TRNG.hash[17] ),
    .X(net3856));
 sg13g2_dlygate4sd3_1 hold2729 (.A(\TRNG.hash[174] ),
    .X(net3857));
 sg13g2_dlygate4sd3_1 hold2730 (.A(\TRNG.hash[15] ),
    .X(net3858));
 sg13g2_dlygate4sd3_1 hold2731 (.A(_03049_),
    .X(net3859));
 sg13g2_dlygate4sd3_1 hold2732 (.A(\TRNG.hash[178] ),
    .X(net3860));
 sg13g2_dlygate4sd3_1 hold2733 (.A(\TRNG.hash[185] ),
    .X(net3861));
 sg13g2_dlygate4sd3_1 hold2734 (.A(\TRNG.hash[30] ),
    .X(net3862));
 sg13g2_dlygate4sd3_1 hold2735 (.A(\TRNG.hash[197] ),
    .X(net3863));
 sg13g2_dlygate4sd3_1 hold2736 (.A(_00567_),
    .X(net3864));
 sg13g2_dlygate4sd3_1 hold2737 (.A(\TRNG.hash[242] ),
    .X(net3865));
 sg13g2_dlygate4sd3_1 hold2738 (.A(\TRNG.hash[220] ),
    .X(net3866));
 sg13g2_dlygate4sd3_1 hold2739 (.A(\TRNG.hash[110] ),
    .X(net3867));
 sg13g2_dlygate4sd3_1 hold2740 (.A(\TRNG.hash[219] ),
    .X(net3868));
 sg13g2_dlygate4sd3_1 hold2741 (.A(_01135_),
    .X(net3869));
 sg13g2_dlygate4sd3_1 hold2742 (.A(\TRNG.state[0] ),
    .X(net3870));
 sg13g2_dlygate4sd3_1 hold2743 (.A(\TRNG.hash[112] ),
    .X(net3871));
 sg13g2_dlygate4sd3_1 hold2744 (.A(\TRNG.hash[196] ),
    .X(net3872));
 sg13g2_dlygate4sd3_1 hold2745 (.A(_00566_),
    .X(net3873));
 sg13g2_dlygate4sd3_1 hold2746 (.A(\TRNG.hash[19] ),
    .X(net3874));
 sg13g2_dlygate4sd3_1 hold2747 (.A(\TRNG.hash[232] ),
    .X(net3875));
 sg13g2_dlygate4sd3_1 hold2748 (.A(_00569_),
    .X(net3876));
 sg13g2_dlygate4sd3_1 hold2749 (.A(\TRNG.hash[104] ),
    .X(net3877));
 sg13g2_dlygate4sd3_1 hold2750 (.A(\TRNG.hash[198] ),
    .X(net3878));
 sg13g2_dlygate4sd3_1 hold2751 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][20] ),
    .X(net3879));
 sg13g2_dlygate4sd3_1 hold2752 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][18] ),
    .X(net3880));
 sg13g2_dlygate4sd3_1 hold2753 (.A(_00073_),
    .X(net3881));
 sg13g2_dlygate4sd3_1 hold2754 (.A(\TRNG.hash[248] ),
    .X(net3882));
 sg13g2_dlygate4sd3_1 hold2755 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][20] ),
    .X(net3883));
 sg13g2_dlygate4sd3_1 hold2756 (.A(_05202_),
    .X(net3884));
 sg13g2_dlygate4sd3_1 hold2757 (.A(_05204_),
    .X(net3885));
 sg13g2_dlygate4sd3_1 hold2758 (.A(_00119_),
    .X(net3886));
 sg13g2_dlygate4sd3_1 hold2759 (.A(\TRNG.hash[221] ),
    .X(net3887));
 sg13g2_dlygate4sd3_1 hold2760 (.A(\TRNG.hash[171] ),
    .X(net3888));
 sg13g2_dlygate4sd3_1 hold2761 (.A(\TRNG.sha256.compress.count[4] ),
    .X(net3889));
 sg13g2_dlygate4sd3_1 hold2762 (.A(\TRNG.sha256.expand.msg_schdl.RAM[1][23] ),
    .X(net3890));
 sg13g2_dlygate4sd3_1 hold2763 (.A(_00079_),
    .X(net3891));
 sg13g2_dlygate4sd3_1 hold2764 (.A(\TRNG.hash[117] ),
    .X(net3892));
 sg13g2_dlygate4sd3_1 hold2765 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][28] ),
    .X(net3893));
 sg13g2_dlygate4sd3_1 hold2766 (.A(_05300_),
    .X(net3894));
 sg13g2_dlygate4sd3_1 hold2767 (.A(\TRNG.hash[109] ),
    .X(net3895));
 sg13g2_dlygate4sd3_1 hold2768 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][12] ),
    .X(net3896));
 sg13g2_dlygate4sd3_1 hold2769 (.A(\TRNG.hash[193] ),
    .X(net3897));
 sg13g2_dlygate4sd3_1 hold2770 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][27] ),
    .X(net3898));
 sg13g2_dlygate4sd3_1 hold2771 (.A(\TRNG.sha256.expand.msg_schdl.RAM[6][30] ),
    .X(net3899));
 sg13g2_dlygate4sd3_1 hold2772 (.A(_05330_),
    .X(net3900));
 sg13g2_dlygate4sd3_1 hold2773 (.A(\TRNG.hash[246] ),
    .X(net3901));
 sg13g2_dlygate4sd3_1 hold2774 (.A(\TRNG.sha256.expand.msg_schdl.RAM[13][6] ),
    .X(net3902));
 sg13g2_dlygate4sd3_1 hold2775 (.A(_05043_),
    .X(net3903));
 sg13g2_dlygate4sd3_1 hold2776 (.A(_05045_),
    .X(net3904));
 sg13g2_dlygate4sd3_1 hold2777 (.A(_00092_),
    .X(net3905));
 sg13g2_dlygate4sd3_1 hold2778 (.A(\TRNG.hash[241] ),
    .X(net3906));
 sg13g2_dlygate4sd3_1 hold2779 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][7] ),
    .X(net3907));
 sg13g2_dlygate4sd3_1 hold2780 (.A(_00093_),
    .X(net3908));
 sg13g2_dlygate4sd3_1 hold2781 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][5] ),
    .X(net3909));
 sg13g2_dlygate4sd3_1 hold2782 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][14] ),
    .X(net3910));
 sg13g2_dlygate4sd3_1 hold2783 (.A(_05139_),
    .X(net3911));
 sg13g2_dlygate4sd3_1 hold2784 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][17] ),
    .X(net3912));
 sg13g2_dlygate4sd3_1 hold2785 (.A(_05177_),
    .X(net3913));
 sg13g2_dlygate4sd3_1 hold2786 (.A(_00072_),
    .X(net3914));
 sg13g2_dlygate4sd3_1 hold2787 (.A(\TRNG.sha256.expand.msg_schdl.RAM[11][1] ),
    .X(net3915));
 sg13g2_dlygate4sd3_1 hold2788 (.A(_04985_),
    .X(net3916));
 sg13g2_dlygate4sd3_1 hold2789 (.A(_00075_),
    .X(net3917));
 sg13g2_dlygate4sd3_1 hold2790 (.A(\TRNG.hash[236] ),
    .X(net3918));
 sg13g2_dlygate4sd3_1 hold2791 (.A(\TRNG.hash[124] ),
    .X(net3919));
 sg13g2_dlygate4sd3_1 hold2792 (.A(\TRNG.sha256.expand.msg_schdl.RAM[14][3] ),
    .X(net3920));
 sg13g2_dlygate4sd3_1 hold2793 (.A(\TRNG.hash[239] ),
    .X(net3921));
 sg13g2_dlygate4sd3_1 hold2794 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][19] ),
    .X(net3922));
 sg13g2_dlygate4sd3_1 hold2795 (.A(_00220_),
    .X(net3923));
 sg13g2_dlygate4sd3_1 hold2796 (.A(_00237_),
    .X(net3924));
 sg13g2_dlygate4sd3_1 hold2797 (.A(\TRNG.sha256.expand.msg_schdl.RAM[2][29] ),
    .X(net3925));
 sg13g2_dlygate4sd3_1 hold2798 (.A(_05318_),
    .X(net3926));
 sg13g2_dlygate4sd3_1 hold2799 (.A(_00085_),
    .X(net3927));
 sg13g2_dlygate4sd3_1 hold2800 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][22] ),
    .X(net3928));
 sg13g2_dlygate4sd3_1 hold2801 (.A(_05237_),
    .X(net3929));
 sg13g2_dlygate4sd3_1 hold2802 (.A(_00078_),
    .X(net3930));
 sg13g2_dlygate4sd3_1 hold2803 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][10] ),
    .X(net3931));
 sg13g2_dlygate4sd3_1 hold2804 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][4] ),
    .X(net3932));
 sg13g2_dlygate4sd3_1 hold2805 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][16] ),
    .X(net3933));
 sg13g2_dlygate4sd3_1 hold2806 (.A(\TRNG.sha256.expand.data1_to_ram[31] ),
    .X(net3934));
 sg13g2_dlygate4sd3_1 hold2807 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][11] ),
    .X(net3935));
 sg13g2_dlygate4sd3_1 hold2808 (.A(\TRNG.sha256.expand.msg_schdl.RAM[7][2] ),
    .X(net3936));
 sg13g2_dlygate4sd3_1 hold2809 (.A(\TRNG.Repetition_Count_Test.prev_bit ),
    .X(net3937));
 sg13g2_dlygate4sd3_1 hold2810 (.A(\TRNG.sha256.expand.msg_schdl.RAM[10][31] ),
    .X(net3938));
 sg13g2_dlygate4sd3_1 hold2811 (.A(\TRNG.hash[53] ),
    .X(net3939));
 sg13g2_dlygate4sd3_1 hold2812 (.A(_00232_),
    .X(net3940));
 sg13g2_dlygate4sd3_1 hold2813 (.A(\TRNG.sha256.expand.msg_schdl.RAM[15][25] ),
    .X(net3941));
 sg13g2_antennanp ANTENNA_1 (.A(_00022_));
 sg13g2_antennanp ANTENNA_2 (.A(_00025_));
 sg13g2_antennanp ANTENNA_3 (.A(_02205_));
 sg13g2_antennanp ANTENNA_4 (.A(_02205_));
 sg13g2_antennanp ANTENNA_5 (.A(_02205_));
 sg13g2_antennanp ANTENNA_6 (.A(_02205_));
 sg13g2_antennanp ANTENNA_7 (.A(_04304_));
 sg13g2_antennanp ANTENNA_8 (.A(_04304_));
 sg13g2_antennanp ANTENNA_9 (.A(_04304_));
 sg13g2_antennanp ANTENNA_10 (.A(_04845_));
 sg13g2_antennanp ANTENNA_11 (.A(_04845_));
 sg13g2_antennanp ANTENNA_12 (.A(_04845_));
 sg13g2_antennanp ANTENNA_13 (.A(_08817_));
 sg13g2_antennanp ANTENNA_14 (.A(clk));
 sg13g2_antennanp ANTENNA_15 (.A(clk));
 sg13g2_antennanp ANTENNA_16 (.A(net5090));
 sg13g2_antennanp ANTENNA_17 (.A(net5090));
 sg13g2_antennanp ANTENNA_18 (.A(net5090));
 sg13g2_antennanp ANTENNA_19 (.A(net5090));
 sg13g2_antennanp ANTENNA_20 (.A(net5090));
 sg13g2_antennanp ANTENNA_21 (.A(net5090));
 sg13g2_antennanp ANTENNA_22 (.A(net5090));
 sg13g2_antennanp ANTENNA_23 (.A(net1));
 sg13g2_antennanp ANTENNA_24 (.A(net1));
 sg13g2_antennanp ANTENNA_25 (.A(net1));
 sg13g2_antennanp ANTENNA_26 (.A(\TRNG.Word_Valid ));
 sg13g2_antennanp ANTENNA_27 (.A(\TRNG.Word_Valid ));
 sg13g2_antennanp ANTENNA_28 (.A(\TRNG.Word_Valid ));
 sg13g2_antennanp ANTENNA_29 (.A(\TRNG.Word_Valid ));
 sg13g2_antennanp ANTENNA_30 (.A(\TRNG.Word_Valid ));
 sg13g2_antennanp ANTENNA_31 (.A(\TRNG.sha256.W[1] ));
 sg13g2_antennanp ANTENNA_32 (.A(\TRNG.sha256.W[1] ));
 sg13g2_antennanp ANTENNA_33 (.A(\TRNG.sha256.W[1] ));
 sg13g2_antennanp ANTENNA_34 (.A(\TRNG.sha256.expand.data1_to_ram[11] ));
 sg13g2_antennanp ANTENNA_35 (.A(\TRNG.sha256.expand.data1_to_ram[11] ));
 sg13g2_antennanp ANTENNA_36 (.A(\TRNG.sha256.expand.data1_to_ram[11] ));
 sg13g2_antennanp ANTENNA_37 (.A(_00002_));
 sg13g2_antennanp ANTENNA_38 (.A(_00022_));
 sg13g2_antennanp ANTENNA_39 (.A(_00030_));
 sg13g2_antennanp ANTENNA_40 (.A(_02205_));
 sg13g2_antennanp ANTENNA_41 (.A(_02205_));
 sg13g2_antennanp ANTENNA_42 (.A(_02205_));
 sg13g2_antennanp ANTENNA_43 (.A(_02205_));
 sg13g2_antennanp ANTENNA_44 (.A(_04845_));
 sg13g2_antennanp ANTENNA_45 (.A(_04845_));
 sg13g2_antennanp ANTENNA_46 (.A(_04845_));
 sg13g2_antennanp ANTENNA_47 (.A(_04845_));
 sg13g2_antennanp ANTENNA_48 (.A(_04845_));
 sg13g2_antennanp ANTENNA_49 (.A(_04845_));
 sg13g2_antennanp ANTENNA_50 (.A(_04845_));
 sg13g2_antennanp ANTENNA_51 (.A(_04845_));
 sg13g2_antennanp ANTENNA_52 (.A(_04845_));
 sg13g2_antennanp ANTENNA_53 (.A(_08817_));
 sg13g2_antennanp ANTENNA_54 (.A(clk));
 sg13g2_antennanp ANTENNA_55 (.A(clk));
 sg13g2_antennanp ANTENNA_56 (.A(net4914));
 sg13g2_antennanp ANTENNA_57 (.A(net4914));
 sg13g2_antennanp ANTENNA_58 (.A(net4914));
 sg13g2_antennanp ANTENNA_59 (.A(net4914));
 sg13g2_antennanp ANTENNA_60 (.A(net4914));
 sg13g2_antennanp ANTENNA_61 (.A(net4914));
 sg13g2_antennanp ANTENNA_62 (.A(net4914));
 sg13g2_antennanp ANTENNA_63 (.A(net4914));
 sg13g2_antennanp ANTENNA_64 (.A(\TRNG.sha256.W[1] ));
 sg13g2_antennanp ANTENNA_65 (.A(\TRNG.sha256.W[1] ));
 sg13g2_antennanp ANTENNA_66 (.A(\TRNG.sha256.W[1] ));
 sg13g2_antennanp ANTENNA_67 (.A(_00002_));
 sg13g2_antennanp ANTENNA_68 (.A(_00030_));
 sg13g2_antennanp ANTENNA_69 (.A(_02205_));
 sg13g2_antennanp ANTENNA_70 (.A(_02205_));
 sg13g2_antennanp ANTENNA_71 (.A(_04845_));
 sg13g2_antennanp ANTENNA_72 (.A(_04845_));
 sg13g2_antennanp ANTENNA_73 (.A(_04845_));
 sg13g2_antennanp ANTENNA_74 (.A(_08817_));
 sg13g2_antennanp ANTENNA_75 (.A(clk));
 sg13g2_antennanp ANTENNA_76 (.A(clk));
 sg13g2_antennanp ANTENNA_77 (.A(net4914));
 sg13g2_antennanp ANTENNA_78 (.A(net4914));
 sg13g2_antennanp ANTENNA_79 (.A(net4914));
 sg13g2_antennanp ANTENNA_80 (.A(net4914));
 sg13g2_antennanp ANTENNA_81 (.A(net4914));
 sg13g2_antennanp ANTENNA_82 (.A(net4914));
 sg13g2_antennanp ANTENNA_83 (.A(net4914));
 sg13g2_antennanp ANTENNA_84 (.A(net4914));
 sg13g2_antennanp ANTENNA_85 (.A(net4914));
 sg13g2_antennanp ANTENNA_86 (.A(net4914));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_decap_8 FILLER_0_896 ();
 sg13g2_decap_8 FILLER_0_903 ();
 sg13g2_decap_8 FILLER_0_910 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_decap_8 FILLER_0_924 ();
 sg13g2_decap_8 FILLER_0_931 ();
 sg13g2_decap_8 FILLER_0_938 ();
 sg13g2_decap_8 FILLER_0_945 ();
 sg13g2_decap_4 FILLER_0_952 ();
 sg13g2_fill_2 FILLER_0_956 ();
 sg13g2_fill_1 FILLER_0_1020 ();
 sg13g2_fill_1 FILLER_0_1078 ();
 sg13g2_fill_2 FILLER_0_1115 ();
 sg13g2_fill_1 FILLER_0_1122 ();
 sg13g2_fill_2 FILLER_0_1132 ();
 sg13g2_fill_1 FILLER_0_1268 ();
 sg13g2_fill_2 FILLER_0_1492 ();
 sg13g2_fill_1 FILLER_0_1558 ();
 sg13g2_decap_8 FILLER_0_1637 ();
 sg13g2_decap_8 FILLER_0_1644 ();
 sg13g2_decap_8 FILLER_0_1651 ();
 sg13g2_decap_8 FILLER_0_1658 ();
 sg13g2_decap_8 FILLER_0_1665 ();
 sg13g2_decap_4 FILLER_0_1672 ();
 sg13g2_fill_1 FILLER_0_1688 ();
 sg13g2_fill_2 FILLER_0_1732 ();
 sg13g2_fill_1 FILLER_0_1734 ();
 sg13g2_decap_4 FILLER_0_1798 ();
 sg13g2_fill_1 FILLER_0_1802 ();
 sg13g2_decap_4 FILLER_0_1813 ();
 sg13g2_fill_1 FILLER_0_1817 ();
 sg13g2_decap_8 FILLER_0_1831 ();
 sg13g2_decap_8 FILLER_0_1838 ();
 sg13g2_decap_8 FILLER_0_1845 ();
 sg13g2_decap_8 FILLER_0_1852 ();
 sg13g2_decap_8 FILLER_0_1859 ();
 sg13g2_decap_8 FILLER_0_1866 ();
 sg13g2_decap_8 FILLER_0_1873 ();
 sg13g2_decap_8 FILLER_0_1880 ();
 sg13g2_fill_2 FILLER_0_1887 ();
 sg13g2_fill_1 FILLER_0_1922 ();
 sg13g2_decap_8 FILLER_0_1971 ();
 sg13g2_decap_8 FILLER_0_1978 ();
 sg13g2_decap_8 FILLER_0_1985 ();
 sg13g2_decap_8 FILLER_0_1992 ();
 sg13g2_decap_8 FILLER_0_1999 ();
 sg13g2_decap_8 FILLER_0_2006 ();
 sg13g2_decap_8 FILLER_0_2013 ();
 sg13g2_decap_8 FILLER_0_2020 ();
 sg13g2_decap_8 FILLER_0_2027 ();
 sg13g2_decap_8 FILLER_0_2034 ();
 sg13g2_decap_8 FILLER_0_2064 ();
 sg13g2_decap_8 FILLER_0_2071 ();
 sg13g2_decap_8 FILLER_0_2078 ();
 sg13g2_decap_8 FILLER_0_2085 ();
 sg13g2_decap_8 FILLER_0_2092 ();
 sg13g2_decap_8 FILLER_0_2099 ();
 sg13g2_decap_8 FILLER_0_2106 ();
 sg13g2_decap_8 FILLER_0_2113 ();
 sg13g2_decap_8 FILLER_0_2120 ();
 sg13g2_decap_8 FILLER_0_2127 ();
 sg13g2_decap_8 FILLER_0_2134 ();
 sg13g2_decap_8 FILLER_0_2141 ();
 sg13g2_decap_8 FILLER_0_2148 ();
 sg13g2_decap_8 FILLER_0_2155 ();
 sg13g2_decap_8 FILLER_0_2162 ();
 sg13g2_decap_8 FILLER_0_2169 ();
 sg13g2_decap_8 FILLER_0_2176 ();
 sg13g2_decap_8 FILLER_0_2183 ();
 sg13g2_decap_8 FILLER_0_2190 ();
 sg13g2_decap_8 FILLER_0_2197 ();
 sg13g2_decap_8 FILLER_0_2204 ();
 sg13g2_decap_8 FILLER_0_2211 ();
 sg13g2_decap_8 FILLER_0_2218 ();
 sg13g2_decap_8 FILLER_0_2225 ();
 sg13g2_decap_8 FILLER_0_2232 ();
 sg13g2_decap_8 FILLER_0_2239 ();
 sg13g2_decap_8 FILLER_0_2246 ();
 sg13g2_decap_8 FILLER_0_2253 ();
 sg13g2_decap_8 FILLER_0_2260 ();
 sg13g2_decap_8 FILLER_0_2267 ();
 sg13g2_decap_8 FILLER_0_2274 ();
 sg13g2_decap_8 FILLER_0_2281 ();
 sg13g2_decap_8 FILLER_0_2288 ();
 sg13g2_decap_8 FILLER_0_2295 ();
 sg13g2_decap_8 FILLER_0_2302 ();
 sg13g2_decap_8 FILLER_0_2309 ();
 sg13g2_decap_8 FILLER_0_2316 ();
 sg13g2_decap_8 FILLER_0_2323 ();
 sg13g2_decap_8 FILLER_0_2330 ();
 sg13g2_decap_8 FILLER_0_2337 ();
 sg13g2_decap_8 FILLER_0_2344 ();
 sg13g2_decap_8 FILLER_0_2351 ();
 sg13g2_decap_8 FILLER_0_2358 ();
 sg13g2_decap_8 FILLER_0_2365 ();
 sg13g2_decap_8 FILLER_0_2372 ();
 sg13g2_decap_8 FILLER_0_2379 ();
 sg13g2_decap_8 FILLER_0_2386 ();
 sg13g2_decap_8 FILLER_0_2393 ();
 sg13g2_decap_8 FILLER_0_2400 ();
 sg13g2_decap_8 FILLER_0_2407 ();
 sg13g2_decap_8 FILLER_0_2414 ();
 sg13g2_decap_8 FILLER_0_2421 ();
 sg13g2_decap_8 FILLER_0_2428 ();
 sg13g2_decap_8 FILLER_0_2435 ();
 sg13g2_decap_8 FILLER_0_2442 ();
 sg13g2_decap_8 FILLER_0_2449 ();
 sg13g2_decap_8 FILLER_0_2456 ();
 sg13g2_decap_8 FILLER_0_2463 ();
 sg13g2_decap_8 FILLER_0_2470 ();
 sg13g2_decap_8 FILLER_0_2477 ();
 sg13g2_decap_8 FILLER_0_2484 ();
 sg13g2_decap_8 FILLER_0_2491 ();
 sg13g2_decap_8 FILLER_0_2498 ();
 sg13g2_decap_8 FILLER_0_2505 ();
 sg13g2_decap_8 FILLER_0_2512 ();
 sg13g2_decap_8 FILLER_0_2519 ();
 sg13g2_decap_8 FILLER_0_2526 ();
 sg13g2_decap_8 FILLER_0_2533 ();
 sg13g2_decap_8 FILLER_0_2540 ();
 sg13g2_decap_8 FILLER_0_2547 ();
 sg13g2_decap_8 FILLER_0_2554 ();
 sg13g2_decap_8 FILLER_0_2561 ();
 sg13g2_decap_8 FILLER_0_2568 ();
 sg13g2_decap_8 FILLER_0_2575 ();
 sg13g2_decap_8 FILLER_0_2582 ();
 sg13g2_decap_8 FILLER_0_2589 ();
 sg13g2_decap_8 FILLER_0_2596 ();
 sg13g2_decap_8 FILLER_0_2603 ();
 sg13g2_decap_8 FILLER_0_2610 ();
 sg13g2_decap_8 FILLER_0_2617 ();
 sg13g2_decap_8 FILLER_0_2624 ();
 sg13g2_decap_8 FILLER_0_2631 ();
 sg13g2_decap_8 FILLER_0_2638 ();
 sg13g2_decap_8 FILLER_0_2645 ();
 sg13g2_decap_8 FILLER_0_2652 ();
 sg13g2_decap_8 FILLER_0_2659 ();
 sg13g2_decap_8 FILLER_0_2666 ();
 sg13g2_fill_1 FILLER_0_2673 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_decap_8 FILLER_1_875 ();
 sg13g2_decap_8 FILLER_1_882 ();
 sg13g2_decap_8 FILLER_1_889 ();
 sg13g2_decap_8 FILLER_1_896 ();
 sg13g2_decap_8 FILLER_1_903 ();
 sg13g2_decap_8 FILLER_1_910 ();
 sg13g2_decap_8 FILLER_1_917 ();
 sg13g2_decap_8 FILLER_1_924 ();
 sg13g2_decap_8 FILLER_1_931 ();
 sg13g2_decap_8 FILLER_1_938 ();
 sg13g2_decap_8 FILLER_1_945 ();
 sg13g2_decap_8 FILLER_1_952 ();
 sg13g2_fill_2 FILLER_1_959 ();
 sg13g2_fill_1 FILLER_1_1236 ();
 sg13g2_fill_1 FILLER_1_1306 ();
 sg13g2_fill_2 FILLER_1_1520 ();
 sg13g2_decap_8 FILLER_1_1651 ();
 sg13g2_decap_8 FILLER_1_1658 ();
 sg13g2_decap_4 FILLER_1_1665 ();
 sg13g2_fill_2 FILLER_1_1783 ();
 sg13g2_fill_1 FILLER_1_1785 ();
 sg13g2_decap_8 FILLER_1_1847 ();
 sg13g2_decap_4 FILLER_1_1864 ();
 sg13g2_decap_8 FILLER_1_1881 ();
 sg13g2_fill_2 FILLER_1_1888 ();
 sg13g2_fill_2 FILLER_1_1946 ();
 sg13g2_decap_4 FILLER_1_1974 ();
 sg13g2_decap_4 FILLER_1_1987 ();
 sg13g2_fill_2 FILLER_1_1991 ();
 sg13g2_decap_8 FILLER_1_2010 ();
 sg13g2_decap_8 FILLER_1_2017 ();
 sg13g2_decap_8 FILLER_1_2024 ();
 sg13g2_decap_8 FILLER_1_2031 ();
 sg13g2_fill_1 FILLER_1_2038 ();
 sg13g2_decap_8 FILLER_1_2087 ();
 sg13g2_decap_8 FILLER_1_2094 ();
 sg13g2_decap_8 FILLER_1_2101 ();
 sg13g2_decap_4 FILLER_1_2108 ();
 sg13g2_fill_1 FILLER_1_2112 ();
 sg13g2_decap_8 FILLER_1_2117 ();
 sg13g2_decap_8 FILLER_1_2124 ();
 sg13g2_decap_8 FILLER_1_2131 ();
 sg13g2_decap_8 FILLER_1_2138 ();
 sg13g2_decap_8 FILLER_1_2145 ();
 sg13g2_decap_8 FILLER_1_2152 ();
 sg13g2_decap_8 FILLER_1_2159 ();
 sg13g2_decap_8 FILLER_1_2166 ();
 sg13g2_decap_8 FILLER_1_2173 ();
 sg13g2_decap_8 FILLER_1_2180 ();
 sg13g2_decap_8 FILLER_1_2187 ();
 sg13g2_decap_8 FILLER_1_2194 ();
 sg13g2_decap_8 FILLER_1_2201 ();
 sg13g2_decap_8 FILLER_1_2208 ();
 sg13g2_decap_8 FILLER_1_2215 ();
 sg13g2_decap_8 FILLER_1_2222 ();
 sg13g2_decap_8 FILLER_1_2229 ();
 sg13g2_decap_8 FILLER_1_2236 ();
 sg13g2_decap_8 FILLER_1_2243 ();
 sg13g2_decap_8 FILLER_1_2250 ();
 sg13g2_decap_8 FILLER_1_2257 ();
 sg13g2_decap_8 FILLER_1_2264 ();
 sg13g2_decap_8 FILLER_1_2271 ();
 sg13g2_decap_8 FILLER_1_2278 ();
 sg13g2_decap_8 FILLER_1_2285 ();
 sg13g2_decap_8 FILLER_1_2292 ();
 sg13g2_decap_8 FILLER_1_2299 ();
 sg13g2_decap_8 FILLER_1_2306 ();
 sg13g2_decap_8 FILLER_1_2313 ();
 sg13g2_decap_8 FILLER_1_2320 ();
 sg13g2_decap_8 FILLER_1_2327 ();
 sg13g2_decap_8 FILLER_1_2334 ();
 sg13g2_decap_8 FILLER_1_2341 ();
 sg13g2_decap_8 FILLER_1_2348 ();
 sg13g2_decap_8 FILLER_1_2355 ();
 sg13g2_decap_8 FILLER_1_2362 ();
 sg13g2_decap_8 FILLER_1_2369 ();
 sg13g2_decap_8 FILLER_1_2376 ();
 sg13g2_decap_8 FILLER_1_2383 ();
 sg13g2_decap_8 FILLER_1_2390 ();
 sg13g2_decap_8 FILLER_1_2397 ();
 sg13g2_decap_8 FILLER_1_2404 ();
 sg13g2_decap_8 FILLER_1_2411 ();
 sg13g2_decap_8 FILLER_1_2418 ();
 sg13g2_decap_8 FILLER_1_2425 ();
 sg13g2_decap_8 FILLER_1_2432 ();
 sg13g2_decap_8 FILLER_1_2439 ();
 sg13g2_decap_8 FILLER_1_2446 ();
 sg13g2_decap_8 FILLER_1_2453 ();
 sg13g2_decap_8 FILLER_1_2460 ();
 sg13g2_decap_8 FILLER_1_2467 ();
 sg13g2_decap_8 FILLER_1_2474 ();
 sg13g2_decap_8 FILLER_1_2481 ();
 sg13g2_decap_8 FILLER_1_2488 ();
 sg13g2_decap_8 FILLER_1_2495 ();
 sg13g2_decap_8 FILLER_1_2502 ();
 sg13g2_decap_8 FILLER_1_2509 ();
 sg13g2_decap_8 FILLER_1_2516 ();
 sg13g2_decap_8 FILLER_1_2523 ();
 sg13g2_decap_8 FILLER_1_2530 ();
 sg13g2_decap_8 FILLER_1_2537 ();
 sg13g2_decap_8 FILLER_1_2544 ();
 sg13g2_decap_8 FILLER_1_2551 ();
 sg13g2_decap_8 FILLER_1_2558 ();
 sg13g2_decap_8 FILLER_1_2565 ();
 sg13g2_decap_8 FILLER_1_2572 ();
 sg13g2_decap_8 FILLER_1_2579 ();
 sg13g2_decap_8 FILLER_1_2586 ();
 sg13g2_decap_8 FILLER_1_2593 ();
 sg13g2_decap_8 FILLER_1_2600 ();
 sg13g2_decap_8 FILLER_1_2607 ();
 sg13g2_decap_8 FILLER_1_2614 ();
 sg13g2_decap_8 FILLER_1_2621 ();
 sg13g2_decap_8 FILLER_1_2628 ();
 sg13g2_decap_8 FILLER_1_2635 ();
 sg13g2_decap_8 FILLER_1_2642 ();
 sg13g2_decap_8 FILLER_1_2649 ();
 sg13g2_decap_8 FILLER_1_2656 ();
 sg13g2_decap_8 FILLER_1_2663 ();
 sg13g2_decap_4 FILLER_1_2670 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_decap_8 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_2_868 ();
 sg13g2_decap_8 FILLER_2_875 ();
 sg13g2_decap_8 FILLER_2_882 ();
 sg13g2_decap_8 FILLER_2_889 ();
 sg13g2_decap_8 FILLER_2_896 ();
 sg13g2_decap_8 FILLER_2_903 ();
 sg13g2_decap_8 FILLER_2_910 ();
 sg13g2_decap_8 FILLER_2_917 ();
 sg13g2_decap_8 FILLER_2_924 ();
 sg13g2_decap_8 FILLER_2_931 ();
 sg13g2_decap_8 FILLER_2_938 ();
 sg13g2_decap_8 FILLER_2_945 ();
 sg13g2_fill_1 FILLER_2_957 ();
 sg13g2_fill_1 FILLER_2_1190 ();
 sg13g2_fill_2 FILLER_2_1321 ();
 sg13g2_fill_1 FILLER_2_1405 ();
 sg13g2_fill_2 FILLER_2_1521 ();
 sg13g2_fill_1 FILLER_2_1537 ();
 sg13g2_decap_4 FILLER_2_1653 ();
 sg13g2_fill_2 FILLER_2_1657 ();
 sg13g2_fill_2 FILLER_2_1707 ();
 sg13g2_fill_2 FILLER_2_1737 ();
 sg13g2_fill_1 FILLER_2_1739 ();
 sg13g2_fill_2 FILLER_2_1757 ();
 sg13g2_fill_2 FILLER_2_1795 ();
 sg13g2_decap_8 FILLER_2_1810 ();
 sg13g2_fill_1 FILLER_2_1817 ();
 sg13g2_decap_4 FILLER_2_1854 ();
 sg13g2_fill_2 FILLER_2_1858 ();
 sg13g2_decap_8 FILLER_2_1886 ();
 sg13g2_decap_8 FILLER_2_1893 ();
 sg13g2_fill_2 FILLER_2_1900 ();
 sg13g2_fill_1 FILLER_2_1902 ();
 sg13g2_fill_2 FILLER_2_1913 ();
 sg13g2_fill_1 FILLER_2_1915 ();
 sg13g2_fill_2 FILLER_2_2004 ();
 sg13g2_decap_4 FILLER_2_2021 ();
 sg13g2_fill_2 FILLER_2_2025 ();
 sg13g2_fill_2 FILLER_2_2040 ();
 sg13g2_decap_8 FILLER_2_2052 ();
 sg13g2_fill_1 FILLER_2_2059 ();
 sg13g2_fill_1 FILLER_2_2096 ();
 sg13g2_fill_2 FILLER_2_2123 ();
 sg13g2_fill_1 FILLER_2_2125 ();
 sg13g2_decap_8 FILLER_2_2152 ();
 sg13g2_decap_8 FILLER_2_2159 ();
 sg13g2_decap_8 FILLER_2_2166 ();
 sg13g2_decap_8 FILLER_2_2173 ();
 sg13g2_decap_8 FILLER_2_2180 ();
 sg13g2_decap_8 FILLER_2_2187 ();
 sg13g2_decap_8 FILLER_2_2194 ();
 sg13g2_decap_8 FILLER_2_2205 ();
 sg13g2_decap_8 FILLER_2_2212 ();
 sg13g2_decap_8 FILLER_2_2219 ();
 sg13g2_decap_8 FILLER_2_2226 ();
 sg13g2_decap_8 FILLER_2_2233 ();
 sg13g2_decap_8 FILLER_2_2240 ();
 sg13g2_decap_8 FILLER_2_2247 ();
 sg13g2_decap_8 FILLER_2_2254 ();
 sg13g2_decap_8 FILLER_2_2261 ();
 sg13g2_decap_8 FILLER_2_2268 ();
 sg13g2_decap_8 FILLER_2_2275 ();
 sg13g2_decap_8 FILLER_2_2282 ();
 sg13g2_decap_8 FILLER_2_2289 ();
 sg13g2_decap_8 FILLER_2_2296 ();
 sg13g2_decap_8 FILLER_2_2303 ();
 sg13g2_decap_8 FILLER_2_2310 ();
 sg13g2_decap_8 FILLER_2_2317 ();
 sg13g2_decap_8 FILLER_2_2324 ();
 sg13g2_decap_8 FILLER_2_2331 ();
 sg13g2_decap_8 FILLER_2_2338 ();
 sg13g2_decap_8 FILLER_2_2345 ();
 sg13g2_decap_8 FILLER_2_2352 ();
 sg13g2_decap_8 FILLER_2_2359 ();
 sg13g2_decap_8 FILLER_2_2366 ();
 sg13g2_decap_8 FILLER_2_2373 ();
 sg13g2_decap_8 FILLER_2_2380 ();
 sg13g2_decap_8 FILLER_2_2387 ();
 sg13g2_decap_8 FILLER_2_2394 ();
 sg13g2_decap_8 FILLER_2_2401 ();
 sg13g2_decap_8 FILLER_2_2408 ();
 sg13g2_decap_8 FILLER_2_2415 ();
 sg13g2_decap_8 FILLER_2_2422 ();
 sg13g2_decap_8 FILLER_2_2429 ();
 sg13g2_decap_8 FILLER_2_2436 ();
 sg13g2_decap_8 FILLER_2_2443 ();
 sg13g2_decap_8 FILLER_2_2450 ();
 sg13g2_decap_8 FILLER_2_2457 ();
 sg13g2_decap_8 FILLER_2_2464 ();
 sg13g2_decap_8 FILLER_2_2471 ();
 sg13g2_decap_8 FILLER_2_2478 ();
 sg13g2_decap_8 FILLER_2_2485 ();
 sg13g2_decap_8 FILLER_2_2492 ();
 sg13g2_decap_8 FILLER_2_2499 ();
 sg13g2_decap_8 FILLER_2_2506 ();
 sg13g2_decap_8 FILLER_2_2513 ();
 sg13g2_decap_8 FILLER_2_2520 ();
 sg13g2_decap_8 FILLER_2_2527 ();
 sg13g2_decap_8 FILLER_2_2534 ();
 sg13g2_decap_8 FILLER_2_2541 ();
 sg13g2_decap_8 FILLER_2_2548 ();
 sg13g2_decap_8 FILLER_2_2555 ();
 sg13g2_decap_8 FILLER_2_2562 ();
 sg13g2_decap_8 FILLER_2_2569 ();
 sg13g2_decap_8 FILLER_2_2576 ();
 sg13g2_decap_8 FILLER_2_2583 ();
 sg13g2_decap_8 FILLER_2_2590 ();
 sg13g2_decap_8 FILLER_2_2597 ();
 sg13g2_decap_8 FILLER_2_2604 ();
 sg13g2_decap_8 FILLER_2_2611 ();
 sg13g2_decap_8 FILLER_2_2618 ();
 sg13g2_decap_8 FILLER_2_2625 ();
 sg13g2_decap_8 FILLER_2_2632 ();
 sg13g2_decap_8 FILLER_2_2639 ();
 sg13g2_decap_8 FILLER_2_2646 ();
 sg13g2_decap_8 FILLER_2_2653 ();
 sg13g2_decap_8 FILLER_2_2660 ();
 sg13g2_decap_8 FILLER_2_2667 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_decap_8 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_3_868 ();
 sg13g2_decap_8 FILLER_3_875 ();
 sg13g2_decap_8 FILLER_3_882 ();
 sg13g2_decap_8 FILLER_3_889 ();
 sg13g2_decap_8 FILLER_3_896 ();
 sg13g2_decap_8 FILLER_3_903 ();
 sg13g2_decap_8 FILLER_3_910 ();
 sg13g2_decap_8 FILLER_3_917 ();
 sg13g2_decap_8 FILLER_3_924 ();
 sg13g2_decap_8 FILLER_3_931 ();
 sg13g2_fill_1 FILLER_3_938 ();
 sg13g2_fill_1 FILLER_3_964 ();
 sg13g2_fill_1 FILLER_3_983 ();
 sg13g2_fill_2 FILLER_3_994 ();
 sg13g2_fill_2 FILLER_3_1061 ();
 sg13g2_fill_1 FILLER_3_1119 ();
 sg13g2_fill_1 FILLER_3_1207 ();
 sg13g2_fill_2 FILLER_3_1291 ();
 sg13g2_fill_1 FILLER_3_1333 ();
 sg13g2_fill_2 FILLER_3_1586 ();
 sg13g2_fill_2 FILLER_3_1779 ();
 sg13g2_fill_2 FILLER_3_1791 ();
 sg13g2_fill_1 FILLER_3_1793 ();
 sg13g2_fill_2 FILLER_3_1807 ();
 sg13g2_fill_1 FILLER_3_1809 ();
 sg13g2_fill_2 FILLER_3_1836 ();
 sg13g2_fill_1 FILLER_3_1838 ();
 sg13g2_decap_8 FILLER_3_1843 ();
 sg13g2_fill_2 FILLER_3_1850 ();
 sg13g2_decap_8 FILLER_3_1862 ();
 sg13g2_fill_1 FILLER_3_1869 ();
 sg13g2_fill_1 FILLER_3_1906 ();
 sg13g2_fill_2 FILLER_3_1938 ();
 sg13g2_fill_2 FILLER_3_1975 ();
 sg13g2_fill_1 FILLER_3_1977 ();
 sg13g2_fill_1 FILLER_3_2047 ();
 sg13g2_decap_4 FILLER_3_2088 ();
 sg13g2_fill_2 FILLER_3_2092 ();
 sg13g2_fill_2 FILLER_3_2104 ();
 sg13g2_fill_1 FILLER_3_2131 ();
 sg13g2_decap_8 FILLER_3_2159 ();
 sg13g2_decap_8 FILLER_3_2166 ();
 sg13g2_decap_8 FILLER_3_2173 ();
 sg13g2_decap_8 FILLER_3_2229 ();
 sg13g2_decap_8 FILLER_3_2236 ();
 sg13g2_decap_8 FILLER_3_2243 ();
 sg13g2_decap_8 FILLER_3_2250 ();
 sg13g2_decap_8 FILLER_3_2257 ();
 sg13g2_decap_8 FILLER_3_2264 ();
 sg13g2_decap_8 FILLER_3_2271 ();
 sg13g2_decap_8 FILLER_3_2278 ();
 sg13g2_decap_8 FILLER_3_2285 ();
 sg13g2_decap_8 FILLER_3_2292 ();
 sg13g2_decap_8 FILLER_3_2299 ();
 sg13g2_decap_8 FILLER_3_2306 ();
 sg13g2_decap_8 FILLER_3_2313 ();
 sg13g2_decap_8 FILLER_3_2320 ();
 sg13g2_decap_8 FILLER_3_2327 ();
 sg13g2_decap_8 FILLER_3_2334 ();
 sg13g2_decap_8 FILLER_3_2341 ();
 sg13g2_decap_8 FILLER_3_2348 ();
 sg13g2_decap_8 FILLER_3_2355 ();
 sg13g2_decap_8 FILLER_3_2362 ();
 sg13g2_decap_8 FILLER_3_2369 ();
 sg13g2_decap_8 FILLER_3_2376 ();
 sg13g2_decap_8 FILLER_3_2383 ();
 sg13g2_decap_8 FILLER_3_2390 ();
 sg13g2_decap_8 FILLER_3_2397 ();
 sg13g2_decap_8 FILLER_3_2404 ();
 sg13g2_decap_8 FILLER_3_2411 ();
 sg13g2_decap_8 FILLER_3_2418 ();
 sg13g2_decap_8 FILLER_3_2425 ();
 sg13g2_decap_8 FILLER_3_2432 ();
 sg13g2_decap_8 FILLER_3_2439 ();
 sg13g2_decap_8 FILLER_3_2446 ();
 sg13g2_decap_8 FILLER_3_2453 ();
 sg13g2_decap_8 FILLER_3_2460 ();
 sg13g2_decap_8 FILLER_3_2467 ();
 sg13g2_decap_8 FILLER_3_2474 ();
 sg13g2_decap_8 FILLER_3_2481 ();
 sg13g2_decap_8 FILLER_3_2488 ();
 sg13g2_decap_8 FILLER_3_2495 ();
 sg13g2_decap_8 FILLER_3_2502 ();
 sg13g2_decap_8 FILLER_3_2509 ();
 sg13g2_decap_8 FILLER_3_2516 ();
 sg13g2_decap_8 FILLER_3_2523 ();
 sg13g2_decap_8 FILLER_3_2530 ();
 sg13g2_decap_8 FILLER_3_2537 ();
 sg13g2_decap_8 FILLER_3_2544 ();
 sg13g2_decap_8 FILLER_3_2551 ();
 sg13g2_decap_8 FILLER_3_2558 ();
 sg13g2_decap_8 FILLER_3_2565 ();
 sg13g2_decap_8 FILLER_3_2572 ();
 sg13g2_decap_8 FILLER_3_2579 ();
 sg13g2_decap_8 FILLER_3_2586 ();
 sg13g2_decap_8 FILLER_3_2593 ();
 sg13g2_decap_8 FILLER_3_2600 ();
 sg13g2_decap_8 FILLER_3_2607 ();
 sg13g2_decap_8 FILLER_3_2614 ();
 sg13g2_decap_8 FILLER_3_2621 ();
 sg13g2_decap_8 FILLER_3_2628 ();
 sg13g2_decap_8 FILLER_3_2635 ();
 sg13g2_decap_8 FILLER_3_2642 ();
 sg13g2_decap_8 FILLER_3_2649 ();
 sg13g2_decap_8 FILLER_3_2656 ();
 sg13g2_decap_8 FILLER_3_2663 ();
 sg13g2_decap_4 FILLER_3_2670 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_decap_8 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_4_868 ();
 sg13g2_decap_8 FILLER_4_875 ();
 sg13g2_decap_8 FILLER_4_882 ();
 sg13g2_decap_8 FILLER_4_889 ();
 sg13g2_decap_8 FILLER_4_896 ();
 sg13g2_decap_8 FILLER_4_903 ();
 sg13g2_decap_8 FILLER_4_910 ();
 sg13g2_decap_8 FILLER_4_917 ();
 sg13g2_decap_8 FILLER_4_924 ();
 sg13g2_fill_1 FILLER_4_946 ();
 sg13g2_fill_1 FILLER_4_952 ();
 sg13g2_fill_2 FILLER_4_992 ();
 sg13g2_fill_2 FILLER_4_1004 ();
 sg13g2_fill_2 FILLER_4_1089 ();
 sg13g2_fill_1 FILLER_4_1267 ();
 sg13g2_fill_1 FILLER_4_1369 ();
 sg13g2_fill_1 FILLER_4_1440 ();
 sg13g2_fill_1 FILLER_4_1538 ();
 sg13g2_fill_1 FILLER_4_1605 ();
 sg13g2_fill_1 FILLER_4_1650 ();
 sg13g2_fill_2 FILLER_4_1738 ();
 sg13g2_fill_2 FILLER_4_1822 ();
 sg13g2_fill_2 FILLER_4_1855 ();
 sg13g2_fill_2 FILLER_4_1892 ();
 sg13g2_fill_2 FILLER_4_1930 ();
 sg13g2_fill_1 FILLER_4_1932 ();
 sg13g2_fill_2 FILLER_4_1956 ();
 sg13g2_decap_8 FILLER_4_1994 ();
 sg13g2_fill_2 FILLER_4_2001 ();
 sg13g2_fill_1 FILLER_4_2003 ();
 sg13g2_fill_2 FILLER_4_2040 ();
 sg13g2_fill_1 FILLER_4_2072 ();
 sg13g2_fill_2 FILLER_4_2108 ();
 sg13g2_fill_1 FILLER_4_2110 ();
 sg13g2_fill_1 FILLER_4_2120 ();
 sg13g2_fill_2 FILLER_4_2157 ();
 sg13g2_fill_1 FILLER_4_2185 ();
 sg13g2_fill_1 FILLER_4_2257 ();
 sg13g2_decap_8 FILLER_4_2262 ();
 sg13g2_decap_8 FILLER_4_2269 ();
 sg13g2_decap_8 FILLER_4_2276 ();
 sg13g2_decap_8 FILLER_4_2283 ();
 sg13g2_decap_8 FILLER_4_2290 ();
 sg13g2_decap_8 FILLER_4_2297 ();
 sg13g2_decap_8 FILLER_4_2304 ();
 sg13g2_decap_8 FILLER_4_2311 ();
 sg13g2_decap_8 FILLER_4_2318 ();
 sg13g2_decap_8 FILLER_4_2325 ();
 sg13g2_decap_8 FILLER_4_2332 ();
 sg13g2_decap_8 FILLER_4_2339 ();
 sg13g2_decap_8 FILLER_4_2346 ();
 sg13g2_decap_8 FILLER_4_2353 ();
 sg13g2_decap_8 FILLER_4_2360 ();
 sg13g2_decap_8 FILLER_4_2367 ();
 sg13g2_decap_8 FILLER_4_2374 ();
 sg13g2_decap_8 FILLER_4_2381 ();
 sg13g2_decap_8 FILLER_4_2388 ();
 sg13g2_decap_8 FILLER_4_2395 ();
 sg13g2_decap_8 FILLER_4_2402 ();
 sg13g2_decap_8 FILLER_4_2409 ();
 sg13g2_decap_8 FILLER_4_2416 ();
 sg13g2_decap_8 FILLER_4_2423 ();
 sg13g2_decap_8 FILLER_4_2430 ();
 sg13g2_decap_8 FILLER_4_2437 ();
 sg13g2_decap_8 FILLER_4_2444 ();
 sg13g2_decap_8 FILLER_4_2451 ();
 sg13g2_decap_8 FILLER_4_2458 ();
 sg13g2_decap_8 FILLER_4_2465 ();
 sg13g2_decap_8 FILLER_4_2472 ();
 sg13g2_decap_8 FILLER_4_2479 ();
 sg13g2_decap_8 FILLER_4_2486 ();
 sg13g2_decap_8 FILLER_4_2493 ();
 sg13g2_decap_8 FILLER_4_2500 ();
 sg13g2_decap_8 FILLER_4_2507 ();
 sg13g2_decap_8 FILLER_4_2514 ();
 sg13g2_decap_8 FILLER_4_2521 ();
 sg13g2_decap_8 FILLER_4_2528 ();
 sg13g2_decap_8 FILLER_4_2535 ();
 sg13g2_decap_8 FILLER_4_2542 ();
 sg13g2_decap_8 FILLER_4_2549 ();
 sg13g2_decap_8 FILLER_4_2556 ();
 sg13g2_decap_8 FILLER_4_2563 ();
 sg13g2_decap_8 FILLER_4_2570 ();
 sg13g2_decap_8 FILLER_4_2577 ();
 sg13g2_decap_8 FILLER_4_2584 ();
 sg13g2_decap_8 FILLER_4_2591 ();
 sg13g2_decap_8 FILLER_4_2598 ();
 sg13g2_decap_8 FILLER_4_2605 ();
 sg13g2_decap_8 FILLER_4_2612 ();
 sg13g2_decap_8 FILLER_4_2619 ();
 sg13g2_decap_8 FILLER_4_2626 ();
 sg13g2_decap_8 FILLER_4_2633 ();
 sg13g2_decap_8 FILLER_4_2640 ();
 sg13g2_decap_8 FILLER_4_2647 ();
 sg13g2_decap_8 FILLER_4_2654 ();
 sg13g2_decap_8 FILLER_4_2661 ();
 sg13g2_decap_4 FILLER_4_2668 ();
 sg13g2_fill_2 FILLER_4_2672 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_326 ();
 sg13g2_decap_8 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_340 ();
 sg13g2_decap_8 FILLER_5_373 ();
 sg13g2_decap_8 FILLER_5_380 ();
 sg13g2_decap_8 FILLER_5_387 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_decap_8 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_5_415 ();
 sg13g2_decap_8 FILLER_5_422 ();
 sg13g2_decap_8 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_5_436 ();
 sg13g2_decap_8 FILLER_5_443 ();
 sg13g2_decap_8 FILLER_5_450 ();
 sg13g2_decap_8 FILLER_5_457 ();
 sg13g2_decap_8 FILLER_5_464 ();
 sg13g2_decap_8 FILLER_5_471 ();
 sg13g2_decap_8 FILLER_5_478 ();
 sg13g2_decap_8 FILLER_5_485 ();
 sg13g2_decap_8 FILLER_5_492 ();
 sg13g2_decap_8 FILLER_5_499 ();
 sg13g2_decap_8 FILLER_5_506 ();
 sg13g2_decap_8 FILLER_5_513 ();
 sg13g2_decap_8 FILLER_5_520 ();
 sg13g2_decap_8 FILLER_5_527 ();
 sg13g2_decap_8 FILLER_5_534 ();
 sg13g2_decap_8 FILLER_5_541 ();
 sg13g2_decap_8 FILLER_5_548 ();
 sg13g2_decap_8 FILLER_5_555 ();
 sg13g2_decap_8 FILLER_5_562 ();
 sg13g2_decap_8 FILLER_5_569 ();
 sg13g2_decap_8 FILLER_5_576 ();
 sg13g2_decap_8 FILLER_5_583 ();
 sg13g2_decap_8 FILLER_5_590 ();
 sg13g2_decap_8 FILLER_5_597 ();
 sg13g2_decap_8 FILLER_5_604 ();
 sg13g2_decap_8 FILLER_5_611 ();
 sg13g2_decap_8 FILLER_5_618 ();
 sg13g2_decap_8 FILLER_5_625 ();
 sg13g2_decap_8 FILLER_5_632 ();
 sg13g2_decap_8 FILLER_5_639 ();
 sg13g2_decap_8 FILLER_5_646 ();
 sg13g2_decap_8 FILLER_5_653 ();
 sg13g2_decap_4 FILLER_5_660 ();
 sg13g2_fill_1 FILLER_5_668 ();
 sg13g2_decap_8 FILLER_5_681 ();
 sg13g2_decap_8 FILLER_5_688 ();
 sg13g2_decap_8 FILLER_5_695 ();
 sg13g2_decap_8 FILLER_5_702 ();
 sg13g2_decap_8 FILLER_5_709 ();
 sg13g2_decap_8 FILLER_5_716 ();
 sg13g2_decap_8 FILLER_5_723 ();
 sg13g2_decap_8 FILLER_5_730 ();
 sg13g2_decap_8 FILLER_5_737 ();
 sg13g2_decap_8 FILLER_5_744 ();
 sg13g2_decap_8 FILLER_5_751 ();
 sg13g2_decap_8 FILLER_5_758 ();
 sg13g2_decap_8 FILLER_5_765 ();
 sg13g2_decap_8 FILLER_5_772 ();
 sg13g2_decap_8 FILLER_5_779 ();
 sg13g2_decap_8 FILLER_5_786 ();
 sg13g2_decap_8 FILLER_5_793 ();
 sg13g2_decap_8 FILLER_5_800 ();
 sg13g2_decap_8 FILLER_5_807 ();
 sg13g2_decap_8 FILLER_5_814 ();
 sg13g2_decap_8 FILLER_5_821 ();
 sg13g2_decap_8 FILLER_5_828 ();
 sg13g2_decap_8 FILLER_5_835 ();
 sg13g2_decap_8 FILLER_5_842 ();
 sg13g2_decap_8 FILLER_5_849 ();
 sg13g2_decap_8 FILLER_5_856 ();
 sg13g2_decap_8 FILLER_5_863 ();
 sg13g2_decap_8 FILLER_5_870 ();
 sg13g2_decap_8 FILLER_5_877 ();
 sg13g2_decap_8 FILLER_5_884 ();
 sg13g2_decap_8 FILLER_5_891 ();
 sg13g2_decap_8 FILLER_5_898 ();
 sg13g2_decap_8 FILLER_5_905 ();
 sg13g2_fill_2 FILLER_5_912 ();
 sg13g2_fill_1 FILLER_5_914 ();
 sg13g2_fill_1 FILLER_5_960 ();
 sg13g2_fill_1 FILLER_5_1010 ();
 sg13g2_fill_2 FILLER_5_1064 ();
 sg13g2_fill_2 FILLER_5_1075 ();
 sg13g2_fill_1 FILLER_5_1118 ();
 sg13g2_fill_2 FILLER_5_1257 ();
 sg13g2_fill_1 FILLER_5_1401 ();
 sg13g2_fill_1 FILLER_5_1442 ();
 sg13g2_fill_1 FILLER_5_1471 ();
 sg13g2_fill_2 FILLER_5_1593 ();
 sg13g2_fill_1 FILLER_5_1609 ();
 sg13g2_fill_1 FILLER_5_1659 ();
 sg13g2_fill_2 FILLER_5_1775 ();
 sg13g2_fill_1 FILLER_5_1777 ();
 sg13g2_fill_1 FILLER_5_1787 ();
 sg13g2_fill_2 FILLER_5_1818 ();
 sg13g2_fill_2 FILLER_5_1859 ();
 sg13g2_fill_2 FILLER_5_1875 ();
 sg13g2_fill_1 FILLER_5_1877 ();
 sg13g2_fill_2 FILLER_5_1887 ();
 sg13g2_fill_1 FILLER_5_1889 ();
 sg13g2_decap_8 FILLER_5_1903 ();
 sg13g2_fill_1 FILLER_5_1927 ();
 sg13g2_decap_4 FILLER_5_1968 ();
 sg13g2_fill_1 FILLER_5_1972 ();
 sg13g2_fill_1 FILLER_5_2017 ();
 sg13g2_fill_2 FILLER_5_2054 ();
 sg13g2_fill_1 FILLER_5_2056 ();
 sg13g2_fill_2 FILLER_5_2129 ();
 sg13g2_fill_2 FILLER_5_2167 ();
 sg13g2_fill_1 FILLER_5_2169 ();
 sg13g2_decap_4 FILLER_5_2196 ();
 sg13g2_fill_1 FILLER_5_2200 ();
 sg13g2_fill_2 FILLER_5_2227 ();
 sg13g2_fill_2 FILLER_5_2262 ();
 sg13g2_decap_4 FILLER_5_2274 ();
 sg13g2_fill_1 FILLER_5_2278 ();
 sg13g2_decap_8 FILLER_5_2292 ();
 sg13g2_decap_8 FILLER_5_2299 ();
 sg13g2_decap_8 FILLER_5_2306 ();
 sg13g2_decap_8 FILLER_5_2313 ();
 sg13g2_decap_8 FILLER_5_2320 ();
 sg13g2_decap_8 FILLER_5_2327 ();
 sg13g2_decap_8 FILLER_5_2334 ();
 sg13g2_decap_8 FILLER_5_2341 ();
 sg13g2_decap_8 FILLER_5_2348 ();
 sg13g2_decap_8 FILLER_5_2355 ();
 sg13g2_decap_8 FILLER_5_2362 ();
 sg13g2_decap_8 FILLER_5_2369 ();
 sg13g2_decap_8 FILLER_5_2376 ();
 sg13g2_decap_8 FILLER_5_2383 ();
 sg13g2_decap_8 FILLER_5_2390 ();
 sg13g2_decap_8 FILLER_5_2397 ();
 sg13g2_decap_8 FILLER_5_2404 ();
 sg13g2_decap_8 FILLER_5_2411 ();
 sg13g2_decap_8 FILLER_5_2418 ();
 sg13g2_decap_8 FILLER_5_2425 ();
 sg13g2_decap_8 FILLER_5_2432 ();
 sg13g2_decap_8 FILLER_5_2439 ();
 sg13g2_decap_8 FILLER_5_2446 ();
 sg13g2_decap_8 FILLER_5_2453 ();
 sg13g2_decap_8 FILLER_5_2460 ();
 sg13g2_decap_8 FILLER_5_2467 ();
 sg13g2_decap_8 FILLER_5_2474 ();
 sg13g2_decap_8 FILLER_5_2481 ();
 sg13g2_decap_8 FILLER_5_2488 ();
 sg13g2_decap_8 FILLER_5_2495 ();
 sg13g2_decap_8 FILLER_5_2502 ();
 sg13g2_decap_8 FILLER_5_2509 ();
 sg13g2_decap_8 FILLER_5_2516 ();
 sg13g2_decap_8 FILLER_5_2523 ();
 sg13g2_decap_8 FILLER_5_2530 ();
 sg13g2_decap_8 FILLER_5_2537 ();
 sg13g2_decap_8 FILLER_5_2544 ();
 sg13g2_decap_8 FILLER_5_2551 ();
 sg13g2_decap_8 FILLER_5_2558 ();
 sg13g2_decap_8 FILLER_5_2565 ();
 sg13g2_decap_8 FILLER_5_2572 ();
 sg13g2_decap_8 FILLER_5_2579 ();
 sg13g2_decap_8 FILLER_5_2586 ();
 sg13g2_decap_8 FILLER_5_2593 ();
 sg13g2_decap_8 FILLER_5_2600 ();
 sg13g2_decap_8 FILLER_5_2607 ();
 sg13g2_decap_8 FILLER_5_2614 ();
 sg13g2_decap_8 FILLER_5_2621 ();
 sg13g2_decap_8 FILLER_5_2628 ();
 sg13g2_decap_8 FILLER_5_2635 ();
 sg13g2_decap_8 FILLER_5_2642 ();
 sg13g2_decap_8 FILLER_5_2649 ();
 sg13g2_decap_8 FILLER_5_2656 ();
 sg13g2_decap_8 FILLER_5_2663 ();
 sg13g2_decap_4 FILLER_5_2670 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_4 FILLER_6_273 ();
 sg13g2_fill_2 FILLER_6_277 ();
 sg13g2_fill_2 FILLER_6_288 ();
 sg13g2_decap_8 FILLER_6_304 ();
 sg13g2_decap_4 FILLER_6_337 ();
 sg13g2_decap_8 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_372 ();
 sg13g2_decap_8 FILLER_6_379 ();
 sg13g2_decap_8 FILLER_6_386 ();
 sg13g2_decap_8 FILLER_6_393 ();
 sg13g2_fill_2 FILLER_6_400 ();
 sg13g2_fill_1 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_fill_1 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_fill_1 FILLER_6_602 ();
 sg13g2_decap_4 FILLER_6_616 ();
 sg13g2_fill_2 FILLER_6_632 ();
 sg13g2_fill_2 FILLER_6_638 ();
 sg13g2_decap_4 FILLER_6_688 ();
 sg13g2_fill_1 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_712 ();
 sg13g2_decap_8 FILLER_6_719 ();
 sg13g2_decap_8 FILLER_6_726 ();
 sg13g2_decap_8 FILLER_6_733 ();
 sg13g2_decap_8 FILLER_6_740 ();
 sg13g2_decap_8 FILLER_6_747 ();
 sg13g2_decap_8 FILLER_6_754 ();
 sg13g2_decap_8 FILLER_6_761 ();
 sg13g2_decap_8 FILLER_6_768 ();
 sg13g2_decap_8 FILLER_6_775 ();
 sg13g2_decap_8 FILLER_6_782 ();
 sg13g2_decap_8 FILLER_6_789 ();
 sg13g2_decap_8 FILLER_6_796 ();
 sg13g2_decap_8 FILLER_6_803 ();
 sg13g2_decap_8 FILLER_6_810 ();
 sg13g2_decap_8 FILLER_6_817 ();
 sg13g2_decap_8 FILLER_6_824 ();
 sg13g2_decap_8 FILLER_6_831 ();
 sg13g2_decap_8 FILLER_6_838 ();
 sg13g2_decap_8 FILLER_6_845 ();
 sg13g2_decap_8 FILLER_6_852 ();
 sg13g2_decap_8 FILLER_6_859 ();
 sg13g2_decap_8 FILLER_6_866 ();
 sg13g2_decap_8 FILLER_6_873 ();
 sg13g2_decap_8 FILLER_6_880 ();
 sg13g2_decap_8 FILLER_6_887 ();
 sg13g2_decap_8 FILLER_6_894 ();
 sg13g2_decap_8 FILLER_6_901 ();
 sg13g2_decap_8 FILLER_6_908 ();
 sg13g2_decap_4 FILLER_6_915 ();
 sg13g2_fill_2 FILLER_6_955 ();
 sg13g2_fill_2 FILLER_6_983 ();
 sg13g2_fill_2 FILLER_6_1157 ();
 sg13g2_fill_1 FILLER_6_1206 ();
 sg13g2_fill_1 FILLER_6_1266 ();
 sg13g2_fill_2 FILLER_6_1285 ();
 sg13g2_fill_2 FILLER_6_1296 ();
 sg13g2_fill_1 FILLER_6_1331 ();
 sg13g2_fill_2 FILLER_6_1389 ();
 sg13g2_fill_1 FILLER_6_1503 ();
 sg13g2_fill_2 FILLER_6_1530 ();
 sg13g2_fill_1 FILLER_6_1578 ();
 sg13g2_fill_2 FILLER_6_1642 ();
 sg13g2_fill_2 FILLER_6_1685 ();
 sg13g2_fill_1 FILLER_6_1706 ();
 sg13g2_fill_1 FILLER_6_1718 ();
 sg13g2_fill_2 FILLER_6_1729 ();
 sg13g2_fill_1 FILLER_6_1731 ();
 sg13g2_fill_1 FILLER_6_1743 ();
 sg13g2_fill_2 FILLER_6_1750 ();
 sg13g2_fill_1 FILLER_6_1752 ();
 sg13g2_fill_1 FILLER_6_1819 ();
 sg13g2_fill_1 FILLER_6_1922 ();
 sg13g2_fill_2 FILLER_6_1933 ();
 sg13g2_fill_1 FILLER_6_1935 ();
 sg13g2_fill_2 FILLER_6_1953 ();
 sg13g2_fill_1 FILLER_6_1955 ();
 sg13g2_fill_1 FILLER_6_1992 ();
 sg13g2_decap_4 FILLER_6_2006 ();
 sg13g2_fill_1 FILLER_6_2010 ();
 sg13g2_decap_4 FILLER_6_2021 ();
 sg13g2_decap_4 FILLER_6_2034 ();
 sg13g2_fill_1 FILLER_6_2038 ();
 sg13g2_decap_4 FILLER_6_2101 ();
 sg13g2_fill_2 FILLER_6_2118 ();
 sg13g2_fill_1 FILLER_6_2120 ();
 sg13g2_fill_1 FILLER_6_2158 ();
 sg13g2_decap_4 FILLER_6_2205 ();
 sg13g2_decap_8 FILLER_6_2222 ();
 sg13g2_fill_1 FILLER_6_2229 ();
 sg13g2_fill_2 FILLER_6_2244 ();
 sg13g2_fill_1 FILLER_6_2246 ();
 sg13g2_decap_8 FILLER_6_2299 ();
 sg13g2_decap_8 FILLER_6_2306 ();
 sg13g2_decap_8 FILLER_6_2313 ();
 sg13g2_decap_8 FILLER_6_2320 ();
 sg13g2_decap_8 FILLER_6_2327 ();
 sg13g2_decap_8 FILLER_6_2334 ();
 sg13g2_decap_8 FILLER_6_2341 ();
 sg13g2_decap_8 FILLER_6_2348 ();
 sg13g2_decap_8 FILLER_6_2355 ();
 sg13g2_decap_8 FILLER_6_2362 ();
 sg13g2_decap_8 FILLER_6_2369 ();
 sg13g2_decap_8 FILLER_6_2376 ();
 sg13g2_decap_8 FILLER_6_2383 ();
 sg13g2_decap_8 FILLER_6_2390 ();
 sg13g2_decap_8 FILLER_6_2397 ();
 sg13g2_decap_8 FILLER_6_2404 ();
 sg13g2_decap_8 FILLER_6_2411 ();
 sg13g2_decap_8 FILLER_6_2418 ();
 sg13g2_decap_8 FILLER_6_2425 ();
 sg13g2_decap_8 FILLER_6_2432 ();
 sg13g2_decap_8 FILLER_6_2439 ();
 sg13g2_decap_8 FILLER_6_2446 ();
 sg13g2_decap_8 FILLER_6_2453 ();
 sg13g2_decap_8 FILLER_6_2460 ();
 sg13g2_decap_8 FILLER_6_2467 ();
 sg13g2_decap_8 FILLER_6_2474 ();
 sg13g2_decap_8 FILLER_6_2481 ();
 sg13g2_decap_8 FILLER_6_2488 ();
 sg13g2_decap_8 FILLER_6_2495 ();
 sg13g2_decap_8 FILLER_6_2502 ();
 sg13g2_decap_8 FILLER_6_2509 ();
 sg13g2_decap_8 FILLER_6_2516 ();
 sg13g2_decap_8 FILLER_6_2523 ();
 sg13g2_decap_8 FILLER_6_2530 ();
 sg13g2_decap_8 FILLER_6_2537 ();
 sg13g2_decap_8 FILLER_6_2544 ();
 sg13g2_decap_8 FILLER_6_2551 ();
 sg13g2_decap_8 FILLER_6_2558 ();
 sg13g2_decap_8 FILLER_6_2565 ();
 sg13g2_decap_8 FILLER_6_2572 ();
 sg13g2_decap_8 FILLER_6_2579 ();
 sg13g2_decap_8 FILLER_6_2586 ();
 sg13g2_decap_8 FILLER_6_2593 ();
 sg13g2_decap_8 FILLER_6_2600 ();
 sg13g2_decap_8 FILLER_6_2607 ();
 sg13g2_decap_8 FILLER_6_2614 ();
 sg13g2_decap_8 FILLER_6_2621 ();
 sg13g2_decap_8 FILLER_6_2628 ();
 sg13g2_decap_8 FILLER_6_2635 ();
 sg13g2_decap_8 FILLER_6_2642 ();
 sg13g2_decap_8 FILLER_6_2649 ();
 sg13g2_decap_8 FILLER_6_2656 ();
 sg13g2_decap_8 FILLER_6_2663 ();
 sg13g2_decap_4 FILLER_6_2670 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_fill_2 FILLER_7_252 ();
 sg13g2_fill_1 FILLER_7_254 ();
 sg13g2_fill_2 FILLER_7_259 ();
 sg13g2_fill_1 FILLER_7_261 ();
 sg13g2_fill_1 FILLER_7_323 ();
 sg13g2_decap_8 FILLER_7_431 ();
 sg13g2_decap_8 FILLER_7_438 ();
 sg13g2_decap_8 FILLER_7_445 ();
 sg13g2_decap_8 FILLER_7_452 ();
 sg13g2_decap_8 FILLER_7_459 ();
 sg13g2_decap_8 FILLER_7_466 ();
 sg13g2_decap_8 FILLER_7_473 ();
 sg13g2_decap_8 FILLER_7_480 ();
 sg13g2_decap_8 FILLER_7_487 ();
 sg13g2_decap_8 FILLER_7_494 ();
 sg13g2_decap_8 FILLER_7_501 ();
 sg13g2_decap_8 FILLER_7_508 ();
 sg13g2_decap_8 FILLER_7_515 ();
 sg13g2_decap_8 FILLER_7_522 ();
 sg13g2_decap_8 FILLER_7_555 ();
 sg13g2_decap_8 FILLER_7_562 ();
 sg13g2_decap_8 FILLER_7_569 ();
 sg13g2_decap_8 FILLER_7_576 ();
 sg13g2_fill_2 FILLER_7_583 ();
 sg13g2_fill_1 FILLER_7_585 ();
 sg13g2_decap_4 FILLER_7_595 ();
 sg13g2_fill_1 FILLER_7_599 ();
 sg13g2_fill_2 FILLER_7_682 ();
 sg13g2_decap_8 FILLER_7_726 ();
 sg13g2_decap_8 FILLER_7_733 ();
 sg13g2_decap_8 FILLER_7_740 ();
 sg13g2_decap_8 FILLER_7_747 ();
 sg13g2_decap_8 FILLER_7_754 ();
 sg13g2_decap_8 FILLER_7_761 ();
 sg13g2_decap_8 FILLER_7_768 ();
 sg13g2_decap_8 FILLER_7_775 ();
 sg13g2_decap_8 FILLER_7_782 ();
 sg13g2_decap_8 FILLER_7_789 ();
 sg13g2_decap_8 FILLER_7_796 ();
 sg13g2_decap_8 FILLER_7_803 ();
 sg13g2_decap_8 FILLER_7_810 ();
 sg13g2_decap_8 FILLER_7_817 ();
 sg13g2_decap_8 FILLER_7_824 ();
 sg13g2_decap_8 FILLER_7_831 ();
 sg13g2_decap_8 FILLER_7_838 ();
 sg13g2_decap_8 FILLER_7_845 ();
 sg13g2_decap_8 FILLER_7_852 ();
 sg13g2_decap_8 FILLER_7_859 ();
 sg13g2_decap_8 FILLER_7_866 ();
 sg13g2_decap_8 FILLER_7_873 ();
 sg13g2_decap_8 FILLER_7_880 ();
 sg13g2_decap_8 FILLER_7_887 ();
 sg13g2_decap_8 FILLER_7_894 ();
 sg13g2_decap_8 FILLER_7_901 ();
 sg13g2_decap_4 FILLER_7_908 ();
 sg13g2_fill_1 FILLER_7_919 ();
 sg13g2_fill_2 FILLER_7_944 ();
 sg13g2_fill_1 FILLER_7_961 ();
 sg13g2_fill_1 FILLER_7_987 ();
 sg13g2_fill_2 FILLER_7_1020 ();
 sg13g2_fill_2 FILLER_7_1105 ();
 sg13g2_fill_2 FILLER_7_1172 ();
 sg13g2_fill_2 FILLER_7_1254 ();
 sg13g2_fill_2 FILLER_7_1265 ();
 sg13g2_fill_1 FILLER_7_1329 ();
 sg13g2_fill_2 FILLER_7_1366 ();
 sg13g2_fill_2 FILLER_7_1373 ();
 sg13g2_fill_1 FILLER_7_1425 ();
 sg13g2_fill_1 FILLER_7_1514 ();
 sg13g2_fill_1 FILLER_7_1724 ();
 sg13g2_fill_2 FILLER_7_1730 ();
 sg13g2_fill_1 FILLER_7_1732 ();
 sg13g2_decap_8 FILLER_7_1767 ();
 sg13g2_decap_4 FILLER_7_1778 ();
 sg13g2_decap_8 FILLER_7_1786 ();
 sg13g2_fill_2 FILLER_7_1793 ();
 sg13g2_fill_1 FILLER_7_1874 ();
 sg13g2_fill_2 FILLER_7_1886 ();
 sg13g2_fill_2 FILLER_7_1900 ();
 sg13g2_fill_2 FILLER_7_1908 ();
 sg13g2_fill_1 FILLER_7_1910 ();
 sg13g2_decap_8 FILLER_7_1921 ();
 sg13g2_fill_2 FILLER_7_1969 ();
 sg13g2_fill_2 FILLER_7_1985 ();
 sg13g2_fill_2 FILLER_7_1997 ();
 sg13g2_fill_2 FILLER_7_2034 ();
 sg13g2_fill_1 FILLER_7_2036 ();
 sg13g2_decap_8 FILLER_7_2047 ();
 sg13g2_decap_4 FILLER_7_2072 ();
 sg13g2_fill_2 FILLER_7_2126 ();
 sg13g2_fill_1 FILLER_7_2128 ();
 sg13g2_decap_4 FILLER_7_2159 ();
 sg13g2_fill_1 FILLER_7_2163 ();
 sg13g2_fill_1 FILLER_7_2168 ();
 sg13g2_decap_8 FILLER_7_2179 ();
 sg13g2_fill_2 FILLER_7_2186 ();
 sg13g2_decap_4 FILLER_7_2224 ();
 sg13g2_fill_2 FILLER_7_2277 ();
 sg13g2_decap_4 FILLER_7_2293 ();
 sg13g2_decap_8 FILLER_7_2310 ();
 sg13g2_decap_8 FILLER_7_2317 ();
 sg13g2_decap_8 FILLER_7_2324 ();
 sg13g2_decap_8 FILLER_7_2331 ();
 sg13g2_decap_8 FILLER_7_2338 ();
 sg13g2_decap_8 FILLER_7_2345 ();
 sg13g2_decap_8 FILLER_7_2352 ();
 sg13g2_decap_8 FILLER_7_2359 ();
 sg13g2_decap_8 FILLER_7_2366 ();
 sg13g2_decap_8 FILLER_7_2373 ();
 sg13g2_decap_8 FILLER_7_2380 ();
 sg13g2_decap_8 FILLER_7_2387 ();
 sg13g2_decap_8 FILLER_7_2394 ();
 sg13g2_decap_8 FILLER_7_2401 ();
 sg13g2_decap_8 FILLER_7_2408 ();
 sg13g2_decap_8 FILLER_7_2415 ();
 sg13g2_decap_8 FILLER_7_2422 ();
 sg13g2_decap_8 FILLER_7_2429 ();
 sg13g2_decap_8 FILLER_7_2436 ();
 sg13g2_decap_8 FILLER_7_2443 ();
 sg13g2_decap_8 FILLER_7_2450 ();
 sg13g2_decap_8 FILLER_7_2457 ();
 sg13g2_decap_8 FILLER_7_2464 ();
 sg13g2_decap_8 FILLER_7_2471 ();
 sg13g2_decap_8 FILLER_7_2478 ();
 sg13g2_decap_8 FILLER_7_2485 ();
 sg13g2_decap_8 FILLER_7_2492 ();
 sg13g2_decap_8 FILLER_7_2499 ();
 sg13g2_decap_8 FILLER_7_2506 ();
 sg13g2_decap_8 FILLER_7_2513 ();
 sg13g2_decap_8 FILLER_7_2520 ();
 sg13g2_decap_8 FILLER_7_2527 ();
 sg13g2_decap_8 FILLER_7_2534 ();
 sg13g2_decap_8 FILLER_7_2541 ();
 sg13g2_decap_8 FILLER_7_2548 ();
 sg13g2_decap_8 FILLER_7_2555 ();
 sg13g2_decap_8 FILLER_7_2562 ();
 sg13g2_decap_8 FILLER_7_2569 ();
 sg13g2_decap_8 FILLER_7_2576 ();
 sg13g2_decap_8 FILLER_7_2583 ();
 sg13g2_decap_8 FILLER_7_2590 ();
 sg13g2_decap_8 FILLER_7_2597 ();
 sg13g2_decap_8 FILLER_7_2604 ();
 sg13g2_decap_8 FILLER_7_2611 ();
 sg13g2_decap_8 FILLER_7_2618 ();
 sg13g2_decap_8 FILLER_7_2625 ();
 sg13g2_decap_8 FILLER_7_2632 ();
 sg13g2_decap_8 FILLER_7_2639 ();
 sg13g2_decap_8 FILLER_7_2646 ();
 sg13g2_decap_8 FILLER_7_2653 ();
 sg13g2_decap_8 FILLER_7_2660 ();
 sg13g2_decap_8 FILLER_7_2667 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_4 FILLER_8_224 ();
 sg13g2_fill_2 FILLER_8_228 ();
 sg13g2_decap_4 FILLER_8_239 ();
 sg13g2_fill_2 FILLER_8_243 ();
 sg13g2_fill_1 FILLER_8_341 ();
 sg13g2_fill_2 FILLER_8_385 ();
 sg13g2_fill_2 FILLER_8_400 ();
 sg13g2_fill_2 FILLER_8_408 ();
 sg13g2_fill_2 FILLER_8_449 ();
 sg13g2_fill_1 FILLER_8_451 ();
 sg13g2_decap_8 FILLER_8_457 ();
 sg13g2_decap_4 FILLER_8_464 ();
 sg13g2_fill_2 FILLER_8_468 ();
 sg13g2_decap_8 FILLER_8_474 ();
 sg13g2_decap_8 FILLER_8_481 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_fill_1 FILLER_8_518 ();
 sg13g2_fill_2 FILLER_8_538 ();
 sg13g2_fill_2 FILLER_8_549 ();
 sg13g2_decap_8 FILLER_8_559 ();
 sg13g2_decap_8 FILLER_8_566 ();
 sg13g2_decap_4 FILLER_8_573 ();
 sg13g2_fill_2 FILLER_8_577 ();
 sg13g2_fill_1 FILLER_8_635 ();
 sg13g2_fill_2 FILLER_8_645 ();
 sg13g2_fill_2 FILLER_8_689 ();
 sg13g2_fill_2 FILLER_8_702 ();
 sg13g2_fill_1 FILLER_8_704 ();
 sg13g2_fill_2 FILLER_8_731 ();
 sg13g2_decap_8 FILLER_8_738 ();
 sg13g2_decap_8 FILLER_8_745 ();
 sg13g2_decap_8 FILLER_8_752 ();
 sg13g2_decap_8 FILLER_8_759 ();
 sg13g2_decap_8 FILLER_8_766 ();
 sg13g2_decap_8 FILLER_8_773 ();
 sg13g2_decap_8 FILLER_8_780 ();
 sg13g2_decap_8 FILLER_8_787 ();
 sg13g2_decap_8 FILLER_8_794 ();
 sg13g2_decap_8 FILLER_8_801 ();
 sg13g2_decap_8 FILLER_8_808 ();
 sg13g2_decap_8 FILLER_8_815 ();
 sg13g2_decap_8 FILLER_8_822 ();
 sg13g2_decap_8 FILLER_8_829 ();
 sg13g2_decap_8 FILLER_8_836 ();
 sg13g2_decap_8 FILLER_8_843 ();
 sg13g2_decap_8 FILLER_8_850 ();
 sg13g2_decap_8 FILLER_8_857 ();
 sg13g2_decap_8 FILLER_8_864 ();
 sg13g2_decap_8 FILLER_8_871 ();
 sg13g2_decap_8 FILLER_8_878 ();
 sg13g2_decap_8 FILLER_8_885 ();
 sg13g2_decap_8 FILLER_8_892 ();
 sg13g2_decap_4 FILLER_8_899 ();
 sg13g2_fill_2 FILLER_8_994 ();
 sg13g2_fill_1 FILLER_8_1005 ();
 sg13g2_fill_2 FILLER_8_1035 ();
 sg13g2_fill_2 FILLER_8_1078 ();
 sg13g2_fill_1 FILLER_8_1169 ();
 sg13g2_fill_2 FILLER_8_1205 ();
 sg13g2_fill_1 FILLER_8_1391 ();
 sg13g2_fill_1 FILLER_8_1401 ();
 sg13g2_fill_1 FILLER_8_1457 ();
 sg13g2_fill_2 FILLER_8_1472 ();
 sg13g2_fill_2 FILLER_8_1530 ();
 sg13g2_fill_1 FILLER_8_1586 ();
 sg13g2_fill_2 FILLER_8_1596 ();
 sg13g2_fill_2 FILLER_8_1617 ();
 sg13g2_fill_1 FILLER_8_1646 ();
 sg13g2_fill_2 FILLER_8_1706 ();
 sg13g2_fill_1 FILLER_8_1708 ();
 sg13g2_fill_2 FILLER_8_1725 ();
 sg13g2_fill_1 FILLER_8_1727 ();
 sg13g2_fill_2 FILLER_8_1741 ();
 sg13g2_fill_2 FILLER_8_1764 ();
 sg13g2_fill_2 FILLER_8_1794 ();
 sg13g2_fill_1 FILLER_8_1804 ();
 sg13g2_decap_4 FILLER_8_1816 ();
 sg13g2_decap_4 FILLER_8_1843 ();
 sg13g2_fill_2 FILLER_8_1899 ();
 sg13g2_fill_1 FILLER_8_1901 ();
 sg13g2_decap_8 FILLER_8_1927 ();
 sg13g2_fill_2 FILLER_8_1934 ();
 sg13g2_fill_2 FILLER_8_1976 ();
 sg13g2_fill_1 FILLER_8_1978 ();
 sg13g2_decap_4 FILLER_8_2006 ();
 sg13g2_fill_1 FILLER_8_2014 ();
 sg13g2_decap_4 FILLER_8_2020 ();
 sg13g2_fill_1 FILLER_8_2138 ();
 sg13g2_fill_2 FILLER_8_2205 ();
 sg13g2_fill_1 FILLER_8_2207 ();
 sg13g2_decap_4 FILLER_8_2221 ();
 sg13g2_fill_2 FILLER_8_2239 ();
 sg13g2_fill_1 FILLER_8_2247 ();
 sg13g2_fill_2 FILLER_8_2284 ();
 sg13g2_decap_8 FILLER_8_2312 ();
 sg13g2_decap_8 FILLER_8_2319 ();
 sg13g2_decap_8 FILLER_8_2326 ();
 sg13g2_decap_8 FILLER_8_2333 ();
 sg13g2_decap_8 FILLER_8_2340 ();
 sg13g2_decap_8 FILLER_8_2347 ();
 sg13g2_decap_8 FILLER_8_2354 ();
 sg13g2_decap_8 FILLER_8_2361 ();
 sg13g2_decap_8 FILLER_8_2368 ();
 sg13g2_decap_8 FILLER_8_2375 ();
 sg13g2_decap_8 FILLER_8_2382 ();
 sg13g2_decap_8 FILLER_8_2389 ();
 sg13g2_decap_8 FILLER_8_2396 ();
 sg13g2_decap_8 FILLER_8_2403 ();
 sg13g2_decap_8 FILLER_8_2410 ();
 sg13g2_decap_8 FILLER_8_2417 ();
 sg13g2_decap_8 FILLER_8_2424 ();
 sg13g2_decap_8 FILLER_8_2431 ();
 sg13g2_decap_8 FILLER_8_2438 ();
 sg13g2_decap_8 FILLER_8_2445 ();
 sg13g2_decap_8 FILLER_8_2452 ();
 sg13g2_decap_8 FILLER_8_2459 ();
 sg13g2_decap_8 FILLER_8_2466 ();
 sg13g2_decap_8 FILLER_8_2473 ();
 sg13g2_decap_8 FILLER_8_2480 ();
 sg13g2_decap_8 FILLER_8_2487 ();
 sg13g2_decap_8 FILLER_8_2494 ();
 sg13g2_decap_8 FILLER_8_2501 ();
 sg13g2_decap_8 FILLER_8_2508 ();
 sg13g2_decap_8 FILLER_8_2515 ();
 sg13g2_decap_8 FILLER_8_2522 ();
 sg13g2_decap_8 FILLER_8_2529 ();
 sg13g2_decap_8 FILLER_8_2536 ();
 sg13g2_decap_8 FILLER_8_2543 ();
 sg13g2_decap_8 FILLER_8_2550 ();
 sg13g2_decap_8 FILLER_8_2557 ();
 sg13g2_decap_8 FILLER_8_2564 ();
 sg13g2_decap_8 FILLER_8_2571 ();
 sg13g2_decap_8 FILLER_8_2578 ();
 sg13g2_decap_8 FILLER_8_2585 ();
 sg13g2_decap_8 FILLER_8_2592 ();
 sg13g2_decap_8 FILLER_8_2599 ();
 sg13g2_decap_8 FILLER_8_2606 ();
 sg13g2_decap_8 FILLER_8_2613 ();
 sg13g2_decap_8 FILLER_8_2620 ();
 sg13g2_decap_8 FILLER_8_2627 ();
 sg13g2_decap_8 FILLER_8_2634 ();
 sg13g2_decap_8 FILLER_8_2641 ();
 sg13g2_decap_8 FILLER_8_2648 ();
 sg13g2_decap_8 FILLER_8_2655 ();
 sg13g2_decap_8 FILLER_8_2662 ();
 sg13g2_decap_4 FILLER_8_2669 ();
 sg13g2_fill_1 FILLER_8_2673 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_4 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_204 ();
 sg13g2_decap_4 FILLER_9_211 ();
 sg13g2_decap_4 FILLER_9_220 ();
 sg13g2_fill_2 FILLER_9_224 ();
 sg13g2_fill_1 FILLER_9_301 ();
 sg13g2_decap_4 FILLER_9_323 ();
 sg13g2_fill_1 FILLER_9_338 ();
 sg13g2_fill_2 FILLER_9_372 ();
 sg13g2_fill_1 FILLER_9_374 ();
 sg13g2_fill_2 FILLER_9_379 ();
 sg13g2_fill_1 FILLER_9_381 ();
 sg13g2_fill_1 FILLER_9_412 ();
 sg13g2_fill_1 FILLER_9_433 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_fill_1 FILLER_9_448 ();
 sg13g2_fill_2 FILLER_9_454 ();
 sg13g2_fill_1 FILLER_9_473 ();
 sg13g2_fill_2 FILLER_9_478 ();
 sg13g2_fill_1 FILLER_9_480 ();
 sg13g2_decap_4 FILLER_9_510 ();
 sg13g2_fill_1 FILLER_9_514 ();
 sg13g2_decap_4 FILLER_9_538 ();
 sg13g2_fill_2 FILLER_9_542 ();
 sg13g2_fill_1 FILLER_9_547 ();
 sg13g2_fill_2 FILLER_9_552 ();
 sg13g2_fill_1 FILLER_9_559 ();
 sg13g2_fill_1 FILLER_9_594 ();
 sg13g2_fill_1 FILLER_9_659 ();
 sg13g2_fill_1 FILLER_9_675 ();
 sg13g2_fill_1 FILLER_9_693 ();
 sg13g2_fill_1 FILLER_9_698 ();
 sg13g2_decap_4 FILLER_9_746 ();
 sg13g2_decap_4 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_771 ();
 sg13g2_decap_8 FILLER_9_778 ();
 sg13g2_decap_8 FILLER_9_785 ();
 sg13g2_decap_8 FILLER_9_792 ();
 sg13g2_decap_8 FILLER_9_799 ();
 sg13g2_decap_8 FILLER_9_806 ();
 sg13g2_decap_8 FILLER_9_813 ();
 sg13g2_decap_8 FILLER_9_820 ();
 sg13g2_fill_1 FILLER_9_827 ();
 sg13g2_decap_8 FILLER_9_837 ();
 sg13g2_decap_8 FILLER_9_844 ();
 sg13g2_decap_8 FILLER_9_851 ();
 sg13g2_decap_8 FILLER_9_858 ();
 sg13g2_decap_8 FILLER_9_865 ();
 sg13g2_decap_8 FILLER_9_872 ();
 sg13g2_decap_8 FILLER_9_879 ();
 sg13g2_decap_8 FILLER_9_886 ();
 sg13g2_decap_4 FILLER_9_893 ();
 sg13g2_fill_1 FILLER_9_954 ();
 sg13g2_fill_2 FILLER_9_1055 ();
 sg13g2_fill_1 FILLER_9_1080 ();
 sg13g2_fill_1 FILLER_9_1107 ();
 sg13g2_fill_2 FILLER_9_1178 ();
 sg13g2_fill_2 FILLER_9_1195 ();
 sg13g2_fill_2 FILLER_9_1244 ();
 sg13g2_fill_1 FILLER_9_1267 ();
 sg13g2_fill_2 FILLER_9_1294 ();
 sg13g2_fill_1 FILLER_9_1341 ();
 sg13g2_fill_2 FILLER_9_1374 ();
 sg13g2_fill_1 FILLER_9_1416 ();
 sg13g2_fill_1 FILLER_9_1532 ();
 sg13g2_fill_1 FILLER_9_1583 ();
 sg13g2_fill_2 FILLER_9_1610 ();
 sg13g2_fill_2 FILLER_9_1756 ();
 sg13g2_fill_1 FILLER_9_1834 ();
 sg13g2_fill_1 FILLER_9_1840 ();
 sg13g2_fill_1 FILLER_9_1876 ();
 sg13g2_decap_4 FILLER_9_1912 ();
 sg13g2_fill_1 FILLER_9_1935 ();
 sg13g2_fill_2 FILLER_9_1955 ();
 sg13g2_fill_1 FILLER_9_1957 ();
 sg13g2_decap_4 FILLER_9_1993 ();
 sg13g2_fill_2 FILLER_9_2006 ();
 sg13g2_fill_1 FILLER_9_2008 ();
 sg13g2_fill_1 FILLER_9_2030 ();
 sg13g2_fill_2 FILLER_9_2042 ();
 sg13g2_fill_1 FILLER_9_2044 ();
 sg13g2_fill_2 FILLER_9_2098 ();
 sg13g2_decap_4 FILLER_9_2136 ();
 sg13g2_fill_2 FILLER_9_2140 ();
 sg13g2_decap_4 FILLER_9_2151 ();
 sg13g2_fill_2 FILLER_9_2160 ();
 sg13g2_fill_1 FILLER_9_2162 ();
 sg13g2_decap_8 FILLER_9_2172 ();
 sg13g2_fill_1 FILLER_9_2179 ();
 sg13g2_decap_4 FILLER_9_2204 ();
 sg13g2_fill_2 FILLER_9_2213 ();
 sg13g2_fill_1 FILLER_9_2250 ();
 sg13g2_decap_4 FILLER_9_2275 ();
 sg13g2_fill_2 FILLER_9_2292 ();
 sg13g2_decap_8 FILLER_9_2320 ();
 sg13g2_decap_8 FILLER_9_2327 ();
 sg13g2_decap_8 FILLER_9_2334 ();
 sg13g2_decap_8 FILLER_9_2341 ();
 sg13g2_decap_8 FILLER_9_2348 ();
 sg13g2_decap_8 FILLER_9_2355 ();
 sg13g2_decap_8 FILLER_9_2362 ();
 sg13g2_decap_8 FILLER_9_2369 ();
 sg13g2_decap_8 FILLER_9_2376 ();
 sg13g2_decap_8 FILLER_9_2383 ();
 sg13g2_decap_8 FILLER_9_2390 ();
 sg13g2_decap_8 FILLER_9_2397 ();
 sg13g2_decap_8 FILLER_9_2404 ();
 sg13g2_decap_8 FILLER_9_2411 ();
 sg13g2_decap_8 FILLER_9_2418 ();
 sg13g2_decap_8 FILLER_9_2425 ();
 sg13g2_decap_8 FILLER_9_2432 ();
 sg13g2_decap_8 FILLER_9_2439 ();
 sg13g2_decap_8 FILLER_9_2446 ();
 sg13g2_decap_8 FILLER_9_2453 ();
 sg13g2_decap_8 FILLER_9_2460 ();
 sg13g2_decap_8 FILLER_9_2467 ();
 sg13g2_decap_8 FILLER_9_2474 ();
 sg13g2_decap_8 FILLER_9_2481 ();
 sg13g2_decap_8 FILLER_9_2488 ();
 sg13g2_decap_8 FILLER_9_2495 ();
 sg13g2_decap_8 FILLER_9_2502 ();
 sg13g2_decap_8 FILLER_9_2509 ();
 sg13g2_decap_8 FILLER_9_2516 ();
 sg13g2_decap_8 FILLER_9_2523 ();
 sg13g2_decap_8 FILLER_9_2530 ();
 sg13g2_decap_8 FILLER_9_2537 ();
 sg13g2_decap_8 FILLER_9_2544 ();
 sg13g2_decap_8 FILLER_9_2551 ();
 sg13g2_decap_8 FILLER_9_2558 ();
 sg13g2_decap_8 FILLER_9_2565 ();
 sg13g2_decap_8 FILLER_9_2572 ();
 sg13g2_decap_8 FILLER_9_2579 ();
 sg13g2_decap_8 FILLER_9_2586 ();
 sg13g2_decap_8 FILLER_9_2593 ();
 sg13g2_decap_8 FILLER_9_2600 ();
 sg13g2_decap_8 FILLER_9_2607 ();
 sg13g2_decap_8 FILLER_9_2614 ();
 sg13g2_decap_8 FILLER_9_2621 ();
 sg13g2_decap_8 FILLER_9_2628 ();
 sg13g2_decap_8 FILLER_9_2635 ();
 sg13g2_decap_8 FILLER_9_2642 ();
 sg13g2_decap_8 FILLER_9_2649 ();
 sg13g2_decap_8 FILLER_9_2656 ();
 sg13g2_decap_8 FILLER_9_2663 ();
 sg13g2_decap_4 FILLER_9_2670 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_fill_1 FILLER_10_234 ();
 sg13g2_fill_2 FILLER_10_239 ();
 sg13g2_decap_4 FILLER_10_245 ();
 sg13g2_fill_1 FILLER_10_249 ();
 sg13g2_fill_2 FILLER_10_286 ();
 sg13g2_fill_1 FILLER_10_288 ();
 sg13g2_fill_1 FILLER_10_294 ();
 sg13g2_fill_2 FILLER_10_299 ();
 sg13g2_fill_2 FILLER_10_306 ();
 sg13g2_fill_1 FILLER_10_356 ();
 sg13g2_fill_1 FILLER_10_401 ();
 sg13g2_fill_2 FILLER_10_421 ();
 sg13g2_fill_2 FILLER_10_454 ();
 sg13g2_decap_4 FILLER_10_487 ();
 sg13g2_fill_1 FILLER_10_491 ();
 sg13g2_fill_2 FILLER_10_505 ();
 sg13g2_fill_2 FILLER_10_535 ();
 sg13g2_fill_2 FILLER_10_575 ();
 sg13g2_fill_1 FILLER_10_595 ();
 sg13g2_fill_1 FILLER_10_637 ();
 sg13g2_fill_1 FILLER_10_716 ();
 sg13g2_fill_1 FILLER_10_730 ();
 sg13g2_fill_2 FILLER_10_759 ();
 sg13g2_fill_1 FILLER_10_761 ();
 sg13g2_decap_8 FILLER_10_783 ();
 sg13g2_decap_4 FILLER_10_790 ();
 sg13g2_decap_8 FILLER_10_802 ();
 sg13g2_decap_8 FILLER_10_809 ();
 sg13g2_decap_8 FILLER_10_816 ();
 sg13g2_decap_8 FILLER_10_823 ();
 sg13g2_decap_8 FILLER_10_830 ();
 sg13g2_decap_8 FILLER_10_837 ();
 sg13g2_decap_8 FILLER_10_844 ();
 sg13g2_decap_8 FILLER_10_851 ();
 sg13g2_decap_8 FILLER_10_858 ();
 sg13g2_decap_8 FILLER_10_865 ();
 sg13g2_decap_8 FILLER_10_872 ();
 sg13g2_decap_8 FILLER_10_879 ();
 sg13g2_fill_2 FILLER_10_886 ();
 sg13g2_fill_1 FILLER_10_888 ();
 sg13g2_fill_1 FILLER_10_917 ();
 sg13g2_fill_1 FILLER_10_933 ();
 sg13g2_fill_2 FILLER_10_965 ();
 sg13g2_fill_2 FILLER_10_976 ();
 sg13g2_fill_1 FILLER_10_1080 ();
 sg13g2_fill_2 FILLER_10_1102 ();
 sg13g2_fill_1 FILLER_10_1184 ();
 sg13g2_fill_1 FILLER_10_1216 ();
 sg13g2_fill_1 FILLER_10_1325 ();
 sg13g2_fill_1 FILLER_10_1394 ();
 sg13g2_fill_1 FILLER_10_1426 ();
 sg13g2_fill_1 FILLER_10_1499 ();
 sg13g2_fill_1 FILLER_10_1548 ();
 sg13g2_fill_1 FILLER_10_1639 ();
 sg13g2_fill_2 FILLER_10_1777 ();
 sg13g2_fill_1 FILLER_10_1779 ();
 sg13g2_fill_2 FILLER_10_1799 ();
 sg13g2_fill_1 FILLER_10_1910 ();
 sg13g2_decap_4 FILLER_10_1926 ();
 sg13g2_fill_2 FILLER_10_1930 ();
 sg13g2_fill_1 FILLER_10_1967 ();
 sg13g2_decap_8 FILLER_10_2027 ();
 sg13g2_fill_1 FILLER_10_2034 ();
 sg13g2_decap_4 FILLER_10_2039 ();
 sg13g2_fill_2 FILLER_10_2043 ();
 sg13g2_decap_4 FILLER_10_2059 ();
 sg13g2_decap_8 FILLER_10_2083 ();
 sg13g2_decap_4 FILLER_10_2090 ();
 sg13g2_fill_2 FILLER_10_2094 ();
 sg13g2_fill_1 FILLER_10_2106 ();
 sg13g2_fill_1 FILLER_10_2131 ();
 sg13g2_fill_2 FILLER_10_2142 ();
 sg13g2_fill_1 FILLER_10_2144 ();
 sg13g2_fill_1 FILLER_10_2165 ();
 sg13g2_fill_2 FILLER_10_2205 ();
 sg13g2_fill_1 FILLER_10_2207 ();
 sg13g2_fill_1 FILLER_10_2228 ();
 sg13g2_fill_1 FILLER_10_2285 ();
 sg13g2_decap_4 FILLER_10_2301 ();
 sg13g2_decap_8 FILLER_10_2318 ();
 sg13g2_decap_8 FILLER_10_2325 ();
 sg13g2_decap_8 FILLER_10_2332 ();
 sg13g2_decap_8 FILLER_10_2339 ();
 sg13g2_decap_8 FILLER_10_2346 ();
 sg13g2_decap_8 FILLER_10_2353 ();
 sg13g2_decap_8 FILLER_10_2360 ();
 sg13g2_decap_8 FILLER_10_2367 ();
 sg13g2_decap_8 FILLER_10_2374 ();
 sg13g2_decap_8 FILLER_10_2381 ();
 sg13g2_decap_8 FILLER_10_2388 ();
 sg13g2_decap_8 FILLER_10_2395 ();
 sg13g2_decap_8 FILLER_10_2402 ();
 sg13g2_decap_8 FILLER_10_2409 ();
 sg13g2_decap_8 FILLER_10_2416 ();
 sg13g2_decap_8 FILLER_10_2423 ();
 sg13g2_decap_8 FILLER_10_2430 ();
 sg13g2_decap_8 FILLER_10_2437 ();
 sg13g2_decap_8 FILLER_10_2444 ();
 sg13g2_decap_8 FILLER_10_2451 ();
 sg13g2_decap_8 FILLER_10_2458 ();
 sg13g2_decap_8 FILLER_10_2465 ();
 sg13g2_decap_8 FILLER_10_2472 ();
 sg13g2_decap_8 FILLER_10_2479 ();
 sg13g2_decap_8 FILLER_10_2486 ();
 sg13g2_decap_8 FILLER_10_2493 ();
 sg13g2_decap_8 FILLER_10_2500 ();
 sg13g2_decap_8 FILLER_10_2507 ();
 sg13g2_decap_8 FILLER_10_2514 ();
 sg13g2_decap_8 FILLER_10_2521 ();
 sg13g2_decap_8 FILLER_10_2528 ();
 sg13g2_decap_8 FILLER_10_2535 ();
 sg13g2_decap_8 FILLER_10_2542 ();
 sg13g2_decap_8 FILLER_10_2549 ();
 sg13g2_decap_8 FILLER_10_2556 ();
 sg13g2_decap_8 FILLER_10_2563 ();
 sg13g2_decap_8 FILLER_10_2570 ();
 sg13g2_decap_8 FILLER_10_2577 ();
 sg13g2_decap_8 FILLER_10_2584 ();
 sg13g2_decap_8 FILLER_10_2591 ();
 sg13g2_decap_8 FILLER_10_2598 ();
 sg13g2_decap_8 FILLER_10_2605 ();
 sg13g2_decap_8 FILLER_10_2612 ();
 sg13g2_decap_8 FILLER_10_2619 ();
 sg13g2_decap_8 FILLER_10_2626 ();
 sg13g2_decap_8 FILLER_10_2633 ();
 sg13g2_decap_8 FILLER_10_2640 ();
 sg13g2_decap_8 FILLER_10_2647 ();
 sg13g2_decap_8 FILLER_10_2654 ();
 sg13g2_decap_8 FILLER_10_2661 ();
 sg13g2_decap_4 FILLER_10_2668 ();
 sg13g2_fill_2 FILLER_10_2672 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_204 ();
 sg13g2_fill_1 FILLER_11_211 ();
 sg13g2_decap_4 FILLER_11_224 ();
 sg13g2_decap_4 FILLER_11_241 ();
 sg13g2_fill_1 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_251 ();
 sg13g2_fill_2 FILLER_11_258 ();
 sg13g2_fill_2 FILLER_11_264 ();
 sg13g2_fill_1 FILLER_11_266 ();
 sg13g2_fill_2 FILLER_11_302 ();
 sg13g2_fill_1 FILLER_11_304 ();
 sg13g2_decap_4 FILLER_11_331 ();
 sg13g2_fill_2 FILLER_11_335 ();
 sg13g2_fill_1 FILLER_11_350 ();
 sg13g2_fill_1 FILLER_11_356 ();
 sg13g2_fill_1 FILLER_11_372 ();
 sg13g2_fill_2 FILLER_11_382 ();
 sg13g2_fill_1 FILLER_11_400 ();
 sg13g2_fill_1 FILLER_11_466 ();
 sg13g2_fill_1 FILLER_11_489 ();
 sg13g2_decap_8 FILLER_11_500 ();
 sg13g2_fill_2 FILLER_11_507 ();
 sg13g2_fill_1 FILLER_11_509 ();
 sg13g2_fill_2 FILLER_11_518 ();
 sg13g2_decap_4 FILLER_11_525 ();
 sg13g2_fill_1 FILLER_11_529 ();
 sg13g2_decap_8 FILLER_11_540 ();
 sg13g2_decap_4 FILLER_11_547 ();
 sg13g2_fill_2 FILLER_11_551 ();
 sg13g2_decap_8 FILLER_11_561 ();
 sg13g2_fill_1 FILLER_11_568 ();
 sg13g2_fill_2 FILLER_11_625 ();
 sg13g2_fill_1 FILLER_11_658 ();
 sg13g2_fill_2 FILLER_11_677 ();
 sg13g2_fill_1 FILLER_11_687 ();
 sg13g2_fill_2 FILLER_11_740 ();
 sg13g2_fill_1 FILLER_11_742 ();
 sg13g2_fill_1 FILLER_11_751 ();
 sg13g2_fill_1 FILLER_11_762 ();
 sg13g2_decap_8 FILLER_11_768 ();
 sg13g2_fill_2 FILLER_11_775 ();
 sg13g2_fill_1 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_809 ();
 sg13g2_decap_8 FILLER_11_816 ();
 sg13g2_decap_8 FILLER_11_823 ();
 sg13g2_decap_8 FILLER_11_830 ();
 sg13g2_decap_8 FILLER_11_837 ();
 sg13g2_decap_8 FILLER_11_844 ();
 sg13g2_decap_8 FILLER_11_851 ();
 sg13g2_decap_8 FILLER_11_858 ();
 sg13g2_decap_8 FILLER_11_865 ();
 sg13g2_decap_8 FILLER_11_872 ();
 sg13g2_fill_2 FILLER_11_1001 ();
 sg13g2_fill_1 FILLER_11_1026 ();
 sg13g2_fill_1 FILLER_11_1084 ();
 sg13g2_fill_2 FILLER_11_1163 ();
 sg13g2_fill_2 FILLER_11_1207 ();
 sg13g2_fill_2 FILLER_11_1325 ();
 sg13g2_fill_1 FILLER_11_1362 ();
 sg13g2_fill_2 FILLER_11_1369 ();
 sg13g2_fill_1 FILLER_11_1412 ();
 sg13g2_fill_2 FILLER_11_1418 ();
 sg13g2_fill_1 FILLER_11_1495 ();
 sg13g2_fill_1 FILLER_11_1558 ();
 sg13g2_fill_1 FILLER_11_1590 ();
 sg13g2_fill_2 FILLER_11_1732 ();
 sg13g2_fill_2 FILLER_11_1761 ();
 sg13g2_fill_1 FILLER_11_1794 ();
 sg13g2_fill_2 FILLER_11_1852 ();
 sg13g2_fill_2 FILLER_11_1869 ();
 sg13g2_fill_1 FILLER_11_1871 ();
 sg13g2_fill_2 FILLER_11_1889 ();
 sg13g2_fill_1 FILLER_11_1891 ();
 sg13g2_decap_8 FILLER_11_1897 ();
 sg13g2_decap_4 FILLER_11_1914 ();
 sg13g2_fill_2 FILLER_11_1944 ();
 sg13g2_fill_2 FILLER_11_1982 ();
 sg13g2_decap_8 FILLER_11_1989 ();
 sg13g2_fill_1 FILLER_11_1996 ();
 sg13g2_fill_2 FILLER_11_2021 ();
 sg13g2_fill_1 FILLER_11_2023 ();
 sg13g2_fill_2 FILLER_11_2050 ();
 sg13g2_fill_2 FILLER_11_2085 ();
 sg13g2_decap_4 FILLER_11_2113 ();
 sg13g2_fill_2 FILLER_11_2117 ();
 sg13g2_decap_4 FILLER_11_2160 ();
 sg13g2_fill_2 FILLER_11_2192 ();
 sg13g2_decap_8 FILLER_11_2203 ();
 sg13g2_fill_1 FILLER_11_2220 ();
 sg13g2_decap_8 FILLER_11_2226 ();
 sg13g2_fill_2 FILLER_11_2233 ();
 sg13g2_fill_2 FILLER_11_2257 ();
 sg13g2_decap_8 FILLER_11_2277 ();
 sg13g2_fill_2 FILLER_11_2284 ();
 sg13g2_fill_1 FILLER_11_2286 ();
 sg13g2_decap_8 FILLER_11_2323 ();
 sg13g2_decap_8 FILLER_11_2330 ();
 sg13g2_decap_8 FILLER_11_2337 ();
 sg13g2_decap_8 FILLER_11_2344 ();
 sg13g2_decap_8 FILLER_11_2351 ();
 sg13g2_decap_8 FILLER_11_2358 ();
 sg13g2_decap_8 FILLER_11_2365 ();
 sg13g2_decap_8 FILLER_11_2372 ();
 sg13g2_decap_8 FILLER_11_2379 ();
 sg13g2_decap_8 FILLER_11_2386 ();
 sg13g2_decap_8 FILLER_11_2393 ();
 sg13g2_decap_8 FILLER_11_2400 ();
 sg13g2_decap_8 FILLER_11_2407 ();
 sg13g2_decap_8 FILLER_11_2414 ();
 sg13g2_decap_8 FILLER_11_2421 ();
 sg13g2_decap_8 FILLER_11_2428 ();
 sg13g2_decap_8 FILLER_11_2435 ();
 sg13g2_decap_8 FILLER_11_2442 ();
 sg13g2_decap_8 FILLER_11_2449 ();
 sg13g2_decap_8 FILLER_11_2456 ();
 sg13g2_decap_8 FILLER_11_2463 ();
 sg13g2_decap_8 FILLER_11_2470 ();
 sg13g2_decap_8 FILLER_11_2477 ();
 sg13g2_decap_8 FILLER_11_2484 ();
 sg13g2_decap_8 FILLER_11_2491 ();
 sg13g2_decap_8 FILLER_11_2498 ();
 sg13g2_decap_8 FILLER_11_2505 ();
 sg13g2_decap_8 FILLER_11_2512 ();
 sg13g2_decap_8 FILLER_11_2519 ();
 sg13g2_decap_8 FILLER_11_2526 ();
 sg13g2_decap_8 FILLER_11_2533 ();
 sg13g2_decap_8 FILLER_11_2540 ();
 sg13g2_decap_8 FILLER_11_2547 ();
 sg13g2_decap_8 FILLER_11_2554 ();
 sg13g2_decap_8 FILLER_11_2561 ();
 sg13g2_decap_8 FILLER_11_2568 ();
 sg13g2_decap_8 FILLER_11_2575 ();
 sg13g2_decap_8 FILLER_11_2582 ();
 sg13g2_decap_8 FILLER_11_2589 ();
 sg13g2_decap_8 FILLER_11_2596 ();
 sg13g2_decap_8 FILLER_11_2603 ();
 sg13g2_decap_8 FILLER_11_2610 ();
 sg13g2_decap_8 FILLER_11_2617 ();
 sg13g2_decap_8 FILLER_11_2624 ();
 sg13g2_decap_8 FILLER_11_2631 ();
 sg13g2_decap_8 FILLER_11_2638 ();
 sg13g2_decap_8 FILLER_11_2645 ();
 sg13g2_decap_8 FILLER_11_2652 ();
 sg13g2_decap_8 FILLER_11_2659 ();
 sg13g2_decap_8 FILLER_11_2666 ();
 sg13g2_fill_1 FILLER_11_2673 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_4 FILLER_12_161 ();
 sg13g2_fill_2 FILLER_12_191 ();
 sg13g2_fill_2 FILLER_12_199 ();
 sg13g2_fill_1 FILLER_12_201 ();
 sg13g2_fill_1 FILLER_12_232 ();
 sg13g2_fill_2 FILLER_12_238 ();
 sg13g2_fill_1 FILLER_12_261 ();
 sg13g2_fill_2 FILLER_12_270 ();
 sg13g2_fill_1 FILLER_12_272 ();
 sg13g2_fill_2 FILLER_12_304 ();
 sg13g2_fill_1 FILLER_12_306 ();
 sg13g2_fill_1 FILLER_12_312 ();
 sg13g2_decap_4 FILLER_12_365 ();
 sg13g2_fill_2 FILLER_12_395 ();
 sg13g2_fill_1 FILLER_12_397 ();
 sg13g2_fill_2 FILLER_12_408 ();
 sg13g2_fill_1 FILLER_12_410 ();
 sg13g2_fill_2 FILLER_12_420 ();
 sg13g2_fill_1 FILLER_12_444 ();
 sg13g2_fill_1 FILLER_12_471 ();
 sg13g2_fill_2 FILLER_12_490 ();
 sg13g2_fill_1 FILLER_12_492 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_fill_2 FILLER_12_521 ();
 sg13g2_fill_1 FILLER_12_523 ();
 sg13g2_decap_4 FILLER_12_529 ();
 sg13g2_fill_1 FILLER_12_533 ();
 sg13g2_fill_2 FILLER_12_539 ();
 sg13g2_fill_1 FILLER_12_541 ();
 sg13g2_fill_2 FILLER_12_584 ();
 sg13g2_fill_1 FILLER_12_595 ();
 sg13g2_fill_2 FILLER_12_663 ();
 sg13g2_fill_2 FILLER_12_702 ();
 sg13g2_fill_1 FILLER_12_704 ();
 sg13g2_fill_2 FILLER_12_719 ();
 sg13g2_fill_1 FILLER_12_721 ();
 sg13g2_fill_2 FILLER_12_753 ();
 sg13g2_fill_1 FILLER_12_755 ();
 sg13g2_decap_8 FILLER_12_773 ();
 sg13g2_decap_8 FILLER_12_780 ();
 sg13g2_fill_1 FILLER_12_787 ();
 sg13g2_decap_8 FILLER_12_792 ();
 sg13g2_decap_8 FILLER_12_799 ();
 sg13g2_decap_8 FILLER_12_806 ();
 sg13g2_decap_8 FILLER_12_813 ();
 sg13g2_decap_8 FILLER_12_820 ();
 sg13g2_decap_8 FILLER_12_827 ();
 sg13g2_decap_8 FILLER_12_834 ();
 sg13g2_decap_8 FILLER_12_841 ();
 sg13g2_decap_8 FILLER_12_848 ();
 sg13g2_decap_8 FILLER_12_855 ();
 sg13g2_decap_8 FILLER_12_862 ();
 sg13g2_decap_4 FILLER_12_869 ();
 sg13g2_fill_1 FILLER_12_873 ();
 sg13g2_fill_1 FILLER_12_987 ();
 sg13g2_fill_1 FILLER_12_1039 ();
 sg13g2_fill_1 FILLER_12_1049 ();
 sg13g2_fill_2 FILLER_12_1109 ();
 sg13g2_fill_2 FILLER_12_1121 ();
 sg13g2_fill_2 FILLER_12_1186 ();
 sg13g2_fill_2 FILLER_12_1197 ();
 sg13g2_fill_1 FILLER_12_1383 ();
 sg13g2_fill_2 FILLER_12_1483 ();
 sg13g2_fill_1 FILLER_12_1583 ();
 sg13g2_fill_2 FILLER_12_1603 ();
 sg13g2_fill_2 FILLER_12_1656 ();
 sg13g2_fill_1 FILLER_12_1725 ();
 sg13g2_fill_2 FILLER_12_1820 ();
 sg13g2_fill_1 FILLER_12_1822 ();
 sg13g2_fill_2 FILLER_12_1859 ();
 sg13g2_decap_4 FILLER_12_1923 ();
 sg13g2_fill_2 FILLER_12_1927 ();
 sg13g2_fill_1 FILLER_12_1933 ();
 sg13g2_fill_2 FILLER_12_1963 ();
 sg13g2_fill_1 FILLER_12_1965 ();
 sg13g2_fill_2 FILLER_12_1999 ();
 sg13g2_fill_1 FILLER_12_2006 ();
 sg13g2_decap_8 FILLER_12_2017 ();
 sg13g2_decap_4 FILLER_12_2024 ();
 sg13g2_fill_1 FILLER_12_2028 ();
 sg13g2_fill_2 FILLER_12_2042 ();
 sg13g2_decap_4 FILLER_12_2077 ();
 sg13g2_decap_8 FILLER_12_2086 ();
 sg13g2_decap_4 FILLER_12_2093 ();
 sg13g2_fill_1 FILLER_12_2097 ();
 sg13g2_fill_2 FILLER_12_2108 ();
 sg13g2_fill_1 FILLER_12_2110 ();
 sg13g2_fill_2 FILLER_12_2137 ();
 sg13g2_decap_4 FILLER_12_2194 ();
 sg13g2_decap_8 FILLER_12_2202 ();
 sg13g2_decap_4 FILLER_12_2214 ();
 sg13g2_fill_1 FILLER_12_2218 ();
 sg13g2_decap_4 FILLER_12_2285 ();
 sg13g2_fill_1 FILLER_12_2289 ();
 sg13g2_fill_2 FILLER_12_2309 ();
 sg13g2_decap_8 FILLER_12_2328 ();
 sg13g2_decap_8 FILLER_12_2335 ();
 sg13g2_decap_8 FILLER_12_2342 ();
 sg13g2_decap_8 FILLER_12_2349 ();
 sg13g2_decap_8 FILLER_12_2356 ();
 sg13g2_decap_8 FILLER_12_2363 ();
 sg13g2_decap_8 FILLER_12_2370 ();
 sg13g2_decap_8 FILLER_12_2377 ();
 sg13g2_decap_8 FILLER_12_2384 ();
 sg13g2_decap_8 FILLER_12_2391 ();
 sg13g2_decap_8 FILLER_12_2398 ();
 sg13g2_decap_8 FILLER_12_2405 ();
 sg13g2_decap_8 FILLER_12_2412 ();
 sg13g2_decap_8 FILLER_12_2419 ();
 sg13g2_decap_8 FILLER_12_2426 ();
 sg13g2_decap_8 FILLER_12_2433 ();
 sg13g2_decap_8 FILLER_12_2440 ();
 sg13g2_decap_8 FILLER_12_2447 ();
 sg13g2_decap_8 FILLER_12_2454 ();
 sg13g2_decap_8 FILLER_12_2461 ();
 sg13g2_decap_8 FILLER_12_2468 ();
 sg13g2_decap_8 FILLER_12_2475 ();
 sg13g2_decap_8 FILLER_12_2482 ();
 sg13g2_decap_8 FILLER_12_2489 ();
 sg13g2_decap_8 FILLER_12_2496 ();
 sg13g2_decap_8 FILLER_12_2503 ();
 sg13g2_decap_8 FILLER_12_2510 ();
 sg13g2_decap_8 FILLER_12_2517 ();
 sg13g2_decap_8 FILLER_12_2524 ();
 sg13g2_decap_8 FILLER_12_2531 ();
 sg13g2_decap_8 FILLER_12_2538 ();
 sg13g2_decap_8 FILLER_12_2545 ();
 sg13g2_decap_8 FILLER_12_2552 ();
 sg13g2_decap_8 FILLER_12_2559 ();
 sg13g2_decap_8 FILLER_12_2566 ();
 sg13g2_decap_8 FILLER_12_2573 ();
 sg13g2_decap_8 FILLER_12_2580 ();
 sg13g2_decap_8 FILLER_12_2587 ();
 sg13g2_decap_8 FILLER_12_2594 ();
 sg13g2_decap_8 FILLER_12_2601 ();
 sg13g2_decap_8 FILLER_12_2608 ();
 sg13g2_decap_8 FILLER_12_2615 ();
 sg13g2_decap_8 FILLER_12_2622 ();
 sg13g2_decap_8 FILLER_12_2629 ();
 sg13g2_decap_8 FILLER_12_2636 ();
 sg13g2_decap_8 FILLER_12_2643 ();
 sg13g2_decap_8 FILLER_12_2650 ();
 sg13g2_decap_8 FILLER_12_2657 ();
 sg13g2_decap_8 FILLER_12_2664 ();
 sg13g2_fill_2 FILLER_12_2671 ();
 sg13g2_fill_1 FILLER_12_2673 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_fill_2 FILLER_13_175 ();
 sg13g2_fill_1 FILLER_13_177 ();
 sg13g2_fill_2 FILLER_13_212 ();
 sg13g2_fill_2 FILLER_13_241 ();
 sg13g2_fill_2 FILLER_13_256 ();
 sg13g2_fill_1 FILLER_13_258 ();
 sg13g2_fill_1 FILLER_13_274 ();
 sg13g2_decap_4 FILLER_13_285 ();
 sg13g2_fill_1 FILLER_13_289 ();
 sg13g2_fill_1 FILLER_13_294 ();
 sg13g2_fill_1 FILLER_13_300 ();
 sg13g2_decap_4 FILLER_13_322 ();
 sg13g2_fill_1 FILLER_13_358 ();
 sg13g2_fill_1 FILLER_13_363 ();
 sg13g2_fill_1 FILLER_13_412 ();
 sg13g2_fill_1 FILLER_13_431 ();
 sg13g2_decap_8 FILLER_13_446 ();
 sg13g2_fill_1 FILLER_13_453 ();
 sg13g2_fill_1 FILLER_13_494 ();
 sg13g2_fill_2 FILLER_13_511 ();
 sg13g2_fill_2 FILLER_13_518 ();
 sg13g2_fill_1 FILLER_13_520 ();
 sg13g2_decap_4 FILLER_13_565 ();
 sg13g2_fill_2 FILLER_13_569 ();
 sg13g2_fill_2 FILLER_13_625 ();
 sg13g2_fill_1 FILLER_13_627 ();
 sg13g2_fill_1 FILLER_13_643 ();
 sg13g2_fill_2 FILLER_13_680 ();
 sg13g2_fill_1 FILLER_13_682 ();
 sg13g2_fill_1 FILLER_13_697 ();
 sg13g2_fill_2 FILLER_13_712 ();
 sg13g2_fill_2 FILLER_13_756 ();
 sg13g2_fill_2 FILLER_13_779 ();
 sg13g2_fill_1 FILLER_13_781 ();
 sg13g2_fill_2 FILLER_13_786 ();
 sg13g2_fill_1 FILLER_13_788 ();
 sg13g2_decap_8 FILLER_13_801 ();
 sg13g2_decap_4 FILLER_13_808 ();
 sg13g2_fill_1 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_816 ();
 sg13g2_decap_8 FILLER_13_823 ();
 sg13g2_decap_8 FILLER_13_830 ();
 sg13g2_decap_8 FILLER_13_837 ();
 sg13g2_decap_8 FILLER_13_844 ();
 sg13g2_decap_8 FILLER_13_851 ();
 sg13g2_decap_8 FILLER_13_858 ();
 sg13g2_decap_8 FILLER_13_865 ();
 sg13g2_decap_4 FILLER_13_872 ();
 sg13g2_fill_2 FILLER_13_876 ();
 sg13g2_fill_2 FILLER_13_960 ();
 sg13g2_fill_1 FILLER_13_1014 ();
 sg13g2_fill_1 FILLER_13_1024 ();
 sg13g2_fill_2 FILLER_13_1045 ();
 sg13g2_fill_1 FILLER_13_1168 ();
 sg13g2_fill_2 FILLER_13_1357 ();
 sg13g2_fill_2 FILLER_13_1385 ();
 sg13g2_fill_1 FILLER_13_1422 ();
 sg13g2_fill_1 FILLER_13_1468 ();
 sg13g2_fill_1 FILLER_13_1631 ();
 sg13g2_fill_1 FILLER_13_1734 ();
 sg13g2_fill_1 FILLER_13_1757 ();
 sg13g2_fill_1 FILLER_13_1782 ();
 sg13g2_fill_1 FILLER_13_1800 ();
 sg13g2_fill_1 FILLER_13_1830 ();
 sg13g2_fill_2 FILLER_13_1881 ();
 sg13g2_fill_1 FILLER_13_1883 ();
 sg13g2_fill_1 FILLER_13_1912 ();
 sg13g2_fill_2 FILLER_13_1926 ();
 sg13g2_fill_2 FILLER_13_1955 ();
 sg13g2_fill_1 FILLER_13_1957 ();
 sg13g2_fill_1 FILLER_13_1967 ();
 sg13g2_fill_1 FILLER_13_1997 ();
 sg13g2_fill_1 FILLER_13_2008 ();
 sg13g2_decap_4 FILLER_13_2067 ();
 sg13g2_fill_1 FILLER_13_2083 ();
 sg13g2_decap_8 FILLER_13_2088 ();
 sg13g2_fill_2 FILLER_13_2112 ();
 sg13g2_fill_1 FILLER_13_2114 ();
 sg13g2_fill_2 FILLER_13_2121 ();
 sg13g2_fill_2 FILLER_13_2166 ();
 sg13g2_fill_2 FILLER_13_2173 ();
 sg13g2_fill_2 FILLER_13_2185 ();
 sg13g2_decap_4 FILLER_13_2213 ();
 sg13g2_fill_2 FILLER_13_2217 ();
 sg13g2_decap_8 FILLER_13_2236 ();
 sg13g2_decap_8 FILLER_13_2243 ();
 sg13g2_fill_2 FILLER_13_2250 ();
 sg13g2_fill_1 FILLER_13_2252 ();
 sg13g2_fill_1 FILLER_13_2270 ();
 sg13g2_decap_8 FILLER_13_2328 ();
 sg13g2_decap_8 FILLER_13_2335 ();
 sg13g2_decap_8 FILLER_13_2342 ();
 sg13g2_decap_8 FILLER_13_2349 ();
 sg13g2_decap_8 FILLER_13_2356 ();
 sg13g2_decap_8 FILLER_13_2363 ();
 sg13g2_decap_8 FILLER_13_2370 ();
 sg13g2_decap_8 FILLER_13_2377 ();
 sg13g2_decap_8 FILLER_13_2384 ();
 sg13g2_decap_8 FILLER_13_2391 ();
 sg13g2_decap_8 FILLER_13_2398 ();
 sg13g2_decap_8 FILLER_13_2405 ();
 sg13g2_decap_8 FILLER_13_2412 ();
 sg13g2_decap_8 FILLER_13_2419 ();
 sg13g2_decap_8 FILLER_13_2426 ();
 sg13g2_decap_8 FILLER_13_2433 ();
 sg13g2_decap_8 FILLER_13_2440 ();
 sg13g2_decap_8 FILLER_13_2447 ();
 sg13g2_decap_8 FILLER_13_2454 ();
 sg13g2_decap_8 FILLER_13_2461 ();
 sg13g2_decap_8 FILLER_13_2468 ();
 sg13g2_decap_8 FILLER_13_2475 ();
 sg13g2_decap_8 FILLER_13_2482 ();
 sg13g2_decap_8 FILLER_13_2489 ();
 sg13g2_decap_8 FILLER_13_2496 ();
 sg13g2_decap_8 FILLER_13_2503 ();
 sg13g2_decap_8 FILLER_13_2510 ();
 sg13g2_decap_8 FILLER_13_2517 ();
 sg13g2_decap_8 FILLER_13_2524 ();
 sg13g2_decap_8 FILLER_13_2531 ();
 sg13g2_decap_8 FILLER_13_2538 ();
 sg13g2_decap_8 FILLER_13_2545 ();
 sg13g2_decap_8 FILLER_13_2552 ();
 sg13g2_decap_8 FILLER_13_2559 ();
 sg13g2_decap_8 FILLER_13_2566 ();
 sg13g2_decap_8 FILLER_13_2573 ();
 sg13g2_decap_8 FILLER_13_2580 ();
 sg13g2_decap_8 FILLER_13_2587 ();
 sg13g2_decap_8 FILLER_13_2594 ();
 sg13g2_decap_8 FILLER_13_2601 ();
 sg13g2_decap_8 FILLER_13_2608 ();
 sg13g2_decap_8 FILLER_13_2615 ();
 sg13g2_decap_8 FILLER_13_2622 ();
 sg13g2_decap_8 FILLER_13_2629 ();
 sg13g2_decap_8 FILLER_13_2636 ();
 sg13g2_decap_8 FILLER_13_2643 ();
 sg13g2_decap_8 FILLER_13_2650 ();
 sg13g2_decap_8 FILLER_13_2657 ();
 sg13g2_decap_8 FILLER_13_2664 ();
 sg13g2_fill_2 FILLER_13_2671 ();
 sg13g2_fill_1 FILLER_13_2673 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_fill_1 FILLER_14_175 ();
 sg13g2_decap_4 FILLER_14_180 ();
 sg13g2_fill_1 FILLER_14_184 ();
 sg13g2_fill_2 FILLER_14_194 ();
 sg13g2_fill_1 FILLER_14_196 ();
 sg13g2_decap_4 FILLER_14_233 ();
 sg13g2_decap_4 FILLER_14_249 ();
 sg13g2_decap_4 FILLER_14_292 ();
 sg13g2_fill_2 FILLER_14_296 ();
 sg13g2_decap_8 FILLER_14_305 ();
 sg13g2_fill_1 FILLER_14_325 ();
 sg13g2_fill_1 FILLER_14_335 ();
 sg13g2_fill_2 FILLER_14_345 ();
 sg13g2_fill_1 FILLER_14_347 ();
 sg13g2_fill_2 FILLER_14_362 ();
 sg13g2_fill_1 FILLER_14_364 ();
 sg13g2_fill_1 FILLER_14_374 ();
 sg13g2_fill_2 FILLER_14_395 ();
 sg13g2_fill_1 FILLER_14_397 ();
 sg13g2_fill_2 FILLER_14_437 ();
 sg13g2_fill_1 FILLER_14_439 ();
 sg13g2_fill_2 FILLER_14_469 ();
 sg13g2_fill_1 FILLER_14_471 ();
 sg13g2_decap_8 FILLER_14_482 ();
 sg13g2_fill_2 FILLER_14_489 ();
 sg13g2_fill_1 FILLER_14_491 ();
 sg13g2_fill_1 FILLER_14_496 ();
 sg13g2_fill_1 FILLER_14_506 ();
 sg13g2_decap_8 FILLER_14_520 ();
 sg13g2_decap_4 FILLER_14_531 ();
 sg13g2_fill_2 FILLER_14_540 ();
 sg13g2_decap_4 FILLER_14_546 ();
 sg13g2_fill_1 FILLER_14_550 ();
 sg13g2_fill_2 FILLER_14_585 ();
 sg13g2_fill_1 FILLER_14_587 ();
 sg13g2_fill_2 FILLER_14_623 ();
 sg13g2_fill_1 FILLER_14_651 ();
 sg13g2_fill_1 FILLER_14_675 ();
 sg13g2_fill_1 FILLER_14_721 ();
 sg13g2_fill_2 FILLER_14_757 ();
 sg13g2_fill_2 FILLER_14_771 ();
 sg13g2_fill_1 FILLER_14_782 ();
 sg13g2_fill_1 FILLER_14_793 ();
 sg13g2_fill_2 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_832 ();
 sg13g2_decap_8 FILLER_14_839 ();
 sg13g2_decap_8 FILLER_14_846 ();
 sg13g2_decap_4 FILLER_14_853 ();
 sg13g2_fill_1 FILLER_14_857 ();
 sg13g2_fill_2 FILLER_14_913 ();
 sg13g2_fill_1 FILLER_14_953 ();
 sg13g2_fill_2 FILLER_14_963 ();
 sg13g2_fill_2 FILLER_14_1063 ();
 sg13g2_fill_1 FILLER_14_1099 ();
 sg13g2_fill_2 FILLER_14_1201 ();
 sg13g2_fill_2 FILLER_14_1233 ();
 sg13g2_fill_2 FILLER_14_1253 ();
 sg13g2_fill_2 FILLER_14_1311 ();
 sg13g2_fill_1 FILLER_14_1521 ();
 sg13g2_fill_1 FILLER_14_1534 ();
 sg13g2_fill_2 FILLER_14_1618 ();
 sg13g2_fill_2 FILLER_14_1676 ();
 sg13g2_fill_2 FILLER_14_1727 ();
 sg13g2_fill_1 FILLER_14_1737 ();
 sg13g2_fill_2 FILLER_14_1820 ();
 sg13g2_fill_1 FILLER_14_1822 ();
 sg13g2_fill_2 FILLER_14_1833 ();
 sg13g2_fill_1 FILLER_14_1835 ();
 sg13g2_decap_8 FILLER_14_1903 ();
 sg13g2_fill_2 FILLER_14_1928 ();
 sg13g2_fill_1 FILLER_14_1935 ();
 sg13g2_fill_2 FILLER_14_1977 ();
 sg13g2_decap_4 FILLER_14_1983 ();
 sg13g2_fill_2 FILLER_14_1987 ();
 sg13g2_fill_1 FILLER_14_2003 ();
 sg13g2_fill_1 FILLER_14_2008 ();
 sg13g2_decap_8 FILLER_14_2019 ();
 sg13g2_fill_2 FILLER_14_2067 ();
 sg13g2_fill_2 FILLER_14_2113 ();
 sg13g2_fill_1 FILLER_14_2174 ();
 sg13g2_fill_1 FILLER_14_2189 ();
 sg13g2_fill_2 FILLER_14_2246 ();
 sg13g2_fill_1 FILLER_14_2248 ();
 sg13g2_fill_1 FILLER_14_2253 ();
 sg13g2_decap_4 FILLER_14_2309 ();
 sg13g2_decap_4 FILLER_14_2328 ();
 sg13g2_decap_8 FILLER_14_2345 ();
 sg13g2_decap_8 FILLER_14_2352 ();
 sg13g2_decap_8 FILLER_14_2359 ();
 sg13g2_decap_8 FILLER_14_2366 ();
 sg13g2_decap_8 FILLER_14_2373 ();
 sg13g2_decap_8 FILLER_14_2380 ();
 sg13g2_decap_8 FILLER_14_2387 ();
 sg13g2_decap_8 FILLER_14_2394 ();
 sg13g2_decap_8 FILLER_14_2401 ();
 sg13g2_decap_8 FILLER_14_2408 ();
 sg13g2_decap_8 FILLER_14_2415 ();
 sg13g2_decap_8 FILLER_14_2422 ();
 sg13g2_decap_8 FILLER_14_2429 ();
 sg13g2_decap_8 FILLER_14_2436 ();
 sg13g2_decap_8 FILLER_14_2443 ();
 sg13g2_decap_8 FILLER_14_2450 ();
 sg13g2_decap_8 FILLER_14_2457 ();
 sg13g2_decap_8 FILLER_14_2464 ();
 sg13g2_decap_8 FILLER_14_2471 ();
 sg13g2_decap_8 FILLER_14_2478 ();
 sg13g2_decap_8 FILLER_14_2485 ();
 sg13g2_decap_8 FILLER_14_2492 ();
 sg13g2_decap_8 FILLER_14_2499 ();
 sg13g2_decap_8 FILLER_14_2506 ();
 sg13g2_decap_8 FILLER_14_2513 ();
 sg13g2_decap_8 FILLER_14_2520 ();
 sg13g2_decap_8 FILLER_14_2527 ();
 sg13g2_decap_8 FILLER_14_2534 ();
 sg13g2_decap_8 FILLER_14_2541 ();
 sg13g2_decap_8 FILLER_14_2548 ();
 sg13g2_decap_8 FILLER_14_2555 ();
 sg13g2_decap_8 FILLER_14_2562 ();
 sg13g2_decap_8 FILLER_14_2569 ();
 sg13g2_decap_8 FILLER_14_2576 ();
 sg13g2_decap_8 FILLER_14_2583 ();
 sg13g2_decap_8 FILLER_14_2590 ();
 sg13g2_decap_8 FILLER_14_2597 ();
 sg13g2_decap_8 FILLER_14_2604 ();
 sg13g2_decap_8 FILLER_14_2611 ();
 sg13g2_decap_8 FILLER_14_2618 ();
 sg13g2_decap_8 FILLER_14_2625 ();
 sg13g2_decap_8 FILLER_14_2632 ();
 sg13g2_decap_8 FILLER_14_2639 ();
 sg13g2_decap_8 FILLER_14_2646 ();
 sg13g2_decap_8 FILLER_14_2653 ();
 sg13g2_decap_8 FILLER_14_2660 ();
 sg13g2_decap_8 FILLER_14_2667 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_fill_1 FILLER_15_147 ();
 sg13g2_decap_4 FILLER_15_152 ();
 sg13g2_fill_1 FILLER_15_156 ();
 sg13g2_fill_2 FILLER_15_188 ();
 sg13g2_fill_1 FILLER_15_190 ();
 sg13g2_decap_4 FILLER_15_196 ();
 sg13g2_fill_1 FILLER_15_200 ();
 sg13g2_decap_8 FILLER_15_206 ();
 sg13g2_fill_2 FILLER_15_213 ();
 sg13g2_fill_1 FILLER_15_215 ();
 sg13g2_fill_1 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_253 ();
 sg13g2_fill_1 FILLER_15_260 ();
 sg13g2_fill_1 FILLER_15_274 ();
 sg13g2_fill_2 FILLER_15_288 ();
 sg13g2_fill_1 FILLER_15_290 ();
 sg13g2_fill_2 FILLER_15_301 ();
 sg13g2_fill_2 FILLER_15_311 ();
 sg13g2_fill_1 FILLER_15_358 ();
 sg13g2_fill_2 FILLER_15_394 ();
 sg13g2_fill_2 FILLER_15_416 ();
 sg13g2_fill_2 FILLER_15_432 ();
 sg13g2_fill_1 FILLER_15_434 ();
 sg13g2_fill_1 FILLER_15_449 ();
 sg13g2_fill_2 FILLER_15_516 ();
 sg13g2_fill_1 FILLER_15_518 ();
 sg13g2_fill_1 FILLER_15_541 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_4 FILLER_15_553 ();
 sg13g2_fill_1 FILLER_15_569 ();
 sg13g2_fill_2 FILLER_15_583 ();
 sg13g2_fill_2 FILLER_15_619 ();
 sg13g2_fill_2 FILLER_15_632 ();
 sg13g2_fill_1 FILLER_15_634 ();
 sg13g2_fill_2 FILLER_15_657 ();
 sg13g2_fill_2 FILLER_15_687 ();
 sg13g2_fill_2 FILLER_15_710 ();
 sg13g2_fill_2 FILLER_15_741 ();
 sg13g2_fill_1 FILLER_15_743 ();
 sg13g2_decap_4 FILLER_15_764 ();
 sg13g2_fill_2 FILLER_15_793 ();
 sg13g2_decap_8 FILLER_15_836 ();
 sg13g2_decap_8 FILLER_15_843 ();
 sg13g2_decap_8 FILLER_15_850 ();
 sg13g2_fill_2 FILLER_15_857 ();
 sg13g2_fill_2 FILLER_15_907 ();
 sg13g2_fill_2 FILLER_15_918 ();
 sg13g2_fill_2 FILLER_15_929 ();
 sg13g2_fill_1 FILLER_15_998 ();
 sg13g2_fill_2 FILLER_15_1140 ();
 sg13g2_fill_2 FILLER_15_1341 ();
 sg13g2_fill_2 FILLER_15_1352 ();
 sg13g2_fill_2 FILLER_15_1459 ();
 sg13g2_fill_1 FILLER_15_1487 ();
 sg13g2_fill_1 FILLER_15_1527 ();
 sg13g2_fill_1 FILLER_15_1537 ();
 sg13g2_fill_1 FILLER_15_1657 ();
 sg13g2_fill_2 FILLER_15_1667 ();
 sg13g2_fill_1 FILLER_15_1747 ();
 sg13g2_fill_2 FILLER_15_1771 ();
 sg13g2_fill_1 FILLER_15_1773 ();
 sg13g2_fill_1 FILLER_15_1783 ();
 sg13g2_fill_2 FILLER_15_1812 ();
 sg13g2_fill_1 FILLER_15_1855 ();
 sg13g2_fill_2 FILLER_15_1895 ();
 sg13g2_decap_8 FILLER_15_1920 ();
 sg13g2_decap_4 FILLER_15_1927 ();
 sg13g2_fill_1 FILLER_15_1939 ();
 sg13g2_fill_2 FILLER_15_1966 ();
 sg13g2_fill_1 FILLER_15_1968 ();
 sg13g2_fill_2 FILLER_15_1973 ();
 sg13g2_decap_4 FILLER_15_1979 ();
 sg13g2_fill_2 FILLER_15_2010 ();
 sg13g2_fill_1 FILLER_15_2073 ();
 sg13g2_fill_1 FILLER_15_2134 ();
 sg13g2_fill_1 FILLER_15_2148 ();
 sg13g2_fill_2 FILLER_15_2228 ();
 sg13g2_fill_1 FILLER_15_2230 ();
 sg13g2_decap_8 FILLER_15_2252 ();
 sg13g2_decap_8 FILLER_15_2259 ();
 sg13g2_decap_4 FILLER_15_2266 ();
 sg13g2_fill_2 FILLER_15_2270 ();
 sg13g2_fill_1 FILLER_15_2277 ();
 sg13g2_fill_1 FILLER_15_2320 ();
 sg13g2_decap_8 FILLER_15_2347 ();
 sg13g2_decap_8 FILLER_15_2354 ();
 sg13g2_decap_8 FILLER_15_2361 ();
 sg13g2_decap_8 FILLER_15_2368 ();
 sg13g2_decap_8 FILLER_15_2375 ();
 sg13g2_decap_8 FILLER_15_2382 ();
 sg13g2_decap_8 FILLER_15_2389 ();
 sg13g2_decap_8 FILLER_15_2396 ();
 sg13g2_decap_8 FILLER_15_2403 ();
 sg13g2_decap_8 FILLER_15_2410 ();
 sg13g2_decap_8 FILLER_15_2417 ();
 sg13g2_decap_8 FILLER_15_2424 ();
 sg13g2_decap_8 FILLER_15_2431 ();
 sg13g2_decap_8 FILLER_15_2438 ();
 sg13g2_decap_8 FILLER_15_2445 ();
 sg13g2_decap_8 FILLER_15_2452 ();
 sg13g2_decap_8 FILLER_15_2459 ();
 sg13g2_decap_8 FILLER_15_2466 ();
 sg13g2_decap_8 FILLER_15_2473 ();
 sg13g2_decap_8 FILLER_15_2480 ();
 sg13g2_decap_8 FILLER_15_2487 ();
 sg13g2_decap_8 FILLER_15_2494 ();
 sg13g2_decap_8 FILLER_15_2501 ();
 sg13g2_decap_8 FILLER_15_2508 ();
 sg13g2_decap_8 FILLER_15_2515 ();
 sg13g2_decap_8 FILLER_15_2522 ();
 sg13g2_decap_8 FILLER_15_2529 ();
 sg13g2_decap_8 FILLER_15_2536 ();
 sg13g2_decap_8 FILLER_15_2543 ();
 sg13g2_decap_8 FILLER_15_2550 ();
 sg13g2_decap_8 FILLER_15_2557 ();
 sg13g2_decap_8 FILLER_15_2564 ();
 sg13g2_decap_8 FILLER_15_2571 ();
 sg13g2_decap_8 FILLER_15_2578 ();
 sg13g2_decap_8 FILLER_15_2585 ();
 sg13g2_decap_8 FILLER_15_2592 ();
 sg13g2_decap_8 FILLER_15_2599 ();
 sg13g2_decap_8 FILLER_15_2606 ();
 sg13g2_decap_8 FILLER_15_2613 ();
 sg13g2_decap_8 FILLER_15_2620 ();
 sg13g2_decap_8 FILLER_15_2627 ();
 sg13g2_decap_8 FILLER_15_2634 ();
 sg13g2_decap_8 FILLER_15_2641 ();
 sg13g2_decap_8 FILLER_15_2648 ();
 sg13g2_decap_8 FILLER_15_2655 ();
 sg13g2_decap_8 FILLER_15_2662 ();
 sg13g2_decap_4 FILLER_15_2669 ();
 sg13g2_fill_1 FILLER_15_2673 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_fill_1 FILLER_16_163 ();
 sg13g2_fill_1 FILLER_16_182 ();
 sg13g2_fill_2 FILLER_16_198 ();
 sg13g2_fill_2 FILLER_16_213 ();
 sg13g2_decap_4 FILLER_16_233 ();
 sg13g2_fill_2 FILLER_16_253 ();
 sg13g2_fill_1 FILLER_16_255 ();
 sg13g2_fill_2 FILLER_16_271 ();
 sg13g2_fill_2 FILLER_16_352 ();
 sg13g2_fill_1 FILLER_16_376 ();
 sg13g2_fill_2 FILLER_16_421 ();
 sg13g2_fill_1 FILLER_16_423 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_fill_2 FILLER_16_439 ();
 sg13g2_fill_1 FILLER_16_441 ();
 sg13g2_fill_2 FILLER_16_463 ();
 sg13g2_fill_1 FILLER_16_530 ();
 sg13g2_decap_4 FILLER_16_557 ();
 sg13g2_fill_2 FILLER_16_561 ();
 sg13g2_fill_2 FILLER_16_577 ();
 sg13g2_fill_1 FILLER_16_579 ();
 sg13g2_fill_2 FILLER_16_606 ();
 sg13g2_fill_1 FILLER_16_608 ();
 sg13g2_fill_1 FILLER_16_652 ();
 sg13g2_fill_1 FILLER_16_713 ();
 sg13g2_fill_1 FILLER_16_749 ();
 sg13g2_decap_4 FILLER_16_762 ();
 sg13g2_fill_2 FILLER_16_766 ();
 sg13g2_fill_1 FILLER_16_789 ();
 sg13g2_decap_8 FILLER_16_810 ();
 sg13g2_decap_4 FILLER_16_817 ();
 sg13g2_fill_1 FILLER_16_821 ();
 sg13g2_decap_8 FILLER_16_843 ();
 sg13g2_decap_8 FILLER_16_850 ();
 sg13g2_fill_1 FILLER_16_857 ();
 sg13g2_fill_1 FILLER_16_968 ();
 sg13g2_fill_2 FILLER_16_998 ();
 sg13g2_fill_1 FILLER_16_1049 ();
 sg13g2_fill_1 FILLER_16_1157 ();
 sg13g2_fill_1 FILLER_16_1199 ();
 sg13g2_fill_2 FILLER_16_1209 ();
 sg13g2_fill_1 FILLER_16_1309 ();
 sg13g2_fill_2 FILLER_16_1350 ();
 sg13g2_fill_1 FILLER_16_1423 ();
 sg13g2_fill_2 FILLER_16_1508 ();
 sg13g2_fill_1 FILLER_16_1652 ();
 sg13g2_fill_2 FILLER_16_1708 ();
 sg13g2_fill_1 FILLER_16_1724 ();
 sg13g2_fill_2 FILLER_16_1730 ();
 sg13g2_fill_2 FILLER_16_1809 ();
 sg13g2_fill_1 FILLER_16_1811 ();
 sg13g2_fill_2 FILLER_16_1879 ();
 sg13g2_fill_2 FILLER_16_1923 ();
 sg13g2_fill_1 FILLER_16_1925 ();
 sg13g2_fill_2 FILLER_16_1934 ();
 sg13g2_fill_1 FILLER_16_1936 ();
 sg13g2_fill_2 FILLER_16_2018 ();
 sg13g2_fill_1 FILLER_16_2020 ();
 sg13g2_fill_2 FILLER_16_2034 ();
 sg13g2_fill_1 FILLER_16_2036 ();
 sg13g2_fill_2 FILLER_16_2092 ();
 sg13g2_decap_4 FILLER_16_2154 ();
 sg13g2_decap_8 FILLER_16_2202 ();
 sg13g2_fill_2 FILLER_16_2209 ();
 sg13g2_fill_1 FILLER_16_2211 ();
 sg13g2_fill_1 FILLER_16_2288 ();
 sg13g2_decap_8 FILLER_16_2353 ();
 sg13g2_decap_8 FILLER_16_2360 ();
 sg13g2_decap_8 FILLER_16_2367 ();
 sg13g2_decap_8 FILLER_16_2374 ();
 sg13g2_decap_8 FILLER_16_2381 ();
 sg13g2_decap_8 FILLER_16_2388 ();
 sg13g2_decap_8 FILLER_16_2395 ();
 sg13g2_decap_8 FILLER_16_2402 ();
 sg13g2_decap_8 FILLER_16_2409 ();
 sg13g2_decap_8 FILLER_16_2416 ();
 sg13g2_decap_8 FILLER_16_2423 ();
 sg13g2_decap_8 FILLER_16_2430 ();
 sg13g2_decap_8 FILLER_16_2437 ();
 sg13g2_decap_8 FILLER_16_2444 ();
 sg13g2_decap_8 FILLER_16_2451 ();
 sg13g2_decap_8 FILLER_16_2458 ();
 sg13g2_decap_8 FILLER_16_2465 ();
 sg13g2_decap_8 FILLER_16_2472 ();
 sg13g2_decap_8 FILLER_16_2479 ();
 sg13g2_decap_8 FILLER_16_2486 ();
 sg13g2_decap_8 FILLER_16_2493 ();
 sg13g2_decap_8 FILLER_16_2500 ();
 sg13g2_decap_8 FILLER_16_2507 ();
 sg13g2_decap_8 FILLER_16_2514 ();
 sg13g2_decap_8 FILLER_16_2521 ();
 sg13g2_decap_8 FILLER_16_2528 ();
 sg13g2_decap_8 FILLER_16_2535 ();
 sg13g2_decap_8 FILLER_16_2542 ();
 sg13g2_decap_8 FILLER_16_2549 ();
 sg13g2_decap_8 FILLER_16_2556 ();
 sg13g2_decap_8 FILLER_16_2563 ();
 sg13g2_decap_8 FILLER_16_2570 ();
 sg13g2_decap_8 FILLER_16_2577 ();
 sg13g2_decap_8 FILLER_16_2584 ();
 sg13g2_decap_8 FILLER_16_2591 ();
 sg13g2_decap_8 FILLER_16_2598 ();
 sg13g2_decap_8 FILLER_16_2605 ();
 sg13g2_decap_8 FILLER_16_2612 ();
 sg13g2_decap_8 FILLER_16_2619 ();
 sg13g2_decap_8 FILLER_16_2626 ();
 sg13g2_decap_8 FILLER_16_2633 ();
 sg13g2_decap_8 FILLER_16_2640 ();
 sg13g2_decap_8 FILLER_16_2647 ();
 sg13g2_decap_8 FILLER_16_2654 ();
 sg13g2_decap_8 FILLER_16_2661 ();
 sg13g2_decap_4 FILLER_16_2668 ();
 sg13g2_fill_2 FILLER_16_2672 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_4 FILLER_17_119 ();
 sg13g2_fill_2 FILLER_17_162 ();
 sg13g2_fill_1 FILLER_17_164 ();
 sg13g2_fill_1 FILLER_17_173 ();
 sg13g2_decap_4 FILLER_17_179 ();
 sg13g2_fill_1 FILLER_17_183 ();
 sg13g2_fill_2 FILLER_17_198 ();
 sg13g2_fill_1 FILLER_17_200 ();
 sg13g2_decap_8 FILLER_17_228 ();
 sg13g2_decap_4 FILLER_17_235 ();
 sg13g2_fill_2 FILLER_17_239 ();
 sg13g2_fill_1 FILLER_17_249 ();
 sg13g2_fill_2 FILLER_17_260 ();
 sg13g2_fill_1 FILLER_17_262 ();
 sg13g2_fill_1 FILLER_17_285 ();
 sg13g2_fill_2 FILLER_17_365 ();
 sg13g2_fill_1 FILLER_17_367 ();
 sg13g2_fill_1 FILLER_17_376 ();
 sg13g2_fill_2 FILLER_17_385 ();
 sg13g2_fill_1 FILLER_17_387 ();
 sg13g2_fill_2 FILLER_17_397 ();
 sg13g2_fill_2 FILLER_17_467 ();
 sg13g2_fill_2 FILLER_17_486 ();
 sg13g2_fill_1 FILLER_17_488 ();
 sg13g2_fill_1 FILLER_17_498 ();
 sg13g2_fill_1 FILLER_17_507 ();
 sg13g2_fill_2 FILLER_17_513 ();
 sg13g2_decap_8 FILLER_17_531 ();
 sg13g2_decap_4 FILLER_17_538 ();
 sg13g2_fill_2 FILLER_17_542 ();
 sg13g2_decap_8 FILLER_17_548 ();
 sg13g2_fill_1 FILLER_17_596 ();
 sg13g2_fill_2 FILLER_17_626 ();
 sg13g2_fill_2 FILLER_17_664 ();
 sg13g2_fill_1 FILLER_17_666 ();
 sg13g2_fill_1 FILLER_17_686 ();
 sg13g2_decap_4 FILLER_17_753 ();
 sg13g2_fill_2 FILLER_17_757 ();
 sg13g2_decap_4 FILLER_17_784 ();
 sg13g2_fill_2 FILLER_17_788 ();
 sg13g2_decap_8 FILLER_17_809 ();
 sg13g2_decap_8 FILLER_17_816 ();
 sg13g2_fill_2 FILLER_17_823 ();
 sg13g2_fill_1 FILLER_17_825 ();
 sg13g2_fill_2 FILLER_17_838 ();
 sg13g2_decap_8 FILLER_17_848 ();
 sg13g2_fill_1 FILLER_17_863 ();
 sg13g2_fill_1 FILLER_17_874 ();
 sg13g2_fill_2 FILLER_17_879 ();
 sg13g2_fill_2 FILLER_17_1081 ();
 sg13g2_fill_2 FILLER_17_1177 ();
 sg13g2_fill_2 FILLER_17_1363 ();
 sg13g2_fill_2 FILLER_17_1403 ();
 sg13g2_fill_2 FILLER_17_1450 ();
 sg13g2_fill_1 FILLER_17_1509 ();
 sg13g2_fill_1 FILLER_17_1524 ();
 sg13g2_fill_1 FILLER_17_1559 ();
 sg13g2_fill_2 FILLER_17_1602 ();
 sg13g2_fill_2 FILLER_17_1627 ();
 sg13g2_fill_2 FILLER_17_1733 ();
 sg13g2_fill_2 FILLER_17_1750 ();
 sg13g2_fill_1 FILLER_17_1765 ();
 sg13g2_fill_1 FILLER_17_1780 ();
 sg13g2_fill_2 FILLER_17_1794 ();
 sg13g2_fill_1 FILLER_17_1806 ();
 sg13g2_fill_1 FILLER_17_1858 ();
 sg13g2_fill_1 FILLER_17_1893 ();
 sg13g2_fill_2 FILLER_17_1912 ();
 sg13g2_fill_2 FILLER_17_1925 ();
 sg13g2_fill_1 FILLER_17_1950 ();
 sg13g2_fill_2 FILLER_17_1960 ();
 sg13g2_fill_2 FILLER_17_1970 ();
 sg13g2_fill_1 FILLER_17_1972 ();
 sg13g2_fill_1 FILLER_17_1992 ();
 sg13g2_fill_2 FILLER_17_2002 ();
 sg13g2_fill_1 FILLER_17_2004 ();
 sg13g2_decap_8 FILLER_17_2041 ();
 sg13g2_decap_8 FILLER_17_2048 ();
 sg13g2_fill_1 FILLER_17_2055 ();
 sg13g2_decap_8 FILLER_17_2070 ();
 sg13g2_fill_2 FILLER_17_2077 ();
 sg13g2_fill_1 FILLER_17_2089 ();
 sg13g2_fill_2 FILLER_17_2108 ();
 sg13g2_fill_1 FILLER_17_2110 ();
 sg13g2_decap_4 FILLER_17_2134 ();
 sg13g2_fill_1 FILLER_17_2138 ();
 sg13g2_decap_8 FILLER_17_2147 ();
 sg13g2_fill_2 FILLER_17_2180 ();
 sg13g2_fill_1 FILLER_17_2182 ();
 sg13g2_fill_2 FILLER_17_2237 ();
 sg13g2_decap_8 FILLER_17_2261 ();
 sg13g2_fill_1 FILLER_17_2283 ();
 sg13g2_fill_1 FILLER_17_2289 ();
 sg13g2_decap_8 FILLER_17_2328 ();
 sg13g2_fill_2 FILLER_17_2335 ();
 sg13g2_decap_8 FILLER_17_2350 ();
 sg13g2_decap_8 FILLER_17_2357 ();
 sg13g2_decap_8 FILLER_17_2364 ();
 sg13g2_decap_8 FILLER_17_2371 ();
 sg13g2_decap_8 FILLER_17_2378 ();
 sg13g2_decap_8 FILLER_17_2385 ();
 sg13g2_decap_8 FILLER_17_2392 ();
 sg13g2_decap_8 FILLER_17_2399 ();
 sg13g2_decap_8 FILLER_17_2406 ();
 sg13g2_decap_8 FILLER_17_2413 ();
 sg13g2_decap_8 FILLER_17_2420 ();
 sg13g2_decap_8 FILLER_17_2427 ();
 sg13g2_decap_8 FILLER_17_2434 ();
 sg13g2_decap_8 FILLER_17_2441 ();
 sg13g2_decap_8 FILLER_17_2448 ();
 sg13g2_decap_8 FILLER_17_2455 ();
 sg13g2_decap_8 FILLER_17_2462 ();
 sg13g2_decap_8 FILLER_17_2469 ();
 sg13g2_decap_8 FILLER_17_2476 ();
 sg13g2_decap_8 FILLER_17_2483 ();
 sg13g2_decap_8 FILLER_17_2490 ();
 sg13g2_decap_8 FILLER_17_2497 ();
 sg13g2_decap_8 FILLER_17_2504 ();
 sg13g2_decap_8 FILLER_17_2511 ();
 sg13g2_decap_8 FILLER_17_2518 ();
 sg13g2_decap_8 FILLER_17_2525 ();
 sg13g2_decap_8 FILLER_17_2532 ();
 sg13g2_decap_8 FILLER_17_2539 ();
 sg13g2_decap_8 FILLER_17_2546 ();
 sg13g2_decap_8 FILLER_17_2553 ();
 sg13g2_decap_8 FILLER_17_2560 ();
 sg13g2_decap_8 FILLER_17_2567 ();
 sg13g2_decap_8 FILLER_17_2574 ();
 sg13g2_decap_8 FILLER_17_2581 ();
 sg13g2_decap_8 FILLER_17_2588 ();
 sg13g2_decap_8 FILLER_17_2595 ();
 sg13g2_decap_8 FILLER_17_2602 ();
 sg13g2_decap_8 FILLER_17_2609 ();
 sg13g2_decap_8 FILLER_17_2616 ();
 sg13g2_decap_8 FILLER_17_2623 ();
 sg13g2_decap_8 FILLER_17_2630 ();
 sg13g2_decap_8 FILLER_17_2637 ();
 sg13g2_decap_8 FILLER_17_2644 ();
 sg13g2_decap_8 FILLER_17_2651 ();
 sg13g2_decap_8 FILLER_17_2658 ();
 sg13g2_decap_8 FILLER_17_2665 ();
 sg13g2_fill_2 FILLER_17_2672 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_4 FILLER_18_126 ();
 sg13g2_fill_1 FILLER_18_130 ();
 sg13g2_fill_2 FILLER_18_162 ();
 sg13g2_decap_8 FILLER_18_174 ();
 sg13g2_decap_4 FILLER_18_181 ();
 sg13g2_fill_1 FILLER_18_217 ();
 sg13g2_decap_4 FILLER_18_228 ();
 sg13g2_fill_2 FILLER_18_244 ();
 sg13g2_fill_2 FILLER_18_260 ();
 sg13g2_fill_2 FILLER_18_282 ();
 sg13g2_fill_1 FILLER_18_284 ();
 sg13g2_fill_2 FILLER_18_293 ();
 sg13g2_decap_4 FILLER_18_304 ();
 sg13g2_fill_1 FILLER_18_308 ();
 sg13g2_decap_4 FILLER_18_313 ();
 sg13g2_fill_1 FILLER_18_317 ();
 sg13g2_fill_1 FILLER_18_355 ();
 sg13g2_fill_2 FILLER_18_370 ();
 sg13g2_fill_2 FILLER_18_386 ();
 sg13g2_fill_1 FILLER_18_388 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_fill_1 FILLER_18_409 ();
 sg13g2_fill_1 FILLER_18_436 ();
 sg13g2_fill_1 FILLER_18_440 ();
 sg13g2_fill_2 FILLER_18_505 ();
 sg13g2_fill_2 FILLER_18_635 ();
 sg13g2_fill_1 FILLER_18_647 ();
 sg13g2_fill_1 FILLER_18_659 ();
 sg13g2_fill_2 FILLER_18_702 ();
 sg13g2_fill_1 FILLER_18_713 ();
 sg13g2_fill_1 FILLER_18_733 ();
 sg13g2_fill_2 FILLER_18_764 ();
 sg13g2_fill_1 FILLER_18_766 ();
 sg13g2_fill_1 FILLER_18_792 ();
 sg13g2_fill_1 FILLER_18_809 ();
 sg13g2_decap_4 FILLER_18_823 ();
 sg13g2_fill_1 FILLER_18_840 ();
 sg13g2_decap_4 FILLER_18_864 ();
 sg13g2_fill_2 FILLER_18_876 ();
 sg13g2_fill_1 FILLER_18_878 ();
 sg13g2_fill_1 FILLER_18_1036 ();
 sg13g2_fill_2 FILLER_18_1043 ();
 sg13g2_fill_1 FILLER_18_1068 ();
 sg13g2_fill_2 FILLER_18_1083 ();
 sg13g2_fill_1 FILLER_18_1130 ();
 sg13g2_fill_2 FILLER_18_1284 ();
 sg13g2_fill_1 FILLER_18_1295 ();
 sg13g2_fill_2 FILLER_18_1349 ();
 sg13g2_fill_1 FILLER_18_1591 ();
 sg13g2_fill_2 FILLER_18_1627 ();
 sg13g2_fill_1 FILLER_18_1690 ();
 sg13g2_fill_1 FILLER_18_1727 ();
 sg13g2_fill_2 FILLER_18_1759 ();
 sg13g2_fill_2 FILLER_18_1805 ();
 sg13g2_fill_1 FILLER_18_1807 ();
 sg13g2_fill_1 FILLER_18_1823 ();
 sg13g2_fill_2 FILLER_18_1838 ();
 sg13g2_fill_1 FILLER_18_1853 ();
 sg13g2_fill_1 FILLER_18_1859 ();
 sg13g2_decap_4 FILLER_18_1864 ();
 sg13g2_fill_2 FILLER_18_1868 ();
 sg13g2_fill_2 FILLER_18_1874 ();
 sg13g2_fill_1 FILLER_18_1876 ();
 sg13g2_fill_1 FILLER_18_1882 ();
 sg13g2_fill_1 FILLER_18_1950 ();
 sg13g2_fill_1 FILLER_18_2027 ();
 sg13g2_fill_2 FILLER_18_2116 ();
 sg13g2_fill_2 FILLER_18_2176 ();
 sg13g2_fill_1 FILLER_18_2289 ();
 sg13g2_decap_8 FILLER_18_2342 ();
 sg13g2_decap_8 FILLER_18_2349 ();
 sg13g2_decap_8 FILLER_18_2356 ();
 sg13g2_decap_8 FILLER_18_2363 ();
 sg13g2_decap_8 FILLER_18_2370 ();
 sg13g2_decap_8 FILLER_18_2377 ();
 sg13g2_decap_8 FILLER_18_2384 ();
 sg13g2_decap_8 FILLER_18_2391 ();
 sg13g2_decap_8 FILLER_18_2398 ();
 sg13g2_decap_8 FILLER_18_2405 ();
 sg13g2_decap_8 FILLER_18_2412 ();
 sg13g2_decap_8 FILLER_18_2419 ();
 sg13g2_decap_8 FILLER_18_2426 ();
 sg13g2_decap_8 FILLER_18_2433 ();
 sg13g2_decap_8 FILLER_18_2440 ();
 sg13g2_decap_8 FILLER_18_2447 ();
 sg13g2_decap_8 FILLER_18_2454 ();
 sg13g2_decap_8 FILLER_18_2461 ();
 sg13g2_decap_8 FILLER_18_2468 ();
 sg13g2_decap_8 FILLER_18_2475 ();
 sg13g2_decap_8 FILLER_18_2482 ();
 sg13g2_decap_8 FILLER_18_2489 ();
 sg13g2_decap_8 FILLER_18_2496 ();
 sg13g2_decap_8 FILLER_18_2503 ();
 sg13g2_decap_8 FILLER_18_2510 ();
 sg13g2_decap_8 FILLER_18_2517 ();
 sg13g2_decap_8 FILLER_18_2524 ();
 sg13g2_decap_8 FILLER_18_2531 ();
 sg13g2_decap_8 FILLER_18_2538 ();
 sg13g2_decap_8 FILLER_18_2545 ();
 sg13g2_decap_8 FILLER_18_2552 ();
 sg13g2_decap_8 FILLER_18_2559 ();
 sg13g2_decap_8 FILLER_18_2566 ();
 sg13g2_decap_8 FILLER_18_2573 ();
 sg13g2_decap_8 FILLER_18_2580 ();
 sg13g2_decap_8 FILLER_18_2587 ();
 sg13g2_decap_8 FILLER_18_2594 ();
 sg13g2_decap_8 FILLER_18_2601 ();
 sg13g2_decap_8 FILLER_18_2608 ();
 sg13g2_decap_8 FILLER_18_2615 ();
 sg13g2_decap_8 FILLER_18_2622 ();
 sg13g2_decap_8 FILLER_18_2629 ();
 sg13g2_decap_8 FILLER_18_2636 ();
 sg13g2_decap_8 FILLER_18_2643 ();
 sg13g2_decap_8 FILLER_18_2650 ();
 sg13g2_decap_8 FILLER_18_2657 ();
 sg13g2_decap_8 FILLER_18_2664 ();
 sg13g2_fill_2 FILLER_18_2671 ();
 sg13g2_fill_1 FILLER_18_2673 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_4 FILLER_19_105 ();
 sg13g2_fill_2 FILLER_19_162 ();
 sg13g2_fill_1 FILLER_19_164 ();
 sg13g2_fill_2 FILLER_19_256 ();
 sg13g2_fill_2 FILLER_19_281 ();
 sg13g2_fill_1 FILLER_19_283 ();
 sg13g2_decap_8 FILLER_19_293 ();
 sg13g2_fill_1 FILLER_19_300 ();
 sg13g2_fill_1 FILLER_19_383 ();
 sg13g2_fill_2 FILLER_19_418 ();
 sg13g2_fill_2 FILLER_19_445 ();
 sg13g2_decap_4 FILLER_19_478 ();
 sg13g2_fill_1 FILLER_19_490 ();
 sg13g2_fill_2 FILLER_19_520 ();
 sg13g2_fill_1 FILLER_19_526 ();
 sg13g2_fill_2 FILLER_19_544 ();
 sg13g2_fill_1 FILLER_19_624 ();
 sg13g2_fill_2 FILLER_19_651 ();
 sg13g2_fill_2 FILLER_19_735 ();
 sg13g2_fill_1 FILLER_19_737 ();
 sg13g2_decap_8 FILLER_19_773 ();
 sg13g2_fill_2 FILLER_19_797 ();
 sg13g2_fill_1 FILLER_19_799 ();
 sg13g2_fill_1 FILLER_19_809 ();
 sg13g2_decap_4 FILLER_19_831 ();
 sg13g2_fill_2 FILLER_19_843 ();
 sg13g2_fill_1 FILLER_19_848 ();
 sg13g2_fill_1 FILLER_19_1143 ();
 sg13g2_fill_1 FILLER_19_1263 ();
 sg13g2_fill_2 FILLER_19_1330 ();
 sg13g2_fill_2 FILLER_19_1371 ();
 sg13g2_fill_2 FILLER_19_1422 ();
 sg13g2_fill_1 FILLER_19_1505 ();
 sg13g2_fill_1 FILLER_19_1580 ();
 sg13g2_fill_1 FILLER_19_1648 ();
 sg13g2_fill_2 FILLER_19_1658 ();
 sg13g2_fill_1 FILLER_19_1674 ();
 sg13g2_fill_2 FILLER_19_1696 ();
 sg13g2_fill_1 FILLER_19_1778 ();
 sg13g2_fill_2 FILLER_19_1788 ();
 sg13g2_fill_1 FILLER_19_1790 ();
 sg13g2_decap_8 FILLER_19_1817 ();
 sg13g2_fill_2 FILLER_19_1824 ();
 sg13g2_fill_2 FILLER_19_1888 ();
 sg13g2_fill_2 FILLER_19_1918 ();
 sg13g2_fill_1 FILLER_19_1920 ();
 sg13g2_fill_2 FILLER_19_1961 ();
 sg13g2_fill_1 FILLER_19_1963 ();
 sg13g2_decap_4 FILLER_19_2009 ();
 sg13g2_fill_1 FILLER_19_2013 ();
 sg13g2_decap_4 FILLER_19_2044 ();
 sg13g2_fill_1 FILLER_19_2074 ();
 sg13g2_fill_2 FILLER_19_2093 ();
 sg13g2_fill_1 FILLER_19_2131 ();
 sg13g2_fill_1 FILLER_19_2137 ();
 sg13g2_fill_2 FILLER_19_2174 ();
 sg13g2_fill_2 FILLER_19_2196 ();
 sg13g2_fill_2 FILLER_19_2207 ();
 sg13g2_fill_1 FILLER_19_2222 ();
 sg13g2_fill_2 FILLER_19_2244 ();
 sg13g2_fill_1 FILLER_19_2246 ();
 sg13g2_fill_1 FILLER_19_2264 ();
 sg13g2_fill_2 FILLER_19_2276 ();
 sg13g2_fill_1 FILLER_19_2293 ();
 sg13g2_fill_1 FILLER_19_2299 ();
 sg13g2_fill_1 FILLER_19_2333 ();
 sg13g2_decap_8 FILLER_19_2351 ();
 sg13g2_decap_8 FILLER_19_2358 ();
 sg13g2_decap_8 FILLER_19_2365 ();
 sg13g2_decap_8 FILLER_19_2372 ();
 sg13g2_decap_8 FILLER_19_2379 ();
 sg13g2_decap_8 FILLER_19_2386 ();
 sg13g2_decap_8 FILLER_19_2393 ();
 sg13g2_decap_8 FILLER_19_2400 ();
 sg13g2_decap_8 FILLER_19_2407 ();
 sg13g2_decap_8 FILLER_19_2414 ();
 sg13g2_decap_8 FILLER_19_2421 ();
 sg13g2_decap_8 FILLER_19_2428 ();
 sg13g2_decap_8 FILLER_19_2435 ();
 sg13g2_decap_8 FILLER_19_2442 ();
 sg13g2_decap_8 FILLER_19_2449 ();
 sg13g2_decap_8 FILLER_19_2456 ();
 sg13g2_decap_8 FILLER_19_2463 ();
 sg13g2_decap_8 FILLER_19_2470 ();
 sg13g2_decap_8 FILLER_19_2477 ();
 sg13g2_decap_8 FILLER_19_2484 ();
 sg13g2_decap_8 FILLER_19_2491 ();
 sg13g2_decap_8 FILLER_19_2498 ();
 sg13g2_decap_8 FILLER_19_2505 ();
 sg13g2_decap_8 FILLER_19_2512 ();
 sg13g2_decap_8 FILLER_19_2519 ();
 sg13g2_decap_8 FILLER_19_2526 ();
 sg13g2_decap_8 FILLER_19_2533 ();
 sg13g2_decap_8 FILLER_19_2540 ();
 sg13g2_decap_8 FILLER_19_2547 ();
 sg13g2_decap_8 FILLER_19_2554 ();
 sg13g2_decap_8 FILLER_19_2561 ();
 sg13g2_decap_8 FILLER_19_2568 ();
 sg13g2_decap_8 FILLER_19_2575 ();
 sg13g2_decap_8 FILLER_19_2582 ();
 sg13g2_decap_8 FILLER_19_2589 ();
 sg13g2_decap_8 FILLER_19_2596 ();
 sg13g2_decap_8 FILLER_19_2603 ();
 sg13g2_decap_8 FILLER_19_2610 ();
 sg13g2_decap_8 FILLER_19_2617 ();
 sg13g2_decap_8 FILLER_19_2624 ();
 sg13g2_decap_8 FILLER_19_2631 ();
 sg13g2_decap_8 FILLER_19_2638 ();
 sg13g2_decap_8 FILLER_19_2645 ();
 sg13g2_decap_8 FILLER_19_2652 ();
 sg13g2_decap_8 FILLER_19_2659 ();
 sg13g2_decap_8 FILLER_19_2666 ();
 sg13g2_fill_1 FILLER_19_2673 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_fill_1 FILLER_20_112 ();
 sg13g2_fill_2 FILLER_20_135 ();
 sg13g2_fill_1 FILLER_20_137 ();
 sg13g2_decap_4 FILLER_20_186 ();
 sg13g2_fill_2 FILLER_20_204 ();
 sg13g2_decap_8 FILLER_20_236 ();
 sg13g2_fill_1 FILLER_20_248 ();
 sg13g2_fill_2 FILLER_20_261 ();
 sg13g2_fill_1 FILLER_20_271 ();
 sg13g2_decap_4 FILLER_20_297 ();
 sg13g2_fill_2 FILLER_20_301 ();
 sg13g2_fill_1 FILLER_20_308 ();
 sg13g2_fill_2 FILLER_20_335 ();
 sg13g2_decap_4 FILLER_20_341 ();
 sg13g2_fill_1 FILLER_20_345 ();
 sg13g2_fill_1 FILLER_20_352 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_403 ();
 sg13g2_decap_4 FILLER_20_410 ();
 sg13g2_fill_1 FILLER_20_414 ();
 sg13g2_decap_4 FILLER_20_437 ();
 sg13g2_fill_2 FILLER_20_441 ();
 sg13g2_fill_2 FILLER_20_451 ();
 sg13g2_decap_8 FILLER_20_458 ();
 sg13g2_decap_4 FILLER_20_465 ();
 sg13g2_decap_4 FILLER_20_474 ();
 sg13g2_fill_1 FILLER_20_490 ();
 sg13g2_fill_2 FILLER_20_511 ();
 sg13g2_decap_4 FILLER_20_535 ();
 sg13g2_decap_4 FILLER_20_551 ();
 sg13g2_fill_1 FILLER_20_555 ();
 sg13g2_fill_1 FILLER_20_588 ();
 sg13g2_fill_1 FILLER_20_628 ();
 sg13g2_fill_1 FILLER_20_642 ();
 sg13g2_fill_2 FILLER_20_737 ();
 sg13g2_fill_1 FILLER_20_739 ();
 sg13g2_fill_2 FILLER_20_766 ();
 sg13g2_fill_1 FILLER_20_768 ();
 sg13g2_fill_1 FILLER_20_805 ();
 sg13g2_fill_1 FILLER_20_838 ();
 sg13g2_fill_1 FILLER_20_927 ();
 sg13g2_fill_2 FILLER_20_1018 ();
 sg13g2_fill_1 FILLER_20_1046 ();
 sg13g2_fill_2 FILLER_20_1120 ();
 sg13g2_fill_1 FILLER_20_1192 ();
 sg13g2_fill_1 FILLER_20_1202 ();
 sg13g2_fill_1 FILLER_20_1278 ();
 sg13g2_fill_1 FILLER_20_1306 ();
 sg13g2_fill_1 FILLER_20_1416 ();
 sg13g2_fill_1 FILLER_20_1593 ();
 sg13g2_fill_1 FILLER_20_1623 ();
 sg13g2_fill_1 FILLER_20_1639 ();
 sg13g2_fill_2 FILLER_20_1645 ();
 sg13g2_fill_1 FILLER_20_1677 ();
 sg13g2_fill_1 FILLER_20_1749 ();
 sg13g2_fill_2 FILLER_20_1799 ();
 sg13g2_fill_1 FILLER_20_1801 ();
 sg13g2_decap_8 FILLER_20_1828 ();
 sg13g2_fill_1 FILLER_20_1835 ();
 sg13g2_fill_2 FILLER_20_1850 ();
 sg13g2_fill_1 FILLER_20_1852 ();
 sg13g2_fill_2 FILLER_20_1895 ();
 sg13g2_fill_1 FILLER_20_1897 ();
 sg13g2_fill_1 FILLER_20_1924 ();
 sg13g2_decap_8 FILLER_20_1935 ();
 sg13g2_fill_1 FILLER_20_2008 ();
 sg13g2_decap_4 FILLER_20_2053 ();
 sg13g2_fill_2 FILLER_20_2086 ();
 sg13g2_fill_1 FILLER_20_2102 ();
 sg13g2_decap_4 FILLER_20_2112 ();
 sg13g2_decap_8 FILLER_20_2120 ();
 sg13g2_fill_2 FILLER_20_2127 ();
 sg13g2_fill_2 FILLER_20_2156 ();
 sg13g2_fill_2 FILLER_20_2162 ();
 sg13g2_fill_2 FILLER_20_2225 ();
 sg13g2_decap_4 FILLER_20_2263 ();
 sg13g2_fill_1 FILLER_20_2272 ();
 sg13g2_decap_8 FILLER_20_2350 ();
 sg13g2_decap_8 FILLER_20_2357 ();
 sg13g2_decap_8 FILLER_20_2364 ();
 sg13g2_decap_8 FILLER_20_2371 ();
 sg13g2_decap_8 FILLER_20_2378 ();
 sg13g2_decap_8 FILLER_20_2385 ();
 sg13g2_decap_8 FILLER_20_2392 ();
 sg13g2_decap_8 FILLER_20_2399 ();
 sg13g2_decap_8 FILLER_20_2406 ();
 sg13g2_decap_8 FILLER_20_2413 ();
 sg13g2_decap_8 FILLER_20_2420 ();
 sg13g2_decap_8 FILLER_20_2427 ();
 sg13g2_decap_8 FILLER_20_2434 ();
 sg13g2_decap_8 FILLER_20_2441 ();
 sg13g2_decap_8 FILLER_20_2448 ();
 sg13g2_decap_8 FILLER_20_2455 ();
 sg13g2_decap_8 FILLER_20_2462 ();
 sg13g2_decap_8 FILLER_20_2469 ();
 sg13g2_decap_8 FILLER_20_2476 ();
 sg13g2_decap_8 FILLER_20_2483 ();
 sg13g2_decap_8 FILLER_20_2490 ();
 sg13g2_decap_8 FILLER_20_2497 ();
 sg13g2_decap_8 FILLER_20_2504 ();
 sg13g2_decap_8 FILLER_20_2511 ();
 sg13g2_decap_8 FILLER_20_2518 ();
 sg13g2_decap_8 FILLER_20_2525 ();
 sg13g2_decap_8 FILLER_20_2532 ();
 sg13g2_decap_8 FILLER_20_2539 ();
 sg13g2_decap_8 FILLER_20_2546 ();
 sg13g2_decap_8 FILLER_20_2553 ();
 sg13g2_decap_8 FILLER_20_2560 ();
 sg13g2_decap_8 FILLER_20_2567 ();
 sg13g2_decap_8 FILLER_20_2574 ();
 sg13g2_decap_8 FILLER_20_2581 ();
 sg13g2_decap_8 FILLER_20_2588 ();
 sg13g2_decap_8 FILLER_20_2595 ();
 sg13g2_decap_8 FILLER_20_2602 ();
 sg13g2_decap_8 FILLER_20_2609 ();
 sg13g2_decap_8 FILLER_20_2616 ();
 sg13g2_decap_8 FILLER_20_2623 ();
 sg13g2_decap_8 FILLER_20_2630 ();
 sg13g2_decap_8 FILLER_20_2637 ();
 sg13g2_decap_8 FILLER_20_2644 ();
 sg13g2_decap_8 FILLER_20_2651 ();
 sg13g2_decap_8 FILLER_20_2658 ();
 sg13g2_decap_8 FILLER_20_2665 ();
 sg13g2_fill_2 FILLER_20_2672 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_fill_1 FILLER_21_112 ();
 sg13g2_fill_2 FILLER_21_139 ();
 sg13g2_fill_1 FILLER_21_141 ();
 sg13g2_decap_4 FILLER_21_151 ();
 sg13g2_decap_4 FILLER_21_182 ();
 sg13g2_fill_2 FILLER_21_194 ();
 sg13g2_fill_1 FILLER_21_196 ();
 sg13g2_fill_2 FILLER_21_214 ();
 sg13g2_fill_1 FILLER_21_216 ();
 sg13g2_decap_4 FILLER_21_221 ();
 sg13g2_fill_1 FILLER_21_225 ();
 sg13g2_decap_4 FILLER_21_231 ();
 sg13g2_fill_1 FILLER_21_235 ();
 sg13g2_fill_1 FILLER_21_249 ();
 sg13g2_fill_2 FILLER_21_267 ();
 sg13g2_fill_2 FILLER_21_281 ();
 sg13g2_fill_1 FILLER_21_283 ();
 sg13g2_decap_8 FILLER_21_289 ();
 sg13g2_decap_4 FILLER_21_336 ();
 sg13g2_decap_4 FILLER_21_348 ();
 sg13g2_fill_1 FILLER_21_392 ();
 sg13g2_fill_1 FILLER_21_405 ();
 sg13g2_fill_1 FILLER_21_459 ();
 sg13g2_decap_4 FILLER_21_477 ();
 sg13g2_fill_2 FILLER_21_486 ();
 sg13g2_fill_1 FILLER_21_488 ();
 sg13g2_fill_1 FILLER_21_590 ();
 sg13g2_fill_2 FILLER_21_600 ();
 sg13g2_fill_1 FILLER_21_611 ();
 sg13g2_fill_1 FILLER_21_626 ();
 sg13g2_fill_2 FILLER_21_648 ();
 sg13g2_fill_1 FILLER_21_650 ();
 sg13g2_fill_1 FILLER_21_665 ();
 sg13g2_fill_2 FILLER_21_682 ();
 sg13g2_fill_1 FILLER_21_684 ();
 sg13g2_fill_1 FILLER_21_702 ();
 sg13g2_fill_1 FILLER_21_768 ();
 sg13g2_fill_2 FILLER_21_779 ();
 sg13g2_fill_1 FILLER_21_781 ();
 sg13g2_fill_2 FILLER_21_826 ();
 sg13g2_fill_1 FILLER_21_841 ();
 sg13g2_fill_1 FILLER_21_869 ();
 sg13g2_fill_2 FILLER_21_940 ();
 sg13g2_fill_1 FILLER_21_1009 ();
 sg13g2_fill_1 FILLER_21_1051 ();
 sg13g2_fill_1 FILLER_21_1391 ();
 sg13g2_fill_1 FILLER_21_1454 ();
 sg13g2_fill_2 FILLER_21_1556 ();
 sg13g2_fill_1 FILLER_21_1584 ();
 sg13g2_fill_1 FILLER_21_1593 ();
 sg13g2_fill_2 FILLER_21_1628 ();
 sg13g2_fill_1 FILLER_21_1664 ();
 sg13g2_fill_2 FILLER_21_1699 ();
 sg13g2_fill_2 FILLER_21_1723 ();
 sg13g2_fill_1 FILLER_21_1753 ();
 sg13g2_fill_1 FILLER_21_1763 ();
 sg13g2_fill_2 FILLER_21_1777 ();
 sg13g2_fill_2 FILLER_21_1797 ();
 sg13g2_decap_8 FILLER_21_1840 ();
 sg13g2_decap_4 FILLER_21_1882 ();
 sg13g2_decap_8 FILLER_21_1922 ();
 sg13g2_decap_4 FILLER_21_1985 ();
 sg13g2_fill_2 FILLER_21_2025 ();
 sg13g2_fill_1 FILLER_21_2039 ();
 sg13g2_fill_2 FILLER_21_2092 ();
 sg13g2_decap_4 FILLER_21_2120 ();
 sg13g2_fill_2 FILLER_21_2124 ();
 sg13g2_decap_4 FILLER_21_2139 ();
 sg13g2_fill_1 FILLER_21_2143 ();
 sg13g2_fill_1 FILLER_21_2179 ();
 sg13g2_fill_2 FILLER_21_2224 ();
 sg13g2_decap_4 FILLER_21_2246 ();
 sg13g2_fill_1 FILLER_21_2250 ();
 sg13g2_fill_2 FILLER_21_2277 ();
 sg13g2_fill_1 FILLER_21_2279 ();
 sg13g2_fill_2 FILLER_21_2290 ();
 sg13g2_fill_1 FILLER_21_2322 ();
 sg13g2_decap_8 FILLER_21_2349 ();
 sg13g2_decap_8 FILLER_21_2356 ();
 sg13g2_decap_8 FILLER_21_2363 ();
 sg13g2_decap_8 FILLER_21_2370 ();
 sg13g2_decap_8 FILLER_21_2377 ();
 sg13g2_decap_8 FILLER_21_2384 ();
 sg13g2_decap_8 FILLER_21_2391 ();
 sg13g2_decap_8 FILLER_21_2398 ();
 sg13g2_decap_8 FILLER_21_2405 ();
 sg13g2_decap_8 FILLER_21_2412 ();
 sg13g2_decap_8 FILLER_21_2419 ();
 sg13g2_decap_8 FILLER_21_2426 ();
 sg13g2_decap_8 FILLER_21_2433 ();
 sg13g2_decap_8 FILLER_21_2440 ();
 sg13g2_decap_8 FILLER_21_2447 ();
 sg13g2_decap_8 FILLER_21_2454 ();
 sg13g2_decap_8 FILLER_21_2461 ();
 sg13g2_decap_8 FILLER_21_2468 ();
 sg13g2_decap_8 FILLER_21_2475 ();
 sg13g2_decap_8 FILLER_21_2482 ();
 sg13g2_decap_8 FILLER_21_2489 ();
 sg13g2_decap_8 FILLER_21_2496 ();
 sg13g2_decap_8 FILLER_21_2503 ();
 sg13g2_decap_8 FILLER_21_2510 ();
 sg13g2_decap_8 FILLER_21_2517 ();
 sg13g2_decap_8 FILLER_21_2524 ();
 sg13g2_decap_8 FILLER_21_2531 ();
 sg13g2_decap_8 FILLER_21_2538 ();
 sg13g2_decap_8 FILLER_21_2545 ();
 sg13g2_decap_8 FILLER_21_2552 ();
 sg13g2_decap_8 FILLER_21_2559 ();
 sg13g2_decap_8 FILLER_21_2566 ();
 sg13g2_decap_8 FILLER_21_2573 ();
 sg13g2_decap_8 FILLER_21_2580 ();
 sg13g2_decap_8 FILLER_21_2587 ();
 sg13g2_decap_8 FILLER_21_2594 ();
 sg13g2_decap_8 FILLER_21_2601 ();
 sg13g2_decap_8 FILLER_21_2608 ();
 sg13g2_decap_8 FILLER_21_2615 ();
 sg13g2_decap_8 FILLER_21_2622 ();
 sg13g2_decap_8 FILLER_21_2629 ();
 sg13g2_decap_8 FILLER_21_2636 ();
 sg13g2_decap_8 FILLER_21_2643 ();
 sg13g2_decap_8 FILLER_21_2650 ();
 sg13g2_decap_8 FILLER_21_2657 ();
 sg13g2_decap_8 FILLER_21_2664 ();
 sg13g2_fill_2 FILLER_21_2671 ();
 sg13g2_fill_1 FILLER_21_2673 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_fill_2 FILLER_22_112 ();
 sg13g2_fill_1 FILLER_22_114 ();
 sg13g2_fill_1 FILLER_22_141 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_4 FILLER_22_198 ();
 sg13g2_fill_2 FILLER_22_202 ();
 sg13g2_fill_1 FILLER_22_216 ();
 sg13g2_fill_2 FILLER_22_224 ();
 sg13g2_fill_2 FILLER_22_231 ();
 sg13g2_fill_1 FILLER_22_233 ();
 sg13g2_fill_2 FILLER_22_256 ();
 sg13g2_decap_4 FILLER_22_270 ();
 sg13g2_decap_8 FILLER_22_279 ();
 sg13g2_fill_2 FILLER_22_286 ();
 sg13g2_fill_1 FILLER_22_288 ();
 sg13g2_decap_4 FILLER_22_293 ();
 sg13g2_decap_4 FILLER_22_312 ();
 sg13g2_fill_1 FILLER_22_316 ();
 sg13g2_decap_8 FILLER_22_333 ();
 sg13g2_decap_4 FILLER_22_340 ();
 sg13g2_fill_1 FILLER_22_344 ();
 sg13g2_fill_1 FILLER_22_369 ();
 sg13g2_fill_2 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_439 ();
 sg13g2_fill_1 FILLER_22_461 ();
 sg13g2_fill_2 FILLER_22_470 ();
 sg13g2_fill_2 FILLER_22_490 ();
 sg13g2_decap_8 FILLER_22_511 ();
 sg13g2_fill_1 FILLER_22_518 ();
 sg13g2_fill_1 FILLER_22_543 ();
 sg13g2_decap_4 FILLER_22_560 ();
 sg13g2_fill_1 FILLER_22_606 ();
 sg13g2_fill_2 FILLER_22_618 ();
 sg13g2_fill_1 FILLER_22_620 ();
 sg13g2_fill_2 FILLER_22_626 ();
 sg13g2_fill_2 FILLER_22_695 ();
 sg13g2_fill_2 FILLER_22_707 ();
 sg13g2_fill_1 FILLER_22_709 ();
 sg13g2_fill_2 FILLER_22_765 ();
 sg13g2_decap_4 FILLER_22_784 ();
 sg13g2_fill_1 FILLER_22_788 ();
 sg13g2_fill_1 FILLER_22_809 ();
 sg13g2_fill_2 FILLER_22_815 ();
 sg13g2_fill_1 FILLER_22_817 ();
 sg13g2_decap_8 FILLER_22_836 ();
 sg13g2_fill_2 FILLER_22_843 ();
 sg13g2_fill_1 FILLER_22_910 ();
 sg13g2_fill_1 FILLER_22_956 ();
 sg13g2_fill_1 FILLER_22_1000 ();
 sg13g2_fill_1 FILLER_22_1108 ();
 sg13g2_fill_1 FILLER_22_1162 ();
 sg13g2_fill_1 FILLER_22_1185 ();
 sg13g2_fill_1 FILLER_22_1217 ();
 sg13g2_fill_1 FILLER_22_1254 ();
 sg13g2_fill_1 FILLER_22_1381 ();
 sg13g2_fill_1 FILLER_22_1451 ();
 sg13g2_fill_1 FILLER_22_1530 ();
 sg13g2_fill_2 FILLER_22_1550 ();
 sg13g2_fill_1 FILLER_22_1593 ();
 sg13g2_fill_1 FILLER_22_1630 ();
 sg13g2_fill_2 FILLER_22_1686 ();
 sg13g2_fill_2 FILLER_22_1727 ();
 sg13g2_fill_2 FILLER_22_1850 ();
 sg13g2_fill_1 FILLER_22_1852 ();
 sg13g2_fill_1 FILLER_22_1871 ();
 sg13g2_fill_2 FILLER_22_1880 ();
 sg13g2_decap_8 FILLER_22_1888 ();
 sg13g2_decap_8 FILLER_22_1895 ();
 sg13g2_decap_4 FILLER_22_1902 ();
 sg13g2_decap_8 FILLER_22_1923 ();
 sg13g2_fill_2 FILLER_22_1930 ();
 sg13g2_fill_1 FILLER_22_1932 ();
 sg13g2_decap_4 FILLER_22_1951 ();
 sg13g2_fill_2 FILLER_22_2037 ();
 sg13g2_fill_1 FILLER_22_2056 ();
 sg13g2_fill_2 FILLER_22_2061 ();
 sg13g2_fill_1 FILLER_22_2063 ();
 sg13g2_fill_1 FILLER_22_2073 ();
 sg13g2_fill_1 FILLER_22_2104 ();
 sg13g2_fill_2 FILLER_22_2123 ();
 sg13g2_fill_1 FILLER_22_2125 ();
 sg13g2_decap_8 FILLER_22_2130 ();
 sg13g2_fill_2 FILLER_22_2137 ();
 sg13g2_fill_2 FILLER_22_2149 ();
 sg13g2_fill_1 FILLER_22_2151 ();
 sg13g2_fill_2 FILLER_22_2165 ();
 sg13g2_fill_1 FILLER_22_2175 ();
 sg13g2_decap_4 FILLER_22_2184 ();
 sg13g2_fill_1 FILLER_22_2207 ();
 sg13g2_fill_1 FILLER_22_2251 ();
 sg13g2_decap_8 FILLER_22_2281 ();
 sg13g2_fill_1 FILLER_22_2292 ();
 sg13g2_decap_4 FILLER_22_2303 ();
 sg13g2_decap_8 FILLER_22_2324 ();
 sg13g2_fill_2 FILLER_22_2331 ();
 sg13g2_decap_8 FILLER_22_2346 ();
 sg13g2_decap_8 FILLER_22_2353 ();
 sg13g2_decap_8 FILLER_22_2360 ();
 sg13g2_decap_8 FILLER_22_2367 ();
 sg13g2_decap_8 FILLER_22_2374 ();
 sg13g2_decap_8 FILLER_22_2381 ();
 sg13g2_decap_8 FILLER_22_2388 ();
 sg13g2_decap_8 FILLER_22_2395 ();
 sg13g2_decap_8 FILLER_22_2402 ();
 sg13g2_decap_8 FILLER_22_2409 ();
 sg13g2_decap_8 FILLER_22_2416 ();
 sg13g2_decap_8 FILLER_22_2423 ();
 sg13g2_decap_8 FILLER_22_2430 ();
 sg13g2_decap_8 FILLER_22_2437 ();
 sg13g2_decap_8 FILLER_22_2444 ();
 sg13g2_decap_8 FILLER_22_2451 ();
 sg13g2_decap_8 FILLER_22_2458 ();
 sg13g2_decap_8 FILLER_22_2465 ();
 sg13g2_decap_8 FILLER_22_2472 ();
 sg13g2_decap_8 FILLER_22_2479 ();
 sg13g2_decap_8 FILLER_22_2486 ();
 sg13g2_decap_8 FILLER_22_2493 ();
 sg13g2_decap_8 FILLER_22_2500 ();
 sg13g2_decap_8 FILLER_22_2507 ();
 sg13g2_decap_8 FILLER_22_2514 ();
 sg13g2_decap_8 FILLER_22_2521 ();
 sg13g2_decap_8 FILLER_22_2528 ();
 sg13g2_decap_8 FILLER_22_2535 ();
 sg13g2_decap_8 FILLER_22_2542 ();
 sg13g2_decap_8 FILLER_22_2549 ();
 sg13g2_decap_8 FILLER_22_2556 ();
 sg13g2_decap_8 FILLER_22_2563 ();
 sg13g2_decap_8 FILLER_22_2570 ();
 sg13g2_decap_8 FILLER_22_2577 ();
 sg13g2_decap_8 FILLER_22_2584 ();
 sg13g2_decap_8 FILLER_22_2591 ();
 sg13g2_decap_8 FILLER_22_2598 ();
 sg13g2_decap_8 FILLER_22_2605 ();
 sg13g2_decap_8 FILLER_22_2612 ();
 sg13g2_decap_8 FILLER_22_2619 ();
 sg13g2_decap_8 FILLER_22_2626 ();
 sg13g2_decap_8 FILLER_22_2633 ();
 sg13g2_decap_8 FILLER_22_2640 ();
 sg13g2_decap_8 FILLER_22_2647 ();
 sg13g2_decap_8 FILLER_22_2654 ();
 sg13g2_decap_8 FILLER_22_2661 ();
 sg13g2_decap_4 FILLER_22_2668 ();
 sg13g2_fill_2 FILLER_22_2672 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_fill_1 FILLER_23_131 ();
 sg13g2_fill_1 FILLER_23_175 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_fill_2 FILLER_23_193 ();
 sg13g2_fill_1 FILLER_23_199 ();
 sg13g2_fill_2 FILLER_23_206 ();
 sg13g2_fill_1 FILLER_23_208 ();
 sg13g2_decap_8 FILLER_23_232 ();
 sg13g2_fill_1 FILLER_23_239 ();
 sg13g2_fill_1 FILLER_23_255 ();
 sg13g2_fill_2 FILLER_23_275 ();
 sg13g2_fill_1 FILLER_23_277 ();
 sg13g2_fill_2 FILLER_23_304 ();
 sg13g2_fill_1 FILLER_23_306 ();
 sg13g2_decap_8 FILLER_23_319 ();
 sg13g2_fill_2 FILLER_23_326 ();
 sg13g2_fill_2 FILLER_23_388 ();
 sg13g2_fill_2 FILLER_23_397 ();
 sg13g2_fill_1 FILLER_23_425 ();
 sg13g2_fill_1 FILLER_23_447 ();
 sg13g2_fill_2 FILLER_23_456 ();
 sg13g2_fill_1 FILLER_23_458 ();
 sg13g2_decap_4 FILLER_23_473 ();
 sg13g2_fill_2 FILLER_23_499 ();
 sg13g2_fill_1 FILLER_23_501 ();
 sg13g2_decap_8 FILLER_23_536 ();
 sg13g2_decap_4 FILLER_23_551 ();
 sg13g2_fill_2 FILLER_23_555 ();
 sg13g2_fill_2 FILLER_23_569 ();
 sg13g2_fill_2 FILLER_23_636 ();
 sg13g2_fill_2 FILLER_23_652 ();
 sg13g2_fill_1 FILLER_23_669 ();
 sg13g2_fill_2 FILLER_23_733 ();
 sg13g2_fill_1 FILLER_23_795 ();
 sg13g2_fill_2 FILLER_23_808 ();
 sg13g2_fill_1 FILLER_23_810 ();
 sg13g2_fill_2 FILLER_23_836 ();
 sg13g2_fill_2 FILLER_23_851 ();
 sg13g2_fill_1 FILLER_23_862 ();
 sg13g2_fill_2 FILLER_23_926 ();
 sg13g2_fill_2 FILLER_23_950 ();
 sg13g2_fill_2 FILLER_23_1015 ();
 sg13g2_fill_2 FILLER_23_1026 ();
 sg13g2_fill_1 FILLER_23_1043 ();
 sg13g2_fill_2 FILLER_23_1144 ();
 sg13g2_fill_1 FILLER_23_1194 ();
 sg13g2_fill_2 FILLER_23_1282 ();
 sg13g2_fill_1 FILLER_23_1476 ();
 sg13g2_fill_2 FILLER_23_1509 ();
 sg13g2_fill_1 FILLER_23_1625 ();
 sg13g2_fill_2 FILLER_23_1664 ();
 sg13g2_fill_1 FILLER_23_1675 ();
 sg13g2_fill_2 FILLER_23_1702 ();
 sg13g2_fill_2 FILLER_23_1755 ();
 sg13g2_fill_2 FILLER_23_1779 ();
 sg13g2_fill_1 FILLER_23_1781 ();
 sg13g2_fill_2 FILLER_23_1839 ();
 sg13g2_decap_4 FILLER_23_1866 ();
 sg13g2_fill_1 FILLER_23_1870 ();
 sg13g2_fill_2 FILLER_23_1882 ();
 sg13g2_decap_8 FILLER_23_1893 ();
 sg13g2_decap_4 FILLER_23_1926 ();
 sg13g2_fill_1 FILLER_23_1930 ();
 sg13g2_decap_8 FILLER_23_1936 ();
 sg13g2_fill_2 FILLER_23_2016 ();
 sg13g2_fill_1 FILLER_23_2018 ();
 sg13g2_fill_1 FILLER_23_2055 ();
 sg13g2_fill_2 FILLER_23_2065 ();
 sg13g2_fill_1 FILLER_23_2067 ();
 sg13g2_fill_2 FILLER_23_2074 ();
 sg13g2_fill_1 FILLER_23_2076 ();
 sg13g2_decap_4 FILLER_23_2088 ();
 sg13g2_fill_1 FILLER_23_2092 ();
 sg13g2_fill_2 FILLER_23_2098 ();
 sg13g2_fill_1 FILLER_23_2100 ();
 sg13g2_fill_2 FILLER_23_2141 ();
 sg13g2_decap_8 FILLER_23_2235 ();
 sg13g2_decap_4 FILLER_23_2242 ();
 sg13g2_fill_1 FILLER_23_2246 ();
 sg13g2_decap_8 FILLER_23_2333 ();
 sg13g2_decap_8 FILLER_23_2340 ();
 sg13g2_decap_8 FILLER_23_2347 ();
 sg13g2_decap_8 FILLER_23_2354 ();
 sg13g2_decap_8 FILLER_23_2361 ();
 sg13g2_decap_8 FILLER_23_2368 ();
 sg13g2_decap_8 FILLER_23_2375 ();
 sg13g2_decap_8 FILLER_23_2382 ();
 sg13g2_decap_8 FILLER_23_2389 ();
 sg13g2_decap_8 FILLER_23_2396 ();
 sg13g2_decap_8 FILLER_23_2403 ();
 sg13g2_decap_8 FILLER_23_2410 ();
 sg13g2_decap_8 FILLER_23_2417 ();
 sg13g2_decap_8 FILLER_23_2424 ();
 sg13g2_decap_8 FILLER_23_2431 ();
 sg13g2_decap_8 FILLER_23_2438 ();
 sg13g2_decap_8 FILLER_23_2445 ();
 sg13g2_decap_8 FILLER_23_2452 ();
 sg13g2_decap_8 FILLER_23_2459 ();
 sg13g2_decap_8 FILLER_23_2466 ();
 sg13g2_decap_8 FILLER_23_2473 ();
 sg13g2_decap_8 FILLER_23_2480 ();
 sg13g2_decap_8 FILLER_23_2487 ();
 sg13g2_decap_8 FILLER_23_2494 ();
 sg13g2_decap_8 FILLER_23_2501 ();
 sg13g2_decap_8 FILLER_23_2508 ();
 sg13g2_decap_8 FILLER_23_2515 ();
 sg13g2_decap_8 FILLER_23_2522 ();
 sg13g2_decap_8 FILLER_23_2529 ();
 sg13g2_decap_8 FILLER_23_2536 ();
 sg13g2_decap_8 FILLER_23_2543 ();
 sg13g2_decap_8 FILLER_23_2550 ();
 sg13g2_decap_8 FILLER_23_2557 ();
 sg13g2_decap_8 FILLER_23_2564 ();
 sg13g2_decap_8 FILLER_23_2571 ();
 sg13g2_decap_8 FILLER_23_2578 ();
 sg13g2_decap_8 FILLER_23_2585 ();
 sg13g2_decap_8 FILLER_23_2592 ();
 sg13g2_decap_8 FILLER_23_2599 ();
 sg13g2_decap_8 FILLER_23_2606 ();
 sg13g2_decap_8 FILLER_23_2613 ();
 sg13g2_decap_8 FILLER_23_2620 ();
 sg13g2_decap_8 FILLER_23_2627 ();
 sg13g2_decap_8 FILLER_23_2634 ();
 sg13g2_decap_8 FILLER_23_2641 ();
 sg13g2_decap_8 FILLER_23_2648 ();
 sg13g2_decap_8 FILLER_23_2655 ();
 sg13g2_decap_8 FILLER_23_2662 ();
 sg13g2_decap_4 FILLER_23_2669 ();
 sg13g2_fill_1 FILLER_23_2673 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_4 FILLER_24_176 ();
 sg13g2_fill_1 FILLER_24_180 ();
 sg13g2_fill_2 FILLER_24_186 ();
 sg13g2_fill_1 FILLER_24_188 ();
 sg13g2_fill_2 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_221 ();
 sg13g2_decap_4 FILLER_24_228 ();
 sg13g2_decap_8 FILLER_24_240 ();
 sg13g2_decap_4 FILLER_24_247 ();
 sg13g2_fill_1 FILLER_24_256 ();
 sg13g2_fill_1 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_fill_1 FILLER_24_287 ();
 sg13g2_fill_1 FILLER_24_296 ();
 sg13g2_decap_4 FILLER_24_313 ();
 sg13g2_fill_1 FILLER_24_317 ();
 sg13g2_decap_8 FILLER_24_331 ();
 sg13g2_fill_1 FILLER_24_338 ();
 sg13g2_fill_2 FILLER_24_368 ();
 sg13g2_fill_1 FILLER_24_375 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_fill_2 FILLER_24_437 ();
 sg13g2_fill_1 FILLER_24_439 ();
 sg13g2_fill_2 FILLER_24_459 ();
 sg13g2_fill_1 FILLER_24_495 ();
 sg13g2_fill_1 FILLER_24_501 ();
 sg13g2_fill_2 FILLER_24_511 ();
 sg13g2_fill_2 FILLER_24_517 ();
 sg13g2_fill_2 FILLER_24_594 ();
 sg13g2_fill_1 FILLER_24_604 ();
 sg13g2_fill_1 FILLER_24_662 ();
 sg13g2_fill_1 FILLER_24_677 ();
 sg13g2_fill_2 FILLER_24_696 ();
 sg13g2_decap_4 FILLER_24_703 ();
 sg13g2_fill_2 FILLER_24_722 ();
 sg13g2_fill_2 FILLER_24_738 ();
 sg13g2_fill_1 FILLER_24_740 ();
 sg13g2_decap_8 FILLER_24_785 ();
 sg13g2_fill_2 FILLER_24_792 ();
 sg13g2_fill_1 FILLER_24_794 ();
 sg13g2_fill_1 FILLER_24_802 ();
 sg13g2_fill_1 FILLER_24_815 ();
 sg13g2_fill_1 FILLER_24_834 ();
 sg13g2_fill_2 FILLER_24_848 ();
 sg13g2_fill_1 FILLER_24_882 ();
 sg13g2_fill_1 FILLER_24_978 ();
 sg13g2_fill_2 FILLER_24_1021 ();
 sg13g2_fill_2 FILLER_24_1058 ();
 sg13g2_fill_2 FILLER_24_1285 ();
 sg13g2_fill_1 FILLER_24_1315 ();
 sg13g2_fill_1 FILLER_24_1334 ();
 sg13g2_fill_2 FILLER_24_1378 ();
 sg13g2_fill_1 FILLER_24_1448 ();
 sg13g2_fill_1 FILLER_24_1475 ();
 sg13g2_fill_1 FILLER_24_1485 ();
 sg13g2_fill_1 FILLER_24_1524 ();
 sg13g2_fill_2 FILLER_24_1553 ();
 sg13g2_fill_2 FILLER_24_1599 ();
 sg13g2_fill_1 FILLER_24_1645 ();
 sg13g2_fill_1 FILLER_24_1719 ();
 sg13g2_fill_2 FILLER_24_1755 ();
 sg13g2_decap_8 FILLER_24_1833 ();
 sg13g2_fill_1 FILLER_24_1840 ();
 sg13g2_fill_2 FILLER_24_1845 ();
 sg13g2_fill_1 FILLER_24_1847 ();
 sg13g2_fill_1 FILLER_24_1940 ();
 sg13g2_decap_8 FILLER_24_1945 ();
 sg13g2_fill_2 FILLER_24_1952 ();
 sg13g2_decap_8 FILLER_24_1958 ();
 sg13g2_decap_8 FILLER_24_1965 ();
 sg13g2_fill_2 FILLER_24_1972 ();
 sg13g2_decap_8 FILLER_24_1983 ();
 sg13g2_decap_4 FILLER_24_1990 ();
 sg13g2_fill_2 FILLER_24_1994 ();
 sg13g2_fill_2 FILLER_24_2009 ();
 sg13g2_fill_1 FILLER_24_2011 ();
 sg13g2_fill_1 FILLER_24_2021 ();
 sg13g2_decap_4 FILLER_24_2032 ();
 sg13g2_decap_4 FILLER_24_2080 ();
 sg13g2_fill_1 FILLER_24_2139 ();
 sg13g2_decap_8 FILLER_24_2149 ();
 sg13g2_decap_4 FILLER_24_2156 ();
 sg13g2_fill_1 FILLER_24_2160 ();
 sg13g2_fill_1 FILLER_24_2205 ();
 sg13g2_decap_4 FILLER_24_2241 ();
 sg13g2_fill_1 FILLER_24_2245 ();
 sg13g2_fill_2 FILLER_24_2250 ();
 sg13g2_decap_8 FILLER_24_2256 ();
 sg13g2_fill_2 FILLER_24_2263 ();
 sg13g2_fill_2 FILLER_24_2274 ();
 sg13g2_fill_2 FILLER_24_2286 ();
 sg13g2_fill_1 FILLER_24_2288 ();
 sg13g2_decap_8 FILLER_24_2330 ();
 sg13g2_decap_8 FILLER_24_2337 ();
 sg13g2_decap_8 FILLER_24_2344 ();
 sg13g2_decap_8 FILLER_24_2351 ();
 sg13g2_decap_8 FILLER_24_2358 ();
 sg13g2_decap_8 FILLER_24_2365 ();
 sg13g2_decap_8 FILLER_24_2372 ();
 sg13g2_decap_8 FILLER_24_2379 ();
 sg13g2_decap_8 FILLER_24_2386 ();
 sg13g2_decap_8 FILLER_24_2393 ();
 sg13g2_decap_8 FILLER_24_2400 ();
 sg13g2_decap_8 FILLER_24_2407 ();
 sg13g2_decap_8 FILLER_24_2414 ();
 sg13g2_decap_8 FILLER_24_2421 ();
 sg13g2_decap_8 FILLER_24_2428 ();
 sg13g2_decap_8 FILLER_24_2435 ();
 sg13g2_decap_8 FILLER_24_2442 ();
 sg13g2_decap_8 FILLER_24_2449 ();
 sg13g2_decap_8 FILLER_24_2456 ();
 sg13g2_decap_8 FILLER_24_2463 ();
 sg13g2_decap_8 FILLER_24_2470 ();
 sg13g2_decap_8 FILLER_24_2477 ();
 sg13g2_decap_8 FILLER_24_2484 ();
 sg13g2_decap_8 FILLER_24_2491 ();
 sg13g2_decap_8 FILLER_24_2498 ();
 sg13g2_decap_8 FILLER_24_2505 ();
 sg13g2_decap_8 FILLER_24_2512 ();
 sg13g2_decap_8 FILLER_24_2519 ();
 sg13g2_decap_8 FILLER_24_2526 ();
 sg13g2_decap_8 FILLER_24_2533 ();
 sg13g2_decap_8 FILLER_24_2540 ();
 sg13g2_decap_8 FILLER_24_2547 ();
 sg13g2_decap_8 FILLER_24_2554 ();
 sg13g2_decap_8 FILLER_24_2561 ();
 sg13g2_decap_8 FILLER_24_2568 ();
 sg13g2_decap_8 FILLER_24_2575 ();
 sg13g2_decap_8 FILLER_24_2582 ();
 sg13g2_decap_8 FILLER_24_2589 ();
 sg13g2_decap_8 FILLER_24_2596 ();
 sg13g2_decap_8 FILLER_24_2603 ();
 sg13g2_decap_8 FILLER_24_2610 ();
 sg13g2_decap_8 FILLER_24_2617 ();
 sg13g2_decap_8 FILLER_24_2624 ();
 sg13g2_decap_8 FILLER_24_2631 ();
 sg13g2_decap_8 FILLER_24_2638 ();
 sg13g2_decap_8 FILLER_24_2645 ();
 sg13g2_decap_8 FILLER_24_2652 ();
 sg13g2_decap_8 FILLER_24_2659 ();
 sg13g2_decap_8 FILLER_24_2666 ();
 sg13g2_fill_1 FILLER_24_2673 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_4 FILLER_25_98 ();
 sg13g2_fill_1 FILLER_25_102 ();
 sg13g2_fill_1 FILLER_25_180 ();
 sg13g2_fill_1 FILLER_25_203 ();
 sg13g2_decap_4 FILLER_25_216 ();
 sg13g2_decap_8 FILLER_25_236 ();
 sg13g2_fill_1 FILLER_25_248 ();
 sg13g2_fill_1 FILLER_25_279 ();
 sg13g2_decap_4 FILLER_25_300 ();
 sg13g2_fill_2 FILLER_25_304 ();
 sg13g2_fill_2 FILLER_25_311 ();
 sg13g2_fill_1 FILLER_25_313 ();
 sg13g2_fill_2 FILLER_25_330 ();
 sg13g2_fill_1 FILLER_25_332 ();
 sg13g2_fill_2 FILLER_25_349 ();
 sg13g2_decap_4 FILLER_25_357 ();
 sg13g2_fill_1 FILLER_25_367 ();
 sg13g2_fill_1 FILLER_25_383 ();
 sg13g2_fill_2 FILLER_25_415 ();
 sg13g2_fill_1 FILLER_25_430 ();
 sg13g2_decap_4 FILLER_25_450 ();
 sg13g2_fill_2 FILLER_25_454 ();
 sg13g2_decap_8 FILLER_25_464 ();
 sg13g2_fill_2 FILLER_25_505 ();
 sg13g2_fill_2 FILLER_25_512 ();
 sg13g2_fill_2 FILLER_25_531 ();
 sg13g2_fill_1 FILLER_25_533 ();
 sg13g2_fill_2 FILLER_25_571 ();
 sg13g2_fill_2 FILLER_25_649 ();
 sg13g2_fill_2 FILLER_25_664 ();
 sg13g2_fill_1 FILLER_25_666 ();
 sg13g2_fill_2 FILLER_25_693 ();
 sg13g2_fill_2 FILLER_25_719 ();
 sg13g2_fill_1 FILLER_25_721 ();
 sg13g2_decap_4 FILLER_25_769 ();
 sg13g2_fill_2 FILLER_25_773 ();
 sg13g2_decap_8 FILLER_25_779 ();
 sg13g2_fill_2 FILLER_25_786 ();
 sg13g2_decap_4 FILLER_25_791 ();
 sg13g2_fill_1 FILLER_25_795 ();
 sg13g2_fill_2 FILLER_25_819 ();
 sg13g2_fill_1 FILLER_25_851 ();
 sg13g2_fill_2 FILLER_25_861 ();
 sg13g2_fill_2 FILLER_25_888 ();
 sg13g2_fill_2 FILLER_25_920 ();
 sg13g2_fill_2 FILLER_25_953 ();
 sg13g2_fill_2 FILLER_25_1003 ();
 sg13g2_fill_1 FILLER_25_1036 ();
 sg13g2_fill_2 FILLER_25_1152 ();
 sg13g2_fill_1 FILLER_25_1194 ();
 sg13g2_fill_1 FILLER_25_1456 ();
 sg13g2_fill_1 FILLER_25_1506 ();
 sg13g2_fill_2 FILLER_25_1715 ();
 sg13g2_fill_1 FILLER_25_1722 ();
 sg13g2_fill_1 FILLER_25_1786 ();
 sg13g2_fill_1 FILLER_25_1815 ();
 sg13g2_decap_8 FILLER_25_1847 ();
 sg13g2_fill_1 FILLER_25_1854 ();
 sg13g2_fill_1 FILLER_25_1907 ();
 sg13g2_decap_8 FILLER_25_1912 ();
 sg13g2_fill_2 FILLER_25_1919 ();
 sg13g2_fill_1 FILLER_25_1921 ();
 sg13g2_decap_4 FILLER_25_1926 ();
 sg13g2_fill_2 FILLER_25_1956 ();
 sg13g2_fill_2 FILLER_25_1966 ();
 sg13g2_fill_1 FILLER_25_1968 ();
 sg13g2_fill_2 FILLER_25_1985 ();
 sg13g2_fill_2 FILLER_25_2063 ();
 sg13g2_fill_1 FILLER_25_2095 ();
 sg13g2_fill_1 FILLER_25_2107 ();
 sg13g2_fill_2 FILLER_25_2127 ();
 sg13g2_fill_1 FILLER_25_2129 ();
 sg13g2_fill_2 FILLER_25_2156 ();
 sg13g2_fill_1 FILLER_25_2158 ();
 sg13g2_fill_2 FILLER_25_2177 ();
 sg13g2_decap_8 FILLER_25_2224 ();
 sg13g2_decap_8 FILLER_25_2334 ();
 sg13g2_decap_8 FILLER_25_2341 ();
 sg13g2_decap_8 FILLER_25_2348 ();
 sg13g2_decap_8 FILLER_25_2355 ();
 sg13g2_decap_8 FILLER_25_2362 ();
 sg13g2_decap_8 FILLER_25_2369 ();
 sg13g2_decap_8 FILLER_25_2376 ();
 sg13g2_decap_8 FILLER_25_2383 ();
 sg13g2_decap_8 FILLER_25_2390 ();
 sg13g2_decap_8 FILLER_25_2397 ();
 sg13g2_decap_8 FILLER_25_2404 ();
 sg13g2_decap_8 FILLER_25_2411 ();
 sg13g2_decap_8 FILLER_25_2418 ();
 sg13g2_decap_8 FILLER_25_2425 ();
 sg13g2_decap_8 FILLER_25_2432 ();
 sg13g2_decap_8 FILLER_25_2439 ();
 sg13g2_decap_8 FILLER_25_2446 ();
 sg13g2_decap_8 FILLER_25_2453 ();
 sg13g2_decap_8 FILLER_25_2460 ();
 sg13g2_decap_8 FILLER_25_2467 ();
 sg13g2_decap_8 FILLER_25_2474 ();
 sg13g2_decap_8 FILLER_25_2481 ();
 sg13g2_decap_8 FILLER_25_2488 ();
 sg13g2_decap_8 FILLER_25_2495 ();
 sg13g2_decap_8 FILLER_25_2502 ();
 sg13g2_decap_8 FILLER_25_2509 ();
 sg13g2_decap_8 FILLER_25_2516 ();
 sg13g2_decap_8 FILLER_25_2523 ();
 sg13g2_decap_8 FILLER_25_2530 ();
 sg13g2_decap_8 FILLER_25_2537 ();
 sg13g2_decap_8 FILLER_25_2544 ();
 sg13g2_decap_8 FILLER_25_2551 ();
 sg13g2_decap_8 FILLER_25_2558 ();
 sg13g2_decap_8 FILLER_25_2565 ();
 sg13g2_decap_8 FILLER_25_2572 ();
 sg13g2_decap_8 FILLER_25_2579 ();
 sg13g2_decap_8 FILLER_25_2586 ();
 sg13g2_decap_8 FILLER_25_2593 ();
 sg13g2_decap_8 FILLER_25_2600 ();
 sg13g2_decap_8 FILLER_25_2607 ();
 sg13g2_decap_8 FILLER_25_2614 ();
 sg13g2_decap_8 FILLER_25_2621 ();
 sg13g2_decap_8 FILLER_25_2628 ();
 sg13g2_decap_8 FILLER_25_2635 ();
 sg13g2_decap_8 FILLER_25_2642 ();
 sg13g2_decap_8 FILLER_25_2649 ();
 sg13g2_decap_8 FILLER_25_2656 ();
 sg13g2_decap_8 FILLER_25_2663 ();
 sg13g2_decap_4 FILLER_25_2670 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_fill_2 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_100 ();
 sg13g2_fill_1 FILLER_26_131 ();
 sg13g2_fill_1 FILLER_26_146 ();
 sg13g2_fill_1 FILLER_26_165 ();
 sg13g2_fill_1 FILLER_26_206 ();
 sg13g2_fill_1 FILLER_26_233 ();
 sg13g2_fill_2 FILLER_26_258 ();
 sg13g2_fill_2 FILLER_26_293 ();
 sg13g2_fill_1 FILLER_26_295 ();
 sg13g2_decap_8 FILLER_26_311 ();
 sg13g2_decap_4 FILLER_26_318 ();
 sg13g2_fill_2 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_fill_1 FILLER_26_399 ();
 sg13g2_fill_1 FILLER_26_404 ();
 sg13g2_fill_2 FILLER_26_423 ();
 sg13g2_decap_8 FILLER_26_455 ();
 sg13g2_decap_4 FILLER_26_462 ();
 sg13g2_fill_1 FILLER_26_470 ();
 sg13g2_fill_2 FILLER_26_476 ();
 sg13g2_fill_1 FILLER_26_478 ();
 sg13g2_decap_4 FILLER_26_487 ();
 sg13g2_fill_1 FILLER_26_499 ();
 sg13g2_fill_2 FILLER_26_505 ();
 sg13g2_decap_4 FILLER_26_516 ();
 sg13g2_fill_1 FILLER_26_546 ();
 sg13g2_fill_2 FILLER_26_589 ();
 sg13g2_fill_1 FILLER_26_591 ();
 sg13g2_fill_2 FILLER_26_639 ();
 sg13g2_fill_2 FILLER_26_652 ();
 sg13g2_fill_1 FILLER_26_654 ();
 sg13g2_fill_1 FILLER_26_664 ();
 sg13g2_fill_2 FILLER_26_679 ();
 sg13g2_fill_1 FILLER_26_698 ();
 sg13g2_fill_1 FILLER_26_707 ();
 sg13g2_fill_2 FILLER_26_716 ();
 sg13g2_fill_1 FILLER_26_718 ();
 sg13g2_fill_1 FILLER_26_725 ();
 sg13g2_fill_2 FILLER_26_744 ();
 sg13g2_fill_1 FILLER_26_746 ();
 sg13g2_fill_2 FILLER_26_790 ();
 sg13g2_fill_1 FILLER_26_818 ();
 sg13g2_decap_8 FILLER_26_832 ();
 sg13g2_fill_2 FILLER_26_839 ();
 sg13g2_fill_1 FILLER_26_841 ();
 sg13g2_fill_2 FILLER_26_880 ();
 sg13g2_fill_2 FILLER_26_886 ();
 sg13g2_fill_2 FILLER_26_915 ();
 sg13g2_fill_2 FILLER_26_922 ();
 sg13g2_fill_1 FILLER_26_1159 ();
 sg13g2_fill_2 FILLER_26_1219 ();
 sg13g2_fill_2 FILLER_26_1267 ();
 sg13g2_fill_1 FILLER_26_1336 ();
 sg13g2_fill_1 FILLER_26_1523 ();
 sg13g2_fill_1 FILLER_26_1583 ();
 sg13g2_fill_2 FILLER_26_1593 ();
 sg13g2_fill_1 FILLER_26_1626 ();
 sg13g2_fill_1 FILLER_26_1664 ();
 sg13g2_fill_1 FILLER_26_1679 ();
 sg13g2_fill_2 FILLER_26_1741 ();
 sg13g2_fill_2 FILLER_26_1752 ();
 sg13g2_decap_4 FILLER_26_1814 ();
 sg13g2_decap_8 FILLER_26_1831 ();
 sg13g2_fill_2 FILLER_26_1838 ();
 sg13g2_decap_4 FILLER_26_1928 ();
 sg13g2_fill_1 FILLER_26_1932 ();
 sg13g2_fill_2 FILLER_26_1957 ();
 sg13g2_decap_8 FILLER_26_1963 ();
 sg13g2_fill_2 FILLER_26_1975 ();
 sg13g2_fill_2 FILLER_26_1991 ();
 sg13g2_fill_2 FILLER_26_1998 ();
 sg13g2_fill_1 FILLER_26_2000 ();
 sg13g2_decap_4 FILLER_26_2018 ();
 sg13g2_decap_4 FILLER_26_2032 ();
 sg13g2_fill_2 FILLER_26_2087 ();
 sg13g2_fill_1 FILLER_26_2089 ();
 sg13g2_fill_2 FILLER_26_2106 ();
 sg13g2_fill_1 FILLER_26_2108 ();
 sg13g2_decap_4 FILLER_26_2202 ();
 sg13g2_fill_2 FILLER_26_2206 ();
 sg13g2_fill_1 FILLER_26_2221 ();
 sg13g2_fill_2 FILLER_26_2231 ();
 sg13g2_fill_1 FILLER_26_2233 ();
 sg13g2_fill_1 FILLER_26_2260 ();
 sg13g2_fill_2 FILLER_26_2309 ();
 sg13g2_fill_1 FILLER_26_2311 ();
 sg13g2_decap_8 FILLER_26_2338 ();
 sg13g2_decap_8 FILLER_26_2345 ();
 sg13g2_decap_8 FILLER_26_2352 ();
 sg13g2_decap_8 FILLER_26_2359 ();
 sg13g2_decap_8 FILLER_26_2366 ();
 sg13g2_decap_8 FILLER_26_2373 ();
 sg13g2_decap_8 FILLER_26_2380 ();
 sg13g2_decap_8 FILLER_26_2387 ();
 sg13g2_decap_8 FILLER_26_2394 ();
 sg13g2_decap_8 FILLER_26_2401 ();
 sg13g2_decap_8 FILLER_26_2408 ();
 sg13g2_decap_8 FILLER_26_2415 ();
 sg13g2_decap_8 FILLER_26_2422 ();
 sg13g2_decap_8 FILLER_26_2429 ();
 sg13g2_decap_8 FILLER_26_2436 ();
 sg13g2_decap_8 FILLER_26_2443 ();
 sg13g2_decap_8 FILLER_26_2450 ();
 sg13g2_decap_8 FILLER_26_2457 ();
 sg13g2_decap_8 FILLER_26_2464 ();
 sg13g2_decap_8 FILLER_26_2471 ();
 sg13g2_decap_8 FILLER_26_2478 ();
 sg13g2_decap_8 FILLER_26_2485 ();
 sg13g2_decap_8 FILLER_26_2492 ();
 sg13g2_decap_8 FILLER_26_2499 ();
 sg13g2_decap_8 FILLER_26_2506 ();
 sg13g2_decap_8 FILLER_26_2513 ();
 sg13g2_decap_8 FILLER_26_2520 ();
 sg13g2_decap_8 FILLER_26_2527 ();
 sg13g2_decap_8 FILLER_26_2534 ();
 sg13g2_decap_8 FILLER_26_2541 ();
 sg13g2_decap_8 FILLER_26_2548 ();
 sg13g2_decap_8 FILLER_26_2555 ();
 sg13g2_decap_8 FILLER_26_2562 ();
 sg13g2_decap_8 FILLER_26_2569 ();
 sg13g2_decap_8 FILLER_26_2576 ();
 sg13g2_decap_8 FILLER_26_2583 ();
 sg13g2_decap_8 FILLER_26_2590 ();
 sg13g2_decap_8 FILLER_26_2597 ();
 sg13g2_decap_8 FILLER_26_2604 ();
 sg13g2_decap_8 FILLER_26_2611 ();
 sg13g2_decap_8 FILLER_26_2618 ();
 sg13g2_decap_8 FILLER_26_2625 ();
 sg13g2_decap_8 FILLER_26_2632 ();
 sg13g2_decap_8 FILLER_26_2639 ();
 sg13g2_decap_8 FILLER_26_2646 ();
 sg13g2_decap_8 FILLER_26_2653 ();
 sg13g2_decap_8 FILLER_26_2660 ();
 sg13g2_decap_8 FILLER_26_2667 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_fill_2 FILLER_27_112 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_fill_2 FILLER_27_119 ();
 sg13g2_fill_1 FILLER_27_165 ();
 sg13g2_fill_1 FILLER_27_190 ();
 sg13g2_decap_4 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_235 ();
 sg13g2_decap_8 FILLER_27_250 ();
 sg13g2_fill_2 FILLER_27_257 ();
 sg13g2_fill_2 FILLER_27_263 ();
 sg13g2_fill_1 FILLER_27_265 ();
 sg13g2_fill_2 FILLER_27_270 ();
 sg13g2_fill_1 FILLER_27_281 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_318 ();
 sg13g2_decap_4 FILLER_27_327 ();
 sg13g2_decap_8 FILLER_27_339 ();
 sg13g2_fill_2 FILLER_27_346 ();
 sg13g2_decap_4 FILLER_27_354 ();
 sg13g2_fill_1 FILLER_27_358 ();
 sg13g2_fill_1 FILLER_27_388 ();
 sg13g2_decap_4 FILLER_27_481 ();
 sg13g2_fill_1 FILLER_27_485 ();
 sg13g2_fill_2 FILLER_27_520 ();
 sg13g2_fill_1 FILLER_27_522 ();
 sg13g2_decap_4 FILLER_27_531 ();
 sg13g2_fill_2 FILLER_27_551 ();
 sg13g2_fill_1 FILLER_27_574 ();
 sg13g2_fill_2 FILLER_27_648 ();
 sg13g2_fill_1 FILLER_27_650 ();
 sg13g2_fill_1 FILLER_27_666 ();
 sg13g2_fill_2 FILLER_27_718 ();
 sg13g2_fill_1 FILLER_27_720 ();
 sg13g2_decap_8 FILLER_27_775 ();
 sg13g2_decap_8 FILLER_27_782 ();
 sg13g2_fill_2 FILLER_27_789 ();
 sg13g2_fill_1 FILLER_27_791 ();
 sg13g2_fill_2 FILLER_27_800 ();
 sg13g2_fill_1 FILLER_27_802 ();
 sg13g2_fill_1 FILLER_27_818 ();
 sg13g2_fill_1 FILLER_27_824 ();
 sg13g2_fill_2 FILLER_27_854 ();
 sg13g2_fill_1 FILLER_27_856 ();
 sg13g2_fill_1 FILLER_27_1085 ();
 sg13g2_fill_2 FILLER_27_1189 ();
 sg13g2_fill_2 FILLER_27_1221 ();
 sg13g2_fill_1 FILLER_27_1228 ();
 sg13g2_fill_1 FILLER_27_1289 ();
 sg13g2_fill_2 FILLER_27_1313 ();
 sg13g2_decap_8 FILLER_27_1340 ();
 sg13g2_decap_4 FILLER_27_1347 ();
 sg13g2_fill_1 FILLER_27_1399 ();
 sg13g2_fill_1 FILLER_27_1498 ();
 sg13g2_fill_1 FILLER_27_1559 ();
 sg13g2_fill_1 FILLER_27_1642 ();
 sg13g2_fill_2 FILLER_27_1680 ();
 sg13g2_fill_1 FILLER_27_1710 ();
 sg13g2_fill_2 FILLER_27_1788 ();
 sg13g2_fill_2 FILLER_27_1795 ();
 sg13g2_fill_1 FILLER_27_1797 ();
 sg13g2_decap_4 FILLER_27_1840 ();
 sg13g2_fill_1 FILLER_27_1880 ();
 sg13g2_fill_2 FILLER_27_1886 ();
 sg13g2_fill_1 FILLER_27_1897 ();
 sg13g2_fill_2 FILLER_27_1911 ();
 sg13g2_fill_2 FILLER_27_1938 ();
 sg13g2_fill_1 FILLER_27_1940 ();
 sg13g2_fill_2 FILLER_27_2048 ();
 sg13g2_fill_1 FILLER_27_2050 ();
 sg13g2_fill_2 FILLER_27_2082 ();
 sg13g2_fill_1 FILLER_27_2089 ();
 sg13g2_fill_2 FILLER_27_2105 ();
 sg13g2_fill_1 FILLER_27_2107 ();
 sg13g2_fill_1 FILLER_27_2144 ();
 sg13g2_fill_1 FILLER_27_2149 ();
 sg13g2_fill_1 FILLER_27_2189 ();
 sg13g2_fill_2 FILLER_27_2275 ();
 sg13g2_fill_1 FILLER_27_2277 ();
 sg13g2_fill_2 FILLER_27_2313 ();
 sg13g2_fill_2 FILLER_27_2333 ();
 sg13g2_decap_8 FILLER_27_2348 ();
 sg13g2_decap_8 FILLER_27_2355 ();
 sg13g2_decap_8 FILLER_27_2362 ();
 sg13g2_decap_8 FILLER_27_2369 ();
 sg13g2_decap_8 FILLER_27_2376 ();
 sg13g2_decap_8 FILLER_27_2383 ();
 sg13g2_decap_8 FILLER_27_2390 ();
 sg13g2_decap_8 FILLER_27_2397 ();
 sg13g2_decap_8 FILLER_27_2404 ();
 sg13g2_decap_8 FILLER_27_2411 ();
 sg13g2_decap_8 FILLER_27_2418 ();
 sg13g2_decap_8 FILLER_27_2425 ();
 sg13g2_decap_8 FILLER_27_2432 ();
 sg13g2_decap_8 FILLER_27_2439 ();
 sg13g2_decap_8 FILLER_27_2446 ();
 sg13g2_decap_8 FILLER_27_2453 ();
 sg13g2_decap_8 FILLER_27_2460 ();
 sg13g2_decap_8 FILLER_27_2467 ();
 sg13g2_decap_8 FILLER_27_2474 ();
 sg13g2_decap_8 FILLER_27_2481 ();
 sg13g2_decap_8 FILLER_27_2488 ();
 sg13g2_decap_8 FILLER_27_2495 ();
 sg13g2_decap_8 FILLER_27_2502 ();
 sg13g2_decap_8 FILLER_27_2509 ();
 sg13g2_decap_8 FILLER_27_2516 ();
 sg13g2_decap_8 FILLER_27_2523 ();
 sg13g2_decap_8 FILLER_27_2530 ();
 sg13g2_decap_8 FILLER_27_2537 ();
 sg13g2_decap_8 FILLER_27_2544 ();
 sg13g2_decap_8 FILLER_27_2551 ();
 sg13g2_decap_8 FILLER_27_2558 ();
 sg13g2_decap_8 FILLER_27_2565 ();
 sg13g2_decap_8 FILLER_27_2572 ();
 sg13g2_decap_8 FILLER_27_2579 ();
 sg13g2_decap_8 FILLER_27_2586 ();
 sg13g2_decap_8 FILLER_27_2593 ();
 sg13g2_decap_8 FILLER_27_2600 ();
 sg13g2_decap_8 FILLER_27_2607 ();
 sg13g2_decap_8 FILLER_27_2614 ();
 sg13g2_decap_8 FILLER_27_2621 ();
 sg13g2_decap_8 FILLER_27_2628 ();
 sg13g2_decap_8 FILLER_27_2635 ();
 sg13g2_decap_8 FILLER_27_2642 ();
 sg13g2_decap_8 FILLER_27_2649 ();
 sg13g2_decap_8 FILLER_27_2656 ();
 sg13g2_decap_8 FILLER_27_2663 ();
 sg13g2_decap_4 FILLER_27_2670 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_4 FILLER_28_105 ();
 sg13g2_fill_2 FILLER_28_109 ();
 sg13g2_fill_1 FILLER_28_137 ();
 sg13g2_fill_1 FILLER_28_143 ();
 sg13g2_fill_1 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_213 ();
 sg13g2_decap_4 FILLER_28_230 ();
 sg13g2_decap_8 FILLER_28_249 ();
 sg13g2_decap_4 FILLER_28_260 ();
 sg13g2_fill_1 FILLER_28_264 ();
 sg13g2_decap_4 FILLER_28_276 ();
 sg13g2_fill_2 FILLER_28_280 ();
 sg13g2_decap_4 FILLER_28_298 ();
 sg13g2_fill_1 FILLER_28_320 ();
 sg13g2_fill_1 FILLER_28_353 ();
 sg13g2_fill_2 FILLER_28_358 ();
 sg13g2_fill_2 FILLER_28_364 ();
 sg13g2_fill_2 FILLER_28_383 ();
 sg13g2_fill_2 FILLER_28_394 ();
 sg13g2_fill_1 FILLER_28_415 ();
 sg13g2_fill_2 FILLER_28_442 ();
 sg13g2_fill_1 FILLER_28_444 ();
 sg13g2_fill_2 FILLER_28_464 ();
 sg13g2_fill_1 FILLER_28_466 ();
 sg13g2_fill_1 FILLER_28_485 ();
 sg13g2_fill_2 FILLER_28_536 ();
 sg13g2_fill_2 FILLER_28_551 ();
 sg13g2_fill_1 FILLER_28_553 ();
 sg13g2_decap_8 FILLER_28_564 ();
 sg13g2_fill_2 FILLER_28_571 ();
 sg13g2_fill_1 FILLER_28_630 ();
 sg13g2_fill_2 FILLER_28_636 ();
 sg13g2_fill_1 FILLER_28_670 ();
 sg13g2_decap_4 FILLER_28_687 ();
 sg13g2_fill_2 FILLER_28_691 ();
 sg13g2_fill_1 FILLER_28_710 ();
 sg13g2_fill_2 FILLER_28_754 ();
 sg13g2_fill_1 FILLER_28_780 ();
 sg13g2_fill_1 FILLER_28_797 ();
 sg13g2_fill_2 FILLER_28_811 ();
 sg13g2_fill_1 FILLER_28_813 ();
 sg13g2_fill_2 FILLER_28_830 ();
 sg13g2_fill_1 FILLER_28_832 ();
 sg13g2_fill_2 FILLER_28_838 ();
 sg13g2_fill_2 FILLER_28_870 ();
 sg13g2_fill_1 FILLER_28_872 ();
 sg13g2_fill_1 FILLER_28_881 ();
 sg13g2_fill_2 FILLER_28_922 ();
 sg13g2_fill_2 FILLER_28_938 ();
 sg13g2_fill_1 FILLER_28_989 ();
 sg13g2_fill_1 FILLER_28_1030 ();
 sg13g2_fill_2 FILLER_28_1159 ();
 sg13g2_fill_1 FILLER_28_1173 ();
 sg13g2_fill_2 FILLER_28_1197 ();
 sg13g2_fill_1 FILLER_28_1204 ();
 sg13g2_fill_2 FILLER_28_1219 ();
 sg13g2_fill_1 FILLER_28_1247 ();
 sg13g2_fill_1 FILLER_28_1259 ();
 sg13g2_fill_1 FILLER_28_1299 ();
 sg13g2_decap_4 FILLER_28_1337 ();
 sg13g2_decap_4 FILLER_28_1349 ();
 sg13g2_fill_2 FILLER_28_1353 ();
 sg13g2_fill_2 FILLER_28_1424 ();
 sg13g2_fill_1 FILLER_28_1456 ();
 sg13g2_fill_1 FILLER_28_1610 ();
 sg13g2_fill_1 FILLER_28_1624 ();
 sg13g2_fill_2 FILLER_28_1628 ();
 sg13g2_fill_2 FILLER_28_1645 ();
 sg13g2_fill_1 FILLER_28_1750 ();
 sg13g2_fill_2 FILLER_28_1796 ();
 sg13g2_fill_2 FILLER_28_1809 ();
 sg13g2_fill_1 FILLER_28_1811 ();
 sg13g2_fill_1 FILLER_28_1825 ();
 sg13g2_fill_1 FILLER_28_1859 ();
 sg13g2_fill_2 FILLER_28_1881 ();
 sg13g2_decap_4 FILLER_28_1891 ();
 sg13g2_fill_1 FILLER_28_1895 ();
 sg13g2_decap_4 FILLER_28_1939 ();
 sg13g2_fill_1 FILLER_28_1943 ();
 sg13g2_fill_2 FILLER_28_1962 ();
 sg13g2_fill_1 FILLER_28_1964 ();
 sg13g2_fill_1 FILLER_28_1975 ();
 sg13g2_decap_8 FILLER_28_1992 ();
 sg13g2_fill_1 FILLER_28_1999 ();
 sg13g2_fill_2 FILLER_28_2008 ();
 sg13g2_fill_2 FILLER_28_2018 ();
 sg13g2_fill_1 FILLER_28_2038 ();
 sg13g2_fill_1 FILLER_28_2100 ();
 sg13g2_fill_2 FILLER_28_2114 ();
 sg13g2_fill_2 FILLER_28_2129 ();
 sg13g2_fill_1 FILLER_28_2131 ();
 sg13g2_fill_2 FILLER_28_2153 ();
 sg13g2_decap_4 FILLER_28_2251 ();
 sg13g2_fill_1 FILLER_28_2255 ();
 sg13g2_fill_2 FILLER_28_2295 ();
 sg13g2_fill_2 FILLER_28_2323 ();
 sg13g2_fill_1 FILLER_28_2325 ();
 sg13g2_decap_8 FILLER_28_2352 ();
 sg13g2_decap_8 FILLER_28_2359 ();
 sg13g2_decap_8 FILLER_28_2366 ();
 sg13g2_decap_8 FILLER_28_2373 ();
 sg13g2_decap_8 FILLER_28_2380 ();
 sg13g2_decap_8 FILLER_28_2387 ();
 sg13g2_decap_8 FILLER_28_2394 ();
 sg13g2_decap_8 FILLER_28_2401 ();
 sg13g2_decap_8 FILLER_28_2408 ();
 sg13g2_decap_8 FILLER_28_2415 ();
 sg13g2_decap_8 FILLER_28_2422 ();
 sg13g2_decap_8 FILLER_28_2429 ();
 sg13g2_decap_8 FILLER_28_2436 ();
 sg13g2_decap_8 FILLER_28_2443 ();
 sg13g2_decap_8 FILLER_28_2450 ();
 sg13g2_decap_8 FILLER_28_2457 ();
 sg13g2_decap_8 FILLER_28_2464 ();
 sg13g2_decap_8 FILLER_28_2471 ();
 sg13g2_decap_8 FILLER_28_2478 ();
 sg13g2_decap_8 FILLER_28_2485 ();
 sg13g2_decap_8 FILLER_28_2492 ();
 sg13g2_decap_8 FILLER_28_2499 ();
 sg13g2_decap_8 FILLER_28_2506 ();
 sg13g2_decap_8 FILLER_28_2513 ();
 sg13g2_decap_8 FILLER_28_2520 ();
 sg13g2_decap_8 FILLER_28_2527 ();
 sg13g2_decap_8 FILLER_28_2534 ();
 sg13g2_decap_8 FILLER_28_2541 ();
 sg13g2_decap_8 FILLER_28_2548 ();
 sg13g2_decap_8 FILLER_28_2555 ();
 sg13g2_decap_8 FILLER_28_2562 ();
 sg13g2_decap_8 FILLER_28_2569 ();
 sg13g2_decap_8 FILLER_28_2576 ();
 sg13g2_decap_8 FILLER_28_2583 ();
 sg13g2_decap_8 FILLER_28_2590 ();
 sg13g2_decap_8 FILLER_28_2597 ();
 sg13g2_decap_8 FILLER_28_2604 ();
 sg13g2_decap_8 FILLER_28_2611 ();
 sg13g2_decap_8 FILLER_28_2618 ();
 sg13g2_decap_8 FILLER_28_2625 ();
 sg13g2_decap_8 FILLER_28_2632 ();
 sg13g2_decap_8 FILLER_28_2639 ();
 sg13g2_decap_8 FILLER_28_2646 ();
 sg13g2_decap_8 FILLER_28_2653 ();
 sg13g2_decap_8 FILLER_28_2660 ();
 sg13g2_decap_8 FILLER_28_2667 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_4 FILLER_29_98 ();
 sg13g2_fill_1 FILLER_29_102 ();
 sg13g2_fill_1 FILLER_29_129 ();
 sg13g2_fill_2 FILLER_29_144 ();
 sg13g2_fill_2 FILLER_29_170 ();
 sg13g2_fill_2 FILLER_29_190 ();
 sg13g2_decap_8 FILLER_29_212 ();
 sg13g2_decap_4 FILLER_29_219 ();
 sg13g2_fill_1 FILLER_29_223 ();
 sg13g2_fill_1 FILLER_29_244 ();
 sg13g2_decap_8 FILLER_29_271 ();
 sg13g2_decap_8 FILLER_29_300 ();
 sg13g2_decap_4 FILLER_29_307 ();
 sg13g2_fill_1 FILLER_29_311 ();
 sg13g2_decap_8 FILLER_29_331 ();
 sg13g2_decap_8 FILLER_29_338 ();
 sg13g2_decap_4 FILLER_29_345 ();
 sg13g2_fill_1 FILLER_29_349 ();
 sg13g2_fill_2 FILLER_29_360 ();
 sg13g2_fill_1 FILLER_29_372 ();
 sg13g2_fill_2 FILLER_29_392 ();
 sg13g2_fill_1 FILLER_29_394 ();
 sg13g2_fill_1 FILLER_29_438 ();
 sg13g2_fill_1 FILLER_29_444 ();
 sg13g2_fill_1 FILLER_29_458 ();
 sg13g2_fill_1 FILLER_29_482 ();
 sg13g2_decap_4 FILLER_29_527 ();
 sg13g2_decap_4 FILLER_29_539 ();
 sg13g2_fill_1 FILLER_29_543 ();
 sg13g2_fill_2 FILLER_29_556 ();
 sg13g2_fill_1 FILLER_29_564 ();
 sg13g2_fill_1 FILLER_29_570 ();
 sg13g2_decap_8 FILLER_29_589 ();
 sg13g2_decap_4 FILLER_29_596 ();
 sg13g2_fill_1 FILLER_29_608 ();
 sg13g2_decap_4 FILLER_29_615 ();
 sg13g2_fill_1 FILLER_29_619 ();
 sg13g2_fill_2 FILLER_29_638 ();
 sg13g2_fill_1 FILLER_29_640 ();
 sg13g2_decap_4 FILLER_29_654 ();
 sg13g2_fill_2 FILLER_29_692 ();
 sg13g2_fill_2 FILLER_29_700 ();
 sg13g2_decap_4 FILLER_29_707 ();
 sg13g2_fill_2 FILLER_29_711 ();
 sg13g2_fill_2 FILLER_29_730 ();
 sg13g2_decap_8 FILLER_29_737 ();
 sg13g2_fill_2 FILLER_29_748 ();
 sg13g2_fill_1 FILLER_29_750 ();
 sg13g2_fill_1 FILLER_29_763 ();
 sg13g2_fill_2 FILLER_29_790 ();
 sg13g2_fill_1 FILLER_29_800 ();
 sg13g2_fill_2 FILLER_29_817 ();
 sg13g2_fill_1 FILLER_29_824 ();
 sg13g2_decap_8 FILLER_29_849 ();
 sg13g2_fill_1 FILLER_29_856 ();
 sg13g2_fill_2 FILLER_29_870 ();
 sg13g2_fill_1 FILLER_29_902 ();
 sg13g2_fill_1 FILLER_29_974 ();
 sg13g2_fill_1 FILLER_29_1006 ();
 sg13g2_fill_1 FILLER_29_1104 ();
 sg13g2_fill_2 FILLER_29_1167 ();
 sg13g2_fill_1 FILLER_29_1169 ();
 sg13g2_fill_1 FILLER_29_1192 ();
 sg13g2_fill_2 FILLER_29_1262 ();
 sg13g2_fill_1 FILLER_29_1272 ();
 sg13g2_fill_1 FILLER_29_1278 ();
 sg13g2_fill_1 FILLER_29_1284 ();
 sg13g2_fill_1 FILLER_29_1381 ();
 sg13g2_fill_1 FILLER_29_1591 ();
 sg13g2_fill_1 FILLER_29_1628 ();
 sg13g2_fill_1 FILLER_29_1651 ();
 sg13g2_fill_1 FILLER_29_1791 ();
 sg13g2_fill_2 FILLER_29_1816 ();
 sg13g2_fill_2 FILLER_29_1826 ();
 sg13g2_fill_1 FILLER_29_1828 ();
 sg13g2_decap_8 FILLER_29_1849 ();
 sg13g2_fill_2 FILLER_29_1856 ();
 sg13g2_fill_1 FILLER_29_1876 ();
 sg13g2_decap_8 FILLER_29_1881 ();
 sg13g2_decap_8 FILLER_29_1888 ();
 sg13g2_decap_4 FILLER_29_1895 ();
 sg13g2_fill_1 FILLER_29_1899 ();
 sg13g2_decap_8 FILLER_29_1917 ();
 sg13g2_decap_4 FILLER_29_1940 ();
 sg13g2_fill_2 FILLER_29_1944 ();
 sg13g2_decap_4 FILLER_29_1954 ();
 sg13g2_fill_2 FILLER_29_1958 ();
 sg13g2_fill_1 FILLER_29_1972 ();
 sg13g2_fill_2 FILLER_29_1977 ();
 sg13g2_fill_1 FILLER_29_1979 ();
 sg13g2_decap_4 FILLER_29_1993 ();
 sg13g2_fill_2 FILLER_29_2049 ();
 sg13g2_fill_2 FILLER_29_2094 ();
 sg13g2_fill_1 FILLER_29_2096 ();
 sg13g2_fill_2 FILLER_29_2136 ();
 sg13g2_fill_1 FILLER_29_2164 ();
 sg13g2_fill_1 FILLER_29_2171 ();
 sg13g2_fill_2 FILLER_29_2187 ();
 sg13g2_decap_4 FILLER_29_2199 ();
 sg13g2_fill_1 FILLER_29_2251 ();
 sg13g2_fill_1 FILLER_29_2256 ();
 sg13g2_fill_2 FILLER_29_2275 ();
 sg13g2_fill_1 FILLER_29_2277 ();
 sg13g2_fill_2 FILLER_29_2310 ();
 sg13g2_fill_1 FILLER_29_2322 ();
 sg13g2_decap_8 FILLER_29_2349 ();
 sg13g2_decap_8 FILLER_29_2356 ();
 sg13g2_decap_8 FILLER_29_2363 ();
 sg13g2_decap_8 FILLER_29_2370 ();
 sg13g2_decap_8 FILLER_29_2377 ();
 sg13g2_decap_8 FILLER_29_2384 ();
 sg13g2_decap_8 FILLER_29_2391 ();
 sg13g2_decap_8 FILLER_29_2398 ();
 sg13g2_decap_8 FILLER_29_2405 ();
 sg13g2_decap_8 FILLER_29_2412 ();
 sg13g2_decap_8 FILLER_29_2419 ();
 sg13g2_decap_8 FILLER_29_2426 ();
 sg13g2_decap_8 FILLER_29_2433 ();
 sg13g2_decap_8 FILLER_29_2440 ();
 sg13g2_decap_8 FILLER_29_2447 ();
 sg13g2_decap_8 FILLER_29_2454 ();
 sg13g2_decap_8 FILLER_29_2461 ();
 sg13g2_decap_8 FILLER_29_2468 ();
 sg13g2_decap_8 FILLER_29_2475 ();
 sg13g2_decap_8 FILLER_29_2482 ();
 sg13g2_decap_8 FILLER_29_2489 ();
 sg13g2_decap_8 FILLER_29_2496 ();
 sg13g2_decap_8 FILLER_29_2503 ();
 sg13g2_decap_8 FILLER_29_2510 ();
 sg13g2_decap_8 FILLER_29_2517 ();
 sg13g2_decap_8 FILLER_29_2524 ();
 sg13g2_decap_8 FILLER_29_2531 ();
 sg13g2_decap_8 FILLER_29_2538 ();
 sg13g2_decap_8 FILLER_29_2545 ();
 sg13g2_decap_8 FILLER_29_2552 ();
 sg13g2_decap_8 FILLER_29_2559 ();
 sg13g2_decap_8 FILLER_29_2566 ();
 sg13g2_decap_8 FILLER_29_2573 ();
 sg13g2_decap_8 FILLER_29_2580 ();
 sg13g2_decap_8 FILLER_29_2587 ();
 sg13g2_decap_8 FILLER_29_2594 ();
 sg13g2_decap_8 FILLER_29_2601 ();
 sg13g2_decap_8 FILLER_29_2608 ();
 sg13g2_decap_8 FILLER_29_2615 ();
 sg13g2_decap_8 FILLER_29_2622 ();
 sg13g2_decap_8 FILLER_29_2629 ();
 sg13g2_decap_8 FILLER_29_2636 ();
 sg13g2_decap_8 FILLER_29_2643 ();
 sg13g2_decap_8 FILLER_29_2650 ();
 sg13g2_decap_8 FILLER_29_2657 ();
 sg13g2_decap_8 FILLER_29_2664 ();
 sg13g2_fill_2 FILLER_29_2671 ();
 sg13g2_fill_1 FILLER_29_2673 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_4 FILLER_30_98 ();
 sg13g2_fill_2 FILLER_30_102 ();
 sg13g2_fill_2 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_118 ();
 sg13g2_fill_2 FILLER_30_138 ();
 sg13g2_fill_1 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_146 ();
 sg13g2_fill_2 FILLER_30_182 ();
 sg13g2_fill_1 FILLER_30_184 ();
 sg13g2_decap_4 FILLER_30_208 ();
 sg13g2_fill_2 FILLER_30_220 ();
 sg13g2_fill_2 FILLER_30_235 ();
 sg13g2_fill_2 FILLER_30_253 ();
 sg13g2_fill_1 FILLER_30_255 ();
 sg13g2_fill_1 FILLER_30_264 ();
 sg13g2_fill_2 FILLER_30_273 ();
 sg13g2_decap_4 FILLER_30_306 ();
 sg13g2_fill_2 FILLER_30_310 ();
 sg13g2_decap_8 FILLER_30_332 ();
 sg13g2_decap_8 FILLER_30_339 ();
 sg13g2_fill_1 FILLER_30_346 ();
 sg13g2_decap_8 FILLER_30_352 ();
 sg13g2_decap_8 FILLER_30_359 ();
 sg13g2_fill_1 FILLER_30_378 ();
 sg13g2_fill_1 FILLER_30_384 ();
 sg13g2_decap_4 FILLER_30_409 ();
 sg13g2_fill_2 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_419 ();
 sg13g2_fill_2 FILLER_30_426 ();
 sg13g2_decap_4 FILLER_30_436 ();
 sg13g2_fill_2 FILLER_30_453 ();
 sg13g2_fill_1 FILLER_30_455 ();
 sg13g2_fill_2 FILLER_30_485 ();
 sg13g2_fill_1 FILLER_30_487 ();
 sg13g2_fill_1 FILLER_30_506 ();
 sg13g2_decap_4 FILLER_30_519 ();
 sg13g2_fill_2 FILLER_30_528 ();
 sg13g2_fill_2 FILLER_30_539 ();
 sg13g2_fill_2 FILLER_30_564 ();
 sg13g2_fill_2 FILLER_30_572 ();
 sg13g2_fill_1 FILLER_30_574 ();
 sg13g2_decap_4 FILLER_30_586 ();
 sg13g2_decap_8 FILLER_30_601 ();
 sg13g2_fill_2 FILLER_30_608 ();
 sg13g2_fill_1 FILLER_30_660 ();
 sg13g2_fill_1 FILLER_30_666 ();
 sg13g2_fill_1 FILLER_30_693 ();
 sg13g2_fill_1 FILLER_30_699 ();
 sg13g2_decap_8 FILLER_30_704 ();
 sg13g2_fill_1 FILLER_30_711 ();
 sg13g2_fill_2 FILLER_30_720 ();
 sg13g2_fill_1 FILLER_30_722 ();
 sg13g2_fill_2 FILLER_30_729 ();
 sg13g2_fill_2 FILLER_30_741 ();
 sg13g2_fill_1 FILLER_30_743 ();
 sg13g2_fill_2 FILLER_30_750 ();
 sg13g2_fill_1 FILLER_30_752 ();
 sg13g2_fill_2 FILLER_30_769 ();
 sg13g2_fill_2 FILLER_30_775 ();
 sg13g2_fill_2 FILLER_30_789 ();
 sg13g2_fill_1 FILLER_30_791 ();
 sg13g2_fill_2 FILLER_30_810 ();
 sg13g2_fill_1 FILLER_30_825 ();
 sg13g2_fill_2 FILLER_30_834 ();
 sg13g2_fill_1 FILLER_30_875 ();
 sg13g2_fill_2 FILLER_30_884 ();
 sg13g2_fill_2 FILLER_30_927 ();
 sg13g2_fill_1 FILLER_30_994 ();
 sg13g2_fill_2 FILLER_30_1063 ();
 sg13g2_fill_2 FILLER_30_1096 ();
 sg13g2_fill_2 FILLER_30_1189 ();
 sg13g2_fill_2 FILLER_30_1223 ();
 sg13g2_fill_1 FILLER_30_1240 ();
 sg13g2_fill_1 FILLER_30_1311 ();
 sg13g2_fill_2 FILLER_30_1331 ();
 sg13g2_fill_2 FILLER_30_1342 ();
 sg13g2_fill_2 FILLER_30_1381 ();
 sg13g2_fill_1 FILLER_30_1440 ();
 sg13g2_fill_1 FILLER_30_1460 ();
 sg13g2_fill_2 FILLER_30_1528 ();
 sg13g2_fill_1 FILLER_30_1613 ();
 sg13g2_fill_1 FILLER_30_1660 ();
 sg13g2_fill_2 FILLER_30_1701 ();
 sg13g2_fill_2 FILLER_30_1748 ();
 sg13g2_fill_1 FILLER_30_1750 ();
 sg13g2_fill_1 FILLER_30_1755 ();
 sg13g2_fill_1 FILLER_30_1796 ();
 sg13g2_fill_1 FILLER_30_1855 ();
 sg13g2_decap_4 FILLER_30_1915 ();
 sg13g2_fill_2 FILLER_30_1919 ();
 sg13g2_decap_8 FILLER_30_1925 ();
 sg13g2_decap_8 FILLER_30_1958 ();
 sg13g2_fill_2 FILLER_30_1978 ();
 sg13g2_fill_1 FILLER_30_1980 ();
 sg13g2_decap_8 FILLER_30_2007 ();
 sg13g2_decap_8 FILLER_30_2014 ();
 sg13g2_decap_4 FILLER_30_2021 ();
 sg13g2_fill_1 FILLER_30_2025 ();
 sg13g2_fill_2 FILLER_30_2035 ();
 sg13g2_fill_2 FILLER_30_2050 ();
 sg13g2_fill_1 FILLER_30_2052 ();
 sg13g2_fill_2 FILLER_30_2079 ();
 sg13g2_fill_1 FILLER_30_2081 ();
 sg13g2_fill_2 FILLER_30_2109 ();
 sg13g2_fill_1 FILLER_30_2111 ();
 sg13g2_fill_2 FILLER_30_2145 ();
 sg13g2_fill_2 FILLER_30_2159 ();
 sg13g2_fill_1 FILLER_30_2161 ();
 sg13g2_fill_2 FILLER_30_2192 ();
 sg13g2_decap_4 FILLER_30_2229 ();
 sg13g2_fill_1 FILLER_30_2267 ();
 sg13g2_fill_2 FILLER_30_2329 ();
 sg13g2_fill_1 FILLER_30_2331 ();
 sg13g2_decap_8 FILLER_30_2345 ();
 sg13g2_decap_8 FILLER_30_2352 ();
 sg13g2_decap_8 FILLER_30_2359 ();
 sg13g2_decap_8 FILLER_30_2366 ();
 sg13g2_decap_8 FILLER_30_2373 ();
 sg13g2_decap_8 FILLER_30_2380 ();
 sg13g2_decap_8 FILLER_30_2387 ();
 sg13g2_decap_8 FILLER_30_2394 ();
 sg13g2_decap_8 FILLER_30_2401 ();
 sg13g2_decap_8 FILLER_30_2408 ();
 sg13g2_decap_8 FILLER_30_2415 ();
 sg13g2_decap_8 FILLER_30_2422 ();
 sg13g2_decap_8 FILLER_30_2429 ();
 sg13g2_decap_8 FILLER_30_2436 ();
 sg13g2_decap_8 FILLER_30_2443 ();
 sg13g2_decap_8 FILLER_30_2450 ();
 sg13g2_decap_8 FILLER_30_2457 ();
 sg13g2_decap_8 FILLER_30_2464 ();
 sg13g2_decap_8 FILLER_30_2471 ();
 sg13g2_decap_8 FILLER_30_2478 ();
 sg13g2_decap_8 FILLER_30_2485 ();
 sg13g2_decap_8 FILLER_30_2492 ();
 sg13g2_decap_8 FILLER_30_2499 ();
 sg13g2_decap_8 FILLER_30_2506 ();
 sg13g2_decap_8 FILLER_30_2513 ();
 sg13g2_decap_8 FILLER_30_2520 ();
 sg13g2_decap_8 FILLER_30_2527 ();
 sg13g2_decap_8 FILLER_30_2534 ();
 sg13g2_decap_8 FILLER_30_2541 ();
 sg13g2_decap_8 FILLER_30_2548 ();
 sg13g2_decap_8 FILLER_30_2555 ();
 sg13g2_decap_8 FILLER_30_2562 ();
 sg13g2_decap_8 FILLER_30_2569 ();
 sg13g2_decap_8 FILLER_30_2576 ();
 sg13g2_decap_8 FILLER_30_2583 ();
 sg13g2_decap_8 FILLER_30_2590 ();
 sg13g2_decap_8 FILLER_30_2597 ();
 sg13g2_decap_8 FILLER_30_2604 ();
 sg13g2_decap_8 FILLER_30_2611 ();
 sg13g2_decap_8 FILLER_30_2618 ();
 sg13g2_decap_8 FILLER_30_2625 ();
 sg13g2_decap_8 FILLER_30_2632 ();
 sg13g2_decap_8 FILLER_30_2639 ();
 sg13g2_decap_8 FILLER_30_2646 ();
 sg13g2_decap_8 FILLER_30_2653 ();
 sg13g2_decap_8 FILLER_30_2660 ();
 sg13g2_decap_8 FILLER_30_2667 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_4 FILLER_31_98 ();
 sg13g2_fill_1 FILLER_31_102 ();
 sg13g2_decap_4 FILLER_31_129 ();
 sg13g2_decap_4 FILLER_31_187 ();
 sg13g2_fill_1 FILLER_31_191 ();
 sg13g2_decap_4 FILLER_31_208 ();
 sg13g2_fill_1 FILLER_31_212 ();
 sg13g2_fill_1 FILLER_31_229 ();
 sg13g2_fill_1 FILLER_31_244 ();
 sg13g2_fill_1 FILLER_31_261 ();
 sg13g2_fill_2 FILLER_31_297 ();
 sg13g2_fill_2 FILLER_31_304 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_fill_2 FILLER_31_321 ();
 sg13g2_fill_1 FILLER_31_323 ();
 sg13g2_fill_2 FILLER_31_335 ();
 sg13g2_fill_1 FILLER_31_337 ();
 sg13g2_fill_2 FILLER_31_350 ();
 sg13g2_fill_1 FILLER_31_352 ();
 sg13g2_decap_4 FILLER_31_365 ();
 sg13g2_fill_2 FILLER_31_377 ();
 sg13g2_decap_4 FILLER_31_387 ();
 sg13g2_fill_2 FILLER_31_391 ();
 sg13g2_fill_2 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_403 ();
 sg13g2_fill_1 FILLER_31_430 ();
 sg13g2_decap_8 FILLER_31_452 ();
 sg13g2_fill_2 FILLER_31_473 ();
 sg13g2_fill_1 FILLER_31_480 ();
 sg13g2_decap_4 FILLER_31_507 ();
 sg13g2_fill_2 FILLER_31_511 ();
 sg13g2_decap_4 FILLER_31_521 ();
 sg13g2_fill_1 FILLER_31_525 ();
 sg13g2_decap_8 FILLER_31_542 ();
 sg13g2_decap_8 FILLER_31_566 ();
 sg13g2_decap_8 FILLER_31_573 ();
 sg13g2_decap_4 FILLER_31_580 ();
 sg13g2_fill_2 FILLER_31_584 ();
 sg13g2_fill_1 FILLER_31_614 ();
 sg13g2_decap_8 FILLER_31_631 ();
 sg13g2_fill_2 FILLER_31_638 ();
 sg13g2_decap_8 FILLER_31_656 ();
 sg13g2_fill_2 FILLER_31_671 ();
 sg13g2_fill_1 FILLER_31_673 ();
 sg13g2_fill_2 FILLER_31_682 ();
 sg13g2_fill_1 FILLER_31_684 ();
 sg13g2_decap_4 FILLER_31_693 ();
 sg13g2_fill_1 FILLER_31_697 ();
 sg13g2_decap_8 FILLER_31_728 ();
 sg13g2_fill_2 FILLER_31_735 ();
 sg13g2_fill_1 FILLER_31_737 ();
 sg13g2_fill_2 FILLER_31_754 ();
 sg13g2_fill_1 FILLER_31_756 ();
 sg13g2_decap_4 FILLER_31_771 ();
 sg13g2_fill_2 FILLER_31_778 ();
 sg13g2_fill_1 FILLER_31_806 ();
 sg13g2_decap_8 FILLER_31_833 ();
 sg13g2_decap_8 FILLER_31_840 ();
 sg13g2_decap_4 FILLER_31_847 ();
 sg13g2_decap_8 FILLER_31_855 ();
 sg13g2_fill_2 FILLER_31_862 ();
 sg13g2_fill_1 FILLER_31_869 ();
 sg13g2_fill_1 FILLER_31_888 ();
 sg13g2_fill_2 FILLER_31_920 ();
 sg13g2_fill_2 FILLER_31_1083 ();
 sg13g2_fill_1 FILLER_31_1194 ();
 sg13g2_fill_1 FILLER_31_1234 ();
 sg13g2_fill_1 FILLER_31_1292 ();
 sg13g2_fill_2 FILLER_31_1312 ();
 sg13g2_fill_1 FILLER_31_1506 ();
 sg13g2_fill_1 FILLER_31_1547 ();
 sg13g2_fill_2 FILLER_31_1557 ();
 sg13g2_fill_1 FILLER_31_1577 ();
 sg13g2_fill_1 FILLER_31_1665 ();
 sg13g2_fill_1 FILLER_31_1728 ();
 sg13g2_fill_2 FILLER_31_1823 ();
 sg13g2_decap_4 FILLER_31_1833 ();
 sg13g2_fill_2 FILLER_31_1837 ();
 sg13g2_fill_2 FILLER_31_1852 ();
 sg13g2_fill_1 FILLER_31_1854 ();
 sg13g2_fill_2 FILLER_31_1867 ();
 sg13g2_fill_1 FILLER_31_1869 ();
 sg13g2_decap_8 FILLER_31_1894 ();
 sg13g2_fill_2 FILLER_31_1901 ();
 sg13g2_fill_2 FILLER_31_1908 ();
 sg13g2_fill_2 FILLER_31_1936 ();
 sg13g2_fill_2 FILLER_31_1968 ();
 sg13g2_fill_1 FILLER_31_1970 ();
 sg13g2_decap_8 FILLER_31_2001 ();
 sg13g2_decap_4 FILLER_31_2012 ();
 sg13g2_fill_2 FILLER_31_2016 ();
 sg13g2_decap_4 FILLER_31_2057 ();
 sg13g2_fill_1 FILLER_31_2061 ();
 sg13g2_fill_2 FILLER_31_2076 ();
 sg13g2_fill_1 FILLER_31_2094 ();
 sg13g2_fill_1 FILLER_31_2112 ();
 sg13g2_fill_2 FILLER_31_2123 ();
 sg13g2_fill_1 FILLER_31_2125 ();
 sg13g2_fill_1 FILLER_31_2156 ();
 sg13g2_decap_8 FILLER_31_2186 ();
 sg13g2_decap_8 FILLER_31_2198 ();
 sg13g2_decap_4 FILLER_31_2234 ();
 sg13g2_decap_8 FILLER_31_2252 ();
 sg13g2_fill_2 FILLER_31_2300 ();
 sg13g2_fill_1 FILLER_31_2302 ();
 sg13g2_fill_2 FILLER_31_2323 ();
 sg13g2_decap_8 FILLER_31_2351 ();
 sg13g2_decap_8 FILLER_31_2358 ();
 sg13g2_decap_8 FILLER_31_2365 ();
 sg13g2_decap_8 FILLER_31_2372 ();
 sg13g2_decap_8 FILLER_31_2379 ();
 sg13g2_decap_8 FILLER_31_2386 ();
 sg13g2_decap_8 FILLER_31_2393 ();
 sg13g2_decap_8 FILLER_31_2400 ();
 sg13g2_decap_8 FILLER_31_2407 ();
 sg13g2_decap_8 FILLER_31_2414 ();
 sg13g2_decap_8 FILLER_31_2421 ();
 sg13g2_decap_8 FILLER_31_2428 ();
 sg13g2_decap_8 FILLER_31_2435 ();
 sg13g2_decap_8 FILLER_31_2442 ();
 sg13g2_decap_8 FILLER_31_2449 ();
 sg13g2_decap_8 FILLER_31_2456 ();
 sg13g2_decap_8 FILLER_31_2463 ();
 sg13g2_decap_8 FILLER_31_2470 ();
 sg13g2_decap_8 FILLER_31_2477 ();
 sg13g2_decap_8 FILLER_31_2484 ();
 sg13g2_decap_8 FILLER_31_2491 ();
 sg13g2_decap_8 FILLER_31_2498 ();
 sg13g2_decap_8 FILLER_31_2505 ();
 sg13g2_decap_8 FILLER_31_2512 ();
 sg13g2_decap_8 FILLER_31_2519 ();
 sg13g2_decap_8 FILLER_31_2526 ();
 sg13g2_decap_8 FILLER_31_2533 ();
 sg13g2_decap_8 FILLER_31_2540 ();
 sg13g2_decap_8 FILLER_31_2547 ();
 sg13g2_decap_8 FILLER_31_2554 ();
 sg13g2_decap_8 FILLER_31_2561 ();
 sg13g2_decap_8 FILLER_31_2568 ();
 sg13g2_decap_8 FILLER_31_2575 ();
 sg13g2_decap_8 FILLER_31_2582 ();
 sg13g2_decap_8 FILLER_31_2589 ();
 sg13g2_decap_8 FILLER_31_2596 ();
 sg13g2_decap_8 FILLER_31_2603 ();
 sg13g2_decap_8 FILLER_31_2610 ();
 sg13g2_decap_8 FILLER_31_2617 ();
 sg13g2_decap_8 FILLER_31_2624 ();
 sg13g2_decap_8 FILLER_31_2631 ();
 sg13g2_decap_8 FILLER_31_2638 ();
 sg13g2_decap_8 FILLER_31_2645 ();
 sg13g2_decap_8 FILLER_31_2652 ();
 sg13g2_decap_8 FILLER_31_2659 ();
 sg13g2_decap_8 FILLER_31_2666 ();
 sg13g2_fill_1 FILLER_31_2673 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_105 ();
 sg13g2_fill_1 FILLER_32_107 ();
 sg13g2_fill_2 FILLER_32_112 ();
 sg13g2_decap_4 FILLER_32_118 ();
 sg13g2_fill_2 FILLER_32_122 ();
 sg13g2_fill_1 FILLER_32_178 ();
 sg13g2_decap_8 FILLER_32_198 ();
 sg13g2_decap_4 FILLER_32_205 ();
 sg13g2_fill_1 FILLER_32_209 ();
 sg13g2_decap_8 FILLER_32_234 ();
 sg13g2_decap_8 FILLER_32_241 ();
 sg13g2_fill_1 FILLER_32_256 ();
 sg13g2_decap_8 FILLER_32_279 ();
 sg13g2_fill_1 FILLER_32_286 ();
 sg13g2_fill_2 FILLER_32_311 ();
 sg13g2_fill_1 FILLER_32_313 ();
 sg13g2_fill_1 FILLER_32_320 ();
 sg13g2_decap_4 FILLER_32_332 ();
 sg13g2_fill_1 FILLER_32_360 ();
 sg13g2_decap_4 FILLER_32_377 ();
 sg13g2_decap_4 FILLER_32_401 ();
 sg13g2_fill_2 FILLER_32_419 ();
 sg13g2_fill_1 FILLER_32_421 ();
 sg13g2_fill_2 FILLER_32_436 ();
 sg13g2_fill_1 FILLER_32_438 ();
 sg13g2_decap_8 FILLER_32_452 ();
 sg13g2_decap_8 FILLER_32_459 ();
 sg13g2_decap_4 FILLER_32_466 ();
 sg13g2_fill_1 FILLER_32_488 ();
 sg13g2_decap_4 FILLER_32_502 ();
 sg13g2_fill_1 FILLER_32_506 ();
 sg13g2_fill_1 FILLER_32_531 ();
 sg13g2_decap_8 FILLER_32_540 ();
 sg13g2_decap_8 FILLER_32_547 ();
 sg13g2_fill_1 FILLER_32_554 ();
 sg13g2_fill_2 FILLER_32_566 ();
 sg13g2_fill_2 FILLER_32_618 ();
 sg13g2_fill_1 FILLER_32_620 ();
 sg13g2_decap_4 FILLER_32_629 ();
 sg13g2_fill_1 FILLER_32_633 ();
 sg13g2_fill_2 FILLER_32_644 ();
 sg13g2_decap_8 FILLER_32_654 ();
 sg13g2_decap_8 FILLER_32_689 ();
 sg13g2_decap_4 FILLER_32_701 ();
 sg13g2_decap_8 FILLER_32_713 ();
 sg13g2_fill_2 FILLER_32_720 ();
 sg13g2_fill_2 FILLER_32_767 ();
 sg13g2_fill_1 FILLER_32_769 ();
 sg13g2_fill_1 FILLER_32_783 ();
 sg13g2_decap_4 FILLER_32_788 ();
 sg13g2_fill_2 FILLER_32_825 ();
 sg13g2_fill_1 FILLER_32_827 ();
 sg13g2_fill_2 FILLER_32_849 ();
 sg13g2_fill_1 FILLER_32_851 ();
 sg13g2_fill_1 FILLER_32_868 ();
 sg13g2_decap_8 FILLER_32_874 ();
 sg13g2_fill_1 FILLER_32_881 ();
 sg13g2_fill_1 FILLER_32_893 ();
 sg13g2_fill_1 FILLER_32_965 ();
 sg13g2_fill_1 FILLER_32_998 ();
 sg13g2_fill_2 FILLER_32_1038 ();
 sg13g2_fill_1 FILLER_32_1144 ();
 sg13g2_fill_1 FILLER_32_1220 ();
 sg13g2_fill_1 FILLER_32_1239 ();
 sg13g2_fill_2 FILLER_32_1275 ();
 sg13g2_fill_2 FILLER_32_1320 ();
 sg13g2_fill_1 FILLER_32_1363 ();
 sg13g2_fill_1 FILLER_32_1399 ();
 sg13g2_fill_1 FILLER_32_1405 ();
 sg13g2_fill_1 FILLER_32_1587 ();
 sg13g2_fill_1 FILLER_32_1614 ();
 sg13g2_fill_1 FILLER_32_1624 ();
 sg13g2_fill_2 FILLER_32_1643 ();
 sg13g2_fill_2 FILLER_32_1659 ();
 sg13g2_fill_2 FILLER_32_1705 ();
 sg13g2_fill_1 FILLER_32_1712 ();
 sg13g2_fill_2 FILLER_32_1758 ();
 sg13g2_decap_8 FILLER_32_1821 ();
 sg13g2_decap_8 FILLER_32_1828 ();
 sg13g2_decap_8 FILLER_32_1835 ();
 sg13g2_fill_1 FILLER_32_1842 ();
 sg13g2_decap_8 FILLER_32_1848 ();
 sg13g2_decap_4 FILLER_32_1855 ();
 sg13g2_decap_8 FILLER_32_1869 ();
 sg13g2_decap_4 FILLER_32_1876 ();
 sg13g2_fill_1 FILLER_32_1905 ();
 sg13g2_fill_1 FILLER_32_1919 ();
 sg13g2_decap_4 FILLER_32_1924 ();
 sg13g2_fill_1 FILLER_32_1928 ();
 sg13g2_decap_4 FILLER_32_1933 ();
 sg13g2_fill_2 FILLER_32_1937 ();
 sg13g2_decap_8 FILLER_32_1943 ();
 sg13g2_fill_2 FILLER_32_1950 ();
 sg13g2_fill_1 FILLER_32_1952 ();
 sg13g2_decap_4 FILLER_32_1957 ();
 sg13g2_fill_1 FILLER_32_1961 ();
 sg13g2_fill_1 FILLER_32_1975 ();
 sg13g2_fill_2 FILLER_32_2002 ();
 sg13g2_fill_1 FILLER_32_2004 ();
 sg13g2_decap_4 FILLER_32_2039 ();
 sg13g2_fill_2 FILLER_32_2043 ();
 sg13g2_decap_4 FILLER_32_2084 ();
 sg13g2_fill_1 FILLER_32_2088 ();
 sg13g2_fill_1 FILLER_32_2101 ();
 sg13g2_fill_1 FILLER_32_2106 ();
 sg13g2_fill_2 FILLER_32_2125 ();
 sg13g2_fill_2 FILLER_32_2221 ();
 sg13g2_fill_2 FILLER_32_2259 ();
 sg13g2_fill_2 FILLER_32_2292 ();
 sg13g2_fill_1 FILLER_32_2294 ();
 sg13g2_decap_8 FILLER_32_2356 ();
 sg13g2_decap_8 FILLER_32_2363 ();
 sg13g2_decap_8 FILLER_32_2370 ();
 sg13g2_decap_8 FILLER_32_2377 ();
 sg13g2_decap_8 FILLER_32_2384 ();
 sg13g2_decap_8 FILLER_32_2391 ();
 sg13g2_decap_8 FILLER_32_2398 ();
 sg13g2_decap_8 FILLER_32_2405 ();
 sg13g2_decap_8 FILLER_32_2412 ();
 sg13g2_decap_8 FILLER_32_2419 ();
 sg13g2_decap_8 FILLER_32_2426 ();
 sg13g2_decap_8 FILLER_32_2433 ();
 sg13g2_decap_8 FILLER_32_2440 ();
 sg13g2_decap_8 FILLER_32_2447 ();
 sg13g2_decap_8 FILLER_32_2454 ();
 sg13g2_decap_8 FILLER_32_2461 ();
 sg13g2_decap_8 FILLER_32_2468 ();
 sg13g2_decap_8 FILLER_32_2475 ();
 sg13g2_decap_8 FILLER_32_2482 ();
 sg13g2_decap_8 FILLER_32_2489 ();
 sg13g2_decap_8 FILLER_32_2496 ();
 sg13g2_decap_8 FILLER_32_2503 ();
 sg13g2_decap_8 FILLER_32_2510 ();
 sg13g2_decap_8 FILLER_32_2517 ();
 sg13g2_decap_8 FILLER_32_2524 ();
 sg13g2_decap_8 FILLER_32_2531 ();
 sg13g2_decap_8 FILLER_32_2538 ();
 sg13g2_decap_8 FILLER_32_2545 ();
 sg13g2_decap_8 FILLER_32_2552 ();
 sg13g2_decap_8 FILLER_32_2559 ();
 sg13g2_decap_8 FILLER_32_2566 ();
 sg13g2_decap_8 FILLER_32_2573 ();
 sg13g2_decap_8 FILLER_32_2580 ();
 sg13g2_decap_8 FILLER_32_2587 ();
 sg13g2_decap_8 FILLER_32_2594 ();
 sg13g2_decap_8 FILLER_32_2601 ();
 sg13g2_decap_8 FILLER_32_2608 ();
 sg13g2_decap_8 FILLER_32_2615 ();
 sg13g2_decap_8 FILLER_32_2622 ();
 sg13g2_decap_8 FILLER_32_2629 ();
 sg13g2_decap_8 FILLER_32_2636 ();
 sg13g2_decap_8 FILLER_32_2643 ();
 sg13g2_decap_8 FILLER_32_2650 ();
 sg13g2_decap_8 FILLER_32_2657 ();
 sg13g2_decap_8 FILLER_32_2664 ();
 sg13g2_fill_2 FILLER_32_2671 ();
 sg13g2_fill_1 FILLER_32_2673 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_4 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_102 ();
 sg13g2_fill_2 FILLER_33_130 ();
 sg13g2_fill_1 FILLER_33_132 ();
 sg13g2_decap_4 FILLER_33_164 ();
 sg13g2_fill_1 FILLER_33_177 ();
 sg13g2_decap_4 FILLER_33_186 ();
 sg13g2_decap_8 FILLER_33_207 ();
 sg13g2_fill_2 FILLER_33_214 ();
 sg13g2_fill_1 FILLER_33_216 ();
 sg13g2_decap_4 FILLER_33_242 ();
 sg13g2_fill_1 FILLER_33_246 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_decap_4 FILLER_33_280 ();
 sg13g2_fill_1 FILLER_33_284 ();
 sg13g2_fill_2 FILLER_33_297 ();
 sg13g2_fill_1 FILLER_33_299 ();
 sg13g2_decap_4 FILLER_33_320 ();
 sg13g2_decap_4 FILLER_33_340 ();
 sg13g2_fill_2 FILLER_33_344 ();
 sg13g2_decap_4 FILLER_33_371 ();
 sg13g2_fill_1 FILLER_33_375 ();
 sg13g2_fill_2 FILLER_33_384 ();
 sg13g2_fill_1 FILLER_33_386 ();
 sg13g2_fill_1 FILLER_33_395 ();
 sg13g2_fill_1 FILLER_33_413 ();
 sg13g2_fill_2 FILLER_33_419 ();
 sg13g2_decap_8 FILLER_33_449 ();
 sg13g2_decap_4 FILLER_33_456 ();
 sg13g2_fill_1 FILLER_33_460 ();
 sg13g2_fill_1 FILLER_33_479 ();
 sg13g2_decap_4 FILLER_33_492 ();
 sg13g2_fill_2 FILLER_33_496 ();
 sg13g2_fill_2 FILLER_33_528 ();
 sg13g2_decap_4 FILLER_33_544 ();
 sg13g2_fill_1 FILLER_33_583 ();
 sg13g2_fill_2 FILLER_33_589 ();
 sg13g2_fill_1 FILLER_33_591 ();
 sg13g2_fill_1 FILLER_33_606 ();
 sg13g2_decap_8 FILLER_33_612 ();
 sg13g2_fill_2 FILLER_33_619 ();
 sg13g2_fill_1 FILLER_33_621 ();
 sg13g2_decap_8 FILLER_33_647 ();
 sg13g2_fill_2 FILLER_33_654 ();
 sg13g2_fill_1 FILLER_33_656 ();
 sg13g2_fill_2 FILLER_33_667 ();
 sg13g2_fill_2 FILLER_33_674 ();
 sg13g2_fill_1 FILLER_33_688 ();
 sg13g2_decap_4 FILLER_33_715 ();
 sg13g2_fill_2 FILLER_33_729 ();
 sg13g2_fill_1 FILLER_33_731 ();
 sg13g2_fill_1 FILLER_33_749 ();
 sg13g2_fill_2 FILLER_33_758 ();
 sg13g2_fill_2 FILLER_33_767 ();
 sg13g2_fill_2 FILLER_33_786 ();
 sg13g2_decap_8 FILLER_33_808 ();
 sg13g2_fill_2 FILLER_33_815 ();
 sg13g2_decap_4 FILLER_33_822 ();
 sg13g2_fill_1 FILLER_33_826 ();
 sg13g2_fill_2 FILLER_33_844 ();
 sg13g2_fill_1 FILLER_33_953 ();
 sg13g2_fill_2 FILLER_33_1075 ();
 sg13g2_fill_2 FILLER_33_1101 ();
 sg13g2_fill_1 FILLER_33_1158 ();
 sg13g2_fill_2 FILLER_33_1198 ();
 sg13g2_fill_1 FILLER_33_1249 ();
 sg13g2_fill_1 FILLER_33_1290 ();
 sg13g2_fill_2 FILLER_33_1354 ();
 sg13g2_fill_2 FILLER_33_1385 ();
 sg13g2_fill_2 FILLER_33_1436 ();
 sg13g2_fill_2 FILLER_33_1607 ();
 sg13g2_fill_2 FILLER_33_1624 ();
 sg13g2_fill_1 FILLER_33_1720 ();
 sg13g2_fill_2 FILLER_33_1755 ();
 sg13g2_decap_8 FILLER_33_1787 ();
 sg13g2_decap_4 FILLER_33_1794 ();
 sg13g2_fill_2 FILLER_33_1798 ();
 sg13g2_decap_4 FILLER_33_1830 ();
 sg13g2_fill_2 FILLER_33_1834 ();
 sg13g2_fill_2 FILLER_33_1898 ();
 sg13g2_fill_1 FILLER_33_1900 ();
 sg13g2_fill_2 FILLER_33_1939 ();
 sg13g2_decap_8 FILLER_33_1957 ();
 sg13g2_fill_1 FILLER_33_1964 ();
 sg13g2_decap_4 FILLER_33_1978 ();
 sg13g2_decap_8 FILLER_33_2002 ();
 sg13g2_decap_8 FILLER_33_2009 ();
 sg13g2_decap_4 FILLER_33_2016 ();
 sg13g2_fill_1 FILLER_33_2020 ();
 sg13g2_fill_2 FILLER_33_2039 ();
 sg13g2_decap_8 FILLER_33_2054 ();
 sg13g2_decap_4 FILLER_33_2061 ();
 sg13g2_fill_2 FILLER_33_2073 ();
 sg13g2_decap_4 FILLER_33_2084 ();
 sg13g2_fill_1 FILLER_33_2088 ();
 sg13g2_fill_2 FILLER_33_2128 ();
 sg13g2_fill_2 FILLER_33_2143 ();
 sg13g2_fill_1 FILLER_33_2145 ();
 sg13g2_fill_2 FILLER_33_2159 ();
 sg13g2_fill_1 FILLER_33_2161 ();
 sg13g2_decap_4 FILLER_33_2200 ();
 sg13g2_fill_1 FILLER_33_2204 ();
 sg13g2_fill_2 FILLER_33_2209 ();
 sg13g2_fill_1 FILLER_33_2211 ();
 sg13g2_decap_8 FILLER_33_2221 ();
 sg13g2_decap_8 FILLER_33_2228 ();
 sg13g2_decap_4 FILLER_33_2235 ();
 sg13g2_decap_4 FILLER_33_2249 ();
 sg13g2_decap_8 FILLER_33_2258 ();
 sg13g2_fill_2 FILLER_33_2265 ();
 sg13g2_fill_2 FILLER_33_2292 ();
 sg13g2_fill_1 FILLER_33_2294 ();
 sg13g2_decap_8 FILLER_33_2317 ();
 sg13g2_decap_8 FILLER_33_2324 ();
 sg13g2_fill_1 FILLER_33_2331 ();
 sg13g2_decap_8 FILLER_33_2349 ();
 sg13g2_decap_8 FILLER_33_2356 ();
 sg13g2_decap_8 FILLER_33_2363 ();
 sg13g2_decap_8 FILLER_33_2370 ();
 sg13g2_decap_8 FILLER_33_2377 ();
 sg13g2_decap_8 FILLER_33_2384 ();
 sg13g2_decap_8 FILLER_33_2391 ();
 sg13g2_decap_8 FILLER_33_2398 ();
 sg13g2_decap_8 FILLER_33_2405 ();
 sg13g2_decap_8 FILLER_33_2412 ();
 sg13g2_decap_8 FILLER_33_2419 ();
 sg13g2_decap_8 FILLER_33_2426 ();
 sg13g2_decap_8 FILLER_33_2433 ();
 sg13g2_decap_8 FILLER_33_2440 ();
 sg13g2_decap_8 FILLER_33_2447 ();
 sg13g2_decap_8 FILLER_33_2454 ();
 sg13g2_decap_8 FILLER_33_2461 ();
 sg13g2_decap_8 FILLER_33_2468 ();
 sg13g2_decap_8 FILLER_33_2475 ();
 sg13g2_decap_8 FILLER_33_2482 ();
 sg13g2_decap_8 FILLER_33_2489 ();
 sg13g2_decap_8 FILLER_33_2496 ();
 sg13g2_decap_8 FILLER_33_2503 ();
 sg13g2_decap_8 FILLER_33_2510 ();
 sg13g2_decap_8 FILLER_33_2517 ();
 sg13g2_decap_8 FILLER_33_2524 ();
 sg13g2_decap_8 FILLER_33_2531 ();
 sg13g2_decap_8 FILLER_33_2538 ();
 sg13g2_decap_8 FILLER_33_2545 ();
 sg13g2_decap_8 FILLER_33_2552 ();
 sg13g2_decap_8 FILLER_33_2559 ();
 sg13g2_decap_8 FILLER_33_2566 ();
 sg13g2_decap_8 FILLER_33_2573 ();
 sg13g2_decap_8 FILLER_33_2580 ();
 sg13g2_decap_8 FILLER_33_2587 ();
 sg13g2_decap_8 FILLER_33_2594 ();
 sg13g2_decap_8 FILLER_33_2601 ();
 sg13g2_decap_8 FILLER_33_2608 ();
 sg13g2_decap_8 FILLER_33_2615 ();
 sg13g2_decap_8 FILLER_33_2622 ();
 sg13g2_decap_8 FILLER_33_2629 ();
 sg13g2_decap_8 FILLER_33_2636 ();
 sg13g2_decap_8 FILLER_33_2643 ();
 sg13g2_decap_8 FILLER_33_2650 ();
 sg13g2_decap_8 FILLER_33_2657 ();
 sg13g2_decap_8 FILLER_33_2664 ();
 sg13g2_fill_2 FILLER_33_2671 ();
 sg13g2_fill_1 FILLER_33_2673 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_fill_2 FILLER_34_112 ();
 sg13g2_fill_1 FILLER_34_114 ();
 sg13g2_decap_4 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_140 ();
 sg13g2_fill_1 FILLER_34_142 ();
 sg13g2_fill_2 FILLER_34_153 ();
 sg13g2_fill_1 FILLER_34_179 ();
 sg13g2_fill_1 FILLER_34_184 ();
 sg13g2_fill_2 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_decap_4 FILLER_34_201 ();
 sg13g2_fill_2 FILLER_34_221 ();
 sg13g2_fill_1 FILLER_34_223 ();
 sg13g2_fill_2 FILLER_34_237 ();
 sg13g2_fill_1 FILLER_34_267 ();
 sg13g2_decap_4 FILLER_34_294 ();
 sg13g2_fill_2 FILLER_34_316 ();
 sg13g2_decap_4 FILLER_34_330 ();
 sg13g2_decap_8 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_fill_2 FILLER_34_413 ();
 sg13g2_fill_1 FILLER_34_415 ();
 sg13g2_decap_4 FILLER_34_422 ();
 sg13g2_fill_1 FILLER_34_435 ();
 sg13g2_decap_4 FILLER_34_456 ();
 sg13g2_fill_2 FILLER_34_460 ();
 sg13g2_decap_8 FILLER_34_467 ();
 sg13g2_decap_4 FILLER_34_474 ();
 sg13g2_fill_2 FILLER_34_508 ();
 sg13g2_fill_1 FILLER_34_510 ();
 sg13g2_fill_2 FILLER_34_551 ();
 sg13g2_fill_1 FILLER_34_553 ();
 sg13g2_decap_8 FILLER_34_562 ();
 sg13g2_fill_2 FILLER_34_574 ();
 sg13g2_decap_4 FILLER_34_587 ();
 sg13g2_fill_2 FILLER_34_597 ();
 sg13g2_fill_1 FILLER_34_619 ();
 sg13g2_fill_2 FILLER_34_628 ();
 sg13g2_fill_1 FILLER_34_630 ();
 sg13g2_fill_2 FILLER_34_674 ();
 sg13g2_fill_1 FILLER_34_676 ();
 sg13g2_fill_2 FILLER_34_700 ();
 sg13g2_fill_1 FILLER_34_702 ();
 sg13g2_fill_2 FILLER_34_712 ();
 sg13g2_fill_1 FILLER_34_714 ();
 sg13g2_fill_2 FILLER_34_731 ();
 sg13g2_fill_2 FILLER_34_754 ();
 sg13g2_decap_4 FILLER_34_766 ();
 sg13g2_fill_2 FILLER_34_770 ();
 sg13g2_decap_8 FILLER_34_777 ();
 sg13g2_fill_2 FILLER_34_784 ();
 sg13g2_fill_1 FILLER_34_786 ();
 sg13g2_decap_8 FILLER_34_844 ();
 sg13g2_decap_8 FILLER_34_851 ();
 sg13g2_fill_1 FILLER_34_858 ();
 sg13g2_decap_8 FILLER_34_863 ();
 sg13g2_fill_2 FILLER_34_870 ();
 sg13g2_fill_1 FILLER_34_872 ();
 sg13g2_fill_1 FILLER_34_957 ();
 sg13g2_fill_2 FILLER_34_1043 ();
 sg13g2_fill_2 FILLER_34_1156 ();
 sg13g2_fill_1 FILLER_34_1227 ();
 sg13g2_fill_1 FILLER_34_1233 ();
 sg13g2_fill_1 FILLER_34_1291 ();
 sg13g2_fill_1 FILLER_34_1343 ();
 sg13g2_fill_2 FILLER_34_1453 ();
 sg13g2_fill_1 FILLER_34_1516 ();
 sg13g2_fill_1 FILLER_34_1543 ();
 sg13g2_fill_2 FILLER_34_1592 ();
 sg13g2_fill_2 FILLER_34_1620 ();
 sg13g2_fill_1 FILLER_34_1630 ();
 sg13g2_fill_1 FILLER_34_1693 ();
 sg13g2_decap_4 FILLER_34_1776 ();
 sg13g2_fill_1 FILLER_34_1810 ();
 sg13g2_fill_2 FILLER_34_1850 ();
 sg13g2_fill_1 FILLER_34_1852 ();
 sg13g2_fill_1 FILLER_34_1858 ();
 sg13g2_decap_8 FILLER_34_1867 ();
 sg13g2_decap_4 FILLER_34_1874 ();
 sg13g2_fill_2 FILLER_34_1878 ();
 sg13g2_fill_1 FILLER_34_1884 ();
 sg13g2_decap_8 FILLER_34_1894 ();
 sg13g2_fill_2 FILLER_34_1901 ();
 sg13g2_fill_1 FILLER_34_1903 ();
 sg13g2_decap_4 FILLER_34_1912 ();
 sg13g2_fill_2 FILLER_34_1916 ();
 sg13g2_decap_4 FILLER_34_1926 ();
 sg13g2_decap_8 FILLER_34_1934 ();
 sg13g2_fill_2 FILLER_34_1941 ();
 sg13g2_fill_1 FILLER_34_1957 ();
 sg13g2_fill_1 FILLER_34_1967 ();
 sg13g2_decap_8 FILLER_34_1989 ();
 sg13g2_decap_4 FILLER_34_1996 ();
 sg13g2_fill_1 FILLER_34_2000 ();
 sg13g2_fill_2 FILLER_34_2006 ();
 sg13g2_fill_1 FILLER_34_2008 ();
 sg13g2_fill_2 FILLER_34_2043 ();
 sg13g2_fill_1 FILLER_34_2045 ();
 sg13g2_decap_8 FILLER_34_2072 ();
 sg13g2_fill_2 FILLER_34_2079 ();
 sg13g2_fill_2 FILLER_34_2108 ();
 sg13g2_fill_2 FILLER_34_2155 ();
 sg13g2_fill_1 FILLER_34_2157 ();
 sg13g2_decap_8 FILLER_34_2183 ();
 sg13g2_decap_8 FILLER_34_2190 ();
 sg13g2_decap_8 FILLER_34_2197 ();
 sg13g2_fill_2 FILLER_34_2204 ();
 sg13g2_fill_1 FILLER_34_2272 ();
 sg13g2_decap_8 FILLER_34_2320 ();
 sg13g2_fill_1 FILLER_34_2327 ();
 sg13g2_decap_8 FILLER_34_2332 ();
 sg13g2_decap_8 FILLER_34_2339 ();
 sg13g2_decap_8 FILLER_34_2346 ();
 sg13g2_decap_8 FILLER_34_2353 ();
 sg13g2_decap_8 FILLER_34_2360 ();
 sg13g2_decap_8 FILLER_34_2367 ();
 sg13g2_decap_8 FILLER_34_2374 ();
 sg13g2_decap_8 FILLER_34_2381 ();
 sg13g2_decap_8 FILLER_34_2388 ();
 sg13g2_decap_8 FILLER_34_2395 ();
 sg13g2_decap_8 FILLER_34_2402 ();
 sg13g2_decap_8 FILLER_34_2409 ();
 sg13g2_decap_8 FILLER_34_2416 ();
 sg13g2_decap_8 FILLER_34_2423 ();
 sg13g2_decap_8 FILLER_34_2430 ();
 sg13g2_decap_8 FILLER_34_2437 ();
 sg13g2_decap_8 FILLER_34_2444 ();
 sg13g2_decap_8 FILLER_34_2451 ();
 sg13g2_decap_8 FILLER_34_2458 ();
 sg13g2_decap_8 FILLER_34_2465 ();
 sg13g2_decap_8 FILLER_34_2472 ();
 sg13g2_decap_8 FILLER_34_2479 ();
 sg13g2_decap_8 FILLER_34_2486 ();
 sg13g2_decap_8 FILLER_34_2493 ();
 sg13g2_decap_8 FILLER_34_2500 ();
 sg13g2_decap_8 FILLER_34_2507 ();
 sg13g2_decap_8 FILLER_34_2514 ();
 sg13g2_decap_8 FILLER_34_2521 ();
 sg13g2_decap_8 FILLER_34_2528 ();
 sg13g2_decap_8 FILLER_34_2535 ();
 sg13g2_decap_8 FILLER_34_2542 ();
 sg13g2_decap_8 FILLER_34_2549 ();
 sg13g2_decap_8 FILLER_34_2556 ();
 sg13g2_decap_8 FILLER_34_2563 ();
 sg13g2_decap_8 FILLER_34_2570 ();
 sg13g2_decap_8 FILLER_34_2577 ();
 sg13g2_decap_8 FILLER_34_2584 ();
 sg13g2_decap_8 FILLER_34_2591 ();
 sg13g2_decap_8 FILLER_34_2598 ();
 sg13g2_decap_8 FILLER_34_2605 ();
 sg13g2_decap_8 FILLER_34_2612 ();
 sg13g2_decap_8 FILLER_34_2619 ();
 sg13g2_decap_8 FILLER_34_2626 ();
 sg13g2_decap_8 FILLER_34_2633 ();
 sg13g2_decap_8 FILLER_34_2640 ();
 sg13g2_decap_8 FILLER_34_2647 ();
 sg13g2_decap_8 FILLER_34_2654 ();
 sg13g2_decap_8 FILLER_34_2661 ();
 sg13g2_decap_4 FILLER_34_2668 ();
 sg13g2_fill_2 FILLER_34_2672 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_4 FILLER_35_105 ();
 sg13g2_fill_2 FILLER_35_135 ();
 sg13g2_fill_1 FILLER_35_146 ();
 sg13g2_fill_1 FILLER_35_163 ();
 sg13g2_fill_2 FILLER_35_205 ();
 sg13g2_fill_2 FILLER_35_217 ();
 sg13g2_fill_1 FILLER_35_219 ();
 sg13g2_decap_4 FILLER_35_238 ();
 sg13g2_decap_4 FILLER_35_257 ();
 sg13g2_fill_2 FILLER_35_261 ();
 sg13g2_decap_8 FILLER_35_277 ();
 sg13g2_fill_1 FILLER_35_289 ();
 sg13g2_fill_1 FILLER_35_295 ();
 sg13g2_decap_8 FILLER_35_306 ();
 sg13g2_fill_2 FILLER_35_313 ();
 sg13g2_fill_2 FILLER_35_331 ();
 sg13g2_fill_1 FILLER_35_333 ();
 sg13g2_fill_2 FILLER_35_358 ();
 sg13g2_fill_1 FILLER_35_360 ();
 sg13g2_fill_2 FILLER_35_369 ();
 sg13g2_fill_1 FILLER_35_376 ();
 sg13g2_fill_2 FILLER_35_402 ();
 sg13g2_fill_2 FILLER_35_433 ();
 sg13g2_fill_2 FILLER_35_452 ();
 sg13g2_fill_2 FILLER_35_481 ();
 sg13g2_fill_1 FILLER_35_483 ();
 sg13g2_decap_8 FILLER_35_493 ();
 sg13g2_fill_1 FILLER_35_500 ();
 sg13g2_fill_1 FILLER_35_536 ();
 sg13g2_fill_1 FILLER_35_549 ();
 sg13g2_decap_4 FILLER_35_597 ();
 sg13g2_fill_2 FILLER_35_601 ();
 sg13g2_decap_4 FILLER_35_612 ();
 sg13g2_fill_2 FILLER_35_616 ();
 sg13g2_fill_1 FILLER_35_623 ();
 sg13g2_fill_2 FILLER_35_633 ();
 sg13g2_fill_1 FILLER_35_700 ();
 sg13g2_fill_2 FILLER_35_709 ();
 sg13g2_decap_4 FILLER_35_763 ();
 sg13g2_fill_2 FILLER_35_783 ();
 sg13g2_fill_1 FILLER_35_801 ();
 sg13g2_fill_1 FILLER_35_806 ();
 sg13g2_fill_2 FILLER_35_815 ();
 sg13g2_fill_2 FILLER_35_822 ();
 sg13g2_fill_1 FILLER_35_824 ();
 sg13g2_decap_8 FILLER_35_841 ();
 sg13g2_fill_2 FILLER_35_848 ();
 sg13g2_fill_1 FILLER_35_850 ();
 sg13g2_fill_2 FILLER_35_891 ();
 sg13g2_fill_1 FILLER_35_893 ();
 sg13g2_fill_1 FILLER_35_1071 ();
 sg13g2_fill_2 FILLER_35_1094 ();
 sg13g2_fill_2 FILLER_35_1102 ();
 sg13g2_fill_2 FILLER_35_1149 ();
 sg13g2_fill_1 FILLER_35_1187 ();
 sg13g2_fill_1 FILLER_35_1233 ();
 sg13g2_fill_2 FILLER_35_1286 ();
 sg13g2_fill_2 FILLER_35_1344 ();
 sg13g2_fill_1 FILLER_35_1394 ();
 sg13g2_fill_1 FILLER_35_1437 ();
 sg13g2_fill_1 FILLER_35_1447 ();
 sg13g2_fill_2 FILLER_35_1494 ();
 sg13g2_fill_2 FILLER_35_1508 ();
 sg13g2_fill_1 FILLER_35_1528 ();
 sg13g2_fill_1 FILLER_35_1538 ();
 sg13g2_fill_1 FILLER_35_1563 ();
 sg13g2_fill_1 FILLER_35_1595 ();
 sg13g2_fill_2 FILLER_35_1601 ();
 sg13g2_fill_1 FILLER_35_1603 ();
 sg13g2_decap_4 FILLER_35_1608 ();
 sg13g2_fill_1 FILLER_35_1612 ();
 sg13g2_fill_1 FILLER_35_1616 ();
 sg13g2_fill_1 FILLER_35_1636 ();
 sg13g2_fill_2 FILLER_35_1646 ();
 sg13g2_fill_2 FILLER_35_1660 ();
 sg13g2_fill_2 FILLER_35_1676 ();
 sg13g2_fill_2 FILLER_35_1721 ();
 sg13g2_decap_4 FILLER_35_1736 ();
 sg13g2_fill_2 FILLER_35_1766 ();
 sg13g2_decap_8 FILLER_35_1785 ();
 sg13g2_fill_2 FILLER_35_1792 ();
 sg13g2_fill_1 FILLER_35_1794 ();
 sg13g2_decap_8 FILLER_35_1799 ();
 sg13g2_fill_2 FILLER_35_1806 ();
 sg13g2_fill_1 FILLER_35_1871 ();
 sg13g2_decap_4 FILLER_35_1945 ();
 sg13g2_fill_1 FILLER_35_1949 ();
 sg13g2_fill_2 FILLER_35_1971 ();
 sg13g2_fill_1 FILLER_35_1973 ();
 sg13g2_fill_2 FILLER_35_2030 ();
 sg13g2_decap_8 FILLER_35_2041 ();
 sg13g2_fill_1 FILLER_35_2048 ();
 sg13g2_fill_2 FILLER_35_2054 ();
 sg13g2_fill_2 FILLER_35_2156 ();
 sg13g2_fill_2 FILLER_35_2209 ();
 sg13g2_fill_1 FILLER_35_2211 ();
 sg13g2_fill_2 FILLER_35_2225 ();
 sg13g2_fill_1 FILLER_35_2240 ();
 sg13g2_fill_2 FILLER_35_2254 ();
 sg13g2_decap_8 FILLER_35_2261 ();
 sg13g2_decap_4 FILLER_35_2298 ();
 sg13g2_fill_1 FILLER_35_2316 ();
 sg13g2_decap_8 FILLER_35_2343 ();
 sg13g2_decap_8 FILLER_35_2350 ();
 sg13g2_decap_8 FILLER_35_2357 ();
 sg13g2_decap_8 FILLER_35_2364 ();
 sg13g2_decap_8 FILLER_35_2371 ();
 sg13g2_decap_8 FILLER_35_2378 ();
 sg13g2_decap_8 FILLER_35_2385 ();
 sg13g2_decap_8 FILLER_35_2392 ();
 sg13g2_decap_8 FILLER_35_2399 ();
 sg13g2_decap_8 FILLER_35_2406 ();
 sg13g2_decap_8 FILLER_35_2413 ();
 sg13g2_decap_8 FILLER_35_2420 ();
 sg13g2_decap_8 FILLER_35_2427 ();
 sg13g2_decap_8 FILLER_35_2434 ();
 sg13g2_decap_8 FILLER_35_2441 ();
 sg13g2_decap_8 FILLER_35_2448 ();
 sg13g2_decap_8 FILLER_35_2455 ();
 sg13g2_decap_8 FILLER_35_2462 ();
 sg13g2_decap_8 FILLER_35_2469 ();
 sg13g2_decap_8 FILLER_35_2476 ();
 sg13g2_decap_8 FILLER_35_2483 ();
 sg13g2_decap_8 FILLER_35_2490 ();
 sg13g2_decap_8 FILLER_35_2497 ();
 sg13g2_decap_8 FILLER_35_2504 ();
 sg13g2_decap_8 FILLER_35_2511 ();
 sg13g2_decap_8 FILLER_35_2518 ();
 sg13g2_decap_8 FILLER_35_2525 ();
 sg13g2_decap_8 FILLER_35_2532 ();
 sg13g2_decap_8 FILLER_35_2539 ();
 sg13g2_decap_8 FILLER_35_2546 ();
 sg13g2_decap_8 FILLER_35_2553 ();
 sg13g2_decap_8 FILLER_35_2560 ();
 sg13g2_decap_8 FILLER_35_2567 ();
 sg13g2_decap_8 FILLER_35_2574 ();
 sg13g2_decap_8 FILLER_35_2581 ();
 sg13g2_decap_8 FILLER_35_2588 ();
 sg13g2_decap_8 FILLER_35_2595 ();
 sg13g2_decap_8 FILLER_35_2602 ();
 sg13g2_decap_8 FILLER_35_2609 ();
 sg13g2_decap_8 FILLER_35_2616 ();
 sg13g2_decap_8 FILLER_35_2623 ();
 sg13g2_decap_8 FILLER_35_2630 ();
 sg13g2_decap_8 FILLER_35_2637 ();
 sg13g2_decap_8 FILLER_35_2644 ();
 sg13g2_decap_8 FILLER_35_2651 ();
 sg13g2_decap_8 FILLER_35_2658 ();
 sg13g2_decap_8 FILLER_35_2665 ();
 sg13g2_fill_2 FILLER_35_2672 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_119 ();
 sg13g2_decap_4 FILLER_36_124 ();
 sg13g2_fill_1 FILLER_36_128 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_decap_4 FILLER_36_185 ();
 sg13g2_fill_1 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_195 ();
 sg13g2_fill_1 FILLER_36_228 ();
 sg13g2_fill_2 FILLER_36_248 ();
 sg13g2_fill_1 FILLER_36_250 ();
 sg13g2_decap_4 FILLER_36_259 ();
 sg13g2_fill_1 FILLER_36_263 ();
 sg13g2_decap_8 FILLER_36_277 ();
 sg13g2_fill_2 FILLER_36_284 ();
 sg13g2_fill_1 FILLER_36_286 ();
 sg13g2_decap_8 FILLER_36_303 ();
 sg13g2_fill_2 FILLER_36_310 ();
 sg13g2_decap_4 FILLER_36_320 ();
 sg13g2_fill_1 FILLER_36_324 ();
 sg13g2_decap_4 FILLER_36_329 ();
 sg13g2_fill_1 FILLER_36_333 ();
 sg13g2_decap_8 FILLER_36_338 ();
 sg13g2_decap_8 FILLER_36_345 ();
 sg13g2_fill_2 FILLER_36_352 ();
 sg13g2_fill_2 FILLER_36_360 ();
 sg13g2_fill_1 FILLER_36_388 ();
 sg13g2_fill_2 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_425 ();
 sg13g2_fill_2 FILLER_36_431 ();
 sg13g2_decap_8 FILLER_36_449 ();
 sg13g2_decap_4 FILLER_36_456 ();
 sg13g2_fill_1 FILLER_36_460 ();
 sg13g2_fill_2 FILLER_36_474 ();
 sg13g2_fill_1 FILLER_36_476 ();
 sg13g2_fill_2 FILLER_36_486 ();
 sg13g2_fill_1 FILLER_36_488 ();
 sg13g2_fill_2 FILLER_36_529 ();
 sg13g2_decap_4 FILLER_36_539 ();
 sg13g2_fill_1 FILLER_36_543 ();
 sg13g2_decap_4 FILLER_36_557 ();
 sg13g2_fill_2 FILLER_36_571 ();
 sg13g2_fill_1 FILLER_36_573 ();
 sg13g2_decap_8 FILLER_36_583 ();
 sg13g2_decap_4 FILLER_36_590 ();
 sg13g2_fill_1 FILLER_36_601 ();
 sg13g2_fill_2 FILLER_36_641 ();
 sg13g2_fill_1 FILLER_36_643 ();
 sg13g2_fill_2 FILLER_36_670 ();
 sg13g2_fill_1 FILLER_36_672 ();
 sg13g2_fill_2 FILLER_36_716 ();
 sg13g2_fill_1 FILLER_36_718 ();
 sg13g2_fill_2 FILLER_36_752 ();
 sg13g2_fill_1 FILLER_36_754 ();
 sg13g2_fill_2 FILLER_36_785 ();
 sg13g2_decap_8 FILLER_36_816 ();
 sg13g2_decap_8 FILLER_36_823 ();
 sg13g2_decap_4 FILLER_36_830 ();
 sg13g2_decap_8 FILLER_36_847 ();
 sg13g2_decap_4 FILLER_36_892 ();
 sg13g2_fill_1 FILLER_36_945 ();
 sg13g2_fill_2 FILLER_36_964 ();
 sg13g2_fill_2 FILLER_36_1022 ();
 sg13g2_fill_1 FILLER_36_1091 ();
 sg13g2_fill_1 FILLER_36_1138 ();
 sg13g2_fill_2 FILLER_36_1174 ();
 sg13g2_fill_2 FILLER_36_1202 ();
 sg13g2_fill_1 FILLER_36_1289 ();
 sg13g2_fill_2 FILLER_36_1358 ();
 sg13g2_fill_2 FILLER_36_1369 ();
 sg13g2_fill_1 FILLER_36_1477 ();
 sg13g2_fill_2 FILLER_36_1485 ();
 sg13g2_fill_1 FILLER_36_1487 ();
 sg13g2_decap_4 FILLER_36_1496 ();
 sg13g2_fill_2 FILLER_36_1500 ();
 sg13g2_fill_2 FILLER_36_1533 ();
 sg13g2_fill_2 FILLER_36_1583 ();
 sg13g2_decap_8 FILLER_36_1595 ();
 sg13g2_fill_2 FILLER_36_1611 ();
 sg13g2_fill_1 FILLER_36_1703 ();
 sg13g2_decap_8 FILLER_36_1764 ();
 sg13g2_fill_1 FILLER_36_1844 ();
 sg13g2_decap_4 FILLER_36_1849 ();
 sg13g2_fill_1 FILLER_36_1853 ();
 sg13g2_fill_2 FILLER_36_1866 ();
 sg13g2_decap_8 FILLER_36_1876 ();
 sg13g2_decap_4 FILLER_36_1883 ();
 sg13g2_fill_2 FILLER_36_1887 ();
 sg13g2_decap_4 FILLER_36_1897 ();
 sg13g2_decap_4 FILLER_36_1905 ();
 sg13g2_decap_8 FILLER_36_1917 ();
 sg13g2_fill_1 FILLER_36_1924 ();
 sg13g2_fill_1 FILLER_36_1946 ();
 sg13g2_decap_4 FILLER_36_1967 ();
 sg13g2_fill_2 FILLER_36_1971 ();
 sg13g2_fill_1 FILLER_36_1985 ();
 sg13g2_fill_1 FILLER_36_2007 ();
 sg13g2_decap_8 FILLER_36_2013 ();
 sg13g2_decap_8 FILLER_36_2020 ();
 sg13g2_fill_1 FILLER_36_2027 ();
 sg13g2_decap_8 FILLER_36_2048 ();
 sg13g2_decap_4 FILLER_36_2055 ();
 sg13g2_decap_8 FILLER_36_2063 ();
 sg13g2_fill_1 FILLER_36_2070 ();
 sg13g2_decap_8 FILLER_36_2075 ();
 sg13g2_decap_4 FILLER_36_2082 ();
 sg13g2_fill_2 FILLER_36_2086 ();
 sg13g2_decap_8 FILLER_36_2092 ();
 sg13g2_fill_2 FILLER_36_2146 ();
 sg13g2_fill_1 FILLER_36_2152 ();
 sg13g2_fill_2 FILLER_36_2157 ();
 sg13g2_fill_1 FILLER_36_2232 ();
 sg13g2_decap_4 FILLER_36_2268 ();
 sg13g2_fill_2 FILLER_36_2272 ();
 sg13g2_fill_2 FILLER_36_2297 ();
 sg13g2_decap_8 FILLER_36_2344 ();
 sg13g2_decap_8 FILLER_36_2351 ();
 sg13g2_decap_8 FILLER_36_2358 ();
 sg13g2_decap_8 FILLER_36_2365 ();
 sg13g2_decap_8 FILLER_36_2372 ();
 sg13g2_decap_8 FILLER_36_2379 ();
 sg13g2_decap_8 FILLER_36_2386 ();
 sg13g2_decap_8 FILLER_36_2393 ();
 sg13g2_decap_8 FILLER_36_2400 ();
 sg13g2_decap_8 FILLER_36_2407 ();
 sg13g2_decap_8 FILLER_36_2414 ();
 sg13g2_decap_8 FILLER_36_2421 ();
 sg13g2_decap_8 FILLER_36_2428 ();
 sg13g2_decap_8 FILLER_36_2435 ();
 sg13g2_decap_8 FILLER_36_2442 ();
 sg13g2_decap_8 FILLER_36_2449 ();
 sg13g2_decap_8 FILLER_36_2456 ();
 sg13g2_decap_8 FILLER_36_2463 ();
 sg13g2_decap_8 FILLER_36_2470 ();
 sg13g2_decap_8 FILLER_36_2477 ();
 sg13g2_decap_8 FILLER_36_2484 ();
 sg13g2_decap_8 FILLER_36_2491 ();
 sg13g2_decap_8 FILLER_36_2498 ();
 sg13g2_decap_8 FILLER_36_2505 ();
 sg13g2_decap_8 FILLER_36_2512 ();
 sg13g2_decap_8 FILLER_36_2519 ();
 sg13g2_decap_8 FILLER_36_2526 ();
 sg13g2_decap_8 FILLER_36_2533 ();
 sg13g2_decap_8 FILLER_36_2540 ();
 sg13g2_decap_8 FILLER_36_2547 ();
 sg13g2_decap_8 FILLER_36_2554 ();
 sg13g2_decap_8 FILLER_36_2561 ();
 sg13g2_decap_8 FILLER_36_2568 ();
 sg13g2_decap_8 FILLER_36_2575 ();
 sg13g2_decap_8 FILLER_36_2582 ();
 sg13g2_decap_8 FILLER_36_2589 ();
 sg13g2_decap_8 FILLER_36_2596 ();
 sg13g2_decap_8 FILLER_36_2603 ();
 sg13g2_decap_8 FILLER_36_2610 ();
 sg13g2_decap_8 FILLER_36_2617 ();
 sg13g2_decap_8 FILLER_36_2624 ();
 sg13g2_decap_8 FILLER_36_2631 ();
 sg13g2_decap_8 FILLER_36_2638 ();
 sg13g2_decap_8 FILLER_36_2645 ();
 sg13g2_decap_8 FILLER_36_2652 ();
 sg13g2_decap_8 FILLER_36_2659 ();
 sg13g2_decap_8 FILLER_36_2666 ();
 sg13g2_fill_1 FILLER_36_2673 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_119 ();
 sg13g2_fill_1 FILLER_37_133 ();
 sg13g2_fill_2 FILLER_37_139 ();
 sg13g2_fill_1 FILLER_37_141 ();
 sg13g2_fill_1 FILLER_37_160 ();
 sg13g2_fill_1 FILLER_37_185 ();
 sg13g2_decap_4 FILLER_37_207 ();
 sg13g2_fill_1 FILLER_37_211 ();
 sg13g2_decap_8 FILLER_37_216 ();
 sg13g2_fill_1 FILLER_37_223 ();
 sg13g2_decap_4 FILLER_37_237 ();
 sg13g2_fill_1 FILLER_37_241 ();
 sg13g2_fill_1 FILLER_37_287 ();
 sg13g2_decap_4 FILLER_37_296 ();
 sg13g2_fill_1 FILLER_37_300 ();
 sg13g2_fill_2 FILLER_37_322 ();
 sg13g2_decap_4 FILLER_37_350 ();
 sg13g2_decap_4 FILLER_37_367 ();
 sg13g2_fill_1 FILLER_37_381 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_fill_2 FILLER_37_449 ();
 sg13g2_fill_2 FILLER_37_465 ();
 sg13g2_fill_1 FILLER_37_467 ();
 sg13g2_fill_2 FILLER_37_494 ();
 sg13g2_fill_1 FILLER_37_496 ();
 sg13g2_fill_2 FILLER_37_520 ();
 sg13g2_fill_2 FILLER_37_572 ();
 sg13g2_fill_1 FILLER_37_574 ();
 sg13g2_fill_1 FILLER_37_597 ();
 sg13g2_decap_8 FILLER_37_614 ();
 sg13g2_decap_4 FILLER_37_621 ();
 sg13g2_fill_1 FILLER_37_625 ();
 sg13g2_fill_1 FILLER_37_638 ();
 sg13g2_fill_2 FILLER_37_683 ();
 sg13g2_fill_1 FILLER_37_685 ();
 sg13g2_decap_4 FILLER_37_700 ();
 sg13g2_fill_2 FILLER_37_704 ();
 sg13g2_decap_4 FILLER_37_714 ();
 sg13g2_fill_2 FILLER_37_727 ();
 sg13g2_fill_1 FILLER_37_735 ();
 sg13g2_fill_1 FILLER_37_796 ();
 sg13g2_fill_1 FILLER_37_848 ();
 sg13g2_fill_2 FILLER_37_857 ();
 sg13g2_fill_2 FILLER_37_885 ();
 sg13g2_fill_1 FILLER_37_887 ();
 sg13g2_fill_2 FILLER_37_1037 ();
 sg13g2_fill_1 FILLER_37_1094 ();
 sg13g2_fill_1 FILLER_37_1163 ();
 sg13g2_fill_2 FILLER_37_1182 ();
 sg13g2_fill_1 FILLER_37_1250 ();
 sg13g2_fill_1 FILLER_37_1354 ();
 sg13g2_fill_2 FILLER_37_1420 ();
 sg13g2_fill_1 FILLER_37_1510 ();
 sg13g2_fill_2 FILLER_37_1571 ();
 sg13g2_decap_8 FILLER_37_1587 ();
 sg13g2_decap_4 FILLER_37_1616 ();
 sg13g2_fill_1 FILLER_37_1620 ();
 sg13g2_fill_2 FILLER_37_1624 ();
 sg13g2_fill_2 FILLER_37_1649 ();
 sg13g2_fill_1 FILLER_37_1669 ();
 sg13g2_decap_8 FILLER_37_1699 ();
 sg13g2_fill_1 FILLER_37_1706 ();
 sg13g2_decap_4 FILLER_37_1733 ();
 sg13g2_fill_2 FILLER_37_1737 ();
 sg13g2_fill_2 FILLER_37_1756 ();
 sg13g2_fill_1 FILLER_37_1758 ();
 sg13g2_fill_2 FILLER_37_1777 ();
 sg13g2_fill_1 FILLER_37_1779 ();
 sg13g2_fill_2 FILLER_37_1785 ();
 sg13g2_decap_4 FILLER_37_1799 ();
 sg13g2_fill_1 FILLER_37_1803 ();
 sg13g2_decap_8 FILLER_37_1808 ();
 sg13g2_fill_2 FILLER_37_1815 ();
 sg13g2_fill_2 FILLER_37_1825 ();
 sg13g2_fill_1 FILLER_37_1827 ();
 sg13g2_decap_8 FILLER_37_1836 ();
 sg13g2_decap_8 FILLER_37_1843 ();
 sg13g2_decap_8 FILLER_37_1858 ();
 sg13g2_decap_4 FILLER_37_1873 ();
 sg13g2_fill_1 FILLER_37_1877 ();
 sg13g2_fill_2 FILLER_37_1910 ();
 sg13g2_fill_1 FILLER_37_1912 ();
 sg13g2_decap_4 FILLER_37_1929 ();
 sg13g2_fill_1 FILLER_37_1933 ();
 sg13g2_decap_4 FILLER_37_1942 ();
 sg13g2_fill_1 FILLER_37_1946 ();
 sg13g2_fill_2 FILLER_37_1963 ();
 sg13g2_fill_1 FILLER_37_1965 ();
 sg13g2_decap_4 FILLER_37_1982 ();
 sg13g2_fill_1 FILLER_37_1986 ();
 sg13g2_decap_4 FILLER_37_1995 ();
 sg13g2_fill_1 FILLER_37_1999 ();
 sg13g2_fill_2 FILLER_37_2029 ();
 sg13g2_fill_2 FILLER_37_2036 ();
 sg13g2_fill_2 FILLER_37_2046 ();
 sg13g2_fill_1 FILLER_37_2048 ();
 sg13g2_decap_8 FILLER_37_2075 ();
 sg13g2_decap_8 FILLER_37_2082 ();
 sg13g2_fill_2 FILLER_37_2089 ();
 sg13g2_fill_1 FILLER_37_2091 ();
 sg13g2_fill_2 FILLER_37_2139 ();
 sg13g2_fill_1 FILLER_37_2141 ();
 sg13g2_decap_8 FILLER_37_2198 ();
 sg13g2_decap_4 FILLER_37_2205 ();
 sg13g2_fill_2 FILLER_37_2213 ();
 sg13g2_fill_1 FILLER_37_2215 ();
 sg13g2_fill_2 FILLER_37_2252 ();
 sg13g2_fill_1 FILLER_37_2280 ();
 sg13g2_fill_2 FILLER_37_2307 ();
 sg13g2_fill_1 FILLER_37_2309 ();
 sg13g2_decap_8 FILLER_37_2337 ();
 sg13g2_decap_8 FILLER_37_2344 ();
 sg13g2_decap_8 FILLER_37_2351 ();
 sg13g2_decap_8 FILLER_37_2358 ();
 sg13g2_decap_8 FILLER_37_2365 ();
 sg13g2_decap_8 FILLER_37_2372 ();
 sg13g2_decap_8 FILLER_37_2379 ();
 sg13g2_decap_8 FILLER_37_2386 ();
 sg13g2_decap_8 FILLER_37_2393 ();
 sg13g2_decap_8 FILLER_37_2400 ();
 sg13g2_decap_8 FILLER_37_2407 ();
 sg13g2_decap_8 FILLER_37_2414 ();
 sg13g2_decap_8 FILLER_37_2421 ();
 sg13g2_decap_8 FILLER_37_2428 ();
 sg13g2_decap_8 FILLER_37_2435 ();
 sg13g2_decap_8 FILLER_37_2442 ();
 sg13g2_decap_8 FILLER_37_2449 ();
 sg13g2_decap_8 FILLER_37_2456 ();
 sg13g2_decap_8 FILLER_37_2463 ();
 sg13g2_decap_8 FILLER_37_2470 ();
 sg13g2_decap_8 FILLER_37_2477 ();
 sg13g2_decap_8 FILLER_37_2484 ();
 sg13g2_decap_8 FILLER_37_2491 ();
 sg13g2_decap_8 FILLER_37_2498 ();
 sg13g2_decap_8 FILLER_37_2505 ();
 sg13g2_decap_8 FILLER_37_2512 ();
 sg13g2_decap_8 FILLER_37_2519 ();
 sg13g2_decap_8 FILLER_37_2526 ();
 sg13g2_decap_8 FILLER_37_2533 ();
 sg13g2_decap_8 FILLER_37_2540 ();
 sg13g2_decap_8 FILLER_37_2547 ();
 sg13g2_decap_8 FILLER_37_2554 ();
 sg13g2_decap_8 FILLER_37_2561 ();
 sg13g2_decap_8 FILLER_37_2568 ();
 sg13g2_decap_8 FILLER_37_2575 ();
 sg13g2_decap_8 FILLER_37_2582 ();
 sg13g2_decap_8 FILLER_37_2589 ();
 sg13g2_decap_8 FILLER_37_2596 ();
 sg13g2_decap_8 FILLER_37_2603 ();
 sg13g2_decap_8 FILLER_37_2610 ();
 sg13g2_decap_8 FILLER_37_2617 ();
 sg13g2_decap_8 FILLER_37_2624 ();
 sg13g2_decap_8 FILLER_37_2631 ();
 sg13g2_decap_8 FILLER_37_2638 ();
 sg13g2_decap_8 FILLER_37_2645 ();
 sg13g2_decap_8 FILLER_37_2652 ();
 sg13g2_decap_8 FILLER_37_2659 ();
 sg13g2_decap_8 FILLER_37_2666 ();
 sg13g2_fill_1 FILLER_37_2673 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_fill_2 FILLER_38_98 ();
 sg13g2_fill_2 FILLER_38_152 ();
 sg13g2_fill_2 FILLER_38_168 ();
 sg13g2_fill_1 FILLER_38_170 ();
 sg13g2_fill_2 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_fill_1 FILLER_38_203 ();
 sg13g2_fill_2 FILLER_38_213 ();
 sg13g2_fill_1 FILLER_38_215 ();
 sg13g2_decap_4 FILLER_38_239 ();
 sg13g2_decap_4 FILLER_38_258 ();
 sg13g2_fill_1 FILLER_38_262 ();
 sg13g2_decap_8 FILLER_38_278 ();
 sg13g2_decap_4 FILLER_38_285 ();
 sg13g2_fill_2 FILLER_38_289 ();
 sg13g2_fill_2 FILLER_38_304 ();
 sg13g2_fill_2 FILLER_38_366 ();
 sg13g2_fill_1 FILLER_38_368 ();
 sg13g2_fill_2 FILLER_38_374 ();
 sg13g2_fill_1 FILLER_38_376 ();
 sg13g2_fill_1 FILLER_38_402 ();
 sg13g2_fill_1 FILLER_38_437 ();
 sg13g2_decap_4 FILLER_38_455 ();
 sg13g2_fill_1 FILLER_38_476 ();
 sg13g2_fill_2 FILLER_38_502 ();
 sg13g2_fill_2 FILLER_38_529 ();
 sg13g2_fill_2 FILLER_38_583 ();
 sg13g2_fill_2 FILLER_38_622 ();
 sg13g2_decap_8 FILLER_38_658 ();
 sg13g2_fill_2 FILLER_38_702 ();
 sg13g2_decap_4 FILLER_38_709 ();
 sg13g2_decap_8 FILLER_38_735 ();
 sg13g2_fill_1 FILLER_38_742 ();
 sg13g2_fill_1 FILLER_38_751 ();
 sg13g2_fill_1 FILLER_38_766 ();
 sg13g2_fill_2 FILLER_38_823 ();
 sg13g2_decap_4 FILLER_38_829 ();
 sg13g2_fill_2 FILLER_38_833 ();
 sg13g2_fill_2 FILLER_38_848 ();
 sg13g2_fill_2 FILLER_38_863 ();
 sg13g2_fill_1 FILLER_38_865 ();
 sg13g2_decap_4 FILLER_38_897 ();
 sg13g2_fill_2 FILLER_38_901 ();
 sg13g2_fill_2 FILLER_38_906 ();
 sg13g2_fill_1 FILLER_38_908 ();
 sg13g2_fill_1 FILLER_38_1011 ();
 sg13g2_fill_2 FILLER_38_1149 ();
 sg13g2_fill_2 FILLER_38_1220 ();
 sg13g2_fill_1 FILLER_38_1235 ();
 sg13g2_fill_1 FILLER_38_1282 ();
 sg13g2_fill_1 FILLER_38_1308 ();
 sg13g2_fill_2 FILLER_38_1313 ();
 sg13g2_fill_2 FILLER_38_1332 ();
 sg13g2_fill_1 FILLER_38_1352 ();
 sg13g2_fill_1 FILLER_38_1396 ();
 sg13g2_fill_1 FILLER_38_1463 ();
 sg13g2_decap_4 FILLER_38_1494 ();
 sg13g2_fill_2 FILLER_38_1498 ();
 sg13g2_fill_1 FILLER_38_1560 ();
 sg13g2_fill_1 FILLER_38_1592 ();
 sg13g2_decap_4 FILLER_38_1635 ();
 sg13g2_fill_2 FILLER_38_1654 ();
 sg13g2_fill_1 FILLER_38_1656 ();
 sg13g2_fill_1 FILLER_38_1665 ();
 sg13g2_fill_1 FILLER_38_1718 ();
 sg13g2_decap_4 FILLER_38_1745 ();
 sg13g2_fill_2 FILLER_38_1749 ();
 sg13g2_fill_2 FILLER_38_1755 ();
 sg13g2_fill_1 FILLER_38_1757 ();
 sg13g2_fill_2 FILLER_38_1766 ();
 sg13g2_fill_2 FILLER_38_1782 ();
 sg13g2_fill_1 FILLER_38_1784 ();
 sg13g2_fill_2 FILLER_38_1793 ();
 sg13g2_fill_1 FILLER_38_1795 ();
 sg13g2_fill_2 FILLER_38_1822 ();
 sg13g2_fill_1 FILLER_38_1824 ();
 sg13g2_fill_2 FILLER_38_1843 ();
 sg13g2_fill_1 FILLER_38_1845 ();
 sg13g2_fill_2 FILLER_38_1862 ();
 sg13g2_fill_1 FILLER_38_1882 ();
 sg13g2_decap_4 FILLER_38_1895 ();
 sg13g2_decap_8 FILLER_38_1915 ();
 sg13g2_decap_4 FILLER_38_1922 ();
 sg13g2_fill_2 FILLER_38_1926 ();
 sg13g2_decap_4 FILLER_38_1948 ();
 sg13g2_fill_1 FILLER_38_1968 ();
 sg13g2_decap_8 FILLER_38_1977 ();
 sg13g2_fill_1 FILLER_38_1984 ();
 sg13g2_decap_4 FILLER_38_2025 ();
 sg13g2_fill_2 FILLER_38_2043 ();
 sg13g2_fill_2 FILLER_38_2055 ();
 sg13g2_fill_2 FILLER_38_2114 ();
 sg13g2_decap_8 FILLER_38_2156 ();
 sg13g2_decap_4 FILLER_38_2163 ();
 sg13g2_decap_4 FILLER_38_2171 ();
 sg13g2_fill_1 FILLER_38_2175 ();
 sg13g2_fill_2 FILLER_38_2234 ();
 sg13g2_decap_8 FILLER_38_2249 ();
 sg13g2_decap_4 FILLER_38_2256 ();
 sg13g2_fill_1 FILLER_38_2260 ();
 sg13g2_decap_8 FILLER_38_2276 ();
 sg13g2_decap_4 FILLER_38_2303 ();
 sg13g2_decap_8 FILLER_38_2333 ();
 sg13g2_decap_8 FILLER_38_2340 ();
 sg13g2_decap_8 FILLER_38_2347 ();
 sg13g2_decap_8 FILLER_38_2354 ();
 sg13g2_decap_8 FILLER_38_2361 ();
 sg13g2_decap_8 FILLER_38_2368 ();
 sg13g2_decap_8 FILLER_38_2375 ();
 sg13g2_decap_8 FILLER_38_2382 ();
 sg13g2_decap_8 FILLER_38_2389 ();
 sg13g2_decap_8 FILLER_38_2396 ();
 sg13g2_decap_8 FILLER_38_2403 ();
 sg13g2_decap_8 FILLER_38_2410 ();
 sg13g2_decap_8 FILLER_38_2417 ();
 sg13g2_decap_8 FILLER_38_2424 ();
 sg13g2_decap_8 FILLER_38_2431 ();
 sg13g2_decap_8 FILLER_38_2438 ();
 sg13g2_decap_8 FILLER_38_2445 ();
 sg13g2_decap_8 FILLER_38_2452 ();
 sg13g2_decap_8 FILLER_38_2459 ();
 sg13g2_decap_8 FILLER_38_2466 ();
 sg13g2_decap_8 FILLER_38_2473 ();
 sg13g2_decap_8 FILLER_38_2480 ();
 sg13g2_decap_8 FILLER_38_2487 ();
 sg13g2_decap_8 FILLER_38_2494 ();
 sg13g2_decap_8 FILLER_38_2501 ();
 sg13g2_decap_8 FILLER_38_2508 ();
 sg13g2_decap_8 FILLER_38_2515 ();
 sg13g2_decap_8 FILLER_38_2522 ();
 sg13g2_decap_8 FILLER_38_2529 ();
 sg13g2_decap_8 FILLER_38_2536 ();
 sg13g2_decap_8 FILLER_38_2543 ();
 sg13g2_decap_8 FILLER_38_2550 ();
 sg13g2_decap_8 FILLER_38_2557 ();
 sg13g2_decap_8 FILLER_38_2564 ();
 sg13g2_decap_8 FILLER_38_2571 ();
 sg13g2_decap_8 FILLER_38_2578 ();
 sg13g2_decap_8 FILLER_38_2585 ();
 sg13g2_decap_8 FILLER_38_2592 ();
 sg13g2_decap_8 FILLER_38_2599 ();
 sg13g2_decap_8 FILLER_38_2606 ();
 sg13g2_decap_8 FILLER_38_2613 ();
 sg13g2_decap_8 FILLER_38_2620 ();
 sg13g2_decap_8 FILLER_38_2627 ();
 sg13g2_decap_8 FILLER_38_2634 ();
 sg13g2_decap_8 FILLER_38_2641 ();
 sg13g2_decap_8 FILLER_38_2648 ();
 sg13g2_decap_8 FILLER_38_2655 ();
 sg13g2_decap_8 FILLER_38_2662 ();
 sg13g2_decap_4 FILLER_38_2669 ();
 sg13g2_fill_1 FILLER_38_2673 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_4 FILLER_39_112 ();
 sg13g2_fill_1 FILLER_39_116 ();
 sg13g2_decap_8 FILLER_39_121 ();
 sg13g2_fill_1 FILLER_39_128 ();
 sg13g2_decap_4 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_145 ();
 sg13g2_decap_8 FILLER_39_152 ();
 sg13g2_fill_2 FILLER_39_159 ();
 sg13g2_fill_2 FILLER_39_183 ();
 sg13g2_fill_2 FILLER_39_210 ();
 sg13g2_decap_4 FILLER_39_220 ();
 sg13g2_decap_8 FILLER_39_265 ();
 sg13g2_decap_4 FILLER_39_285 ();
 sg13g2_fill_1 FILLER_39_289 ();
 sg13g2_fill_1 FILLER_39_325 ();
 sg13g2_fill_2 FILLER_39_355 ();
 sg13g2_fill_1 FILLER_39_357 ();
 sg13g2_fill_1 FILLER_39_363 ();
 sg13g2_fill_2 FILLER_39_381 ();
 sg13g2_fill_2 FILLER_39_389 ();
 sg13g2_fill_1 FILLER_39_391 ();
 sg13g2_decap_4 FILLER_39_435 ();
 sg13g2_decap_4 FILLER_39_449 ();
 sg13g2_fill_1 FILLER_39_453 ();
 sg13g2_fill_1 FILLER_39_485 ();
 sg13g2_fill_1 FILLER_39_502 ();
 sg13g2_fill_1 FILLER_39_544 ();
 sg13g2_fill_2 FILLER_39_568 ();
 sg13g2_fill_2 FILLER_39_587 ();
 sg13g2_fill_2 FILLER_39_601 ();
 sg13g2_fill_1 FILLER_39_611 ();
 sg13g2_fill_2 FILLER_39_625 ();
 sg13g2_fill_2 FILLER_39_639 ();
 sg13g2_fill_1 FILLER_39_641 ();
 sg13g2_fill_1 FILLER_39_677 ();
 sg13g2_fill_1 FILLER_39_695 ();
 sg13g2_fill_2 FILLER_39_704 ();
 sg13g2_decap_4 FILLER_39_724 ();
 sg13g2_fill_1 FILLER_39_766 ();
 sg13g2_fill_1 FILLER_39_786 ();
 sg13g2_fill_2 FILLER_39_801 ();
 sg13g2_decap_4 FILLER_39_816 ();
 sg13g2_fill_2 FILLER_39_820 ();
 sg13g2_decap_8 FILLER_39_853 ();
 sg13g2_decap_8 FILLER_39_860 ();
 sg13g2_fill_2 FILLER_39_867 ();
 sg13g2_fill_1 FILLER_39_869 ();
 sg13g2_decap_8 FILLER_39_874 ();
 sg13g2_decap_8 FILLER_39_913 ();
 sg13g2_decap_8 FILLER_39_920 ();
 sg13g2_decap_4 FILLER_39_927 ();
 sg13g2_fill_2 FILLER_39_989 ();
 sg13g2_fill_2 FILLER_39_1040 ();
 sg13g2_fill_1 FILLER_39_1047 ();
 sg13g2_fill_1 FILLER_39_1074 ();
 sg13g2_fill_1 FILLER_39_1118 ();
 sg13g2_fill_2 FILLER_39_1206 ();
 sg13g2_fill_1 FILLER_39_1270 ();
 sg13g2_fill_2 FILLER_39_1289 ();
 sg13g2_fill_2 FILLER_39_1300 ();
 sg13g2_fill_1 FILLER_39_1343 ();
 sg13g2_fill_1 FILLER_39_1449 ();
 sg13g2_fill_2 FILLER_39_1508 ();
 sg13g2_fill_1 FILLER_39_1549 ();
 sg13g2_decap_4 FILLER_39_1559 ();
 sg13g2_fill_2 FILLER_39_1563 ();
 sg13g2_fill_2 FILLER_39_1644 ();
 sg13g2_fill_1 FILLER_39_1665 ();
 sg13g2_decap_4 FILLER_39_1705 ();
 sg13g2_fill_1 FILLER_39_1713 ();
 sg13g2_fill_1 FILLER_39_1722 ();
 sg13g2_fill_2 FILLER_39_1728 ();
 sg13g2_decap_4 FILLER_39_1734 ();
 sg13g2_fill_2 FILLER_39_1738 ();
 sg13g2_fill_1 FILLER_39_1766 ();
 sg13g2_decap_8 FILLER_39_1779 ();
 sg13g2_fill_2 FILLER_39_1786 ();
 sg13g2_decap_8 FILLER_39_1793 ();
 sg13g2_decap_8 FILLER_39_1800 ();
 sg13g2_fill_2 FILLER_39_1811 ();
 sg13g2_fill_1 FILLER_39_1813 ();
 sg13g2_decap_8 FILLER_39_1840 ();
 sg13g2_fill_1 FILLER_39_1863 ();
 sg13g2_fill_2 FILLER_39_1880 ();
 sg13g2_fill_1 FILLER_39_1904 ();
 sg13g2_fill_2 FILLER_39_1937 ();
 sg13g2_fill_1 FILLER_39_1939 ();
 sg13g2_decap_8 FILLER_39_1945 ();
 sg13g2_decap_4 FILLER_39_1952 ();
 sg13g2_fill_1 FILLER_39_1956 ();
 sg13g2_decap_8 FILLER_39_1965 ();
 sg13g2_decap_8 FILLER_39_1972 ();
 sg13g2_decap_8 FILLER_39_1979 ();
 sg13g2_fill_2 FILLER_39_1986 ();
 sg13g2_fill_1 FILLER_39_1988 ();
 sg13g2_fill_2 FILLER_39_2002 ();
 sg13g2_fill_2 FILLER_39_2016 ();
 sg13g2_fill_1 FILLER_39_2018 ();
 sg13g2_fill_2 FILLER_39_2058 ();
 sg13g2_decap_4 FILLER_39_2073 ();
 sg13g2_fill_2 FILLER_39_2077 ();
 sg13g2_fill_2 FILLER_39_2087 ();
 sg13g2_decap_4 FILLER_39_2093 ();
 sg13g2_fill_1 FILLER_39_2097 ();
 sg13g2_decap_4 FILLER_39_2106 ();
 sg13g2_fill_2 FILLER_39_2110 ();
 sg13g2_decap_4 FILLER_39_2169 ();
 sg13g2_fill_2 FILLER_39_2173 ();
 sg13g2_fill_2 FILLER_39_2209 ();
 sg13g2_fill_1 FILLER_39_2229 ();
 sg13g2_fill_2 FILLER_39_2251 ();
 sg13g2_fill_2 FILLER_39_2304 ();
 sg13g2_decap_8 FILLER_39_2332 ();
 sg13g2_decap_8 FILLER_39_2339 ();
 sg13g2_decap_8 FILLER_39_2346 ();
 sg13g2_decap_8 FILLER_39_2353 ();
 sg13g2_decap_8 FILLER_39_2360 ();
 sg13g2_decap_8 FILLER_39_2367 ();
 sg13g2_decap_8 FILLER_39_2374 ();
 sg13g2_decap_8 FILLER_39_2381 ();
 sg13g2_decap_8 FILLER_39_2388 ();
 sg13g2_decap_8 FILLER_39_2395 ();
 sg13g2_decap_8 FILLER_39_2402 ();
 sg13g2_decap_8 FILLER_39_2409 ();
 sg13g2_decap_8 FILLER_39_2416 ();
 sg13g2_decap_8 FILLER_39_2423 ();
 sg13g2_decap_8 FILLER_39_2430 ();
 sg13g2_decap_8 FILLER_39_2437 ();
 sg13g2_decap_8 FILLER_39_2444 ();
 sg13g2_decap_8 FILLER_39_2451 ();
 sg13g2_decap_8 FILLER_39_2458 ();
 sg13g2_decap_8 FILLER_39_2465 ();
 sg13g2_decap_8 FILLER_39_2472 ();
 sg13g2_decap_8 FILLER_39_2479 ();
 sg13g2_decap_8 FILLER_39_2486 ();
 sg13g2_decap_8 FILLER_39_2493 ();
 sg13g2_decap_8 FILLER_39_2500 ();
 sg13g2_decap_8 FILLER_39_2507 ();
 sg13g2_decap_8 FILLER_39_2514 ();
 sg13g2_decap_8 FILLER_39_2521 ();
 sg13g2_decap_8 FILLER_39_2528 ();
 sg13g2_decap_8 FILLER_39_2535 ();
 sg13g2_decap_8 FILLER_39_2542 ();
 sg13g2_decap_8 FILLER_39_2549 ();
 sg13g2_decap_8 FILLER_39_2556 ();
 sg13g2_decap_8 FILLER_39_2563 ();
 sg13g2_decap_8 FILLER_39_2570 ();
 sg13g2_decap_8 FILLER_39_2577 ();
 sg13g2_decap_8 FILLER_39_2584 ();
 sg13g2_decap_8 FILLER_39_2591 ();
 sg13g2_decap_8 FILLER_39_2598 ();
 sg13g2_decap_8 FILLER_39_2605 ();
 sg13g2_decap_8 FILLER_39_2612 ();
 sg13g2_decap_8 FILLER_39_2619 ();
 sg13g2_decap_8 FILLER_39_2626 ();
 sg13g2_decap_8 FILLER_39_2633 ();
 sg13g2_decap_8 FILLER_39_2640 ();
 sg13g2_decap_8 FILLER_39_2647 ();
 sg13g2_decap_8 FILLER_39_2654 ();
 sg13g2_decap_8 FILLER_39_2661 ();
 sg13g2_decap_4 FILLER_39_2668 ();
 sg13g2_fill_2 FILLER_39_2672 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_fill_1 FILLER_40_133 ();
 sg13g2_fill_2 FILLER_40_160 ();
 sg13g2_decap_4 FILLER_40_171 ();
 sg13g2_fill_2 FILLER_40_202 ();
 sg13g2_fill_1 FILLER_40_204 ();
 sg13g2_decap_8 FILLER_40_209 ();
 sg13g2_fill_2 FILLER_40_228 ();
 sg13g2_fill_1 FILLER_40_248 ();
 sg13g2_decap_8 FILLER_40_275 ();
 sg13g2_fill_1 FILLER_40_282 ();
 sg13g2_fill_2 FILLER_40_288 ();
 sg13g2_fill_1 FILLER_40_290 ();
 sg13g2_fill_2 FILLER_40_370 ();
 sg13g2_fill_1 FILLER_40_372 ();
 sg13g2_fill_2 FILLER_40_378 ();
 sg13g2_fill_1 FILLER_40_390 ();
 sg13g2_fill_2 FILLER_40_400 ();
 sg13g2_decap_8 FILLER_40_406 ();
 sg13g2_decap_8 FILLER_40_420 ();
 sg13g2_fill_1 FILLER_40_427 ();
 sg13g2_decap_4 FILLER_40_458 ();
 sg13g2_fill_1 FILLER_40_462 ();
 sg13g2_fill_2 FILLER_40_484 ();
 sg13g2_fill_1 FILLER_40_486 ();
 sg13g2_decap_8 FILLER_40_504 ();
 sg13g2_fill_2 FILLER_40_511 ();
 sg13g2_fill_1 FILLER_40_513 ();
 sg13g2_fill_1 FILLER_40_522 ();
 sg13g2_fill_1 FILLER_40_533 ();
 sg13g2_fill_1 FILLER_40_574 ();
 sg13g2_fill_1 FILLER_40_614 ();
 sg13g2_decap_8 FILLER_40_623 ();
 sg13g2_fill_2 FILLER_40_630 ();
 sg13g2_fill_1 FILLER_40_632 ();
 sg13g2_decap_8 FILLER_40_641 ();
 sg13g2_decap_8 FILLER_40_648 ();
 sg13g2_fill_1 FILLER_40_655 ();
 sg13g2_fill_2 FILLER_40_666 ();
 sg13g2_fill_2 FILLER_40_689 ();
 sg13g2_fill_1 FILLER_40_691 ();
 sg13g2_fill_2 FILLER_40_722 ();
 sg13g2_fill_2 FILLER_40_738 ();
 sg13g2_fill_2 FILLER_40_780 ();
 sg13g2_fill_1 FILLER_40_782 ();
 sg13g2_fill_2 FILLER_40_791 ();
 sg13g2_fill_1 FILLER_40_823 ();
 sg13g2_fill_1 FILLER_40_844 ();
 sg13g2_decap_4 FILLER_40_867 ();
 sg13g2_fill_2 FILLER_40_871 ();
 sg13g2_decap_8 FILLER_40_885 ();
 sg13g2_fill_2 FILLER_40_892 ();
 sg13g2_decap_4 FILLER_40_898 ();
 sg13g2_fill_2 FILLER_40_902 ();
 sg13g2_decap_8 FILLER_40_915 ();
 sg13g2_fill_1 FILLER_40_922 ();
 sg13g2_decap_8 FILLER_40_932 ();
 sg13g2_fill_1 FILLER_40_939 ();
 sg13g2_fill_1 FILLER_40_945 ();
 sg13g2_fill_1 FILLER_40_963 ();
 sg13g2_fill_1 FILLER_40_1020 ();
 sg13g2_fill_1 FILLER_40_1039 ();
 sg13g2_fill_2 FILLER_40_1095 ();
 sg13g2_fill_1 FILLER_40_1124 ();
 sg13g2_fill_1 FILLER_40_1155 ();
 sg13g2_fill_1 FILLER_40_1224 ();
 sg13g2_fill_2 FILLER_40_1243 ();
 sg13g2_fill_2 FILLER_40_1271 ();
 sg13g2_fill_2 FILLER_40_1282 ();
 sg13g2_fill_2 FILLER_40_1310 ();
 sg13g2_fill_1 FILLER_40_1363 ();
 sg13g2_fill_1 FILLER_40_1390 ();
 sg13g2_fill_2 FILLER_40_1436 ();
 sg13g2_fill_1 FILLER_40_1463 ();
 sg13g2_fill_2 FILLER_40_1562 ();
 sg13g2_fill_1 FILLER_40_1564 ();
 sg13g2_fill_2 FILLER_40_1570 ();
 sg13g2_decap_4 FILLER_40_1585 ();
 sg13g2_fill_2 FILLER_40_1604 ();
 sg13g2_fill_1 FILLER_40_1623 ();
 sg13g2_fill_1 FILLER_40_1629 ();
 sg13g2_fill_1 FILLER_40_1636 ();
 sg13g2_fill_2 FILLER_40_1645 ();
 sg13g2_decap_4 FILLER_40_1699 ();
 sg13g2_decap_8 FILLER_40_1729 ();
 sg13g2_decap_8 FILLER_40_1736 ();
 sg13g2_decap_8 FILLER_40_1743 ();
 sg13g2_fill_2 FILLER_40_1763 ();
 sg13g2_fill_1 FILLER_40_1765 ();
 sg13g2_fill_1 FILLER_40_1775 ();
 sg13g2_decap_8 FILLER_40_1802 ();
 sg13g2_decap_4 FILLER_40_1809 ();
 sg13g2_fill_1 FILLER_40_1813 ();
 sg13g2_decap_8 FILLER_40_1839 ();
 sg13g2_fill_2 FILLER_40_1846 ();
 sg13g2_fill_1 FILLER_40_1848 ();
 sg13g2_decap_8 FILLER_40_1866 ();
 sg13g2_decap_8 FILLER_40_1873 ();
 sg13g2_decap_4 FILLER_40_1880 ();
 sg13g2_fill_1 FILLER_40_1898 ();
 sg13g2_fill_2 FILLER_40_1907 ();
 sg13g2_fill_1 FILLER_40_1909 ();
 sg13g2_fill_1 FILLER_40_1928 ();
 sg13g2_decap_4 FILLER_40_1958 ();
 sg13g2_fill_2 FILLER_40_1962 ();
 sg13g2_decap_8 FILLER_40_2002 ();
 sg13g2_decap_8 FILLER_40_2022 ();
 sg13g2_fill_1 FILLER_40_2029 ();
 sg13g2_decap_8 FILLER_40_2034 ();
 sg13g2_decap_4 FILLER_40_2041 ();
 sg13g2_fill_1 FILLER_40_2045 ();
 sg13g2_fill_2 FILLER_40_2050 ();
 sg13g2_decap_4 FILLER_40_2057 ();
 sg13g2_fill_1 FILLER_40_2061 ();
 sg13g2_decap_4 FILLER_40_2088 ();
 sg13g2_fill_1 FILLER_40_2092 ();
 sg13g2_decap_8 FILLER_40_2111 ();
 sg13g2_decap_4 FILLER_40_2118 ();
 sg13g2_fill_1 FILLER_40_2122 ();
 sg13g2_decap_8 FILLER_40_2127 ();
 sg13g2_fill_2 FILLER_40_2134 ();
 sg13g2_fill_1 FILLER_40_2136 ();
 sg13g2_decap_4 FILLER_40_2145 ();
 sg13g2_fill_2 FILLER_40_2149 ();
 sg13g2_fill_1 FILLER_40_2198 ();
 sg13g2_decap_4 FILLER_40_2233 ();
 sg13g2_fill_2 FILLER_40_2251 ();
 sg13g2_fill_1 FILLER_40_2253 ();
 sg13g2_fill_2 FILLER_40_2285 ();
 sg13g2_fill_1 FILLER_40_2287 ();
 sg13g2_decap_4 FILLER_40_2292 ();
 sg13g2_fill_1 FILLER_40_2296 ();
 sg13g2_decap_4 FILLER_40_2310 ();
 sg13g2_decap_8 FILLER_40_2331 ();
 sg13g2_decap_8 FILLER_40_2338 ();
 sg13g2_decap_8 FILLER_40_2345 ();
 sg13g2_decap_8 FILLER_40_2352 ();
 sg13g2_decap_8 FILLER_40_2359 ();
 sg13g2_decap_8 FILLER_40_2366 ();
 sg13g2_decap_8 FILLER_40_2373 ();
 sg13g2_decap_8 FILLER_40_2380 ();
 sg13g2_decap_8 FILLER_40_2387 ();
 sg13g2_decap_8 FILLER_40_2394 ();
 sg13g2_decap_8 FILLER_40_2401 ();
 sg13g2_decap_8 FILLER_40_2408 ();
 sg13g2_decap_8 FILLER_40_2415 ();
 sg13g2_decap_8 FILLER_40_2422 ();
 sg13g2_decap_8 FILLER_40_2429 ();
 sg13g2_decap_8 FILLER_40_2436 ();
 sg13g2_decap_8 FILLER_40_2443 ();
 sg13g2_decap_8 FILLER_40_2450 ();
 sg13g2_decap_8 FILLER_40_2457 ();
 sg13g2_decap_8 FILLER_40_2464 ();
 sg13g2_decap_8 FILLER_40_2471 ();
 sg13g2_decap_8 FILLER_40_2478 ();
 sg13g2_decap_8 FILLER_40_2485 ();
 sg13g2_decap_8 FILLER_40_2492 ();
 sg13g2_decap_8 FILLER_40_2499 ();
 sg13g2_decap_8 FILLER_40_2506 ();
 sg13g2_decap_8 FILLER_40_2513 ();
 sg13g2_decap_8 FILLER_40_2520 ();
 sg13g2_decap_8 FILLER_40_2527 ();
 sg13g2_decap_8 FILLER_40_2534 ();
 sg13g2_decap_8 FILLER_40_2541 ();
 sg13g2_decap_8 FILLER_40_2548 ();
 sg13g2_decap_8 FILLER_40_2555 ();
 sg13g2_decap_8 FILLER_40_2562 ();
 sg13g2_decap_8 FILLER_40_2569 ();
 sg13g2_decap_8 FILLER_40_2576 ();
 sg13g2_decap_8 FILLER_40_2583 ();
 sg13g2_decap_8 FILLER_40_2590 ();
 sg13g2_decap_8 FILLER_40_2597 ();
 sg13g2_decap_8 FILLER_40_2604 ();
 sg13g2_decap_8 FILLER_40_2611 ();
 sg13g2_decap_8 FILLER_40_2618 ();
 sg13g2_decap_8 FILLER_40_2625 ();
 sg13g2_decap_8 FILLER_40_2632 ();
 sg13g2_decap_8 FILLER_40_2639 ();
 sg13g2_decap_8 FILLER_40_2646 ();
 sg13g2_decap_8 FILLER_40_2653 ();
 sg13g2_decap_8 FILLER_40_2660 ();
 sg13g2_decap_8 FILLER_40_2667 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_4 FILLER_41_133 ();
 sg13g2_fill_2 FILLER_41_137 ();
 sg13g2_fill_1 FILLER_41_169 ();
 sg13g2_fill_1 FILLER_41_176 ();
 sg13g2_fill_2 FILLER_41_192 ();
 sg13g2_fill_2 FILLER_41_237 ();
 sg13g2_fill_1 FILLER_41_239 ();
 sg13g2_fill_2 FILLER_41_250 ();
 sg13g2_decap_4 FILLER_41_260 ();
 sg13g2_fill_1 FILLER_41_264 ();
 sg13g2_decap_4 FILLER_41_295 ();
 sg13g2_decap_8 FILLER_41_311 ();
 sg13g2_decap_4 FILLER_41_318 ();
 sg13g2_decap_4 FILLER_41_328 ();
 sg13g2_fill_2 FILLER_41_354 ();
 sg13g2_fill_1 FILLER_41_376 ();
 sg13g2_fill_1 FILLER_41_395 ();
 sg13g2_fill_2 FILLER_41_415 ();
 sg13g2_fill_1 FILLER_41_417 ();
 sg13g2_fill_1 FILLER_41_429 ();
 sg13g2_fill_2 FILLER_41_451 ();
 sg13g2_decap_8 FILLER_41_461 ();
 sg13g2_fill_1 FILLER_41_468 ();
 sg13g2_decap_4 FILLER_41_520 ();
 sg13g2_decap_8 FILLER_41_529 ();
 sg13g2_fill_2 FILLER_41_536 ();
 sg13g2_fill_2 FILLER_41_591 ();
 sg13g2_fill_2 FILLER_41_607 ();
 sg13g2_fill_2 FILLER_41_627 ();
 sg13g2_fill_1 FILLER_41_629 ();
 sg13g2_fill_2 FILLER_41_669 ();
 sg13g2_fill_1 FILLER_41_671 ();
 sg13g2_fill_1 FILLER_41_712 ();
 sg13g2_fill_2 FILLER_41_719 ();
 sg13g2_decap_4 FILLER_41_727 ();
 sg13g2_fill_1 FILLER_41_731 ();
 sg13g2_fill_2 FILLER_41_740 ();
 sg13g2_fill_1 FILLER_41_768 ();
 sg13g2_fill_2 FILLER_41_782 ();
 sg13g2_fill_2 FILLER_41_798 ();
 sg13g2_fill_1 FILLER_41_800 ();
 sg13g2_fill_1 FILLER_41_814 ();
 sg13g2_fill_2 FILLER_41_828 ();
 sg13g2_decap_4 FILLER_41_834 ();
 sg13g2_fill_2 FILLER_41_838 ();
 sg13g2_decap_8 FILLER_41_844 ();
 sg13g2_decap_8 FILLER_41_855 ();
 sg13g2_decap_4 FILLER_41_862 ();
 sg13g2_fill_2 FILLER_41_866 ();
 sg13g2_decap_4 FILLER_41_872 ();
 sg13g2_decap_8 FILLER_41_889 ();
 sg13g2_decap_8 FILLER_41_896 ();
 sg13g2_decap_4 FILLER_41_903 ();
 sg13g2_decap_8 FILLER_41_910 ();
 sg13g2_decap_4 FILLER_41_917 ();
 sg13g2_fill_2 FILLER_41_921 ();
 sg13g2_decap_8 FILLER_41_928 ();
 sg13g2_decap_4 FILLER_41_935 ();
 sg13g2_fill_1 FILLER_41_939 ();
 sg13g2_fill_1 FILLER_41_1017 ();
 sg13g2_fill_2 FILLER_41_1053 ();
 sg13g2_fill_1 FILLER_41_1090 ();
 sg13g2_fill_2 FILLER_41_1171 ();
 sg13g2_fill_2 FILLER_41_1346 ();
 sg13g2_fill_2 FILLER_41_1542 ();
 sg13g2_decap_8 FILLER_41_1579 ();
 sg13g2_fill_2 FILLER_41_1617 ();
 sg13g2_fill_1 FILLER_41_1619 ();
 sg13g2_fill_2 FILLER_41_1623 ();
 sg13g2_fill_1 FILLER_41_1649 ();
 sg13g2_fill_2 FILLER_41_1668 ();
 sg13g2_fill_1 FILLER_41_1670 ();
 sg13g2_decap_4 FILLER_41_1762 ();
 sg13g2_fill_2 FILLER_41_1786 ();
 sg13g2_fill_1 FILLER_41_1788 ();
 sg13g2_fill_1 FILLER_41_1810 ();
 sg13g2_decap_8 FILLER_41_1815 ();
 sg13g2_decap_4 FILLER_41_1822 ();
 sg13g2_fill_2 FILLER_41_1841 ();
 sg13g2_fill_2 FILLER_41_1864 ();
 sg13g2_fill_1 FILLER_41_1866 ();
 sg13g2_decap_8 FILLER_41_1922 ();
 sg13g2_fill_1 FILLER_41_1929 ();
 sg13g2_fill_2 FILLER_41_1937 ();
 sg13g2_fill_1 FILLER_41_1939 ();
 sg13g2_decap_8 FILLER_41_1945 ();
 sg13g2_fill_2 FILLER_41_2023 ();
 sg13g2_decap_4 FILLER_41_2067 ();
 sg13g2_fill_2 FILLER_41_2071 ();
 sg13g2_fill_2 FILLER_41_2077 ();
 sg13g2_fill_1 FILLER_41_2079 ();
 sg13g2_decap_8 FILLER_41_2152 ();
 sg13g2_decap_8 FILLER_41_2159 ();
 sg13g2_fill_2 FILLER_41_2166 ();
 sg13g2_decap_8 FILLER_41_2177 ();
 sg13g2_fill_1 FILLER_41_2184 ();
 sg13g2_fill_1 FILLER_41_2190 ();
 sg13g2_decap_8 FILLER_41_2200 ();
 sg13g2_decap_8 FILLER_41_2207 ();
 sg13g2_decap_8 FILLER_41_2214 ();
 sg13g2_decap_8 FILLER_41_2221 ();
 sg13g2_fill_1 FILLER_41_2228 ();
 sg13g2_fill_2 FILLER_41_2245 ();
 sg13g2_decap_8 FILLER_41_2252 ();
 sg13g2_fill_2 FILLER_41_2259 ();
 sg13g2_fill_1 FILLER_41_2315 ();
 sg13g2_decap_8 FILLER_41_2342 ();
 sg13g2_decap_8 FILLER_41_2349 ();
 sg13g2_decap_8 FILLER_41_2356 ();
 sg13g2_decap_8 FILLER_41_2363 ();
 sg13g2_decap_8 FILLER_41_2370 ();
 sg13g2_decap_8 FILLER_41_2377 ();
 sg13g2_decap_8 FILLER_41_2384 ();
 sg13g2_decap_8 FILLER_41_2391 ();
 sg13g2_decap_8 FILLER_41_2398 ();
 sg13g2_decap_8 FILLER_41_2405 ();
 sg13g2_decap_8 FILLER_41_2412 ();
 sg13g2_decap_8 FILLER_41_2419 ();
 sg13g2_decap_8 FILLER_41_2426 ();
 sg13g2_decap_8 FILLER_41_2433 ();
 sg13g2_decap_8 FILLER_41_2440 ();
 sg13g2_decap_8 FILLER_41_2447 ();
 sg13g2_decap_8 FILLER_41_2454 ();
 sg13g2_decap_8 FILLER_41_2461 ();
 sg13g2_decap_8 FILLER_41_2468 ();
 sg13g2_decap_8 FILLER_41_2475 ();
 sg13g2_decap_8 FILLER_41_2482 ();
 sg13g2_decap_8 FILLER_41_2489 ();
 sg13g2_decap_8 FILLER_41_2496 ();
 sg13g2_decap_8 FILLER_41_2503 ();
 sg13g2_decap_8 FILLER_41_2510 ();
 sg13g2_decap_8 FILLER_41_2517 ();
 sg13g2_decap_8 FILLER_41_2524 ();
 sg13g2_decap_8 FILLER_41_2531 ();
 sg13g2_decap_8 FILLER_41_2538 ();
 sg13g2_decap_8 FILLER_41_2545 ();
 sg13g2_decap_8 FILLER_41_2552 ();
 sg13g2_decap_8 FILLER_41_2559 ();
 sg13g2_decap_8 FILLER_41_2566 ();
 sg13g2_decap_8 FILLER_41_2573 ();
 sg13g2_decap_8 FILLER_41_2580 ();
 sg13g2_decap_8 FILLER_41_2587 ();
 sg13g2_decap_8 FILLER_41_2594 ();
 sg13g2_decap_8 FILLER_41_2601 ();
 sg13g2_decap_8 FILLER_41_2608 ();
 sg13g2_decap_8 FILLER_41_2615 ();
 sg13g2_decap_8 FILLER_41_2622 ();
 sg13g2_decap_8 FILLER_41_2629 ();
 sg13g2_decap_8 FILLER_41_2636 ();
 sg13g2_decap_8 FILLER_41_2643 ();
 sg13g2_decap_8 FILLER_41_2650 ();
 sg13g2_decap_8 FILLER_41_2657 ();
 sg13g2_decap_8 FILLER_41_2664 ();
 sg13g2_fill_2 FILLER_41_2671 ();
 sg13g2_fill_1 FILLER_41_2673 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_4 FILLER_42_158 ();
 sg13g2_decap_4 FILLER_42_180 ();
 sg13g2_fill_2 FILLER_42_184 ();
 sg13g2_fill_2 FILLER_42_204 ();
 sg13g2_fill_1 FILLER_42_206 ();
 sg13g2_decap_4 FILLER_42_223 ();
 sg13g2_fill_1 FILLER_42_227 ();
 sg13g2_fill_1 FILLER_42_232 ();
 sg13g2_fill_2 FILLER_42_253 ();
 sg13g2_decap_8 FILLER_42_260 ();
 sg13g2_fill_1 FILLER_42_267 ();
 sg13g2_fill_2 FILLER_42_276 ();
 sg13g2_fill_2 FILLER_42_309 ();
 sg13g2_fill_1 FILLER_42_332 ();
 sg13g2_fill_2 FILLER_42_383 ();
 sg13g2_decap_8 FILLER_42_396 ();
 sg13g2_decap_8 FILLER_42_403 ();
 sg13g2_fill_2 FILLER_42_410 ();
 sg13g2_decap_8 FILLER_42_429 ();
 sg13g2_fill_1 FILLER_42_436 ();
 sg13g2_decap_8 FILLER_42_465 ();
 sg13g2_fill_2 FILLER_42_472 ();
 sg13g2_fill_1 FILLER_42_474 ();
 sg13g2_fill_2 FILLER_42_479 ();
 sg13g2_fill_1 FILLER_42_502 ();
 sg13g2_fill_2 FILLER_42_514 ();
 sg13g2_fill_1 FILLER_42_516 ();
 sg13g2_decap_8 FILLER_42_537 ();
 sg13g2_fill_1 FILLER_42_557 ();
 sg13g2_decap_4 FILLER_42_598 ();
 sg13g2_fill_1 FILLER_42_602 ();
 sg13g2_fill_2 FILLER_42_608 ();
 sg13g2_fill_2 FILLER_42_618 ();
 sg13g2_decap_8 FILLER_42_625 ();
 sg13g2_fill_1 FILLER_42_632 ();
 sg13g2_decap_8 FILLER_42_638 ();
 sg13g2_fill_1 FILLER_42_645 ();
 sg13g2_fill_1 FILLER_42_666 ();
 sg13g2_fill_2 FILLER_42_675 ();
 sg13g2_fill_2 FILLER_42_686 ();
 sg13g2_fill_1 FILLER_42_688 ();
 sg13g2_fill_1 FILLER_42_708 ();
 sg13g2_decap_8 FILLER_42_717 ();
 sg13g2_fill_1 FILLER_42_724 ();
 sg13g2_decap_4 FILLER_42_733 ();
 sg13g2_fill_2 FILLER_42_831 ();
 sg13g2_fill_1 FILLER_42_833 ();
 sg13g2_decap_4 FILLER_42_851 ();
 sg13g2_fill_2 FILLER_42_855 ();
 sg13g2_decap_8 FILLER_42_883 ();
 sg13g2_decap_8 FILLER_42_890 ();
 sg13g2_decap_8 FILLER_42_897 ();
 sg13g2_decap_8 FILLER_42_904 ();
 sg13g2_decap_8 FILLER_42_911 ();
 sg13g2_fill_2 FILLER_42_918 ();
 sg13g2_fill_1 FILLER_42_946 ();
 sg13g2_fill_1 FILLER_42_973 ();
 sg13g2_fill_2 FILLER_42_1080 ();
 sg13g2_fill_1 FILLER_42_1122 ();
 sg13g2_fill_1 FILLER_42_1142 ();
 sg13g2_fill_1 FILLER_42_1161 ();
 sg13g2_fill_2 FILLER_42_1215 ();
 sg13g2_fill_1 FILLER_42_1276 ();
 sg13g2_fill_1 FILLER_42_1313 ();
 sg13g2_fill_2 FILLER_42_1328 ();
 sg13g2_fill_1 FILLER_42_1356 ();
 sg13g2_fill_1 FILLER_42_1362 ();
 sg13g2_fill_1 FILLER_42_1421 ();
 sg13g2_fill_2 FILLER_42_1492 ();
 sg13g2_fill_1 FILLER_42_1494 ();
 sg13g2_decap_8 FILLER_42_1500 ();
 sg13g2_fill_2 FILLER_42_1507 ();
 sg13g2_fill_1 FILLER_42_1563 ();
 sg13g2_decap_4 FILLER_42_1568 ();
 sg13g2_fill_1 FILLER_42_1572 ();
 sg13g2_fill_1 FILLER_42_1578 ();
 sg13g2_fill_1 FILLER_42_1587 ();
 sg13g2_decap_4 FILLER_42_1598 ();
 sg13g2_decap_8 FILLER_42_1606 ();
 sg13g2_fill_2 FILLER_42_1613 ();
 sg13g2_fill_1 FILLER_42_1615 ();
 sg13g2_fill_2 FILLER_42_1676 ();
 sg13g2_fill_1 FILLER_42_1716 ();
 sg13g2_decap_4 FILLER_42_1722 ();
 sg13g2_fill_2 FILLER_42_1726 ();
 sg13g2_fill_1 FILLER_42_1732 ();
 sg13g2_fill_2 FILLER_42_1769 ();
 sg13g2_decap_8 FILLER_42_1779 ();
 sg13g2_decap_4 FILLER_42_1790 ();
 sg13g2_fill_1 FILLER_42_1799 ();
 sg13g2_fill_1 FILLER_42_1830 ();
 sg13g2_decap_8 FILLER_42_1839 ();
 sg13g2_decap_8 FILLER_42_1867 ();
 sg13g2_decap_8 FILLER_42_1874 ();
 sg13g2_decap_8 FILLER_42_1881 ();
 sg13g2_fill_2 FILLER_42_1888 ();
 sg13g2_decap_8 FILLER_42_1895 ();
 sg13g2_fill_2 FILLER_42_1906 ();
 sg13g2_fill_1 FILLER_42_1908 ();
 sg13g2_decap_4 FILLER_42_1938 ();
 sg13g2_fill_2 FILLER_42_1942 ();
 sg13g2_decap_4 FILLER_42_1960 ();
 sg13g2_fill_1 FILLER_42_1964 ();
 sg13g2_decap_8 FILLER_42_1973 ();
 sg13g2_decap_4 FILLER_42_1980 ();
 sg13g2_decap_4 FILLER_42_2001 ();
 sg13g2_fill_2 FILLER_42_2005 ();
 sg13g2_fill_1 FILLER_42_2019 ();
 sg13g2_decap_8 FILLER_42_2028 ();
 sg13g2_fill_2 FILLER_42_2035 ();
 sg13g2_decap_4 FILLER_42_2049 ();
 sg13g2_fill_1 FILLER_42_2053 ();
 sg13g2_fill_1 FILLER_42_2062 ();
 sg13g2_decap_8 FILLER_42_2089 ();
 sg13g2_fill_2 FILLER_42_2114 ();
 sg13g2_decap_4 FILLER_42_2126 ();
 sg13g2_fill_1 FILLER_42_2130 ();
 sg13g2_fill_1 FILLER_42_2145 ();
 sg13g2_decap_8 FILLER_42_2228 ();
 sg13g2_fill_2 FILLER_42_2251 ();
 sg13g2_fill_1 FILLER_42_2253 ();
 sg13g2_fill_1 FILLER_42_2270 ();
 sg13g2_decap_8 FILLER_42_2294 ();
 sg13g2_decap_8 FILLER_42_2301 ();
 sg13g2_decap_4 FILLER_42_2308 ();
 sg13g2_decap_8 FILLER_42_2338 ();
 sg13g2_decap_8 FILLER_42_2345 ();
 sg13g2_decap_8 FILLER_42_2352 ();
 sg13g2_decap_8 FILLER_42_2359 ();
 sg13g2_decap_8 FILLER_42_2366 ();
 sg13g2_decap_8 FILLER_42_2373 ();
 sg13g2_decap_8 FILLER_42_2380 ();
 sg13g2_decap_8 FILLER_42_2387 ();
 sg13g2_decap_8 FILLER_42_2394 ();
 sg13g2_decap_8 FILLER_42_2401 ();
 sg13g2_decap_8 FILLER_42_2408 ();
 sg13g2_decap_8 FILLER_42_2415 ();
 sg13g2_decap_8 FILLER_42_2422 ();
 sg13g2_decap_8 FILLER_42_2429 ();
 sg13g2_decap_8 FILLER_42_2436 ();
 sg13g2_decap_8 FILLER_42_2443 ();
 sg13g2_decap_8 FILLER_42_2450 ();
 sg13g2_decap_8 FILLER_42_2457 ();
 sg13g2_decap_8 FILLER_42_2464 ();
 sg13g2_decap_8 FILLER_42_2471 ();
 sg13g2_decap_8 FILLER_42_2478 ();
 sg13g2_decap_8 FILLER_42_2485 ();
 sg13g2_decap_8 FILLER_42_2492 ();
 sg13g2_decap_8 FILLER_42_2499 ();
 sg13g2_decap_8 FILLER_42_2506 ();
 sg13g2_decap_8 FILLER_42_2513 ();
 sg13g2_decap_8 FILLER_42_2520 ();
 sg13g2_decap_8 FILLER_42_2527 ();
 sg13g2_decap_8 FILLER_42_2534 ();
 sg13g2_decap_8 FILLER_42_2541 ();
 sg13g2_decap_8 FILLER_42_2548 ();
 sg13g2_decap_8 FILLER_42_2555 ();
 sg13g2_decap_8 FILLER_42_2562 ();
 sg13g2_decap_8 FILLER_42_2569 ();
 sg13g2_decap_8 FILLER_42_2576 ();
 sg13g2_decap_8 FILLER_42_2583 ();
 sg13g2_decap_8 FILLER_42_2590 ();
 sg13g2_decap_8 FILLER_42_2597 ();
 sg13g2_decap_8 FILLER_42_2604 ();
 sg13g2_decap_8 FILLER_42_2611 ();
 sg13g2_decap_8 FILLER_42_2618 ();
 sg13g2_decap_8 FILLER_42_2625 ();
 sg13g2_decap_8 FILLER_42_2632 ();
 sg13g2_decap_8 FILLER_42_2639 ();
 sg13g2_decap_8 FILLER_42_2646 ();
 sg13g2_decap_8 FILLER_42_2653 ();
 sg13g2_decap_8 FILLER_42_2660 ();
 sg13g2_decap_8 FILLER_42_2667 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_4 FILLER_43_161 ();
 sg13g2_fill_2 FILLER_43_165 ();
 sg13g2_fill_1 FILLER_43_210 ();
 sg13g2_fill_1 FILLER_43_244 ();
 sg13g2_fill_1 FILLER_43_254 ();
 sg13g2_decap_4 FILLER_43_281 ();
 sg13g2_decap_4 FILLER_43_293 ();
 sg13g2_fill_2 FILLER_43_297 ();
 sg13g2_decap_4 FILLER_43_315 ();
 sg13g2_fill_1 FILLER_43_319 ();
 sg13g2_decap_8 FILLER_43_346 ();
 sg13g2_fill_2 FILLER_43_353 ();
 sg13g2_fill_1 FILLER_43_370 ();
 sg13g2_decap_8 FILLER_43_424 ();
 sg13g2_decap_8 FILLER_43_456 ();
 sg13g2_fill_2 FILLER_43_463 ();
 sg13g2_fill_2 FILLER_43_483 ();
 sg13g2_fill_1 FILLER_43_485 ();
 sg13g2_decap_8 FILLER_43_499 ();
 sg13g2_fill_2 FILLER_43_506 ();
 sg13g2_fill_2 FILLER_43_527 ();
 sg13g2_fill_2 FILLER_43_582 ();
 sg13g2_fill_1 FILLER_43_584 ();
 sg13g2_decap_4 FILLER_43_635 ();
 sg13g2_decap_4 FILLER_43_647 ();
 sg13g2_fill_2 FILLER_43_651 ();
 sg13g2_decap_8 FILLER_43_657 ();
 sg13g2_fill_1 FILLER_43_664 ();
 sg13g2_fill_1 FILLER_43_678 ();
 sg13g2_decap_4 FILLER_43_705 ();
 sg13g2_fill_1 FILLER_43_709 ();
 sg13g2_fill_2 FILLER_43_718 ();
 sg13g2_fill_1 FILLER_43_720 ();
 sg13g2_fill_2 FILLER_43_742 ();
 sg13g2_fill_1 FILLER_43_744 ();
 sg13g2_fill_1 FILLER_43_750 ();
 sg13g2_fill_2 FILLER_43_769 ();
 sg13g2_fill_1 FILLER_43_797 ();
 sg13g2_fill_2 FILLER_43_807 ();
 sg13g2_decap_4 FILLER_43_895 ();
 sg13g2_fill_2 FILLER_43_899 ();
 sg13g2_decap_4 FILLER_43_906 ();
 sg13g2_decap_8 FILLER_43_914 ();
 sg13g2_decap_8 FILLER_43_921 ();
 sg13g2_fill_1 FILLER_43_928 ();
 sg13g2_fill_2 FILLER_43_958 ();
 sg13g2_fill_1 FILLER_43_991 ();
 sg13g2_fill_1 FILLER_43_1015 ();
 sg13g2_fill_1 FILLER_43_1032 ();
 sg13g2_fill_1 FILLER_43_1068 ();
 sg13g2_fill_1 FILLER_43_1078 ();
 sg13g2_fill_2 FILLER_43_1112 ();
 sg13g2_fill_1 FILLER_43_1213 ();
 sg13g2_fill_1 FILLER_43_1254 ();
 sg13g2_fill_2 FILLER_43_1328 ();
 sg13g2_fill_1 FILLER_43_1374 ();
 sg13g2_fill_1 FILLER_43_1393 ();
 sg13g2_fill_2 FILLER_43_1431 ();
 sg13g2_fill_2 FILLER_43_1490 ();
 sg13g2_fill_1 FILLER_43_1492 ();
 sg13g2_fill_1 FILLER_43_1553 ();
 sg13g2_decap_4 FILLER_43_1585 ();
 sg13g2_fill_2 FILLER_43_1589 ();
 sg13g2_decap_8 FILLER_43_1606 ();
 sg13g2_decap_4 FILLER_43_1613 ();
 sg13g2_decap_8 FILLER_43_1621 ();
 sg13g2_fill_2 FILLER_43_1663 ();
 sg13g2_fill_1 FILLER_43_1665 ();
 sg13g2_fill_2 FILLER_43_1697 ();
 sg13g2_fill_2 FILLER_43_1751 ();
 sg13g2_fill_2 FILLER_43_1762 ();
 sg13g2_fill_2 FILLER_43_1832 ();
 sg13g2_decap_4 FILLER_43_1847 ();
 sg13g2_fill_2 FILLER_43_1851 ();
 sg13g2_fill_1 FILLER_43_1861 ();
 sg13g2_fill_1 FILLER_43_1870 ();
 sg13g2_fill_2 FILLER_43_1887 ();
 sg13g2_fill_1 FILLER_43_1889 ();
 sg13g2_decap_8 FILLER_43_1914 ();
 sg13g2_decap_8 FILLER_43_1921 ();
 sg13g2_fill_1 FILLER_43_1928 ();
 sg13g2_decap_4 FILLER_43_1945 ();
 sg13g2_fill_2 FILLER_43_1949 ();
 sg13g2_decap_8 FILLER_43_1959 ();
 sg13g2_decap_4 FILLER_43_1966 ();
 sg13g2_fill_1 FILLER_43_1970 ();
 sg13g2_decap_4 FILLER_43_2011 ();
 sg13g2_decap_8 FILLER_43_2031 ();
 sg13g2_fill_2 FILLER_43_2054 ();
 sg13g2_fill_2 FILLER_43_2086 ();
 sg13g2_decap_4 FILLER_43_2158 ();
 sg13g2_fill_2 FILLER_43_2203 ();
 sg13g2_fill_1 FILLER_43_2241 ();
 sg13g2_fill_1 FILLER_43_2250 ();
 sg13g2_fill_2 FILLER_43_2313 ();
 sg13g2_fill_1 FILLER_43_2315 ();
 sg13g2_decap_8 FILLER_43_2347 ();
 sg13g2_decap_8 FILLER_43_2354 ();
 sg13g2_decap_8 FILLER_43_2361 ();
 sg13g2_decap_8 FILLER_43_2368 ();
 sg13g2_decap_8 FILLER_43_2375 ();
 sg13g2_decap_8 FILLER_43_2382 ();
 sg13g2_decap_8 FILLER_43_2389 ();
 sg13g2_decap_8 FILLER_43_2396 ();
 sg13g2_decap_8 FILLER_43_2403 ();
 sg13g2_decap_8 FILLER_43_2410 ();
 sg13g2_decap_8 FILLER_43_2417 ();
 sg13g2_decap_8 FILLER_43_2424 ();
 sg13g2_decap_8 FILLER_43_2431 ();
 sg13g2_decap_8 FILLER_43_2438 ();
 sg13g2_decap_8 FILLER_43_2445 ();
 sg13g2_decap_8 FILLER_43_2452 ();
 sg13g2_decap_8 FILLER_43_2459 ();
 sg13g2_decap_8 FILLER_43_2466 ();
 sg13g2_decap_8 FILLER_43_2473 ();
 sg13g2_decap_8 FILLER_43_2480 ();
 sg13g2_decap_8 FILLER_43_2487 ();
 sg13g2_decap_8 FILLER_43_2494 ();
 sg13g2_decap_8 FILLER_43_2501 ();
 sg13g2_decap_8 FILLER_43_2508 ();
 sg13g2_decap_8 FILLER_43_2515 ();
 sg13g2_decap_8 FILLER_43_2522 ();
 sg13g2_decap_8 FILLER_43_2529 ();
 sg13g2_decap_8 FILLER_43_2536 ();
 sg13g2_decap_8 FILLER_43_2543 ();
 sg13g2_decap_8 FILLER_43_2550 ();
 sg13g2_decap_8 FILLER_43_2557 ();
 sg13g2_decap_8 FILLER_43_2564 ();
 sg13g2_decap_8 FILLER_43_2571 ();
 sg13g2_decap_8 FILLER_43_2578 ();
 sg13g2_decap_8 FILLER_43_2585 ();
 sg13g2_decap_8 FILLER_43_2592 ();
 sg13g2_decap_8 FILLER_43_2599 ();
 sg13g2_decap_8 FILLER_43_2606 ();
 sg13g2_decap_8 FILLER_43_2613 ();
 sg13g2_decap_8 FILLER_43_2620 ();
 sg13g2_decap_8 FILLER_43_2627 ();
 sg13g2_decap_8 FILLER_43_2634 ();
 sg13g2_decap_8 FILLER_43_2641 ();
 sg13g2_decap_8 FILLER_43_2648 ();
 sg13g2_decap_8 FILLER_43_2655 ();
 sg13g2_decap_8 FILLER_43_2662 ();
 sg13g2_decap_4 FILLER_43_2669 ();
 sg13g2_fill_1 FILLER_43_2673 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_decap_4 FILLER_44_168 ();
 sg13g2_fill_1 FILLER_44_190 ();
 sg13g2_decap_4 FILLER_44_211 ();
 sg13g2_fill_2 FILLER_44_231 ();
 sg13g2_decap_4 FILLER_44_259 ();
 sg13g2_fill_1 FILLER_44_263 ();
 sg13g2_decap_8 FILLER_44_293 ();
 sg13g2_decap_8 FILLER_44_308 ();
 sg13g2_decap_8 FILLER_44_315 ();
 sg13g2_decap_4 FILLER_44_322 ();
 sg13g2_fill_2 FILLER_44_339 ();
 sg13g2_fill_1 FILLER_44_367 ();
 sg13g2_fill_2 FILLER_44_372 ();
 sg13g2_fill_2 FILLER_44_405 ();
 sg13g2_fill_2 FILLER_44_421 ();
 sg13g2_decap_4 FILLER_44_431 ();
 sg13g2_fill_2 FILLER_44_441 ();
 sg13g2_fill_1 FILLER_44_443 ();
 sg13g2_fill_2 FILLER_44_461 ();
 sg13g2_fill_1 FILLER_44_463 ();
 sg13g2_decap_4 FILLER_44_477 ();
 sg13g2_fill_1 FILLER_44_481 ();
 sg13g2_fill_2 FILLER_44_487 ();
 sg13g2_fill_2 FILLER_44_495 ();
 sg13g2_fill_1 FILLER_44_497 ();
 sg13g2_fill_2 FILLER_44_572 ();
 sg13g2_fill_1 FILLER_44_574 ();
 sg13g2_decap_4 FILLER_44_597 ();
 sg13g2_fill_2 FILLER_44_622 ();
 sg13g2_fill_1 FILLER_44_624 ();
 sg13g2_decap_4 FILLER_44_640 ();
 sg13g2_fill_2 FILLER_44_649 ();
 sg13g2_fill_1 FILLER_44_651 ();
 sg13g2_decap_4 FILLER_44_660 ();
 sg13g2_decap_4 FILLER_44_682 ();
 sg13g2_fill_2 FILLER_44_686 ();
 sg13g2_fill_2 FILLER_44_693 ();
 sg13g2_fill_2 FILLER_44_700 ();
 sg13g2_decap_8 FILLER_44_719 ();
 sg13g2_decap_8 FILLER_44_726 ();
 sg13g2_fill_2 FILLER_44_733 ();
 sg13g2_fill_2 FILLER_44_768 ();
 sg13g2_fill_1 FILLER_44_770 ();
 sg13g2_fill_2 FILLER_44_801 ();
 sg13g2_fill_1 FILLER_44_803 ();
 sg13g2_fill_2 FILLER_44_813 ();
 sg13g2_fill_1 FILLER_44_815 ();
 sg13g2_decap_4 FILLER_44_851 ();
 sg13g2_fill_1 FILLER_44_855 ();
 sg13g2_decap_8 FILLER_44_860 ();
 sg13g2_decap_8 FILLER_44_867 ();
 sg13g2_decap_4 FILLER_44_874 ();
 sg13g2_fill_2 FILLER_44_878 ();
 sg13g2_fill_2 FILLER_44_884 ();
 sg13g2_fill_1 FILLER_44_886 ();
 sg13g2_fill_1 FILLER_44_922 ();
 sg13g2_fill_1 FILLER_44_928 ();
 sg13g2_fill_2 FILLER_44_965 ();
 sg13g2_fill_2 FILLER_44_972 ();
 sg13g2_fill_2 FILLER_44_1100 ();
 sg13g2_fill_2 FILLER_44_1133 ();
 sg13g2_fill_2 FILLER_44_1166 ();
 sg13g2_fill_2 FILLER_44_1319 ();
 sg13g2_fill_1 FILLER_44_1326 ();
 sg13g2_fill_2 FILLER_44_1357 ();
 sg13g2_fill_1 FILLER_44_1404 ();
 sg13g2_fill_2 FILLER_44_1567 ();
 sg13g2_fill_2 FILLER_44_1578 ();
 sg13g2_decap_4 FILLER_44_1593 ();
 sg13g2_decap_4 FILLER_44_1602 ();
 sg13g2_fill_1 FILLER_44_1632 ();
 sg13g2_decap_4 FILLER_44_1646 ();
 sg13g2_fill_1 FILLER_44_1689 ();
 sg13g2_decap_4 FILLER_44_1729 ();
 sg13g2_fill_1 FILLER_44_1733 ();
 sg13g2_decap_8 FILLER_44_1780 ();
 sg13g2_fill_2 FILLER_44_1787 ();
 sg13g2_fill_1 FILLER_44_1789 ();
 sg13g2_decap_8 FILLER_44_1799 ();
 sg13g2_fill_1 FILLER_44_1806 ();
 sg13g2_decap_4 FILLER_44_1832 ();
 sg13g2_fill_1 FILLER_44_1836 ();
 sg13g2_decap_4 FILLER_44_1842 ();
 sg13g2_fill_1 FILLER_44_1850 ();
 sg13g2_decap_4 FILLER_44_1872 ();
 sg13g2_fill_2 FILLER_44_1876 ();
 sg13g2_fill_1 FILLER_44_1918 ();
 sg13g2_fill_2 FILLER_44_1932 ();
 sg13g2_fill_2 FILLER_44_1950 ();
 sg13g2_fill_1 FILLER_44_1952 ();
 sg13g2_decap_4 FILLER_44_1969 ();
 sg13g2_fill_1 FILLER_44_1973 ();
 sg13g2_fill_2 FILLER_44_1998 ();
 sg13g2_decap_8 FILLER_44_2008 ();
 sg13g2_fill_2 FILLER_44_2015 ();
 sg13g2_fill_1 FILLER_44_2017 ();
 sg13g2_decap_4 FILLER_44_2030 ();
 sg13g2_fill_1 FILLER_44_2034 ();
 sg13g2_decap_4 FILLER_44_2060 ();
 sg13g2_fill_2 FILLER_44_2064 ();
 sg13g2_decap_8 FILLER_44_2070 ();
 sg13g2_decap_4 FILLER_44_2077 ();
 sg13g2_fill_1 FILLER_44_2081 ();
 sg13g2_decap_4 FILLER_44_2092 ();
 sg13g2_decap_8 FILLER_44_2109 ();
 sg13g2_fill_1 FILLER_44_2116 ();
 sg13g2_decap_4 FILLER_44_2143 ();
 sg13g2_fill_1 FILLER_44_2157 ();
 sg13g2_fill_2 FILLER_44_2174 ();
 sg13g2_fill_1 FILLER_44_2176 ();
 sg13g2_decap_4 FILLER_44_2194 ();
 sg13g2_decap_4 FILLER_44_2273 ();
 sg13g2_fill_1 FILLER_44_2286 ();
 sg13g2_decap_8 FILLER_44_2304 ();
 sg13g2_fill_1 FILLER_44_2311 ();
 sg13g2_decap_8 FILLER_44_2338 ();
 sg13g2_decap_8 FILLER_44_2345 ();
 sg13g2_decap_8 FILLER_44_2352 ();
 sg13g2_decap_8 FILLER_44_2359 ();
 sg13g2_decap_8 FILLER_44_2366 ();
 sg13g2_decap_8 FILLER_44_2373 ();
 sg13g2_decap_8 FILLER_44_2380 ();
 sg13g2_decap_8 FILLER_44_2387 ();
 sg13g2_decap_8 FILLER_44_2394 ();
 sg13g2_decap_8 FILLER_44_2401 ();
 sg13g2_decap_8 FILLER_44_2408 ();
 sg13g2_decap_8 FILLER_44_2415 ();
 sg13g2_decap_8 FILLER_44_2422 ();
 sg13g2_decap_8 FILLER_44_2429 ();
 sg13g2_decap_8 FILLER_44_2436 ();
 sg13g2_decap_8 FILLER_44_2443 ();
 sg13g2_decap_8 FILLER_44_2450 ();
 sg13g2_decap_8 FILLER_44_2457 ();
 sg13g2_decap_8 FILLER_44_2464 ();
 sg13g2_decap_8 FILLER_44_2471 ();
 sg13g2_decap_8 FILLER_44_2478 ();
 sg13g2_decap_8 FILLER_44_2485 ();
 sg13g2_decap_8 FILLER_44_2492 ();
 sg13g2_decap_8 FILLER_44_2499 ();
 sg13g2_decap_8 FILLER_44_2506 ();
 sg13g2_decap_8 FILLER_44_2513 ();
 sg13g2_decap_8 FILLER_44_2520 ();
 sg13g2_decap_8 FILLER_44_2527 ();
 sg13g2_decap_8 FILLER_44_2534 ();
 sg13g2_decap_8 FILLER_44_2541 ();
 sg13g2_decap_8 FILLER_44_2548 ();
 sg13g2_decap_8 FILLER_44_2555 ();
 sg13g2_decap_8 FILLER_44_2562 ();
 sg13g2_decap_8 FILLER_44_2569 ();
 sg13g2_decap_8 FILLER_44_2576 ();
 sg13g2_decap_8 FILLER_44_2583 ();
 sg13g2_decap_8 FILLER_44_2590 ();
 sg13g2_decap_8 FILLER_44_2597 ();
 sg13g2_decap_8 FILLER_44_2604 ();
 sg13g2_decap_8 FILLER_44_2611 ();
 sg13g2_decap_8 FILLER_44_2618 ();
 sg13g2_decap_8 FILLER_44_2625 ();
 sg13g2_decap_8 FILLER_44_2632 ();
 sg13g2_decap_8 FILLER_44_2639 ();
 sg13g2_decap_8 FILLER_44_2646 ();
 sg13g2_decap_8 FILLER_44_2653 ();
 sg13g2_decap_8 FILLER_44_2660 ();
 sg13g2_decap_8 FILLER_44_2667 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_decap_4 FILLER_45_182 ();
 sg13g2_fill_1 FILLER_45_186 ();
 sg13g2_fill_2 FILLER_45_192 ();
 sg13g2_fill_2 FILLER_45_220 ();
 sg13g2_decap_8 FILLER_45_235 ();
 sg13g2_decap_8 FILLER_45_242 ();
 sg13g2_fill_2 FILLER_45_249 ();
 sg13g2_decap_8 FILLER_45_277 ();
 sg13g2_fill_1 FILLER_45_296 ();
 sg13g2_fill_1 FILLER_45_315 ();
 sg13g2_fill_2 FILLER_45_319 ();
 sg13g2_fill_1 FILLER_45_321 ();
 sg13g2_fill_2 FILLER_45_330 ();
 sg13g2_fill_2 FILLER_45_372 ();
 sg13g2_fill_1 FILLER_45_374 ();
 sg13g2_fill_2 FILLER_45_389 ();
 sg13g2_fill_1 FILLER_45_391 ();
 sg13g2_fill_2 FILLER_45_402 ();
 sg13g2_fill_1 FILLER_45_404 ();
 sg13g2_fill_2 FILLER_45_413 ();
 sg13g2_fill_2 FILLER_45_424 ();
 sg13g2_fill_1 FILLER_45_426 ();
 sg13g2_fill_1 FILLER_45_432 ();
 sg13g2_fill_2 FILLER_45_453 ();
 sg13g2_fill_2 FILLER_45_468 ();
 sg13g2_fill_2 FILLER_45_478 ();
 sg13g2_fill_1 FILLER_45_480 ();
 sg13g2_fill_1 FILLER_45_489 ();
 sg13g2_fill_1 FILLER_45_524 ();
 sg13g2_fill_2 FILLER_45_537 ();
 sg13g2_fill_1 FILLER_45_539 ();
 sg13g2_fill_2 FILLER_45_557 ();
 sg13g2_fill_2 FILLER_45_606 ();
 sg13g2_fill_1 FILLER_45_608 ();
 sg13g2_decap_8 FILLER_45_626 ();
 sg13g2_decap_4 FILLER_45_633 ();
 sg13g2_fill_2 FILLER_45_650 ();
 sg13g2_fill_1 FILLER_45_652 ();
 sg13g2_decap_4 FILLER_45_666 ();
 sg13g2_fill_2 FILLER_45_670 ();
 sg13g2_fill_2 FILLER_45_684 ();
 sg13g2_fill_1 FILLER_45_694 ();
 sg13g2_fill_2 FILLER_45_738 ();
 sg13g2_fill_2 FILLER_45_756 ();
 sg13g2_fill_1 FILLER_45_758 ();
 sg13g2_fill_1 FILLER_45_785 ();
 sg13g2_decap_8 FILLER_45_820 ();
 sg13g2_decap_8 FILLER_45_831 ();
 sg13g2_decap_4 FILLER_45_838 ();
 sg13g2_fill_1 FILLER_45_873 ();
 sg13g2_decap_8 FILLER_45_883 ();
 sg13g2_decap_8 FILLER_45_890 ();
 sg13g2_fill_1 FILLER_45_897 ();
 sg13g2_fill_1 FILLER_45_902 ();
 sg13g2_fill_1 FILLER_45_1057 ();
 sg13g2_fill_2 FILLER_45_1098 ();
 sg13g2_fill_2 FILLER_45_1109 ();
 sg13g2_fill_2 FILLER_45_1120 ();
 sg13g2_fill_1 FILLER_45_1154 ();
 sg13g2_fill_2 FILLER_45_1164 ();
 sg13g2_fill_2 FILLER_45_1195 ();
 sg13g2_fill_1 FILLER_45_1211 ();
 sg13g2_fill_2 FILLER_45_1308 ();
 sg13g2_fill_2 FILLER_45_1357 ();
 sg13g2_fill_2 FILLER_45_1437 ();
 sg13g2_fill_2 FILLER_45_1448 ();
 sg13g2_fill_2 FILLER_45_1524 ();
 sg13g2_fill_2 FILLER_45_1595 ();
 sg13g2_fill_2 FILLER_45_1632 ();
 sg13g2_fill_1 FILLER_45_1643 ();
 sg13g2_fill_2 FILLER_45_1715 ();
 sg13g2_fill_2 FILLER_45_1743 ();
 sg13g2_fill_1 FILLER_45_1745 ();
 sg13g2_fill_1 FILLER_45_1765 ();
 sg13g2_fill_1 FILLER_45_1800 ();
 sg13g2_fill_2 FILLER_45_1832 ();
 sg13g2_fill_1 FILLER_45_1834 ();
 sg13g2_decap_4 FILLER_45_1861 ();
 sg13g2_fill_1 FILLER_45_1870 ();
 sg13g2_decap_8 FILLER_45_1887 ();
 sg13g2_fill_2 FILLER_45_1894 ();
 sg13g2_fill_1 FILLER_45_1896 ();
 sg13g2_decap_8 FILLER_45_1905 ();
 sg13g2_decap_8 FILLER_45_1912 ();
 sg13g2_fill_2 FILLER_45_1919 ();
 sg13g2_fill_2 FILLER_45_1952 ();
 sg13g2_fill_2 FILLER_45_1970 ();
 sg13g2_fill_1 FILLER_45_1972 ();
 sg13g2_decap_8 FILLER_45_1986 ();
 sg13g2_fill_2 FILLER_45_1993 ();
 sg13g2_fill_1 FILLER_45_1995 ();
 sg13g2_fill_2 FILLER_45_2027 ();
 sg13g2_fill_1 FILLER_45_2029 ();
 sg13g2_fill_2 FILLER_45_2049 ();
 sg13g2_fill_1 FILLER_45_2051 ();
 sg13g2_fill_2 FILLER_45_2056 ();
 sg13g2_decap_4 FILLER_45_2084 ();
 sg13g2_fill_1 FILLER_45_2146 ();
 sg13g2_fill_2 FILLER_45_2157 ();
 sg13g2_fill_1 FILLER_45_2169 ();
 sg13g2_fill_2 FILLER_45_2258 ();
 sg13g2_fill_1 FILLER_45_2260 ();
 sg13g2_fill_2 FILLER_45_2273 ();
 sg13g2_fill_1 FILLER_45_2275 ();
 sg13g2_decap_4 FILLER_45_2286 ();
 sg13g2_fill_1 FILLER_45_2290 ();
 sg13g2_decap_4 FILLER_45_2296 ();
 sg13g2_fill_1 FILLER_45_2300 ();
 sg13g2_decap_4 FILLER_45_2311 ();
 sg13g2_fill_2 FILLER_45_2315 ();
 sg13g2_decap_8 FILLER_45_2343 ();
 sg13g2_decap_8 FILLER_45_2350 ();
 sg13g2_decap_8 FILLER_45_2357 ();
 sg13g2_decap_8 FILLER_45_2364 ();
 sg13g2_decap_8 FILLER_45_2371 ();
 sg13g2_decap_8 FILLER_45_2378 ();
 sg13g2_decap_8 FILLER_45_2385 ();
 sg13g2_decap_8 FILLER_45_2392 ();
 sg13g2_decap_8 FILLER_45_2399 ();
 sg13g2_decap_8 FILLER_45_2406 ();
 sg13g2_decap_8 FILLER_45_2413 ();
 sg13g2_decap_8 FILLER_45_2420 ();
 sg13g2_decap_8 FILLER_45_2427 ();
 sg13g2_decap_8 FILLER_45_2434 ();
 sg13g2_decap_8 FILLER_45_2441 ();
 sg13g2_decap_8 FILLER_45_2448 ();
 sg13g2_decap_8 FILLER_45_2455 ();
 sg13g2_decap_8 FILLER_45_2462 ();
 sg13g2_decap_8 FILLER_45_2469 ();
 sg13g2_decap_8 FILLER_45_2476 ();
 sg13g2_decap_8 FILLER_45_2483 ();
 sg13g2_decap_8 FILLER_45_2490 ();
 sg13g2_decap_8 FILLER_45_2497 ();
 sg13g2_decap_8 FILLER_45_2504 ();
 sg13g2_decap_8 FILLER_45_2511 ();
 sg13g2_decap_8 FILLER_45_2518 ();
 sg13g2_decap_8 FILLER_45_2525 ();
 sg13g2_decap_8 FILLER_45_2532 ();
 sg13g2_decap_8 FILLER_45_2539 ();
 sg13g2_decap_8 FILLER_45_2546 ();
 sg13g2_decap_8 FILLER_45_2553 ();
 sg13g2_decap_8 FILLER_45_2560 ();
 sg13g2_decap_8 FILLER_45_2567 ();
 sg13g2_decap_8 FILLER_45_2574 ();
 sg13g2_decap_8 FILLER_45_2581 ();
 sg13g2_decap_8 FILLER_45_2588 ();
 sg13g2_decap_8 FILLER_45_2595 ();
 sg13g2_decap_8 FILLER_45_2602 ();
 sg13g2_decap_8 FILLER_45_2609 ();
 sg13g2_decap_8 FILLER_45_2616 ();
 sg13g2_decap_8 FILLER_45_2623 ();
 sg13g2_decap_8 FILLER_45_2630 ();
 sg13g2_decap_8 FILLER_45_2637 ();
 sg13g2_decap_8 FILLER_45_2644 ();
 sg13g2_decap_8 FILLER_45_2651 ();
 sg13g2_decap_8 FILLER_45_2658 ();
 sg13g2_decap_8 FILLER_45_2665 ();
 sg13g2_fill_2 FILLER_45_2672 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_fill_2 FILLER_46_168 ();
 sg13g2_fill_1 FILLER_46_223 ();
 sg13g2_decap_8 FILLER_46_242 ();
 sg13g2_fill_2 FILLER_46_259 ();
 sg13g2_fill_1 FILLER_46_261 ();
 sg13g2_fill_2 FILLER_46_266 ();
 sg13g2_fill_1 FILLER_46_268 ();
 sg13g2_decap_8 FILLER_46_281 ();
 sg13g2_decap_8 FILLER_46_288 ();
 sg13g2_fill_2 FILLER_46_295 ();
 sg13g2_fill_1 FILLER_46_297 ();
 sg13g2_fill_2 FILLER_46_303 ();
 sg13g2_fill_1 FILLER_46_310 ();
 sg13g2_fill_1 FILLER_46_324 ();
 sg13g2_fill_1 FILLER_46_340 ();
 sg13g2_fill_2 FILLER_46_358 ();
 sg13g2_decap_4 FILLER_46_370 ();
 sg13g2_fill_1 FILLER_46_374 ();
 sg13g2_fill_1 FILLER_46_379 ();
 sg13g2_fill_2 FILLER_46_402 ();
 sg13g2_fill_2 FILLER_46_457 ();
 sg13g2_decap_4 FILLER_46_467 ();
 sg13g2_fill_2 FILLER_46_552 ();
 sg13g2_fill_1 FILLER_46_554 ();
 sg13g2_fill_2 FILLER_46_608 ();
 sg13g2_decap_4 FILLER_46_639 ();
 sg13g2_fill_1 FILLER_46_643 ();
 sg13g2_decap_8 FILLER_46_668 ();
 sg13g2_fill_2 FILLER_46_675 ();
 sg13g2_fill_1 FILLER_46_677 ();
 sg13g2_fill_1 FILLER_46_709 ();
 sg13g2_fill_2 FILLER_46_748 ();
 sg13g2_decap_4 FILLER_46_763 ();
 sg13g2_fill_1 FILLER_46_767 ();
 sg13g2_decap_8 FILLER_46_797 ();
 sg13g2_decap_8 FILLER_46_804 ();
 sg13g2_decap_8 FILLER_46_811 ();
 sg13g2_fill_2 FILLER_46_818 ();
 sg13g2_fill_1 FILLER_46_820 ();
 sg13g2_decap_4 FILLER_46_847 ();
 sg13g2_fill_2 FILLER_46_851 ();
 sg13g2_fill_2 FILLER_46_857 ();
 sg13g2_fill_1 FILLER_46_859 ();
 sg13g2_fill_2 FILLER_46_886 ();
 sg13g2_fill_2 FILLER_46_977 ();
 sg13g2_fill_1 FILLER_46_1028 ();
 sg13g2_fill_2 FILLER_46_1065 ();
 sg13g2_fill_2 FILLER_46_1098 ();
 sg13g2_fill_2 FILLER_46_1165 ();
 sg13g2_fill_1 FILLER_46_1191 ();
 sg13g2_fill_2 FILLER_46_1218 ();
 sg13g2_fill_1 FILLER_46_1283 ();
 sg13g2_fill_1 FILLER_46_1315 ();
 sg13g2_fill_2 FILLER_46_1325 ();
 sg13g2_decap_8 FILLER_46_1362 ();
 sg13g2_fill_2 FILLER_46_1433 ();
 sg13g2_fill_2 FILLER_46_1491 ();
 sg13g2_fill_2 FILLER_46_1522 ();
 sg13g2_fill_1 FILLER_46_1563 ();
 sg13g2_fill_2 FILLER_46_1568 ();
 sg13g2_fill_1 FILLER_46_1591 ();
 sg13g2_decap_4 FILLER_46_1614 ();
 sg13g2_fill_2 FILLER_46_1618 ();
 sg13g2_decap_4 FILLER_46_1786 ();
 sg13g2_fill_1 FILLER_46_1790 ();
 sg13g2_decap_8 FILLER_46_1796 ();
 sg13g2_decap_8 FILLER_46_1813 ();
 sg13g2_fill_2 FILLER_46_1820 ();
 sg13g2_fill_2 FILLER_46_1831 ();
 sg13g2_decap_8 FILLER_46_1842 ();
 sg13g2_decap_8 FILLER_46_1849 ();
 sg13g2_fill_2 FILLER_46_1889 ();
 sg13g2_fill_1 FILLER_46_1891 ();
 sg13g2_fill_2 FILLER_46_1940 ();
 sg13g2_decap_4 FILLER_46_1957 ();
 sg13g2_decap_4 FILLER_46_1988 ();
 sg13g2_fill_1 FILLER_46_1992 ();
 sg13g2_decap_8 FILLER_46_1997 ();
 sg13g2_fill_2 FILLER_46_2004 ();
 sg13g2_fill_1 FILLER_46_2006 ();
 sg13g2_decap_4 FILLER_46_2023 ();
 sg13g2_decap_8 FILLER_46_2032 ();
 sg13g2_fill_2 FILLER_46_2039 ();
 sg13g2_fill_2 FILLER_46_2067 ();
 sg13g2_decap_8 FILLER_46_2073 ();
 sg13g2_fill_2 FILLER_46_2080 ();
 sg13g2_fill_2 FILLER_46_2131 ();
 sg13g2_fill_2 FILLER_46_2178 ();
 sg13g2_fill_1 FILLER_46_2180 ();
 sg13g2_fill_2 FILLER_46_2190 ();
 sg13g2_fill_1 FILLER_46_2192 ();
 sg13g2_fill_1 FILLER_46_2208 ();
 sg13g2_fill_2 FILLER_46_2243 ();
 sg13g2_fill_2 FILLER_46_2255 ();
 sg13g2_fill_2 FILLER_46_2262 ();
 sg13g2_fill_1 FILLER_46_2264 ();
 sg13g2_fill_2 FILLER_46_2280 ();
 sg13g2_fill_1 FILLER_46_2282 ();
 sg13g2_decap_8 FILLER_46_2345 ();
 sg13g2_decap_8 FILLER_46_2352 ();
 sg13g2_decap_8 FILLER_46_2359 ();
 sg13g2_decap_8 FILLER_46_2366 ();
 sg13g2_decap_8 FILLER_46_2373 ();
 sg13g2_decap_8 FILLER_46_2380 ();
 sg13g2_decap_8 FILLER_46_2387 ();
 sg13g2_decap_8 FILLER_46_2394 ();
 sg13g2_decap_8 FILLER_46_2401 ();
 sg13g2_decap_8 FILLER_46_2408 ();
 sg13g2_decap_8 FILLER_46_2415 ();
 sg13g2_decap_8 FILLER_46_2422 ();
 sg13g2_decap_8 FILLER_46_2429 ();
 sg13g2_decap_8 FILLER_46_2436 ();
 sg13g2_decap_8 FILLER_46_2443 ();
 sg13g2_decap_8 FILLER_46_2450 ();
 sg13g2_decap_8 FILLER_46_2457 ();
 sg13g2_decap_8 FILLER_46_2464 ();
 sg13g2_decap_8 FILLER_46_2471 ();
 sg13g2_decap_8 FILLER_46_2478 ();
 sg13g2_decap_8 FILLER_46_2485 ();
 sg13g2_decap_8 FILLER_46_2492 ();
 sg13g2_decap_8 FILLER_46_2499 ();
 sg13g2_decap_8 FILLER_46_2506 ();
 sg13g2_decap_8 FILLER_46_2513 ();
 sg13g2_decap_8 FILLER_46_2520 ();
 sg13g2_decap_8 FILLER_46_2527 ();
 sg13g2_decap_8 FILLER_46_2534 ();
 sg13g2_decap_8 FILLER_46_2541 ();
 sg13g2_decap_8 FILLER_46_2548 ();
 sg13g2_decap_8 FILLER_46_2555 ();
 sg13g2_decap_8 FILLER_46_2562 ();
 sg13g2_decap_8 FILLER_46_2569 ();
 sg13g2_decap_8 FILLER_46_2576 ();
 sg13g2_decap_8 FILLER_46_2583 ();
 sg13g2_decap_8 FILLER_46_2590 ();
 sg13g2_decap_8 FILLER_46_2597 ();
 sg13g2_decap_8 FILLER_46_2604 ();
 sg13g2_decap_8 FILLER_46_2611 ();
 sg13g2_decap_8 FILLER_46_2618 ();
 sg13g2_decap_8 FILLER_46_2625 ();
 sg13g2_decap_8 FILLER_46_2632 ();
 sg13g2_decap_8 FILLER_46_2639 ();
 sg13g2_decap_8 FILLER_46_2646 ();
 sg13g2_decap_8 FILLER_46_2653 ();
 sg13g2_decap_8 FILLER_46_2660 ();
 sg13g2_decap_8 FILLER_46_2667 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_fill_2 FILLER_47_175 ();
 sg13g2_fill_2 FILLER_47_191 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_fill_2 FILLER_47_238 ();
 sg13g2_fill_1 FILLER_47_261 ();
 sg13g2_decap_4 FILLER_47_286 ();
 sg13g2_fill_1 FILLER_47_303 ();
 sg13g2_fill_1 FILLER_47_309 ();
 sg13g2_decap_4 FILLER_47_315 ();
 sg13g2_fill_2 FILLER_47_319 ();
 sg13g2_fill_1 FILLER_47_390 ();
 sg13g2_fill_2 FILLER_47_438 ();
 sg13g2_fill_1 FILLER_47_440 ();
 sg13g2_fill_1 FILLER_47_450 ();
 sg13g2_fill_2 FILLER_47_456 ();
 sg13g2_fill_2 FILLER_47_464 ();
 sg13g2_fill_1 FILLER_47_466 ();
 sg13g2_fill_1 FILLER_47_475 ();
 sg13g2_decap_8 FILLER_47_528 ();
 sg13g2_fill_2 FILLER_47_535 ();
 sg13g2_decap_4 FILLER_47_541 ();
 sg13g2_fill_1 FILLER_47_545 ();
 sg13g2_fill_2 FILLER_47_576 ();
 sg13g2_fill_1 FILLER_47_578 ();
 sg13g2_decap_8 FILLER_47_631 ();
 sg13g2_decap_4 FILLER_47_638 ();
 sg13g2_fill_2 FILLER_47_642 ();
 sg13g2_fill_1 FILLER_47_652 ();
 sg13g2_fill_2 FILLER_47_657 ();
 sg13g2_fill_2 FILLER_47_712 ();
 sg13g2_fill_2 FILLER_47_722 ();
 sg13g2_fill_2 FILLER_47_744 ();
 sg13g2_fill_1 FILLER_47_746 ();
 sg13g2_fill_2 FILLER_47_773 ();
 sg13g2_fill_2 FILLER_47_783 ();
 sg13g2_fill_1 FILLER_47_785 ();
 sg13g2_decap_8 FILLER_47_791 ();
 sg13g2_fill_2 FILLER_47_811 ();
 sg13g2_fill_2 FILLER_47_839 ();
 sg13g2_fill_1 FILLER_47_841 ();
 sg13g2_fill_2 FILLER_47_868 ();
 sg13g2_fill_1 FILLER_47_905 ();
 sg13g2_fill_2 FILLER_47_973 ();
 sg13g2_fill_1 FILLER_47_1020 ();
 sg13g2_fill_2 FILLER_47_1136 ();
 sg13g2_fill_1 FILLER_47_1230 ();
 sg13g2_fill_2 FILLER_47_1256 ();
 sg13g2_fill_2 FILLER_47_1289 ();
 sg13g2_fill_2 FILLER_47_1299 ();
 sg13g2_fill_1 FILLER_47_1354 ();
 sg13g2_fill_1 FILLER_47_1414 ();
 sg13g2_fill_2 FILLER_47_1573 ();
 sg13g2_fill_1 FILLER_47_1605 ();
 sg13g2_decap_4 FILLER_47_1623 ();
 sg13g2_fill_1 FILLER_47_1627 ();
 sg13g2_fill_2 FILLER_47_1636 ();
 sg13g2_fill_2 FILLER_47_1709 ();
 sg13g2_fill_1 FILLER_47_1711 ();
 sg13g2_fill_1 FILLER_47_1738 ();
 sg13g2_fill_2 FILLER_47_1749 ();
 sg13g2_fill_1 FILLER_47_1786 ();
 sg13g2_fill_2 FILLER_47_1813 ();
 sg13g2_fill_1 FILLER_47_1815 ();
 sg13g2_fill_1 FILLER_47_1820 ();
 sg13g2_fill_2 FILLER_47_1873 ();
 sg13g2_fill_1 FILLER_47_1875 ();
 sg13g2_fill_2 FILLER_47_1892 ();
 sg13g2_decap_8 FILLER_47_1902 ();
 sg13g2_fill_2 FILLER_47_1909 ();
 sg13g2_fill_1 FILLER_47_1911 ();
 sg13g2_fill_2 FILLER_47_1933 ();
 sg13g2_decap_8 FILLER_47_1950 ();
 sg13g2_decap_8 FILLER_47_1961 ();
 sg13g2_decap_4 FILLER_47_1968 ();
 sg13g2_fill_1 FILLER_47_1972 ();
 sg13g2_fill_2 FILLER_47_1981 ();
 sg13g2_decap_8 FILLER_47_2014 ();
 sg13g2_fill_2 FILLER_47_2021 ();
 sg13g2_decap_4 FILLER_47_2056 ();
 sg13g2_fill_1 FILLER_47_2060 ();
 sg13g2_fill_2 FILLER_47_2065 ();
 sg13g2_fill_1 FILLER_47_2067 ();
 sg13g2_decap_4 FILLER_47_2125 ();
 sg13g2_fill_2 FILLER_47_2144 ();
 sg13g2_fill_1 FILLER_47_2146 ();
 sg13g2_fill_2 FILLER_47_2172 ();
 sg13g2_fill_2 FILLER_47_2200 ();
 sg13g2_fill_1 FILLER_47_2202 ();
 sg13g2_fill_2 FILLER_47_2240 ();
 sg13g2_fill_1 FILLER_47_2242 ();
 sg13g2_fill_1 FILLER_47_2253 ();
 sg13g2_fill_2 FILLER_47_2279 ();
 sg13g2_fill_1 FILLER_47_2281 ();
 sg13g2_decap_4 FILLER_47_2299 ();
 sg13g2_fill_2 FILLER_47_2303 ();
 sg13g2_fill_2 FILLER_47_2315 ();
 sg13g2_decap_8 FILLER_47_2343 ();
 sg13g2_decap_8 FILLER_47_2350 ();
 sg13g2_decap_8 FILLER_47_2357 ();
 sg13g2_decap_8 FILLER_47_2364 ();
 sg13g2_decap_8 FILLER_47_2371 ();
 sg13g2_decap_8 FILLER_47_2378 ();
 sg13g2_decap_8 FILLER_47_2385 ();
 sg13g2_decap_8 FILLER_47_2392 ();
 sg13g2_decap_8 FILLER_47_2399 ();
 sg13g2_decap_8 FILLER_47_2406 ();
 sg13g2_decap_8 FILLER_47_2413 ();
 sg13g2_decap_8 FILLER_47_2420 ();
 sg13g2_decap_8 FILLER_47_2427 ();
 sg13g2_decap_8 FILLER_47_2434 ();
 sg13g2_decap_8 FILLER_47_2441 ();
 sg13g2_decap_8 FILLER_47_2448 ();
 sg13g2_decap_8 FILLER_47_2455 ();
 sg13g2_decap_8 FILLER_47_2462 ();
 sg13g2_decap_8 FILLER_47_2469 ();
 sg13g2_decap_8 FILLER_47_2476 ();
 sg13g2_decap_8 FILLER_47_2483 ();
 sg13g2_decap_8 FILLER_47_2490 ();
 sg13g2_decap_8 FILLER_47_2497 ();
 sg13g2_decap_8 FILLER_47_2504 ();
 sg13g2_decap_8 FILLER_47_2511 ();
 sg13g2_decap_8 FILLER_47_2518 ();
 sg13g2_decap_8 FILLER_47_2525 ();
 sg13g2_decap_8 FILLER_47_2532 ();
 sg13g2_decap_8 FILLER_47_2539 ();
 sg13g2_decap_8 FILLER_47_2546 ();
 sg13g2_decap_8 FILLER_47_2553 ();
 sg13g2_decap_8 FILLER_47_2560 ();
 sg13g2_decap_8 FILLER_47_2567 ();
 sg13g2_decap_8 FILLER_47_2574 ();
 sg13g2_decap_8 FILLER_47_2581 ();
 sg13g2_decap_8 FILLER_47_2588 ();
 sg13g2_decap_8 FILLER_47_2595 ();
 sg13g2_decap_8 FILLER_47_2602 ();
 sg13g2_decap_8 FILLER_47_2609 ();
 sg13g2_decap_8 FILLER_47_2616 ();
 sg13g2_decap_8 FILLER_47_2623 ();
 sg13g2_decap_8 FILLER_47_2630 ();
 sg13g2_decap_8 FILLER_47_2637 ();
 sg13g2_decap_8 FILLER_47_2644 ();
 sg13g2_decap_8 FILLER_47_2651 ();
 sg13g2_decap_8 FILLER_47_2658 ();
 sg13g2_decap_8 FILLER_47_2665 ();
 sg13g2_fill_2 FILLER_47_2672 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_4 FILLER_48_168 ();
 sg13g2_fill_1 FILLER_48_172 ();
 sg13g2_fill_2 FILLER_48_177 ();
 sg13g2_fill_1 FILLER_48_179 ();
 sg13g2_fill_2 FILLER_48_202 ();
 sg13g2_decap_4 FILLER_48_213 ();
 sg13g2_fill_2 FILLER_48_217 ();
 sg13g2_fill_2 FILLER_48_241 ();
 sg13g2_fill_1 FILLER_48_243 ();
 sg13g2_decap_8 FILLER_48_261 ();
 sg13g2_fill_2 FILLER_48_281 ();
 sg13g2_fill_1 FILLER_48_283 ();
 sg13g2_fill_2 FILLER_48_308 ();
 sg13g2_fill_2 FILLER_48_319 ();
 sg13g2_fill_2 FILLER_48_337 ();
 sg13g2_fill_1 FILLER_48_370 ();
 sg13g2_fill_2 FILLER_48_385 ();
 sg13g2_fill_1 FILLER_48_387 ();
 sg13g2_fill_1 FILLER_48_437 ();
 sg13g2_fill_2 FILLER_48_463 ();
 sg13g2_fill_1 FILLER_48_465 ();
 sg13g2_fill_1 FILLER_48_506 ();
 sg13g2_decap_4 FILLER_48_512 ();
 sg13g2_fill_2 FILLER_48_516 ();
 sg13g2_fill_1 FILLER_48_595 ();
 sg13g2_fill_1 FILLER_48_631 ();
 sg13g2_fill_2 FILLER_48_653 ();
 sg13g2_decap_8 FILLER_48_676 ();
 sg13g2_fill_2 FILLER_48_730 ();
 sg13g2_fill_1 FILLER_48_732 ();
 sg13g2_fill_2 FILLER_48_746 ();
 sg13g2_decap_8 FILLER_48_769 ();
 sg13g2_fill_1 FILLER_48_785 ();
 sg13g2_decap_8 FILLER_48_812 ();
 sg13g2_fill_1 FILLER_48_819 ();
 sg13g2_fill_2 FILLER_48_837 ();
 sg13g2_fill_1 FILLER_48_839 ();
 sg13g2_fill_2 FILLER_48_849 ();
 sg13g2_fill_1 FILLER_48_943 ();
 sg13g2_fill_2 FILLER_48_1055 ();
 sg13g2_fill_1 FILLER_48_1118 ();
 sg13g2_fill_1 FILLER_48_1125 ();
 sg13g2_fill_1 FILLER_48_1140 ();
 sg13g2_fill_2 FILLER_48_1439 ();
 sg13g2_fill_1 FILLER_48_1447 ();
 sg13g2_fill_1 FILLER_48_1488 ();
 sg13g2_fill_2 FILLER_48_1565 ();
 sg13g2_fill_1 FILLER_48_1577 ();
 sg13g2_fill_1 FILLER_48_1632 ();
 sg13g2_fill_2 FILLER_48_1679 ();
 sg13g2_fill_1 FILLER_48_1681 ();
 sg13g2_fill_1 FILLER_48_1708 ();
 sg13g2_fill_2 FILLER_48_1796 ();
 sg13g2_decap_8 FILLER_48_1802 ();
 sg13g2_fill_2 FILLER_48_1809 ();
 sg13g2_decap_8 FILLER_48_1832 ();
 sg13g2_fill_1 FILLER_48_1859 ();
 sg13g2_decap_8 FILLER_48_1873 ();
 sg13g2_decap_8 FILLER_48_1885 ();
 sg13g2_decap_4 FILLER_48_1892 ();
 sg13g2_decap_8 FILLER_48_1909 ();
 sg13g2_decap_8 FILLER_48_1920 ();
 sg13g2_fill_2 FILLER_48_1927 ();
 sg13g2_decap_8 FILLER_48_1977 ();
 sg13g2_decap_4 FILLER_48_1984 ();
 sg13g2_fill_2 FILLER_48_1988 ();
 sg13g2_fill_2 FILLER_48_1994 ();
 sg13g2_fill_1 FILLER_48_1996 ();
 sg13g2_fill_2 FILLER_48_2010 ();
 sg13g2_fill_2 FILLER_48_2038 ();
 sg13g2_fill_1 FILLER_48_2040 ();
 sg13g2_decap_4 FILLER_48_2076 ();
 sg13g2_fill_1 FILLER_48_2101 ();
 sg13g2_fill_2 FILLER_48_2123 ();
 sg13g2_fill_2 FILLER_48_2135 ();
 sg13g2_fill_1 FILLER_48_2145 ();
 sg13g2_fill_1 FILLER_48_2160 ();
 sg13g2_fill_2 FILLER_48_2186 ();
 sg13g2_fill_1 FILLER_48_2188 ();
 sg13g2_fill_1 FILLER_48_2198 ();
 sg13g2_decap_8 FILLER_48_2204 ();
 sg13g2_fill_2 FILLER_48_2211 ();
 sg13g2_decap_4 FILLER_48_2218 ();
 sg13g2_decap_4 FILLER_48_2302 ();
 sg13g2_fill_1 FILLER_48_2306 ();
 sg13g2_decap_8 FILLER_48_2346 ();
 sg13g2_decap_8 FILLER_48_2353 ();
 sg13g2_decap_8 FILLER_48_2360 ();
 sg13g2_decap_8 FILLER_48_2367 ();
 sg13g2_decap_8 FILLER_48_2374 ();
 sg13g2_decap_8 FILLER_48_2381 ();
 sg13g2_decap_8 FILLER_48_2388 ();
 sg13g2_decap_8 FILLER_48_2395 ();
 sg13g2_decap_8 FILLER_48_2402 ();
 sg13g2_decap_8 FILLER_48_2409 ();
 sg13g2_decap_8 FILLER_48_2416 ();
 sg13g2_decap_8 FILLER_48_2423 ();
 sg13g2_decap_8 FILLER_48_2430 ();
 sg13g2_decap_8 FILLER_48_2437 ();
 sg13g2_decap_8 FILLER_48_2444 ();
 sg13g2_decap_8 FILLER_48_2451 ();
 sg13g2_decap_8 FILLER_48_2458 ();
 sg13g2_decap_8 FILLER_48_2465 ();
 sg13g2_decap_8 FILLER_48_2472 ();
 sg13g2_decap_8 FILLER_48_2479 ();
 sg13g2_decap_8 FILLER_48_2486 ();
 sg13g2_decap_8 FILLER_48_2493 ();
 sg13g2_decap_8 FILLER_48_2500 ();
 sg13g2_decap_8 FILLER_48_2507 ();
 sg13g2_decap_8 FILLER_48_2514 ();
 sg13g2_decap_8 FILLER_48_2521 ();
 sg13g2_decap_8 FILLER_48_2528 ();
 sg13g2_decap_8 FILLER_48_2535 ();
 sg13g2_decap_8 FILLER_48_2542 ();
 sg13g2_decap_8 FILLER_48_2549 ();
 sg13g2_decap_8 FILLER_48_2556 ();
 sg13g2_decap_8 FILLER_48_2563 ();
 sg13g2_decap_8 FILLER_48_2570 ();
 sg13g2_decap_8 FILLER_48_2577 ();
 sg13g2_decap_8 FILLER_48_2584 ();
 sg13g2_decap_8 FILLER_48_2591 ();
 sg13g2_decap_8 FILLER_48_2598 ();
 sg13g2_decap_8 FILLER_48_2605 ();
 sg13g2_decap_8 FILLER_48_2612 ();
 sg13g2_decap_8 FILLER_48_2619 ();
 sg13g2_decap_8 FILLER_48_2626 ();
 sg13g2_decap_8 FILLER_48_2633 ();
 sg13g2_decap_8 FILLER_48_2640 ();
 sg13g2_decap_8 FILLER_48_2647 ();
 sg13g2_decap_8 FILLER_48_2654 ();
 sg13g2_decap_8 FILLER_48_2661 ();
 sg13g2_decap_4 FILLER_48_2668 ();
 sg13g2_fill_2 FILLER_48_2672 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_decap_8 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_154 ();
 sg13g2_fill_1 FILLER_49_161 ();
 sg13g2_fill_2 FILLER_49_188 ();
 sg13g2_fill_1 FILLER_49_190 ();
 sg13g2_fill_2 FILLER_49_215 ();
 sg13g2_fill_2 FILLER_49_235 ();
 sg13g2_fill_1 FILLER_49_237 ();
 sg13g2_decap_4 FILLER_49_243 ();
 sg13g2_decap_8 FILLER_49_260 ();
 sg13g2_fill_1 FILLER_49_267 ();
 sg13g2_fill_1 FILLER_49_272 ();
 sg13g2_decap_4 FILLER_49_286 ();
 sg13g2_fill_2 FILLER_49_290 ();
 sg13g2_fill_2 FILLER_49_297 ();
 sg13g2_fill_1 FILLER_49_334 ();
 sg13g2_fill_1 FILLER_49_348 ();
 sg13g2_fill_2 FILLER_49_364 ();
 sg13g2_fill_2 FILLER_49_396 ();
 sg13g2_fill_1 FILLER_49_407 ();
 sg13g2_fill_2 FILLER_49_463 ();
 sg13g2_fill_1 FILLER_49_473 ();
 sg13g2_fill_2 FILLER_49_594 ();
 sg13g2_fill_2 FILLER_49_604 ();
 sg13g2_fill_1 FILLER_49_623 ();
 sg13g2_fill_2 FILLER_49_634 ();
 sg13g2_fill_2 FILLER_49_674 ();
 sg13g2_fill_1 FILLER_49_676 ();
 sg13g2_decap_4 FILLER_49_685 ();
 sg13g2_fill_1 FILLER_49_689 ();
 sg13g2_decap_8 FILLER_49_695 ();
 sg13g2_decap_8 FILLER_49_702 ();
 sg13g2_fill_2 FILLER_49_709 ();
 sg13g2_fill_1 FILLER_49_711 ();
 sg13g2_fill_2 FILLER_49_717 ();
 sg13g2_fill_1 FILLER_49_719 ();
 sg13g2_decap_8 FILLER_49_762 ();
 sg13g2_fill_2 FILLER_49_795 ();
 sg13g2_decap_8 FILLER_49_801 ();
 sg13g2_fill_2 FILLER_49_808 ();
 sg13g2_fill_1 FILLER_49_810 ();
 sg13g2_decap_4 FILLER_49_816 ();
 sg13g2_fill_2 FILLER_49_820 ();
 sg13g2_fill_2 FILLER_49_837 ();
 sg13g2_fill_1 FILLER_49_839 ();
 sg13g2_fill_2 FILLER_49_858 ();
 sg13g2_fill_1 FILLER_49_877 ();
 sg13g2_fill_1 FILLER_49_891 ();
 sg13g2_fill_2 FILLER_49_942 ();
 sg13g2_fill_1 FILLER_49_953 ();
 sg13g2_fill_1 FILLER_49_994 ();
 sg13g2_fill_2 FILLER_49_1028 ();
 sg13g2_fill_1 FILLER_49_1048 ();
 sg13g2_fill_2 FILLER_49_1069 ();
 sg13g2_fill_2 FILLER_49_1085 ();
 sg13g2_fill_1 FILLER_49_1096 ();
 sg13g2_fill_1 FILLER_49_1111 ();
 sg13g2_fill_1 FILLER_49_1152 ();
 sg13g2_fill_1 FILLER_49_1191 ();
 sg13g2_fill_2 FILLER_49_1201 ();
 sg13g2_fill_1 FILLER_49_1203 ();
 sg13g2_fill_1 FILLER_49_1305 ();
 sg13g2_fill_2 FILLER_49_1367 ();
 sg13g2_fill_2 FILLER_49_1408 ();
 sg13g2_fill_1 FILLER_49_1518 ();
 sg13g2_fill_1 FILLER_49_1571 ();
 sg13g2_fill_1 FILLER_49_1613 ();
 sg13g2_fill_1 FILLER_49_1628 ();
 sg13g2_fill_1 FILLER_49_1638 ();
 sg13g2_fill_2 FILLER_49_1737 ();
 sg13g2_fill_1 FILLER_49_1739 ();
 sg13g2_fill_1 FILLER_49_1768 ();
 sg13g2_decap_4 FILLER_49_1817 ();
 sg13g2_fill_1 FILLER_49_1821 ();
 sg13g2_fill_2 FILLER_49_1830 ();
 sg13g2_fill_1 FILLER_49_1837 ();
 sg13g2_decap_4 FILLER_49_1873 ();
 sg13g2_fill_2 FILLER_49_1877 ();
 sg13g2_fill_2 FILLER_49_1948 ();
 sg13g2_fill_1 FILLER_49_1950 ();
 sg13g2_fill_1 FILLER_49_1958 ();
 sg13g2_fill_2 FILLER_49_1963 ();
 sg13g2_fill_1 FILLER_49_1965 ();
 sg13g2_decap_8 FILLER_49_2013 ();
 sg13g2_decap_8 FILLER_49_2020 ();
 sg13g2_decap_4 FILLER_49_2027 ();
 sg13g2_decap_4 FILLER_49_2057 ();
 sg13g2_fill_2 FILLER_49_2061 ();
 sg13g2_decap_4 FILLER_49_2071 ();
 sg13g2_fill_1 FILLER_49_2075 ();
 sg13g2_fill_2 FILLER_49_2116 ();
 sg13g2_fill_1 FILLER_49_2118 ();
 sg13g2_fill_2 FILLER_49_2127 ();
 sg13g2_fill_1 FILLER_49_2129 ();
 sg13g2_fill_2 FILLER_49_2181 ();
 sg13g2_decap_8 FILLER_49_2212 ();
 sg13g2_fill_2 FILLER_49_2223 ();
 sg13g2_fill_1 FILLER_49_2225 ();
 sg13g2_decap_8 FILLER_49_2243 ();
 sg13g2_fill_2 FILLER_49_2283 ();
 sg13g2_fill_1 FILLER_49_2285 ();
 sg13g2_fill_1 FILLER_49_2306 ();
 sg13g2_decap_8 FILLER_49_2333 ();
 sg13g2_decap_8 FILLER_49_2340 ();
 sg13g2_decap_8 FILLER_49_2347 ();
 sg13g2_decap_8 FILLER_49_2354 ();
 sg13g2_decap_8 FILLER_49_2361 ();
 sg13g2_decap_8 FILLER_49_2368 ();
 sg13g2_decap_8 FILLER_49_2375 ();
 sg13g2_decap_8 FILLER_49_2382 ();
 sg13g2_decap_8 FILLER_49_2389 ();
 sg13g2_decap_8 FILLER_49_2396 ();
 sg13g2_decap_8 FILLER_49_2403 ();
 sg13g2_decap_8 FILLER_49_2410 ();
 sg13g2_decap_8 FILLER_49_2417 ();
 sg13g2_decap_8 FILLER_49_2424 ();
 sg13g2_decap_8 FILLER_49_2431 ();
 sg13g2_decap_8 FILLER_49_2438 ();
 sg13g2_decap_8 FILLER_49_2445 ();
 sg13g2_decap_8 FILLER_49_2452 ();
 sg13g2_decap_8 FILLER_49_2459 ();
 sg13g2_decap_8 FILLER_49_2466 ();
 sg13g2_decap_8 FILLER_49_2473 ();
 sg13g2_decap_8 FILLER_49_2480 ();
 sg13g2_decap_8 FILLER_49_2487 ();
 sg13g2_decap_8 FILLER_49_2494 ();
 sg13g2_decap_8 FILLER_49_2501 ();
 sg13g2_decap_8 FILLER_49_2508 ();
 sg13g2_decap_8 FILLER_49_2515 ();
 sg13g2_decap_8 FILLER_49_2522 ();
 sg13g2_decap_8 FILLER_49_2529 ();
 sg13g2_decap_8 FILLER_49_2536 ();
 sg13g2_decap_8 FILLER_49_2543 ();
 sg13g2_decap_8 FILLER_49_2550 ();
 sg13g2_decap_8 FILLER_49_2557 ();
 sg13g2_decap_8 FILLER_49_2564 ();
 sg13g2_decap_8 FILLER_49_2571 ();
 sg13g2_decap_8 FILLER_49_2578 ();
 sg13g2_decap_8 FILLER_49_2585 ();
 sg13g2_decap_8 FILLER_49_2592 ();
 sg13g2_decap_8 FILLER_49_2599 ();
 sg13g2_decap_8 FILLER_49_2606 ();
 sg13g2_decap_8 FILLER_49_2613 ();
 sg13g2_decap_8 FILLER_49_2620 ();
 sg13g2_decap_8 FILLER_49_2627 ();
 sg13g2_decap_8 FILLER_49_2634 ();
 sg13g2_decap_8 FILLER_49_2641 ();
 sg13g2_decap_8 FILLER_49_2648 ();
 sg13g2_decap_8 FILLER_49_2655 ();
 sg13g2_decap_8 FILLER_49_2662 ();
 sg13g2_decap_4 FILLER_49_2669 ();
 sg13g2_fill_1 FILLER_49_2673 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_8 FILLER_50_126 ();
 sg13g2_decap_8 FILLER_50_133 ();
 sg13g2_decap_8 FILLER_50_140 ();
 sg13g2_decap_8 FILLER_50_147 ();
 sg13g2_decap_8 FILLER_50_154 ();
 sg13g2_decap_8 FILLER_50_161 ();
 sg13g2_fill_1 FILLER_50_168 ();
 sg13g2_fill_2 FILLER_50_182 ();
 sg13g2_fill_1 FILLER_50_184 ();
 sg13g2_fill_2 FILLER_50_198 ();
 sg13g2_fill_1 FILLER_50_200 ();
 sg13g2_fill_2 FILLER_50_206 ();
 sg13g2_fill_1 FILLER_50_216 ();
 sg13g2_fill_2 FILLER_50_226 ();
 sg13g2_fill_1 FILLER_50_228 ();
 sg13g2_fill_2 FILLER_50_302 ();
 sg13g2_fill_1 FILLER_50_304 ();
 sg13g2_fill_2 FILLER_50_314 ();
 sg13g2_fill_2 FILLER_50_366 ();
 sg13g2_fill_1 FILLER_50_368 ();
 sg13g2_fill_2 FILLER_50_397 ();
 sg13g2_fill_2 FILLER_50_409 ();
 sg13g2_fill_1 FILLER_50_416 ();
 sg13g2_fill_2 FILLER_50_422 ();
 sg13g2_fill_1 FILLER_50_424 ();
 sg13g2_fill_2 FILLER_50_451 ();
 sg13g2_decap_4 FILLER_50_458 ();
 sg13g2_fill_1 FILLER_50_503 ();
 sg13g2_decap_8 FILLER_50_517 ();
 sg13g2_fill_1 FILLER_50_552 ();
 sg13g2_fill_1 FILLER_50_563 ();
 sg13g2_fill_1 FILLER_50_602 ();
 sg13g2_decap_8 FILLER_50_634 ();
 sg13g2_decap_4 FILLER_50_641 ();
 sg13g2_fill_2 FILLER_50_649 ();
 sg13g2_fill_1 FILLER_50_651 ();
 sg13g2_decap_4 FILLER_50_662 ();
 sg13g2_fill_2 FILLER_50_666 ();
 sg13g2_decap_4 FILLER_50_673 ();
 sg13g2_fill_2 FILLER_50_697 ();
 sg13g2_fill_2 FILLER_50_749 ();
 sg13g2_decap_4 FILLER_50_772 ();
 sg13g2_fill_2 FILLER_50_785 ();
 sg13g2_fill_1 FILLER_50_787 ();
 sg13g2_decap_4 FILLER_50_794 ();
 sg13g2_fill_1 FILLER_50_798 ();
 sg13g2_fill_2 FILLER_50_818 ();
 sg13g2_fill_2 FILLER_50_833 ();
 sg13g2_fill_1 FILLER_50_835 ();
 sg13g2_fill_2 FILLER_50_846 ();
 sg13g2_fill_1 FILLER_50_848 ();
 sg13g2_fill_2 FILLER_50_862 ();
 sg13g2_fill_1 FILLER_50_872 ();
 sg13g2_fill_2 FILLER_50_881 ();
 sg13g2_fill_2 FILLER_50_911 ();
 sg13g2_fill_2 FILLER_50_939 ();
 sg13g2_fill_1 FILLER_50_1011 ();
 sg13g2_fill_2 FILLER_50_1032 ();
 sg13g2_fill_1 FILLER_50_1097 ();
 sg13g2_fill_1 FILLER_50_1124 ();
 sg13g2_fill_1 FILLER_50_1179 ();
 sg13g2_fill_1 FILLER_50_1241 ();
 sg13g2_fill_1 FILLER_50_1316 ();
 sg13g2_fill_1 FILLER_50_1336 ();
 sg13g2_fill_2 FILLER_50_1346 ();
 sg13g2_fill_1 FILLER_50_1374 ();
 sg13g2_fill_1 FILLER_50_1447 ();
 sg13g2_fill_1 FILLER_50_1510 ();
 sg13g2_fill_1 FILLER_50_1553 ();
 sg13g2_fill_1 FILLER_50_1567 ();
 sg13g2_fill_1 FILLER_50_1582 ();
 sg13g2_fill_2 FILLER_50_1604 ();
 sg13g2_fill_2 FILLER_50_1632 ();
 sg13g2_fill_1 FILLER_50_1719 ();
 sg13g2_fill_2 FILLER_50_1759 ();
 sg13g2_fill_1 FILLER_50_1766 ();
 sg13g2_fill_1 FILLER_50_1778 ();
 sg13g2_decap_4 FILLER_50_1816 ();
 sg13g2_fill_1 FILLER_50_1820 ();
 sg13g2_decap_4 FILLER_50_1829 ();
 sg13g2_fill_1 FILLER_50_1833 ();
 sg13g2_decap_4 FILLER_50_1839 ();
 sg13g2_fill_1 FILLER_50_1843 ();
 sg13g2_fill_2 FILLER_50_1849 ();
 sg13g2_fill_1 FILLER_50_1851 ();
 sg13g2_decap_8 FILLER_50_1856 ();
 sg13g2_decap_4 FILLER_50_1863 ();
 sg13g2_decap_8 FILLER_50_1871 ();
 sg13g2_fill_1 FILLER_50_1878 ();
 sg13g2_fill_2 FILLER_50_1892 ();
 sg13g2_fill_1 FILLER_50_1894 ();
 sg13g2_fill_2 FILLER_50_1898 ();
 sg13g2_decap_4 FILLER_50_1908 ();
 sg13g2_decap_8 FILLER_50_1920 ();
 sg13g2_fill_2 FILLER_50_1927 ();
 sg13g2_fill_1 FILLER_50_1942 ();
 sg13g2_fill_2 FILLER_50_1969 ();
 sg13g2_decap_4 FILLER_50_1983 ();
 sg13g2_decap_4 FILLER_50_1991 ();
 sg13g2_fill_2 FILLER_50_2008 ();
 sg13g2_fill_1 FILLER_50_2010 ();
 sg13g2_decap_4 FILLER_50_2019 ();
 sg13g2_fill_2 FILLER_50_2036 ();
 sg13g2_decap_8 FILLER_50_2128 ();
 sg13g2_fill_2 FILLER_50_2135 ();
 sg13g2_fill_1 FILLER_50_2137 ();
 sg13g2_fill_1 FILLER_50_2142 ();
 sg13g2_fill_1 FILLER_50_2180 ();
 sg13g2_fill_1 FILLER_50_2244 ();
 sg13g2_decap_8 FILLER_50_2336 ();
 sg13g2_decap_8 FILLER_50_2343 ();
 sg13g2_decap_8 FILLER_50_2350 ();
 sg13g2_decap_8 FILLER_50_2357 ();
 sg13g2_decap_8 FILLER_50_2364 ();
 sg13g2_decap_8 FILLER_50_2371 ();
 sg13g2_decap_8 FILLER_50_2378 ();
 sg13g2_decap_8 FILLER_50_2385 ();
 sg13g2_decap_8 FILLER_50_2392 ();
 sg13g2_decap_8 FILLER_50_2399 ();
 sg13g2_decap_8 FILLER_50_2406 ();
 sg13g2_decap_8 FILLER_50_2413 ();
 sg13g2_decap_8 FILLER_50_2420 ();
 sg13g2_decap_8 FILLER_50_2427 ();
 sg13g2_decap_8 FILLER_50_2434 ();
 sg13g2_decap_8 FILLER_50_2441 ();
 sg13g2_decap_8 FILLER_50_2448 ();
 sg13g2_decap_8 FILLER_50_2455 ();
 sg13g2_decap_8 FILLER_50_2462 ();
 sg13g2_decap_8 FILLER_50_2469 ();
 sg13g2_decap_8 FILLER_50_2476 ();
 sg13g2_decap_8 FILLER_50_2483 ();
 sg13g2_decap_8 FILLER_50_2490 ();
 sg13g2_decap_8 FILLER_50_2497 ();
 sg13g2_decap_8 FILLER_50_2504 ();
 sg13g2_decap_8 FILLER_50_2511 ();
 sg13g2_decap_8 FILLER_50_2518 ();
 sg13g2_decap_8 FILLER_50_2525 ();
 sg13g2_decap_8 FILLER_50_2532 ();
 sg13g2_decap_8 FILLER_50_2539 ();
 sg13g2_decap_8 FILLER_50_2546 ();
 sg13g2_decap_8 FILLER_50_2553 ();
 sg13g2_decap_8 FILLER_50_2560 ();
 sg13g2_decap_8 FILLER_50_2567 ();
 sg13g2_decap_8 FILLER_50_2574 ();
 sg13g2_decap_8 FILLER_50_2581 ();
 sg13g2_decap_8 FILLER_50_2588 ();
 sg13g2_decap_8 FILLER_50_2595 ();
 sg13g2_decap_8 FILLER_50_2602 ();
 sg13g2_decap_8 FILLER_50_2609 ();
 sg13g2_decap_8 FILLER_50_2616 ();
 sg13g2_decap_8 FILLER_50_2623 ();
 sg13g2_decap_8 FILLER_50_2630 ();
 sg13g2_decap_8 FILLER_50_2637 ();
 sg13g2_decap_8 FILLER_50_2644 ();
 sg13g2_decap_8 FILLER_50_2651 ();
 sg13g2_decap_8 FILLER_50_2658 ();
 sg13g2_decap_8 FILLER_50_2665 ();
 sg13g2_fill_2 FILLER_50_2672 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_8 FILLER_51_119 ();
 sg13g2_decap_8 FILLER_51_126 ();
 sg13g2_decap_8 FILLER_51_133 ();
 sg13g2_decap_8 FILLER_51_140 ();
 sg13g2_decap_8 FILLER_51_147 ();
 sg13g2_decap_4 FILLER_51_154 ();
 sg13g2_fill_1 FILLER_51_158 ();
 sg13g2_fill_1 FILLER_51_227 ();
 sg13g2_fill_1 FILLER_51_258 ();
 sg13g2_fill_2 FILLER_51_268 ();
 sg13g2_fill_1 FILLER_51_270 ();
 sg13g2_fill_2 FILLER_51_280 ();
 sg13g2_fill_1 FILLER_51_282 ();
 sg13g2_fill_2 FILLER_51_299 ();
 sg13g2_fill_1 FILLER_51_301 ();
 sg13g2_fill_1 FILLER_51_310 ();
 sg13g2_fill_2 FILLER_51_337 ();
 sg13g2_fill_1 FILLER_51_339 ();
 sg13g2_fill_1 FILLER_51_379 ();
 sg13g2_fill_1 FILLER_51_443 ();
 sg13g2_decap_4 FILLER_51_460 ();
 sg13g2_fill_1 FILLER_51_464 ();
 sg13g2_decap_4 FILLER_51_470 ();
 sg13g2_fill_2 FILLER_51_489 ();
 sg13g2_fill_1 FILLER_51_491 ();
 sg13g2_decap_8 FILLER_51_500 ();
 sg13g2_decap_4 FILLER_51_507 ();
 sg13g2_fill_2 FILLER_51_541 ();
 sg13g2_fill_1 FILLER_51_543 ();
 sg13g2_fill_1 FILLER_51_553 ();
 sg13g2_fill_2 FILLER_51_563 ();
 sg13g2_fill_1 FILLER_51_565 ();
 sg13g2_fill_2 FILLER_51_594 ();
 sg13g2_fill_1 FILLER_51_596 ();
 sg13g2_fill_2 FILLER_51_610 ();
 sg13g2_fill_1 FILLER_51_612 ();
 sg13g2_fill_2 FILLER_51_631 ();
 sg13g2_fill_1 FILLER_51_648 ();
 sg13g2_decap_4 FILLER_51_654 ();
 sg13g2_decap_4 FILLER_51_674 ();
 sg13g2_fill_2 FILLER_51_686 ();
 sg13g2_fill_1 FILLER_51_688 ();
 sg13g2_decap_4 FILLER_51_706 ();
 sg13g2_decap_8 FILLER_51_737 ();
 sg13g2_fill_2 FILLER_51_744 ();
 sg13g2_fill_1 FILLER_51_746 ();
 sg13g2_fill_1 FILLER_51_768 ();
 sg13g2_fill_2 FILLER_51_786 ();
 sg13g2_decap_4 FILLER_51_797 ();
 sg13g2_fill_1 FILLER_51_816 ();
 sg13g2_fill_1 FILLER_51_835 ();
 sg13g2_fill_2 FILLER_51_869 ();
 sg13g2_fill_2 FILLER_51_893 ();
 sg13g2_fill_1 FILLER_51_906 ();
 sg13g2_fill_2 FILLER_51_990 ();
 sg13g2_fill_1 FILLER_51_1018 ();
 sg13g2_fill_2 FILLER_51_1050 ();
 sg13g2_fill_2 FILLER_51_1095 ();
 sg13g2_fill_2 FILLER_51_1134 ();
 sg13g2_fill_2 FILLER_51_1178 ();
 sg13g2_fill_2 FILLER_51_1193 ();
 sg13g2_fill_2 FILLER_51_1295 ();
 sg13g2_fill_1 FILLER_51_1309 ();
 sg13g2_fill_2 FILLER_51_1332 ();
 sg13g2_fill_1 FILLER_51_1373 ();
 sg13g2_fill_2 FILLER_51_1432 ();
 sg13g2_fill_2 FILLER_51_1496 ();
 sg13g2_fill_1 FILLER_51_1516 ();
 sg13g2_fill_1 FILLER_51_1536 ();
 sg13g2_fill_2 FILLER_51_1631 ();
 sg13g2_fill_1 FILLER_51_1715 ();
 sg13g2_fill_2 FILLER_51_1742 ();
 sg13g2_fill_2 FILLER_51_1801 ();
 sg13g2_decap_8 FILLER_51_1829 ();
 sg13g2_decap_4 FILLER_51_1836 ();
 sg13g2_fill_2 FILLER_51_1890 ();
 sg13g2_fill_1 FILLER_51_1892 ();
 sg13g2_fill_2 FILLER_51_1927 ();
 sg13g2_decap_8 FILLER_51_1960 ();
 sg13g2_decap_8 FILLER_51_1967 ();
 sg13g2_fill_1 FILLER_51_1974 ();
 sg13g2_fill_1 FILLER_51_2024 ();
 sg13g2_fill_2 FILLER_51_2038 ();
 sg13g2_decap_4 FILLER_51_2057 ();
 sg13g2_decap_4 FILLER_51_2071 ();
 sg13g2_decap_8 FILLER_51_2088 ();
 sg13g2_fill_2 FILLER_51_2177 ();
 sg13g2_fill_1 FILLER_51_2179 ();
 sg13g2_fill_1 FILLER_51_2225 ();
 sg13g2_fill_1 FILLER_51_2235 ();
 sg13g2_fill_1 FILLER_51_2290 ();
 sg13g2_decap_8 FILLER_51_2295 ();
 sg13g2_decap_4 FILLER_51_2302 ();
 sg13g2_fill_1 FILLER_51_2306 ();
 sg13g2_decap_8 FILLER_51_2329 ();
 sg13g2_decap_8 FILLER_51_2336 ();
 sg13g2_decap_8 FILLER_51_2343 ();
 sg13g2_decap_8 FILLER_51_2350 ();
 sg13g2_decap_8 FILLER_51_2357 ();
 sg13g2_decap_8 FILLER_51_2364 ();
 sg13g2_decap_8 FILLER_51_2371 ();
 sg13g2_decap_8 FILLER_51_2378 ();
 sg13g2_decap_8 FILLER_51_2385 ();
 sg13g2_decap_8 FILLER_51_2392 ();
 sg13g2_decap_8 FILLER_51_2399 ();
 sg13g2_decap_8 FILLER_51_2406 ();
 sg13g2_decap_8 FILLER_51_2413 ();
 sg13g2_decap_8 FILLER_51_2420 ();
 sg13g2_decap_8 FILLER_51_2427 ();
 sg13g2_decap_8 FILLER_51_2434 ();
 sg13g2_decap_8 FILLER_51_2441 ();
 sg13g2_decap_8 FILLER_51_2448 ();
 sg13g2_decap_8 FILLER_51_2455 ();
 sg13g2_decap_8 FILLER_51_2462 ();
 sg13g2_decap_8 FILLER_51_2469 ();
 sg13g2_decap_8 FILLER_51_2476 ();
 sg13g2_decap_8 FILLER_51_2483 ();
 sg13g2_decap_8 FILLER_51_2490 ();
 sg13g2_decap_8 FILLER_51_2497 ();
 sg13g2_decap_8 FILLER_51_2504 ();
 sg13g2_decap_8 FILLER_51_2511 ();
 sg13g2_decap_8 FILLER_51_2518 ();
 sg13g2_decap_8 FILLER_51_2525 ();
 sg13g2_decap_8 FILLER_51_2532 ();
 sg13g2_decap_8 FILLER_51_2539 ();
 sg13g2_decap_8 FILLER_51_2546 ();
 sg13g2_decap_8 FILLER_51_2553 ();
 sg13g2_decap_8 FILLER_51_2560 ();
 sg13g2_decap_8 FILLER_51_2567 ();
 sg13g2_decap_8 FILLER_51_2574 ();
 sg13g2_decap_8 FILLER_51_2581 ();
 sg13g2_decap_8 FILLER_51_2588 ();
 sg13g2_decap_8 FILLER_51_2595 ();
 sg13g2_decap_8 FILLER_51_2602 ();
 sg13g2_decap_8 FILLER_51_2609 ();
 sg13g2_decap_8 FILLER_51_2616 ();
 sg13g2_decap_8 FILLER_51_2623 ();
 sg13g2_decap_8 FILLER_51_2630 ();
 sg13g2_decap_8 FILLER_51_2637 ();
 sg13g2_decap_8 FILLER_51_2644 ();
 sg13g2_decap_8 FILLER_51_2651 ();
 sg13g2_decap_8 FILLER_51_2658 ();
 sg13g2_decap_8 FILLER_51_2665 ();
 sg13g2_fill_2 FILLER_51_2672 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_119 ();
 sg13g2_decap_8 FILLER_52_126 ();
 sg13g2_decap_8 FILLER_52_133 ();
 sg13g2_decap_8 FILLER_52_140 ();
 sg13g2_decap_8 FILLER_52_147 ();
 sg13g2_decap_8 FILLER_52_154 ();
 sg13g2_decap_8 FILLER_52_161 ();
 sg13g2_decap_4 FILLER_52_168 ();
 sg13g2_fill_2 FILLER_52_224 ();
 sg13g2_fill_1 FILLER_52_226 ();
 sg13g2_fill_1 FILLER_52_236 ();
 sg13g2_decap_4 FILLER_52_276 ();
 sg13g2_fill_2 FILLER_52_280 ();
 sg13g2_fill_1 FILLER_52_286 ();
 sg13g2_fill_2 FILLER_52_292 ();
 sg13g2_fill_1 FILLER_52_294 ();
 sg13g2_fill_2 FILLER_52_306 ();
 sg13g2_fill_1 FILLER_52_308 ();
 sg13g2_fill_1 FILLER_52_318 ();
 sg13g2_fill_2 FILLER_52_345 ();
 sg13g2_fill_2 FILLER_52_363 ();
 sg13g2_fill_1 FILLER_52_397 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_fill_1 FILLER_52_426 ();
 sg13g2_fill_2 FILLER_52_440 ();
 sg13g2_fill_1 FILLER_52_442 ();
 sg13g2_fill_1 FILLER_52_460 ();
 sg13g2_fill_2 FILLER_52_492 ();
 sg13g2_fill_1 FILLER_52_504 ();
 sg13g2_fill_2 FILLER_52_558 ();
 sg13g2_fill_1 FILLER_52_560 ();
 sg13g2_fill_2 FILLER_52_571 ();
 sg13g2_decap_4 FILLER_52_656 ();
 sg13g2_fill_2 FILLER_52_678 ();
 sg13g2_fill_1 FILLER_52_680 ();
 sg13g2_fill_1 FILLER_52_686 ();
 sg13g2_fill_1 FILLER_52_699 ();
 sg13g2_decap_4 FILLER_52_759 ();
 sg13g2_fill_1 FILLER_52_763 ();
 sg13g2_decap_4 FILLER_52_805 ();
 sg13g2_fill_2 FILLER_52_812 ();
 sg13g2_decap_8 FILLER_52_819 ();
 sg13g2_fill_1 FILLER_52_826 ();
 sg13g2_decap_4 FILLER_52_845 ();
 sg13g2_fill_1 FILLER_52_849 ();
 sg13g2_decap_4 FILLER_52_860 ();
 sg13g2_fill_2 FILLER_52_864 ();
 sg13g2_fill_2 FILLER_52_876 ();
 sg13g2_fill_1 FILLER_52_883 ();
 sg13g2_fill_2 FILLER_52_941 ();
 sg13g2_fill_2 FILLER_52_952 ();
 sg13g2_fill_1 FILLER_52_1022 ();
 sg13g2_fill_1 FILLER_52_1078 ();
 sg13g2_fill_2 FILLER_52_1136 ();
 sg13g2_fill_2 FILLER_52_1176 ();
 sg13g2_fill_1 FILLER_52_1226 ();
 sg13g2_fill_2 FILLER_52_1313 ();
 sg13g2_fill_2 FILLER_52_1393 ();
 sg13g2_fill_2 FILLER_52_1493 ();
 sg13g2_fill_1 FILLER_52_1582 ();
 sg13g2_decap_4 FILLER_52_1606 ();
 sg13g2_fill_1 FILLER_52_1636 ();
 sg13g2_fill_1 FILLER_52_1651 ();
 sg13g2_fill_1 FILLER_52_1705 ();
 sg13g2_fill_1 FILLER_52_1715 ();
 sg13g2_fill_2 FILLER_52_1729 ();
 sg13g2_decap_4 FILLER_52_1778 ();
 sg13g2_decap_8 FILLER_52_1850 ();
 sg13g2_decap_8 FILLER_52_1857 ();
 sg13g2_decap_8 FILLER_52_1864 ();
 sg13g2_decap_8 FILLER_52_1871 ();
 sg13g2_fill_1 FILLER_52_1878 ();
 sg13g2_decap_8 FILLER_52_1892 ();
 sg13g2_fill_1 FILLER_52_1899 ();
 sg13g2_decap_8 FILLER_52_1912 ();
 sg13g2_decap_8 FILLER_52_1919 ();
 sg13g2_decap_8 FILLER_52_1926 ();
 sg13g2_fill_2 FILLER_52_1933 ();
 sg13g2_fill_1 FILLER_52_1943 ();
 sg13g2_decap_8 FILLER_52_1948 ();
 sg13g2_fill_2 FILLER_52_1968 ();
 sg13g2_decap_8 FILLER_52_1987 ();
 sg13g2_decap_8 FILLER_52_1994 ();
 sg13g2_fill_2 FILLER_52_2013 ();
 sg13g2_decap_4 FILLER_52_2059 ();
 sg13g2_fill_2 FILLER_52_2063 ();
 sg13g2_decap_4 FILLER_52_2069 ();
 sg13g2_decap_8 FILLER_52_2115 ();
 sg13g2_decap_4 FILLER_52_2138 ();
 sg13g2_fill_1 FILLER_52_2142 ();
 sg13g2_decap_8 FILLER_52_2153 ();
 sg13g2_fill_1 FILLER_52_2160 ();
 sg13g2_fill_2 FILLER_52_2273 ();
 sg13g2_decap_8 FILLER_52_2279 ();
 sg13g2_decap_8 FILLER_52_2286 ();
 sg13g2_fill_1 FILLER_52_2303 ();
 sg13g2_decap_8 FILLER_52_2330 ();
 sg13g2_decap_8 FILLER_52_2337 ();
 sg13g2_decap_8 FILLER_52_2344 ();
 sg13g2_decap_8 FILLER_52_2351 ();
 sg13g2_decap_8 FILLER_52_2358 ();
 sg13g2_decap_8 FILLER_52_2365 ();
 sg13g2_decap_8 FILLER_52_2372 ();
 sg13g2_decap_8 FILLER_52_2379 ();
 sg13g2_decap_8 FILLER_52_2386 ();
 sg13g2_decap_8 FILLER_52_2393 ();
 sg13g2_decap_8 FILLER_52_2400 ();
 sg13g2_decap_8 FILLER_52_2407 ();
 sg13g2_decap_8 FILLER_52_2414 ();
 sg13g2_decap_8 FILLER_52_2421 ();
 sg13g2_decap_8 FILLER_52_2428 ();
 sg13g2_decap_8 FILLER_52_2435 ();
 sg13g2_decap_8 FILLER_52_2442 ();
 sg13g2_decap_8 FILLER_52_2449 ();
 sg13g2_decap_8 FILLER_52_2456 ();
 sg13g2_decap_8 FILLER_52_2463 ();
 sg13g2_decap_8 FILLER_52_2470 ();
 sg13g2_decap_8 FILLER_52_2477 ();
 sg13g2_decap_8 FILLER_52_2484 ();
 sg13g2_decap_8 FILLER_52_2491 ();
 sg13g2_decap_8 FILLER_52_2498 ();
 sg13g2_decap_8 FILLER_52_2505 ();
 sg13g2_decap_8 FILLER_52_2512 ();
 sg13g2_decap_8 FILLER_52_2519 ();
 sg13g2_decap_8 FILLER_52_2526 ();
 sg13g2_decap_8 FILLER_52_2533 ();
 sg13g2_decap_8 FILLER_52_2540 ();
 sg13g2_decap_8 FILLER_52_2547 ();
 sg13g2_decap_8 FILLER_52_2554 ();
 sg13g2_decap_8 FILLER_52_2561 ();
 sg13g2_decap_8 FILLER_52_2568 ();
 sg13g2_decap_8 FILLER_52_2575 ();
 sg13g2_decap_8 FILLER_52_2582 ();
 sg13g2_decap_8 FILLER_52_2589 ();
 sg13g2_decap_8 FILLER_52_2596 ();
 sg13g2_decap_8 FILLER_52_2603 ();
 sg13g2_decap_8 FILLER_52_2610 ();
 sg13g2_decap_8 FILLER_52_2617 ();
 sg13g2_decap_8 FILLER_52_2624 ();
 sg13g2_decap_8 FILLER_52_2631 ();
 sg13g2_decap_8 FILLER_52_2638 ();
 sg13g2_decap_8 FILLER_52_2645 ();
 sg13g2_decap_8 FILLER_52_2652 ();
 sg13g2_decap_8 FILLER_52_2659 ();
 sg13g2_decap_8 FILLER_52_2666 ();
 sg13g2_fill_1 FILLER_52_2673 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_decap_8 FILLER_53_133 ();
 sg13g2_decap_8 FILLER_53_140 ();
 sg13g2_decap_8 FILLER_53_147 ();
 sg13g2_decap_8 FILLER_53_154 ();
 sg13g2_fill_2 FILLER_53_161 ();
 sg13g2_fill_1 FILLER_53_163 ();
 sg13g2_fill_1 FILLER_53_223 ();
 sg13g2_fill_1 FILLER_53_257 ();
 sg13g2_fill_1 FILLER_53_298 ();
 sg13g2_fill_2 FILLER_53_334 ();
 sg13g2_fill_1 FILLER_53_336 ();
 sg13g2_fill_2 FILLER_53_348 ();
 sg13g2_fill_2 FILLER_53_357 ();
 sg13g2_fill_1 FILLER_53_382 ();
 sg13g2_fill_1 FILLER_53_394 ();
 sg13g2_fill_1 FILLER_53_413 ();
 sg13g2_fill_2 FILLER_53_448 ();
 sg13g2_fill_1 FILLER_53_450 ();
 sg13g2_fill_2 FILLER_53_456 ();
 sg13g2_fill_1 FILLER_53_458 ();
 sg13g2_decap_8 FILLER_53_468 ();
 sg13g2_fill_2 FILLER_53_475 ();
 sg13g2_fill_2 FILLER_53_501 ();
 sg13g2_fill_1 FILLER_53_503 ();
 sg13g2_fill_1 FILLER_53_550 ();
 sg13g2_fill_2 FILLER_53_579 ();
 sg13g2_fill_1 FILLER_53_581 ();
 sg13g2_decap_4 FILLER_53_651 ();
 sg13g2_fill_1 FILLER_53_676 ();
 sg13g2_fill_2 FILLER_53_693 ();
 sg13g2_fill_2 FILLER_53_715 ();
 sg13g2_fill_1 FILLER_53_717 ();
 sg13g2_fill_2 FILLER_53_727 ();
 sg13g2_fill_2 FILLER_53_742 ();
 sg13g2_fill_1 FILLER_53_744 ();
 sg13g2_fill_1 FILLER_53_753 ();
 sg13g2_decap_4 FILLER_53_762 ();
 sg13g2_fill_1 FILLER_53_815 ();
 sg13g2_fill_1 FILLER_53_830 ();
 sg13g2_decap_8 FILLER_53_836 ();
 sg13g2_fill_2 FILLER_53_843 ();
 sg13g2_fill_1 FILLER_53_894 ();
 sg13g2_fill_2 FILLER_53_912 ();
 sg13g2_fill_1 FILLER_53_998 ();
 sg13g2_fill_1 FILLER_53_1023 ();
 sg13g2_fill_1 FILLER_53_1061 ();
 sg13g2_fill_1 FILLER_53_1116 ();
 sg13g2_fill_1 FILLER_53_1172 ();
 sg13g2_fill_1 FILLER_53_1192 ();
 sg13g2_fill_1 FILLER_53_1312 ();
 sg13g2_fill_2 FILLER_53_1440 ();
 sg13g2_fill_2 FILLER_53_1492 ();
 sg13g2_fill_2 FILLER_53_1523 ();
 sg13g2_fill_1 FILLER_53_1591 ();
 sg13g2_fill_2 FILLER_53_1633 ();
 sg13g2_fill_1 FILLER_53_1676 ();
 sg13g2_fill_2 FILLER_53_1796 ();
 sg13g2_fill_1 FILLER_53_1826 ();
 sg13g2_decap_8 FILLER_53_1831 ();
 sg13g2_decap_4 FILLER_53_1838 ();
 sg13g2_fill_1 FILLER_53_1842 ();
 sg13g2_fill_2 FILLER_53_1851 ();
 sg13g2_decap_8 FILLER_53_1879 ();
 sg13g2_decap_4 FILLER_53_1899 ();
 sg13g2_fill_1 FILLER_53_1914 ();
 sg13g2_fill_2 FILLER_53_1951 ();
 sg13g2_fill_1 FILLER_53_1953 ();
 sg13g2_fill_2 FILLER_53_1967 ();
 sg13g2_fill_1 FILLER_53_1969 ();
 sg13g2_decap_8 FILLER_53_1990 ();
 sg13g2_decap_8 FILLER_53_2010 ();
 sg13g2_decap_4 FILLER_53_2017 ();
 sg13g2_fill_1 FILLER_53_2021 ();
 sg13g2_fill_2 FILLER_53_2039 ();
 sg13g2_fill_1 FILLER_53_2053 ();
 sg13g2_decap_4 FILLER_53_2084 ();
 sg13g2_decap_8 FILLER_53_2106 ();
 sg13g2_fill_1 FILLER_53_2113 ();
 sg13g2_decap_4 FILLER_53_2128 ();
 sg13g2_fill_2 FILLER_53_2132 ();
 sg13g2_fill_2 FILLER_53_2169 ();
 sg13g2_decap_4 FILLER_53_2184 ();
 sg13g2_fill_1 FILLER_53_2188 ();
 sg13g2_fill_2 FILLER_53_2207 ();
 sg13g2_fill_1 FILLER_53_2227 ();
 sg13g2_fill_2 FILLER_53_2237 ();
 sg13g2_fill_2 FILLER_53_2265 ();
 sg13g2_fill_1 FILLER_53_2267 ();
 sg13g2_decap_4 FILLER_53_2299 ();
 sg13g2_fill_2 FILLER_53_2303 ();
 sg13g2_decap_8 FILLER_53_2331 ();
 sg13g2_decap_8 FILLER_53_2338 ();
 sg13g2_decap_8 FILLER_53_2345 ();
 sg13g2_decap_8 FILLER_53_2352 ();
 sg13g2_decap_8 FILLER_53_2359 ();
 sg13g2_decap_8 FILLER_53_2366 ();
 sg13g2_decap_8 FILLER_53_2373 ();
 sg13g2_decap_8 FILLER_53_2380 ();
 sg13g2_decap_8 FILLER_53_2387 ();
 sg13g2_decap_8 FILLER_53_2394 ();
 sg13g2_decap_8 FILLER_53_2401 ();
 sg13g2_decap_8 FILLER_53_2408 ();
 sg13g2_decap_8 FILLER_53_2415 ();
 sg13g2_decap_8 FILLER_53_2422 ();
 sg13g2_decap_8 FILLER_53_2429 ();
 sg13g2_decap_8 FILLER_53_2436 ();
 sg13g2_decap_8 FILLER_53_2443 ();
 sg13g2_decap_8 FILLER_53_2450 ();
 sg13g2_decap_8 FILLER_53_2457 ();
 sg13g2_decap_8 FILLER_53_2464 ();
 sg13g2_decap_8 FILLER_53_2471 ();
 sg13g2_decap_8 FILLER_53_2478 ();
 sg13g2_decap_8 FILLER_53_2485 ();
 sg13g2_decap_8 FILLER_53_2492 ();
 sg13g2_decap_8 FILLER_53_2499 ();
 sg13g2_decap_8 FILLER_53_2506 ();
 sg13g2_decap_8 FILLER_53_2513 ();
 sg13g2_decap_8 FILLER_53_2520 ();
 sg13g2_decap_8 FILLER_53_2527 ();
 sg13g2_decap_8 FILLER_53_2534 ();
 sg13g2_decap_8 FILLER_53_2541 ();
 sg13g2_decap_8 FILLER_53_2548 ();
 sg13g2_decap_8 FILLER_53_2555 ();
 sg13g2_decap_8 FILLER_53_2562 ();
 sg13g2_decap_8 FILLER_53_2569 ();
 sg13g2_decap_8 FILLER_53_2576 ();
 sg13g2_decap_8 FILLER_53_2583 ();
 sg13g2_decap_8 FILLER_53_2590 ();
 sg13g2_decap_8 FILLER_53_2597 ();
 sg13g2_decap_8 FILLER_53_2604 ();
 sg13g2_decap_8 FILLER_53_2611 ();
 sg13g2_decap_8 FILLER_53_2618 ();
 sg13g2_decap_8 FILLER_53_2625 ();
 sg13g2_decap_8 FILLER_53_2632 ();
 sg13g2_decap_8 FILLER_53_2639 ();
 sg13g2_decap_8 FILLER_53_2646 ();
 sg13g2_decap_8 FILLER_53_2653 ();
 sg13g2_decap_8 FILLER_53_2660 ();
 sg13g2_decap_8 FILLER_53_2667 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_decap_8 FILLER_54_119 ();
 sg13g2_decap_8 FILLER_54_126 ();
 sg13g2_decap_8 FILLER_54_133 ();
 sg13g2_decap_8 FILLER_54_140 ();
 sg13g2_decap_8 FILLER_54_147 ();
 sg13g2_decap_8 FILLER_54_154 ();
 sg13g2_decap_8 FILLER_54_161 ();
 sg13g2_decap_8 FILLER_54_168 ();
 sg13g2_fill_2 FILLER_54_175 ();
 sg13g2_fill_1 FILLER_54_177 ();
 sg13g2_fill_2 FILLER_54_191 ();
 sg13g2_fill_1 FILLER_54_193 ();
 sg13g2_fill_1 FILLER_54_210 ();
 sg13g2_decap_4 FILLER_54_224 ();
 sg13g2_fill_2 FILLER_54_228 ();
 sg13g2_fill_2 FILLER_54_238 ();
 sg13g2_fill_1 FILLER_54_240 ();
 sg13g2_fill_2 FILLER_54_250 ();
 sg13g2_fill_1 FILLER_54_252 ();
 sg13g2_decap_8 FILLER_54_257 ();
 sg13g2_decap_4 FILLER_54_264 ();
 sg13g2_decap_4 FILLER_54_273 ();
 sg13g2_fill_1 FILLER_54_277 ();
 sg13g2_fill_1 FILLER_54_292 ();
 sg13g2_fill_2 FILLER_54_310 ();
 sg13g2_fill_1 FILLER_54_312 ();
 sg13g2_fill_1 FILLER_54_318 ();
 sg13g2_fill_1 FILLER_54_335 ();
 sg13g2_fill_1 FILLER_54_350 ();
 sg13g2_fill_2 FILLER_54_387 ();
 sg13g2_fill_2 FILLER_54_423 ();
 sg13g2_fill_1 FILLER_54_429 ();
 sg13g2_decap_4 FILLER_54_455 ();
 sg13g2_fill_2 FILLER_54_466 ();
 sg13g2_fill_1 FILLER_54_472 ();
 sg13g2_fill_2 FILLER_54_487 ();
 sg13g2_fill_1 FILLER_54_625 ();
 sg13g2_decap_4 FILLER_54_644 ();
 sg13g2_fill_1 FILLER_54_648 ();
 sg13g2_decap_8 FILLER_54_671 ();
 sg13g2_fill_2 FILLER_54_678 ();
 sg13g2_fill_1 FILLER_54_696 ();
 sg13g2_fill_2 FILLER_54_707 ();
 sg13g2_fill_1 FILLER_54_735 ();
 sg13g2_fill_1 FILLER_54_752 ();
 sg13g2_decap_4 FILLER_54_766 ();
 sg13g2_decap_4 FILLER_54_774 ();
 sg13g2_fill_1 FILLER_54_778 ();
 sg13g2_decap_4 FILLER_54_785 ();
 sg13g2_fill_1 FILLER_54_789 ();
 sg13g2_fill_1 FILLER_54_796 ();
 sg13g2_fill_1 FILLER_54_804 ();
 sg13g2_fill_2 FILLER_54_816 ();
 sg13g2_fill_2 FILLER_54_823 ();
 sg13g2_fill_1 FILLER_54_825 ();
 sg13g2_fill_1 FILLER_54_837 ();
 sg13g2_decap_4 FILLER_54_856 ();
 sg13g2_fill_1 FILLER_54_860 ();
 sg13g2_fill_2 FILLER_54_875 ();
 sg13g2_fill_1 FILLER_54_992 ();
 sg13g2_fill_1 FILLER_54_998 ();
 sg13g2_fill_2 FILLER_54_1086 ();
 sg13g2_fill_2 FILLER_54_1134 ();
 sg13g2_fill_2 FILLER_54_1145 ();
 sg13g2_fill_2 FILLER_54_1156 ();
 sg13g2_fill_1 FILLER_54_1173 ();
 sg13g2_fill_1 FILLER_54_1313 ();
 sg13g2_fill_2 FILLER_54_1386 ();
 sg13g2_fill_1 FILLER_54_1449 ();
 sg13g2_fill_2 FILLER_54_1523 ();
 sg13g2_fill_1 FILLER_54_1599 ();
 sg13g2_decap_4 FILLER_54_1633 ();
 sg13g2_fill_2 FILLER_54_1723 ();
 sg13g2_fill_1 FILLER_54_1725 ();
 sg13g2_fill_2 FILLER_54_1736 ();
 sg13g2_fill_1 FILLER_54_1748 ();
 sg13g2_fill_1 FILLER_54_1785 ();
 sg13g2_fill_1 FILLER_54_1822 ();
 sg13g2_fill_2 FILLER_54_1861 ();
 sg13g2_fill_1 FILLER_54_1863 ();
 sg13g2_decap_8 FILLER_54_1868 ();
 sg13g2_fill_1 FILLER_54_1875 ();
 sg13g2_decap_8 FILLER_54_1884 ();
 sg13g2_fill_2 FILLER_54_1891 ();
 sg13g2_fill_2 FILLER_54_1901 ();
 sg13g2_fill_1 FILLER_54_1903 ();
 sg13g2_fill_1 FILLER_54_1933 ();
 sg13g2_decap_8 FILLER_54_1967 ();
 sg13g2_fill_2 FILLER_54_1974 ();
 sg13g2_fill_2 FILLER_54_1985 ();
 sg13g2_fill_1 FILLER_54_1987 ();
 sg13g2_decap_4 FILLER_54_2013 ();
 sg13g2_fill_1 FILLER_54_2017 ();
 sg13g2_fill_2 FILLER_54_2031 ();
 sg13g2_fill_1 FILLER_54_2033 ();
 sg13g2_fill_2 FILLER_54_2079 ();
 sg13g2_fill_2 FILLER_54_2187 ();
 sg13g2_fill_1 FILLER_54_2189 ();
 sg13g2_decap_8 FILLER_54_2226 ();
 sg13g2_fill_2 FILLER_54_2243 ();
 sg13g2_decap_4 FILLER_54_2276 ();
 sg13g2_fill_2 FILLER_54_2293 ();
 sg13g2_fill_1 FILLER_54_2295 ();
 sg13g2_decap_8 FILLER_54_2306 ();
 sg13g2_fill_2 FILLER_54_2313 ();
 sg13g2_decap_8 FILLER_54_2332 ();
 sg13g2_decap_8 FILLER_54_2339 ();
 sg13g2_decap_8 FILLER_54_2346 ();
 sg13g2_decap_8 FILLER_54_2353 ();
 sg13g2_decap_8 FILLER_54_2360 ();
 sg13g2_decap_8 FILLER_54_2367 ();
 sg13g2_decap_8 FILLER_54_2374 ();
 sg13g2_decap_8 FILLER_54_2381 ();
 sg13g2_decap_8 FILLER_54_2388 ();
 sg13g2_decap_8 FILLER_54_2395 ();
 sg13g2_decap_8 FILLER_54_2402 ();
 sg13g2_decap_8 FILLER_54_2409 ();
 sg13g2_decap_8 FILLER_54_2416 ();
 sg13g2_decap_8 FILLER_54_2423 ();
 sg13g2_decap_8 FILLER_54_2430 ();
 sg13g2_decap_8 FILLER_54_2437 ();
 sg13g2_decap_8 FILLER_54_2444 ();
 sg13g2_decap_8 FILLER_54_2451 ();
 sg13g2_decap_8 FILLER_54_2458 ();
 sg13g2_decap_8 FILLER_54_2465 ();
 sg13g2_decap_8 FILLER_54_2472 ();
 sg13g2_decap_8 FILLER_54_2479 ();
 sg13g2_decap_8 FILLER_54_2486 ();
 sg13g2_decap_8 FILLER_54_2493 ();
 sg13g2_decap_8 FILLER_54_2500 ();
 sg13g2_decap_8 FILLER_54_2507 ();
 sg13g2_decap_8 FILLER_54_2514 ();
 sg13g2_decap_8 FILLER_54_2521 ();
 sg13g2_decap_8 FILLER_54_2528 ();
 sg13g2_decap_8 FILLER_54_2535 ();
 sg13g2_decap_8 FILLER_54_2542 ();
 sg13g2_decap_8 FILLER_54_2549 ();
 sg13g2_decap_8 FILLER_54_2556 ();
 sg13g2_decap_8 FILLER_54_2563 ();
 sg13g2_decap_8 FILLER_54_2570 ();
 sg13g2_decap_8 FILLER_54_2577 ();
 sg13g2_decap_8 FILLER_54_2584 ();
 sg13g2_decap_8 FILLER_54_2591 ();
 sg13g2_decap_8 FILLER_54_2598 ();
 sg13g2_decap_8 FILLER_54_2605 ();
 sg13g2_decap_8 FILLER_54_2612 ();
 sg13g2_decap_8 FILLER_54_2619 ();
 sg13g2_decap_8 FILLER_54_2626 ();
 sg13g2_decap_8 FILLER_54_2633 ();
 sg13g2_decap_8 FILLER_54_2640 ();
 sg13g2_decap_8 FILLER_54_2647 ();
 sg13g2_decap_8 FILLER_54_2654 ();
 sg13g2_decap_8 FILLER_54_2661 ();
 sg13g2_decap_4 FILLER_54_2668 ();
 sg13g2_fill_2 FILLER_54_2672 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_decap_8 FILLER_55_126 ();
 sg13g2_decap_8 FILLER_55_133 ();
 sg13g2_decap_8 FILLER_55_140 ();
 sg13g2_decap_8 FILLER_55_147 ();
 sg13g2_decap_8 FILLER_55_154 ();
 sg13g2_decap_8 FILLER_55_161 ();
 sg13g2_fill_1 FILLER_55_168 ();
 sg13g2_fill_2 FILLER_55_214 ();
 sg13g2_fill_1 FILLER_55_221 ();
 sg13g2_decap_8 FILLER_55_239 ();
 sg13g2_fill_1 FILLER_55_246 ();
 sg13g2_fill_1 FILLER_55_260 ();
 sg13g2_fill_2 FILLER_55_269 ();
 sg13g2_fill_1 FILLER_55_271 ();
 sg13g2_decap_8 FILLER_55_288 ();
 sg13g2_decap_4 FILLER_55_295 ();
 sg13g2_fill_2 FILLER_55_299 ();
 sg13g2_fill_2 FILLER_55_318 ();
 sg13g2_fill_1 FILLER_55_320 ();
 sg13g2_fill_2 FILLER_55_334 ();
 sg13g2_fill_1 FILLER_55_336 ();
 sg13g2_fill_2 FILLER_55_342 ();
 sg13g2_fill_1 FILLER_55_344 ();
 sg13g2_fill_1 FILLER_55_375 ();
 sg13g2_decap_8 FILLER_55_380 ();
 sg13g2_fill_1 FILLER_55_387 ();
 sg13g2_fill_2 FILLER_55_414 ();
 sg13g2_fill_1 FILLER_55_416 ();
 sg13g2_fill_2 FILLER_55_455 ();
 sg13g2_decap_4 FILLER_55_488 ();
 sg13g2_fill_2 FILLER_55_492 ();
 sg13g2_fill_2 FILLER_55_507 ();
 sg13g2_fill_1 FILLER_55_509 ();
 sg13g2_fill_2 FILLER_55_579 ();
 sg13g2_fill_1 FILLER_55_652 ();
 sg13g2_fill_2 FILLER_55_658 ();
 sg13g2_fill_1 FILLER_55_660 ();
 sg13g2_fill_2 FILLER_55_669 ();
 sg13g2_fill_1 FILLER_55_671 ();
 sg13g2_fill_2 FILLER_55_677 ();
 sg13g2_decap_8 FILLER_55_693 ();
 sg13g2_decap_4 FILLER_55_700 ();
 sg13g2_fill_1 FILLER_55_704 ();
 sg13g2_decap_8 FILLER_55_709 ();
 sg13g2_fill_2 FILLER_55_716 ();
 sg13g2_decap_8 FILLER_55_739 ();
 sg13g2_fill_2 FILLER_55_746 ();
 sg13g2_fill_1 FILLER_55_748 ();
 sg13g2_decap_8 FILLER_55_757 ();
 sg13g2_decap_8 FILLER_55_764 ();
 sg13g2_fill_1 FILLER_55_771 ();
 sg13g2_fill_1 FILLER_55_790 ();
 sg13g2_fill_2 FILLER_55_802 ();
 sg13g2_fill_1 FILLER_55_814 ();
 sg13g2_fill_2 FILLER_55_820 ();
 sg13g2_fill_1 FILLER_55_822 ();
 sg13g2_fill_2 FILLER_55_828 ();
 sg13g2_decap_8 FILLER_55_834 ();
 sg13g2_fill_2 FILLER_55_851 ();
 sg13g2_fill_1 FILLER_55_853 ();
 sg13g2_fill_1 FILLER_55_874 ();
 sg13g2_fill_2 FILLER_55_880 ();
 sg13g2_fill_1 FILLER_55_882 ();
 sg13g2_fill_1 FILLER_55_957 ();
 sg13g2_fill_1 FILLER_55_1028 ();
 sg13g2_fill_1 FILLER_55_1047 ();
 sg13g2_fill_1 FILLER_55_1116 ();
 sg13g2_fill_2 FILLER_55_1252 ();
 sg13g2_fill_1 FILLER_55_1264 ();
 sg13g2_fill_2 FILLER_55_1274 ();
 sg13g2_fill_1 FILLER_55_1302 ();
 sg13g2_fill_1 FILLER_55_1410 ();
 sg13g2_fill_1 FILLER_55_1449 ();
 sg13g2_fill_1 FILLER_55_1520 ();
 sg13g2_fill_2 FILLER_55_1535 ();
 sg13g2_fill_1 FILLER_55_1537 ();
 sg13g2_decap_4 FILLER_55_1567 ();
 sg13g2_fill_1 FILLER_55_1571 ();
 sg13g2_fill_2 FILLER_55_1579 ();
 sg13g2_decap_4 FILLER_55_1590 ();
 sg13g2_fill_2 FILLER_55_1594 ();
 sg13g2_decap_4 FILLER_55_1626 ();
 sg13g2_fill_2 FILLER_55_1634 ();
 sg13g2_fill_1 FILLER_55_1636 ();
 sg13g2_fill_2 FILLER_55_1650 ();
 sg13g2_decap_4 FILLER_55_1709 ();
 sg13g2_fill_2 FILLER_55_1765 ();
 sg13g2_decap_4 FILLER_55_1875 ();
 sg13g2_fill_1 FILLER_55_1879 ();
 sg13g2_decap_4 FILLER_55_1893 ();
 sg13g2_fill_2 FILLER_55_1897 ();
 sg13g2_fill_2 FILLER_55_1912 ();
 sg13g2_fill_1 FILLER_55_1914 ();
 sg13g2_fill_2 FILLER_55_1921 ();
 sg13g2_fill_1 FILLER_55_1923 ();
 sg13g2_fill_1 FILLER_55_1932 ();
 sg13g2_fill_2 FILLER_55_1948 ();
 sg13g2_fill_2 FILLER_55_1990 ();
 sg13g2_fill_2 FILLER_55_2000 ();
 sg13g2_decap_8 FILLER_55_2028 ();
 sg13g2_fill_2 FILLER_55_2035 ();
 sg13g2_fill_2 FILLER_55_2047 ();
 sg13g2_fill_1 FILLER_55_2049 ();
 sg13g2_fill_1 FILLER_55_2091 ();
 sg13g2_fill_2 FILLER_55_2119 ();
 sg13g2_fill_2 FILLER_55_2126 ();
 sg13g2_fill_2 FILLER_55_2164 ();
 sg13g2_fill_1 FILLER_55_2166 ();
 sg13g2_decap_8 FILLER_55_2199 ();
 sg13g2_fill_1 FILLER_55_2250 ();
 sg13g2_fill_2 FILLER_55_2278 ();
 sg13g2_fill_1 FILLER_55_2280 ();
 sg13g2_fill_2 FILLER_55_2296 ();
 sg13g2_fill_1 FILLER_55_2308 ();
 sg13g2_decap_8 FILLER_55_2335 ();
 sg13g2_decap_8 FILLER_55_2342 ();
 sg13g2_decap_8 FILLER_55_2349 ();
 sg13g2_decap_8 FILLER_55_2356 ();
 sg13g2_decap_8 FILLER_55_2363 ();
 sg13g2_decap_8 FILLER_55_2370 ();
 sg13g2_decap_8 FILLER_55_2377 ();
 sg13g2_decap_8 FILLER_55_2384 ();
 sg13g2_decap_8 FILLER_55_2391 ();
 sg13g2_decap_8 FILLER_55_2398 ();
 sg13g2_decap_8 FILLER_55_2405 ();
 sg13g2_decap_8 FILLER_55_2412 ();
 sg13g2_decap_8 FILLER_55_2419 ();
 sg13g2_decap_8 FILLER_55_2426 ();
 sg13g2_decap_8 FILLER_55_2433 ();
 sg13g2_decap_8 FILLER_55_2440 ();
 sg13g2_decap_8 FILLER_55_2447 ();
 sg13g2_decap_8 FILLER_55_2454 ();
 sg13g2_decap_8 FILLER_55_2461 ();
 sg13g2_decap_8 FILLER_55_2468 ();
 sg13g2_decap_8 FILLER_55_2475 ();
 sg13g2_decap_8 FILLER_55_2482 ();
 sg13g2_decap_8 FILLER_55_2489 ();
 sg13g2_decap_8 FILLER_55_2496 ();
 sg13g2_decap_8 FILLER_55_2503 ();
 sg13g2_decap_8 FILLER_55_2510 ();
 sg13g2_decap_8 FILLER_55_2517 ();
 sg13g2_decap_8 FILLER_55_2524 ();
 sg13g2_decap_8 FILLER_55_2531 ();
 sg13g2_decap_8 FILLER_55_2538 ();
 sg13g2_decap_8 FILLER_55_2545 ();
 sg13g2_decap_8 FILLER_55_2552 ();
 sg13g2_decap_8 FILLER_55_2559 ();
 sg13g2_decap_8 FILLER_55_2566 ();
 sg13g2_decap_8 FILLER_55_2573 ();
 sg13g2_decap_8 FILLER_55_2580 ();
 sg13g2_decap_8 FILLER_55_2587 ();
 sg13g2_decap_8 FILLER_55_2594 ();
 sg13g2_decap_8 FILLER_55_2601 ();
 sg13g2_decap_8 FILLER_55_2608 ();
 sg13g2_decap_8 FILLER_55_2615 ();
 sg13g2_decap_8 FILLER_55_2622 ();
 sg13g2_decap_8 FILLER_55_2629 ();
 sg13g2_decap_8 FILLER_55_2636 ();
 sg13g2_decap_8 FILLER_55_2643 ();
 sg13g2_decap_8 FILLER_55_2650 ();
 sg13g2_decap_8 FILLER_55_2657 ();
 sg13g2_decap_8 FILLER_55_2664 ();
 sg13g2_fill_2 FILLER_55_2671 ();
 sg13g2_fill_1 FILLER_55_2673 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_decap_8 FILLER_56_119 ();
 sg13g2_decap_8 FILLER_56_126 ();
 sg13g2_decap_8 FILLER_56_133 ();
 sg13g2_decap_8 FILLER_56_140 ();
 sg13g2_decap_8 FILLER_56_147 ();
 sg13g2_decap_8 FILLER_56_154 ();
 sg13g2_decap_8 FILLER_56_161 ();
 sg13g2_decap_8 FILLER_56_168 ();
 sg13g2_decap_8 FILLER_56_175 ();
 sg13g2_fill_1 FILLER_56_204 ();
 sg13g2_fill_1 FILLER_56_210 ();
 sg13g2_decap_8 FILLER_56_251 ();
 sg13g2_fill_1 FILLER_56_258 ();
 sg13g2_fill_2 FILLER_56_271 ();
 sg13g2_fill_1 FILLER_56_316 ();
 sg13g2_fill_1 FILLER_56_366 ();
 sg13g2_fill_1 FILLER_56_380 ();
 sg13g2_fill_2 FILLER_56_386 ();
 sg13g2_fill_1 FILLER_56_388 ();
 sg13g2_fill_1 FILLER_56_401 ();
 sg13g2_fill_1 FILLER_56_415 ();
 sg13g2_fill_1 FILLER_56_425 ();
 sg13g2_fill_1 FILLER_56_439 ();
 sg13g2_decap_4 FILLER_56_475 ();
 sg13g2_fill_2 FILLER_56_479 ();
 sg13g2_fill_1 FILLER_56_489 ();
 sg13g2_fill_2 FILLER_56_560 ();
 sg13g2_fill_2 FILLER_56_579 ();
 sg13g2_fill_2 FILLER_56_598 ();
 sg13g2_fill_1 FILLER_56_600 ();
 sg13g2_fill_2 FILLER_56_634 ();
 sg13g2_fill_1 FILLER_56_636 ();
 sg13g2_fill_1 FILLER_56_689 ();
 sg13g2_decap_4 FILLER_56_703 ();
 sg13g2_decap_4 FILLER_56_764 ();
 sg13g2_decap_4 FILLER_56_783 ();
 sg13g2_fill_2 FILLER_56_787 ();
 sg13g2_decap_8 FILLER_56_794 ();
 sg13g2_decap_4 FILLER_56_801 ();
 sg13g2_fill_1 FILLER_56_805 ();
 sg13g2_fill_1 FILLER_56_828 ();
 sg13g2_fill_2 FILLER_56_841 ();
 sg13g2_fill_1 FILLER_56_843 ();
 sg13g2_decap_4 FILLER_56_855 ();
 sg13g2_fill_2 FILLER_56_859 ();
 sg13g2_fill_2 FILLER_56_872 ();
 sg13g2_fill_1 FILLER_56_874 ();
 sg13g2_fill_1 FILLER_56_891 ();
 sg13g2_fill_2 FILLER_56_898 ();
 sg13g2_fill_1 FILLER_56_1047 ();
 sg13g2_fill_1 FILLER_56_1098 ();
 sg13g2_fill_1 FILLER_56_1141 ();
 sg13g2_fill_1 FILLER_56_1159 ();
 sg13g2_fill_1 FILLER_56_1175 ();
 sg13g2_fill_1 FILLER_56_1266 ();
 sg13g2_fill_2 FILLER_56_1307 ();
 sg13g2_fill_2 FILLER_56_1357 ();
 sg13g2_fill_2 FILLER_56_1425 ();
 sg13g2_fill_1 FILLER_56_1560 ();
 sg13g2_fill_1 FILLER_56_1569 ();
 sg13g2_fill_1 FILLER_56_1583 ();
 sg13g2_fill_1 FILLER_56_1603 ();
 sg13g2_fill_1 FILLER_56_1645 ();
 sg13g2_fill_1 FILLER_56_1660 ();
 sg13g2_fill_2 FILLER_56_1704 ();
 sg13g2_fill_1 FILLER_56_1725 ();
 sg13g2_fill_2 FILLER_56_1740 ();
 sg13g2_fill_1 FILLER_56_1742 ();
 sg13g2_fill_2 FILLER_56_1752 ();
 sg13g2_fill_1 FILLER_56_1768 ();
 sg13g2_decap_8 FILLER_56_1788 ();
 sg13g2_decap_4 FILLER_56_1795 ();
 sg13g2_fill_1 FILLER_56_1799 ();
 sg13g2_fill_2 FILLER_56_1821 ();
 sg13g2_fill_2 FILLER_56_1858 ();
 sg13g2_decap_4 FILLER_56_1880 ();
 sg13g2_decap_4 FILLER_56_1913 ();
 sg13g2_decap_8 FILLER_56_1943 ();
 sg13g2_fill_2 FILLER_56_1950 ();
 sg13g2_fill_1 FILLER_56_1952 ();
 sg13g2_decap_8 FILLER_56_1965 ();
 sg13g2_fill_1 FILLER_56_1972 ();
 sg13g2_fill_1 FILLER_56_1987 ();
 sg13g2_decap_8 FILLER_56_2004 ();
 sg13g2_fill_2 FILLER_56_2011 ();
 sg13g2_decap_4 FILLER_56_2017 ();
 sg13g2_fill_2 FILLER_56_2082 ();
 sg13g2_fill_2 FILLER_56_2094 ();
 sg13g2_fill_1 FILLER_56_2096 ();
 sg13g2_fill_2 FILLER_56_2123 ();
 sg13g2_fill_1 FILLER_56_2131 ();
 sg13g2_fill_2 FILLER_56_2160 ();
 sg13g2_fill_2 FILLER_56_2206 ();
 sg13g2_fill_1 FILLER_56_2208 ();
 sg13g2_fill_2 FILLER_56_2217 ();
 sg13g2_fill_1 FILLER_56_2229 ();
 sg13g2_fill_1 FILLER_56_2247 ();
 sg13g2_fill_2 FILLER_56_2292 ();
 sg13g2_decap_8 FILLER_56_2328 ();
 sg13g2_decap_8 FILLER_56_2335 ();
 sg13g2_decap_8 FILLER_56_2342 ();
 sg13g2_decap_8 FILLER_56_2349 ();
 sg13g2_decap_8 FILLER_56_2356 ();
 sg13g2_decap_8 FILLER_56_2363 ();
 sg13g2_decap_8 FILLER_56_2370 ();
 sg13g2_decap_8 FILLER_56_2377 ();
 sg13g2_decap_8 FILLER_56_2384 ();
 sg13g2_decap_8 FILLER_56_2391 ();
 sg13g2_decap_8 FILLER_56_2398 ();
 sg13g2_decap_8 FILLER_56_2405 ();
 sg13g2_decap_8 FILLER_56_2412 ();
 sg13g2_decap_8 FILLER_56_2419 ();
 sg13g2_decap_8 FILLER_56_2426 ();
 sg13g2_decap_8 FILLER_56_2433 ();
 sg13g2_decap_8 FILLER_56_2440 ();
 sg13g2_decap_8 FILLER_56_2447 ();
 sg13g2_decap_8 FILLER_56_2454 ();
 sg13g2_decap_8 FILLER_56_2461 ();
 sg13g2_decap_8 FILLER_56_2468 ();
 sg13g2_decap_8 FILLER_56_2475 ();
 sg13g2_decap_8 FILLER_56_2482 ();
 sg13g2_decap_8 FILLER_56_2489 ();
 sg13g2_decap_8 FILLER_56_2496 ();
 sg13g2_decap_8 FILLER_56_2503 ();
 sg13g2_decap_8 FILLER_56_2510 ();
 sg13g2_decap_8 FILLER_56_2517 ();
 sg13g2_decap_8 FILLER_56_2524 ();
 sg13g2_decap_8 FILLER_56_2531 ();
 sg13g2_decap_8 FILLER_56_2538 ();
 sg13g2_decap_8 FILLER_56_2545 ();
 sg13g2_decap_8 FILLER_56_2552 ();
 sg13g2_decap_8 FILLER_56_2559 ();
 sg13g2_decap_8 FILLER_56_2566 ();
 sg13g2_decap_8 FILLER_56_2573 ();
 sg13g2_decap_8 FILLER_56_2580 ();
 sg13g2_decap_8 FILLER_56_2587 ();
 sg13g2_decap_8 FILLER_56_2594 ();
 sg13g2_decap_8 FILLER_56_2601 ();
 sg13g2_decap_8 FILLER_56_2608 ();
 sg13g2_decap_8 FILLER_56_2615 ();
 sg13g2_decap_8 FILLER_56_2622 ();
 sg13g2_decap_8 FILLER_56_2629 ();
 sg13g2_decap_8 FILLER_56_2636 ();
 sg13g2_decap_8 FILLER_56_2643 ();
 sg13g2_decap_8 FILLER_56_2650 ();
 sg13g2_decap_8 FILLER_56_2657 ();
 sg13g2_decap_8 FILLER_56_2664 ();
 sg13g2_fill_2 FILLER_56_2671 ();
 sg13g2_fill_1 FILLER_56_2673 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_decap_8 FILLER_57_126 ();
 sg13g2_decap_8 FILLER_57_133 ();
 sg13g2_decap_8 FILLER_57_140 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_decap_8 FILLER_57_154 ();
 sg13g2_decap_8 FILLER_57_161 ();
 sg13g2_decap_8 FILLER_57_168 ();
 sg13g2_fill_1 FILLER_57_175 ();
 sg13g2_fill_1 FILLER_57_266 ();
 sg13g2_decap_4 FILLER_57_272 ();
 sg13g2_decap_8 FILLER_57_311 ();
 sg13g2_decap_4 FILLER_57_327 ();
 sg13g2_fill_1 FILLER_57_331 ();
 sg13g2_fill_2 FILLER_57_340 ();
 sg13g2_fill_1 FILLER_57_389 ();
 sg13g2_fill_2 FILLER_57_563 ();
 sg13g2_fill_2 FILLER_57_579 ();
 sg13g2_fill_2 FILLER_57_591 ();
 sg13g2_fill_2 FILLER_57_620 ();
 sg13g2_fill_2 FILLER_57_659 ();
 sg13g2_fill_2 FILLER_57_682 ();
 sg13g2_fill_2 FILLER_57_689 ();
 sg13g2_fill_1 FILLER_57_702 ();
 sg13g2_decap_4 FILLER_57_745 ();
 sg13g2_fill_2 FILLER_57_749 ();
 sg13g2_fill_2 FILLER_57_768 ();
 sg13g2_fill_1 FILLER_57_770 ();
 sg13g2_fill_2 FILLER_57_785 ();
 sg13g2_fill_1 FILLER_57_787 ();
 sg13g2_fill_1 FILLER_57_798 ();
 sg13g2_fill_2 FILLER_57_809 ();
 sg13g2_fill_1 FILLER_57_816 ();
 sg13g2_fill_1 FILLER_57_826 ();
 sg13g2_decap_4 FILLER_57_831 ();
 sg13g2_fill_1 FILLER_57_835 ();
 sg13g2_decap_4 FILLER_57_850 ();
 sg13g2_fill_2 FILLER_57_854 ();
 sg13g2_fill_1 FILLER_57_861 ();
 sg13g2_fill_1 FILLER_57_874 ();
 sg13g2_fill_1 FILLER_57_944 ();
 sg13g2_fill_2 FILLER_57_1025 ();
 sg13g2_fill_1 FILLER_57_1058 ();
 sg13g2_fill_2 FILLER_57_1136 ();
 sg13g2_fill_1 FILLER_57_1197 ();
 sg13g2_fill_1 FILLER_57_1203 ();
 sg13g2_fill_2 FILLER_57_1239 ();
 sg13g2_fill_2 FILLER_57_1321 ();
 sg13g2_fill_1 FILLER_57_1323 ();
 sg13g2_fill_1 FILLER_57_1364 ();
 sg13g2_fill_1 FILLER_57_1452 ();
 sg13g2_fill_1 FILLER_57_1494 ();
 sg13g2_fill_1 FILLER_57_1528 ();
 sg13g2_fill_2 FILLER_57_1616 ();
 sg13g2_fill_1 FILLER_57_1618 ();
 sg13g2_fill_2 FILLER_57_1633 ();
 sg13g2_fill_1 FILLER_57_1635 ();
 sg13g2_fill_1 FILLER_57_1710 ();
 sg13g2_fill_2 FILLER_57_1745 ();
 sg13g2_fill_1 FILLER_57_1747 ();
 sg13g2_fill_1 FILLER_57_1758 ();
 sg13g2_fill_2 FILLER_57_1786 ();
 sg13g2_fill_2 FILLER_57_1793 ();
 sg13g2_fill_1 FILLER_57_1805 ();
 sg13g2_fill_2 FILLER_57_1827 ();
 sg13g2_fill_1 FILLER_57_1838 ();
 sg13g2_fill_2 FILLER_57_1849 ();
 sg13g2_decap_4 FILLER_57_1877 ();
 sg13g2_fill_2 FILLER_57_1881 ();
 sg13g2_decap_4 FILLER_57_1896 ();
 sg13g2_decap_8 FILLER_57_1922 ();
 sg13g2_decap_8 FILLER_57_1929 ();
 sg13g2_fill_2 FILLER_57_1936 ();
 sg13g2_fill_1 FILLER_57_1938 ();
 sg13g2_decap_4 FILLER_57_1965 ();
 sg13g2_fill_2 FILLER_57_1969 ();
 sg13g2_fill_2 FILLER_57_1984 ();
 sg13g2_fill_1 FILLER_57_1986 ();
 sg13g2_fill_2 FILLER_57_2000 ();
 sg13g2_decap_4 FILLER_57_2041 ();
 sg13g2_fill_1 FILLER_57_2045 ();
 sg13g2_decap_8 FILLER_57_2117 ();
 sg13g2_fill_2 FILLER_57_2129 ();
 sg13g2_fill_1 FILLER_57_2137 ();
 sg13g2_fill_2 FILLER_57_2164 ();
 sg13g2_fill_1 FILLER_57_2166 ();
 sg13g2_fill_2 FILLER_57_2197 ();
 sg13g2_fill_2 FILLER_57_2225 ();
 sg13g2_fill_2 FILLER_57_2253 ();
 sg13g2_fill_2 FILLER_57_2303 ();
 sg13g2_fill_1 FILLER_57_2305 ();
 sg13g2_decap_8 FILLER_57_2341 ();
 sg13g2_decap_8 FILLER_57_2348 ();
 sg13g2_decap_8 FILLER_57_2355 ();
 sg13g2_decap_8 FILLER_57_2362 ();
 sg13g2_decap_8 FILLER_57_2369 ();
 sg13g2_decap_8 FILLER_57_2376 ();
 sg13g2_decap_8 FILLER_57_2383 ();
 sg13g2_decap_8 FILLER_57_2390 ();
 sg13g2_decap_8 FILLER_57_2397 ();
 sg13g2_decap_8 FILLER_57_2404 ();
 sg13g2_decap_8 FILLER_57_2411 ();
 sg13g2_decap_8 FILLER_57_2418 ();
 sg13g2_decap_8 FILLER_57_2425 ();
 sg13g2_decap_8 FILLER_57_2432 ();
 sg13g2_decap_8 FILLER_57_2439 ();
 sg13g2_decap_8 FILLER_57_2446 ();
 sg13g2_decap_8 FILLER_57_2453 ();
 sg13g2_decap_8 FILLER_57_2460 ();
 sg13g2_decap_8 FILLER_57_2467 ();
 sg13g2_decap_8 FILLER_57_2474 ();
 sg13g2_decap_8 FILLER_57_2481 ();
 sg13g2_decap_8 FILLER_57_2488 ();
 sg13g2_decap_8 FILLER_57_2495 ();
 sg13g2_decap_8 FILLER_57_2502 ();
 sg13g2_decap_8 FILLER_57_2509 ();
 sg13g2_decap_8 FILLER_57_2516 ();
 sg13g2_decap_8 FILLER_57_2523 ();
 sg13g2_decap_8 FILLER_57_2530 ();
 sg13g2_decap_8 FILLER_57_2537 ();
 sg13g2_decap_8 FILLER_57_2544 ();
 sg13g2_decap_8 FILLER_57_2551 ();
 sg13g2_decap_8 FILLER_57_2558 ();
 sg13g2_decap_8 FILLER_57_2565 ();
 sg13g2_decap_8 FILLER_57_2572 ();
 sg13g2_decap_8 FILLER_57_2579 ();
 sg13g2_decap_8 FILLER_57_2586 ();
 sg13g2_decap_8 FILLER_57_2593 ();
 sg13g2_decap_8 FILLER_57_2600 ();
 sg13g2_decap_8 FILLER_57_2607 ();
 sg13g2_decap_8 FILLER_57_2614 ();
 sg13g2_decap_8 FILLER_57_2621 ();
 sg13g2_decap_8 FILLER_57_2628 ();
 sg13g2_decap_8 FILLER_57_2635 ();
 sg13g2_decap_8 FILLER_57_2642 ();
 sg13g2_decap_8 FILLER_57_2649 ();
 sg13g2_decap_8 FILLER_57_2656 ();
 sg13g2_decap_8 FILLER_57_2663 ();
 sg13g2_decap_4 FILLER_57_2670 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_8 FILLER_58_133 ();
 sg13g2_decap_8 FILLER_58_140 ();
 sg13g2_decap_8 FILLER_58_147 ();
 sg13g2_decap_8 FILLER_58_154 ();
 sg13g2_decap_8 FILLER_58_161 ();
 sg13g2_decap_8 FILLER_58_168 ();
 sg13g2_decap_8 FILLER_58_175 ();
 sg13g2_decap_4 FILLER_58_182 ();
 sg13g2_fill_1 FILLER_58_186 ();
 sg13g2_fill_2 FILLER_58_191 ();
 sg13g2_fill_1 FILLER_58_210 ();
 sg13g2_fill_2 FILLER_58_216 ();
 sg13g2_fill_1 FILLER_58_218 ();
 sg13g2_fill_2 FILLER_58_227 ();
 sg13g2_fill_2 FILLER_58_260 ();
 sg13g2_decap_4 FILLER_58_267 ();
 sg13g2_fill_2 FILLER_58_271 ();
 sg13g2_fill_2 FILLER_58_291 ();
 sg13g2_fill_1 FILLER_58_330 ();
 sg13g2_fill_2 FILLER_58_344 ();
 sg13g2_fill_1 FILLER_58_346 ();
 sg13g2_fill_2 FILLER_58_373 ();
 sg13g2_fill_1 FILLER_58_375 ();
 sg13g2_fill_2 FILLER_58_381 ();
 sg13g2_fill_1 FILLER_58_383 ();
 sg13g2_decap_8 FILLER_58_419 ();
 sg13g2_fill_1 FILLER_58_426 ();
 sg13g2_decap_4 FILLER_58_446 ();
 sg13g2_fill_2 FILLER_58_454 ();
 sg13g2_fill_1 FILLER_58_456 ();
 sg13g2_fill_2 FILLER_58_549 ();
 sg13g2_fill_1 FILLER_58_565 ();
 sg13g2_fill_1 FILLER_58_627 ();
 sg13g2_fill_1 FILLER_58_633 ();
 sg13g2_fill_2 FILLER_58_666 ();
 sg13g2_fill_1 FILLER_58_676 ();
 sg13g2_fill_2 FILLER_58_732 ();
 sg13g2_fill_2 FILLER_58_783 ();
 sg13g2_fill_1 FILLER_58_785 ();
 sg13g2_fill_2 FILLER_58_791 ();
 sg13g2_fill_1 FILLER_58_793 ();
 sg13g2_fill_2 FILLER_58_809 ();
 sg13g2_fill_1 FILLER_58_811 ();
 sg13g2_fill_2 FILLER_58_823 ();
 sg13g2_fill_1 FILLER_58_825 ();
 sg13g2_fill_2 FILLER_58_830 ();
 sg13g2_fill_1 FILLER_58_842 ();
 sg13g2_fill_2 FILLER_58_872 ();
 sg13g2_fill_1 FILLER_58_880 ();
 sg13g2_fill_2 FILLER_58_1064 ();
 sg13g2_fill_1 FILLER_58_1132 ();
 sg13g2_fill_2 FILLER_58_1224 ();
 sg13g2_fill_2 FILLER_58_1235 ();
 sg13g2_fill_2 FILLER_58_1283 ();
 sg13g2_fill_2 FILLER_58_1348 ();
 sg13g2_fill_2 FILLER_58_1364 ();
 sg13g2_fill_1 FILLER_58_1401 ();
 sg13g2_fill_2 FILLER_58_1419 ();
 sg13g2_fill_2 FILLER_58_1453 ();
 sg13g2_fill_2 FILLER_58_1498 ();
 sg13g2_fill_1 FILLER_58_1548 ();
 sg13g2_fill_2 FILLER_58_1584 ();
 sg13g2_fill_2 FILLER_58_1654 ();
 sg13g2_fill_2 FILLER_58_1666 ();
 sg13g2_fill_1 FILLER_58_1668 ();
 sg13g2_fill_2 FILLER_58_1699 ();
 sg13g2_fill_2 FILLER_58_1789 ();
 sg13g2_decap_8 FILLER_58_1867 ();
 sg13g2_fill_1 FILLER_58_1874 ();
 sg13g2_decap_8 FILLER_58_1883 ();
 sg13g2_fill_2 FILLER_58_1890 ();
 sg13g2_fill_1 FILLER_58_1892 ();
 sg13g2_fill_2 FILLER_58_1902 ();
 sg13g2_decap_8 FILLER_58_1935 ();
 sg13g2_decap_4 FILLER_58_1959 ();
 sg13g2_fill_1 FILLER_58_1963 ();
 sg13g2_fill_2 FILLER_58_1976 ();
 sg13g2_fill_1 FILLER_58_1978 ();
 sg13g2_fill_1 FILLER_58_1996 ();
 sg13g2_fill_1 FILLER_58_2001 ();
 sg13g2_fill_2 FILLER_58_2010 ();
 sg13g2_decap_8 FILLER_58_2016 ();
 sg13g2_decap_4 FILLER_58_2023 ();
 sg13g2_decap_4 FILLER_58_2036 ();
 sg13g2_fill_1 FILLER_58_2040 ();
 sg13g2_fill_2 FILLER_58_2097 ();
 sg13g2_fill_1 FILLER_58_2099 ();
 sg13g2_fill_1 FILLER_58_2105 ();
 sg13g2_fill_1 FILLER_58_2140 ();
 sg13g2_fill_2 FILLER_58_2176 ();
 sg13g2_fill_1 FILLER_58_2178 ();
 sg13g2_fill_2 FILLER_58_2209 ();
 sg13g2_fill_2 FILLER_58_2236 ();
 sg13g2_fill_1 FILLER_58_2265 ();
 sg13g2_fill_2 FILLER_58_2272 ();
 sg13g2_fill_1 FILLER_58_2274 ();
 sg13g2_fill_2 FILLER_58_2290 ();
 sg13g2_fill_2 FILLER_58_2302 ();
 sg13g2_fill_1 FILLER_58_2304 ();
 sg13g2_decap_4 FILLER_58_2320 ();
 sg13g2_fill_1 FILLER_58_2324 ();
 sg13g2_decap_8 FILLER_58_2338 ();
 sg13g2_decap_8 FILLER_58_2345 ();
 sg13g2_decap_8 FILLER_58_2352 ();
 sg13g2_decap_8 FILLER_58_2359 ();
 sg13g2_decap_8 FILLER_58_2366 ();
 sg13g2_decap_8 FILLER_58_2373 ();
 sg13g2_decap_8 FILLER_58_2380 ();
 sg13g2_decap_8 FILLER_58_2387 ();
 sg13g2_decap_8 FILLER_58_2394 ();
 sg13g2_decap_8 FILLER_58_2401 ();
 sg13g2_decap_8 FILLER_58_2408 ();
 sg13g2_decap_8 FILLER_58_2415 ();
 sg13g2_decap_8 FILLER_58_2422 ();
 sg13g2_decap_8 FILLER_58_2429 ();
 sg13g2_decap_8 FILLER_58_2436 ();
 sg13g2_decap_8 FILLER_58_2443 ();
 sg13g2_decap_8 FILLER_58_2450 ();
 sg13g2_decap_8 FILLER_58_2457 ();
 sg13g2_decap_8 FILLER_58_2464 ();
 sg13g2_decap_8 FILLER_58_2471 ();
 sg13g2_decap_8 FILLER_58_2478 ();
 sg13g2_decap_8 FILLER_58_2485 ();
 sg13g2_decap_8 FILLER_58_2492 ();
 sg13g2_decap_8 FILLER_58_2499 ();
 sg13g2_decap_8 FILLER_58_2506 ();
 sg13g2_decap_8 FILLER_58_2513 ();
 sg13g2_decap_8 FILLER_58_2520 ();
 sg13g2_decap_8 FILLER_58_2527 ();
 sg13g2_decap_8 FILLER_58_2534 ();
 sg13g2_decap_8 FILLER_58_2541 ();
 sg13g2_decap_8 FILLER_58_2548 ();
 sg13g2_decap_8 FILLER_58_2555 ();
 sg13g2_decap_8 FILLER_58_2562 ();
 sg13g2_decap_8 FILLER_58_2569 ();
 sg13g2_decap_8 FILLER_58_2576 ();
 sg13g2_decap_8 FILLER_58_2583 ();
 sg13g2_decap_8 FILLER_58_2590 ();
 sg13g2_decap_8 FILLER_58_2597 ();
 sg13g2_decap_8 FILLER_58_2604 ();
 sg13g2_decap_8 FILLER_58_2611 ();
 sg13g2_decap_8 FILLER_58_2618 ();
 sg13g2_decap_8 FILLER_58_2625 ();
 sg13g2_decap_8 FILLER_58_2632 ();
 sg13g2_decap_8 FILLER_58_2639 ();
 sg13g2_decap_8 FILLER_58_2646 ();
 sg13g2_decap_8 FILLER_58_2653 ();
 sg13g2_decap_8 FILLER_58_2660 ();
 sg13g2_decap_8 FILLER_58_2667 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_8 FILLER_59_126 ();
 sg13g2_decap_8 FILLER_59_133 ();
 sg13g2_decap_8 FILLER_59_140 ();
 sg13g2_decap_8 FILLER_59_147 ();
 sg13g2_decap_8 FILLER_59_154 ();
 sg13g2_decap_8 FILLER_59_161 ();
 sg13g2_decap_8 FILLER_59_168 ();
 sg13g2_decap_8 FILLER_59_175 ();
 sg13g2_decap_8 FILLER_59_182 ();
 sg13g2_decap_8 FILLER_59_189 ();
 sg13g2_decap_4 FILLER_59_196 ();
 sg13g2_fill_2 FILLER_59_200 ();
 sg13g2_fill_2 FILLER_59_230 ();
 sg13g2_decap_4 FILLER_59_242 ();
 sg13g2_fill_2 FILLER_59_246 ();
 sg13g2_fill_2 FILLER_59_262 ();
 sg13g2_decap_4 FILLER_59_278 ();
 sg13g2_fill_2 FILLER_59_305 ();
 sg13g2_fill_1 FILLER_59_329 ();
 sg13g2_fill_1 FILLER_59_363 ();
 sg13g2_decap_8 FILLER_59_403 ();
 sg13g2_decap_8 FILLER_59_410 ();
 sg13g2_decap_4 FILLER_59_417 ();
 sg13g2_fill_1 FILLER_59_421 ();
 sg13g2_fill_1 FILLER_59_438 ();
 sg13g2_fill_1 FILLER_59_516 ();
 sg13g2_fill_1 FILLER_59_526 ();
 sg13g2_fill_1 FILLER_59_546 ();
 sg13g2_fill_2 FILLER_59_595 ();
 sg13g2_fill_1 FILLER_59_597 ();
 sg13g2_fill_1 FILLER_59_603 ();
 sg13g2_fill_2 FILLER_59_617 ();
 sg13g2_fill_2 FILLER_59_697 ();
 sg13g2_decap_8 FILLER_59_733 ();
 sg13g2_decap_4 FILLER_59_740 ();
 sg13g2_fill_1 FILLER_59_744 ();
 sg13g2_decap_8 FILLER_59_749 ();
 sg13g2_fill_2 FILLER_59_756 ();
 sg13g2_fill_1 FILLER_59_762 ();
 sg13g2_fill_1 FILLER_59_794 ();
 sg13g2_fill_2 FILLER_59_808 ();
 sg13g2_fill_1 FILLER_59_810 ();
 sg13g2_fill_1 FILLER_59_827 ();
 sg13g2_fill_2 FILLER_59_838 ();
 sg13g2_fill_1 FILLER_59_867 ();
 sg13g2_fill_1 FILLER_59_884 ();
 sg13g2_fill_2 FILLER_59_890 ();
 sg13g2_fill_2 FILLER_59_971 ();
 sg13g2_fill_2 FILLER_59_999 ();
 sg13g2_fill_2 FILLER_59_1088 ();
 sg13g2_fill_1 FILLER_59_1114 ();
 sg13g2_fill_2 FILLER_59_1190 ();
 sg13g2_fill_1 FILLER_59_1206 ();
 sg13g2_fill_2 FILLER_59_1252 ();
 sg13g2_fill_1 FILLER_59_1387 ();
 sg13g2_fill_2 FILLER_59_1414 ();
 sg13g2_fill_1 FILLER_59_1439 ();
 sg13g2_fill_1 FILLER_59_1528 ();
 sg13g2_fill_1 FILLER_59_1567 ();
 sg13g2_fill_2 FILLER_59_1578 ();
 sg13g2_fill_2 FILLER_59_1592 ();
 sg13g2_fill_1 FILLER_59_1604 ();
 sg13g2_fill_2 FILLER_59_1666 ();
 sg13g2_fill_2 FILLER_59_1711 ();
 sg13g2_fill_1 FILLER_59_1713 ();
 sg13g2_fill_1 FILLER_59_1750 ();
 sg13g2_fill_2 FILLER_59_1770 ();
 sg13g2_fill_2 FILLER_59_1811 ();
 sg13g2_fill_1 FILLER_59_1813 ();
 sg13g2_fill_2 FILLER_59_1824 ();
 sg13g2_fill_1 FILLER_59_1826 ();
 sg13g2_fill_2 FILLER_59_1837 ();
 sg13g2_fill_1 FILLER_59_1861 ();
 sg13g2_decap_8 FILLER_59_1866 ();
 sg13g2_fill_2 FILLER_59_1873 ();
 sg13g2_decap_4 FILLER_59_1888 ();
 sg13g2_fill_1 FILLER_59_1892 ();
 sg13g2_fill_2 FILLER_59_1907 ();
 sg13g2_fill_2 FILLER_59_1913 ();
 sg13g2_fill_1 FILLER_59_1915 ();
 sg13g2_fill_1 FILLER_59_1922 ();
 sg13g2_fill_2 FILLER_59_1936 ();
 sg13g2_fill_1 FILLER_59_1964 ();
 sg13g2_fill_2 FILLER_59_1973 ();
 sg13g2_fill_1 FILLER_59_1975 ();
 sg13g2_fill_2 FILLER_59_1989 ();
 sg13g2_fill_1 FILLER_59_1991 ();
 sg13g2_decap_8 FILLER_59_2052 ();
 sg13g2_fill_2 FILLER_59_2059 ();
 sg13g2_fill_1 FILLER_59_2061 ();
 sg13g2_fill_2 FILLER_59_2098 ();
 sg13g2_fill_1 FILLER_59_2100 ();
 sg13g2_fill_2 FILLER_59_2113 ();
 sg13g2_fill_1 FILLER_59_2115 ();
 sg13g2_fill_1 FILLER_59_2121 ();
 sg13g2_fill_1 FILLER_59_2144 ();
 sg13g2_fill_1 FILLER_59_2220 ();
 sg13g2_fill_2 FILLER_59_2267 ();
 sg13g2_fill_1 FILLER_59_2269 ();
 sg13g2_decap_8 FILLER_59_2352 ();
 sg13g2_decap_8 FILLER_59_2359 ();
 sg13g2_decap_8 FILLER_59_2366 ();
 sg13g2_decap_8 FILLER_59_2373 ();
 sg13g2_decap_8 FILLER_59_2380 ();
 sg13g2_decap_8 FILLER_59_2387 ();
 sg13g2_decap_8 FILLER_59_2394 ();
 sg13g2_decap_8 FILLER_59_2401 ();
 sg13g2_decap_8 FILLER_59_2408 ();
 sg13g2_decap_8 FILLER_59_2415 ();
 sg13g2_decap_8 FILLER_59_2422 ();
 sg13g2_decap_8 FILLER_59_2429 ();
 sg13g2_decap_8 FILLER_59_2436 ();
 sg13g2_decap_8 FILLER_59_2443 ();
 sg13g2_decap_8 FILLER_59_2450 ();
 sg13g2_decap_8 FILLER_59_2457 ();
 sg13g2_decap_8 FILLER_59_2464 ();
 sg13g2_decap_8 FILLER_59_2471 ();
 sg13g2_decap_8 FILLER_59_2478 ();
 sg13g2_decap_8 FILLER_59_2485 ();
 sg13g2_decap_8 FILLER_59_2492 ();
 sg13g2_decap_8 FILLER_59_2499 ();
 sg13g2_decap_8 FILLER_59_2506 ();
 sg13g2_decap_8 FILLER_59_2513 ();
 sg13g2_decap_8 FILLER_59_2520 ();
 sg13g2_decap_8 FILLER_59_2527 ();
 sg13g2_decap_8 FILLER_59_2534 ();
 sg13g2_decap_8 FILLER_59_2541 ();
 sg13g2_decap_8 FILLER_59_2548 ();
 sg13g2_decap_8 FILLER_59_2555 ();
 sg13g2_decap_8 FILLER_59_2562 ();
 sg13g2_decap_8 FILLER_59_2569 ();
 sg13g2_decap_8 FILLER_59_2576 ();
 sg13g2_decap_8 FILLER_59_2583 ();
 sg13g2_decap_8 FILLER_59_2590 ();
 sg13g2_decap_8 FILLER_59_2597 ();
 sg13g2_decap_8 FILLER_59_2604 ();
 sg13g2_decap_8 FILLER_59_2611 ();
 sg13g2_decap_8 FILLER_59_2618 ();
 sg13g2_decap_8 FILLER_59_2625 ();
 sg13g2_decap_8 FILLER_59_2632 ();
 sg13g2_decap_8 FILLER_59_2639 ();
 sg13g2_decap_8 FILLER_59_2646 ();
 sg13g2_decap_8 FILLER_59_2653 ();
 sg13g2_decap_8 FILLER_59_2660 ();
 sg13g2_decap_8 FILLER_59_2667 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_112 ();
 sg13g2_decap_8 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_126 ();
 sg13g2_decap_8 FILLER_60_133 ();
 sg13g2_decap_8 FILLER_60_140 ();
 sg13g2_decap_8 FILLER_60_147 ();
 sg13g2_decap_8 FILLER_60_154 ();
 sg13g2_decap_8 FILLER_60_161 ();
 sg13g2_decap_8 FILLER_60_168 ();
 sg13g2_decap_8 FILLER_60_175 ();
 sg13g2_decap_8 FILLER_60_182 ();
 sg13g2_decap_8 FILLER_60_189 ();
 sg13g2_decap_8 FILLER_60_196 ();
 sg13g2_decap_4 FILLER_60_203 ();
 sg13g2_fill_2 FILLER_60_207 ();
 sg13g2_fill_2 FILLER_60_235 ();
 sg13g2_fill_2 FILLER_60_241 ();
 sg13g2_fill_2 FILLER_60_269 ();
 sg13g2_fill_2 FILLER_60_332 ();
 sg13g2_fill_1 FILLER_60_334 ();
 sg13g2_decap_4 FILLER_60_370 ();
 sg13g2_fill_1 FILLER_60_374 ();
 sg13g2_decap_8 FILLER_60_379 ();
 sg13g2_decap_8 FILLER_60_386 ();
 sg13g2_decap_8 FILLER_60_393 ();
 sg13g2_decap_8 FILLER_60_400 ();
 sg13g2_decap_8 FILLER_60_407 ();
 sg13g2_decap_4 FILLER_60_414 ();
 sg13g2_fill_2 FILLER_60_418 ();
 sg13g2_fill_2 FILLER_60_440 ();
 sg13g2_fill_1 FILLER_60_468 ();
 sg13g2_fill_1 FILLER_60_535 ();
 sg13g2_fill_2 FILLER_60_545 ();
 sg13g2_fill_1 FILLER_60_561 ();
 sg13g2_fill_2 FILLER_60_578 ();
 sg13g2_fill_1 FILLER_60_580 ();
 sg13g2_fill_1 FILLER_60_589 ();
 sg13g2_fill_2 FILLER_60_595 ();
 sg13g2_fill_2 FILLER_60_628 ();
 sg13g2_fill_1 FILLER_60_634 ();
 sg13g2_fill_2 FILLER_60_639 ();
 sg13g2_decap_4 FILLER_60_667 ();
 sg13g2_fill_1 FILLER_60_671 ();
 sg13g2_fill_2 FILLER_60_680 ();
 sg13g2_fill_1 FILLER_60_682 ();
 sg13g2_fill_2 FILLER_60_756 ();
 sg13g2_fill_1 FILLER_60_758 ();
 sg13g2_fill_2 FILLER_60_775 ();
 sg13g2_fill_1 FILLER_60_777 ();
 sg13g2_fill_2 FILLER_60_789 ();
 sg13g2_fill_2 FILLER_60_804 ();
 sg13g2_fill_2 FILLER_60_811 ();
 sg13g2_fill_1 FILLER_60_822 ();
 sg13g2_fill_2 FILLER_60_843 ();
 sg13g2_fill_2 FILLER_60_940 ();
 sg13g2_fill_1 FILLER_60_1011 ();
 sg13g2_fill_2 FILLER_60_1095 ();
 sg13g2_fill_1 FILLER_60_1158 ();
 sg13g2_fill_1 FILLER_60_1168 ();
 sg13g2_fill_1 FILLER_60_1178 ();
 sg13g2_fill_1 FILLER_60_1252 ();
 sg13g2_fill_1 FILLER_60_1423 ();
 sg13g2_fill_1 FILLER_60_1439 ();
 sg13g2_fill_1 FILLER_60_1492 ();
 sg13g2_fill_2 FILLER_60_1498 ();
 sg13g2_fill_1 FILLER_60_1571 ();
 sg13g2_fill_2 FILLER_60_1623 ();
 sg13g2_fill_1 FILLER_60_1634 ();
 sg13g2_fill_1 FILLER_60_1700 ();
 sg13g2_fill_1 FILLER_60_1710 ();
 sg13g2_fill_1 FILLER_60_1721 ();
 sg13g2_fill_2 FILLER_60_1726 ();
 sg13g2_fill_1 FILLER_60_1728 ();
 sg13g2_fill_1 FILLER_60_1791 ();
 sg13g2_decap_4 FILLER_60_1799 ();
 sg13g2_fill_1 FILLER_60_1808 ();
 sg13g2_fill_2 FILLER_60_1821 ();
 sg13g2_fill_2 FILLER_60_1831 ();
 sg13g2_fill_1 FILLER_60_1833 ();
 sg13g2_decap_4 FILLER_60_1870 ();
 sg13g2_fill_2 FILLER_60_1893 ();
 sg13g2_fill_2 FILLER_60_1903 ();
 sg13g2_fill_1 FILLER_60_1905 ();
 sg13g2_fill_2 FILLER_60_1918 ();
 sg13g2_fill_1 FILLER_60_1920 ();
 sg13g2_decap_4 FILLER_60_1931 ();
 sg13g2_fill_2 FILLER_60_1935 ();
 sg13g2_decap_4 FILLER_60_1945 ();
 sg13g2_decap_8 FILLER_60_1953 ();
 sg13g2_fill_1 FILLER_60_1960 ();
 sg13g2_decap_4 FILLER_60_1969 ();
 sg13g2_fill_1 FILLER_60_1973 ();
 sg13g2_decap_8 FILLER_60_1983 ();
 sg13g2_decap_4 FILLER_60_1990 ();
 sg13g2_fill_1 FILLER_60_1994 ();
 sg13g2_fill_2 FILLER_60_2001 ();
 sg13g2_decap_8 FILLER_60_2007 ();
 sg13g2_fill_2 FILLER_60_2014 ();
 sg13g2_decap_8 FILLER_60_2029 ();
 sg13g2_decap_8 FILLER_60_2062 ();
 sg13g2_fill_2 FILLER_60_2069 ();
 sg13g2_fill_1 FILLER_60_2071 ();
 sg13g2_decap_8 FILLER_60_2076 ();
 sg13g2_fill_2 FILLER_60_2106 ();
 sg13g2_decap_4 FILLER_60_2173 ();
 sg13g2_fill_1 FILLER_60_2177 ();
 sg13g2_fill_1 FILLER_60_2191 ();
 sg13g2_decap_8 FILLER_60_2233 ();
 sg13g2_decap_8 FILLER_60_2240 ();
 sg13g2_decap_4 FILLER_60_2247 ();
 sg13g2_decap_8 FILLER_60_2319 ();
 sg13g2_decap_8 FILLER_60_2339 ();
 sg13g2_decap_8 FILLER_60_2346 ();
 sg13g2_decap_8 FILLER_60_2353 ();
 sg13g2_decap_8 FILLER_60_2360 ();
 sg13g2_decap_8 FILLER_60_2367 ();
 sg13g2_decap_8 FILLER_60_2374 ();
 sg13g2_decap_8 FILLER_60_2381 ();
 sg13g2_decap_8 FILLER_60_2388 ();
 sg13g2_decap_8 FILLER_60_2395 ();
 sg13g2_decap_8 FILLER_60_2402 ();
 sg13g2_decap_8 FILLER_60_2409 ();
 sg13g2_decap_8 FILLER_60_2416 ();
 sg13g2_decap_8 FILLER_60_2423 ();
 sg13g2_decap_8 FILLER_60_2430 ();
 sg13g2_decap_8 FILLER_60_2437 ();
 sg13g2_decap_8 FILLER_60_2444 ();
 sg13g2_decap_8 FILLER_60_2451 ();
 sg13g2_decap_8 FILLER_60_2458 ();
 sg13g2_decap_8 FILLER_60_2465 ();
 sg13g2_decap_8 FILLER_60_2472 ();
 sg13g2_decap_8 FILLER_60_2479 ();
 sg13g2_decap_8 FILLER_60_2486 ();
 sg13g2_decap_8 FILLER_60_2493 ();
 sg13g2_decap_8 FILLER_60_2500 ();
 sg13g2_decap_8 FILLER_60_2507 ();
 sg13g2_decap_8 FILLER_60_2514 ();
 sg13g2_decap_8 FILLER_60_2521 ();
 sg13g2_decap_8 FILLER_60_2528 ();
 sg13g2_decap_8 FILLER_60_2535 ();
 sg13g2_decap_8 FILLER_60_2542 ();
 sg13g2_decap_8 FILLER_60_2549 ();
 sg13g2_decap_8 FILLER_60_2556 ();
 sg13g2_decap_8 FILLER_60_2563 ();
 sg13g2_decap_8 FILLER_60_2570 ();
 sg13g2_decap_8 FILLER_60_2577 ();
 sg13g2_decap_8 FILLER_60_2584 ();
 sg13g2_decap_8 FILLER_60_2591 ();
 sg13g2_decap_8 FILLER_60_2598 ();
 sg13g2_decap_8 FILLER_60_2605 ();
 sg13g2_decap_8 FILLER_60_2612 ();
 sg13g2_decap_8 FILLER_60_2619 ();
 sg13g2_decap_8 FILLER_60_2626 ();
 sg13g2_decap_8 FILLER_60_2633 ();
 sg13g2_decap_8 FILLER_60_2640 ();
 sg13g2_decap_8 FILLER_60_2647 ();
 sg13g2_decap_8 FILLER_60_2654 ();
 sg13g2_decap_8 FILLER_60_2661 ();
 sg13g2_decap_4 FILLER_60_2668 ();
 sg13g2_fill_2 FILLER_60_2672 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_decap_8 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_126 ();
 sg13g2_decap_8 FILLER_61_133 ();
 sg13g2_decap_8 FILLER_61_140 ();
 sg13g2_decap_8 FILLER_61_147 ();
 sg13g2_decap_8 FILLER_61_154 ();
 sg13g2_decap_8 FILLER_61_161 ();
 sg13g2_decap_8 FILLER_61_168 ();
 sg13g2_decap_8 FILLER_61_175 ();
 sg13g2_decap_8 FILLER_61_182 ();
 sg13g2_decap_8 FILLER_61_189 ();
 sg13g2_decap_8 FILLER_61_196 ();
 sg13g2_decap_8 FILLER_61_203 ();
 sg13g2_decap_8 FILLER_61_210 ();
 sg13g2_fill_1 FILLER_61_217 ();
 sg13g2_decap_4 FILLER_61_252 ();
 sg13g2_fill_2 FILLER_61_286 ();
 sg13g2_fill_2 FILLER_61_349 ();
 sg13g2_decap_8 FILLER_61_364 ();
 sg13g2_decap_8 FILLER_61_371 ();
 sg13g2_decap_8 FILLER_61_378 ();
 sg13g2_decap_8 FILLER_61_385 ();
 sg13g2_decap_8 FILLER_61_392 ();
 sg13g2_decap_8 FILLER_61_399 ();
 sg13g2_decap_8 FILLER_61_406 ();
 sg13g2_decap_8 FILLER_61_413 ();
 sg13g2_fill_2 FILLER_61_420 ();
 sg13g2_decap_8 FILLER_61_438 ();
 sg13g2_decap_8 FILLER_61_445 ();
 sg13g2_fill_1 FILLER_61_452 ();
 sg13g2_fill_1 FILLER_61_457 ();
 sg13g2_fill_1 FILLER_61_505 ();
 sg13g2_fill_1 FILLER_61_579 ();
 sg13g2_fill_2 FILLER_61_623 ();
 sg13g2_fill_1 FILLER_61_631 ();
 sg13g2_decap_8 FILLER_61_641 ();
 sg13g2_decap_4 FILLER_61_648 ();
 sg13g2_decap_4 FILLER_61_656 ();
 sg13g2_fill_1 FILLER_61_660 ();
 sg13g2_fill_2 FILLER_61_723 ();
 sg13g2_decap_8 FILLER_61_730 ();
 sg13g2_decap_4 FILLER_61_737 ();
 sg13g2_decap_8 FILLER_61_745 ();
 sg13g2_decap_4 FILLER_61_752 ();
 sg13g2_fill_2 FILLER_61_766 ();
 sg13g2_fill_1 FILLER_61_768 ();
 sg13g2_fill_1 FILLER_61_780 ();
 sg13g2_decap_4 FILLER_61_794 ();
 sg13g2_decap_8 FILLER_61_816 ();
 sg13g2_fill_2 FILLER_61_837 ();
 sg13g2_fill_1 FILLER_61_839 ();
 sg13g2_decap_4 FILLER_61_853 ();
 sg13g2_fill_1 FILLER_61_868 ();
 sg13g2_fill_1 FILLER_61_892 ();
 sg13g2_fill_2 FILLER_61_908 ();
 sg13g2_fill_1 FILLER_61_916 ();
 sg13g2_fill_2 FILLER_61_927 ();
 sg13g2_fill_1 FILLER_61_985 ();
 sg13g2_fill_1 FILLER_61_1040 ();
 sg13g2_fill_1 FILLER_61_1060 ();
 sg13g2_fill_1 FILLER_61_1075 ();
 sg13g2_fill_1 FILLER_61_1241 ();
 sg13g2_fill_2 FILLER_61_1299 ();
 sg13g2_fill_2 FILLER_61_1304 ();
 sg13g2_fill_1 FILLER_61_1435 ();
 sg13g2_fill_2 FILLER_61_1472 ();
 sg13g2_fill_2 FILLER_61_1561 ();
 sg13g2_fill_2 FILLER_61_1567 ();
 sg13g2_fill_2 FILLER_61_1615 ();
 sg13g2_fill_1 FILLER_61_1675 ();
 sg13g2_fill_1 FILLER_61_1750 ();
 sg13g2_fill_2 FILLER_61_1864 ();
 sg13g2_decap_4 FILLER_61_1879 ();
 sg13g2_decap_4 FILLER_61_1896 ();
 sg13g2_fill_1 FILLER_61_1926 ();
 sg13g2_decap_8 FILLER_61_1957 ();
 sg13g2_decap_8 FILLER_61_1978 ();
 sg13g2_fill_1 FILLER_61_1985 ();
 sg13g2_decap_4 FILLER_61_1990 ();
 sg13g2_fill_2 FILLER_61_1994 ();
 sg13g2_fill_2 FILLER_61_2022 ();
 sg13g2_fill_2 FILLER_61_2054 ();
 sg13g2_decap_8 FILLER_61_2082 ();
 sg13g2_fill_2 FILLER_61_2089 ();
 sg13g2_fill_2 FILLER_61_2134 ();
 sg13g2_decap_8 FILLER_61_2158 ();
 sg13g2_decap_8 FILLER_61_2165 ();
 sg13g2_decap_8 FILLER_61_2172 ();
 sg13g2_decap_4 FILLER_61_2179 ();
 sg13g2_fill_1 FILLER_61_2183 ();
 sg13g2_fill_1 FILLER_61_2197 ();
 sg13g2_fill_2 FILLER_61_2204 ();
 sg13g2_fill_1 FILLER_61_2211 ();
 sg13g2_fill_2 FILLER_61_2226 ();
 sg13g2_fill_2 FILLER_61_2236 ();
 sg13g2_decap_4 FILLER_61_2251 ();
 sg13g2_fill_1 FILLER_61_2255 ();
 sg13g2_decap_4 FILLER_61_2287 ();
 sg13g2_fill_2 FILLER_61_2300 ();
 sg13g2_fill_2 FILLER_61_2317 ();
 sg13g2_fill_1 FILLER_61_2319 ();
 sg13g2_decap_8 FILLER_61_2333 ();
 sg13g2_decap_8 FILLER_61_2340 ();
 sg13g2_decap_8 FILLER_61_2347 ();
 sg13g2_decap_8 FILLER_61_2354 ();
 sg13g2_decap_8 FILLER_61_2361 ();
 sg13g2_decap_8 FILLER_61_2368 ();
 sg13g2_decap_8 FILLER_61_2375 ();
 sg13g2_decap_8 FILLER_61_2382 ();
 sg13g2_decap_8 FILLER_61_2389 ();
 sg13g2_decap_8 FILLER_61_2396 ();
 sg13g2_decap_8 FILLER_61_2403 ();
 sg13g2_decap_8 FILLER_61_2410 ();
 sg13g2_decap_8 FILLER_61_2417 ();
 sg13g2_decap_8 FILLER_61_2424 ();
 sg13g2_decap_8 FILLER_61_2431 ();
 sg13g2_decap_8 FILLER_61_2438 ();
 sg13g2_decap_8 FILLER_61_2445 ();
 sg13g2_decap_8 FILLER_61_2452 ();
 sg13g2_decap_8 FILLER_61_2459 ();
 sg13g2_decap_8 FILLER_61_2466 ();
 sg13g2_decap_8 FILLER_61_2473 ();
 sg13g2_decap_8 FILLER_61_2480 ();
 sg13g2_decap_8 FILLER_61_2487 ();
 sg13g2_decap_8 FILLER_61_2494 ();
 sg13g2_decap_8 FILLER_61_2501 ();
 sg13g2_decap_8 FILLER_61_2508 ();
 sg13g2_decap_8 FILLER_61_2515 ();
 sg13g2_decap_8 FILLER_61_2522 ();
 sg13g2_decap_8 FILLER_61_2529 ();
 sg13g2_decap_8 FILLER_61_2536 ();
 sg13g2_decap_8 FILLER_61_2543 ();
 sg13g2_decap_8 FILLER_61_2550 ();
 sg13g2_decap_8 FILLER_61_2557 ();
 sg13g2_decap_8 FILLER_61_2564 ();
 sg13g2_decap_8 FILLER_61_2571 ();
 sg13g2_decap_8 FILLER_61_2578 ();
 sg13g2_decap_8 FILLER_61_2585 ();
 sg13g2_decap_8 FILLER_61_2592 ();
 sg13g2_decap_8 FILLER_61_2599 ();
 sg13g2_decap_8 FILLER_61_2606 ();
 sg13g2_decap_8 FILLER_61_2613 ();
 sg13g2_decap_8 FILLER_61_2620 ();
 sg13g2_decap_8 FILLER_61_2627 ();
 sg13g2_decap_8 FILLER_61_2634 ();
 sg13g2_decap_8 FILLER_61_2641 ();
 sg13g2_decap_8 FILLER_61_2648 ();
 sg13g2_decap_8 FILLER_61_2655 ();
 sg13g2_decap_8 FILLER_61_2662 ();
 sg13g2_decap_4 FILLER_61_2669 ();
 sg13g2_fill_1 FILLER_61_2673 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_decap_8 FILLER_62_126 ();
 sg13g2_decap_8 FILLER_62_133 ();
 sg13g2_decap_8 FILLER_62_140 ();
 sg13g2_decap_8 FILLER_62_147 ();
 sg13g2_decap_8 FILLER_62_154 ();
 sg13g2_decap_8 FILLER_62_161 ();
 sg13g2_decap_8 FILLER_62_168 ();
 sg13g2_decap_8 FILLER_62_175 ();
 sg13g2_decap_8 FILLER_62_182 ();
 sg13g2_decap_8 FILLER_62_189 ();
 sg13g2_decap_8 FILLER_62_196 ();
 sg13g2_decap_8 FILLER_62_203 ();
 sg13g2_decap_8 FILLER_62_210 ();
 sg13g2_decap_8 FILLER_62_217 ();
 sg13g2_decap_8 FILLER_62_224 ();
 sg13g2_decap_8 FILLER_62_231 ();
 sg13g2_decap_8 FILLER_62_238 ();
 sg13g2_decap_8 FILLER_62_245 ();
 sg13g2_decap_8 FILLER_62_252 ();
 sg13g2_decap_8 FILLER_62_259 ();
 sg13g2_decap_4 FILLER_62_266 ();
 sg13g2_decap_8 FILLER_62_283 ();
 sg13g2_decap_8 FILLER_62_290 ();
 sg13g2_decap_8 FILLER_62_297 ();
 sg13g2_decap_8 FILLER_62_308 ();
 sg13g2_decap_8 FILLER_62_315 ();
 sg13g2_decap_4 FILLER_62_322 ();
 sg13g2_fill_1 FILLER_62_326 ();
 sg13g2_fill_2 FILLER_62_336 ();
 sg13g2_decap_8 FILLER_62_343 ();
 sg13g2_decap_8 FILLER_62_350 ();
 sg13g2_decap_8 FILLER_62_357 ();
 sg13g2_decap_8 FILLER_62_364 ();
 sg13g2_decap_8 FILLER_62_371 ();
 sg13g2_decap_8 FILLER_62_378 ();
 sg13g2_decap_8 FILLER_62_385 ();
 sg13g2_decap_8 FILLER_62_392 ();
 sg13g2_decap_8 FILLER_62_399 ();
 sg13g2_decap_8 FILLER_62_406 ();
 sg13g2_decap_8 FILLER_62_413 ();
 sg13g2_decap_8 FILLER_62_420 ();
 sg13g2_decap_8 FILLER_62_427 ();
 sg13g2_fill_1 FILLER_62_434 ();
 sg13g2_fill_1 FILLER_62_474 ();
 sg13g2_fill_2 FILLER_62_485 ();
 sg13g2_fill_1 FILLER_62_487 ();
 sg13g2_fill_1 FILLER_62_493 ();
 sg13g2_fill_1 FILLER_62_499 ();
 sg13g2_fill_2 FILLER_62_510 ();
 sg13g2_fill_2 FILLER_62_526 ();
 sg13g2_fill_1 FILLER_62_533 ();
 sg13g2_fill_2 FILLER_62_544 ();
 sg13g2_fill_2 FILLER_62_560 ();
 sg13g2_fill_2 FILLER_62_579 ();
 sg13g2_fill_2 FILLER_62_595 ();
 sg13g2_decap_8 FILLER_62_663 ();
 sg13g2_fill_1 FILLER_62_670 ();
 sg13g2_fill_2 FILLER_62_714 ();
 sg13g2_fill_2 FILLER_62_742 ();
 sg13g2_fill_1 FILLER_62_744 ();
 sg13g2_fill_2 FILLER_62_753 ();
 sg13g2_fill_1 FILLER_62_755 ();
 sg13g2_fill_2 FILLER_62_771 ();
 sg13g2_fill_1 FILLER_62_791 ();
 sg13g2_fill_2 FILLER_62_803 ();
 sg13g2_fill_1 FILLER_62_805 ();
 sg13g2_fill_2 FILLER_62_810 ();
 sg13g2_fill_1 FILLER_62_812 ();
 sg13g2_decap_4 FILLER_62_826 ();
 sg13g2_decap_4 FILLER_62_835 ();
 sg13g2_fill_1 FILLER_62_839 ();
 sg13g2_fill_1 FILLER_62_849 ();
 sg13g2_fill_1 FILLER_62_865 ();
 sg13g2_fill_2 FILLER_62_881 ();
 sg13g2_fill_1 FILLER_62_891 ();
 sg13g2_fill_2 FILLER_62_948 ();
 sg13g2_fill_1 FILLER_62_1028 ();
 sg13g2_fill_1 FILLER_62_1309 ();
 sg13g2_fill_2 FILLER_62_1450 ();
 sg13g2_fill_2 FILLER_62_1549 ();
 sg13g2_fill_1 FILLER_62_1621 ();
 sg13g2_fill_2 FILLER_62_1641 ();
 sg13g2_fill_2 FILLER_62_1693 ();
 sg13g2_fill_1 FILLER_62_1695 ();
 sg13g2_fill_2 FILLER_62_1722 ();
 sg13g2_fill_1 FILLER_62_1789 ();
 sg13g2_fill_1 FILLER_62_1804 ();
 sg13g2_decap_4 FILLER_62_1820 ();
 sg13g2_fill_1 FILLER_62_1824 ();
 sg13g2_decap_4 FILLER_62_1870 ();
 sg13g2_fill_1 FILLER_62_1874 ();
 sg13g2_decap_8 FILLER_62_1880 ();
 sg13g2_decap_4 FILLER_62_1887 ();
 sg13g2_fill_2 FILLER_62_1891 ();
 sg13g2_fill_2 FILLER_62_1908 ();
 sg13g2_fill_1 FILLER_62_1910 ();
 sg13g2_fill_2 FILLER_62_1924 ();
 sg13g2_fill_1 FILLER_62_1926 ();
 sg13g2_fill_1 FILLER_62_1936 ();
 sg13g2_decap_8 FILLER_62_2024 ();
 sg13g2_decap_4 FILLER_62_2031 ();
 sg13g2_decap_8 FILLER_62_2039 ();
 sg13g2_decap_8 FILLER_62_2046 ();
 sg13g2_fill_2 FILLER_62_2053 ();
 sg13g2_fill_1 FILLER_62_2055 ();
 sg13g2_fill_1 FILLER_62_2060 ();
 sg13g2_fill_2 FILLER_62_2119 ();
 sg13g2_fill_2 FILLER_62_2126 ();
 sg13g2_decap_8 FILLER_62_2230 ();
 sg13g2_fill_1 FILLER_62_2237 ();
 sg13g2_decap_8 FILLER_62_2242 ();
 sg13g2_fill_2 FILLER_62_2249 ();
 sg13g2_fill_1 FILLER_62_2251 ();
 sg13g2_fill_2 FILLER_62_2262 ();
 sg13g2_fill_1 FILLER_62_2264 ();
 sg13g2_decap_8 FILLER_62_2343 ();
 sg13g2_decap_8 FILLER_62_2350 ();
 sg13g2_decap_8 FILLER_62_2357 ();
 sg13g2_decap_8 FILLER_62_2364 ();
 sg13g2_decap_8 FILLER_62_2371 ();
 sg13g2_decap_8 FILLER_62_2378 ();
 sg13g2_decap_8 FILLER_62_2385 ();
 sg13g2_decap_8 FILLER_62_2392 ();
 sg13g2_decap_8 FILLER_62_2399 ();
 sg13g2_decap_8 FILLER_62_2406 ();
 sg13g2_decap_8 FILLER_62_2413 ();
 sg13g2_decap_8 FILLER_62_2420 ();
 sg13g2_decap_8 FILLER_62_2427 ();
 sg13g2_decap_8 FILLER_62_2434 ();
 sg13g2_decap_8 FILLER_62_2441 ();
 sg13g2_decap_8 FILLER_62_2448 ();
 sg13g2_decap_8 FILLER_62_2455 ();
 sg13g2_decap_8 FILLER_62_2462 ();
 sg13g2_decap_8 FILLER_62_2469 ();
 sg13g2_decap_8 FILLER_62_2476 ();
 sg13g2_decap_8 FILLER_62_2483 ();
 sg13g2_decap_8 FILLER_62_2490 ();
 sg13g2_decap_8 FILLER_62_2497 ();
 sg13g2_decap_8 FILLER_62_2504 ();
 sg13g2_decap_8 FILLER_62_2511 ();
 sg13g2_decap_8 FILLER_62_2518 ();
 sg13g2_decap_8 FILLER_62_2525 ();
 sg13g2_decap_8 FILLER_62_2532 ();
 sg13g2_decap_8 FILLER_62_2539 ();
 sg13g2_decap_8 FILLER_62_2546 ();
 sg13g2_decap_8 FILLER_62_2553 ();
 sg13g2_decap_8 FILLER_62_2560 ();
 sg13g2_decap_8 FILLER_62_2567 ();
 sg13g2_decap_8 FILLER_62_2574 ();
 sg13g2_decap_8 FILLER_62_2581 ();
 sg13g2_decap_8 FILLER_62_2588 ();
 sg13g2_decap_8 FILLER_62_2595 ();
 sg13g2_decap_8 FILLER_62_2602 ();
 sg13g2_decap_8 FILLER_62_2609 ();
 sg13g2_decap_8 FILLER_62_2616 ();
 sg13g2_decap_8 FILLER_62_2623 ();
 sg13g2_decap_8 FILLER_62_2630 ();
 sg13g2_decap_8 FILLER_62_2637 ();
 sg13g2_decap_8 FILLER_62_2644 ();
 sg13g2_decap_8 FILLER_62_2651 ();
 sg13g2_decap_8 FILLER_62_2658 ();
 sg13g2_decap_8 FILLER_62_2665 ();
 sg13g2_fill_2 FILLER_62_2672 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_8 FILLER_63_126 ();
 sg13g2_decap_8 FILLER_63_133 ();
 sg13g2_decap_8 FILLER_63_140 ();
 sg13g2_decap_8 FILLER_63_147 ();
 sg13g2_decap_8 FILLER_63_154 ();
 sg13g2_decap_8 FILLER_63_161 ();
 sg13g2_decap_8 FILLER_63_168 ();
 sg13g2_decap_8 FILLER_63_175 ();
 sg13g2_decap_8 FILLER_63_182 ();
 sg13g2_decap_8 FILLER_63_189 ();
 sg13g2_decap_8 FILLER_63_196 ();
 sg13g2_decap_8 FILLER_63_203 ();
 sg13g2_decap_8 FILLER_63_210 ();
 sg13g2_decap_8 FILLER_63_217 ();
 sg13g2_decap_8 FILLER_63_224 ();
 sg13g2_decap_8 FILLER_63_231 ();
 sg13g2_decap_8 FILLER_63_238 ();
 sg13g2_decap_8 FILLER_63_245 ();
 sg13g2_decap_8 FILLER_63_252 ();
 sg13g2_decap_8 FILLER_63_259 ();
 sg13g2_decap_8 FILLER_63_266 ();
 sg13g2_decap_8 FILLER_63_273 ();
 sg13g2_decap_8 FILLER_63_280 ();
 sg13g2_decap_8 FILLER_63_287 ();
 sg13g2_decap_8 FILLER_63_294 ();
 sg13g2_decap_8 FILLER_63_301 ();
 sg13g2_decap_8 FILLER_63_308 ();
 sg13g2_decap_8 FILLER_63_315 ();
 sg13g2_decap_8 FILLER_63_322 ();
 sg13g2_decap_8 FILLER_63_329 ();
 sg13g2_decap_8 FILLER_63_336 ();
 sg13g2_decap_8 FILLER_63_343 ();
 sg13g2_decap_8 FILLER_63_350 ();
 sg13g2_decap_8 FILLER_63_357 ();
 sg13g2_decap_8 FILLER_63_364 ();
 sg13g2_decap_8 FILLER_63_371 ();
 sg13g2_decap_8 FILLER_63_378 ();
 sg13g2_decap_8 FILLER_63_385 ();
 sg13g2_decap_8 FILLER_63_392 ();
 sg13g2_decap_8 FILLER_63_399 ();
 sg13g2_decap_8 FILLER_63_406 ();
 sg13g2_decap_8 FILLER_63_413 ();
 sg13g2_decap_8 FILLER_63_420 ();
 sg13g2_decap_8 FILLER_63_427 ();
 sg13g2_decap_8 FILLER_63_434 ();
 sg13g2_decap_4 FILLER_63_441 ();
 sg13g2_fill_1 FILLER_63_497 ();
 sg13g2_fill_2 FILLER_63_534 ();
 sg13g2_fill_1 FILLER_63_566 ();
 sg13g2_fill_2 FILLER_63_629 ();
 sg13g2_fill_1 FILLER_63_631 ();
 sg13g2_fill_2 FILLER_63_645 ();
 sg13g2_fill_1 FILLER_63_647 ();
 sg13g2_fill_2 FILLER_63_678 ();
 sg13g2_fill_1 FILLER_63_680 ();
 sg13g2_decap_4 FILLER_63_685 ();
 sg13g2_fill_2 FILLER_63_715 ();
 sg13g2_fill_1 FILLER_63_717 ();
 sg13g2_decap_8 FILLER_63_748 ();
 sg13g2_fill_1 FILLER_63_755 ();
 sg13g2_fill_1 FILLER_63_769 ();
 sg13g2_decap_4 FILLER_63_775 ();
 sg13g2_fill_2 FILLER_63_789 ();
 sg13g2_fill_1 FILLER_63_791 ();
 sg13g2_fill_2 FILLER_63_798 ();
 sg13g2_fill_1 FILLER_63_800 ();
 sg13g2_fill_1 FILLER_63_806 ();
 sg13g2_fill_2 FILLER_63_819 ();
 sg13g2_fill_1 FILLER_63_852 ();
 sg13g2_fill_1 FILLER_63_914 ();
 sg13g2_fill_2 FILLER_63_949 ();
 sg13g2_fill_2 FILLER_63_1011 ();
 sg13g2_fill_2 FILLER_63_1078 ();
 sg13g2_fill_2 FILLER_63_1106 ();
 sg13g2_fill_2 FILLER_63_1131 ();
 sg13g2_fill_2 FILLER_63_1203 ();
 sg13g2_fill_1 FILLER_63_1300 ();
 sg13g2_fill_2 FILLER_63_1360 ();
 sg13g2_fill_2 FILLER_63_1419 ();
 sg13g2_fill_2 FILLER_63_1507 ();
 sg13g2_fill_2 FILLER_63_1622 ();
 sg13g2_fill_2 FILLER_63_1663 ();
 sg13g2_fill_2 FILLER_63_1719 ();
 sg13g2_fill_1 FILLER_63_1721 ();
 sg13g2_fill_2 FILLER_63_1765 ();
 sg13g2_fill_1 FILLER_63_1767 ();
 sg13g2_fill_1 FILLER_63_1860 ();
 sg13g2_fill_2 FILLER_63_1897 ();
 sg13g2_fill_2 FILLER_63_1961 ();
 sg13g2_fill_1 FILLER_63_1963 ();
 sg13g2_decap_8 FILLER_63_1973 ();
 sg13g2_decap_4 FILLER_63_1980 ();
 sg13g2_fill_2 FILLER_63_1984 ();
 sg13g2_decap_4 FILLER_63_2104 ();
 sg13g2_fill_2 FILLER_63_2114 ();
 sg13g2_fill_1 FILLER_63_2116 ();
 sg13g2_fill_2 FILLER_63_2137 ();
 sg13g2_fill_1 FILLER_63_2139 ();
 sg13g2_fill_2 FILLER_63_2144 ();
 sg13g2_fill_1 FILLER_63_2146 ();
 sg13g2_fill_1 FILLER_63_2183 ();
 sg13g2_fill_1 FILLER_63_2199 ();
 sg13g2_decap_8 FILLER_63_2209 ();
 sg13g2_fill_1 FILLER_63_2216 ();
 sg13g2_decap_4 FILLER_63_2253 ();
 sg13g2_fill_2 FILLER_63_2257 ();
 sg13g2_fill_2 FILLER_63_2264 ();
 sg13g2_fill_2 FILLER_63_2271 ();
 sg13g2_decap_4 FILLER_63_2290 ();
 sg13g2_fill_1 FILLER_63_2294 ();
 sg13g2_decap_8 FILLER_63_2312 ();
 sg13g2_decap_8 FILLER_63_2319 ();
 sg13g2_decap_8 FILLER_63_2326 ();
 sg13g2_decap_8 FILLER_63_2333 ();
 sg13g2_decap_8 FILLER_63_2340 ();
 sg13g2_decap_8 FILLER_63_2347 ();
 sg13g2_decap_8 FILLER_63_2354 ();
 sg13g2_decap_8 FILLER_63_2361 ();
 sg13g2_decap_8 FILLER_63_2368 ();
 sg13g2_decap_8 FILLER_63_2375 ();
 sg13g2_decap_8 FILLER_63_2382 ();
 sg13g2_decap_8 FILLER_63_2389 ();
 sg13g2_decap_8 FILLER_63_2396 ();
 sg13g2_decap_8 FILLER_63_2403 ();
 sg13g2_decap_8 FILLER_63_2410 ();
 sg13g2_decap_8 FILLER_63_2417 ();
 sg13g2_decap_8 FILLER_63_2424 ();
 sg13g2_decap_8 FILLER_63_2431 ();
 sg13g2_decap_8 FILLER_63_2438 ();
 sg13g2_decap_8 FILLER_63_2445 ();
 sg13g2_decap_8 FILLER_63_2452 ();
 sg13g2_decap_8 FILLER_63_2459 ();
 sg13g2_decap_8 FILLER_63_2466 ();
 sg13g2_decap_8 FILLER_63_2473 ();
 sg13g2_decap_8 FILLER_63_2480 ();
 sg13g2_decap_8 FILLER_63_2487 ();
 sg13g2_decap_8 FILLER_63_2494 ();
 sg13g2_decap_8 FILLER_63_2501 ();
 sg13g2_decap_8 FILLER_63_2508 ();
 sg13g2_decap_8 FILLER_63_2515 ();
 sg13g2_decap_8 FILLER_63_2522 ();
 sg13g2_decap_8 FILLER_63_2529 ();
 sg13g2_decap_8 FILLER_63_2536 ();
 sg13g2_decap_8 FILLER_63_2543 ();
 sg13g2_decap_8 FILLER_63_2550 ();
 sg13g2_decap_8 FILLER_63_2557 ();
 sg13g2_decap_8 FILLER_63_2564 ();
 sg13g2_decap_8 FILLER_63_2571 ();
 sg13g2_decap_8 FILLER_63_2578 ();
 sg13g2_decap_8 FILLER_63_2585 ();
 sg13g2_decap_8 FILLER_63_2592 ();
 sg13g2_decap_8 FILLER_63_2599 ();
 sg13g2_decap_8 FILLER_63_2606 ();
 sg13g2_decap_8 FILLER_63_2613 ();
 sg13g2_decap_8 FILLER_63_2620 ();
 sg13g2_decap_8 FILLER_63_2627 ();
 sg13g2_decap_8 FILLER_63_2634 ();
 sg13g2_decap_8 FILLER_63_2641 ();
 sg13g2_decap_8 FILLER_63_2648 ();
 sg13g2_decap_8 FILLER_63_2655 ();
 sg13g2_decap_8 FILLER_63_2662 ();
 sg13g2_decap_4 FILLER_63_2669 ();
 sg13g2_fill_1 FILLER_63_2673 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_147 ();
 sg13g2_decap_8 FILLER_64_154 ();
 sg13g2_decap_8 FILLER_64_161 ();
 sg13g2_decap_8 FILLER_64_168 ();
 sg13g2_decap_8 FILLER_64_175 ();
 sg13g2_decap_8 FILLER_64_182 ();
 sg13g2_decap_8 FILLER_64_189 ();
 sg13g2_decap_8 FILLER_64_196 ();
 sg13g2_decap_8 FILLER_64_203 ();
 sg13g2_decap_8 FILLER_64_210 ();
 sg13g2_decap_8 FILLER_64_217 ();
 sg13g2_decap_8 FILLER_64_224 ();
 sg13g2_decap_8 FILLER_64_231 ();
 sg13g2_decap_8 FILLER_64_238 ();
 sg13g2_decap_8 FILLER_64_245 ();
 sg13g2_decap_8 FILLER_64_252 ();
 sg13g2_decap_8 FILLER_64_259 ();
 sg13g2_decap_8 FILLER_64_266 ();
 sg13g2_decap_8 FILLER_64_273 ();
 sg13g2_decap_8 FILLER_64_280 ();
 sg13g2_decap_8 FILLER_64_287 ();
 sg13g2_decap_8 FILLER_64_294 ();
 sg13g2_decap_8 FILLER_64_301 ();
 sg13g2_decap_8 FILLER_64_308 ();
 sg13g2_decap_8 FILLER_64_315 ();
 sg13g2_decap_8 FILLER_64_322 ();
 sg13g2_decap_8 FILLER_64_329 ();
 sg13g2_decap_8 FILLER_64_336 ();
 sg13g2_decap_8 FILLER_64_343 ();
 sg13g2_decap_8 FILLER_64_350 ();
 sg13g2_fill_1 FILLER_64_357 ();
 sg13g2_decap_8 FILLER_64_369 ();
 sg13g2_decap_8 FILLER_64_376 ();
 sg13g2_decap_8 FILLER_64_383 ();
 sg13g2_decap_8 FILLER_64_390 ();
 sg13g2_decap_8 FILLER_64_397 ();
 sg13g2_decap_8 FILLER_64_404 ();
 sg13g2_decap_8 FILLER_64_411 ();
 sg13g2_decap_8 FILLER_64_418 ();
 sg13g2_decap_8 FILLER_64_425 ();
 sg13g2_fill_2 FILLER_64_432 ();
 sg13g2_fill_2 FILLER_64_470 ();
 sg13g2_fill_2 FILLER_64_532 ();
 sg13g2_fill_1 FILLER_64_619 ();
 sg13g2_fill_2 FILLER_64_630 ();
 sg13g2_fill_2 FILLER_64_672 ();
 sg13g2_decap_8 FILLER_64_687 ();
 sg13g2_fill_2 FILLER_64_694 ();
 sg13g2_fill_1 FILLER_64_696 ();
 sg13g2_fill_1 FILLER_64_705 ();
 sg13g2_decap_8 FILLER_64_712 ();
 sg13g2_decap_8 FILLER_64_719 ();
 sg13g2_decap_4 FILLER_64_726 ();
 sg13g2_fill_2 FILLER_64_730 ();
 sg13g2_fill_2 FILLER_64_758 ();
 sg13g2_fill_1 FILLER_64_765 ();
 sg13g2_fill_2 FILLER_64_779 ();
 sg13g2_fill_1 FILLER_64_781 ();
 sg13g2_fill_1 FILLER_64_798 ();
 sg13g2_decap_4 FILLER_64_804 ();
 sg13g2_fill_1 FILLER_64_808 ();
 sg13g2_decap_8 FILLER_64_823 ();
 sg13g2_decap_8 FILLER_64_834 ();
 sg13g2_decap_8 FILLER_64_841 ();
 sg13g2_fill_2 FILLER_64_863 ();
 sg13g2_fill_2 FILLER_64_879 ();
 sg13g2_fill_2 FILLER_64_986 ();
 sg13g2_fill_1 FILLER_64_1088 ();
 sg13g2_fill_1 FILLER_64_1191 ();
 sg13g2_fill_1 FILLER_64_1284 ();
 sg13g2_fill_1 FILLER_64_1309 ();
 sg13g2_fill_1 FILLER_64_1324 ();
 sg13g2_fill_1 FILLER_64_1417 ();
 sg13g2_fill_2 FILLER_64_1424 ();
 sg13g2_fill_1 FILLER_64_1532 ();
 sg13g2_fill_1 FILLER_64_1572 ();
 sg13g2_fill_2 FILLER_64_1714 ();
 sg13g2_fill_1 FILLER_64_1716 ();
 sg13g2_fill_2 FILLER_64_1783 ();
 sg13g2_fill_2 FILLER_64_1804 ();
 sg13g2_fill_1 FILLER_64_1806 ();
 sg13g2_fill_2 FILLER_64_1820 ();
 sg13g2_fill_1 FILLER_64_1822 ();
 sg13g2_decap_8 FILLER_64_1870 ();
 sg13g2_decap_4 FILLER_64_1877 ();
 sg13g2_fill_2 FILLER_64_1904 ();
 sg13g2_decap_4 FILLER_64_1990 ();
 sg13g2_fill_1 FILLER_64_2007 ();
 sg13g2_decap_8 FILLER_64_2044 ();
 sg13g2_fill_2 FILLER_64_2051 ();
 sg13g2_fill_2 FILLER_64_2072 ();
 sg13g2_decap_4 FILLER_64_2107 ();
 sg13g2_fill_1 FILLER_64_2116 ();
 sg13g2_fill_2 FILLER_64_2127 ();
 sg13g2_fill_2 FILLER_64_2160 ();
 sg13g2_fill_1 FILLER_64_2185 ();
 sg13g2_fill_2 FILLER_64_2279 ();
 sg13g2_fill_1 FILLER_64_2281 ();
 sg13g2_decap_8 FILLER_64_2323 ();
 sg13g2_decap_8 FILLER_64_2330 ();
 sg13g2_decap_8 FILLER_64_2337 ();
 sg13g2_decap_8 FILLER_64_2344 ();
 sg13g2_decap_8 FILLER_64_2351 ();
 sg13g2_decap_8 FILLER_64_2358 ();
 sg13g2_decap_8 FILLER_64_2365 ();
 sg13g2_decap_8 FILLER_64_2372 ();
 sg13g2_decap_8 FILLER_64_2379 ();
 sg13g2_decap_8 FILLER_64_2386 ();
 sg13g2_decap_8 FILLER_64_2393 ();
 sg13g2_decap_8 FILLER_64_2400 ();
 sg13g2_decap_8 FILLER_64_2407 ();
 sg13g2_decap_8 FILLER_64_2414 ();
 sg13g2_decap_8 FILLER_64_2421 ();
 sg13g2_decap_8 FILLER_64_2428 ();
 sg13g2_decap_8 FILLER_64_2435 ();
 sg13g2_decap_8 FILLER_64_2442 ();
 sg13g2_decap_8 FILLER_64_2449 ();
 sg13g2_decap_8 FILLER_64_2456 ();
 sg13g2_decap_8 FILLER_64_2463 ();
 sg13g2_decap_8 FILLER_64_2470 ();
 sg13g2_decap_8 FILLER_64_2477 ();
 sg13g2_decap_8 FILLER_64_2484 ();
 sg13g2_decap_8 FILLER_64_2491 ();
 sg13g2_decap_8 FILLER_64_2498 ();
 sg13g2_decap_8 FILLER_64_2505 ();
 sg13g2_decap_8 FILLER_64_2512 ();
 sg13g2_decap_8 FILLER_64_2519 ();
 sg13g2_decap_8 FILLER_64_2526 ();
 sg13g2_decap_8 FILLER_64_2533 ();
 sg13g2_decap_8 FILLER_64_2540 ();
 sg13g2_decap_8 FILLER_64_2547 ();
 sg13g2_decap_8 FILLER_64_2554 ();
 sg13g2_decap_8 FILLER_64_2561 ();
 sg13g2_decap_8 FILLER_64_2568 ();
 sg13g2_decap_8 FILLER_64_2575 ();
 sg13g2_decap_8 FILLER_64_2582 ();
 sg13g2_decap_8 FILLER_64_2589 ();
 sg13g2_decap_8 FILLER_64_2596 ();
 sg13g2_decap_8 FILLER_64_2603 ();
 sg13g2_decap_8 FILLER_64_2610 ();
 sg13g2_decap_8 FILLER_64_2617 ();
 sg13g2_decap_8 FILLER_64_2624 ();
 sg13g2_decap_8 FILLER_64_2631 ();
 sg13g2_decap_8 FILLER_64_2638 ();
 sg13g2_decap_8 FILLER_64_2645 ();
 sg13g2_decap_8 FILLER_64_2652 ();
 sg13g2_decap_8 FILLER_64_2659 ();
 sg13g2_decap_8 FILLER_64_2666 ();
 sg13g2_fill_1 FILLER_64_2673 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_decap_8 FILLER_65_140 ();
 sg13g2_decap_8 FILLER_65_147 ();
 sg13g2_decap_8 FILLER_65_154 ();
 sg13g2_decap_8 FILLER_65_161 ();
 sg13g2_decap_8 FILLER_65_168 ();
 sg13g2_decap_8 FILLER_65_175 ();
 sg13g2_decap_8 FILLER_65_182 ();
 sg13g2_decap_8 FILLER_65_189 ();
 sg13g2_decap_8 FILLER_65_196 ();
 sg13g2_decap_8 FILLER_65_203 ();
 sg13g2_decap_8 FILLER_65_210 ();
 sg13g2_decap_8 FILLER_65_217 ();
 sg13g2_decap_8 FILLER_65_224 ();
 sg13g2_decap_8 FILLER_65_231 ();
 sg13g2_decap_8 FILLER_65_238 ();
 sg13g2_decap_8 FILLER_65_245 ();
 sg13g2_decap_8 FILLER_65_252 ();
 sg13g2_decap_8 FILLER_65_259 ();
 sg13g2_decap_8 FILLER_65_266 ();
 sg13g2_decap_8 FILLER_65_273 ();
 sg13g2_decap_8 FILLER_65_280 ();
 sg13g2_decap_8 FILLER_65_287 ();
 sg13g2_decap_8 FILLER_65_294 ();
 sg13g2_decap_8 FILLER_65_301 ();
 sg13g2_decap_8 FILLER_65_308 ();
 sg13g2_decap_8 FILLER_65_315 ();
 sg13g2_decap_8 FILLER_65_322 ();
 sg13g2_decap_8 FILLER_65_329 ();
 sg13g2_decap_8 FILLER_65_336 ();
 sg13g2_decap_8 FILLER_65_343 ();
 sg13g2_decap_8 FILLER_65_350 ();
 sg13g2_decap_8 FILLER_65_357 ();
 sg13g2_decap_8 FILLER_65_364 ();
 sg13g2_decap_8 FILLER_65_371 ();
 sg13g2_decap_8 FILLER_65_378 ();
 sg13g2_decap_8 FILLER_65_385 ();
 sg13g2_decap_8 FILLER_65_392 ();
 sg13g2_decap_8 FILLER_65_399 ();
 sg13g2_decap_8 FILLER_65_406 ();
 sg13g2_decap_8 FILLER_65_413 ();
 sg13g2_decap_4 FILLER_65_420 ();
 sg13g2_fill_2 FILLER_65_463 ();
 sg13g2_fill_2 FILLER_65_489 ();
 sg13g2_fill_1 FILLER_65_491 ();
 sg13g2_fill_1 FILLER_65_501 ();
 sg13g2_fill_2 FILLER_65_512 ();
 sg13g2_fill_2 FILLER_65_545 ();
 sg13g2_fill_2 FILLER_65_552 ();
 sg13g2_fill_1 FILLER_65_554 ();
 sg13g2_fill_1 FILLER_65_584 ();
 sg13g2_fill_1 FILLER_65_591 ();
 sg13g2_fill_2 FILLER_65_613 ();
 sg13g2_fill_1 FILLER_65_615 ();
 sg13g2_fill_2 FILLER_65_632 ();
 sg13g2_fill_1 FILLER_65_634 ();
 sg13g2_fill_2 FILLER_65_656 ();
 sg13g2_fill_2 FILLER_65_666 ();
 sg13g2_fill_1 FILLER_65_668 ();
 sg13g2_decap_8 FILLER_65_700 ();
 sg13g2_decap_8 FILLER_65_707 ();
 sg13g2_decap_4 FILLER_65_714 ();
 sg13g2_fill_2 FILLER_65_718 ();
 sg13g2_decap_8 FILLER_65_725 ();
 sg13g2_decap_4 FILLER_65_732 ();
 sg13g2_fill_1 FILLER_65_736 ();
 sg13g2_fill_2 FILLER_65_763 ();
 sg13g2_fill_1 FILLER_65_765 ();
 sg13g2_decap_4 FILLER_65_772 ();
 sg13g2_fill_1 FILLER_65_796 ();
 sg13g2_fill_1 FILLER_65_819 ();
 sg13g2_fill_1 FILLER_65_838 ();
 sg13g2_fill_2 FILLER_65_873 ();
 sg13g2_fill_1 FILLER_65_899 ();
 sg13g2_fill_1 FILLER_65_1051 ();
 sg13g2_fill_1 FILLER_65_1066 ();
 sg13g2_fill_1 FILLER_65_1139 ();
 sg13g2_fill_2 FILLER_65_1174 ();
 sg13g2_fill_1 FILLER_65_1200 ();
 sg13g2_fill_1 FILLER_65_1215 ();
 sg13g2_fill_1 FILLER_65_1225 ();
 sg13g2_fill_1 FILLER_65_1266 ();
 sg13g2_fill_1 FILLER_65_1279 ();
 sg13g2_fill_2 FILLER_65_1290 ();
 sg13g2_fill_2 FILLER_65_1413 ();
 sg13g2_fill_2 FILLER_65_1647 ();
 sg13g2_fill_2 FILLER_65_1655 ();
 sg13g2_fill_2 FILLER_65_1675 ();
 sg13g2_fill_2 FILLER_65_1691 ();
 sg13g2_fill_2 FILLER_65_1738 ();
 sg13g2_fill_1 FILLER_65_1740 ();
 sg13g2_fill_1 FILLER_65_1813 ();
 sg13g2_fill_2 FILLER_65_1906 ();
 sg13g2_fill_1 FILLER_65_1908 ();
 sg13g2_fill_2 FILLER_65_1940 ();
 sg13g2_fill_1 FILLER_65_1950 ();
 sg13g2_fill_2 FILLER_65_1972 ();
 sg13g2_fill_1 FILLER_65_1974 ();
 sg13g2_fill_2 FILLER_65_2015 ();
 sg13g2_fill_2 FILLER_65_2118 ();
 sg13g2_fill_2 FILLER_65_2145 ();
 sg13g2_fill_2 FILLER_65_2191 ();
 sg13g2_fill_1 FILLER_65_2214 ();
 sg13g2_fill_2 FILLER_65_2225 ();
 sg13g2_fill_1 FILLER_65_2227 ();
 sg13g2_fill_1 FILLER_65_2291 ();
 sg13g2_fill_1 FILLER_65_2297 ();
 sg13g2_decap_8 FILLER_65_2311 ();
 sg13g2_decap_8 FILLER_65_2318 ();
 sg13g2_decap_8 FILLER_65_2325 ();
 sg13g2_decap_8 FILLER_65_2332 ();
 sg13g2_decap_8 FILLER_65_2339 ();
 sg13g2_decap_8 FILLER_65_2346 ();
 sg13g2_decap_8 FILLER_65_2353 ();
 sg13g2_decap_8 FILLER_65_2360 ();
 sg13g2_decap_8 FILLER_65_2367 ();
 sg13g2_decap_8 FILLER_65_2374 ();
 sg13g2_decap_8 FILLER_65_2381 ();
 sg13g2_decap_8 FILLER_65_2388 ();
 sg13g2_decap_8 FILLER_65_2395 ();
 sg13g2_decap_8 FILLER_65_2402 ();
 sg13g2_decap_8 FILLER_65_2409 ();
 sg13g2_decap_8 FILLER_65_2416 ();
 sg13g2_decap_8 FILLER_65_2423 ();
 sg13g2_decap_8 FILLER_65_2430 ();
 sg13g2_decap_8 FILLER_65_2437 ();
 sg13g2_decap_8 FILLER_65_2444 ();
 sg13g2_decap_8 FILLER_65_2451 ();
 sg13g2_decap_8 FILLER_65_2458 ();
 sg13g2_decap_8 FILLER_65_2465 ();
 sg13g2_decap_8 FILLER_65_2472 ();
 sg13g2_decap_8 FILLER_65_2479 ();
 sg13g2_decap_8 FILLER_65_2486 ();
 sg13g2_decap_8 FILLER_65_2493 ();
 sg13g2_decap_8 FILLER_65_2500 ();
 sg13g2_decap_8 FILLER_65_2507 ();
 sg13g2_decap_8 FILLER_65_2514 ();
 sg13g2_decap_8 FILLER_65_2521 ();
 sg13g2_decap_8 FILLER_65_2528 ();
 sg13g2_decap_8 FILLER_65_2535 ();
 sg13g2_decap_8 FILLER_65_2542 ();
 sg13g2_decap_8 FILLER_65_2549 ();
 sg13g2_decap_8 FILLER_65_2556 ();
 sg13g2_decap_8 FILLER_65_2563 ();
 sg13g2_decap_8 FILLER_65_2570 ();
 sg13g2_decap_8 FILLER_65_2577 ();
 sg13g2_decap_8 FILLER_65_2584 ();
 sg13g2_decap_8 FILLER_65_2591 ();
 sg13g2_decap_8 FILLER_65_2598 ();
 sg13g2_decap_8 FILLER_65_2605 ();
 sg13g2_decap_8 FILLER_65_2612 ();
 sg13g2_decap_8 FILLER_65_2619 ();
 sg13g2_decap_8 FILLER_65_2626 ();
 sg13g2_decap_8 FILLER_65_2633 ();
 sg13g2_decap_8 FILLER_65_2640 ();
 sg13g2_decap_8 FILLER_65_2647 ();
 sg13g2_decap_8 FILLER_65_2654 ();
 sg13g2_decap_8 FILLER_65_2661 ();
 sg13g2_decap_4 FILLER_65_2668 ();
 sg13g2_fill_2 FILLER_65_2672 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_126 ();
 sg13g2_decap_8 FILLER_66_133 ();
 sg13g2_decap_8 FILLER_66_140 ();
 sg13g2_decap_8 FILLER_66_147 ();
 sg13g2_decap_8 FILLER_66_154 ();
 sg13g2_decap_8 FILLER_66_161 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_decap_8 FILLER_66_175 ();
 sg13g2_decap_8 FILLER_66_182 ();
 sg13g2_decap_8 FILLER_66_189 ();
 sg13g2_decap_8 FILLER_66_196 ();
 sg13g2_decap_8 FILLER_66_203 ();
 sg13g2_decap_8 FILLER_66_210 ();
 sg13g2_decap_8 FILLER_66_217 ();
 sg13g2_decap_8 FILLER_66_224 ();
 sg13g2_decap_8 FILLER_66_231 ();
 sg13g2_decap_8 FILLER_66_238 ();
 sg13g2_decap_8 FILLER_66_245 ();
 sg13g2_decap_8 FILLER_66_252 ();
 sg13g2_decap_8 FILLER_66_259 ();
 sg13g2_decap_8 FILLER_66_266 ();
 sg13g2_decap_8 FILLER_66_273 ();
 sg13g2_decap_8 FILLER_66_280 ();
 sg13g2_decap_8 FILLER_66_287 ();
 sg13g2_decap_8 FILLER_66_294 ();
 sg13g2_decap_8 FILLER_66_301 ();
 sg13g2_decap_8 FILLER_66_308 ();
 sg13g2_decap_8 FILLER_66_315 ();
 sg13g2_decap_8 FILLER_66_322 ();
 sg13g2_decap_8 FILLER_66_329 ();
 sg13g2_decap_8 FILLER_66_336 ();
 sg13g2_decap_8 FILLER_66_343 ();
 sg13g2_decap_8 FILLER_66_350 ();
 sg13g2_decap_8 FILLER_66_357 ();
 sg13g2_decap_8 FILLER_66_364 ();
 sg13g2_decap_8 FILLER_66_371 ();
 sg13g2_decap_8 FILLER_66_378 ();
 sg13g2_decap_8 FILLER_66_385 ();
 sg13g2_decap_8 FILLER_66_392 ();
 sg13g2_decap_8 FILLER_66_399 ();
 sg13g2_decap_8 FILLER_66_406 ();
 sg13g2_decap_8 FILLER_66_413 ();
 sg13g2_decap_8 FILLER_66_420 ();
 sg13g2_fill_1 FILLER_66_427 ();
 sg13g2_fill_2 FILLER_66_481 ();
 sg13g2_fill_1 FILLER_66_483 ();
 sg13g2_fill_1 FILLER_66_517 ();
 sg13g2_fill_1 FILLER_66_537 ();
 sg13g2_fill_2 FILLER_66_547 ();
 sg13g2_fill_1 FILLER_66_549 ();
 sg13g2_fill_1 FILLER_66_559 ();
 sg13g2_fill_2 FILLER_66_631 ();
 sg13g2_fill_2 FILLER_66_643 ();
 sg13g2_fill_1 FILLER_66_645 ();
 sg13g2_fill_2 FILLER_66_651 ();
 sg13g2_fill_1 FILLER_66_653 ();
 sg13g2_fill_2 FILLER_66_664 ();
 sg13g2_fill_1 FILLER_66_666 ();
 sg13g2_fill_2 FILLER_66_672 ();
 sg13g2_fill_1 FILLER_66_674 ();
 sg13g2_decap_8 FILLER_66_701 ();
 sg13g2_decap_4 FILLER_66_708 ();
 sg13g2_fill_2 FILLER_66_712 ();
 sg13g2_fill_2 FILLER_66_740 ();
 sg13g2_fill_2 FILLER_66_746 ();
 sg13g2_decap_8 FILLER_66_752 ();
 sg13g2_decap_8 FILLER_66_759 ();
 sg13g2_decap_8 FILLER_66_785 ();
 sg13g2_fill_1 FILLER_66_792 ();
 sg13g2_fill_1 FILLER_66_805 ();
 sg13g2_fill_2 FILLER_66_812 ();
 sg13g2_decap_4 FILLER_66_819 ();
 sg13g2_decap_4 FILLER_66_843 ();
 sg13g2_fill_2 FILLER_66_847 ();
 sg13g2_fill_1 FILLER_66_875 ();
 sg13g2_fill_1 FILLER_66_915 ();
 sg13g2_fill_1 FILLER_66_995 ();
 sg13g2_fill_2 FILLER_66_1063 ();
 sg13g2_fill_2 FILLER_66_1098 ();
 sg13g2_fill_1 FILLER_66_1196 ();
 sg13g2_fill_1 FILLER_66_1256 ();
 sg13g2_fill_2 FILLER_66_1295 ();
 sg13g2_fill_1 FILLER_66_1374 ();
 sg13g2_fill_1 FILLER_66_1483 ();
 sg13g2_fill_1 FILLER_66_1595 ();
 sg13g2_fill_2 FILLER_66_1690 ();
 sg13g2_fill_1 FILLER_66_1692 ();
 sg13g2_fill_1 FILLER_66_1702 ();
 sg13g2_fill_2 FILLER_66_1789 ();
 sg13g2_fill_1 FILLER_66_1811 ();
 sg13g2_fill_2 FILLER_66_1846 ();
 sg13g2_fill_1 FILLER_66_1848 ();
 sg13g2_fill_2 FILLER_66_1875 ();
 sg13g2_fill_1 FILLER_66_1877 ();
 sg13g2_fill_2 FILLER_66_1933 ();
 sg13g2_fill_1 FILLER_66_1935 ();
 sg13g2_fill_2 FILLER_66_1954 ();
 sg13g2_fill_2 FILLER_66_1971 ();
 sg13g2_fill_2 FILLER_66_2009 ();
 sg13g2_fill_1 FILLER_66_2011 ();
 sg13g2_fill_2 FILLER_66_2048 ();
 sg13g2_fill_1 FILLER_66_2050 ();
 sg13g2_fill_1 FILLER_66_2060 ();
 sg13g2_fill_2 FILLER_66_2080 ();
 sg13g2_fill_2 FILLER_66_2140 ();
 sg13g2_fill_1 FILLER_66_2142 ();
 sg13g2_fill_2 FILLER_66_2178 ();
 sg13g2_fill_1 FILLER_66_2180 ();
 sg13g2_fill_2 FILLER_66_2248 ();
 sg13g2_fill_2 FILLER_66_2284 ();
 sg13g2_fill_1 FILLER_66_2286 ();
 sg13g2_decap_8 FILLER_66_2326 ();
 sg13g2_decap_8 FILLER_66_2333 ();
 sg13g2_decap_8 FILLER_66_2340 ();
 sg13g2_decap_8 FILLER_66_2347 ();
 sg13g2_decap_8 FILLER_66_2354 ();
 sg13g2_decap_8 FILLER_66_2361 ();
 sg13g2_decap_8 FILLER_66_2368 ();
 sg13g2_decap_8 FILLER_66_2375 ();
 sg13g2_decap_8 FILLER_66_2382 ();
 sg13g2_decap_8 FILLER_66_2389 ();
 sg13g2_decap_8 FILLER_66_2396 ();
 sg13g2_decap_8 FILLER_66_2403 ();
 sg13g2_decap_8 FILLER_66_2410 ();
 sg13g2_decap_8 FILLER_66_2417 ();
 sg13g2_decap_8 FILLER_66_2424 ();
 sg13g2_decap_8 FILLER_66_2431 ();
 sg13g2_decap_8 FILLER_66_2438 ();
 sg13g2_decap_8 FILLER_66_2445 ();
 sg13g2_decap_8 FILLER_66_2452 ();
 sg13g2_decap_8 FILLER_66_2459 ();
 sg13g2_decap_8 FILLER_66_2466 ();
 sg13g2_decap_8 FILLER_66_2473 ();
 sg13g2_decap_8 FILLER_66_2480 ();
 sg13g2_decap_8 FILLER_66_2487 ();
 sg13g2_decap_8 FILLER_66_2494 ();
 sg13g2_decap_8 FILLER_66_2501 ();
 sg13g2_decap_8 FILLER_66_2508 ();
 sg13g2_decap_8 FILLER_66_2515 ();
 sg13g2_decap_8 FILLER_66_2522 ();
 sg13g2_decap_8 FILLER_66_2529 ();
 sg13g2_decap_8 FILLER_66_2536 ();
 sg13g2_decap_8 FILLER_66_2543 ();
 sg13g2_decap_8 FILLER_66_2550 ();
 sg13g2_decap_8 FILLER_66_2557 ();
 sg13g2_decap_8 FILLER_66_2564 ();
 sg13g2_decap_8 FILLER_66_2571 ();
 sg13g2_decap_8 FILLER_66_2578 ();
 sg13g2_decap_8 FILLER_66_2585 ();
 sg13g2_decap_8 FILLER_66_2592 ();
 sg13g2_decap_8 FILLER_66_2599 ();
 sg13g2_decap_8 FILLER_66_2606 ();
 sg13g2_decap_8 FILLER_66_2613 ();
 sg13g2_decap_8 FILLER_66_2620 ();
 sg13g2_decap_8 FILLER_66_2627 ();
 sg13g2_decap_8 FILLER_66_2634 ();
 sg13g2_decap_8 FILLER_66_2641 ();
 sg13g2_decap_8 FILLER_66_2648 ();
 sg13g2_decap_8 FILLER_66_2655 ();
 sg13g2_decap_8 FILLER_66_2662 ();
 sg13g2_decap_4 FILLER_66_2669 ();
 sg13g2_fill_1 FILLER_66_2673 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_decap_8 FILLER_67_154 ();
 sg13g2_decap_8 FILLER_67_161 ();
 sg13g2_decap_8 FILLER_67_168 ();
 sg13g2_decap_8 FILLER_67_175 ();
 sg13g2_decap_8 FILLER_67_182 ();
 sg13g2_decap_8 FILLER_67_189 ();
 sg13g2_decap_8 FILLER_67_196 ();
 sg13g2_decap_8 FILLER_67_203 ();
 sg13g2_decap_8 FILLER_67_210 ();
 sg13g2_decap_8 FILLER_67_217 ();
 sg13g2_decap_8 FILLER_67_224 ();
 sg13g2_decap_8 FILLER_67_231 ();
 sg13g2_decap_8 FILLER_67_238 ();
 sg13g2_decap_8 FILLER_67_245 ();
 sg13g2_decap_8 FILLER_67_252 ();
 sg13g2_decap_8 FILLER_67_259 ();
 sg13g2_decap_8 FILLER_67_266 ();
 sg13g2_decap_8 FILLER_67_273 ();
 sg13g2_decap_8 FILLER_67_280 ();
 sg13g2_decap_8 FILLER_67_287 ();
 sg13g2_decap_8 FILLER_67_294 ();
 sg13g2_decap_8 FILLER_67_301 ();
 sg13g2_decap_8 FILLER_67_308 ();
 sg13g2_decap_8 FILLER_67_315 ();
 sg13g2_decap_8 FILLER_67_322 ();
 sg13g2_decap_8 FILLER_67_329 ();
 sg13g2_decap_8 FILLER_67_336 ();
 sg13g2_decap_8 FILLER_67_343 ();
 sg13g2_decap_8 FILLER_67_350 ();
 sg13g2_decap_8 FILLER_67_357 ();
 sg13g2_decap_8 FILLER_67_364 ();
 sg13g2_decap_8 FILLER_67_371 ();
 sg13g2_decap_8 FILLER_67_378 ();
 sg13g2_decap_8 FILLER_67_385 ();
 sg13g2_decap_8 FILLER_67_392 ();
 sg13g2_decap_8 FILLER_67_399 ();
 sg13g2_decap_8 FILLER_67_406 ();
 sg13g2_decap_8 FILLER_67_413 ();
 sg13g2_decap_8 FILLER_67_420 ();
 sg13g2_decap_8 FILLER_67_427 ();
 sg13g2_fill_2 FILLER_67_496 ();
 sg13g2_fill_1 FILLER_67_547 ();
 sg13g2_fill_2 FILLER_67_574 ();
 sg13g2_fill_1 FILLER_67_630 ();
 sg13g2_fill_2 FILLER_67_653 ();
 sg13g2_fill_1 FILLER_67_655 ();
 sg13g2_fill_2 FILLER_67_661 ();
 sg13g2_fill_1 FILLER_67_663 ();
 sg13g2_fill_2 FILLER_67_707 ();
 sg13g2_decap_4 FILLER_67_718 ();
 sg13g2_fill_2 FILLER_67_722 ();
 sg13g2_decap_8 FILLER_67_728 ();
 sg13g2_decap_4 FILLER_67_735 ();
 sg13g2_fill_2 FILLER_67_739 ();
 sg13g2_fill_2 FILLER_67_767 ();
 sg13g2_fill_2 FILLER_67_779 ();
 sg13g2_fill_1 FILLER_67_781 ();
 sg13g2_decap_4 FILLER_67_799 ();
 sg13g2_fill_1 FILLER_67_839 ();
 sg13g2_fill_2 FILLER_67_853 ();
 sg13g2_fill_1 FILLER_67_868 ();
 sg13g2_fill_2 FILLER_67_914 ();
 sg13g2_fill_1 FILLER_67_921 ();
 sg13g2_fill_2 FILLER_67_948 ();
 sg13g2_fill_1 FILLER_67_1100 ();
 sg13g2_fill_2 FILLER_67_1115 ();
 sg13g2_fill_1 FILLER_67_1144 ();
 sg13g2_fill_1 FILLER_67_1190 ();
 sg13g2_fill_2 FILLER_67_1295 ();
 sg13g2_fill_2 FILLER_67_1302 ();
 sg13g2_fill_1 FILLER_67_1309 ();
 sg13g2_fill_2 FILLER_67_1457 ();
 sg13g2_fill_2 FILLER_67_1468 ();
 sg13g2_fill_1 FILLER_67_1510 ();
 sg13g2_fill_1 FILLER_67_1559 ();
 sg13g2_fill_2 FILLER_67_1585 ();
 sg13g2_fill_2 FILLER_67_1622 ();
 sg13g2_fill_2 FILLER_67_1675 ();
 sg13g2_fill_1 FILLER_67_1711 ();
 sg13g2_fill_1 FILLER_67_1722 ();
 sg13g2_fill_2 FILLER_67_1776 ();
 sg13g2_fill_1 FILLER_67_1778 ();
 sg13g2_fill_2 FILLER_67_1821 ();
 sg13g2_fill_1 FILLER_67_1823 ();
 sg13g2_fill_2 FILLER_67_1863 ();
 sg13g2_fill_1 FILLER_67_1865 ();
 sg13g2_fill_2 FILLER_67_1932 ();
 sg13g2_decap_4 FILLER_67_1943 ();
 sg13g2_fill_2 FILLER_67_1947 ();
 sg13g2_decap_4 FILLER_67_1959 ();
 sg13g2_fill_2 FILLER_67_2018 ();
 sg13g2_decap_4 FILLER_67_2046 ();
 sg13g2_fill_1 FILLER_67_2050 ();
 sg13g2_fill_1 FILLER_67_2132 ();
 sg13g2_fill_2 FILLER_67_2174 ();
 sg13g2_fill_2 FILLER_67_2199 ();
 sg13g2_decap_8 FILLER_67_2216 ();
 sg13g2_fill_1 FILLER_67_2223 ();
 sg13g2_fill_1 FILLER_67_2241 ();
 sg13g2_decap_8 FILLER_67_2247 ();
 sg13g2_fill_2 FILLER_67_2275 ();
 sg13g2_fill_2 FILLER_67_2282 ();
 sg13g2_fill_2 FILLER_67_2309 ();
 sg13g2_decap_8 FILLER_67_2337 ();
 sg13g2_decap_8 FILLER_67_2344 ();
 sg13g2_decap_8 FILLER_67_2351 ();
 sg13g2_decap_8 FILLER_67_2358 ();
 sg13g2_decap_8 FILLER_67_2365 ();
 sg13g2_decap_8 FILLER_67_2372 ();
 sg13g2_decap_8 FILLER_67_2379 ();
 sg13g2_decap_8 FILLER_67_2386 ();
 sg13g2_decap_8 FILLER_67_2393 ();
 sg13g2_decap_8 FILLER_67_2400 ();
 sg13g2_decap_8 FILLER_67_2407 ();
 sg13g2_decap_8 FILLER_67_2414 ();
 sg13g2_decap_8 FILLER_67_2421 ();
 sg13g2_decap_8 FILLER_67_2428 ();
 sg13g2_decap_8 FILLER_67_2435 ();
 sg13g2_decap_8 FILLER_67_2442 ();
 sg13g2_decap_8 FILLER_67_2449 ();
 sg13g2_decap_8 FILLER_67_2456 ();
 sg13g2_decap_8 FILLER_67_2463 ();
 sg13g2_decap_8 FILLER_67_2470 ();
 sg13g2_decap_8 FILLER_67_2477 ();
 sg13g2_decap_8 FILLER_67_2484 ();
 sg13g2_decap_8 FILLER_67_2491 ();
 sg13g2_decap_8 FILLER_67_2498 ();
 sg13g2_decap_8 FILLER_67_2505 ();
 sg13g2_decap_8 FILLER_67_2512 ();
 sg13g2_decap_8 FILLER_67_2519 ();
 sg13g2_decap_8 FILLER_67_2526 ();
 sg13g2_decap_8 FILLER_67_2533 ();
 sg13g2_decap_8 FILLER_67_2540 ();
 sg13g2_decap_8 FILLER_67_2547 ();
 sg13g2_decap_8 FILLER_67_2554 ();
 sg13g2_decap_8 FILLER_67_2561 ();
 sg13g2_decap_8 FILLER_67_2568 ();
 sg13g2_decap_8 FILLER_67_2575 ();
 sg13g2_decap_8 FILLER_67_2582 ();
 sg13g2_decap_8 FILLER_67_2589 ();
 sg13g2_decap_8 FILLER_67_2596 ();
 sg13g2_decap_8 FILLER_67_2603 ();
 sg13g2_decap_8 FILLER_67_2610 ();
 sg13g2_decap_8 FILLER_67_2617 ();
 sg13g2_decap_8 FILLER_67_2624 ();
 sg13g2_decap_8 FILLER_67_2631 ();
 sg13g2_decap_8 FILLER_67_2638 ();
 sg13g2_decap_8 FILLER_67_2645 ();
 sg13g2_decap_8 FILLER_67_2652 ();
 sg13g2_decap_8 FILLER_67_2659 ();
 sg13g2_decap_8 FILLER_67_2666 ();
 sg13g2_fill_1 FILLER_67_2673 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_decap_8 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_decap_8 FILLER_68_147 ();
 sg13g2_decap_8 FILLER_68_154 ();
 sg13g2_decap_8 FILLER_68_161 ();
 sg13g2_decap_8 FILLER_68_168 ();
 sg13g2_decap_8 FILLER_68_175 ();
 sg13g2_decap_8 FILLER_68_182 ();
 sg13g2_decap_8 FILLER_68_189 ();
 sg13g2_decap_8 FILLER_68_196 ();
 sg13g2_decap_8 FILLER_68_203 ();
 sg13g2_decap_8 FILLER_68_210 ();
 sg13g2_decap_8 FILLER_68_217 ();
 sg13g2_decap_8 FILLER_68_224 ();
 sg13g2_decap_8 FILLER_68_231 ();
 sg13g2_decap_8 FILLER_68_238 ();
 sg13g2_decap_8 FILLER_68_245 ();
 sg13g2_decap_8 FILLER_68_252 ();
 sg13g2_decap_8 FILLER_68_259 ();
 sg13g2_decap_8 FILLER_68_266 ();
 sg13g2_decap_8 FILLER_68_273 ();
 sg13g2_decap_8 FILLER_68_280 ();
 sg13g2_decap_8 FILLER_68_287 ();
 sg13g2_decap_8 FILLER_68_294 ();
 sg13g2_decap_8 FILLER_68_301 ();
 sg13g2_decap_8 FILLER_68_308 ();
 sg13g2_decap_8 FILLER_68_315 ();
 sg13g2_decap_8 FILLER_68_322 ();
 sg13g2_decap_8 FILLER_68_329 ();
 sg13g2_decap_8 FILLER_68_336 ();
 sg13g2_decap_8 FILLER_68_343 ();
 sg13g2_decap_8 FILLER_68_350 ();
 sg13g2_decap_8 FILLER_68_357 ();
 sg13g2_decap_8 FILLER_68_364 ();
 sg13g2_decap_8 FILLER_68_371 ();
 sg13g2_decap_8 FILLER_68_378 ();
 sg13g2_decap_8 FILLER_68_385 ();
 sg13g2_decap_8 FILLER_68_392 ();
 sg13g2_decap_8 FILLER_68_399 ();
 sg13g2_decap_8 FILLER_68_406 ();
 sg13g2_decap_8 FILLER_68_413 ();
 sg13g2_decap_4 FILLER_68_420 ();
 sg13g2_fill_1 FILLER_68_424 ();
 sg13g2_fill_2 FILLER_68_462 ();
 sg13g2_fill_2 FILLER_68_482 ();
 sg13g2_fill_1 FILLER_68_484 ();
 sg13g2_fill_1 FILLER_68_518 ();
 sg13g2_fill_2 FILLER_68_545 ();
 sg13g2_fill_2 FILLER_68_651 ();
 sg13g2_decap_8 FILLER_68_721 ();
 sg13g2_decap_8 FILLER_68_728 ();
 sg13g2_decap_8 FILLER_68_735 ();
 sg13g2_decap_8 FILLER_68_742 ();
 sg13g2_fill_2 FILLER_68_749 ();
 sg13g2_fill_1 FILLER_68_751 ();
 sg13g2_decap_8 FILLER_68_756 ();
 sg13g2_decap_8 FILLER_68_763 ();
 sg13g2_decap_8 FILLER_68_770 ();
 sg13g2_fill_2 FILLER_68_777 ();
 sg13g2_decap_4 FILLER_68_797 ();
 sg13g2_fill_2 FILLER_68_816 ();
 sg13g2_fill_2 FILLER_68_823 ();
 sg13g2_fill_2 FILLER_68_829 ();
 sg13g2_fill_2 FILLER_68_842 ();
 sg13g2_fill_1 FILLER_68_844 ();
 sg13g2_fill_1 FILLER_68_874 ();
 sg13g2_fill_2 FILLER_68_883 ();
 sg13g2_fill_2 FILLER_68_1018 ();
 sg13g2_fill_2 FILLER_68_1062 ();
 sg13g2_fill_1 FILLER_68_1073 ();
 sg13g2_fill_1 FILLER_68_1115 ();
 sg13g2_fill_1 FILLER_68_1125 ();
 sg13g2_fill_2 FILLER_68_1131 ();
 sg13g2_fill_2 FILLER_68_1201 ();
 sg13g2_fill_1 FILLER_68_1212 ();
 sg13g2_fill_1 FILLER_68_1232 ();
 sg13g2_fill_2 FILLER_68_1404 ();
 sg13g2_fill_2 FILLER_68_1486 ();
 sg13g2_fill_1 FILLER_68_1515 ();
 sg13g2_fill_2 FILLER_68_1545 ();
 sg13g2_fill_2 FILLER_68_1567 ();
 sg13g2_fill_1 FILLER_68_1569 ();
 sg13g2_decap_4 FILLER_68_1587 ();
 sg13g2_fill_1 FILLER_68_1591 ();
 sg13g2_decap_4 FILLER_68_1597 ();
 sg13g2_fill_1 FILLER_68_1601 ();
 sg13g2_fill_2 FILLER_68_1693 ();
 sg13g2_fill_1 FILLER_68_1695 ();
 sg13g2_fill_2 FILLER_68_1730 ();
 sg13g2_fill_1 FILLER_68_1732 ();
 sg13g2_fill_1 FILLER_68_1743 ();
 sg13g2_fill_2 FILLER_68_1771 ();
 sg13g2_fill_1 FILLER_68_1784 ();
 sg13g2_decap_4 FILLER_68_1797 ();
 sg13g2_fill_2 FILLER_68_1809 ();
 sg13g2_fill_1 FILLER_68_1811 ();
 sg13g2_fill_2 FILLER_68_1863 ();
 sg13g2_fill_1 FILLER_68_1891 ();
 sg13g2_fill_2 FILLER_68_1926 ();
 sg13g2_fill_1 FILLER_68_1928 ();
 sg13g2_fill_1 FILLER_68_1976 ();
 sg13g2_fill_2 FILLER_68_1995 ();
 sg13g2_fill_2 FILLER_68_2013 ();
 sg13g2_fill_1 FILLER_68_2015 ();
 sg13g2_fill_1 FILLER_68_2052 ();
 sg13g2_decap_8 FILLER_68_2057 ();
 sg13g2_fill_2 FILLER_68_2074 ();
 sg13g2_fill_2 FILLER_68_2099 ();
 sg13g2_fill_1 FILLER_68_2148 ();
 sg13g2_fill_1 FILLER_68_2176 ();
 sg13g2_fill_2 FILLER_68_2191 ();
 sg13g2_decap_4 FILLER_68_2208 ();
 sg13g2_fill_1 FILLER_68_2233 ();
 sg13g2_fill_2 FILLER_68_2254 ();
 sg13g2_fill_1 FILLER_68_2256 ();
 sg13g2_decap_4 FILLER_68_2269 ();
 sg13g2_fill_1 FILLER_68_2273 ();
 sg13g2_fill_2 FILLER_68_2279 ();
 sg13g2_fill_1 FILLER_68_2281 ();
 sg13g2_fill_2 FILLER_68_2287 ();
 sg13g2_decap_4 FILLER_68_2315 ();
 sg13g2_fill_1 FILLER_68_2319 ();
 sg13g2_decap_8 FILLER_68_2333 ();
 sg13g2_decap_8 FILLER_68_2340 ();
 sg13g2_decap_8 FILLER_68_2347 ();
 sg13g2_decap_8 FILLER_68_2354 ();
 sg13g2_decap_8 FILLER_68_2361 ();
 sg13g2_decap_8 FILLER_68_2368 ();
 sg13g2_decap_8 FILLER_68_2375 ();
 sg13g2_decap_8 FILLER_68_2382 ();
 sg13g2_decap_8 FILLER_68_2389 ();
 sg13g2_decap_8 FILLER_68_2396 ();
 sg13g2_decap_8 FILLER_68_2403 ();
 sg13g2_decap_8 FILLER_68_2410 ();
 sg13g2_decap_8 FILLER_68_2417 ();
 sg13g2_decap_8 FILLER_68_2424 ();
 sg13g2_decap_8 FILLER_68_2431 ();
 sg13g2_decap_8 FILLER_68_2438 ();
 sg13g2_decap_8 FILLER_68_2445 ();
 sg13g2_decap_8 FILLER_68_2452 ();
 sg13g2_decap_8 FILLER_68_2459 ();
 sg13g2_decap_8 FILLER_68_2466 ();
 sg13g2_decap_8 FILLER_68_2473 ();
 sg13g2_decap_8 FILLER_68_2480 ();
 sg13g2_decap_8 FILLER_68_2487 ();
 sg13g2_decap_8 FILLER_68_2494 ();
 sg13g2_decap_8 FILLER_68_2501 ();
 sg13g2_decap_8 FILLER_68_2508 ();
 sg13g2_decap_8 FILLER_68_2515 ();
 sg13g2_decap_8 FILLER_68_2522 ();
 sg13g2_decap_8 FILLER_68_2529 ();
 sg13g2_decap_8 FILLER_68_2536 ();
 sg13g2_decap_8 FILLER_68_2543 ();
 sg13g2_decap_8 FILLER_68_2550 ();
 sg13g2_decap_8 FILLER_68_2557 ();
 sg13g2_decap_8 FILLER_68_2564 ();
 sg13g2_decap_8 FILLER_68_2571 ();
 sg13g2_decap_8 FILLER_68_2578 ();
 sg13g2_decap_8 FILLER_68_2585 ();
 sg13g2_decap_8 FILLER_68_2592 ();
 sg13g2_decap_8 FILLER_68_2599 ();
 sg13g2_decap_8 FILLER_68_2606 ();
 sg13g2_decap_8 FILLER_68_2613 ();
 sg13g2_decap_8 FILLER_68_2620 ();
 sg13g2_decap_8 FILLER_68_2627 ();
 sg13g2_decap_8 FILLER_68_2634 ();
 sg13g2_decap_8 FILLER_68_2641 ();
 sg13g2_decap_8 FILLER_68_2648 ();
 sg13g2_decap_8 FILLER_68_2655 ();
 sg13g2_decap_8 FILLER_68_2662 ();
 sg13g2_decap_4 FILLER_68_2669 ();
 sg13g2_fill_1 FILLER_68_2673 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_decap_8 FILLER_69_133 ();
 sg13g2_decap_8 FILLER_69_140 ();
 sg13g2_decap_8 FILLER_69_147 ();
 sg13g2_decap_8 FILLER_69_154 ();
 sg13g2_decap_8 FILLER_69_161 ();
 sg13g2_decap_8 FILLER_69_168 ();
 sg13g2_decap_8 FILLER_69_175 ();
 sg13g2_decap_8 FILLER_69_182 ();
 sg13g2_decap_8 FILLER_69_189 ();
 sg13g2_decap_8 FILLER_69_196 ();
 sg13g2_decap_8 FILLER_69_203 ();
 sg13g2_decap_8 FILLER_69_210 ();
 sg13g2_decap_8 FILLER_69_217 ();
 sg13g2_decap_8 FILLER_69_224 ();
 sg13g2_decap_8 FILLER_69_231 ();
 sg13g2_decap_8 FILLER_69_238 ();
 sg13g2_decap_8 FILLER_69_245 ();
 sg13g2_decap_8 FILLER_69_252 ();
 sg13g2_decap_8 FILLER_69_259 ();
 sg13g2_decap_8 FILLER_69_266 ();
 sg13g2_decap_8 FILLER_69_273 ();
 sg13g2_decap_8 FILLER_69_280 ();
 sg13g2_decap_8 FILLER_69_287 ();
 sg13g2_decap_8 FILLER_69_294 ();
 sg13g2_decap_8 FILLER_69_301 ();
 sg13g2_decap_8 FILLER_69_308 ();
 sg13g2_decap_8 FILLER_69_315 ();
 sg13g2_decap_8 FILLER_69_322 ();
 sg13g2_decap_8 FILLER_69_329 ();
 sg13g2_decap_8 FILLER_69_336 ();
 sg13g2_decap_8 FILLER_69_343 ();
 sg13g2_decap_8 FILLER_69_350 ();
 sg13g2_decap_8 FILLER_69_357 ();
 sg13g2_decap_8 FILLER_69_364 ();
 sg13g2_decap_8 FILLER_69_371 ();
 sg13g2_decap_8 FILLER_69_378 ();
 sg13g2_decap_8 FILLER_69_385 ();
 sg13g2_decap_8 FILLER_69_392 ();
 sg13g2_decap_8 FILLER_69_399 ();
 sg13g2_decap_8 FILLER_69_406 ();
 sg13g2_decap_8 FILLER_69_413 ();
 sg13g2_decap_8 FILLER_69_420 ();
 sg13g2_decap_4 FILLER_69_427 ();
 sg13g2_fill_2 FILLER_69_431 ();
 sg13g2_fill_2 FILLER_69_529 ();
 sg13g2_fill_1 FILLER_69_555 ();
 sg13g2_fill_2 FILLER_69_596 ();
 sg13g2_fill_1 FILLER_69_607 ();
 sg13g2_fill_1 FILLER_69_644 ();
 sg13g2_fill_1 FILLER_69_658 ();
 sg13g2_fill_2 FILLER_69_668 ();
 sg13g2_fill_2 FILLER_69_701 ();
 sg13g2_decap_8 FILLER_69_711 ();
 sg13g2_decap_8 FILLER_69_718 ();
 sg13g2_decap_8 FILLER_69_725 ();
 sg13g2_decap_8 FILLER_69_732 ();
 sg13g2_decap_8 FILLER_69_739 ();
 sg13g2_decap_8 FILLER_69_746 ();
 sg13g2_decap_8 FILLER_69_753 ();
 sg13g2_decap_8 FILLER_69_760 ();
 sg13g2_decap_8 FILLER_69_767 ();
 sg13g2_decap_8 FILLER_69_774 ();
 sg13g2_decap_4 FILLER_69_820 ();
 sg13g2_fill_2 FILLER_69_824 ();
 sg13g2_decap_4 FILLER_69_841 ();
 sg13g2_fill_2 FILLER_69_845 ();
 sg13g2_fill_1 FILLER_69_850 ();
 sg13g2_fill_1 FILLER_69_855 ();
 sg13g2_fill_2 FILLER_69_869 ();
 sg13g2_fill_2 FILLER_69_910 ();
 sg13g2_fill_1 FILLER_69_924 ();
 sg13g2_fill_2 FILLER_69_937 ();
 sg13g2_fill_1 FILLER_69_985 ();
 sg13g2_fill_1 FILLER_69_1099 ();
 sg13g2_fill_2 FILLER_69_1126 ();
 sg13g2_fill_2 FILLER_69_1379 ();
 sg13g2_fill_2 FILLER_69_1433 ();
 sg13g2_fill_1 FILLER_69_1471 ();
 sg13g2_fill_2 FILLER_69_1493 ();
 sg13g2_fill_1 FILLER_69_1504 ();
 sg13g2_fill_1 FILLER_69_1547 ();
 sg13g2_fill_2 FILLER_69_1553 ();
 sg13g2_fill_1 FILLER_69_1564 ();
 sg13g2_decap_4 FILLER_69_1587 ();
 sg13g2_decap_8 FILLER_69_1614 ();
 sg13g2_decap_4 FILLER_69_1625 ();
 sg13g2_fill_2 FILLER_69_1629 ();
 sg13g2_fill_2 FILLER_69_1664 ();
 sg13g2_decap_4 FILLER_69_1761 ();
 sg13g2_fill_1 FILLER_69_1765 ();
 sg13g2_fill_1 FILLER_69_1787 ();
 sg13g2_fill_2 FILLER_69_1793 ();
 sg13g2_fill_2 FILLER_69_1808 ();
 sg13g2_decap_4 FILLER_69_1820 ();
 sg13g2_fill_1 FILLER_69_1833 ();
 sg13g2_decap_4 FILLER_69_1856 ();
 sg13g2_fill_1 FILLER_69_1860 ();
 sg13g2_fill_2 FILLER_69_1871 ();
 sg13g2_fill_2 FILLER_69_1914 ();
 sg13g2_decap_8 FILLER_69_1932 ();
 sg13g2_fill_1 FILLER_69_1939 ();
 sg13g2_decap_4 FILLER_69_1953 ();
 sg13g2_fill_1 FILLER_69_1957 ();
 sg13g2_fill_2 FILLER_69_1963 ();
 sg13g2_decap_4 FILLER_69_1970 ();
 sg13g2_decap_8 FILLER_69_1982 ();
 sg13g2_fill_1 FILLER_69_1989 ();
 sg13g2_fill_1 FILLER_69_2000 ();
 sg13g2_fill_2 FILLER_69_2007 ();
 sg13g2_fill_2 FILLER_69_2117 ();
 sg13g2_fill_1 FILLER_69_2119 ();
 sg13g2_fill_2 FILLER_69_2160 ();
 sg13g2_fill_1 FILLER_69_2162 ();
 sg13g2_fill_2 FILLER_69_2176 ();
 sg13g2_fill_1 FILLER_69_2178 ();
 sg13g2_fill_2 FILLER_69_2256 ();
 sg13g2_fill_2 FILLER_69_2289 ();
 sg13g2_decap_8 FILLER_69_2336 ();
 sg13g2_decap_8 FILLER_69_2343 ();
 sg13g2_decap_8 FILLER_69_2350 ();
 sg13g2_decap_8 FILLER_69_2357 ();
 sg13g2_decap_8 FILLER_69_2364 ();
 sg13g2_decap_8 FILLER_69_2371 ();
 sg13g2_decap_8 FILLER_69_2378 ();
 sg13g2_decap_8 FILLER_69_2385 ();
 sg13g2_decap_8 FILLER_69_2392 ();
 sg13g2_decap_8 FILLER_69_2399 ();
 sg13g2_decap_8 FILLER_69_2406 ();
 sg13g2_decap_8 FILLER_69_2413 ();
 sg13g2_decap_8 FILLER_69_2420 ();
 sg13g2_decap_8 FILLER_69_2427 ();
 sg13g2_decap_8 FILLER_69_2434 ();
 sg13g2_decap_8 FILLER_69_2441 ();
 sg13g2_decap_8 FILLER_69_2448 ();
 sg13g2_decap_8 FILLER_69_2455 ();
 sg13g2_decap_8 FILLER_69_2462 ();
 sg13g2_decap_8 FILLER_69_2469 ();
 sg13g2_decap_8 FILLER_69_2476 ();
 sg13g2_decap_8 FILLER_69_2483 ();
 sg13g2_decap_8 FILLER_69_2490 ();
 sg13g2_decap_8 FILLER_69_2497 ();
 sg13g2_decap_8 FILLER_69_2504 ();
 sg13g2_decap_8 FILLER_69_2511 ();
 sg13g2_decap_8 FILLER_69_2518 ();
 sg13g2_decap_8 FILLER_69_2525 ();
 sg13g2_decap_8 FILLER_69_2532 ();
 sg13g2_decap_8 FILLER_69_2539 ();
 sg13g2_decap_8 FILLER_69_2546 ();
 sg13g2_decap_8 FILLER_69_2553 ();
 sg13g2_decap_8 FILLER_69_2560 ();
 sg13g2_decap_8 FILLER_69_2567 ();
 sg13g2_decap_8 FILLER_69_2574 ();
 sg13g2_decap_8 FILLER_69_2581 ();
 sg13g2_decap_8 FILLER_69_2588 ();
 sg13g2_decap_8 FILLER_69_2595 ();
 sg13g2_decap_8 FILLER_69_2602 ();
 sg13g2_decap_8 FILLER_69_2609 ();
 sg13g2_decap_8 FILLER_69_2616 ();
 sg13g2_decap_8 FILLER_69_2623 ();
 sg13g2_decap_8 FILLER_69_2630 ();
 sg13g2_decap_8 FILLER_69_2637 ();
 sg13g2_decap_8 FILLER_69_2644 ();
 sg13g2_decap_8 FILLER_69_2651 ();
 sg13g2_decap_8 FILLER_69_2658 ();
 sg13g2_decap_8 FILLER_69_2665 ();
 sg13g2_fill_2 FILLER_69_2672 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_decap_8 FILLER_70_161 ();
 sg13g2_decap_8 FILLER_70_168 ();
 sg13g2_decap_8 FILLER_70_175 ();
 sg13g2_decap_8 FILLER_70_182 ();
 sg13g2_decap_8 FILLER_70_189 ();
 sg13g2_decap_8 FILLER_70_196 ();
 sg13g2_decap_8 FILLER_70_203 ();
 sg13g2_decap_8 FILLER_70_210 ();
 sg13g2_decap_8 FILLER_70_217 ();
 sg13g2_decap_8 FILLER_70_224 ();
 sg13g2_decap_8 FILLER_70_231 ();
 sg13g2_decap_8 FILLER_70_238 ();
 sg13g2_decap_8 FILLER_70_245 ();
 sg13g2_decap_8 FILLER_70_252 ();
 sg13g2_decap_8 FILLER_70_259 ();
 sg13g2_decap_8 FILLER_70_266 ();
 sg13g2_decap_8 FILLER_70_273 ();
 sg13g2_decap_8 FILLER_70_280 ();
 sg13g2_decap_8 FILLER_70_287 ();
 sg13g2_decap_8 FILLER_70_294 ();
 sg13g2_decap_8 FILLER_70_301 ();
 sg13g2_decap_8 FILLER_70_308 ();
 sg13g2_decap_8 FILLER_70_315 ();
 sg13g2_decap_8 FILLER_70_322 ();
 sg13g2_decap_8 FILLER_70_329 ();
 sg13g2_decap_8 FILLER_70_336 ();
 sg13g2_decap_8 FILLER_70_343 ();
 sg13g2_decap_8 FILLER_70_350 ();
 sg13g2_decap_8 FILLER_70_357 ();
 sg13g2_decap_8 FILLER_70_364 ();
 sg13g2_decap_8 FILLER_70_371 ();
 sg13g2_decap_8 FILLER_70_378 ();
 sg13g2_decap_8 FILLER_70_385 ();
 sg13g2_decap_8 FILLER_70_392 ();
 sg13g2_decap_8 FILLER_70_399 ();
 sg13g2_decap_8 FILLER_70_406 ();
 sg13g2_decap_8 FILLER_70_413 ();
 sg13g2_decap_4 FILLER_70_420 ();
 sg13g2_fill_2 FILLER_70_499 ();
 sg13g2_fill_2 FILLER_70_559 ();
 sg13g2_fill_1 FILLER_70_582 ();
 sg13g2_fill_2 FILLER_70_635 ();
 sg13g2_fill_2 FILLER_70_689 ();
 sg13g2_decap_8 FILLER_70_722 ();
 sg13g2_decap_8 FILLER_70_729 ();
 sg13g2_decap_8 FILLER_70_736 ();
 sg13g2_decap_8 FILLER_70_743 ();
 sg13g2_decap_8 FILLER_70_750 ();
 sg13g2_decap_8 FILLER_70_757 ();
 sg13g2_decap_8 FILLER_70_764 ();
 sg13g2_decap_8 FILLER_70_771 ();
 sg13g2_decap_8 FILLER_70_778 ();
 sg13g2_decap_8 FILLER_70_785 ();
 sg13g2_decap_8 FILLER_70_798 ();
 sg13g2_decap_8 FILLER_70_805 ();
 sg13g2_fill_2 FILLER_70_812 ();
 sg13g2_decap_8 FILLER_70_820 ();
 sg13g2_fill_1 FILLER_70_835 ();
 sg13g2_fill_1 FILLER_70_842 ();
 sg13g2_fill_1 FILLER_70_864 ();
 sg13g2_fill_2 FILLER_70_928 ();
 sg13g2_fill_2 FILLER_70_936 ();
 sg13g2_fill_1 FILLER_70_978 ();
 sg13g2_fill_2 FILLER_70_1014 ();
 sg13g2_fill_2 FILLER_70_1045 ();
 sg13g2_fill_1 FILLER_70_1061 ();
 sg13g2_fill_2 FILLER_70_1071 ();
 sg13g2_fill_2 FILLER_70_1144 ();
 sg13g2_fill_1 FILLER_70_1177 ();
 sg13g2_fill_1 FILLER_70_1209 ();
 sg13g2_fill_2 FILLER_70_1255 ();
 sg13g2_fill_1 FILLER_70_1315 ();
 sg13g2_fill_2 FILLER_70_1325 ();
 sg13g2_fill_1 FILLER_70_1356 ();
 sg13g2_fill_1 FILLER_70_1394 ();
 sg13g2_fill_1 FILLER_70_1421 ();
 sg13g2_fill_1 FILLER_70_1450 ();
 sg13g2_fill_1 FILLER_70_1503 ();
 sg13g2_fill_2 FILLER_70_1533 ();
 sg13g2_fill_1 FILLER_70_1556 ();
 sg13g2_fill_2 FILLER_70_1565 ();
 sg13g2_fill_2 FILLER_70_1577 ();
 sg13g2_fill_1 FILLER_70_1579 ();
 sg13g2_decap_4 FILLER_70_1590 ();
 sg13g2_fill_2 FILLER_70_1594 ();
 sg13g2_decap_4 FILLER_70_1606 ();
 sg13g2_fill_1 FILLER_70_1610 ();
 sg13g2_decap_4 FILLER_70_1721 ();
 sg13g2_fill_1 FILLER_70_1725 ();
 sg13g2_fill_1 FILLER_70_1758 ();
 sg13g2_decap_4 FILLER_70_1768 ();
 sg13g2_fill_2 FILLER_70_1782 ();
 sg13g2_decap_4 FILLER_70_1789 ();
 sg13g2_fill_1 FILLER_70_1793 ();
 sg13g2_decap_4 FILLER_70_1810 ();
 sg13g2_fill_2 FILLER_70_1855 ();
 sg13g2_fill_1 FILLER_70_1857 ();
 sg13g2_decap_4 FILLER_70_1884 ();
 sg13g2_fill_1 FILLER_70_1888 ();
 sg13g2_fill_2 FILLER_70_1936 ();
 sg13g2_fill_1 FILLER_70_1938 ();
 sg13g2_decap_8 FILLER_70_1973 ();
 sg13g2_fill_1 FILLER_70_1980 ();
 sg13g2_decap_4 FILLER_70_1991 ();
 sg13g2_decap_8 FILLER_70_2021 ();
 sg13g2_fill_1 FILLER_70_2028 ();
 sg13g2_decap_8 FILLER_70_2042 ();
 sg13g2_fill_2 FILLER_70_2049 ();
 sg13g2_fill_1 FILLER_70_2051 ();
 sg13g2_decap_4 FILLER_70_2056 ();
 sg13g2_fill_1 FILLER_70_2060 ();
 sg13g2_fill_1 FILLER_70_2071 ();
 sg13g2_decap_4 FILLER_70_2091 ();
 sg13g2_fill_1 FILLER_70_2095 ();
 sg13g2_decap_4 FILLER_70_2117 ();
 sg13g2_fill_2 FILLER_70_2138 ();
 sg13g2_fill_1 FILLER_70_2140 ();
 sg13g2_fill_2 FILLER_70_2156 ();
 sg13g2_fill_1 FILLER_70_2158 ();
 sg13g2_fill_2 FILLER_70_2169 ();
 sg13g2_decap_8 FILLER_70_2176 ();
 sg13g2_decap_8 FILLER_70_2183 ();
 sg13g2_fill_2 FILLER_70_2194 ();
 sg13g2_fill_2 FILLER_70_2206 ();
 sg13g2_fill_1 FILLER_70_2208 ();
 sg13g2_decap_8 FILLER_70_2214 ();
 sg13g2_decap_8 FILLER_70_2221 ();
 sg13g2_decap_4 FILLER_70_2228 ();
 sg13g2_decap_8 FILLER_70_2237 ();
 sg13g2_fill_2 FILLER_70_2244 ();
 sg13g2_fill_2 FILLER_70_2272 ();
 sg13g2_fill_1 FILLER_70_2274 ();
 sg13g2_decap_8 FILLER_70_2311 ();
 sg13g2_fill_2 FILLER_70_2318 ();
 sg13g2_decap_8 FILLER_70_2329 ();
 sg13g2_decap_8 FILLER_70_2336 ();
 sg13g2_decap_8 FILLER_70_2343 ();
 sg13g2_decap_8 FILLER_70_2350 ();
 sg13g2_decap_8 FILLER_70_2357 ();
 sg13g2_decap_8 FILLER_70_2364 ();
 sg13g2_decap_8 FILLER_70_2371 ();
 sg13g2_decap_8 FILLER_70_2378 ();
 sg13g2_decap_8 FILLER_70_2385 ();
 sg13g2_decap_8 FILLER_70_2392 ();
 sg13g2_decap_8 FILLER_70_2399 ();
 sg13g2_decap_8 FILLER_70_2406 ();
 sg13g2_decap_8 FILLER_70_2413 ();
 sg13g2_decap_8 FILLER_70_2420 ();
 sg13g2_decap_8 FILLER_70_2427 ();
 sg13g2_decap_8 FILLER_70_2434 ();
 sg13g2_decap_8 FILLER_70_2441 ();
 sg13g2_decap_8 FILLER_70_2448 ();
 sg13g2_decap_8 FILLER_70_2455 ();
 sg13g2_decap_8 FILLER_70_2462 ();
 sg13g2_decap_8 FILLER_70_2469 ();
 sg13g2_decap_8 FILLER_70_2476 ();
 sg13g2_decap_8 FILLER_70_2483 ();
 sg13g2_decap_8 FILLER_70_2490 ();
 sg13g2_decap_8 FILLER_70_2497 ();
 sg13g2_decap_8 FILLER_70_2504 ();
 sg13g2_decap_8 FILLER_70_2511 ();
 sg13g2_decap_8 FILLER_70_2518 ();
 sg13g2_decap_8 FILLER_70_2525 ();
 sg13g2_decap_8 FILLER_70_2532 ();
 sg13g2_decap_8 FILLER_70_2539 ();
 sg13g2_decap_8 FILLER_70_2546 ();
 sg13g2_decap_8 FILLER_70_2553 ();
 sg13g2_decap_8 FILLER_70_2560 ();
 sg13g2_decap_8 FILLER_70_2567 ();
 sg13g2_decap_8 FILLER_70_2574 ();
 sg13g2_decap_8 FILLER_70_2581 ();
 sg13g2_decap_8 FILLER_70_2588 ();
 sg13g2_decap_8 FILLER_70_2595 ();
 sg13g2_decap_8 FILLER_70_2602 ();
 sg13g2_decap_8 FILLER_70_2609 ();
 sg13g2_decap_8 FILLER_70_2616 ();
 sg13g2_decap_8 FILLER_70_2623 ();
 sg13g2_decap_8 FILLER_70_2630 ();
 sg13g2_decap_8 FILLER_70_2637 ();
 sg13g2_decap_8 FILLER_70_2644 ();
 sg13g2_decap_8 FILLER_70_2651 ();
 sg13g2_decap_8 FILLER_70_2658 ();
 sg13g2_decap_8 FILLER_70_2665 ();
 sg13g2_fill_2 FILLER_70_2672 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_decap_8 FILLER_71_147 ();
 sg13g2_decap_8 FILLER_71_154 ();
 sg13g2_decap_8 FILLER_71_161 ();
 sg13g2_decap_8 FILLER_71_168 ();
 sg13g2_decap_8 FILLER_71_175 ();
 sg13g2_decap_8 FILLER_71_182 ();
 sg13g2_decap_8 FILLER_71_189 ();
 sg13g2_decap_8 FILLER_71_196 ();
 sg13g2_decap_8 FILLER_71_203 ();
 sg13g2_decap_8 FILLER_71_210 ();
 sg13g2_decap_8 FILLER_71_217 ();
 sg13g2_decap_8 FILLER_71_224 ();
 sg13g2_decap_8 FILLER_71_231 ();
 sg13g2_decap_8 FILLER_71_238 ();
 sg13g2_decap_8 FILLER_71_245 ();
 sg13g2_decap_8 FILLER_71_252 ();
 sg13g2_decap_8 FILLER_71_259 ();
 sg13g2_decap_8 FILLER_71_266 ();
 sg13g2_decap_8 FILLER_71_273 ();
 sg13g2_decap_8 FILLER_71_280 ();
 sg13g2_decap_8 FILLER_71_287 ();
 sg13g2_decap_8 FILLER_71_294 ();
 sg13g2_decap_8 FILLER_71_301 ();
 sg13g2_decap_8 FILLER_71_308 ();
 sg13g2_decap_8 FILLER_71_315 ();
 sg13g2_decap_8 FILLER_71_322 ();
 sg13g2_decap_8 FILLER_71_329 ();
 sg13g2_decap_8 FILLER_71_336 ();
 sg13g2_decap_8 FILLER_71_343 ();
 sg13g2_decap_8 FILLER_71_350 ();
 sg13g2_decap_8 FILLER_71_357 ();
 sg13g2_decap_8 FILLER_71_364 ();
 sg13g2_decap_8 FILLER_71_371 ();
 sg13g2_decap_8 FILLER_71_378 ();
 sg13g2_decap_8 FILLER_71_385 ();
 sg13g2_decap_8 FILLER_71_392 ();
 sg13g2_decap_8 FILLER_71_399 ();
 sg13g2_decap_8 FILLER_71_406 ();
 sg13g2_decap_8 FILLER_71_413 ();
 sg13g2_decap_8 FILLER_71_420 ();
 sg13g2_decap_4 FILLER_71_427 ();
 sg13g2_fill_1 FILLER_71_431 ();
 sg13g2_fill_2 FILLER_71_463 ();
 sg13g2_fill_2 FILLER_71_499 ();
 sg13g2_fill_1 FILLER_71_501 ();
 sg13g2_fill_1 FILLER_71_515 ();
 sg13g2_fill_1 FILLER_71_534 ();
 sg13g2_fill_2 FILLER_71_640 ();
 sg13g2_fill_1 FILLER_71_660 ();
 sg13g2_fill_1 FILLER_71_696 ();
 sg13g2_fill_1 FILLER_71_702 ();
 sg13g2_fill_1 FILLER_71_712 ();
 sg13g2_decap_8 FILLER_71_726 ();
 sg13g2_decap_8 FILLER_71_733 ();
 sg13g2_decap_8 FILLER_71_740 ();
 sg13g2_decap_8 FILLER_71_747 ();
 sg13g2_decap_8 FILLER_71_754 ();
 sg13g2_decap_8 FILLER_71_761 ();
 sg13g2_decap_8 FILLER_71_768 ();
 sg13g2_decap_8 FILLER_71_780 ();
 sg13g2_decap_8 FILLER_71_787 ();
 sg13g2_decap_8 FILLER_71_794 ();
 sg13g2_decap_8 FILLER_71_801 ();
 sg13g2_decap_8 FILLER_71_808 ();
 sg13g2_decap_8 FILLER_71_815 ();
 sg13g2_decap_8 FILLER_71_822 ();
 sg13g2_decap_8 FILLER_71_829 ();
 sg13g2_decap_4 FILLER_71_836 ();
 sg13g2_decap_8 FILLER_71_845 ();
 sg13g2_decap_4 FILLER_71_852 ();
 sg13g2_fill_1 FILLER_71_856 ();
 sg13g2_fill_1 FILLER_71_873 ();
 sg13g2_fill_1 FILLER_71_917 ();
 sg13g2_fill_2 FILLER_71_1046 ();
 sg13g2_fill_2 FILLER_71_1057 ();
 sg13g2_fill_1 FILLER_71_1105 ();
 sg13g2_fill_2 FILLER_71_1133 ();
 sg13g2_fill_2 FILLER_71_1304 ();
 sg13g2_fill_2 FILLER_71_1332 ();
 sg13g2_fill_2 FILLER_71_1414 ();
 sg13g2_fill_2 FILLER_71_1442 ();
 sg13g2_fill_2 FILLER_71_1486 ();
 sg13g2_fill_1 FILLER_71_1609 ();
 sg13g2_fill_1 FILLER_71_1659 ();
 sg13g2_fill_2 FILLER_71_1665 ();
 sg13g2_fill_1 FILLER_71_1667 ();
 sg13g2_fill_2 FILLER_71_1705 ();
 sg13g2_fill_1 FILLER_71_1707 ();
 sg13g2_decap_8 FILLER_71_1734 ();
 sg13g2_fill_1 FILLER_71_1792 ();
 sg13g2_decap_4 FILLER_71_1819 ();
 sg13g2_fill_1 FILLER_71_1823 ();
 sg13g2_decap_4 FILLER_71_1850 ();
 sg13g2_fill_2 FILLER_71_1854 ();
 sg13g2_fill_2 FILLER_71_1866 ();
 sg13g2_decap_4 FILLER_71_1885 ();
 sg13g2_fill_1 FILLER_71_1889 ();
 sg13g2_fill_2 FILLER_71_1899 ();
 sg13g2_fill_1 FILLER_71_1901 ();
 sg13g2_fill_1 FILLER_71_1915 ();
 sg13g2_decap_4 FILLER_71_1927 ();
 sg13g2_fill_1 FILLER_71_1931 ();
 sg13g2_fill_2 FILLER_71_1956 ();
 sg13g2_fill_2 FILLER_71_1962 ();
 sg13g2_fill_1 FILLER_71_1964 ();
 sg13g2_fill_2 FILLER_71_1973 ();
 sg13g2_fill_1 FILLER_71_1975 ();
 sg13g2_decap_4 FILLER_71_1987 ();
 sg13g2_fill_2 FILLER_71_1996 ();
 sg13g2_fill_1 FILLER_71_1998 ();
 sg13g2_fill_1 FILLER_71_2020 ();
 sg13g2_decap_4 FILLER_71_2118 ();
 sg13g2_fill_1 FILLER_71_2122 ();
 sg13g2_fill_1 FILLER_71_2138 ();
 sg13g2_decap_4 FILLER_71_2176 ();
 sg13g2_fill_2 FILLER_71_2190 ();
 sg13g2_fill_1 FILLER_71_2192 ();
 sg13g2_fill_2 FILLER_71_2206 ();
 sg13g2_fill_2 FILLER_71_2254 ();
 sg13g2_decap_8 FILLER_71_2310 ();
 sg13g2_decap_8 FILLER_71_2317 ();
 sg13g2_decap_8 FILLER_71_2324 ();
 sg13g2_decap_8 FILLER_71_2331 ();
 sg13g2_decap_8 FILLER_71_2338 ();
 sg13g2_decap_8 FILLER_71_2345 ();
 sg13g2_decap_8 FILLER_71_2352 ();
 sg13g2_decap_8 FILLER_71_2359 ();
 sg13g2_decap_8 FILLER_71_2366 ();
 sg13g2_decap_8 FILLER_71_2373 ();
 sg13g2_decap_8 FILLER_71_2380 ();
 sg13g2_decap_8 FILLER_71_2387 ();
 sg13g2_decap_8 FILLER_71_2394 ();
 sg13g2_decap_8 FILLER_71_2401 ();
 sg13g2_decap_8 FILLER_71_2408 ();
 sg13g2_decap_8 FILLER_71_2415 ();
 sg13g2_decap_8 FILLER_71_2422 ();
 sg13g2_decap_8 FILLER_71_2429 ();
 sg13g2_decap_8 FILLER_71_2436 ();
 sg13g2_decap_8 FILLER_71_2443 ();
 sg13g2_decap_8 FILLER_71_2450 ();
 sg13g2_decap_8 FILLER_71_2457 ();
 sg13g2_decap_8 FILLER_71_2464 ();
 sg13g2_decap_8 FILLER_71_2471 ();
 sg13g2_decap_8 FILLER_71_2478 ();
 sg13g2_decap_8 FILLER_71_2485 ();
 sg13g2_decap_8 FILLER_71_2492 ();
 sg13g2_decap_8 FILLER_71_2499 ();
 sg13g2_decap_8 FILLER_71_2506 ();
 sg13g2_decap_8 FILLER_71_2513 ();
 sg13g2_decap_8 FILLER_71_2520 ();
 sg13g2_decap_8 FILLER_71_2527 ();
 sg13g2_decap_8 FILLER_71_2534 ();
 sg13g2_decap_8 FILLER_71_2541 ();
 sg13g2_decap_8 FILLER_71_2548 ();
 sg13g2_decap_8 FILLER_71_2555 ();
 sg13g2_decap_8 FILLER_71_2562 ();
 sg13g2_decap_8 FILLER_71_2569 ();
 sg13g2_decap_8 FILLER_71_2576 ();
 sg13g2_decap_8 FILLER_71_2583 ();
 sg13g2_decap_8 FILLER_71_2590 ();
 sg13g2_decap_8 FILLER_71_2597 ();
 sg13g2_decap_8 FILLER_71_2604 ();
 sg13g2_decap_8 FILLER_71_2611 ();
 sg13g2_decap_8 FILLER_71_2618 ();
 sg13g2_decap_8 FILLER_71_2625 ();
 sg13g2_decap_8 FILLER_71_2632 ();
 sg13g2_decap_8 FILLER_71_2639 ();
 sg13g2_decap_8 FILLER_71_2646 ();
 sg13g2_decap_8 FILLER_71_2653 ();
 sg13g2_decap_8 FILLER_71_2660 ();
 sg13g2_decap_8 FILLER_71_2667 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_decap_8 FILLER_72_161 ();
 sg13g2_decap_8 FILLER_72_168 ();
 sg13g2_decap_8 FILLER_72_175 ();
 sg13g2_decap_8 FILLER_72_182 ();
 sg13g2_decap_8 FILLER_72_189 ();
 sg13g2_decap_8 FILLER_72_196 ();
 sg13g2_decap_8 FILLER_72_203 ();
 sg13g2_decap_8 FILLER_72_210 ();
 sg13g2_decap_8 FILLER_72_217 ();
 sg13g2_decap_8 FILLER_72_224 ();
 sg13g2_decap_8 FILLER_72_231 ();
 sg13g2_decap_8 FILLER_72_238 ();
 sg13g2_decap_8 FILLER_72_245 ();
 sg13g2_decap_8 FILLER_72_252 ();
 sg13g2_decap_8 FILLER_72_259 ();
 sg13g2_decap_8 FILLER_72_266 ();
 sg13g2_decap_8 FILLER_72_273 ();
 sg13g2_decap_8 FILLER_72_280 ();
 sg13g2_decap_8 FILLER_72_287 ();
 sg13g2_decap_8 FILLER_72_294 ();
 sg13g2_decap_8 FILLER_72_301 ();
 sg13g2_decap_8 FILLER_72_308 ();
 sg13g2_decap_8 FILLER_72_315 ();
 sg13g2_decap_8 FILLER_72_322 ();
 sg13g2_decap_8 FILLER_72_329 ();
 sg13g2_decap_8 FILLER_72_336 ();
 sg13g2_decap_8 FILLER_72_343 ();
 sg13g2_decap_8 FILLER_72_350 ();
 sg13g2_decap_8 FILLER_72_357 ();
 sg13g2_decap_8 FILLER_72_364 ();
 sg13g2_decap_8 FILLER_72_371 ();
 sg13g2_decap_8 FILLER_72_378 ();
 sg13g2_decap_8 FILLER_72_385 ();
 sg13g2_decap_8 FILLER_72_392 ();
 sg13g2_decap_8 FILLER_72_399 ();
 sg13g2_decap_8 FILLER_72_406 ();
 sg13g2_decap_8 FILLER_72_413 ();
 sg13g2_decap_8 FILLER_72_420 ();
 sg13g2_decap_8 FILLER_72_427 ();
 sg13g2_fill_2 FILLER_72_434 ();
 sg13g2_fill_2 FILLER_72_484 ();
 sg13g2_fill_1 FILLER_72_486 ();
 sg13g2_fill_2 FILLER_72_536 ();
 sg13g2_fill_1 FILLER_72_551 ();
 sg13g2_fill_2 FILLER_72_586 ();
 sg13g2_fill_1 FILLER_72_588 ();
 sg13g2_fill_1 FILLER_72_597 ();
 sg13g2_fill_2 FILLER_72_658 ();
 sg13g2_fill_1 FILLER_72_679 ();
 sg13g2_decap_8 FILLER_72_720 ();
 sg13g2_decap_8 FILLER_72_727 ();
 sg13g2_decap_8 FILLER_72_734 ();
 sg13g2_decap_8 FILLER_72_741 ();
 sg13g2_decap_8 FILLER_72_748 ();
 sg13g2_decap_8 FILLER_72_755 ();
 sg13g2_decap_8 FILLER_72_762 ();
 sg13g2_decap_8 FILLER_72_769 ();
 sg13g2_decap_8 FILLER_72_776 ();
 sg13g2_decap_8 FILLER_72_783 ();
 sg13g2_decap_8 FILLER_72_790 ();
 sg13g2_decap_8 FILLER_72_797 ();
 sg13g2_decap_8 FILLER_72_804 ();
 sg13g2_decap_8 FILLER_72_811 ();
 sg13g2_decap_8 FILLER_72_818 ();
 sg13g2_decap_8 FILLER_72_825 ();
 sg13g2_decap_8 FILLER_72_832 ();
 sg13g2_decap_8 FILLER_72_839 ();
 sg13g2_decap_8 FILLER_72_846 ();
 sg13g2_decap_8 FILLER_72_853 ();
 sg13g2_fill_1 FILLER_72_860 ();
 sg13g2_fill_1 FILLER_72_865 ();
 sg13g2_fill_2 FILLER_72_882 ();
 sg13g2_fill_1 FILLER_72_884 ();
 sg13g2_fill_1 FILLER_72_939 ();
 sg13g2_fill_2 FILLER_72_1014 ();
 sg13g2_fill_1 FILLER_72_1081 ();
 sg13g2_fill_1 FILLER_72_1172 ();
 sg13g2_fill_2 FILLER_72_1246 ();
 sg13g2_fill_1 FILLER_72_1351 ();
 sg13g2_fill_2 FILLER_72_1443 ();
 sg13g2_fill_1 FILLER_72_1524 ();
 sg13g2_fill_1 FILLER_72_1619 ();
 sg13g2_fill_1 FILLER_72_1643 ();
 sg13g2_fill_1 FILLER_72_1695 ();
 sg13g2_fill_2 FILLER_72_1724 ();
 sg13g2_fill_2 FILLER_72_1786 ();
 sg13g2_fill_2 FILLER_72_1815 ();
 sg13g2_fill_2 FILLER_72_1972 ();
 sg13g2_decap_8 FILLER_72_2013 ();
 sg13g2_fill_1 FILLER_72_2069 ();
 sg13g2_fill_1 FILLER_72_2106 ();
 sg13g2_decap_8 FILLER_72_2136 ();
 sg13g2_fill_2 FILLER_72_2152 ();
 sg13g2_fill_1 FILLER_72_2154 ();
 sg13g2_fill_2 FILLER_72_2182 ();
 sg13g2_decap_4 FILLER_72_2210 ();
 sg13g2_fill_2 FILLER_72_2214 ();
 sg13g2_fill_1 FILLER_72_2246 ();
 sg13g2_fill_1 FILLER_72_2281 ();
 sg13g2_decap_8 FILLER_72_2308 ();
 sg13g2_decap_8 FILLER_72_2315 ();
 sg13g2_decap_8 FILLER_72_2322 ();
 sg13g2_decap_8 FILLER_72_2329 ();
 sg13g2_decap_8 FILLER_72_2336 ();
 sg13g2_decap_8 FILLER_72_2343 ();
 sg13g2_decap_8 FILLER_72_2350 ();
 sg13g2_decap_8 FILLER_72_2357 ();
 sg13g2_decap_8 FILLER_72_2364 ();
 sg13g2_decap_8 FILLER_72_2371 ();
 sg13g2_decap_8 FILLER_72_2378 ();
 sg13g2_decap_8 FILLER_72_2385 ();
 sg13g2_decap_8 FILLER_72_2392 ();
 sg13g2_decap_8 FILLER_72_2399 ();
 sg13g2_decap_8 FILLER_72_2406 ();
 sg13g2_decap_8 FILLER_72_2413 ();
 sg13g2_decap_8 FILLER_72_2420 ();
 sg13g2_decap_8 FILLER_72_2427 ();
 sg13g2_decap_8 FILLER_72_2434 ();
 sg13g2_decap_8 FILLER_72_2441 ();
 sg13g2_decap_8 FILLER_72_2448 ();
 sg13g2_decap_8 FILLER_72_2455 ();
 sg13g2_decap_8 FILLER_72_2462 ();
 sg13g2_decap_8 FILLER_72_2469 ();
 sg13g2_decap_8 FILLER_72_2476 ();
 sg13g2_decap_8 FILLER_72_2483 ();
 sg13g2_decap_8 FILLER_72_2490 ();
 sg13g2_decap_8 FILLER_72_2497 ();
 sg13g2_decap_8 FILLER_72_2504 ();
 sg13g2_decap_8 FILLER_72_2511 ();
 sg13g2_decap_8 FILLER_72_2518 ();
 sg13g2_decap_8 FILLER_72_2525 ();
 sg13g2_decap_8 FILLER_72_2532 ();
 sg13g2_decap_8 FILLER_72_2539 ();
 sg13g2_decap_8 FILLER_72_2546 ();
 sg13g2_decap_8 FILLER_72_2553 ();
 sg13g2_decap_8 FILLER_72_2560 ();
 sg13g2_decap_8 FILLER_72_2567 ();
 sg13g2_decap_8 FILLER_72_2574 ();
 sg13g2_decap_8 FILLER_72_2581 ();
 sg13g2_decap_8 FILLER_72_2588 ();
 sg13g2_decap_8 FILLER_72_2595 ();
 sg13g2_decap_8 FILLER_72_2602 ();
 sg13g2_decap_8 FILLER_72_2609 ();
 sg13g2_decap_8 FILLER_72_2616 ();
 sg13g2_decap_8 FILLER_72_2623 ();
 sg13g2_decap_8 FILLER_72_2630 ();
 sg13g2_decap_8 FILLER_72_2637 ();
 sg13g2_decap_8 FILLER_72_2644 ();
 sg13g2_decap_8 FILLER_72_2651 ();
 sg13g2_decap_8 FILLER_72_2658 ();
 sg13g2_decap_8 FILLER_72_2665 ();
 sg13g2_fill_2 FILLER_72_2672 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_decap_8 FILLER_73_168 ();
 sg13g2_decap_8 FILLER_73_175 ();
 sg13g2_decap_8 FILLER_73_182 ();
 sg13g2_decap_8 FILLER_73_189 ();
 sg13g2_decap_8 FILLER_73_196 ();
 sg13g2_decap_8 FILLER_73_203 ();
 sg13g2_decap_8 FILLER_73_210 ();
 sg13g2_decap_8 FILLER_73_217 ();
 sg13g2_decap_8 FILLER_73_224 ();
 sg13g2_decap_8 FILLER_73_231 ();
 sg13g2_decap_8 FILLER_73_238 ();
 sg13g2_decap_8 FILLER_73_245 ();
 sg13g2_decap_8 FILLER_73_252 ();
 sg13g2_decap_8 FILLER_73_259 ();
 sg13g2_decap_8 FILLER_73_266 ();
 sg13g2_decap_8 FILLER_73_273 ();
 sg13g2_decap_8 FILLER_73_280 ();
 sg13g2_decap_8 FILLER_73_287 ();
 sg13g2_decap_8 FILLER_73_294 ();
 sg13g2_decap_8 FILLER_73_301 ();
 sg13g2_decap_8 FILLER_73_308 ();
 sg13g2_decap_8 FILLER_73_315 ();
 sg13g2_decap_8 FILLER_73_322 ();
 sg13g2_decap_8 FILLER_73_329 ();
 sg13g2_decap_8 FILLER_73_336 ();
 sg13g2_decap_8 FILLER_73_343 ();
 sg13g2_decap_8 FILLER_73_350 ();
 sg13g2_decap_8 FILLER_73_357 ();
 sg13g2_decap_8 FILLER_73_364 ();
 sg13g2_decap_8 FILLER_73_371 ();
 sg13g2_decap_8 FILLER_73_378 ();
 sg13g2_decap_8 FILLER_73_385 ();
 sg13g2_decap_8 FILLER_73_392 ();
 sg13g2_decap_8 FILLER_73_399 ();
 sg13g2_decap_8 FILLER_73_406 ();
 sg13g2_decap_8 FILLER_73_413 ();
 sg13g2_decap_8 FILLER_73_420 ();
 sg13g2_decap_8 FILLER_73_427 ();
 sg13g2_decap_4 FILLER_73_434 ();
 sg13g2_fill_2 FILLER_73_486 ();
 sg13g2_fill_1 FILLER_73_497 ();
 sg13g2_fill_2 FILLER_73_577 ();
 sg13g2_fill_2 FILLER_73_627 ();
 sg13g2_fill_2 FILLER_73_686 ();
 sg13g2_decap_4 FILLER_73_711 ();
 sg13g2_decap_8 FILLER_73_725 ();
 sg13g2_decap_8 FILLER_73_732 ();
 sg13g2_decap_8 FILLER_73_739 ();
 sg13g2_decap_8 FILLER_73_746 ();
 sg13g2_decap_8 FILLER_73_753 ();
 sg13g2_decap_8 FILLER_73_760 ();
 sg13g2_decap_8 FILLER_73_767 ();
 sg13g2_decap_8 FILLER_73_774 ();
 sg13g2_decap_8 FILLER_73_781 ();
 sg13g2_decap_8 FILLER_73_788 ();
 sg13g2_decap_8 FILLER_73_795 ();
 sg13g2_decap_8 FILLER_73_802 ();
 sg13g2_decap_8 FILLER_73_809 ();
 sg13g2_decap_8 FILLER_73_816 ();
 sg13g2_decap_8 FILLER_73_823 ();
 sg13g2_decap_8 FILLER_73_830 ();
 sg13g2_decap_8 FILLER_73_837 ();
 sg13g2_decap_8 FILLER_73_844 ();
 sg13g2_decap_8 FILLER_73_851 ();
 sg13g2_decap_8 FILLER_73_858 ();
 sg13g2_fill_1 FILLER_73_865 ();
 sg13g2_fill_2 FILLER_73_944 ();
 sg13g2_fill_1 FILLER_73_985 ();
 sg13g2_fill_2 FILLER_73_1020 ();
 sg13g2_fill_2 FILLER_73_1080 ();
 sg13g2_fill_1 FILLER_73_1100 ();
 sg13g2_fill_2 FILLER_73_1132 ();
 sg13g2_fill_1 FILLER_73_1153 ();
 sg13g2_fill_1 FILLER_73_1159 ();
 sg13g2_fill_2 FILLER_73_1223 ();
 sg13g2_fill_1 FILLER_73_1247 ();
 sg13g2_fill_1 FILLER_73_1346 ();
 sg13g2_fill_1 FILLER_73_1362 ();
 sg13g2_fill_2 FILLER_73_1443 ();
 sg13g2_fill_2 FILLER_73_1471 ();
 sg13g2_fill_1 FILLER_73_1508 ();
 sg13g2_decap_4 FILLER_73_1547 ();
 sg13g2_fill_1 FILLER_73_1654 ();
 sg13g2_fill_2 FILLER_73_1659 ();
 sg13g2_fill_2 FILLER_73_1686 ();
 sg13g2_fill_1 FILLER_73_1688 ();
 sg13g2_fill_2 FILLER_73_1694 ();
 sg13g2_fill_2 FILLER_73_1722 ();
 sg13g2_fill_1 FILLER_73_1724 ();
 sg13g2_decap_4 FILLER_73_1742 ();
 sg13g2_fill_2 FILLER_73_1760 ();
 sg13g2_fill_1 FILLER_73_1787 ();
 sg13g2_fill_2 FILLER_73_1802 ();
 sg13g2_fill_1 FILLER_73_1804 ();
 sg13g2_decap_8 FILLER_73_1869 ();
 sg13g2_decap_4 FILLER_73_1910 ();
 sg13g2_fill_1 FILLER_73_1914 ();
 sg13g2_fill_1 FILLER_73_1931 ();
 sg13g2_decap_4 FILLER_73_1956 ();
 sg13g2_decap_4 FILLER_73_1968 ();
 sg13g2_fill_2 FILLER_73_1986 ();
 sg13g2_fill_1 FILLER_73_1988 ();
 sg13g2_fill_1 FILLER_73_1999 ();
 sg13g2_fill_2 FILLER_73_2029 ();
 sg13g2_fill_1 FILLER_73_2035 ();
 sg13g2_decap_4 FILLER_73_2072 ();
 sg13g2_decap_4 FILLER_73_2080 ();
 sg13g2_fill_2 FILLER_73_2084 ();
 sg13g2_fill_2 FILLER_73_2114 ();
 sg13g2_fill_1 FILLER_73_2116 ();
 sg13g2_fill_1 FILLER_73_2142 ();
 sg13g2_fill_1 FILLER_73_2161 ();
 sg13g2_fill_1 FILLER_73_2171 ();
 sg13g2_fill_2 FILLER_73_2245 ();
 sg13g2_fill_1 FILLER_73_2247 ();
 sg13g2_fill_2 FILLER_73_2258 ();
 sg13g2_fill_1 FILLER_73_2260 ();
 sg13g2_decap_8 FILLER_73_2301 ();
 sg13g2_decap_8 FILLER_73_2308 ();
 sg13g2_decap_8 FILLER_73_2315 ();
 sg13g2_decap_8 FILLER_73_2322 ();
 sg13g2_decap_8 FILLER_73_2329 ();
 sg13g2_decap_8 FILLER_73_2336 ();
 sg13g2_decap_8 FILLER_73_2343 ();
 sg13g2_decap_8 FILLER_73_2350 ();
 sg13g2_decap_8 FILLER_73_2357 ();
 sg13g2_decap_8 FILLER_73_2364 ();
 sg13g2_decap_8 FILLER_73_2371 ();
 sg13g2_decap_8 FILLER_73_2378 ();
 sg13g2_decap_8 FILLER_73_2385 ();
 sg13g2_decap_8 FILLER_73_2392 ();
 sg13g2_decap_8 FILLER_73_2399 ();
 sg13g2_decap_8 FILLER_73_2406 ();
 sg13g2_decap_8 FILLER_73_2413 ();
 sg13g2_decap_8 FILLER_73_2420 ();
 sg13g2_decap_8 FILLER_73_2427 ();
 sg13g2_decap_8 FILLER_73_2434 ();
 sg13g2_decap_8 FILLER_73_2441 ();
 sg13g2_decap_8 FILLER_73_2448 ();
 sg13g2_decap_8 FILLER_73_2455 ();
 sg13g2_decap_8 FILLER_73_2462 ();
 sg13g2_decap_8 FILLER_73_2469 ();
 sg13g2_decap_8 FILLER_73_2476 ();
 sg13g2_decap_8 FILLER_73_2483 ();
 sg13g2_decap_8 FILLER_73_2490 ();
 sg13g2_decap_8 FILLER_73_2497 ();
 sg13g2_decap_8 FILLER_73_2504 ();
 sg13g2_decap_8 FILLER_73_2511 ();
 sg13g2_decap_8 FILLER_73_2518 ();
 sg13g2_decap_8 FILLER_73_2525 ();
 sg13g2_decap_8 FILLER_73_2532 ();
 sg13g2_decap_8 FILLER_73_2539 ();
 sg13g2_decap_8 FILLER_73_2546 ();
 sg13g2_decap_8 FILLER_73_2553 ();
 sg13g2_decap_8 FILLER_73_2560 ();
 sg13g2_decap_8 FILLER_73_2567 ();
 sg13g2_decap_8 FILLER_73_2574 ();
 sg13g2_decap_8 FILLER_73_2581 ();
 sg13g2_decap_8 FILLER_73_2588 ();
 sg13g2_decap_8 FILLER_73_2595 ();
 sg13g2_decap_8 FILLER_73_2602 ();
 sg13g2_decap_8 FILLER_73_2609 ();
 sg13g2_decap_8 FILLER_73_2616 ();
 sg13g2_decap_8 FILLER_73_2623 ();
 sg13g2_decap_8 FILLER_73_2630 ();
 sg13g2_decap_8 FILLER_73_2637 ();
 sg13g2_decap_8 FILLER_73_2644 ();
 sg13g2_decap_8 FILLER_73_2651 ();
 sg13g2_decap_8 FILLER_73_2658 ();
 sg13g2_decap_8 FILLER_73_2665 ();
 sg13g2_fill_2 FILLER_73_2672 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_168 ();
 sg13g2_decap_8 FILLER_74_175 ();
 sg13g2_decap_8 FILLER_74_182 ();
 sg13g2_decap_8 FILLER_74_189 ();
 sg13g2_decap_8 FILLER_74_196 ();
 sg13g2_decap_8 FILLER_74_203 ();
 sg13g2_decap_8 FILLER_74_210 ();
 sg13g2_decap_8 FILLER_74_217 ();
 sg13g2_decap_8 FILLER_74_224 ();
 sg13g2_decap_8 FILLER_74_231 ();
 sg13g2_decap_8 FILLER_74_238 ();
 sg13g2_decap_8 FILLER_74_245 ();
 sg13g2_decap_8 FILLER_74_252 ();
 sg13g2_decap_8 FILLER_74_259 ();
 sg13g2_decap_8 FILLER_74_266 ();
 sg13g2_decap_8 FILLER_74_273 ();
 sg13g2_decap_8 FILLER_74_280 ();
 sg13g2_decap_8 FILLER_74_287 ();
 sg13g2_decap_8 FILLER_74_294 ();
 sg13g2_decap_8 FILLER_74_301 ();
 sg13g2_decap_8 FILLER_74_308 ();
 sg13g2_decap_8 FILLER_74_315 ();
 sg13g2_decap_8 FILLER_74_322 ();
 sg13g2_decap_8 FILLER_74_329 ();
 sg13g2_decap_8 FILLER_74_336 ();
 sg13g2_decap_8 FILLER_74_343 ();
 sg13g2_decap_8 FILLER_74_350 ();
 sg13g2_decap_8 FILLER_74_357 ();
 sg13g2_decap_8 FILLER_74_364 ();
 sg13g2_decap_8 FILLER_74_371 ();
 sg13g2_decap_8 FILLER_74_378 ();
 sg13g2_decap_8 FILLER_74_385 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_decap_8 FILLER_74_399 ();
 sg13g2_decap_8 FILLER_74_406 ();
 sg13g2_decap_8 FILLER_74_413 ();
 sg13g2_decap_8 FILLER_74_420 ();
 sg13g2_decap_8 FILLER_74_427 ();
 sg13g2_decap_8 FILLER_74_434 ();
 sg13g2_decap_4 FILLER_74_441 ();
 sg13g2_fill_1 FILLER_74_445 ();
 sg13g2_fill_2 FILLER_74_525 ();
 sg13g2_fill_1 FILLER_74_671 ();
 sg13g2_fill_2 FILLER_74_689 ();
 sg13g2_decap_8 FILLER_74_717 ();
 sg13g2_decap_8 FILLER_74_724 ();
 sg13g2_decap_8 FILLER_74_731 ();
 sg13g2_decap_8 FILLER_74_738 ();
 sg13g2_decap_8 FILLER_74_745 ();
 sg13g2_decap_8 FILLER_74_752 ();
 sg13g2_decap_8 FILLER_74_759 ();
 sg13g2_decap_8 FILLER_74_766 ();
 sg13g2_decap_8 FILLER_74_773 ();
 sg13g2_decap_8 FILLER_74_780 ();
 sg13g2_decap_8 FILLER_74_787 ();
 sg13g2_decap_8 FILLER_74_794 ();
 sg13g2_decap_8 FILLER_74_801 ();
 sg13g2_decap_8 FILLER_74_808 ();
 sg13g2_decap_8 FILLER_74_815 ();
 sg13g2_decap_8 FILLER_74_822 ();
 sg13g2_decap_8 FILLER_74_829 ();
 sg13g2_decap_8 FILLER_74_836 ();
 sg13g2_decap_8 FILLER_74_843 ();
 sg13g2_decap_8 FILLER_74_850 ();
 sg13g2_decap_8 FILLER_74_857 ();
 sg13g2_decap_8 FILLER_74_864 ();
 sg13g2_decap_8 FILLER_74_871 ();
 sg13g2_decap_8 FILLER_74_878 ();
 sg13g2_decap_8 FILLER_74_885 ();
 sg13g2_decap_8 FILLER_74_892 ();
 sg13g2_fill_2 FILLER_74_899 ();
 sg13g2_fill_1 FILLER_74_901 ();
 sg13g2_fill_2 FILLER_74_911 ();
 sg13g2_fill_2 FILLER_74_1153 ();
 sg13g2_fill_1 FILLER_74_1301 ();
 sg13g2_fill_1 FILLER_74_1415 ();
 sg13g2_fill_2 FILLER_74_1466 ();
 sg13g2_fill_2 FILLER_74_1524 ();
 sg13g2_decap_8 FILLER_74_1562 ();
 sg13g2_fill_1 FILLER_74_1588 ();
 sg13g2_fill_2 FILLER_74_1704 ();
 sg13g2_fill_1 FILLER_74_1706 ();
 sg13g2_decap_4 FILLER_74_1747 ();
 sg13g2_fill_2 FILLER_74_1751 ();
 sg13g2_fill_2 FILLER_74_1810 ();
 sg13g2_fill_1 FILLER_74_1812 ();
 sg13g2_fill_2 FILLER_74_1841 ();
 sg13g2_fill_2 FILLER_74_1869 ();
 sg13g2_fill_1 FILLER_74_1871 ();
 sg13g2_decap_8 FILLER_74_1904 ();
 sg13g2_decap_4 FILLER_74_1911 ();
 sg13g2_fill_2 FILLER_74_1932 ();
 sg13g2_fill_1 FILLER_74_1956 ();
 sg13g2_decap_4 FILLER_74_1971 ();
 sg13g2_fill_1 FILLER_74_1986 ();
 sg13g2_fill_1 FILLER_74_2016 ();
 sg13g2_fill_1 FILLER_74_2043 ();
 sg13g2_decap_4 FILLER_74_2053 ();
 sg13g2_decap_4 FILLER_74_2061 ();
 sg13g2_fill_1 FILLER_74_2065 ();
 sg13g2_fill_2 FILLER_74_2199 ();
 sg13g2_fill_1 FILLER_74_2201 ();
 sg13g2_fill_1 FILLER_74_2238 ();
 sg13g2_decap_8 FILLER_74_2274 ();
 sg13g2_decap_8 FILLER_74_2294 ();
 sg13g2_decap_8 FILLER_74_2301 ();
 sg13g2_decap_8 FILLER_74_2308 ();
 sg13g2_decap_8 FILLER_74_2315 ();
 sg13g2_decap_8 FILLER_74_2322 ();
 sg13g2_decap_8 FILLER_74_2329 ();
 sg13g2_decap_8 FILLER_74_2336 ();
 sg13g2_decap_8 FILLER_74_2343 ();
 sg13g2_decap_8 FILLER_74_2350 ();
 sg13g2_decap_8 FILLER_74_2357 ();
 sg13g2_decap_8 FILLER_74_2364 ();
 sg13g2_decap_8 FILLER_74_2371 ();
 sg13g2_decap_8 FILLER_74_2378 ();
 sg13g2_decap_8 FILLER_74_2385 ();
 sg13g2_decap_8 FILLER_74_2392 ();
 sg13g2_decap_8 FILLER_74_2399 ();
 sg13g2_decap_8 FILLER_74_2406 ();
 sg13g2_decap_8 FILLER_74_2413 ();
 sg13g2_decap_8 FILLER_74_2420 ();
 sg13g2_decap_8 FILLER_74_2427 ();
 sg13g2_decap_8 FILLER_74_2434 ();
 sg13g2_decap_8 FILLER_74_2441 ();
 sg13g2_decap_8 FILLER_74_2448 ();
 sg13g2_decap_8 FILLER_74_2455 ();
 sg13g2_decap_8 FILLER_74_2462 ();
 sg13g2_decap_8 FILLER_74_2469 ();
 sg13g2_decap_8 FILLER_74_2476 ();
 sg13g2_decap_8 FILLER_74_2483 ();
 sg13g2_decap_8 FILLER_74_2490 ();
 sg13g2_decap_8 FILLER_74_2497 ();
 sg13g2_decap_8 FILLER_74_2504 ();
 sg13g2_decap_8 FILLER_74_2511 ();
 sg13g2_decap_8 FILLER_74_2518 ();
 sg13g2_decap_8 FILLER_74_2525 ();
 sg13g2_decap_8 FILLER_74_2532 ();
 sg13g2_decap_8 FILLER_74_2539 ();
 sg13g2_decap_8 FILLER_74_2546 ();
 sg13g2_decap_8 FILLER_74_2553 ();
 sg13g2_decap_8 FILLER_74_2560 ();
 sg13g2_decap_8 FILLER_74_2567 ();
 sg13g2_decap_8 FILLER_74_2574 ();
 sg13g2_decap_8 FILLER_74_2581 ();
 sg13g2_decap_8 FILLER_74_2588 ();
 sg13g2_decap_8 FILLER_74_2595 ();
 sg13g2_decap_8 FILLER_74_2602 ();
 sg13g2_decap_8 FILLER_74_2609 ();
 sg13g2_decap_8 FILLER_74_2616 ();
 sg13g2_decap_8 FILLER_74_2623 ();
 sg13g2_decap_8 FILLER_74_2630 ();
 sg13g2_decap_8 FILLER_74_2637 ();
 sg13g2_decap_8 FILLER_74_2644 ();
 sg13g2_decap_8 FILLER_74_2651 ();
 sg13g2_decap_8 FILLER_74_2658 ();
 sg13g2_decap_8 FILLER_74_2665 ();
 sg13g2_fill_2 FILLER_74_2672 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_8 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_182 ();
 sg13g2_decap_8 FILLER_75_189 ();
 sg13g2_decap_8 FILLER_75_196 ();
 sg13g2_decap_8 FILLER_75_203 ();
 sg13g2_decap_8 FILLER_75_210 ();
 sg13g2_decap_8 FILLER_75_217 ();
 sg13g2_decap_8 FILLER_75_224 ();
 sg13g2_decap_8 FILLER_75_231 ();
 sg13g2_decap_8 FILLER_75_238 ();
 sg13g2_decap_8 FILLER_75_245 ();
 sg13g2_decap_8 FILLER_75_252 ();
 sg13g2_decap_8 FILLER_75_259 ();
 sg13g2_decap_8 FILLER_75_266 ();
 sg13g2_decap_8 FILLER_75_273 ();
 sg13g2_decap_8 FILLER_75_280 ();
 sg13g2_decap_8 FILLER_75_287 ();
 sg13g2_decap_8 FILLER_75_294 ();
 sg13g2_decap_8 FILLER_75_301 ();
 sg13g2_decap_8 FILLER_75_308 ();
 sg13g2_decap_8 FILLER_75_315 ();
 sg13g2_decap_8 FILLER_75_322 ();
 sg13g2_decap_8 FILLER_75_329 ();
 sg13g2_decap_8 FILLER_75_336 ();
 sg13g2_decap_8 FILLER_75_343 ();
 sg13g2_decap_8 FILLER_75_350 ();
 sg13g2_decap_8 FILLER_75_357 ();
 sg13g2_decap_8 FILLER_75_364 ();
 sg13g2_decap_8 FILLER_75_371 ();
 sg13g2_decap_8 FILLER_75_378 ();
 sg13g2_decap_8 FILLER_75_385 ();
 sg13g2_decap_8 FILLER_75_392 ();
 sg13g2_decap_8 FILLER_75_399 ();
 sg13g2_decap_8 FILLER_75_406 ();
 sg13g2_decap_8 FILLER_75_413 ();
 sg13g2_decap_8 FILLER_75_420 ();
 sg13g2_decap_8 FILLER_75_427 ();
 sg13g2_decap_8 FILLER_75_434 ();
 sg13g2_decap_8 FILLER_75_441 ();
 sg13g2_fill_2 FILLER_75_448 ();
 sg13g2_fill_2 FILLER_75_453 ();
 sg13g2_fill_2 FILLER_75_552 ();
 sg13g2_fill_1 FILLER_75_554 ();
 sg13g2_fill_1 FILLER_75_562 ();
 sg13g2_decap_4 FILLER_75_647 ();
 sg13g2_fill_1 FILLER_75_683 ();
 sg13g2_decap_8 FILLER_75_707 ();
 sg13g2_decap_8 FILLER_75_714 ();
 sg13g2_decap_8 FILLER_75_721 ();
 sg13g2_decap_8 FILLER_75_728 ();
 sg13g2_decap_8 FILLER_75_735 ();
 sg13g2_decap_8 FILLER_75_742 ();
 sg13g2_decap_8 FILLER_75_749 ();
 sg13g2_decap_8 FILLER_75_756 ();
 sg13g2_decap_8 FILLER_75_763 ();
 sg13g2_decap_8 FILLER_75_770 ();
 sg13g2_decap_8 FILLER_75_777 ();
 sg13g2_decap_8 FILLER_75_784 ();
 sg13g2_decap_8 FILLER_75_791 ();
 sg13g2_decap_8 FILLER_75_798 ();
 sg13g2_decap_8 FILLER_75_805 ();
 sg13g2_decap_8 FILLER_75_812 ();
 sg13g2_decap_8 FILLER_75_819 ();
 sg13g2_decap_8 FILLER_75_826 ();
 sg13g2_decap_8 FILLER_75_833 ();
 sg13g2_decap_8 FILLER_75_840 ();
 sg13g2_decap_8 FILLER_75_847 ();
 sg13g2_decap_8 FILLER_75_854 ();
 sg13g2_decap_8 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_75_868 ();
 sg13g2_decap_8 FILLER_75_875 ();
 sg13g2_decap_8 FILLER_75_882 ();
 sg13g2_decap_8 FILLER_75_889 ();
 sg13g2_decap_8 FILLER_75_896 ();
 sg13g2_decap_8 FILLER_75_903 ();
 sg13g2_decap_8 FILLER_75_910 ();
 sg13g2_fill_2 FILLER_75_917 ();
 sg13g2_fill_1 FILLER_75_919 ();
 sg13g2_fill_1 FILLER_75_933 ();
 sg13g2_fill_1 FILLER_75_957 ();
 sg13g2_fill_1 FILLER_75_987 ();
 sg13g2_fill_1 FILLER_75_1042 ();
 sg13g2_fill_1 FILLER_75_1187 ();
 sg13g2_fill_1 FILLER_75_1287 ();
 sg13g2_fill_1 FILLER_75_1357 ();
 sg13g2_fill_1 FILLER_75_1376 ();
 sg13g2_fill_1 FILLER_75_1394 ();
 sg13g2_fill_2 FILLER_75_1481 ();
 sg13g2_fill_1 FILLER_75_1509 ();
 sg13g2_fill_1 FILLER_75_1583 ();
 sg13g2_fill_2 FILLER_75_1597 ();
 sg13g2_fill_2 FILLER_75_1604 ();
 sg13g2_fill_1 FILLER_75_1632 ();
 sg13g2_fill_1 FILLER_75_1647 ();
 sg13g2_fill_2 FILLER_75_1657 ();
 sg13g2_fill_1 FILLER_75_1659 ();
 sg13g2_fill_1 FILLER_75_1695 ();
 sg13g2_fill_2 FILLER_75_1705 ();
 sg13g2_fill_1 FILLER_75_1731 ();
 sg13g2_fill_1 FILLER_75_1767 ();
 sg13g2_fill_2 FILLER_75_1795 ();
 sg13g2_fill_2 FILLER_75_1851 ();
 sg13g2_fill_1 FILLER_75_1853 ();
 sg13g2_decap_4 FILLER_75_1912 ();
 sg13g2_decap_4 FILLER_75_2072 ();
 sg13g2_fill_1 FILLER_75_2076 ();
 sg13g2_fill_2 FILLER_75_2086 ();
 sg13g2_fill_1 FILLER_75_2088 ();
 sg13g2_fill_2 FILLER_75_2103 ();
 sg13g2_fill_1 FILLER_75_2105 ();
 sg13g2_fill_1 FILLER_75_2115 ();
 sg13g2_decap_8 FILLER_75_2145 ();
 sg13g2_fill_2 FILLER_75_2175 ();
 sg13g2_decap_8 FILLER_75_2213 ();
 sg13g2_fill_2 FILLER_75_2220 ();
 sg13g2_fill_1 FILLER_75_2236 ();
 sg13g2_fill_2 FILLER_75_2251 ();
 sg13g2_fill_1 FILLER_75_2253 ();
 sg13g2_decap_8 FILLER_75_2290 ();
 sg13g2_decap_8 FILLER_75_2297 ();
 sg13g2_decap_8 FILLER_75_2304 ();
 sg13g2_decap_8 FILLER_75_2311 ();
 sg13g2_decap_8 FILLER_75_2318 ();
 sg13g2_decap_8 FILLER_75_2325 ();
 sg13g2_decap_8 FILLER_75_2332 ();
 sg13g2_decap_8 FILLER_75_2339 ();
 sg13g2_decap_8 FILLER_75_2346 ();
 sg13g2_decap_8 FILLER_75_2353 ();
 sg13g2_decap_8 FILLER_75_2360 ();
 sg13g2_decap_8 FILLER_75_2367 ();
 sg13g2_decap_8 FILLER_75_2374 ();
 sg13g2_decap_8 FILLER_75_2381 ();
 sg13g2_decap_8 FILLER_75_2388 ();
 sg13g2_decap_8 FILLER_75_2395 ();
 sg13g2_decap_8 FILLER_75_2402 ();
 sg13g2_decap_8 FILLER_75_2409 ();
 sg13g2_decap_8 FILLER_75_2416 ();
 sg13g2_decap_8 FILLER_75_2423 ();
 sg13g2_decap_8 FILLER_75_2430 ();
 sg13g2_decap_8 FILLER_75_2437 ();
 sg13g2_decap_8 FILLER_75_2444 ();
 sg13g2_decap_8 FILLER_75_2451 ();
 sg13g2_decap_8 FILLER_75_2458 ();
 sg13g2_decap_8 FILLER_75_2465 ();
 sg13g2_decap_8 FILLER_75_2472 ();
 sg13g2_decap_8 FILLER_75_2479 ();
 sg13g2_decap_8 FILLER_75_2486 ();
 sg13g2_decap_8 FILLER_75_2493 ();
 sg13g2_decap_8 FILLER_75_2500 ();
 sg13g2_decap_8 FILLER_75_2507 ();
 sg13g2_decap_8 FILLER_75_2514 ();
 sg13g2_decap_8 FILLER_75_2521 ();
 sg13g2_decap_8 FILLER_75_2528 ();
 sg13g2_decap_8 FILLER_75_2535 ();
 sg13g2_decap_8 FILLER_75_2542 ();
 sg13g2_decap_8 FILLER_75_2549 ();
 sg13g2_decap_8 FILLER_75_2556 ();
 sg13g2_decap_8 FILLER_75_2563 ();
 sg13g2_decap_8 FILLER_75_2570 ();
 sg13g2_decap_8 FILLER_75_2577 ();
 sg13g2_decap_8 FILLER_75_2584 ();
 sg13g2_decap_8 FILLER_75_2591 ();
 sg13g2_decap_8 FILLER_75_2598 ();
 sg13g2_decap_8 FILLER_75_2605 ();
 sg13g2_decap_8 FILLER_75_2612 ();
 sg13g2_decap_8 FILLER_75_2619 ();
 sg13g2_decap_8 FILLER_75_2626 ();
 sg13g2_decap_8 FILLER_75_2633 ();
 sg13g2_decap_8 FILLER_75_2640 ();
 sg13g2_decap_8 FILLER_75_2647 ();
 sg13g2_decap_8 FILLER_75_2654 ();
 sg13g2_decap_8 FILLER_75_2661 ();
 sg13g2_decap_4 FILLER_75_2668 ();
 sg13g2_fill_2 FILLER_75_2672 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_8 FILLER_76_189 ();
 sg13g2_decap_8 FILLER_76_196 ();
 sg13g2_decap_8 FILLER_76_203 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_decap_8 FILLER_76_217 ();
 sg13g2_decap_8 FILLER_76_224 ();
 sg13g2_decap_8 FILLER_76_231 ();
 sg13g2_decap_8 FILLER_76_238 ();
 sg13g2_decap_8 FILLER_76_245 ();
 sg13g2_decap_8 FILLER_76_252 ();
 sg13g2_decap_8 FILLER_76_259 ();
 sg13g2_decap_8 FILLER_76_266 ();
 sg13g2_decap_8 FILLER_76_273 ();
 sg13g2_decap_8 FILLER_76_280 ();
 sg13g2_decap_8 FILLER_76_287 ();
 sg13g2_decap_8 FILLER_76_294 ();
 sg13g2_decap_8 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_308 ();
 sg13g2_decap_8 FILLER_76_315 ();
 sg13g2_decap_8 FILLER_76_322 ();
 sg13g2_decap_8 FILLER_76_329 ();
 sg13g2_decap_8 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_decap_8 FILLER_76_357 ();
 sg13g2_decap_8 FILLER_76_364 ();
 sg13g2_decap_8 FILLER_76_371 ();
 sg13g2_decap_8 FILLER_76_378 ();
 sg13g2_decap_8 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_392 ();
 sg13g2_decap_8 FILLER_76_399 ();
 sg13g2_decap_8 FILLER_76_406 ();
 sg13g2_decap_8 FILLER_76_413 ();
 sg13g2_decap_8 FILLER_76_420 ();
 sg13g2_decap_8 FILLER_76_427 ();
 sg13g2_decap_8 FILLER_76_434 ();
 sg13g2_decap_8 FILLER_76_441 ();
 sg13g2_decap_8 FILLER_76_448 ();
 sg13g2_decap_8 FILLER_76_455 ();
 sg13g2_fill_2 FILLER_76_462 ();
 sg13g2_fill_1 FILLER_76_507 ();
 sg13g2_fill_1 FILLER_76_534 ();
 sg13g2_decap_4 FILLER_76_646 ();
 sg13g2_fill_2 FILLER_76_650 ();
 sg13g2_decap_8 FILLER_76_661 ();
 sg13g2_fill_2 FILLER_76_668 ();
 sg13g2_decap_4 FILLER_76_674 ();
 sg13g2_decap_8 FILLER_76_681 ();
 sg13g2_decap_4 FILLER_76_688 ();
 sg13g2_decap_8 FILLER_76_701 ();
 sg13g2_decap_8 FILLER_76_708 ();
 sg13g2_decap_8 FILLER_76_715 ();
 sg13g2_decap_8 FILLER_76_722 ();
 sg13g2_decap_8 FILLER_76_729 ();
 sg13g2_decap_8 FILLER_76_736 ();
 sg13g2_decap_8 FILLER_76_743 ();
 sg13g2_decap_8 FILLER_76_750 ();
 sg13g2_decap_8 FILLER_76_757 ();
 sg13g2_decap_8 FILLER_76_764 ();
 sg13g2_decap_8 FILLER_76_771 ();
 sg13g2_decap_8 FILLER_76_778 ();
 sg13g2_decap_8 FILLER_76_785 ();
 sg13g2_decap_8 FILLER_76_792 ();
 sg13g2_decap_8 FILLER_76_799 ();
 sg13g2_decap_8 FILLER_76_806 ();
 sg13g2_decap_8 FILLER_76_813 ();
 sg13g2_decap_8 FILLER_76_820 ();
 sg13g2_decap_8 FILLER_76_827 ();
 sg13g2_decap_8 FILLER_76_834 ();
 sg13g2_decap_8 FILLER_76_841 ();
 sg13g2_decap_8 FILLER_76_848 ();
 sg13g2_decap_8 FILLER_76_855 ();
 sg13g2_decap_8 FILLER_76_862 ();
 sg13g2_decap_8 FILLER_76_869 ();
 sg13g2_decap_8 FILLER_76_876 ();
 sg13g2_decap_8 FILLER_76_883 ();
 sg13g2_decap_8 FILLER_76_890 ();
 sg13g2_decap_8 FILLER_76_897 ();
 sg13g2_decap_8 FILLER_76_904 ();
 sg13g2_decap_8 FILLER_76_911 ();
 sg13g2_decap_4 FILLER_76_918 ();
 sg13g2_fill_2 FILLER_76_922 ();
 sg13g2_fill_2 FILLER_76_939 ();
 sg13g2_fill_2 FILLER_76_953 ();
 sg13g2_fill_1 FILLER_76_1011 ();
 sg13g2_fill_1 FILLER_76_1114 ();
 sg13g2_fill_1 FILLER_76_1141 ();
 sg13g2_fill_2 FILLER_76_1200 ();
 sg13g2_fill_1 FILLER_76_1271 ();
 sg13g2_fill_2 FILLER_76_1344 ();
 sg13g2_fill_2 FILLER_76_1355 ();
 sg13g2_fill_2 FILLER_76_1371 ();
 sg13g2_fill_1 FILLER_76_1444 ();
 sg13g2_decap_4 FILLER_76_1525 ();
 sg13g2_fill_2 FILLER_76_1529 ();
 sg13g2_fill_1 FILLER_76_1599 ();
 sg13g2_fill_1 FILLER_76_1616 ();
 sg13g2_fill_1 FILLER_76_1636 ();
 sg13g2_fill_1 FILLER_76_1673 ();
 sg13g2_fill_2 FILLER_76_1711 ();
 sg13g2_fill_2 FILLER_76_1739 ();
 sg13g2_fill_1 FILLER_76_1885 ();
 sg13g2_fill_1 FILLER_76_1900 ();
 sg13g2_fill_2 FILLER_76_1936 ();
 sg13g2_fill_1 FILLER_76_1970 ();
 sg13g2_fill_2 FILLER_76_1990 ();
 sg13g2_fill_2 FILLER_76_2002 ();
 sg13g2_fill_2 FILLER_76_2054 ();
 sg13g2_fill_1 FILLER_76_2056 ();
 sg13g2_fill_1 FILLER_76_2093 ();
 sg13g2_fill_2 FILLER_76_2120 ();
 sg13g2_fill_1 FILLER_76_2122 ();
 sg13g2_fill_2 FILLER_76_2238 ();
 sg13g2_fill_1 FILLER_76_2240 ();
 sg13g2_decap_8 FILLER_76_2267 ();
 sg13g2_decap_8 FILLER_76_2287 ();
 sg13g2_decap_8 FILLER_76_2294 ();
 sg13g2_decap_8 FILLER_76_2301 ();
 sg13g2_decap_8 FILLER_76_2308 ();
 sg13g2_decap_8 FILLER_76_2315 ();
 sg13g2_decap_8 FILLER_76_2322 ();
 sg13g2_decap_8 FILLER_76_2329 ();
 sg13g2_decap_8 FILLER_76_2336 ();
 sg13g2_decap_8 FILLER_76_2343 ();
 sg13g2_decap_8 FILLER_76_2350 ();
 sg13g2_decap_8 FILLER_76_2357 ();
 sg13g2_decap_8 FILLER_76_2364 ();
 sg13g2_decap_8 FILLER_76_2371 ();
 sg13g2_decap_8 FILLER_76_2378 ();
 sg13g2_decap_8 FILLER_76_2385 ();
 sg13g2_decap_8 FILLER_76_2392 ();
 sg13g2_decap_8 FILLER_76_2399 ();
 sg13g2_decap_8 FILLER_76_2406 ();
 sg13g2_decap_8 FILLER_76_2413 ();
 sg13g2_decap_8 FILLER_76_2420 ();
 sg13g2_decap_8 FILLER_76_2427 ();
 sg13g2_decap_8 FILLER_76_2434 ();
 sg13g2_decap_8 FILLER_76_2441 ();
 sg13g2_decap_8 FILLER_76_2448 ();
 sg13g2_decap_8 FILLER_76_2455 ();
 sg13g2_decap_8 FILLER_76_2462 ();
 sg13g2_decap_8 FILLER_76_2469 ();
 sg13g2_decap_8 FILLER_76_2476 ();
 sg13g2_decap_8 FILLER_76_2483 ();
 sg13g2_decap_8 FILLER_76_2490 ();
 sg13g2_decap_8 FILLER_76_2497 ();
 sg13g2_decap_8 FILLER_76_2504 ();
 sg13g2_decap_8 FILLER_76_2511 ();
 sg13g2_decap_8 FILLER_76_2518 ();
 sg13g2_decap_8 FILLER_76_2525 ();
 sg13g2_decap_8 FILLER_76_2532 ();
 sg13g2_decap_8 FILLER_76_2539 ();
 sg13g2_decap_8 FILLER_76_2546 ();
 sg13g2_decap_8 FILLER_76_2553 ();
 sg13g2_decap_8 FILLER_76_2560 ();
 sg13g2_decap_8 FILLER_76_2567 ();
 sg13g2_decap_8 FILLER_76_2574 ();
 sg13g2_decap_8 FILLER_76_2581 ();
 sg13g2_decap_8 FILLER_76_2588 ();
 sg13g2_decap_8 FILLER_76_2595 ();
 sg13g2_decap_8 FILLER_76_2602 ();
 sg13g2_decap_8 FILLER_76_2609 ();
 sg13g2_decap_8 FILLER_76_2616 ();
 sg13g2_decap_8 FILLER_76_2623 ();
 sg13g2_decap_8 FILLER_76_2630 ();
 sg13g2_decap_8 FILLER_76_2637 ();
 sg13g2_decap_8 FILLER_76_2644 ();
 sg13g2_decap_8 FILLER_76_2651 ();
 sg13g2_decap_8 FILLER_76_2658 ();
 sg13g2_decap_8 FILLER_76_2665 ();
 sg13g2_fill_2 FILLER_76_2672 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_8 FILLER_77_217 ();
 sg13g2_decap_8 FILLER_77_224 ();
 sg13g2_decap_8 FILLER_77_231 ();
 sg13g2_decap_8 FILLER_77_238 ();
 sg13g2_decap_8 FILLER_77_245 ();
 sg13g2_decap_8 FILLER_77_252 ();
 sg13g2_decap_8 FILLER_77_259 ();
 sg13g2_decap_8 FILLER_77_266 ();
 sg13g2_decap_8 FILLER_77_273 ();
 sg13g2_decap_8 FILLER_77_280 ();
 sg13g2_decap_8 FILLER_77_287 ();
 sg13g2_decap_8 FILLER_77_294 ();
 sg13g2_decap_8 FILLER_77_301 ();
 sg13g2_decap_8 FILLER_77_308 ();
 sg13g2_decap_8 FILLER_77_315 ();
 sg13g2_decap_8 FILLER_77_322 ();
 sg13g2_decap_8 FILLER_77_329 ();
 sg13g2_decap_8 FILLER_77_336 ();
 sg13g2_decap_8 FILLER_77_343 ();
 sg13g2_decap_8 FILLER_77_350 ();
 sg13g2_decap_8 FILLER_77_357 ();
 sg13g2_decap_8 FILLER_77_364 ();
 sg13g2_decap_8 FILLER_77_371 ();
 sg13g2_decap_8 FILLER_77_378 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_decap_8 FILLER_77_406 ();
 sg13g2_decap_8 FILLER_77_413 ();
 sg13g2_decap_8 FILLER_77_420 ();
 sg13g2_decap_8 FILLER_77_427 ();
 sg13g2_decap_8 FILLER_77_434 ();
 sg13g2_decap_8 FILLER_77_441 ();
 sg13g2_decap_8 FILLER_77_448 ();
 sg13g2_decap_8 FILLER_77_455 ();
 sg13g2_decap_8 FILLER_77_462 ();
 sg13g2_decap_4 FILLER_77_469 ();
 sg13g2_fill_2 FILLER_77_473 ();
 sg13g2_fill_1 FILLER_77_511 ();
 sg13g2_fill_2 FILLER_77_542 ();
 sg13g2_fill_2 FILLER_77_550 ();
 sg13g2_decap_8 FILLER_77_645 ();
 sg13g2_decap_8 FILLER_77_652 ();
 sg13g2_decap_8 FILLER_77_659 ();
 sg13g2_decap_8 FILLER_77_666 ();
 sg13g2_decap_8 FILLER_77_673 ();
 sg13g2_decap_8 FILLER_77_680 ();
 sg13g2_decap_8 FILLER_77_687 ();
 sg13g2_decap_8 FILLER_77_694 ();
 sg13g2_decap_8 FILLER_77_701 ();
 sg13g2_decap_8 FILLER_77_708 ();
 sg13g2_decap_8 FILLER_77_715 ();
 sg13g2_decap_8 FILLER_77_722 ();
 sg13g2_decap_8 FILLER_77_729 ();
 sg13g2_decap_8 FILLER_77_736 ();
 sg13g2_decap_8 FILLER_77_743 ();
 sg13g2_decap_8 FILLER_77_750 ();
 sg13g2_decap_8 FILLER_77_757 ();
 sg13g2_decap_8 FILLER_77_764 ();
 sg13g2_decap_8 FILLER_77_771 ();
 sg13g2_decap_8 FILLER_77_778 ();
 sg13g2_decap_8 FILLER_77_785 ();
 sg13g2_decap_8 FILLER_77_792 ();
 sg13g2_decap_8 FILLER_77_799 ();
 sg13g2_decap_8 FILLER_77_806 ();
 sg13g2_decap_8 FILLER_77_813 ();
 sg13g2_decap_8 FILLER_77_820 ();
 sg13g2_decap_8 FILLER_77_827 ();
 sg13g2_decap_8 FILLER_77_834 ();
 sg13g2_decap_8 FILLER_77_841 ();
 sg13g2_decap_8 FILLER_77_848 ();
 sg13g2_decap_8 FILLER_77_855 ();
 sg13g2_decap_8 FILLER_77_862 ();
 sg13g2_decap_8 FILLER_77_869 ();
 sg13g2_decap_8 FILLER_77_876 ();
 sg13g2_decap_8 FILLER_77_883 ();
 sg13g2_decap_8 FILLER_77_890 ();
 sg13g2_decap_8 FILLER_77_897 ();
 sg13g2_decap_8 FILLER_77_904 ();
 sg13g2_decap_8 FILLER_77_911 ();
 sg13g2_decap_8 FILLER_77_918 ();
 sg13g2_decap_4 FILLER_77_925 ();
 sg13g2_fill_1 FILLER_77_935 ();
 sg13g2_fill_1 FILLER_77_947 ();
 sg13g2_fill_1 FILLER_77_978 ();
 sg13g2_fill_2 FILLER_77_1055 ();
 sg13g2_fill_2 FILLER_77_1093 ();
 sg13g2_fill_1 FILLER_77_1267 ();
 sg13g2_fill_2 FILLER_77_1355 ();
 sg13g2_fill_2 FILLER_77_1446 ();
 sg13g2_decap_8 FILLER_77_1518 ();
 sg13g2_decap_4 FILLER_77_1525 ();
 sg13g2_fill_1 FILLER_77_1529 ();
 sg13g2_fill_1 FILLER_77_1565 ();
 sg13g2_fill_2 FILLER_77_1580 ();
 sg13g2_fill_2 FILLER_77_1707 ();
 sg13g2_fill_1 FILLER_77_1709 ();
 sg13g2_fill_1 FILLER_77_1724 ();
 sg13g2_decap_4 FILLER_77_1747 ();
 sg13g2_fill_2 FILLER_77_1793 ();
 sg13g2_fill_1 FILLER_77_1809 ();
 sg13g2_fill_1 FILLER_77_1834 ();
 sg13g2_fill_2 FILLER_77_1864 ();
 sg13g2_fill_1 FILLER_77_1866 ();
 sg13g2_fill_2 FILLER_77_1908 ();
 sg13g2_fill_1 FILLER_77_1910 ();
 sg13g2_decap_4 FILLER_77_1973 ();
 sg13g2_fill_2 FILLER_77_2079 ();
 sg13g2_fill_1 FILLER_77_2081 ();
 sg13g2_fill_2 FILLER_77_2118 ();
 sg13g2_fill_1 FILLER_77_2120 ();
 sg13g2_fill_2 FILLER_77_2131 ();
 sg13g2_fill_1 FILLER_77_2133 ();
 sg13g2_decap_8 FILLER_77_2147 ();
 sg13g2_fill_1 FILLER_77_2154 ();
 sg13g2_decap_8 FILLER_77_2159 ();
 sg13g2_decap_4 FILLER_77_2166 ();
 sg13g2_fill_2 FILLER_77_2170 ();
 sg13g2_decap_8 FILLER_77_2198 ();
 sg13g2_decap_8 FILLER_77_2205 ();
 sg13g2_decap_8 FILLER_77_2212 ();
 sg13g2_fill_2 FILLER_77_2219 ();
 sg13g2_fill_1 FILLER_77_2221 ();
 sg13g2_decap_8 FILLER_77_2235 ();
 sg13g2_fill_2 FILLER_77_2242 ();
 sg13g2_fill_1 FILLER_77_2244 ();
 sg13g2_fill_1 FILLER_77_2253 ();
 sg13g2_decap_8 FILLER_77_2263 ();
 sg13g2_decap_8 FILLER_77_2270 ();
 sg13g2_decap_8 FILLER_77_2277 ();
 sg13g2_decap_8 FILLER_77_2284 ();
 sg13g2_decap_8 FILLER_77_2291 ();
 sg13g2_decap_8 FILLER_77_2298 ();
 sg13g2_decap_8 FILLER_77_2305 ();
 sg13g2_decap_8 FILLER_77_2312 ();
 sg13g2_decap_8 FILLER_77_2319 ();
 sg13g2_decap_8 FILLER_77_2326 ();
 sg13g2_decap_8 FILLER_77_2333 ();
 sg13g2_decap_8 FILLER_77_2340 ();
 sg13g2_decap_8 FILLER_77_2347 ();
 sg13g2_decap_8 FILLER_77_2354 ();
 sg13g2_decap_8 FILLER_77_2361 ();
 sg13g2_decap_8 FILLER_77_2368 ();
 sg13g2_decap_8 FILLER_77_2375 ();
 sg13g2_decap_8 FILLER_77_2382 ();
 sg13g2_decap_8 FILLER_77_2389 ();
 sg13g2_decap_8 FILLER_77_2396 ();
 sg13g2_decap_8 FILLER_77_2403 ();
 sg13g2_decap_8 FILLER_77_2410 ();
 sg13g2_decap_8 FILLER_77_2417 ();
 sg13g2_decap_8 FILLER_77_2424 ();
 sg13g2_decap_8 FILLER_77_2431 ();
 sg13g2_decap_8 FILLER_77_2438 ();
 sg13g2_decap_8 FILLER_77_2445 ();
 sg13g2_decap_8 FILLER_77_2452 ();
 sg13g2_decap_8 FILLER_77_2459 ();
 sg13g2_decap_8 FILLER_77_2466 ();
 sg13g2_decap_8 FILLER_77_2473 ();
 sg13g2_decap_8 FILLER_77_2480 ();
 sg13g2_decap_8 FILLER_77_2487 ();
 sg13g2_decap_8 FILLER_77_2494 ();
 sg13g2_decap_8 FILLER_77_2501 ();
 sg13g2_decap_8 FILLER_77_2508 ();
 sg13g2_decap_8 FILLER_77_2515 ();
 sg13g2_decap_8 FILLER_77_2522 ();
 sg13g2_decap_8 FILLER_77_2529 ();
 sg13g2_decap_8 FILLER_77_2536 ();
 sg13g2_decap_8 FILLER_77_2543 ();
 sg13g2_decap_8 FILLER_77_2550 ();
 sg13g2_decap_8 FILLER_77_2557 ();
 sg13g2_decap_8 FILLER_77_2564 ();
 sg13g2_decap_8 FILLER_77_2571 ();
 sg13g2_decap_8 FILLER_77_2578 ();
 sg13g2_decap_8 FILLER_77_2585 ();
 sg13g2_decap_8 FILLER_77_2592 ();
 sg13g2_decap_8 FILLER_77_2599 ();
 sg13g2_decap_8 FILLER_77_2606 ();
 sg13g2_decap_8 FILLER_77_2613 ();
 sg13g2_decap_8 FILLER_77_2620 ();
 sg13g2_decap_8 FILLER_77_2627 ();
 sg13g2_decap_8 FILLER_77_2634 ();
 sg13g2_decap_8 FILLER_77_2641 ();
 sg13g2_decap_8 FILLER_77_2648 ();
 sg13g2_decap_8 FILLER_77_2655 ();
 sg13g2_decap_8 FILLER_77_2662 ();
 sg13g2_decap_4 FILLER_77_2669 ();
 sg13g2_fill_1 FILLER_77_2673 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_203 ();
 sg13g2_decap_8 FILLER_78_210 ();
 sg13g2_decap_8 FILLER_78_217 ();
 sg13g2_decap_8 FILLER_78_224 ();
 sg13g2_decap_8 FILLER_78_231 ();
 sg13g2_decap_8 FILLER_78_238 ();
 sg13g2_decap_8 FILLER_78_245 ();
 sg13g2_decap_8 FILLER_78_252 ();
 sg13g2_decap_8 FILLER_78_259 ();
 sg13g2_decap_8 FILLER_78_266 ();
 sg13g2_decap_8 FILLER_78_273 ();
 sg13g2_decap_8 FILLER_78_280 ();
 sg13g2_decap_8 FILLER_78_287 ();
 sg13g2_decap_8 FILLER_78_294 ();
 sg13g2_decap_8 FILLER_78_301 ();
 sg13g2_decap_8 FILLER_78_308 ();
 sg13g2_decap_8 FILLER_78_315 ();
 sg13g2_decap_8 FILLER_78_322 ();
 sg13g2_decap_8 FILLER_78_329 ();
 sg13g2_decap_8 FILLER_78_336 ();
 sg13g2_decap_8 FILLER_78_343 ();
 sg13g2_decap_8 FILLER_78_350 ();
 sg13g2_decap_8 FILLER_78_357 ();
 sg13g2_decap_8 FILLER_78_364 ();
 sg13g2_decap_8 FILLER_78_371 ();
 sg13g2_decap_8 FILLER_78_378 ();
 sg13g2_decap_8 FILLER_78_385 ();
 sg13g2_decap_8 FILLER_78_392 ();
 sg13g2_decap_8 FILLER_78_399 ();
 sg13g2_decap_8 FILLER_78_406 ();
 sg13g2_decap_8 FILLER_78_413 ();
 sg13g2_decap_8 FILLER_78_420 ();
 sg13g2_decap_8 FILLER_78_427 ();
 sg13g2_decap_8 FILLER_78_434 ();
 sg13g2_decap_8 FILLER_78_441 ();
 sg13g2_decap_8 FILLER_78_448 ();
 sg13g2_decap_8 FILLER_78_455 ();
 sg13g2_decap_8 FILLER_78_462 ();
 sg13g2_decap_8 FILLER_78_469 ();
 sg13g2_decap_4 FILLER_78_476 ();
 sg13g2_fill_2 FILLER_78_480 ();
 sg13g2_fill_1 FILLER_78_570 ();
 sg13g2_fill_2 FILLER_78_583 ();
 sg13g2_fill_1 FILLER_78_585 ();
 sg13g2_fill_1 FILLER_78_594 ();
 sg13g2_decap_8 FILLER_78_644 ();
 sg13g2_decap_8 FILLER_78_651 ();
 sg13g2_decap_8 FILLER_78_658 ();
 sg13g2_decap_8 FILLER_78_665 ();
 sg13g2_decap_8 FILLER_78_672 ();
 sg13g2_decap_8 FILLER_78_679 ();
 sg13g2_decap_8 FILLER_78_686 ();
 sg13g2_decap_8 FILLER_78_693 ();
 sg13g2_decap_8 FILLER_78_700 ();
 sg13g2_decap_8 FILLER_78_707 ();
 sg13g2_decap_8 FILLER_78_714 ();
 sg13g2_decap_8 FILLER_78_721 ();
 sg13g2_decap_8 FILLER_78_728 ();
 sg13g2_decap_8 FILLER_78_735 ();
 sg13g2_decap_8 FILLER_78_742 ();
 sg13g2_decap_8 FILLER_78_749 ();
 sg13g2_decap_8 FILLER_78_756 ();
 sg13g2_decap_8 FILLER_78_763 ();
 sg13g2_decap_8 FILLER_78_770 ();
 sg13g2_decap_8 FILLER_78_777 ();
 sg13g2_decap_8 FILLER_78_784 ();
 sg13g2_decap_8 FILLER_78_791 ();
 sg13g2_decap_8 FILLER_78_798 ();
 sg13g2_decap_8 FILLER_78_805 ();
 sg13g2_decap_8 FILLER_78_812 ();
 sg13g2_decap_8 FILLER_78_819 ();
 sg13g2_decap_8 FILLER_78_826 ();
 sg13g2_decap_8 FILLER_78_833 ();
 sg13g2_decap_8 FILLER_78_840 ();
 sg13g2_decap_8 FILLER_78_847 ();
 sg13g2_decap_8 FILLER_78_854 ();
 sg13g2_decap_8 FILLER_78_861 ();
 sg13g2_decap_8 FILLER_78_868 ();
 sg13g2_decap_8 FILLER_78_875 ();
 sg13g2_decap_8 FILLER_78_882 ();
 sg13g2_decap_8 FILLER_78_889 ();
 sg13g2_decap_8 FILLER_78_896 ();
 sg13g2_decap_8 FILLER_78_903 ();
 sg13g2_decap_8 FILLER_78_910 ();
 sg13g2_decap_8 FILLER_78_917 ();
 sg13g2_decap_8 FILLER_78_924 ();
 sg13g2_fill_1 FILLER_78_931 ();
 sg13g2_fill_1 FILLER_78_948 ();
 sg13g2_fill_1 FILLER_78_978 ();
 sg13g2_fill_1 FILLER_78_1156 ();
 sg13g2_fill_1 FILLER_78_1269 ();
 sg13g2_fill_1 FILLER_78_1289 ();
 sg13g2_fill_2 FILLER_78_1340 ();
 sg13g2_fill_1 FILLER_78_1412 ();
 sg13g2_fill_1 FILLER_78_1439 ();
 sg13g2_fill_2 FILLER_78_1454 ();
 sg13g2_decap_8 FILLER_78_1511 ();
 sg13g2_decap_8 FILLER_78_1518 ();
 sg13g2_decap_8 FILLER_78_1525 ();
 sg13g2_decap_8 FILLER_78_1532 ();
 sg13g2_decap_8 FILLER_78_1539 ();
 sg13g2_decap_8 FILLER_78_1546 ();
 sg13g2_fill_1 FILLER_78_1604 ();
 sg13g2_fill_1 FILLER_78_1614 ();
 sg13g2_fill_2 FILLER_78_1690 ();
 sg13g2_fill_1 FILLER_78_1692 ();
 sg13g2_fill_2 FILLER_78_1724 ();
 sg13g2_fill_1 FILLER_78_1726 ();
 sg13g2_decap_8 FILLER_78_1763 ();
 sg13g2_fill_1 FILLER_78_1832 ();
 sg13g2_fill_1 FILLER_78_1843 ();
 sg13g2_decap_8 FILLER_78_1874 ();
 sg13g2_fill_2 FILLER_78_1881 ();
 sg13g2_fill_2 FILLER_78_1910 ();
 sg13g2_fill_2 FILLER_78_1961 ();
 sg13g2_fill_2 FILLER_78_1987 ();
 sg13g2_fill_1 FILLER_78_1998 ();
 sg13g2_fill_2 FILLER_78_2060 ();
 sg13g2_decap_8 FILLER_78_2098 ();
 sg13g2_decap_8 FILLER_78_2157 ();
 sg13g2_decap_8 FILLER_78_2164 ();
 sg13g2_decap_4 FILLER_78_2171 ();
 sg13g2_fill_1 FILLER_78_2175 ();
 sg13g2_decap_8 FILLER_78_2194 ();
 sg13g2_decap_8 FILLER_78_2201 ();
 sg13g2_decap_8 FILLER_78_2208 ();
 sg13g2_decap_8 FILLER_78_2215 ();
 sg13g2_decap_8 FILLER_78_2222 ();
 sg13g2_decap_8 FILLER_78_2229 ();
 sg13g2_decap_8 FILLER_78_2236 ();
 sg13g2_decap_8 FILLER_78_2243 ();
 sg13g2_decap_8 FILLER_78_2250 ();
 sg13g2_decap_8 FILLER_78_2257 ();
 sg13g2_decap_8 FILLER_78_2264 ();
 sg13g2_decap_8 FILLER_78_2271 ();
 sg13g2_decap_8 FILLER_78_2278 ();
 sg13g2_decap_8 FILLER_78_2285 ();
 sg13g2_decap_8 FILLER_78_2292 ();
 sg13g2_decap_8 FILLER_78_2299 ();
 sg13g2_decap_8 FILLER_78_2306 ();
 sg13g2_decap_8 FILLER_78_2313 ();
 sg13g2_decap_8 FILLER_78_2320 ();
 sg13g2_decap_8 FILLER_78_2327 ();
 sg13g2_decap_8 FILLER_78_2334 ();
 sg13g2_decap_8 FILLER_78_2341 ();
 sg13g2_decap_8 FILLER_78_2348 ();
 sg13g2_decap_8 FILLER_78_2355 ();
 sg13g2_decap_8 FILLER_78_2362 ();
 sg13g2_decap_8 FILLER_78_2369 ();
 sg13g2_decap_8 FILLER_78_2376 ();
 sg13g2_decap_8 FILLER_78_2383 ();
 sg13g2_decap_8 FILLER_78_2390 ();
 sg13g2_decap_8 FILLER_78_2397 ();
 sg13g2_decap_8 FILLER_78_2404 ();
 sg13g2_decap_8 FILLER_78_2411 ();
 sg13g2_decap_8 FILLER_78_2418 ();
 sg13g2_decap_8 FILLER_78_2425 ();
 sg13g2_decap_8 FILLER_78_2432 ();
 sg13g2_decap_8 FILLER_78_2439 ();
 sg13g2_decap_8 FILLER_78_2446 ();
 sg13g2_decap_8 FILLER_78_2453 ();
 sg13g2_decap_8 FILLER_78_2460 ();
 sg13g2_decap_8 FILLER_78_2467 ();
 sg13g2_decap_8 FILLER_78_2474 ();
 sg13g2_decap_8 FILLER_78_2481 ();
 sg13g2_decap_8 FILLER_78_2488 ();
 sg13g2_decap_8 FILLER_78_2495 ();
 sg13g2_decap_8 FILLER_78_2502 ();
 sg13g2_decap_8 FILLER_78_2509 ();
 sg13g2_decap_8 FILLER_78_2516 ();
 sg13g2_decap_8 FILLER_78_2523 ();
 sg13g2_decap_8 FILLER_78_2530 ();
 sg13g2_decap_8 FILLER_78_2537 ();
 sg13g2_decap_8 FILLER_78_2544 ();
 sg13g2_decap_8 FILLER_78_2551 ();
 sg13g2_decap_8 FILLER_78_2558 ();
 sg13g2_decap_8 FILLER_78_2565 ();
 sg13g2_decap_8 FILLER_78_2572 ();
 sg13g2_decap_8 FILLER_78_2579 ();
 sg13g2_decap_8 FILLER_78_2586 ();
 sg13g2_decap_8 FILLER_78_2593 ();
 sg13g2_decap_8 FILLER_78_2600 ();
 sg13g2_decap_8 FILLER_78_2607 ();
 sg13g2_decap_8 FILLER_78_2614 ();
 sg13g2_decap_8 FILLER_78_2621 ();
 sg13g2_decap_8 FILLER_78_2628 ();
 sg13g2_decap_8 FILLER_78_2635 ();
 sg13g2_decap_8 FILLER_78_2642 ();
 sg13g2_decap_8 FILLER_78_2649 ();
 sg13g2_decap_8 FILLER_78_2656 ();
 sg13g2_decap_8 FILLER_78_2663 ();
 sg13g2_decap_4 FILLER_78_2670 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_decap_8 FILLER_79_231 ();
 sg13g2_decap_8 FILLER_79_238 ();
 sg13g2_decap_8 FILLER_79_245 ();
 sg13g2_decap_8 FILLER_79_252 ();
 sg13g2_decap_8 FILLER_79_259 ();
 sg13g2_decap_8 FILLER_79_266 ();
 sg13g2_decap_8 FILLER_79_273 ();
 sg13g2_decap_8 FILLER_79_280 ();
 sg13g2_decap_8 FILLER_79_287 ();
 sg13g2_decap_8 FILLER_79_294 ();
 sg13g2_decap_8 FILLER_79_301 ();
 sg13g2_decap_8 FILLER_79_308 ();
 sg13g2_decap_8 FILLER_79_315 ();
 sg13g2_decap_8 FILLER_79_322 ();
 sg13g2_decap_8 FILLER_79_329 ();
 sg13g2_decap_8 FILLER_79_336 ();
 sg13g2_decap_8 FILLER_79_343 ();
 sg13g2_decap_8 FILLER_79_350 ();
 sg13g2_decap_8 FILLER_79_357 ();
 sg13g2_decap_8 FILLER_79_364 ();
 sg13g2_decap_8 FILLER_79_371 ();
 sg13g2_decap_8 FILLER_79_378 ();
 sg13g2_decap_8 FILLER_79_385 ();
 sg13g2_decap_8 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_decap_8 FILLER_79_406 ();
 sg13g2_decap_8 FILLER_79_413 ();
 sg13g2_decap_8 FILLER_79_420 ();
 sg13g2_decap_8 FILLER_79_427 ();
 sg13g2_decap_8 FILLER_79_434 ();
 sg13g2_decap_8 FILLER_79_441 ();
 sg13g2_decap_8 FILLER_79_448 ();
 sg13g2_decap_8 FILLER_79_455 ();
 sg13g2_decap_8 FILLER_79_462 ();
 sg13g2_decap_8 FILLER_79_469 ();
 sg13g2_decap_8 FILLER_79_476 ();
 sg13g2_decap_8 FILLER_79_483 ();
 sg13g2_fill_1 FILLER_79_529 ();
 sg13g2_fill_1 FILLER_79_547 ();
 sg13g2_decap_8 FILLER_79_583 ();
 sg13g2_decap_8 FILLER_79_590 ();
 sg13g2_decap_4 FILLER_79_597 ();
 sg13g2_fill_2 FILLER_79_601 ();
 sg13g2_decap_8 FILLER_79_632 ();
 sg13g2_decap_8 FILLER_79_639 ();
 sg13g2_decap_8 FILLER_79_646 ();
 sg13g2_decap_8 FILLER_79_653 ();
 sg13g2_decap_8 FILLER_79_660 ();
 sg13g2_decap_8 FILLER_79_667 ();
 sg13g2_decap_8 FILLER_79_674 ();
 sg13g2_decap_8 FILLER_79_681 ();
 sg13g2_decap_8 FILLER_79_688 ();
 sg13g2_decap_8 FILLER_79_695 ();
 sg13g2_decap_8 FILLER_79_702 ();
 sg13g2_decap_8 FILLER_79_709 ();
 sg13g2_decap_8 FILLER_79_716 ();
 sg13g2_decap_8 FILLER_79_723 ();
 sg13g2_decap_8 FILLER_79_730 ();
 sg13g2_decap_8 FILLER_79_737 ();
 sg13g2_decap_8 FILLER_79_744 ();
 sg13g2_decap_8 FILLER_79_751 ();
 sg13g2_decap_8 FILLER_79_758 ();
 sg13g2_decap_8 FILLER_79_765 ();
 sg13g2_decap_8 FILLER_79_772 ();
 sg13g2_decap_8 FILLER_79_779 ();
 sg13g2_decap_8 FILLER_79_786 ();
 sg13g2_decap_8 FILLER_79_793 ();
 sg13g2_decap_8 FILLER_79_800 ();
 sg13g2_decap_8 FILLER_79_807 ();
 sg13g2_decap_8 FILLER_79_814 ();
 sg13g2_decap_8 FILLER_79_821 ();
 sg13g2_decap_8 FILLER_79_828 ();
 sg13g2_decap_8 FILLER_79_835 ();
 sg13g2_decap_8 FILLER_79_842 ();
 sg13g2_decap_8 FILLER_79_849 ();
 sg13g2_decap_8 FILLER_79_856 ();
 sg13g2_decap_8 FILLER_79_863 ();
 sg13g2_decap_8 FILLER_79_870 ();
 sg13g2_decap_8 FILLER_79_877 ();
 sg13g2_decap_8 FILLER_79_884 ();
 sg13g2_decap_8 FILLER_79_891 ();
 sg13g2_decap_8 FILLER_79_898 ();
 sg13g2_decap_8 FILLER_79_905 ();
 sg13g2_decap_8 FILLER_79_912 ();
 sg13g2_decap_8 FILLER_79_919 ();
 sg13g2_decap_8 FILLER_79_926 ();
 sg13g2_decap_4 FILLER_79_933 ();
 sg13g2_fill_2 FILLER_79_937 ();
 sg13g2_fill_2 FILLER_79_1012 ();
 sg13g2_fill_2 FILLER_79_1168 ();
 sg13g2_fill_1 FILLER_79_1283 ();
 sg13g2_fill_1 FILLER_79_1385 ();
 sg13g2_decap_8 FILLER_79_1503 ();
 sg13g2_decap_8 FILLER_79_1510 ();
 sg13g2_decap_8 FILLER_79_1517 ();
 sg13g2_decap_8 FILLER_79_1524 ();
 sg13g2_decap_8 FILLER_79_1531 ();
 sg13g2_decap_8 FILLER_79_1538 ();
 sg13g2_decap_8 FILLER_79_1545 ();
 sg13g2_decap_8 FILLER_79_1552 ();
 sg13g2_fill_2 FILLER_79_1559 ();
 sg13g2_fill_1 FILLER_79_1579 ();
 sg13g2_fill_1 FILLER_79_1613 ();
 sg13g2_decap_8 FILLER_79_1653 ();
 sg13g2_decap_8 FILLER_79_1660 ();
 sg13g2_decap_8 FILLER_79_1667 ();
 sg13g2_decap_4 FILLER_79_1674 ();
 sg13g2_fill_2 FILLER_79_1722 ();
 sg13g2_fill_1 FILLER_79_1724 ();
 sg13g2_decap_4 FILLER_79_1735 ();
 sg13g2_decap_4 FILLER_79_1762 ();
 sg13g2_fill_2 FILLER_79_1783 ();
 sg13g2_fill_2 FILLER_79_1800 ();
 sg13g2_fill_1 FILLER_79_1811 ();
 sg13g2_fill_1 FILLER_79_1817 ();
 sg13g2_fill_1 FILLER_79_1870 ();
 sg13g2_fill_2 FILLER_79_2021 ();
 sg13g2_decap_8 FILLER_79_2067 ();
 sg13g2_decap_8 FILLER_79_2074 ();
 sg13g2_decap_8 FILLER_79_2081 ();
 sg13g2_decap_8 FILLER_79_2088 ();
 sg13g2_decap_8 FILLER_79_2095 ();
 sg13g2_decap_8 FILLER_79_2102 ();
 sg13g2_fill_2 FILLER_79_2126 ();
 sg13g2_fill_1 FILLER_79_2128 ();
 sg13g2_decap_8 FILLER_79_2142 ();
 sg13g2_decap_8 FILLER_79_2149 ();
 sg13g2_decap_8 FILLER_79_2156 ();
 sg13g2_decap_8 FILLER_79_2163 ();
 sg13g2_decap_8 FILLER_79_2170 ();
 sg13g2_decap_4 FILLER_79_2177 ();
 sg13g2_fill_2 FILLER_79_2181 ();
 sg13g2_decap_8 FILLER_79_2187 ();
 sg13g2_decap_8 FILLER_79_2194 ();
 sg13g2_decap_8 FILLER_79_2201 ();
 sg13g2_decap_8 FILLER_79_2208 ();
 sg13g2_decap_8 FILLER_79_2215 ();
 sg13g2_decap_8 FILLER_79_2222 ();
 sg13g2_decap_8 FILLER_79_2229 ();
 sg13g2_decap_8 FILLER_79_2236 ();
 sg13g2_decap_8 FILLER_79_2243 ();
 sg13g2_decap_8 FILLER_79_2250 ();
 sg13g2_decap_8 FILLER_79_2257 ();
 sg13g2_decap_8 FILLER_79_2264 ();
 sg13g2_decap_8 FILLER_79_2271 ();
 sg13g2_decap_8 FILLER_79_2278 ();
 sg13g2_decap_8 FILLER_79_2285 ();
 sg13g2_decap_8 FILLER_79_2292 ();
 sg13g2_decap_8 FILLER_79_2299 ();
 sg13g2_decap_8 FILLER_79_2306 ();
 sg13g2_decap_8 FILLER_79_2313 ();
 sg13g2_decap_8 FILLER_79_2320 ();
 sg13g2_decap_8 FILLER_79_2327 ();
 sg13g2_decap_8 FILLER_79_2334 ();
 sg13g2_decap_8 FILLER_79_2341 ();
 sg13g2_decap_8 FILLER_79_2348 ();
 sg13g2_decap_8 FILLER_79_2355 ();
 sg13g2_decap_8 FILLER_79_2362 ();
 sg13g2_decap_8 FILLER_79_2369 ();
 sg13g2_decap_8 FILLER_79_2376 ();
 sg13g2_decap_8 FILLER_79_2383 ();
 sg13g2_decap_8 FILLER_79_2390 ();
 sg13g2_decap_8 FILLER_79_2397 ();
 sg13g2_decap_8 FILLER_79_2404 ();
 sg13g2_decap_8 FILLER_79_2411 ();
 sg13g2_decap_8 FILLER_79_2418 ();
 sg13g2_decap_8 FILLER_79_2425 ();
 sg13g2_decap_8 FILLER_79_2432 ();
 sg13g2_decap_8 FILLER_79_2439 ();
 sg13g2_decap_8 FILLER_79_2446 ();
 sg13g2_decap_8 FILLER_79_2453 ();
 sg13g2_decap_8 FILLER_79_2460 ();
 sg13g2_decap_8 FILLER_79_2467 ();
 sg13g2_decap_8 FILLER_79_2474 ();
 sg13g2_decap_8 FILLER_79_2481 ();
 sg13g2_decap_8 FILLER_79_2488 ();
 sg13g2_decap_8 FILLER_79_2495 ();
 sg13g2_decap_8 FILLER_79_2502 ();
 sg13g2_decap_8 FILLER_79_2509 ();
 sg13g2_decap_8 FILLER_79_2516 ();
 sg13g2_decap_8 FILLER_79_2523 ();
 sg13g2_decap_8 FILLER_79_2530 ();
 sg13g2_decap_8 FILLER_79_2537 ();
 sg13g2_decap_8 FILLER_79_2544 ();
 sg13g2_decap_8 FILLER_79_2551 ();
 sg13g2_decap_8 FILLER_79_2558 ();
 sg13g2_decap_8 FILLER_79_2565 ();
 sg13g2_decap_8 FILLER_79_2572 ();
 sg13g2_decap_8 FILLER_79_2579 ();
 sg13g2_decap_8 FILLER_79_2586 ();
 sg13g2_decap_8 FILLER_79_2593 ();
 sg13g2_decap_8 FILLER_79_2600 ();
 sg13g2_decap_8 FILLER_79_2607 ();
 sg13g2_decap_8 FILLER_79_2614 ();
 sg13g2_decap_8 FILLER_79_2621 ();
 sg13g2_decap_8 FILLER_79_2628 ();
 sg13g2_decap_8 FILLER_79_2635 ();
 sg13g2_decap_8 FILLER_79_2642 ();
 sg13g2_decap_8 FILLER_79_2649 ();
 sg13g2_decap_8 FILLER_79_2656 ();
 sg13g2_decap_8 FILLER_79_2663 ();
 sg13g2_decap_4 FILLER_79_2670 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_4 FILLER_80_180 ();
 sg13g2_decap_4 FILLER_80_188 ();
 sg13g2_decap_4 FILLER_80_196 ();
 sg13g2_decap_4 FILLER_80_204 ();
 sg13g2_decap_4 FILLER_80_212 ();
 sg13g2_decap_8 FILLER_80_220 ();
 sg13g2_decap_8 FILLER_80_227 ();
 sg13g2_decap_8 FILLER_80_234 ();
 sg13g2_decap_8 FILLER_80_241 ();
 sg13g2_decap_8 FILLER_80_248 ();
 sg13g2_decap_8 FILLER_80_255 ();
 sg13g2_decap_8 FILLER_80_262 ();
 sg13g2_decap_8 FILLER_80_269 ();
 sg13g2_decap_8 FILLER_80_276 ();
 sg13g2_decap_8 FILLER_80_283 ();
 sg13g2_decap_8 FILLER_80_290 ();
 sg13g2_decap_8 FILLER_80_297 ();
 sg13g2_decap_8 FILLER_80_304 ();
 sg13g2_decap_8 FILLER_80_311 ();
 sg13g2_decap_8 FILLER_80_318 ();
 sg13g2_decap_8 FILLER_80_325 ();
 sg13g2_decap_8 FILLER_80_332 ();
 sg13g2_decap_8 FILLER_80_339 ();
 sg13g2_decap_8 FILLER_80_346 ();
 sg13g2_decap_8 FILLER_80_353 ();
 sg13g2_decap_8 FILLER_80_364 ();
 sg13g2_decap_8 FILLER_80_371 ();
 sg13g2_decap_8 FILLER_80_378 ();
 sg13g2_decap_8 FILLER_80_385 ();
 sg13g2_decap_8 FILLER_80_392 ();
 sg13g2_decap_8 FILLER_80_399 ();
 sg13g2_decap_8 FILLER_80_406 ();
 sg13g2_decap_8 FILLER_80_413 ();
 sg13g2_decap_8 FILLER_80_420 ();
 sg13g2_decap_8 FILLER_80_427 ();
 sg13g2_decap_8 FILLER_80_434 ();
 sg13g2_decap_8 FILLER_80_441 ();
 sg13g2_decap_8 FILLER_80_448 ();
 sg13g2_decap_8 FILLER_80_455 ();
 sg13g2_decap_8 FILLER_80_462 ();
 sg13g2_decap_8 FILLER_80_469 ();
 sg13g2_decap_8 FILLER_80_476 ();
 sg13g2_decap_4 FILLER_80_483 ();
 sg13g2_fill_1 FILLER_80_487 ();
 sg13g2_fill_2 FILLER_80_537 ();
 sg13g2_fill_2 FILLER_80_574 ();
 sg13g2_decap_8 FILLER_80_592 ();
 sg13g2_decap_8 FILLER_80_599 ();
 sg13g2_decap_8 FILLER_80_606 ();
 sg13g2_decap_8 FILLER_80_613 ();
 sg13g2_decap_8 FILLER_80_620 ();
 sg13g2_decap_8 FILLER_80_627 ();
 sg13g2_decap_8 FILLER_80_634 ();
 sg13g2_decap_8 FILLER_80_641 ();
 sg13g2_decap_8 FILLER_80_648 ();
 sg13g2_decap_8 FILLER_80_655 ();
 sg13g2_decap_8 FILLER_80_662 ();
 sg13g2_decap_8 FILLER_80_669 ();
 sg13g2_decap_8 FILLER_80_676 ();
 sg13g2_decap_8 FILLER_80_683 ();
 sg13g2_decap_8 FILLER_80_690 ();
 sg13g2_decap_8 FILLER_80_697 ();
 sg13g2_decap_8 FILLER_80_704 ();
 sg13g2_decap_8 FILLER_80_711 ();
 sg13g2_decap_8 FILLER_80_718 ();
 sg13g2_decap_8 FILLER_80_725 ();
 sg13g2_decap_8 FILLER_80_732 ();
 sg13g2_decap_8 FILLER_80_739 ();
 sg13g2_decap_8 FILLER_80_746 ();
 sg13g2_decap_8 FILLER_80_753 ();
 sg13g2_decap_8 FILLER_80_760 ();
 sg13g2_decap_8 FILLER_80_767 ();
 sg13g2_decap_8 FILLER_80_774 ();
 sg13g2_decap_8 FILLER_80_781 ();
 sg13g2_decap_8 FILLER_80_788 ();
 sg13g2_decap_8 FILLER_80_795 ();
 sg13g2_decap_8 FILLER_80_802 ();
 sg13g2_decap_8 FILLER_80_809 ();
 sg13g2_decap_8 FILLER_80_816 ();
 sg13g2_decap_8 FILLER_80_823 ();
 sg13g2_decap_8 FILLER_80_830 ();
 sg13g2_decap_8 FILLER_80_837 ();
 sg13g2_decap_8 FILLER_80_844 ();
 sg13g2_decap_8 FILLER_80_851 ();
 sg13g2_decap_8 FILLER_80_858 ();
 sg13g2_decap_8 FILLER_80_865 ();
 sg13g2_decap_8 FILLER_80_872 ();
 sg13g2_decap_8 FILLER_80_879 ();
 sg13g2_decap_8 FILLER_80_886 ();
 sg13g2_decap_8 FILLER_80_893 ();
 sg13g2_decap_8 FILLER_80_900 ();
 sg13g2_decap_8 FILLER_80_907 ();
 sg13g2_decap_8 FILLER_80_914 ();
 sg13g2_decap_8 FILLER_80_921 ();
 sg13g2_decap_8 FILLER_80_928 ();
 sg13g2_decap_8 FILLER_80_935 ();
 sg13g2_decap_8 FILLER_80_942 ();
 sg13g2_decap_4 FILLER_80_949 ();
 sg13g2_fill_1 FILLER_80_1039 ();
 sg13g2_fill_2 FILLER_80_1110 ();
 sg13g2_fill_2 FILLER_80_1135 ();
 sg13g2_fill_2 FILLER_80_1195 ();
 sg13g2_fill_2 FILLER_80_1234 ();
 sg13g2_fill_1 FILLER_80_1265 ();
 sg13g2_fill_1 FILLER_80_1274 ();
 sg13g2_fill_1 FILLER_80_1314 ();
 sg13g2_fill_1 FILLER_80_1324 ();
 sg13g2_fill_2 FILLER_80_1360 ();
 sg13g2_fill_1 FILLER_80_1385 ();
 sg13g2_fill_2 FILLER_80_1414 ();
 sg13g2_fill_1 FILLER_80_1479 ();
 sg13g2_decap_8 FILLER_80_1508 ();
 sg13g2_decap_8 FILLER_80_1515 ();
 sg13g2_decap_8 FILLER_80_1522 ();
 sg13g2_decap_8 FILLER_80_1529 ();
 sg13g2_decap_8 FILLER_80_1536 ();
 sg13g2_decap_8 FILLER_80_1543 ();
 sg13g2_decap_8 FILLER_80_1550 ();
 sg13g2_decap_8 FILLER_80_1557 ();
 sg13g2_decap_8 FILLER_80_1569 ();
 sg13g2_fill_1 FILLER_80_1576 ();
 sg13g2_decap_8 FILLER_80_1644 ();
 sg13g2_decap_8 FILLER_80_1651 ();
 sg13g2_decap_8 FILLER_80_1658 ();
 sg13g2_decap_8 FILLER_80_1665 ();
 sg13g2_decap_8 FILLER_80_1672 ();
 sg13g2_decap_8 FILLER_80_1679 ();
 sg13g2_fill_1 FILLER_80_1690 ();
 sg13g2_fill_1 FILLER_80_1699 ();
 sg13g2_decap_8 FILLER_80_1704 ();
 sg13g2_decap_8 FILLER_80_1711 ();
 sg13g2_fill_2 FILLER_80_1718 ();
 sg13g2_fill_1 FILLER_80_1720 ();
 sg13g2_fill_2 FILLER_80_1756 ();
 sg13g2_fill_1 FILLER_80_1758 ();
 sg13g2_fill_1 FILLER_80_1789 ();
 sg13g2_fill_1 FILLER_80_1820 ();
 sg13g2_fill_2 FILLER_80_1831 ();
 sg13g2_fill_2 FILLER_80_1851 ();
 sg13g2_decap_8 FILLER_80_1870 ();
 sg13g2_decap_8 FILLER_80_1877 ();
 sg13g2_decap_8 FILLER_80_1884 ();
 sg13g2_decap_4 FILLER_80_1904 ();
 sg13g2_fill_1 FILLER_80_1916 ();
 sg13g2_fill_2 FILLER_80_1927 ();
 sg13g2_fill_1 FILLER_80_1929 ();
 sg13g2_decap_4 FILLER_80_1943 ();
 sg13g2_fill_2 FILLER_80_1947 ();
 sg13g2_decap_8 FILLER_80_1966 ();
 sg13g2_decap_4 FILLER_80_1973 ();
 sg13g2_fill_2 FILLER_80_1990 ();
 sg13g2_fill_1 FILLER_80_1992 ();
 sg13g2_decap_8 FILLER_80_2024 ();
 sg13g2_fill_2 FILLER_80_2031 ();
 sg13g2_fill_1 FILLER_80_2033 ();
 sg13g2_decap_8 FILLER_80_2056 ();
 sg13g2_decap_8 FILLER_80_2063 ();
 sg13g2_decap_8 FILLER_80_2070 ();
 sg13g2_decap_8 FILLER_80_2077 ();
 sg13g2_decap_8 FILLER_80_2084 ();
 sg13g2_decap_8 FILLER_80_2091 ();
 sg13g2_decap_8 FILLER_80_2098 ();
 sg13g2_decap_8 FILLER_80_2105 ();
 sg13g2_decap_8 FILLER_80_2112 ();
 sg13g2_decap_8 FILLER_80_2119 ();
 sg13g2_decap_8 FILLER_80_2126 ();
 sg13g2_decap_8 FILLER_80_2133 ();
 sg13g2_decap_8 FILLER_80_2140 ();
 sg13g2_decap_8 FILLER_80_2147 ();
 sg13g2_decap_8 FILLER_80_2154 ();
 sg13g2_decap_8 FILLER_80_2161 ();
 sg13g2_decap_8 FILLER_80_2168 ();
 sg13g2_decap_8 FILLER_80_2175 ();
 sg13g2_decap_8 FILLER_80_2182 ();
 sg13g2_decap_8 FILLER_80_2189 ();
 sg13g2_decap_8 FILLER_80_2196 ();
 sg13g2_decap_8 FILLER_80_2203 ();
 sg13g2_decap_8 FILLER_80_2210 ();
 sg13g2_decap_8 FILLER_80_2217 ();
 sg13g2_decap_8 FILLER_80_2224 ();
 sg13g2_decap_8 FILLER_80_2231 ();
 sg13g2_decap_8 FILLER_80_2238 ();
 sg13g2_decap_8 FILLER_80_2245 ();
 sg13g2_decap_8 FILLER_80_2252 ();
 sg13g2_decap_8 FILLER_80_2259 ();
 sg13g2_decap_8 FILLER_80_2266 ();
 sg13g2_decap_8 FILLER_80_2273 ();
 sg13g2_decap_8 FILLER_80_2280 ();
 sg13g2_decap_8 FILLER_80_2287 ();
 sg13g2_decap_8 FILLER_80_2294 ();
 sg13g2_decap_8 FILLER_80_2301 ();
 sg13g2_decap_8 FILLER_80_2308 ();
 sg13g2_decap_8 FILLER_80_2315 ();
 sg13g2_decap_8 FILLER_80_2322 ();
 sg13g2_decap_8 FILLER_80_2329 ();
 sg13g2_decap_8 FILLER_80_2336 ();
 sg13g2_decap_8 FILLER_80_2343 ();
 sg13g2_decap_8 FILLER_80_2350 ();
 sg13g2_decap_8 FILLER_80_2357 ();
 sg13g2_decap_8 FILLER_80_2364 ();
 sg13g2_decap_8 FILLER_80_2371 ();
 sg13g2_decap_8 FILLER_80_2378 ();
 sg13g2_decap_8 FILLER_80_2385 ();
 sg13g2_decap_8 FILLER_80_2392 ();
 sg13g2_decap_8 FILLER_80_2399 ();
 sg13g2_decap_8 FILLER_80_2406 ();
 sg13g2_decap_8 FILLER_80_2413 ();
 sg13g2_decap_8 FILLER_80_2420 ();
 sg13g2_decap_8 FILLER_80_2427 ();
 sg13g2_decap_8 FILLER_80_2434 ();
 sg13g2_decap_8 FILLER_80_2441 ();
 sg13g2_decap_8 FILLER_80_2448 ();
 sg13g2_decap_8 FILLER_80_2455 ();
 sg13g2_decap_8 FILLER_80_2462 ();
 sg13g2_decap_8 FILLER_80_2469 ();
 sg13g2_decap_8 FILLER_80_2476 ();
 sg13g2_decap_8 FILLER_80_2483 ();
 sg13g2_decap_8 FILLER_80_2490 ();
 sg13g2_decap_8 FILLER_80_2497 ();
 sg13g2_decap_8 FILLER_80_2504 ();
 sg13g2_decap_8 FILLER_80_2511 ();
 sg13g2_decap_8 FILLER_80_2518 ();
 sg13g2_decap_8 FILLER_80_2525 ();
 sg13g2_decap_8 FILLER_80_2532 ();
 sg13g2_decap_8 FILLER_80_2539 ();
 sg13g2_decap_8 FILLER_80_2546 ();
 sg13g2_decap_8 FILLER_80_2553 ();
 sg13g2_decap_8 FILLER_80_2560 ();
 sg13g2_decap_8 FILLER_80_2567 ();
 sg13g2_decap_8 FILLER_80_2574 ();
 sg13g2_decap_8 FILLER_80_2581 ();
 sg13g2_decap_8 FILLER_80_2588 ();
 sg13g2_decap_8 FILLER_80_2595 ();
 sg13g2_decap_8 FILLER_80_2602 ();
 sg13g2_decap_8 FILLER_80_2609 ();
 sg13g2_decap_8 FILLER_80_2616 ();
 sg13g2_decap_8 FILLER_80_2623 ();
 sg13g2_decap_8 FILLER_80_2630 ();
 sg13g2_decap_8 FILLER_80_2637 ();
 sg13g2_decap_8 FILLER_80_2644 ();
 sg13g2_decap_8 FILLER_80_2651 ();
 sg13g2_decap_8 FILLER_80_2658 ();
 sg13g2_decap_8 FILLER_80_2665 ();
 sg13g2_fill_2 FILLER_80_2672 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
 assign uo_out[3] = net18;
 assign uo_out[4] = net19;
 assign uo_out[5] = net20;
 assign uo_out[6] = net21;
 assign uo_out[7] = net22;
endmodule

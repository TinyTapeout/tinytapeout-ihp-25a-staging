module tt_um_gus16 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \GUScpu0.IR[0] ;
 wire \GUScpu0.IR[10] ;
 wire \GUScpu0.IR[11] ;
 wire \GUScpu0.IR[12] ;
 wire \GUScpu0.IR[13] ;
 wire \GUScpu0.IR[14] ;
 wire \GUScpu0.IR[15] ;
 wire \GUScpu0.IR[1] ;
 wire \GUScpu0.IR[2] ;
 wire \GUScpu0.IR[3] ;
 wire \GUScpu0.IR[4] ;
 wire \GUScpu0.IR[5] ;
 wire \GUScpu0.IR[6] ;
 wire \GUScpu0.IR[7] ;
 wire \GUScpu0.IR[8] ;
 wire \GUScpu0.IR[9] ;
 wire \GUScpu0.PC0[0] ;
 wire \GUScpu0.PC0[10] ;
 wire \GUScpu0.PC0[11] ;
 wire \GUScpu0.PC0[12] ;
 wire \GUScpu0.PC0[13] ;
 wire \GUScpu0.PC0[14] ;
 wire \GUScpu0.PC0[15] ;
 wire \GUScpu0.PC0[1] ;
 wire \GUScpu0.PC0[2] ;
 wire \GUScpu0.PC0[3] ;
 wire \GUScpu0.PC0[4] ;
 wire \GUScpu0.PC0[5] ;
 wire \GUScpu0.PC0[6] ;
 wire \GUScpu0.PC0[7] ;
 wire \GUScpu0.PC0[8] ;
 wire \GUScpu0.PC0[9] ;
 wire \GUScpu0.PC1[0] ;
 wire \GUScpu0.PC1[10] ;
 wire \GUScpu0.PC1[11] ;
 wire \GUScpu0.PC1[12] ;
 wire \GUScpu0.PC1[13] ;
 wire \GUScpu0.PC1[14] ;
 wire \GUScpu0.PC1[15] ;
 wire \GUScpu0.PC1[1] ;
 wire \GUScpu0.PC1[2] ;
 wire \GUScpu0.PC1[3] ;
 wire \GUScpu0.PC1[4] ;
 wire \GUScpu0.PC1[5] ;
 wire \GUScpu0.PC1[6] ;
 wire \GUScpu0.PC1[7] ;
 wire \GUScpu0.PC1[8] ;
 wire \GUScpu0.PC1[9] ;
 wire \GUScpu0.cdi[0] ;
 wire \GUScpu0.cdi[10] ;
 wire \GUScpu0.cdi[11] ;
 wire \GUScpu0.cdi[12] ;
 wire \GUScpu0.cdi[13] ;
 wire \GUScpu0.cdi[14] ;
 wire \GUScpu0.cdi[15] ;
 wire \GUScpu0.cdi[1] ;
 wire \GUScpu0.cdi[2] ;
 wire \GUScpu0.cdi[3] ;
 wire \GUScpu0.cdi[4] ;
 wire \GUScpu0.cdi[5] ;
 wire \GUScpu0.cdi[6] ;
 wire \GUScpu0.cdi[7] ;
 wire \GUScpu0.cdi[8] ;
 wire \GUScpu0.cdi[9] ;
 wire \GUScpu0.clk ;
 wire \GUScpu0.cv[0][0] ;
 wire \GUScpu0.cv[0][1] ;
 wire \GUScpu0.cv[1][0] ;
 wire \GUScpu0.cv[1][1] ;
 wire \GUScpu0.flag0[0] ;
 wire \GUScpu0.flag0[2] ;
 wire \GUScpu0.imode ;
 wire \GUScpu0.irqq0 ;
 wire \GUScpu0.opval ;
 wire \GUScpu0.opvali ;
 wire \GUScpu0.regs[0][0] ;
 wire \GUScpu0.regs[0][10] ;
 wire \GUScpu0.regs[0][11] ;
 wire \GUScpu0.regs[0][12] ;
 wire \GUScpu0.regs[0][13] ;
 wire \GUScpu0.regs[0][14] ;
 wire \GUScpu0.regs[0][15] ;
 wire \GUScpu0.regs[0][1] ;
 wire \GUScpu0.regs[0][2] ;
 wire \GUScpu0.regs[0][3] ;
 wire \GUScpu0.regs[0][4] ;
 wire \GUScpu0.regs[0][5] ;
 wire \GUScpu0.regs[0][6] ;
 wire \GUScpu0.regs[0][7] ;
 wire \GUScpu0.regs[0][8] ;
 wire \GUScpu0.regs[0][9] ;
 wire \GUScpu0.regs[1][0] ;
 wire \GUScpu0.regs[1][10] ;
 wire \GUScpu0.regs[1][11] ;
 wire \GUScpu0.regs[1][12] ;
 wire \GUScpu0.regs[1][13] ;
 wire \GUScpu0.regs[1][14] ;
 wire \GUScpu0.regs[1][15] ;
 wire \GUScpu0.regs[1][1] ;
 wire \GUScpu0.regs[1][2] ;
 wire \GUScpu0.regs[1][3] ;
 wire \GUScpu0.regs[1][4] ;
 wire \GUScpu0.regs[1][5] ;
 wire \GUScpu0.regs[1][6] ;
 wire \GUScpu0.regs[1][7] ;
 wire \GUScpu0.regs[1][8] ;
 wire \GUScpu0.regs[1][9] ;
 wire \GUScpu0.regs[2][0] ;
 wire \GUScpu0.regs[2][10] ;
 wire \GUScpu0.regs[2][11] ;
 wire \GUScpu0.regs[2][12] ;
 wire \GUScpu0.regs[2][13] ;
 wire \GUScpu0.regs[2][14] ;
 wire \GUScpu0.regs[2][15] ;
 wire \GUScpu0.regs[2][1] ;
 wire \GUScpu0.regs[2][2] ;
 wire \GUScpu0.regs[2][3] ;
 wire \GUScpu0.regs[2][4] ;
 wire \GUScpu0.regs[2][5] ;
 wire \GUScpu0.regs[2][6] ;
 wire \GUScpu0.regs[2][7] ;
 wire \GUScpu0.regs[2][8] ;
 wire \GUScpu0.regs[2][9] ;
 wire \GUScpu0.regs[3][0] ;
 wire \GUScpu0.regs[3][10] ;
 wire \GUScpu0.regs[3][11] ;
 wire \GUScpu0.regs[3][12] ;
 wire \GUScpu0.regs[3][13] ;
 wire \GUScpu0.regs[3][14] ;
 wire \GUScpu0.regs[3][15] ;
 wire \GUScpu0.regs[3][1] ;
 wire \GUScpu0.regs[3][2] ;
 wire \GUScpu0.regs[3][3] ;
 wire \GUScpu0.regs[3][4] ;
 wire \GUScpu0.regs[3][5] ;
 wire \GUScpu0.regs[3][6] ;
 wire \GUScpu0.regs[3][7] ;
 wire \GUScpu0.regs[3][8] ;
 wire \GUScpu0.regs[3][9] ;
 wire \GUScpu0.regs[4][0] ;
 wire \GUScpu0.regs[4][10] ;
 wire \GUScpu0.regs[4][11] ;
 wire \GUScpu0.regs[4][12] ;
 wire \GUScpu0.regs[4][13] ;
 wire \GUScpu0.regs[4][14] ;
 wire \GUScpu0.regs[4][15] ;
 wire \GUScpu0.regs[4][1] ;
 wire \GUScpu0.regs[4][2] ;
 wire \GUScpu0.regs[4][3] ;
 wire \GUScpu0.regs[4][4] ;
 wire \GUScpu0.regs[4][5] ;
 wire \GUScpu0.regs[4][6] ;
 wire \GUScpu0.regs[4][7] ;
 wire \GUScpu0.regs[4][8] ;
 wire \GUScpu0.regs[4][9] ;
 wire \GUScpu0.regs[5][0] ;
 wire \GUScpu0.regs[5][10] ;
 wire \GUScpu0.regs[5][11] ;
 wire \GUScpu0.regs[5][12] ;
 wire \GUScpu0.regs[5][13] ;
 wire \GUScpu0.regs[5][14] ;
 wire \GUScpu0.regs[5][15] ;
 wire \GUScpu0.regs[5][1] ;
 wire \GUScpu0.regs[5][2] ;
 wire \GUScpu0.regs[5][3] ;
 wire \GUScpu0.regs[5][4] ;
 wire \GUScpu0.regs[5][5] ;
 wire \GUScpu0.regs[5][6] ;
 wire \GUScpu0.regs[5][7] ;
 wire \GUScpu0.regs[5][8] ;
 wire \GUScpu0.regs[5][9] ;
 wire \GUScpu0.regs[6][0] ;
 wire \GUScpu0.regs[6][10] ;
 wire \GUScpu0.regs[6][11] ;
 wire \GUScpu0.regs[6][12] ;
 wire \GUScpu0.regs[6][13] ;
 wire \GUScpu0.regs[6][14] ;
 wire \GUScpu0.regs[6][15] ;
 wire \GUScpu0.regs[6][1] ;
 wire \GUScpu0.regs[6][2] ;
 wire \GUScpu0.regs[6][3] ;
 wire \GUScpu0.regs[6][4] ;
 wire \GUScpu0.regs[6][5] ;
 wire \GUScpu0.regs[6][6] ;
 wire \GUScpu0.regs[6][7] ;
 wire \GUScpu0.regs[6][8] ;
 wire \GUScpu0.regs[6][9] ;
 wire \GUScpu0.regs[7][0] ;
 wire \GUScpu0.regs[7][10] ;
 wire \GUScpu0.regs[7][11] ;
 wire \GUScpu0.regs[7][12] ;
 wire \GUScpu0.regs[7][13] ;
 wire \GUScpu0.regs[7][14] ;
 wire \GUScpu0.regs[7][15] ;
 wire \GUScpu0.regs[7][1] ;
 wire \GUScpu0.regs[7][2] ;
 wire \GUScpu0.regs[7][3] ;
 wire \GUScpu0.regs[7][4] ;
 wire \GUScpu0.regs[7][5] ;
 wire \GUScpu0.regs[7][6] ;
 wire \GUScpu0.regs[7][7] ;
 wire \GUScpu0.regs[7][8] ;
 wire \GUScpu0.regs[7][9] ;
 wire \GUScpu0.zn[1][0] ;
 wire \GUScpu0.zn[1][1] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire clk_regs;
 wire net18;
 wire \ckd[0] ;
 wire \ckd[1] ;
 wire gpo;
 wire \irqen[0] ;
 wire \irqen[1] ;
 wire \irqen[2] ;
 wire \irqen[3] ;
 wire \irqen[4] ;
 wire \pwmbuf[0] ;
 wire \pwmbuf[1] ;
 wire \pwmbuf[2] ;
 wire \pwmbuf[3] ;
 wire \pwmbuf[4] ;
 wire \pwmbuf[5] ;
 wire \pwmbuf[6] ;
 wire \pwmbuf[7] ;
 wire \pwmc[0] ;
 wire \pwmc[1] ;
 wire \pwmc[2] ;
 wire \pwmc[3] ;
 wire \pwmc[4] ;
 wire \pwmc[5] ;
 wire \pwmc[6] ;
 wire \pwmc[7] ;
 wire \pwmhold[0] ;
 wire \pwmhold[1] ;
 wire \pwmhold[2] ;
 wire \pwmhold[3] ;
 wire \pwmhold[4] ;
 wire \pwmhold[5] ;
 wire \pwmhold[6] ;
 wire \pwmhold[7] ;
 wire pwmirq;
 wire pwmout;
 wire sdty;
 wire txd;
 wire \uart0.q[0] ;
 wire \uart0.q[1] ;
 wire \uart0.q[2] ;
 wire \uart0.q[3] ;
 wire \uart0.q[4] ;
 wire \uart0.q[5] ;
 wire \uart0.q[6] ;
 wire \uart0.q[7] ;
 wire \uart0.rxdiv[0] ;
 wire \uart0.rxdiv[1] ;
 wire \uart0.rxdiv[2] ;
 wire \uart0.rxdiv[3] ;
 wire \uart0.rxdiv[4] ;
 wire \uart0.rxdiv[5] ;
 wire \uart0.rxoverr ;
 wire \uart0.rxreg[0] ;
 wire \uart0.rxreg[1] ;
 wire \uart0.rxvalid ;
 wire \uart0.txbitcnt[0] ;
 wire \uart0.txbitcnt[1] ;
 wire \uart0.txbitcnt[2] ;
 wire \uart0.txbitcnt[3] ;
 wire \uart0.txdiv[0] ;
 wire \uart0.txdiv[1] ;
 wire \uart0.txdiv[2] ;
 wire \uart0.txdiv[3] ;
 wire \uart0.txdiv[4] ;
 wire \uart0.txdiv[5] ;
 wire \uart0.txsh[1] ;
 wire \uart0.txsh[2] ;
 wire \uart0.txsh[3] ;
 wire \uart0.txsh[4] ;
 wire \uart0.txsh[5] ;
 wire \uart0.txsh[6] ;
 wire \uart0.txsh[7] ;
 wire \uart0.txsh[8] ;
 wire \uart0.urxbuffer[8] ;
 wire \uart0.urxsh[0] ;
 wire \uart0.urxsh[1] ;
 wire \uart0.urxsh[2] ;
 wire \uart0.urxsh[3] ;
 wire \uart0.urxsh[4] ;
 wire \uart0.urxsh[5] ;
 wire \uart0.urxsh[6] ;
 wire \uart0.urxsh[7] ;
 wire \uart0.urxsh[8] ;
 wire \uart0.urxsh[9] ;
 wire \xdi[0] ;
 wire \xdi[1] ;
 wire \xdi[2] ;
 wire \xdi[3] ;
 wire \xdi[4] ;
 wire \xdi[5] ;
 wire \xdi[6] ;
 wire \xdi[7] ;
 wire xlah;
 wire xlal;
 wire xoeb;
 wire xweb;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_1_0__leaf_clk_regs;
 wire clknet_1_1__leaf_clk_regs;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;

 sg13g2_inv_1 _2028_ (.Y(_1460_),
    .A(\uart0.rxvalid ));
 sg13g2_inv_1 _2029_ (.Y(_1461_),
    .A(\uart0.txbitcnt[3] ));
 sg13g2_inv_1 _2030_ (.Y(_1462_),
    .A(pwmirq));
 sg13g2_inv_1 _2031_ (.Y(_1463_),
    .A(pwmout));
 sg13g2_inv_1 _2032_ (.Y(_1464_),
    .A(\pwmbuf[4] ));
 sg13g2_inv_1 _2033_ (.Y(_1465_),
    .A(\pwmbuf[1] ));
 sg13g2_inv_1 _2034_ (.Y(_1466_),
    .A(\pwmc[3] ));
 sg13g2_inv_1 _2035_ (.Y(_1467_),
    .A(\pwmc[2] ));
 sg13g2_inv_1 _2036_ (.Y(_1468_),
    .A(\ckd[1] ));
 sg13g2_inv_1 _2037_ (.Y(_1469_),
    .A(net880));
 sg13g2_inv_1 _2038_ (.Y(_1470_),
    .A(\GUScpu0.IR[15] ));
 sg13g2_inv_1 _2039_ (.Y(_1471_),
    .A(\GUScpu0.opval ));
 sg13g2_inv_4 _2040_ (.A(net870),
    .Y(_1472_));
 sg13g2_inv_1 _2041_ (.Y(_1473_),
    .A(_0087_));
 sg13g2_inv_1 _2042_ (.Y(_1474_),
    .A(_0090_));
 sg13g2_inv_2 _2043_ (.Y(_1475_),
    .A(_0089_));
 sg13g2_inv_1 _2044_ (.Y(_1476_),
    .A(_0095_));
 sg13g2_inv_1 _2045_ (.Y(_1477_),
    .A(net884));
 sg13g2_inv_1 _2046_ (.Y(_1478_),
    .A(\GUScpu0.IR[7] ));
 sg13g2_inv_1 _2047_ (.Y(_1479_),
    .A(_0099_));
 sg13g2_inv_1 _2048_ (.Y(_1480_),
    .A(_0100_));
 sg13g2_inv_1 _2049_ (.Y(_1481_),
    .A(_0108_));
 sg13g2_inv_1 _2050_ (.Y(_1482_),
    .A(_0112_));
 sg13g2_inv_1 _2051_ (.Y(_1483_),
    .A(_0115_));
 sg13g2_inv_1 _2052_ (.Y(_1484_),
    .A(_0124_));
 sg13g2_inv_1 _2053_ (.Y(_1485_),
    .A(_0128_));
 sg13g2_inv_1 _2054_ (.Y(_1486_),
    .A(_0131_));
 sg13g2_inv_1 _2055_ (.Y(_1487_),
    .A(_0132_));
 sg13g2_inv_1 _2056_ (.Y(_1488_),
    .A(_0137_));
 sg13g2_inv_1 _2057_ (.Y(_1489_),
    .A(_0141_));
 sg13g2_inv_1 _2058_ (.Y(_1490_),
    .A(_0145_));
 sg13g2_inv_1 _2059_ (.Y(_1491_),
    .A(_0153_));
 sg13g2_inv_1 _2060_ (.Y(_1492_),
    .A(_0156_));
 sg13g2_inv_1 _2061_ (.Y(_1493_),
    .A(_0047_));
 sg13g2_inv_1 _2062_ (.Y(_1494_),
    .A(_0055_));
 sg13g2_inv_1 _2063_ (.Y(_1495_),
    .A(_0063_));
 sg13g2_inv_1 _2064_ (.Y(_1496_),
    .A(_0068_));
 sg13g2_inv_1 _2065_ (.Y(_1497_),
    .A(_0077_));
 sg13g2_inv_1 _2066_ (.Y(_1498_),
    .A(\uart0.rxdiv[1] ));
 sg13g2_inv_1 _2067_ (.Y(_1499_),
    .A(net221));
 sg13g2_inv_1 _2068_ (.Y(_1500_),
    .A(net226));
 sg13g2_inv_1 _2069_ (.Y(_1501_),
    .A(\irqen[3] ));
 sg13g2_inv_1 _2070_ (.Y(_1502_),
    .A(\xdi[5] ));
 sg13g2_inv_1 _2071_ (.Y(_1503_),
    .A(net14));
 sg13g2_inv_1 _2072_ (.Y(_1504_),
    .A(net15));
 sg13g2_nor2b_1 _2073_ (.A(net880),
    .B_N(net882),
    .Y(_1505_));
 sg13g2_nand2b_2 _2074_ (.Y(_1506_),
    .B(net882),
    .A_N(net881));
 sg13g2_nor2b_1 _2075_ (.A(\GUScpu0.IR[15] ),
    .B_N(\GUScpu0.IR[14] ),
    .Y(_1507_));
 sg13g2_nand3b_1 _2076_ (.B(net879),
    .C(\GUScpu0.IR[14] ),
    .Y(_1508_),
    .A_N(\GUScpu0.IR[15] ));
 sg13g2_nor2_2 _2077_ (.A(_1506_),
    .B(_1508_),
    .Y(_1509_));
 sg13g2_nor3_1 _2078_ (.A(_1471_),
    .B(_1506_),
    .C(_1508_),
    .Y(_1510_));
 sg13g2_nand2_2 _2079_ (.Y(_1511_),
    .A(\GUScpu0.opval ),
    .B(_1509_));
 sg13g2_nor2_2 _2080_ (.A(net880),
    .B(net882),
    .Y(_1512_));
 sg13g2_nand2_1 _2081_ (.Y(_1513_),
    .A(\GUScpu0.IR[14] ),
    .B(_0084_));
 sg13g2_nand3_1 _2082_ (.B(net879),
    .C(_0084_),
    .A(\GUScpu0.IR[14] ),
    .Y(_1514_));
 sg13g2_nor3_2 _2083_ (.A(net881),
    .B(net882),
    .C(_1514_),
    .Y(_1515_));
 sg13g2_nor4_2 _2084_ (.A(net881),
    .B(net882),
    .C(_0083_),
    .Y(_1516_),
    .D(_1514_));
 sg13g2_nor2_1 _2085_ (.A(net865),
    .B(_1516_),
    .Y(_1517_));
 sg13g2_or2_2 _2086_ (.X(_1518_),
    .B(_1516_),
    .A(net865));
 sg13g2_and2_1 _2087_ (.A(net880),
    .B(net882),
    .X(_1519_));
 sg13g2_nand2_2 _2088_ (.Y(_1520_),
    .A(net880),
    .B(net882));
 sg13g2_nand3b_1 _2089_ (.B(_1507_),
    .C(_1519_),
    .Y(_1521_),
    .A_N(net879));
 sg13g2_and2_1 _2090_ (.A(_1477_),
    .B(_1507_),
    .X(_1522_));
 sg13g2_nor4_1 _2091_ (.A(net879),
    .B(\GUScpu0.IR[6] ),
    .C(_1478_),
    .D(_1520_),
    .Y(_1523_));
 sg13g2_nor2b_1 _2092_ (.A(\GUScpu0.IR[5] ),
    .B_N(_1523_),
    .Y(_1524_));
 sg13g2_nor2b_1 _2093_ (.A(\GUScpu0.IR[0] ),
    .B_N(_1507_),
    .Y(_1525_));
 sg13g2_and2_1 _2094_ (.A(_1524_),
    .B(_1525_),
    .X(_1526_));
 sg13g2_o21ai_1 _2095_ (.B1(_1524_),
    .Y(_1527_),
    .A1(_1522_),
    .A2(_1525_));
 sg13g2_o21ai_1 _2096_ (.B1(_1527_),
    .Y(_1528_),
    .A1(\GUScpu0.IR[7] ),
    .A2(_1521_));
 sg13g2_nor2_2 _2097_ (.A(net884),
    .B(\GUScpu0.IR[0] ),
    .Y(_1529_));
 sg13g2_nand2_1 _2098_ (.Y(_1530_),
    .A(\GUScpu0.IR[5] ),
    .B(\GUScpu0.IR[6] ));
 sg13g2_nand3_1 _2099_ (.B(\GUScpu0.IR[6] ),
    .C(\GUScpu0.IR[7] ),
    .A(\GUScpu0.IR[5] ),
    .Y(_1531_));
 sg13g2_nor4_1 _2100_ (.A(net884),
    .B(\GUScpu0.IR[0] ),
    .C(_1521_),
    .D(_1531_),
    .Y(_1532_));
 sg13g2_nor2_2 _2101_ (.A(net879),
    .B(_1513_),
    .Y(_1533_));
 sg13g2_inv_1 _2102_ (.Y(_1534_),
    .A(_1533_));
 sg13g2_nor4_1 _2103_ (.A(_1477_),
    .B(_1520_),
    .C(_1531_),
    .D(_1534_),
    .Y(_1535_));
 sg13g2_or2_1 _2104_ (.X(_1536_),
    .B(_1535_),
    .A(_1532_));
 sg13g2_nor2b_1 _2105_ (.A(\GUScpu0.IR[14] ),
    .B_N(_0084_),
    .Y(_1537_));
 sg13g2_nor2b_2 _2106_ (.A(net879),
    .B_N(_1537_),
    .Y(_1538_));
 sg13g2_and2_1 _2107_ (.A(_1505_),
    .B(_1538_),
    .X(_1539_));
 sg13g2_and2_1 _2108_ (.A(\GUScpu0.IR[0] ),
    .B(_1539_),
    .X(_1540_));
 sg13g2_and2_1 _2109_ (.A(net879),
    .B(_1537_),
    .X(_1541_));
 sg13g2_nand3b_1 _2110_ (.B(net879),
    .C(_0084_),
    .Y(_1542_),
    .A_N(\GUScpu0.IR[14] ));
 sg13g2_nor2_1 _2111_ (.A(_1520_),
    .B(_1542_),
    .Y(_1543_));
 sg13g2_nor2_1 _2112_ (.A(_1469_),
    .B(net882),
    .Y(_1544_));
 sg13g2_and2_1 _2113_ (.A(_1533_),
    .B(_1544_),
    .X(_1545_));
 sg13g2_nor3_1 _2114_ (.A(_1540_),
    .B(_1543_),
    .C(_1545_),
    .Y(_1546_));
 sg13g2_a22oi_1 _2115_ (.Y(_1547_),
    .B1(_1541_),
    .B2(_1544_),
    .A2(_1539_),
    .A1(_1529_));
 sg13g2_and3_1 _2116_ (.X(_1548_),
    .A(\GUScpu0.IR[5] ),
    .B(_1522_),
    .C(_1523_));
 sg13g2_nand2b_1 _2117_ (.Y(_1549_),
    .B(_1548_),
    .A_N(\GUScpu0.IR[0] ));
 sg13g2_nor2_1 _2118_ (.A(_1528_),
    .B(_1536_),
    .Y(_1550_));
 sg13g2_nand4_1 _2119_ (.B(_1547_),
    .C(_1549_),
    .A(_1546_),
    .Y(_1551_),
    .D(_1550_));
 sg13g2_inv_1 _2120_ (.Y(_1552_),
    .A(net766));
 sg13g2_a22oi_1 _2121_ (.Y(_1553_),
    .B1(_1539_),
    .B2(net884),
    .A2(_1533_),
    .A1(_1512_));
 sg13g2_and2_2 _2122_ (.A(_1547_),
    .B(_1553_),
    .X(_1554_));
 sg13g2_nor2b_1 _2123_ (.A(net766),
    .B_N(_1554_),
    .Y(_1555_));
 sg13g2_nand2_1 _2124_ (.Y(_1556_),
    .A(_1552_),
    .B(_1554_));
 sg13g2_a22oi_1 _2125_ (.Y(_1557_),
    .B1(_1541_),
    .B2(_1520_),
    .A2(_1538_),
    .A1(net880));
 sg13g2_or2_1 _2126_ (.X(_1558_),
    .B(_1508_),
    .A(_1469_));
 sg13g2_and2_1 _2127_ (.A(_1470_),
    .B(_1558_),
    .X(_1559_));
 sg13g2_o21ai_1 _2128_ (.B1(_1470_),
    .Y(_1560_),
    .A1(_1469_),
    .A2(_1508_));
 sg13g2_nor3_2 _2129_ (.A(_1509_),
    .B(_1515_),
    .C(net862),
    .Y(_1561_));
 sg13g2_a21oi_1 _2130_ (.A1(_1520_),
    .A2(_1533_),
    .Y(_1562_),
    .B1(_1543_));
 sg13g2_and3_2 _2131_ (.X(_1563_),
    .A(_1557_),
    .B(_1561_),
    .C(_1562_));
 sg13g2_nand3_1 _2132_ (.B(_1561_),
    .C(_1562_),
    .A(_1557_),
    .Y(_1564_));
 sg13g2_nor3_2 _2133_ (.A(_0083_),
    .B(net857),
    .C(net863),
    .Y(_1565_));
 sg13g2_nand2_2 _2134_ (.Y(_1566_),
    .A(net830),
    .B(_1565_));
 sg13g2_mux2_2 _2135_ (.A0(_1473_),
    .A1(_1479_),
    .S(_1566_),
    .X(_1567_));
 sg13g2_mux2_1 _2136_ (.A0(_0087_),
    .A1(_0099_),
    .S(_1566_),
    .X(_1568_));
 sg13g2_mux2_1 _2137_ (.A0(_0089_),
    .A1(_0100_),
    .S(_1566_),
    .X(_1569_));
 sg13g2_mux2_1 _2138_ (.A0(_1475_),
    .A1(_1480_),
    .S(_1566_),
    .X(_1570_));
 sg13g2_mux2_1 _2139_ (.A0(_0074_),
    .A1(_0073_),
    .S(net790),
    .X(_1571_));
 sg13g2_nand2b_1 _2140_ (.Y(_1572_),
    .B(_1566_),
    .A_N(_0101_));
 sg13g2_mux2_1 _2141_ (.A0(net883),
    .A1(_0101_),
    .S(_1566_),
    .X(_1573_));
 sg13g2_o21ai_1 _2142_ (.B1(_1572_),
    .Y(_1574_),
    .A1(net883),
    .A2(_1566_));
 sg13g2_nor2_1 _2143_ (.A(_0076_),
    .B(net790),
    .Y(_1575_));
 sg13g2_o21ai_1 _2144_ (.B1(net780),
    .Y(_1576_),
    .A1(_0075_),
    .A2(net799));
 sg13g2_o21ai_1 _2145_ (.B1(net764),
    .Y(_1577_),
    .A1(_1575_),
    .A2(_1576_));
 sg13g2_a21oi_1 _2146_ (.A1(net783),
    .A2(_1571_),
    .Y(_1578_),
    .B1(_1577_));
 sg13g2_mux2_1 _2147_ (.A0(_0070_),
    .A1(_0069_),
    .S(net791),
    .X(_1579_));
 sg13g2_nor2_1 _2148_ (.A(_0072_),
    .B(net790),
    .Y(_1580_));
 sg13g2_o21ai_1 _2149_ (.B1(net780),
    .Y(_1581_),
    .A1(_0071_),
    .A2(net799));
 sg13g2_o21ai_1 _2150_ (.B1(net775),
    .Y(_1582_),
    .A1(_1580_),
    .A2(_1581_));
 sg13g2_a21oi_1 _2151_ (.A1(net783),
    .A2(_1579_),
    .Y(_1583_),
    .B1(_1582_));
 sg13g2_nor3_2 _2152_ (.A(net863),
    .B(_1578_),
    .C(_1583_),
    .Y(_1584_));
 sg13g2_nand3b_1 _2153_ (.B(_1561_),
    .C(_1562_),
    .Y(_1585_),
    .A_N(_1536_));
 sg13g2_inv_1 _2154_ (.Y(_1586_),
    .A(_1585_));
 sg13g2_nand3_1 _2155_ (.B(_1512_),
    .C(_1538_),
    .A(net884),
    .Y(_1587_));
 sg13g2_nand3_1 _2156_ (.B(_1512_),
    .C(_1538_),
    .A(\GUScpu0.IR[0] ),
    .Y(_1588_));
 sg13g2_nor2b_1 _2157_ (.A(_1539_),
    .B_N(_1557_),
    .Y(_1589_));
 sg13g2_nand3_1 _2158_ (.B(_1588_),
    .C(_1589_),
    .A(_1587_),
    .Y(_1590_));
 sg13g2_or4_1 _2159_ (.A(_1528_),
    .B(_1548_),
    .C(_1585_),
    .D(_1590_),
    .X(_1591_));
 sg13g2_a21oi_1 _2160_ (.A1(_1512_),
    .A2(_1533_),
    .Y(_1592_),
    .B1(_1543_));
 sg13g2_o21ai_1 _2161_ (.B1(_1592_),
    .Y(_1593_),
    .A1(_1506_),
    .A2(_1534_));
 sg13g2_nor2_1 _2162_ (.A(_1590_),
    .B(_1593_),
    .Y(_1594_));
 sg13g2_and3_2 _2163_ (.X(_1595_),
    .A(_1561_),
    .B(_1591_),
    .C(_1594_));
 sg13g2_nand3_1 _2164_ (.B(_1591_),
    .C(_1594_),
    .A(_1561_),
    .Y(_1596_));
 sg13g2_mux2_2 _2165_ (.A0(\GUScpu0.PC0[15] ),
    .A1(\GUScpu0.PC1[15] ),
    .S(net875),
    .X(_1597_));
 sg13g2_o21ai_1 _2166_ (.B1(net757),
    .Y(_1598_),
    .A1(net855),
    .A2(_1597_));
 sg13g2_o21ai_1 _2167_ (.B1(_1505_),
    .Y(_1599_),
    .A1(_1533_),
    .A2(_1541_));
 sg13g2_nand2_1 _2168_ (.Y(_1600_),
    .A(_1588_),
    .B(_1599_));
 sg13g2_a221oi_1 _2169_ (.B2(net884),
    .C1(_1548_),
    .B1(_1540_),
    .A1(_1519_),
    .Y(_1601_),
    .A2(_1538_));
 sg13g2_nand2b_2 _2170_ (.Y(_1602_),
    .B(_1601_),
    .A_N(_1600_));
 sg13g2_or2_1 _2171_ (.X(_1603_),
    .B(_1558_),
    .A(_0083_));
 sg13g2_nand2_2 _2172_ (.Y(_1604_),
    .A(_0084_),
    .B(net848));
 sg13g2_a21oi_2 _2173_ (.B1(net832),
    .Y(_1605_),
    .A2(_1604_),
    .A1(\GUScpu0.IR[11] ));
 sg13g2_nand2_1 _2174_ (.Y(_1606_),
    .A(_1473_),
    .B(net866));
 sg13g2_mux2_1 _2175_ (.A0(_0088_),
    .A1(_0087_),
    .S(net866),
    .X(_1607_));
 sg13g2_o21ai_1 _2176_ (.B1(_1606_),
    .Y(_1608_),
    .A1(_0088_),
    .A2(net865));
 sg13g2_nor2_1 _2177_ (.A(_0090_),
    .B(net865),
    .Y(_1609_));
 sg13g2_a21oi_1 _2178_ (.A1(_1475_),
    .A2(net865),
    .Y(_1610_),
    .B1(_1609_));
 sg13g2_mux2_2 _2179_ (.A0(_1474_),
    .A1(_1475_),
    .S(net865),
    .X(_1611_));
 sg13g2_mux2_1 _2180_ (.A0(_0074_),
    .A1(_0073_),
    .S(net843),
    .X(_1612_));
 sg13g2_o21ai_1 _2181_ (.B1(net837),
    .Y(_1613_),
    .A1(_0076_),
    .A2(net843));
 sg13g2_inv_1 _2182_ (.Y(_1614_),
    .A(_1613_));
 sg13g2_o21ai_1 _2183_ (.B1(_1614_),
    .Y(_1615_),
    .A1(_0075_),
    .A2(net828));
 sg13g2_nor2_1 _2184_ (.A(_0094_),
    .B(net865),
    .Y(_1616_));
 sg13g2_nand2b_1 _2185_ (.Y(_1617_),
    .B(net865),
    .A_N(net883));
 sg13g2_nor2b_1 _2186_ (.A(_1616_),
    .B_N(_1617_),
    .Y(_1618_));
 sg13g2_nand2b_2 _2187_ (.Y(_1619_),
    .B(_1617_),
    .A_N(_1616_));
 sg13g2_a21oi_1 _2188_ (.A1(net826),
    .A2(_1612_),
    .Y(_1620_),
    .B1(net823));
 sg13g2_mux4_1 _2189_ (.S0(net843),
    .A0(_0070_),
    .A1(_0069_),
    .A2(_0072_),
    .A3(_0071_),
    .S1(net837),
    .X(_1621_));
 sg13g2_inv_1 _2190_ (.Y(_1622_),
    .A(_1621_));
 sg13g2_a22oi_1 _2191_ (.Y(_1623_),
    .B1(_1622_),
    .B2(net823),
    .A2(_1620_),
    .A1(_1615_));
 sg13g2_a21oi_1 _2192_ (.A1(net832),
    .A2(_1623_),
    .Y(_1624_),
    .B1(_1605_));
 sg13g2_xnor2_1 _2193_ (.Y(_1625_),
    .A(net774),
    .B(_1624_));
 sg13g2_nor3_2 _2194_ (.A(_1584_),
    .B(_1598_),
    .C(_1625_),
    .Y(_1626_));
 sg13g2_inv_1 _2195_ (.Y(_1627_),
    .A(_1626_));
 sg13g2_o21ai_1 _2196_ (.B1(_1625_),
    .Y(_1628_),
    .A1(_1584_),
    .A2(_1598_));
 sg13g2_inv_1 _2197_ (.Y(_1629_),
    .A(_1628_));
 sg13g2_nand2_1 _2198_ (.Y(_1630_),
    .A(_1627_),
    .B(_1628_));
 sg13g2_nor2_1 _2199_ (.A(_0065_),
    .B(net800),
    .Y(_1631_));
 sg13g2_o21ai_1 _2200_ (.B1(net785),
    .Y(_1632_),
    .A1(_0066_),
    .A2(net796));
 sg13g2_nand2_1 _2201_ (.Y(_1633_),
    .A(_0067_),
    .B(net796));
 sg13g2_o21ai_1 _2202_ (.B1(_1633_),
    .Y(_1634_),
    .A1(_1496_),
    .A2(net796));
 sg13g2_a21oi_1 _2203_ (.A1(net779),
    .A2(_1634_),
    .Y(_1635_),
    .B1(net776));
 sg13g2_o21ai_1 _2204_ (.B1(_1635_),
    .Y(_1636_),
    .A1(_1631_),
    .A2(_1632_));
 sg13g2_mux2_1 _2205_ (.A0(_0062_),
    .A1(_0061_),
    .S(net796),
    .X(_1637_));
 sg13g2_a21oi_1 _2206_ (.A1(_1495_),
    .A2(net796),
    .Y(_1638_),
    .B1(net785));
 sg13g2_o21ai_1 _2207_ (.B1(_1638_),
    .Y(_1639_),
    .A1(_0064_),
    .A2(net796));
 sg13g2_a21oi_1 _2208_ (.A1(net785),
    .A2(_1637_),
    .Y(_1640_),
    .B1(_1574_));
 sg13g2_a21oi_1 _2209_ (.A1(_1639_),
    .A2(_1640_),
    .Y(_1641_),
    .B1(net864));
 sg13g2_mux2_2 _2210_ (.A0(\GUScpu0.PC0[14] ),
    .A1(\GUScpu0.PC1[14] ),
    .S(net876),
    .X(_1642_));
 sg13g2_o21ai_1 _2211_ (.B1(_1596_),
    .Y(_1643_),
    .A1(net856),
    .A2(_1642_));
 sg13g2_a21oi_1 _2212_ (.A1(_1636_),
    .A2(_1641_),
    .Y(_1644_),
    .B1(_1643_));
 sg13g2_mux2_1 _2213_ (.A0(_0066_),
    .A1(_0065_),
    .S(net846),
    .X(_1645_));
 sg13g2_a21oi_1 _2214_ (.A1(_1496_),
    .A2(net829),
    .Y(_1646_),
    .B1(net827));
 sg13g2_o21ai_1 _2215_ (.B1(_1646_),
    .Y(_1647_),
    .A1(_0067_),
    .A2(net829));
 sg13g2_a21oi_1 _2216_ (.A1(net827),
    .A2(_1645_),
    .Y(_1648_),
    .B1(net825));
 sg13g2_mux4_1 _2217_ (.S0(net846),
    .A0(_0062_),
    .A1(_0061_),
    .A2(_0064_),
    .A3(_0063_),
    .S1(net839),
    .X(_1649_));
 sg13g2_inv_1 _2218_ (.Y(_1650_),
    .A(_1649_));
 sg13g2_a22oi_1 _2219_ (.Y(_1651_),
    .B1(_1650_),
    .B2(net825),
    .A2(_1648_),
    .A1(_1647_));
 sg13g2_a21oi_1 _2220_ (.A1(_1563_),
    .A2(_1651_),
    .Y(_1652_),
    .B1(_1605_));
 sg13g2_xnor2_1 _2221_ (.Y(_1653_),
    .A(_1602_),
    .B(_1652_));
 sg13g2_nor2b_1 _2222_ (.A(_1653_),
    .B_N(_1644_),
    .Y(_1654_));
 sg13g2_inv_1 _2223_ (.Y(_1655_),
    .A(_1654_));
 sg13g2_xor2_1 _2224_ (.B(_1653_),
    .A(_1644_),
    .X(_1656_));
 sg13g2_inv_1 _2225_ (.Y(_1657_),
    .A(_1656_));
 sg13g2_nor2_1 _2226_ (.A(_0057_),
    .B(net801),
    .Y(_1658_));
 sg13g2_o21ai_1 _2227_ (.B1(net784),
    .Y(_1659_),
    .A1(_0058_),
    .A2(net796));
 sg13g2_mux2_1 _2228_ (.A0(_0060_),
    .A1(_0059_),
    .S(net794),
    .X(_1660_));
 sg13g2_a21oi_1 _2229_ (.A1(net779),
    .A2(_1660_),
    .Y(_1661_),
    .B1(net776));
 sg13g2_o21ai_1 _2230_ (.B1(_1661_),
    .Y(_1662_),
    .A1(_1658_),
    .A2(_1659_));
 sg13g2_mux2_1 _2231_ (.A0(_0054_),
    .A1(_0053_),
    .S(net793),
    .X(_1663_));
 sg13g2_a21oi_1 _2232_ (.A1(_1494_),
    .A2(net794),
    .Y(_1664_),
    .B1(net784));
 sg13g2_o21ai_1 _2233_ (.B1(_1664_),
    .Y(_1665_),
    .A1(_0056_),
    .A2(net794));
 sg13g2_a21oi_1 _2234_ (.A1(net785),
    .A2(_1663_),
    .Y(_1666_),
    .B1(net765));
 sg13g2_a21oi_1 _2235_ (.A1(_1665_),
    .A2(_1666_),
    .Y(_1667_),
    .B1(net864));
 sg13g2_mux2_2 _2236_ (.A0(\GUScpu0.PC0[13] ),
    .A1(\GUScpu0.PC1[13] ),
    .S(net876),
    .X(_1668_));
 sg13g2_o21ai_1 _2237_ (.B1(_1596_),
    .Y(_1669_),
    .A1(net856),
    .A2(_1668_));
 sg13g2_a21oi_1 _2238_ (.A1(_1662_),
    .A2(_1667_),
    .Y(_1670_),
    .B1(_1669_));
 sg13g2_mux2_1 _2239_ (.A0(_0058_),
    .A1(_0057_),
    .S(net846),
    .X(_1671_));
 sg13g2_o21ai_1 _2240_ (.B1(net838),
    .Y(_1672_),
    .A1(_0060_),
    .A2(net846));
 sg13g2_inv_1 _2241_ (.Y(_1673_),
    .A(_1672_));
 sg13g2_o21ai_1 _2242_ (.B1(_1673_),
    .Y(_1674_),
    .A1(_0059_),
    .A2(net829));
 sg13g2_a21oi_1 _2243_ (.A1(net827),
    .A2(_1671_),
    .Y(_1675_),
    .B1(net824));
 sg13g2_mux4_1 _2244_ (.S0(net845),
    .A0(_0054_),
    .A1(_0053_),
    .A2(_0056_),
    .A3(_0055_),
    .S1(net838),
    .X(_1676_));
 sg13g2_inv_1 _2245_ (.Y(_1677_),
    .A(_1676_));
 sg13g2_a22oi_1 _2246_ (.Y(_1678_),
    .B1(_1677_),
    .B2(net824),
    .A2(_1675_),
    .A1(_1674_));
 sg13g2_a21oi_1 _2247_ (.A1(net832),
    .A2(_1678_),
    .Y(_1679_),
    .B1(_1605_));
 sg13g2_xor2_1 _2248_ (.B(_1679_),
    .A(net774),
    .X(_1680_));
 sg13g2_and2_1 _2249_ (.A(_1670_),
    .B(_1680_),
    .X(_1681_));
 sg13g2_xor2_1 _2250_ (.B(_1680_),
    .A(_1670_),
    .X(_1682_));
 sg13g2_nor2_1 _2251_ (.A(_0049_),
    .B(net800),
    .Y(_1683_));
 sg13g2_o21ai_1 _2252_ (.B1(net784),
    .Y(_1684_),
    .A1(_0050_),
    .A2(net794));
 sg13g2_mux2_1 _2253_ (.A0(_0052_),
    .A1(_0051_),
    .S(net793),
    .X(_1685_));
 sg13g2_a21oi_1 _2254_ (.A1(net779),
    .A2(_1685_),
    .Y(_1686_),
    .B1(net776));
 sg13g2_o21ai_1 _2255_ (.B1(_1686_),
    .Y(_1687_),
    .A1(_1683_),
    .A2(_1684_));
 sg13g2_mux2_1 _2256_ (.A0(_0046_),
    .A1(_0045_),
    .S(net793),
    .X(_1688_));
 sg13g2_a21oi_1 _2257_ (.A1(_1493_),
    .A2(net793),
    .Y(_1689_),
    .B1(net784));
 sg13g2_o21ai_1 _2258_ (.B1(_1689_),
    .Y(_1690_),
    .A1(_0048_),
    .A2(net793));
 sg13g2_a21oi_1 _2259_ (.A1(net784),
    .A2(_1688_),
    .Y(_1691_),
    .B1(net765));
 sg13g2_a21oi_1 _2260_ (.A1(_1690_),
    .A2(_1691_),
    .Y(_1692_),
    .B1(net864));
 sg13g2_mux2_2 _2261_ (.A0(\GUScpu0.PC0[12] ),
    .A1(\GUScpu0.PC1[12] ),
    .S(net876),
    .X(_1693_));
 sg13g2_o21ai_1 _2262_ (.B1(_1596_),
    .Y(_1694_),
    .A1(net856),
    .A2(_1693_));
 sg13g2_a21oi_1 _2263_ (.A1(_1687_),
    .A2(_1692_),
    .Y(_1695_),
    .B1(_1694_));
 sg13g2_mux2_1 _2264_ (.A0(_0050_),
    .A1(_0049_),
    .S(net845),
    .X(_1696_));
 sg13g2_o21ai_1 _2265_ (.B1(net838),
    .Y(_1697_),
    .A1(_0052_),
    .A2(net846));
 sg13g2_inv_1 _2266_ (.Y(_1698_),
    .A(_1697_));
 sg13g2_o21ai_1 _2267_ (.B1(_1698_),
    .Y(_1699_),
    .A1(_0051_),
    .A2(net829));
 sg13g2_a21oi_1 _2268_ (.A1(net827),
    .A2(_1696_),
    .Y(_1700_),
    .B1(net824));
 sg13g2_mux4_1 _2269_ (.S0(net845),
    .A0(_0046_),
    .A1(_0045_),
    .A2(_0048_),
    .A3(_0047_),
    .S1(net838),
    .X(_1701_));
 sg13g2_inv_1 _2270_ (.Y(_1702_),
    .A(_1701_));
 sg13g2_a22oi_1 _2271_ (.Y(_1703_),
    .B1(_1702_),
    .B2(net824),
    .A2(_1700_),
    .A1(_1699_));
 sg13g2_a21oi_1 _2272_ (.A1(_1563_),
    .A2(_1703_),
    .Y(_1704_),
    .B1(_1605_));
 sg13g2_xnor2_1 _2273_ (.Y(_1705_),
    .A(net774),
    .B(_1704_));
 sg13g2_nor2b_1 _2274_ (.A(_1705_),
    .B_N(_1695_),
    .Y(_1706_));
 sg13g2_a21oi_1 _2275_ (.A1(_1486_),
    .A2(net799),
    .Y(_1707_),
    .B1(net780));
 sg13g2_o21ai_1 _2276_ (.B1(_1707_),
    .Y(_1708_),
    .A1(_0130_),
    .A2(net799));
 sg13g2_a21oi_1 _2277_ (.A1(_1487_),
    .A2(net791),
    .Y(_1709_),
    .B1(net783));
 sg13g2_o21ai_1 _2278_ (.B1(_1709_),
    .Y(_1710_),
    .A1(_0133_),
    .A2(net791));
 sg13g2_nand3_1 _2279_ (.B(_1708_),
    .C(_1710_),
    .A(net765),
    .Y(_1711_));
 sg13g2_mux2_1 _2280_ (.A0(_0127_),
    .A1(_0126_),
    .S(net788),
    .X(_0423_));
 sg13g2_a21oi_1 _2281_ (.A1(_1485_),
    .A2(net788),
    .Y(_0424_),
    .B1(net782));
 sg13g2_o21ai_1 _2282_ (.B1(_0424_),
    .Y(_0425_),
    .A1(_0129_),
    .A2(net788));
 sg13g2_a21oi_1 _2283_ (.A1(net782),
    .A2(_0423_),
    .Y(_0426_),
    .B1(net764));
 sg13g2_a21oi_1 _2284_ (.A1(_0425_),
    .A2(_0426_),
    .Y(_0427_),
    .B1(net862));
 sg13g2_mux2_2 _2285_ (.A0(\GUScpu0.PC0[1] ),
    .A1(\GUScpu0.PC1[1] ),
    .S(net872),
    .X(_0428_));
 sg13g2_inv_2 _2286_ (.Y(_0429_),
    .A(_0428_));
 sg13g2_a221oi_1 _2287_ (.B2(net862),
    .C1(_1595_),
    .B1(_0429_),
    .A1(_1711_),
    .Y(_0430_),
    .A2(_0427_));
 sg13g2_nor2_1 _2288_ (.A(_0130_),
    .B(net828),
    .Y(_0431_));
 sg13g2_o21ai_1 _2289_ (.B1(net826),
    .Y(_0432_),
    .A1(_0131_),
    .A2(net844));
 sg13g2_o21ai_1 _2290_ (.B1(net837),
    .Y(_0433_),
    .A1(_0133_),
    .A2(net844));
 sg13g2_a21oi_1 _2291_ (.A1(_1487_),
    .A2(net844),
    .Y(_0434_),
    .B1(_0433_));
 sg13g2_nor2_1 _2292_ (.A(net822),
    .B(_0434_),
    .Y(_0435_));
 sg13g2_o21ai_1 _2293_ (.B1(_0435_),
    .Y(_0436_),
    .A1(_0431_),
    .A2(_0432_));
 sg13g2_mux4_1 _2294_ (.S0(net841),
    .A0(_0127_),
    .A1(_0126_),
    .A2(_0129_),
    .A3(_0128_),
    .S1(net836),
    .X(_0437_));
 sg13g2_o21ai_1 _2295_ (.B1(_0436_),
    .Y(_0438_),
    .A1(_1619_),
    .A2(_0437_));
 sg13g2_inv_4 _2296_ (.A(_0438_),
    .Y(_0439_));
 sg13g2_nand2_1 _2297_ (.Y(_0440_),
    .A(_1477_),
    .B(net830));
 sg13g2_o21ai_1 _2298_ (.B1(_0440_),
    .Y(_0441_),
    .A1(net830),
    .A2(_0438_));
 sg13g2_xor2_1 _2299_ (.B(_0441_),
    .A(net773),
    .X(_0442_));
 sg13g2_nor2b_1 _2300_ (.A(_0442_),
    .B_N(_0430_),
    .Y(_0443_));
 sg13g2_xnor2_1 _2301_ (.Y(_0444_),
    .A(_0430_),
    .B(_0442_));
 sg13g2_mux2_1 _2302_ (.A0(_0140_),
    .A1(_0139_),
    .S(net789),
    .X(_0445_));
 sg13g2_nand2b_1 _2303_ (.Y(_0446_),
    .B(net798),
    .A_N(_0142_));
 sg13g2_a21oi_1 _2304_ (.A1(_1489_),
    .A2(net789),
    .Y(_0447_),
    .B1(net782));
 sg13g2_a221oi_1 _2305_ (.B2(_0447_),
    .C1(net775),
    .B1(_0446_),
    .A1(net782),
    .Y(_0448_),
    .A2(_0445_));
 sg13g2_mux2_1 _2306_ (.A0(_0136_),
    .A1(_0135_),
    .S(net789),
    .X(_0449_));
 sg13g2_nand2b_1 _2307_ (.Y(_0450_),
    .B(net798),
    .A_N(_0138_));
 sg13g2_a21oi_1 _2308_ (.A1(_1488_),
    .A2(net789),
    .Y(_0451_),
    .B1(net782));
 sg13g2_a221oi_1 _2309_ (.B2(_0451_),
    .C1(net764),
    .B1(_0450_),
    .A1(net782),
    .Y(_0452_),
    .A2(_0449_));
 sg13g2_nor3_2 _2310_ (.A(net862),
    .B(_0448_),
    .C(_0452_),
    .Y(_0453_));
 sg13g2_mux2_2 _2311_ (.A0(\GUScpu0.PC0[0] ),
    .A1(\GUScpu0.PC1[0] ),
    .S(net870),
    .X(_0454_));
 sg13g2_o21ai_1 _2312_ (.B1(net757),
    .Y(_0455_),
    .A1(net855),
    .A2(_0454_));
 sg13g2_nor2_1 _2313_ (.A(_0134_),
    .B(net832),
    .Y(_0456_));
 sg13g2_nor2_1 _2314_ (.A(_0139_),
    .B(net828),
    .Y(_0457_));
 sg13g2_o21ai_1 _2315_ (.B1(net826),
    .Y(_0458_),
    .A1(_0140_),
    .A2(net842));
 sg13g2_mux2_1 _2316_ (.A0(_0142_),
    .A1(_0141_),
    .S(net842),
    .X(_0459_));
 sg13g2_a21oi_1 _2317_ (.A1(net835),
    .A2(_0459_),
    .Y(_0460_),
    .B1(net822));
 sg13g2_o21ai_1 _2318_ (.B1(_0460_),
    .Y(_0461_),
    .A1(_0457_),
    .A2(_0458_));
 sg13g2_mux4_1 _2319_ (.S0(net842),
    .A0(_0136_),
    .A1(_0135_),
    .A2(_0138_),
    .A3(_0137_),
    .S1(net835),
    .X(_0462_));
 sg13g2_o21ai_1 _2320_ (.B1(_0461_),
    .Y(_0463_),
    .A1(_1619_),
    .A2(_0462_));
 sg13g2_a21oi_1 _2321_ (.A1(net832),
    .A2(_0463_),
    .Y(_0464_),
    .B1(_0456_));
 sg13g2_xor2_1 _2322_ (.B(_0464_),
    .A(net773),
    .X(_0465_));
 sg13g2_nor3_1 _2323_ (.A(_0453_),
    .B(_0455_),
    .C(_0465_),
    .Y(_0466_));
 sg13g2_o21ai_1 _2324_ (.B1(_0465_),
    .Y(_0467_),
    .A1(_0453_),
    .A2(_0455_));
 sg13g2_nor2b_1 _2325_ (.A(_0466_),
    .B_N(_0467_),
    .Y(_0468_));
 sg13g2_nand2_1 _2326_ (.Y(_0469_),
    .A(_1512_),
    .B(_1541_));
 sg13g2_o21ai_1 _2327_ (.B1(_1587_),
    .Y(_0470_),
    .A1(net880),
    .A2(_1542_));
 sg13g2_a21oi_1 _2328_ (.A1(_1477_),
    .A2(_1526_),
    .Y(_0471_),
    .B1(_0470_));
 sg13g2_mux2_1 _2329_ (.A0(\GUScpu0.cv[0][1] ),
    .A1(\GUScpu0.cv[1][1] ),
    .S(net870),
    .X(_0472_));
 sg13g2_mux2_1 _2330_ (.A0(_0472_),
    .A1(net773),
    .S(_0471_),
    .X(_0473_));
 sg13g2_a21o_1 _2331_ (.A2(_0473_),
    .A1(_0467_),
    .B1(_0466_),
    .X(_0474_));
 sg13g2_a21oi_1 _2332_ (.A1(_0444_),
    .A2(_0474_),
    .Y(_0475_),
    .B1(_0443_));
 sg13g2_a21o_1 _2333_ (.A2(_0474_),
    .A1(_0444_),
    .B1(_0443_),
    .X(_0476_));
 sg13g2_mux2_1 _2334_ (.A0(_0123_),
    .A1(_0122_),
    .S(net788),
    .X(_0477_));
 sg13g2_nand2b_1 _2335_ (.Y(_0478_),
    .B(net798),
    .A_N(_0125_));
 sg13g2_a21oi_1 _2336_ (.A1(_1484_),
    .A2(net787),
    .Y(_0479_),
    .B1(net781));
 sg13g2_a221oi_1 _2337_ (.B2(_0479_),
    .C1(net775),
    .B1(_0478_),
    .A1(net781),
    .Y(_0480_),
    .A2(_0477_));
 sg13g2_nor2_1 _2338_ (.A(_0118_),
    .B(net798),
    .Y(_0481_));
 sg13g2_o21ai_1 _2339_ (.B1(net781),
    .Y(_0482_),
    .A1(_0119_),
    .A2(net787));
 sg13g2_mux2_1 _2340_ (.A0(_0121_),
    .A1(_0120_),
    .S(net787),
    .X(_0483_));
 sg13g2_a21oi_1 _2341_ (.A1(net777),
    .A2(_0483_),
    .Y(_0484_),
    .B1(net764));
 sg13g2_o21ai_1 _2342_ (.B1(_0484_),
    .Y(_0485_),
    .A1(_0481_),
    .A2(_0482_));
 sg13g2_nor2_1 _2343_ (.A(net862),
    .B(_0480_),
    .Y(_0486_));
 sg13g2_and2_1 _2344_ (.A(net872),
    .B(\GUScpu0.PC1[2] ),
    .X(_0487_));
 sg13g2_a21oi_2 _2345_ (.B1(_0487_),
    .Y(_0488_),
    .A2(\GUScpu0.PC0[2] ),
    .A1(_1472_));
 sg13g2_a21o_2 _2346_ (.A2(\GUScpu0.PC0[2] ),
    .A1(_1472_),
    .B1(_0487_),
    .X(_0489_));
 sg13g2_a221oi_1 _2347_ (.B2(net862),
    .C1(_1595_),
    .B1(_0488_),
    .A1(_0485_),
    .Y(_0490_),
    .A2(_0486_));
 sg13g2_mux2_1 _2348_ (.A0(_0123_),
    .A1(_0122_),
    .S(net840),
    .X(_0491_));
 sg13g2_o21ai_1 _2349_ (.B1(net836),
    .Y(_0492_),
    .A1(_0125_),
    .A2(net840));
 sg13g2_a21o_1 _2350_ (.A2(net840),
    .A1(_1484_),
    .B1(_0492_),
    .X(_0493_));
 sg13g2_a21oi_1 _2351_ (.A1(net826),
    .A2(_0491_),
    .Y(_0494_),
    .B1(net823));
 sg13g2_mux4_1 _2352_ (.S0(net841),
    .A0(_0119_),
    .A1(_0118_),
    .A2(_0121_),
    .A3(_0120_),
    .S1(net836),
    .X(_0495_));
 sg13g2_inv_1 _2353_ (.Y(_0496_),
    .A(_0495_));
 sg13g2_a22oi_1 _2354_ (.Y(_0497_),
    .B1(_0496_),
    .B2(net822),
    .A2(_0494_),
    .A1(_0493_));
 sg13g2_mux2_1 _2355_ (.A0(_0088_),
    .A1(_0497_),
    .S(net832),
    .X(_0498_));
 sg13g2_xnor2_1 _2356_ (.Y(_0499_),
    .A(net773),
    .B(_0498_));
 sg13g2_and2_1 _2357_ (.A(_0490_),
    .B(_0499_),
    .X(_0500_));
 sg13g2_xor2_1 _2358_ (.B(_0499_),
    .A(_0490_),
    .X(_0501_));
 sg13g2_a21oi_1 _2359_ (.A1(_1483_),
    .A2(net798),
    .Y(_0502_),
    .B1(net777));
 sg13g2_o21ai_1 _2360_ (.B1(_0502_),
    .Y(_0503_),
    .A1(_0114_),
    .A2(net798));
 sg13g2_mux2_1 _2361_ (.A0(_0117_),
    .A1(_0116_),
    .S(net788),
    .X(_0504_));
 sg13g2_a21oi_1 _2362_ (.A1(net777),
    .A2(_0504_),
    .Y(_0505_),
    .B1(net775));
 sg13g2_mux2_1 _2363_ (.A0(_0111_),
    .A1(_0110_),
    .S(net787),
    .X(_0506_));
 sg13g2_a21oi_1 _2364_ (.A1(_1482_),
    .A2(net788),
    .Y(_0507_),
    .B1(net781));
 sg13g2_o21ai_1 _2365_ (.B1(_0507_),
    .Y(_0508_),
    .A1(_0113_),
    .A2(net788));
 sg13g2_a21oi_1 _2366_ (.A1(net781),
    .A2(_0506_),
    .Y(_0509_),
    .B1(net764));
 sg13g2_a221oi_1 _2367_ (.B2(_0509_),
    .C1(net863),
    .B1(_0508_),
    .A1(_0503_),
    .Y(_0510_),
    .A2(_0505_));
 sg13g2_mux2_2 _2368_ (.A0(\GUScpu0.PC0[3] ),
    .A1(\GUScpu0.PC1[3] ),
    .S(net873),
    .X(_0511_));
 sg13g2_o21ai_1 _2369_ (.B1(net757),
    .Y(_0512_),
    .A1(net855),
    .A2(_0511_));
 sg13g2_mux2_1 _2370_ (.A0(_0115_),
    .A1(_0114_),
    .S(net840),
    .X(_0513_));
 sg13g2_o21ai_1 _2371_ (.B1(net836),
    .Y(_0514_),
    .A1(_0117_),
    .A2(net841));
 sg13g2_inv_1 _2372_ (.Y(_0515_),
    .A(_0514_));
 sg13g2_o21ai_1 _2373_ (.B1(_0515_),
    .Y(_0516_),
    .A1(_0116_),
    .A2(net828));
 sg13g2_a21oi_1 _2374_ (.A1(net826),
    .A2(_0513_),
    .Y(_0517_),
    .B1(net822));
 sg13g2_mux4_1 _2375_ (.S0(net841),
    .A0(_0111_),
    .A1(_0110_),
    .A2(_0113_),
    .A3(_0112_),
    .S1(net835),
    .X(_0518_));
 sg13g2_nor2_1 _2376_ (.A(_1619_),
    .B(_0518_),
    .Y(_0519_));
 sg13g2_a21oi_2 _2377_ (.B1(_0519_),
    .Y(_0520_),
    .A2(_0517_),
    .A1(_0516_));
 sg13g2_a21o_2 _2378_ (.A2(_0517_),
    .A1(_0516_),
    .B1(_0519_),
    .X(_0521_));
 sg13g2_nand2_1 _2379_ (.Y(_0522_),
    .A(_1474_),
    .B(net830));
 sg13g2_o21ai_1 _2380_ (.B1(_0522_),
    .Y(_0523_),
    .A1(net830),
    .A2(_0520_));
 sg13g2_xnor2_1 _2381_ (.Y(_0524_),
    .A(net773),
    .B(_0523_));
 sg13g2_nor3_2 _2382_ (.A(_0510_),
    .B(_0512_),
    .C(_0524_),
    .Y(_0525_));
 sg13g2_o21ai_1 _2383_ (.B1(_0524_),
    .Y(_0526_),
    .A1(_0510_),
    .A2(_0512_));
 sg13g2_nor2b_1 _2384_ (.A(_0525_),
    .B_N(_0526_),
    .Y(_0527_));
 sg13g2_nand2b_1 _2385_ (.Y(_0528_),
    .B(_0526_),
    .A_N(_0525_));
 sg13g2_nand2_1 _2386_ (.Y(_0529_),
    .A(_0501_),
    .B(_0527_));
 sg13g2_o21ai_1 _2387_ (.B1(_0526_),
    .Y(_0530_),
    .A1(_0500_),
    .A2(_0525_));
 sg13g2_o21ai_1 _2388_ (.B1(_0530_),
    .Y(_0531_),
    .A1(_0475_),
    .A2(_0529_));
 sg13g2_nor2_1 _2389_ (.A(_0147_),
    .B(net801),
    .Y(_0532_));
 sg13g2_o21ai_1 _2390_ (.B1(net786),
    .Y(_0533_),
    .A1(_0148_),
    .A2(net792));
 sg13g2_mux2_1 _2391_ (.A0(_0150_),
    .A1(_0149_),
    .S(net791),
    .X(_0534_));
 sg13g2_a21oi_1 _2392_ (.A1(net778),
    .A2(_0534_),
    .Y(_0535_),
    .B1(net775));
 sg13g2_o21ai_1 _2393_ (.B1(_0535_),
    .Y(_0536_),
    .A1(_0532_),
    .A2(_0533_));
 sg13g2_mux2_1 _2394_ (.A0(_0144_),
    .A1(_0143_),
    .S(net790),
    .X(_0537_));
 sg13g2_a21oi_1 _2395_ (.A1(_1490_),
    .A2(net791),
    .Y(_0538_),
    .B1(net783));
 sg13g2_o21ai_1 _2396_ (.B1(_0538_),
    .Y(_0539_),
    .A1(_0146_),
    .A2(net791));
 sg13g2_a21oi_1 _2397_ (.A1(net783),
    .A2(_0537_),
    .Y(_0540_),
    .B1(net764));
 sg13g2_a21oi_2 _2398_ (.B1(net863),
    .Y(_0541_),
    .A2(_0540_),
    .A1(_0539_));
 sg13g2_mux2_2 _2399_ (.A0(\GUScpu0.PC0[6] ),
    .A1(\GUScpu0.PC1[6] ),
    .S(net874),
    .X(_0542_));
 sg13g2_inv_1 _2400_ (.Y(_0543_),
    .A(_0542_));
 sg13g2_a221oi_1 _2401_ (.B2(net864),
    .C1(_1595_),
    .B1(_0543_),
    .A1(_0536_),
    .Y(_0544_),
    .A2(_0541_));
 sg13g2_mux2_1 _2402_ (.A0(_0148_),
    .A1(_0147_),
    .S(net847),
    .X(_0545_));
 sg13g2_nor2_1 _2403_ (.A(_0149_),
    .B(net828),
    .Y(_0546_));
 sg13g2_o21ai_1 _2404_ (.B1(net837),
    .Y(_0547_),
    .A1(_0150_),
    .A2(net843));
 sg13g2_a21oi_1 _2405_ (.A1(net826),
    .A2(_0545_),
    .Y(_0548_),
    .B1(net823));
 sg13g2_o21ai_1 _2406_ (.B1(_0548_),
    .Y(_0549_),
    .A1(_0546_),
    .A2(_0547_));
 sg13g2_mux4_1 _2407_ (.S0(net843),
    .A0(_0144_),
    .A1(_0143_),
    .A2(_0146_),
    .A3(_0145_),
    .S1(net837),
    .X(_0550_));
 sg13g2_o21ai_1 _2408_ (.B1(_0549_),
    .Y(_0551_),
    .A1(_1619_),
    .A2(_0550_));
 sg13g2_and2_1 _2409_ (.A(net831),
    .B(_1604_),
    .X(_0552_));
 sg13g2_o21ai_1 _2410_ (.B1(net830),
    .Y(_0553_),
    .A1(_1565_),
    .A2(_1604_));
 sg13g2_nor2_1 _2411_ (.A(_0100_),
    .B(_0553_),
    .Y(_0554_));
 sg13g2_a21oi_1 _2412_ (.A1(net832),
    .A2(_0551_),
    .Y(_0555_),
    .B1(_0554_));
 sg13g2_xnor2_1 _2413_ (.Y(_0556_),
    .A(net774),
    .B(_0555_));
 sg13g2_and2_1 _2414_ (.A(_0544_),
    .B(_0556_),
    .X(_0557_));
 sg13g2_xor2_1 _2415_ (.B(_0556_),
    .A(_0544_),
    .X(_0558_));
 sg13g2_inv_1 _2416_ (.Y(_0559_),
    .A(_0558_));
 sg13g2_a21oi_1 _2417_ (.A1(_1492_),
    .A2(net799),
    .Y(_0560_),
    .B1(net777));
 sg13g2_o21ai_1 _2418_ (.B1(_0560_),
    .Y(_0561_),
    .A1(_0155_),
    .A2(net799));
 sg13g2_mux2_1 _2419_ (.A0(_0158_),
    .A1(_0157_),
    .S(net790),
    .X(_0562_));
 sg13g2_a21oi_1 _2420_ (.A1(net777),
    .A2(_0562_),
    .Y(_0563_),
    .B1(net775));
 sg13g2_mux2_1 _2421_ (.A0(_0152_),
    .A1(_0151_),
    .S(net790),
    .X(_0564_));
 sg13g2_a21oi_1 _2422_ (.A1(_1491_),
    .A2(net790),
    .Y(_0565_),
    .B1(net783));
 sg13g2_o21ai_1 _2423_ (.B1(_0565_),
    .Y(_0566_),
    .A1(_0154_),
    .A2(net790));
 sg13g2_a21oi_1 _2424_ (.A1(net783),
    .A2(_0564_),
    .Y(_0567_),
    .B1(net765));
 sg13g2_a221oi_1 _2425_ (.B2(_0567_),
    .C1(net862),
    .B1(_0566_),
    .A1(_0561_),
    .Y(_0568_),
    .A2(_0563_));
 sg13g2_mux2_2 _2426_ (.A0(\GUScpu0.PC0[7] ),
    .A1(\GUScpu0.PC1[7] ),
    .S(net874),
    .X(_0569_));
 sg13g2_o21ai_1 _2427_ (.B1(net757),
    .Y(_0570_),
    .A1(net856),
    .A2(_0569_));
 sg13g2_or2_1 _2428_ (.X(_0571_),
    .B(_0553_),
    .A(_0101_));
 sg13g2_mux2_1 _2429_ (.A0(_0156_),
    .A1(_0155_),
    .S(net843),
    .X(_0572_));
 sg13g2_o21ai_1 _2430_ (.B1(net837),
    .Y(_0573_),
    .A1(_0158_),
    .A2(net843));
 sg13g2_inv_1 _2431_ (.Y(_0574_),
    .A(_0573_));
 sg13g2_o21ai_1 _2432_ (.B1(_0574_),
    .Y(_0575_),
    .A1(_0157_),
    .A2(net828));
 sg13g2_a21oi_1 _2433_ (.A1(net826),
    .A2(_0572_),
    .Y(_0576_),
    .B1(net822));
 sg13g2_mux4_1 _2434_ (.S0(net843),
    .A0(_0152_),
    .A1(_0151_),
    .A2(_0154_),
    .A3(_0153_),
    .S1(_1611_),
    .X(_0577_));
 sg13g2_nor2_1 _2435_ (.A(_1619_),
    .B(_0577_),
    .Y(_0578_));
 sg13g2_a21oi_2 _2436_ (.B1(_0578_),
    .Y(_0579_),
    .A2(_0576_),
    .A1(_0575_));
 sg13g2_o21ai_1 _2437_ (.B1(_0571_),
    .Y(_0580_),
    .A1(net831),
    .A2(_0579_));
 sg13g2_xnor2_1 _2438_ (.Y(_0581_),
    .A(net773),
    .B(_0580_));
 sg13g2_nor3_2 _2439_ (.A(_0568_),
    .B(_0570_),
    .C(_0581_),
    .Y(_0582_));
 sg13g2_o21ai_1 _2440_ (.B1(_0581_),
    .Y(_0583_),
    .A1(_0568_),
    .A2(_0570_));
 sg13g2_nor2b_2 _2441_ (.A(_0582_),
    .B_N(_0583_),
    .Y(_0584_));
 sg13g2_nand2_1 _2442_ (.Y(_0585_),
    .A(_0558_),
    .B(_0584_));
 sg13g2_mux2_1 _2443_ (.A0(_0107_),
    .A1(_0106_),
    .S(net787),
    .X(_0586_));
 sg13g2_nand2b_1 _2444_ (.Y(_0587_),
    .B(net798),
    .A_N(_0109_));
 sg13g2_a21oi_1 _2445_ (.A1(_1481_),
    .A2(net787),
    .Y(_0588_),
    .B1(net781));
 sg13g2_a221oi_1 _2446_ (.B2(_0588_),
    .C1(net775),
    .B1(_0587_),
    .A1(net781),
    .Y(_0589_),
    .A2(_0586_));
 sg13g2_nor2_1 _2447_ (.A(_0102_),
    .B(net798),
    .Y(_0590_));
 sg13g2_o21ai_1 _2448_ (.B1(net781),
    .Y(_0591_),
    .A1(_0103_),
    .A2(net787));
 sg13g2_mux2_1 _2449_ (.A0(_0105_),
    .A1(_0104_),
    .S(net787),
    .X(_0592_));
 sg13g2_a21oi_1 _2450_ (.A1(net777),
    .A2(_0592_),
    .Y(_0593_),
    .B1(net764));
 sg13g2_o21ai_1 _2451_ (.B1(_0593_),
    .Y(_0594_),
    .A1(_0590_),
    .A2(_0591_));
 sg13g2_nor2_1 _2452_ (.A(net862),
    .B(_0589_),
    .Y(_0595_));
 sg13g2_mux2_2 _2453_ (.A0(\GUScpu0.PC0[4] ),
    .A1(\GUScpu0.PC1[4] ),
    .S(net872),
    .X(_0596_));
 sg13g2_o21ai_1 _2454_ (.B1(net757),
    .Y(_0597_),
    .A1(net855),
    .A2(_0596_));
 sg13g2_a21oi_2 _2455_ (.B1(_0597_),
    .Y(_0598_),
    .A2(_0595_),
    .A1(_0594_));
 sg13g2_mux2_1 _2456_ (.A0(_0107_),
    .A1(_0106_),
    .S(net840),
    .X(_0599_));
 sg13g2_o21ai_1 _2457_ (.B1(net835),
    .Y(_0600_),
    .A1(_0109_),
    .A2(net840));
 sg13g2_a21o_1 _2458_ (.A2(net840),
    .A1(_1481_),
    .B1(_0600_),
    .X(_0601_));
 sg13g2_a21oi_1 _2459_ (.A1(net826),
    .A2(_0599_),
    .Y(_0602_),
    .B1(net822));
 sg13g2_mux4_1 _2460_ (.S0(net840),
    .A0(_0103_),
    .A1(_0102_),
    .A2(_0105_),
    .A3(_0104_),
    .S1(net835),
    .X(_0603_));
 sg13g2_inv_1 _2461_ (.Y(_0604_),
    .A(_0603_));
 sg13g2_a22oi_1 _2462_ (.Y(_0605_),
    .B1(_0604_),
    .B2(net822),
    .A2(_0602_),
    .A1(_0601_));
 sg13g2_mux2_1 _2463_ (.A0(_0094_),
    .A1(_0605_),
    .S(net832),
    .X(_0606_));
 sg13g2_xnor2_1 _2464_ (.Y(_0607_),
    .A(net773),
    .B(_0606_));
 sg13g2_and2_1 _2465_ (.A(_0598_),
    .B(_0607_),
    .X(_0608_));
 sg13g2_xor2_1 _2466_ (.B(_0607_),
    .A(_0598_),
    .X(_0609_));
 sg13g2_mux4_1 _2467_ (.S0(net789),
    .A0(_0096_),
    .A1(_0095_),
    .A2(_0098_),
    .A3(_0097_),
    .S1(net777),
    .X(_0610_));
 sg13g2_nor2_2 _2468_ (.A(net775),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_mux4_1 _2469_ (.S0(net789),
    .A0(_0086_),
    .A1(_0085_),
    .A2(_0092_),
    .A3(_0091_),
    .S1(net777),
    .X(_0612_));
 sg13g2_o21ai_1 _2470_ (.B1(net855),
    .Y(_0613_),
    .A1(net764),
    .A2(_0612_));
 sg13g2_nor2_1 _2471_ (.A(_0611_),
    .B(_0613_),
    .Y(_0614_));
 sg13g2_mux2_2 _2472_ (.A0(\GUScpu0.PC0[5] ),
    .A1(\GUScpu0.PC1[5] ),
    .S(net872),
    .X(_0615_));
 sg13g2_nor2_1 _2473_ (.A(net855),
    .B(_0615_),
    .Y(_0616_));
 sg13g2_or2_1 _2474_ (.X(_0617_),
    .B(_0616_),
    .A(_1595_));
 sg13g2_a21oi_1 _2475_ (.A1(_1476_),
    .A2(net842),
    .Y(_0618_),
    .B1(net835));
 sg13g2_o21ai_1 _2476_ (.B1(_0618_),
    .Y(_0619_),
    .A1(_0096_),
    .A2(net842));
 sg13g2_mux2_1 _2477_ (.A0(_0098_),
    .A1(_0097_),
    .S(net842),
    .X(_0620_));
 sg13g2_a21oi_1 _2478_ (.A1(net835),
    .A2(_0620_),
    .Y(_0621_),
    .B1(net822));
 sg13g2_mux4_1 _2479_ (.S0(net842),
    .A0(_0086_),
    .A1(_0085_),
    .A2(_0092_),
    .A3(_0091_),
    .S1(net835),
    .X(_0622_));
 sg13g2_nor2_1 _2480_ (.A(_1619_),
    .B(_0622_),
    .Y(_0623_));
 sg13g2_a21oi_2 _2481_ (.B1(_0623_),
    .Y(_0624_),
    .A2(_0621_),
    .A1(_0619_));
 sg13g2_nand2b_1 _2482_ (.Y(_0625_),
    .B(\GUScpu0.IR[5] ),
    .A_N(_0553_));
 sg13g2_o21ai_1 _2483_ (.B1(_0625_),
    .Y(_0626_),
    .A1(net830),
    .A2(_0624_));
 sg13g2_xnor2_1 _2484_ (.Y(_0627_),
    .A(net773),
    .B(_0626_));
 sg13g2_o21ai_1 _2485_ (.B1(_0627_),
    .Y(_0628_),
    .A1(_0614_),
    .A2(_0617_));
 sg13g2_or4_1 _2486_ (.A(_1595_),
    .B(_0614_),
    .C(_0616_),
    .D(_0627_),
    .X(_0629_));
 sg13g2_inv_1 _2487_ (.Y(_0630_),
    .A(_0629_));
 sg13g2_and2_1 _2488_ (.A(_0628_),
    .B(_0629_),
    .X(_0631_));
 sg13g2_and4_1 _2489_ (.A(_0558_),
    .B(_0584_),
    .C(_0609_),
    .D(_0631_),
    .X(_0632_));
 sg13g2_o21ai_1 _2490_ (.B1(_0628_),
    .Y(_0633_),
    .A1(_0608_),
    .A2(_0630_));
 sg13g2_a21oi_1 _2491_ (.A1(_0557_),
    .A2(_0583_),
    .Y(_0634_),
    .B1(_0582_));
 sg13g2_o21ai_1 _2492_ (.B1(_0634_),
    .Y(_0635_),
    .A1(_0585_),
    .A2(_0633_));
 sg13g2_a21oi_2 _2493_ (.B1(_0635_),
    .Y(_0636_),
    .A2(_0632_),
    .A1(_0531_));
 sg13g2_mux2_1 _2494_ (.A0(_0164_),
    .A1(_0163_),
    .S(net792),
    .X(_0637_));
 sg13g2_nor2_1 _2495_ (.A(_0166_),
    .B(net792),
    .Y(_0638_));
 sg13g2_o21ai_1 _2496_ (.B1(net778),
    .Y(_0639_),
    .A1(_0165_),
    .A2(net801));
 sg13g2_o21ai_1 _2497_ (.B1(_1574_),
    .Y(_0640_),
    .A1(_0638_),
    .A2(_0639_));
 sg13g2_a21oi_1 _2498_ (.A1(net786),
    .A2(_0637_),
    .Y(_0641_),
    .B1(_0640_));
 sg13g2_mux2_1 _2499_ (.A0(_0160_),
    .A1(_0159_),
    .S(net792),
    .X(_0642_));
 sg13g2_nor2_1 _2500_ (.A(_0162_),
    .B(net792),
    .Y(_0643_));
 sg13g2_o21ai_1 _2501_ (.B1(net778),
    .Y(_0644_),
    .A1(_0161_),
    .A2(net801));
 sg13g2_o21ai_1 _2502_ (.B1(net776),
    .Y(_0645_),
    .A1(_0643_),
    .A2(_0644_));
 sg13g2_a21oi_1 _2503_ (.A1(net786),
    .A2(_0642_),
    .Y(_0646_),
    .B1(_0645_));
 sg13g2_nor3_2 _2504_ (.A(_1560_),
    .B(_0641_),
    .C(_0646_),
    .Y(_0647_));
 sg13g2_mux2_2 _2505_ (.A0(\GUScpu0.PC0[8] ),
    .A1(\GUScpu0.PC1[8] ),
    .S(net875),
    .X(_0648_));
 sg13g2_nor2_1 _2506_ (.A(net856),
    .B(_0648_),
    .Y(_0649_));
 sg13g2_nor3_1 _2507_ (.A(_1595_),
    .B(_0647_),
    .C(_0649_),
    .Y(_0650_));
 sg13g2_nand2_1 _2508_ (.Y(_0651_),
    .A(_1473_),
    .B(_0552_));
 sg13g2_mux2_1 _2509_ (.A0(_0164_),
    .A1(_0163_),
    .S(net847),
    .X(_0652_));
 sg13g2_o21ai_1 _2510_ (.B1(net839),
    .Y(_0653_),
    .A1(_0166_),
    .A2(net847));
 sg13g2_inv_1 _2511_ (.Y(_0654_),
    .A(_0653_));
 sg13g2_o21ai_1 _2512_ (.B1(_0654_),
    .Y(_0655_),
    .A1(_0165_),
    .A2(net829));
 sg13g2_a21oi_1 _2513_ (.A1(net827),
    .A2(_0652_),
    .Y(_0656_),
    .B1(net825));
 sg13g2_mux4_1 _2514_ (.S0(net847),
    .A0(_0160_),
    .A1(_0159_),
    .A2(_0162_),
    .A3(_0161_),
    .S1(net839),
    .X(_0657_));
 sg13g2_inv_1 _2515_ (.Y(_0658_),
    .A(_0657_));
 sg13g2_a22oi_1 _2516_ (.Y(_0659_),
    .B1(_0658_),
    .B2(net825),
    .A2(_0656_),
    .A1(_0655_));
 sg13g2_o21ai_1 _2517_ (.B1(_0651_),
    .Y(_0660_),
    .A1(net831),
    .A2(_0659_));
 sg13g2_xnor2_1 _2518_ (.Y(_0661_),
    .A(_1602_),
    .B(_0660_));
 sg13g2_nor4_2 _2519_ (.A(_1595_),
    .B(_0647_),
    .C(_0649_),
    .Y(_0662_),
    .D(_0661_));
 sg13g2_inv_1 _2520_ (.Y(_0663_),
    .A(_0662_));
 sg13g2_xor2_1 _2521_ (.B(_0661_),
    .A(_0650_),
    .X(_0664_));
 sg13g2_inv_1 _2522_ (.Y(_0665_),
    .A(_0664_));
 sg13g2_mux2_1 _2523_ (.A0(_0026_),
    .A1(_0025_),
    .S(net795),
    .X(_0666_));
 sg13g2_nor2_1 _2524_ (.A(_0028_),
    .B(net795),
    .Y(_0667_));
 sg13g2_o21ai_1 _2525_ (.B1(net778),
    .Y(_0668_),
    .A1(_0027_),
    .A2(net800));
 sg13g2_o21ai_1 _2526_ (.B1(net765),
    .Y(_0669_),
    .A1(_0667_),
    .A2(_0668_));
 sg13g2_a21oi_1 _2527_ (.A1(net784),
    .A2(_0666_),
    .Y(_0670_),
    .B1(_0669_));
 sg13g2_mux2_1 _2528_ (.A0(_0168_),
    .A1(_0167_),
    .S(net795),
    .X(_0671_));
 sg13g2_nor2_1 _2529_ (.A(_0170_),
    .B(net795),
    .Y(_0672_));
 sg13g2_o21ai_1 _2530_ (.B1(net778),
    .Y(_0673_),
    .A1(_0169_),
    .A2(net800));
 sg13g2_o21ai_1 _2531_ (.B1(net776),
    .Y(_0674_),
    .A1(_0672_),
    .A2(_0673_));
 sg13g2_a21oi_1 _2532_ (.A1(net784),
    .A2(_0671_),
    .Y(_0675_),
    .B1(_0674_));
 sg13g2_nor3_2 _2533_ (.A(net864),
    .B(_0670_),
    .C(_0675_),
    .Y(_0676_));
 sg13g2_mux2_2 _2534_ (.A0(\GUScpu0.PC0[9] ),
    .A1(\GUScpu0.PC1[9] ),
    .S(net878),
    .X(_0677_));
 sg13g2_o21ai_1 _2535_ (.B1(net757),
    .Y(_0678_),
    .A1(net856),
    .A2(_0677_));
 sg13g2_mux2_1 _2536_ (.A0(_0026_),
    .A1(_0025_),
    .S(net845),
    .X(_0679_));
 sg13g2_o21ai_1 _2537_ (.B1(net838),
    .Y(_0680_),
    .A1(_0028_),
    .A2(net845));
 sg13g2_inv_1 _2538_ (.Y(_0681_),
    .A(_0680_));
 sg13g2_o21ai_1 _2539_ (.B1(_0681_),
    .Y(_0682_),
    .A1(_0027_),
    .A2(net828));
 sg13g2_a21oi_1 _2540_ (.A1(net827),
    .A2(_0679_),
    .Y(_0683_),
    .B1(net824));
 sg13g2_mux4_1 _2541_ (.S0(net845),
    .A0(_0168_),
    .A1(_0167_),
    .A2(_0170_),
    .A3(_0169_),
    .S1(net838),
    .X(_0684_));
 sg13g2_inv_1 _2542_ (.Y(_0685_),
    .A(_0684_));
 sg13g2_a22oi_1 _2543_ (.Y(_0686_),
    .B1(_0685_),
    .B2(net824),
    .A2(_0683_),
    .A1(_0682_));
 sg13g2_nand2_1 _2544_ (.Y(_0687_),
    .A(_1475_),
    .B(_0552_));
 sg13g2_o21ai_1 _2545_ (.B1(_0687_),
    .Y(_0688_),
    .A1(net831),
    .A2(_0686_));
 sg13g2_xnor2_1 _2546_ (.Y(_0689_),
    .A(net774),
    .B(_0688_));
 sg13g2_nor3_1 _2547_ (.A(_0676_),
    .B(_0678_),
    .C(_0689_),
    .Y(_0690_));
 sg13g2_o21ai_1 _2548_ (.B1(_0689_),
    .Y(_0691_),
    .A1(_0676_),
    .A2(_0678_));
 sg13g2_nand2b_1 _2549_ (.Y(_0692_),
    .B(_0691_),
    .A_N(_0690_));
 sg13g2_or2_1 _2550_ (.X(_0693_),
    .B(_0692_),
    .A(_0664_));
 sg13g2_mux2_1 _2551_ (.A0(_0042_),
    .A1(_0041_),
    .S(net792),
    .X(_0694_));
 sg13g2_nor2_1 _2552_ (.A(_0044_),
    .B(net797),
    .Y(_0695_));
 sg13g2_o21ai_1 _2553_ (.B1(net779),
    .Y(_0696_),
    .A1(_0043_),
    .A2(net800));
 sg13g2_o21ai_1 _2554_ (.B1(net765),
    .Y(_0697_),
    .A1(_0695_),
    .A2(_0696_));
 sg13g2_a21oi_1 _2555_ (.A1(net786),
    .A2(_0694_),
    .Y(_0698_),
    .B1(_0697_));
 sg13g2_mux2_1 _2556_ (.A0(_0038_),
    .A1(_0037_),
    .S(net792),
    .X(_0699_));
 sg13g2_nor2_1 _2557_ (.A(_0040_),
    .B(net792),
    .Y(_0700_));
 sg13g2_o21ai_1 _2558_ (.B1(net778),
    .Y(_0701_),
    .A1(_0039_),
    .A2(net800));
 sg13g2_o21ai_1 _2559_ (.B1(net776),
    .Y(_0702_),
    .A1(_0700_),
    .A2(_0701_));
 sg13g2_a21oi_1 _2560_ (.A1(net786),
    .A2(_0699_),
    .Y(_0703_),
    .B1(_0702_));
 sg13g2_nor3_1 _2561_ (.A(net864),
    .B(_0698_),
    .C(_0703_),
    .Y(_0704_));
 sg13g2_mux2_2 _2562_ (.A0(\GUScpu0.PC0[11] ),
    .A1(\GUScpu0.PC1[11] ),
    .S(net877),
    .X(_0705_));
 sg13g2_o21ai_1 _2563_ (.B1(net757),
    .Y(_0706_),
    .A1(net855),
    .A2(_0705_));
 sg13g2_mux2_1 _2564_ (.A0(_0042_),
    .A1(_0041_),
    .S(net847),
    .X(_0707_));
 sg13g2_o21ai_1 _2565_ (.B1(net839),
    .Y(_0708_),
    .A1(_0044_),
    .A2(net847));
 sg13g2_inv_1 _2566_ (.Y(_0709_),
    .A(_0708_));
 sg13g2_o21ai_1 _2567_ (.B1(_0709_),
    .Y(_0710_),
    .A1(_0043_),
    .A2(net829));
 sg13g2_a21oi_1 _2568_ (.A1(net827),
    .A2(_0707_),
    .Y(_0711_),
    .B1(net825));
 sg13g2_mux4_1 _2569_ (.S0(net847),
    .A0(_0038_),
    .A1(_0037_),
    .A2(_0040_),
    .A3(_0039_),
    .S1(net839),
    .X(_0712_));
 sg13g2_inv_1 _2570_ (.Y(_0713_),
    .A(_0712_));
 sg13g2_a22oi_1 _2571_ (.Y(_0714_),
    .B1(_0713_),
    .B2(net825),
    .A2(_0711_),
    .A1(_0710_));
 sg13g2_a21oi_1 _2572_ (.A1(_1563_),
    .A2(_0714_),
    .Y(_0715_),
    .B1(_1605_));
 sg13g2_xnor2_1 _2573_ (.Y(_0716_),
    .A(net774),
    .B(_0715_));
 sg13g2_nor3_1 _2574_ (.A(_0704_),
    .B(_0706_),
    .C(_0716_),
    .Y(_0717_));
 sg13g2_o21ai_1 _2575_ (.B1(_0716_),
    .Y(_0718_),
    .A1(_0704_),
    .A2(_0706_));
 sg13g2_nor2b_1 _2576_ (.A(_0717_),
    .B_N(_0718_),
    .Y(_0719_));
 sg13g2_mux2_1 _2577_ (.A0(_0034_),
    .A1(_0033_),
    .S(net795),
    .X(_0720_));
 sg13g2_nor2_1 _2578_ (.A(_0036_),
    .B(net793),
    .Y(_0721_));
 sg13g2_o21ai_1 _2579_ (.B1(net778),
    .Y(_0722_),
    .A1(_0035_),
    .A2(net800));
 sg13g2_o21ai_1 _2580_ (.B1(net765),
    .Y(_0723_),
    .A1(_0721_),
    .A2(_0722_));
 sg13g2_a21oi_1 _2581_ (.A1(net785),
    .A2(_0720_),
    .Y(_0724_),
    .B1(_0723_));
 sg13g2_mux2_1 _2582_ (.A0(_0030_),
    .A1(_0029_),
    .S(net793),
    .X(_0725_));
 sg13g2_nor2_1 _2583_ (.A(_0032_),
    .B(net793),
    .Y(_0726_));
 sg13g2_o21ai_1 _2584_ (.B1(net778),
    .Y(_0727_),
    .A1(_0031_),
    .A2(net800));
 sg13g2_o21ai_1 _2585_ (.B1(net776),
    .Y(_0728_),
    .A1(_0726_),
    .A2(_0727_));
 sg13g2_a21oi_1 _2586_ (.A1(net784),
    .A2(_0725_),
    .Y(_0729_),
    .B1(_0728_));
 sg13g2_nor3_2 _2587_ (.A(net864),
    .B(_0724_),
    .C(_0729_),
    .Y(_0730_));
 sg13g2_mux2_2 _2588_ (.A0(\GUScpu0.PC0[10] ),
    .A1(\GUScpu0.PC1[10] ),
    .S(net877),
    .X(_0731_));
 sg13g2_o21ai_1 _2589_ (.B1(net757),
    .Y(_0732_),
    .A1(net855),
    .A2(_0731_));
 sg13g2_nand2b_1 _2590_ (.Y(_0733_),
    .B(_0552_),
    .A_N(_0093_));
 sg13g2_mux2_1 _2591_ (.A0(_0034_),
    .A1(_0033_),
    .S(net845),
    .X(_0734_));
 sg13g2_o21ai_1 _2592_ (.B1(net838),
    .Y(_0735_),
    .A1(_0036_),
    .A2(net846));
 sg13g2_inv_1 _2593_ (.Y(_0736_),
    .A(_0735_));
 sg13g2_o21ai_1 _2594_ (.B1(_0736_),
    .Y(_0737_),
    .A1(_0035_),
    .A2(net828));
 sg13g2_a21oi_1 _2595_ (.A1(net827),
    .A2(_0734_),
    .Y(_0738_),
    .B1(net824));
 sg13g2_mux4_1 _2596_ (.S0(net845),
    .A0(_0030_),
    .A1(_0029_),
    .A2(_0032_),
    .A3(_0031_),
    .S1(net838),
    .X(_0739_));
 sg13g2_inv_1 _2597_ (.Y(_0740_),
    .A(_0739_));
 sg13g2_a22oi_1 _2598_ (.Y(_0741_),
    .B1(_0740_),
    .B2(net824),
    .A2(_0738_),
    .A1(_0737_));
 sg13g2_o21ai_1 _2599_ (.B1(_0733_),
    .Y(_0742_),
    .A1(net830),
    .A2(_0741_));
 sg13g2_xnor2_1 _2600_ (.Y(_0743_),
    .A(net774),
    .B(_0742_));
 sg13g2_nor3_2 _2601_ (.A(_0730_),
    .B(_0732_),
    .C(_0743_),
    .Y(_0744_));
 sg13g2_o21ai_1 _2602_ (.B1(_0743_),
    .Y(_0745_),
    .A1(_0730_),
    .A2(_0732_));
 sg13g2_inv_1 _2603_ (.Y(_0746_),
    .A(_0745_));
 sg13g2_nor2_2 _2604_ (.A(_0744_),
    .B(_0746_),
    .Y(_0747_));
 sg13g2_nand3b_1 _2605_ (.B(_0719_),
    .C(_0747_),
    .Y(_0748_),
    .A_N(_0693_));
 sg13g2_a21oi_1 _2606_ (.A1(_0662_),
    .A2(_0691_),
    .Y(_0749_),
    .B1(_0690_));
 sg13g2_nor2_1 _2607_ (.A(_0717_),
    .B(_0744_),
    .Y(_0750_));
 sg13g2_o21ai_1 _2608_ (.B1(_0750_),
    .Y(_0751_),
    .A1(_0746_),
    .A2(_0749_));
 sg13g2_nand2_1 _2609_ (.Y(_0752_),
    .A(_0718_),
    .B(_0751_));
 sg13g2_o21ai_1 _2610_ (.B1(_0752_),
    .Y(_0753_),
    .A1(_0636_),
    .A2(_0748_));
 sg13g2_xor2_1 _2611_ (.B(_1705_),
    .A(_1695_),
    .X(_0754_));
 sg13g2_inv_1 _2612_ (.Y(_0755_),
    .A(_0754_));
 sg13g2_and2_1 _2613_ (.A(_1682_),
    .B(_0755_),
    .X(_0756_));
 sg13g2_a21o_1 _2614_ (.A2(_0755_),
    .A1(_0753_),
    .B1(_1706_),
    .X(_0757_));
 sg13g2_a221oi_1 _2615_ (.B2(_0756_),
    .C1(_1681_),
    .B1(_0753_),
    .A1(_1682_),
    .Y(_0758_),
    .A2(_1706_));
 sg13g2_o21ai_1 _2616_ (.B1(_1655_),
    .Y(_0759_),
    .A1(_1656_),
    .A2(_0758_));
 sg13g2_xnor2_1 _2617_ (.Y(_0760_),
    .A(_1630_),
    .B(_0759_));
 sg13g2_nand2_1 _2618_ (.Y(_0761_),
    .A(net766),
    .B(_1626_));
 sg13g2_nor2_1 _2619_ (.A(_1552_),
    .B(_1554_),
    .Y(_0762_));
 sg13g2_nor2_1 _2620_ (.A(net758),
    .B(_0762_),
    .Y(_0763_));
 sg13g2_inv_1 _2621_ (.Y(_0764_),
    .A(net753));
 sg13g2_o21ai_1 _2622_ (.B1(_0761_),
    .Y(_0765_),
    .A1(_1630_),
    .A2(_0764_));
 sg13g2_a21o_2 _2623_ (.A2(_0760_),
    .A1(net758),
    .B1(_0765_),
    .X(_0766_));
 sg13g2_mux2_2 _2624_ (.A0(_1597_),
    .A1(_0766_),
    .S(net858),
    .X(_0767_));
 sg13g2_xnor2_1 _2625_ (.Y(_0768_),
    .A(_1656_),
    .B(_0758_));
 sg13g2_a22oi_1 _2626_ (.Y(_0769_),
    .B1(_1657_),
    .B2(net754),
    .A2(_1654_),
    .A1(net768));
 sg13g2_o21ai_1 _2627_ (.B1(_0769_),
    .Y(_0770_),
    .A1(net756),
    .A2(_0768_));
 sg13g2_or2_1 _2628_ (.X(_0771_),
    .B(_1642_),
    .A(net859));
 sg13g2_o21ai_1 _2629_ (.B1(_0771_),
    .Y(_0772_),
    .A1(net860),
    .A2(_0770_));
 sg13g2_o21ai_1 _2630_ (.B1(_0749_),
    .Y(_0773_),
    .A1(_0636_),
    .A2(_0693_));
 sg13g2_a21oi_1 _2631_ (.A1(_0747_),
    .A2(_0773_),
    .Y(_0774_),
    .B1(_0744_));
 sg13g2_xor2_1 _2632_ (.B(_0774_),
    .A(_0719_),
    .X(_0775_));
 sg13g2_a22oi_1 _2633_ (.Y(_0776_),
    .B1(_0719_),
    .B2(net754),
    .A2(_0717_),
    .A1(net767));
 sg13g2_o21ai_1 _2634_ (.B1(_0776_),
    .Y(_0777_),
    .A1(net756),
    .A2(_0775_));
 sg13g2_and2_1 _2635_ (.A(net858),
    .B(_0777_),
    .X(_0778_));
 sg13g2_and2_1 _2636_ (.A(net860),
    .B(_0705_),
    .X(_0779_));
 sg13g2_xnor2_1 _2637_ (.Y(_0780_),
    .A(_0753_),
    .B(_0755_));
 sg13g2_a22oi_1 _2638_ (.Y(_0781_),
    .B1(_0755_),
    .B2(net754),
    .A2(_1706_),
    .A1(net767));
 sg13g2_o21ai_1 _2639_ (.B1(_0781_),
    .Y(_0782_),
    .A1(net756),
    .A2(_0780_));
 sg13g2_mux2_1 _2640_ (.A0(_1693_),
    .A1(_0782_),
    .S(net858),
    .X(_0783_));
 sg13g2_and2_1 _2641_ (.A(_0531_),
    .B(_0609_),
    .X(_0784_));
 sg13g2_nand3_1 _2642_ (.B(_0609_),
    .C(_0631_),
    .A(_0531_),
    .Y(_0785_));
 sg13g2_a21oi_1 _2643_ (.A1(_0633_),
    .A2(_0785_),
    .Y(_0786_),
    .B1(_0559_));
 sg13g2_and3_1 _2644_ (.X(_0787_),
    .A(_0559_),
    .B(_0633_),
    .C(_0785_));
 sg13g2_nor3_1 _2645_ (.A(net756),
    .B(_0786_),
    .C(_0787_),
    .Y(_0788_));
 sg13g2_a22oi_1 _2646_ (.Y(_0789_),
    .B1(_0558_),
    .B2(net754),
    .A2(_0557_),
    .A1(net767));
 sg13g2_inv_1 _2647_ (.Y(_0790_),
    .A(_0789_));
 sg13g2_nor2_1 _2648_ (.A(_0788_),
    .B(_0790_),
    .Y(_0791_));
 sg13g2_o21ai_1 _2649_ (.B1(_1518_),
    .Y(_0792_),
    .A1(_0788_),
    .A2(_0790_));
 sg13g2_nand2_1 _2650_ (.Y(_0793_),
    .A(net860),
    .B(_0542_));
 sg13g2_nand2_1 _2651_ (.Y(_0794_),
    .A(_0792_),
    .B(_0793_));
 sg13g2_xnor2_1 _2652_ (.Y(_0795_),
    .A(_0636_),
    .B(_0664_));
 sg13g2_a22oi_1 _2653_ (.Y(_0796_),
    .B1(_0665_),
    .B2(net754),
    .A2(_0662_),
    .A1(net767));
 sg13g2_o21ai_1 _2654_ (.B1(_0796_),
    .Y(_0797_),
    .A1(net755),
    .A2(_0795_));
 sg13g2_or2_1 _2655_ (.X(_0798_),
    .B(_0648_),
    .A(net859));
 sg13g2_o21ai_1 _2656_ (.B1(_0798_),
    .Y(_0799_),
    .A1(net860),
    .A2(_0797_));
 sg13g2_nand3_1 _2657_ (.B(_0793_),
    .C(_0799_),
    .A(_0792_),
    .Y(_0800_));
 sg13g2_xnor2_1 _2658_ (.Y(_0801_),
    .A(_0747_),
    .B(_0773_));
 sg13g2_a22oi_1 _2659_ (.Y(_0802_),
    .B1(_0747_),
    .B2(net753),
    .A2(_0744_),
    .A1(net767));
 sg13g2_o21ai_1 _2660_ (.B1(_0802_),
    .Y(_0803_),
    .A1(net755),
    .A2(_0801_));
 sg13g2_mux2_1 _2661_ (.A0(_0731_),
    .A1(_0803_),
    .S(net858),
    .X(_0804_));
 sg13g2_o21ai_1 _2662_ (.B1(_0663_),
    .Y(_0805_),
    .A1(_0636_),
    .A2(_0664_));
 sg13g2_xnor2_1 _2663_ (.Y(_0806_),
    .A(_0692_),
    .B(_0805_));
 sg13g2_nor2_1 _2664_ (.A(_0692_),
    .B(_0764_),
    .Y(_0807_));
 sg13g2_a221oi_1 _2665_ (.B2(net758),
    .C1(_0807_),
    .B1(_0806_),
    .A1(net767),
    .Y(_0808_),
    .A2(_0690_));
 sg13g2_nor2_1 _2666_ (.A(net858),
    .B(_0677_),
    .Y(_0809_));
 sg13g2_a21oi_1 _2667_ (.A1(net859),
    .A2(_0808_),
    .Y(_0810_),
    .B1(_0809_));
 sg13g2_nor4_1 _2668_ (.A(_0783_),
    .B(_0800_),
    .C(_0804_),
    .D(_0810_),
    .Y(_0811_));
 sg13g2_a221oi_1 _2669_ (.B2(_0756_),
    .C1(net755),
    .B1(_0753_),
    .A1(_1682_),
    .Y(_0812_),
    .A2(_1706_));
 sg13g2_o21ai_1 _2670_ (.B1(_0812_),
    .Y(_0813_),
    .A1(_1682_),
    .A2(_0757_));
 sg13g2_nand2_1 _2671_ (.Y(_0814_),
    .A(net767),
    .B(_1681_));
 sg13g2_nand2_1 _2672_ (.Y(_0815_),
    .A(_1682_),
    .B(net753));
 sg13g2_nand3_1 _2673_ (.B(_0814_),
    .C(_0815_),
    .A(_0813_),
    .Y(_0816_));
 sg13g2_or2_1 _2674_ (.X(_0817_),
    .B(_1668_),
    .A(net858));
 sg13g2_o21ai_1 _2675_ (.B1(_0817_),
    .Y(_0818_),
    .A1(net860),
    .A2(_0816_));
 sg13g2_o21ai_1 _2676_ (.B1(_0584_),
    .Y(_0819_),
    .A1(_0557_),
    .A2(_0786_));
 sg13g2_or3_1 _2677_ (.A(_0557_),
    .B(_0584_),
    .C(_0786_),
    .X(_0820_));
 sg13g2_nand3_1 _2678_ (.B(_0819_),
    .C(_0820_),
    .A(net758),
    .Y(_0821_));
 sg13g2_a22oi_1 _2679_ (.Y(_0822_),
    .B1(_0584_),
    .B2(net754),
    .A2(_0582_),
    .A1(net767));
 sg13g2_nand2_1 _2680_ (.Y(_0823_),
    .A(_0821_),
    .B(_0822_));
 sg13g2_nand3_1 _2681_ (.B(_0821_),
    .C(_0822_),
    .A(net857),
    .Y(_0824_));
 sg13g2_or2_1 _2682_ (.X(_0825_),
    .B(_0569_),
    .A(net858));
 sg13g2_nand2_1 _2683_ (.Y(_0826_),
    .A(_0824_),
    .B(_0825_));
 sg13g2_a221oi_1 _2684_ (.B2(_0825_),
    .C1(_0779_),
    .B1(_0824_),
    .A1(net858),
    .Y(_0827_),
    .A2(_0777_));
 sg13g2_nand4_1 _2685_ (.B(_0811_),
    .C(_0818_),
    .A(_0772_),
    .Y(_0828_),
    .D(_0827_));
 sg13g2_or2_1 _2686_ (.X(_0829_),
    .B(_0828_),
    .A(_0767_));
 sg13g2_nor2_1 _2687_ (.A(net857),
    .B(_0615_),
    .Y(_0830_));
 sg13g2_o21ai_1 _2688_ (.B1(_0631_),
    .Y(_0831_),
    .A1(_0608_),
    .A2(_0784_));
 sg13g2_or3_1 _2689_ (.A(_0608_),
    .B(_0631_),
    .C(_0784_),
    .X(_0832_));
 sg13g2_and3_1 _2690_ (.X(_0833_),
    .A(_1555_),
    .B(_0831_),
    .C(_0832_));
 sg13g2_a221oi_1 _2691_ (.B2(net753),
    .C1(_0833_),
    .B1(_0631_),
    .A1(net766),
    .Y(_0834_),
    .A2(_0630_));
 sg13g2_a21oi_2 _2692_ (.B1(_0830_),
    .Y(_0835_),
    .A2(_0834_),
    .A1(net857));
 sg13g2_inv_1 _2693_ (.Y(_0836_),
    .A(_0835_));
 sg13g2_nor3_1 _2694_ (.A(_0767_),
    .B(_0828_),
    .C(_0836_),
    .Y(_0837_));
 sg13g2_a21oi_1 _2695_ (.A1(_0468_),
    .A2(_0473_),
    .Y(_0838_),
    .B1(net755));
 sg13g2_o21ai_1 _2696_ (.B1(_0838_),
    .Y(_0839_),
    .A1(_0468_),
    .A2(_0473_));
 sg13g2_a22oi_1 _2697_ (.Y(_0840_),
    .B1(_0468_),
    .B2(net753),
    .A2(_0466_),
    .A1(net766));
 sg13g2_nand2_1 _2698_ (.Y(_0841_),
    .A(_0839_),
    .B(_0840_));
 sg13g2_a21oi_2 _2699_ (.B1(net861),
    .Y(_0842_),
    .A2(_0840_),
    .A1(_0839_));
 sg13g2_nand2_2 _2700_ (.Y(_0843_),
    .A(net861),
    .B(_0454_));
 sg13g2_nand2b_2 _2701_ (.Y(_0844_),
    .B(_0843_),
    .A_N(_0842_));
 sg13g2_nor2b_2 _2702_ (.A(_0842_),
    .B_N(_0843_),
    .Y(_0845_));
 sg13g2_xnor2_1 _2703_ (.Y(_0846_),
    .A(_0475_),
    .B(_0501_));
 sg13g2_and2_1 _2704_ (.A(_0501_),
    .B(net753),
    .X(_0847_));
 sg13g2_a221oi_1 _2705_ (.B2(net758),
    .C1(_0847_),
    .B1(_0846_),
    .A1(net766),
    .Y(_0848_),
    .A2(_0500_));
 sg13g2_nor2_1 _2706_ (.A(net861),
    .B(_0848_),
    .Y(_0849_));
 sg13g2_nand2_1 _2707_ (.Y(_0850_),
    .A(net860),
    .B(_0489_));
 sg13g2_nor2b_2 _2708_ (.A(_0849_),
    .B_N(_0850_),
    .Y(_0851_));
 sg13g2_o21ai_1 _2709_ (.B1(_0850_),
    .Y(_0852_),
    .A1(net861),
    .A2(_0848_));
 sg13g2_xnor2_1 _2710_ (.Y(_0853_),
    .A(_0444_),
    .B(_0474_));
 sg13g2_a22oi_1 _2711_ (.Y(_0854_),
    .B1(_0444_),
    .B2(net753),
    .A2(_0443_),
    .A1(net766));
 sg13g2_o21ai_1 _2712_ (.B1(_0854_),
    .Y(_0855_),
    .A1(net755),
    .A2(_0853_));
 sg13g2_nor2_1 _2713_ (.A(net857),
    .B(_0429_),
    .Y(_0856_));
 sg13g2_a21oi_2 _2714_ (.B1(_0856_),
    .Y(_0857_),
    .A2(_0855_),
    .A1(net857));
 sg13g2_inv_2 _2715_ (.Y(_0858_),
    .A(net736));
 sg13g2_nor2_1 _2716_ (.A(net735),
    .B(net736),
    .Y(_0859_));
 sg13g2_nand2_1 _2717_ (.Y(_0860_),
    .A(_0845_),
    .B(_0858_));
 sg13g2_nor2_1 _2718_ (.A(net735),
    .B(_0860_),
    .Y(_0861_));
 sg13g2_nand4_1 _2719_ (.B(_1511_),
    .C(net722),
    .A(_0077_),
    .Y(_0862_),
    .D(net733));
 sg13g2_nor4_2 _2720_ (.A(\uart0.txbitcnt[3] ),
    .B(\uart0.txbitcnt[2] ),
    .C(\uart0.txbitcnt[1] ),
    .Y(_0863_),
    .D(\uart0.txbitcnt[0] ));
 sg13g2_and2_2 _2721_ (.A(net867),
    .B(net723),
    .X(_0864_));
 sg13g2_nand2b_1 _2722_ (.Y(_0865_),
    .B(_0864_),
    .A_N(_0860_));
 sg13g2_or2_1 _2723_ (.X(_0866_),
    .B(_0865_),
    .A(net735));
 sg13g2_o21ai_1 _2724_ (.B1(_0862_),
    .Y(_0867_),
    .A1(_0863_),
    .A2(_0866_));
 sg13g2_nand4_1 _2725_ (.B(_1511_),
    .C(net722),
    .A(_1497_),
    .Y(_0868_),
    .D(net733));
 sg13g2_nand3_1 _2726_ (.B(net886),
    .C(_0868_),
    .A(\uart0.rxoverr ),
    .Y(_0869_));
 sg13g2_o21ai_1 _2727_ (.B1(_0869_),
    .Y(_0390_),
    .A1(_1460_),
    .A2(net886));
 sg13g2_nand2_1 _2728_ (.Y(_0870_),
    .A(\uart0.rxvalid ),
    .B(_0868_));
 sg13g2_nand2_1 _2729_ (.Y(_0389_),
    .A(net886),
    .B(_0870_));
 sg13g2_mux2_1 _2730_ (.A0(\uart0.urxsh[9] ),
    .A1(\uart0.urxbuffer[8] ),
    .S(net887),
    .X(_0388_));
 sg13g2_mux2_1 _2731_ (.A0(\uart0.urxsh[8] ),
    .A1(\uart0.q[7] ),
    .S(net887),
    .X(_0387_));
 sg13g2_mux2_1 _2732_ (.A0(\uart0.urxsh[7] ),
    .A1(\uart0.q[6] ),
    .S(net887),
    .X(_0386_));
 sg13g2_mux2_1 _2733_ (.A0(\uart0.urxsh[6] ),
    .A1(\uart0.q[5] ),
    .S(net887),
    .X(_0385_));
 sg13g2_mux2_1 _2734_ (.A0(\uart0.urxsh[5] ),
    .A1(\uart0.q[4] ),
    .S(net887),
    .X(_0384_));
 sg13g2_mux2_1 _2735_ (.A0(\uart0.urxsh[4] ),
    .A1(\uart0.q[3] ),
    .S(net886),
    .X(_0383_));
 sg13g2_mux2_1 _2736_ (.A0(\uart0.urxsh[3] ),
    .A1(\uart0.q[2] ),
    .S(net886),
    .X(_0382_));
 sg13g2_mux2_1 _2737_ (.A0(\uart0.urxsh[2] ),
    .A1(\uart0.q[1] ),
    .S(net886),
    .X(_0381_));
 sg13g2_mux2_1 _2738_ (.A0(\uart0.urxsh[1] ),
    .A1(\uart0.q[0] ),
    .S(net886),
    .X(_0380_));
 sg13g2_and2_1 _2739_ (.A(\uart0.txdiv[0] ),
    .B(\uart0.txdiv[1] ),
    .X(_0871_));
 sg13g2_nor2_1 _2740_ (.A(\uart0.txdiv[3] ),
    .B(\uart0.txdiv[2] ),
    .Y(_0872_));
 sg13g2_and4_1 _2741_ (.A(\uart0.txdiv[4] ),
    .B(\uart0.txdiv[5] ),
    .C(_0871_),
    .D(_0872_),
    .X(_0873_));
 sg13g2_nand4_1 _2742_ (.B(\uart0.txdiv[5] ),
    .C(_0871_),
    .A(\uart0.txdiv[4] ),
    .Y(_0874_),
    .D(_0872_));
 sg13g2_nor3_1 _2743_ (.A(\uart0.txbitcnt[1] ),
    .B(\uart0.txbitcnt[0] ),
    .C(_0874_),
    .Y(_0875_));
 sg13g2_nor2b_1 _2744_ (.A(\uart0.txbitcnt[2] ),
    .B_N(_0875_),
    .Y(_0876_));
 sg13g2_and4_1 _2745_ (.A(net867),
    .B(net722),
    .C(net733),
    .D(_0863_),
    .X(_0877_));
 sg13g2_nand4_1 _2746_ (.B(net722),
    .C(net733),
    .A(net867),
    .Y(_0878_),
    .D(_0863_));
 sg13g2_o21ai_1 _2747_ (.B1(_0878_),
    .Y(_0379_),
    .A1(_1461_),
    .A2(_0876_));
 sg13g2_nor2b_1 _2748_ (.A(_0875_),
    .B_N(\uart0.txbitcnt[2] ),
    .Y(_0879_));
 sg13g2_a21o_1 _2749_ (.A2(_0876_),
    .A1(\uart0.txbitcnt[3] ),
    .B1(_0879_),
    .X(_0378_));
 sg13g2_nor2_2 _2750_ (.A(net868),
    .B(net719),
    .Y(_0880_));
 sg13g2_nand2_1 _2751_ (.Y(_0881_),
    .A(_0874_),
    .B(_0878_));
 sg13g2_o21ai_1 _2752_ (.B1(_0878_),
    .Y(_0882_),
    .A1(_0863_),
    .A2(_0874_));
 sg13g2_nand2b_1 _2753_ (.Y(_0883_),
    .B(_0882_),
    .A_N(\uart0.txbitcnt[0] ));
 sg13g2_xnor2_1 _2754_ (.Y(_0377_),
    .A(\uart0.txbitcnt[1] ),
    .B(_0883_));
 sg13g2_nand2b_1 _2755_ (.Y(_0884_),
    .B(\uart0.txbitcnt[0] ),
    .A_N(_0882_));
 sg13g2_o21ai_1 _2756_ (.B1(_0884_),
    .Y(_0376_),
    .A1(net719),
    .A2(_0883_));
 sg13g2_nand4_1 _2757_ (.B(\uart0.rxdiv[0] ),
    .C(\uart0.rxdiv[3] ),
    .A(_1498_),
    .Y(_0885_),
    .D(\uart0.rxdiv[4] ));
 sg13g2_nor3_1 _2758_ (.A(\uart0.rxdiv[2] ),
    .B(\uart0.rxdiv[5] ),
    .C(_0885_),
    .Y(_0886_));
 sg13g2_nor2b_1 _2759_ (.A(_0886_),
    .B_N(net887),
    .Y(_0887_));
 sg13g2_nand2_1 _2760_ (.Y(_0888_),
    .A(_0190_),
    .B(net834));
 sg13g2_nand2_1 _2761_ (.Y(_0889_),
    .A(net886),
    .B(_0886_));
 sg13g2_o21ai_1 _2762_ (.B1(_0888_),
    .Y(_0375_),
    .A1(\uart0.rxreg[1] ),
    .A2(net833));
 sg13g2_nand2_1 _2763_ (.Y(_0890_),
    .A(_0189_),
    .B(_0887_));
 sg13g2_o21ai_1 _2764_ (.B1(_0890_),
    .Y(_0374_),
    .A1(\uart0.urxsh[9] ),
    .A2(_0889_));
 sg13g2_nand2_1 _2765_ (.Y(_0891_),
    .A(_0188_),
    .B(net834));
 sg13g2_o21ai_1 _2766_ (.B1(_0891_),
    .Y(_0373_),
    .A1(\uart0.urxsh[8] ),
    .A2(net833));
 sg13g2_nand2_1 _2767_ (.Y(_0892_),
    .A(_0187_),
    .B(net834));
 sg13g2_o21ai_1 _2768_ (.B1(_0892_),
    .Y(_0372_),
    .A1(\uart0.urxsh[7] ),
    .A2(net833));
 sg13g2_nand2_1 _2769_ (.Y(_0893_),
    .A(_0186_),
    .B(net834));
 sg13g2_o21ai_1 _2770_ (.B1(_0893_),
    .Y(_0371_),
    .A1(\uart0.urxsh[6] ),
    .A2(_0889_));
 sg13g2_nand2_1 _2771_ (.Y(_0894_),
    .A(_0185_),
    .B(net834));
 sg13g2_o21ai_1 _2772_ (.B1(_0894_),
    .Y(_0370_),
    .A1(\uart0.urxsh[5] ),
    .A2(net833));
 sg13g2_nand2_1 _2773_ (.Y(_0895_),
    .A(_0184_),
    .B(net834));
 sg13g2_o21ai_1 _2774_ (.B1(_0895_),
    .Y(_0369_),
    .A1(\uart0.urxsh[4] ),
    .A2(net833));
 sg13g2_nand2_1 _2775_ (.Y(_0896_),
    .A(_0183_),
    .B(net834));
 sg13g2_o21ai_1 _2776_ (.B1(_0896_),
    .Y(_0368_),
    .A1(\uart0.urxsh[3] ),
    .A2(net833));
 sg13g2_nand2_1 _2777_ (.Y(_0897_),
    .A(_0182_),
    .B(net834));
 sg13g2_o21ai_1 _2778_ (.B1(_0897_),
    .Y(_0367_),
    .A1(\uart0.urxsh[2] ),
    .A2(net833));
 sg13g2_nor2_1 _2779_ (.A(\uart0.urxsh[1] ),
    .B(net833),
    .Y(_0191_));
 sg13g2_nor4_1 _2780_ (.A(\pwmc[5] ),
    .B(\pwmc[4] ),
    .C(\pwmc[7] ),
    .D(\pwmc[6] ),
    .Y(_0898_));
 sg13g2_nor2_1 _2781_ (.A(\pwmc[0] ),
    .B(\pwmc[1] ),
    .Y(_0899_));
 sg13g2_nand4_1 _2782_ (.B(_1467_),
    .C(_0898_),
    .A(_1466_),
    .Y(_0900_),
    .D(_0899_));
 sg13g2_nor2_2 _2783_ (.A(_0845_),
    .B(_0852_),
    .Y(_0901_));
 sg13g2_and2_2 _2784_ (.A(net736),
    .B(_0901_),
    .X(_0902_));
 sg13g2_nand2_1 _2785_ (.Y(_0903_),
    .A(_0857_),
    .B(_0901_));
 sg13g2_and2_1 _2786_ (.A(_0864_),
    .B(_0902_),
    .X(_0904_));
 sg13g2_o21ai_1 _2787_ (.B1(_0900_),
    .Y(_0272_),
    .A1(_1462_),
    .A2(_0904_));
 sg13g2_nand2b_1 _2788_ (.Y(_0905_),
    .B(\pwmc[2] ),
    .A_N(\pwmbuf[2] ));
 sg13g2_xnor2_1 _2789_ (.Y(_0906_),
    .A(\pwmbuf[7] ),
    .B(\pwmc[7] ));
 sg13g2_a22oi_1 _2790_ (.Y(_0907_),
    .B1(_1467_),
    .B2(\pwmbuf[2] ),
    .A2(_1466_),
    .A1(\pwmbuf[3] ));
 sg13g2_nand2b_1 _2791_ (.Y(_0908_),
    .B(\pwmbuf[4] ),
    .A_N(\pwmc[4] ));
 sg13g2_nand2b_1 _2792_ (.Y(_0909_),
    .B(\pwmc[3] ),
    .A_N(\pwmbuf[3] ));
 sg13g2_o21ai_1 _2793_ (.B1(_0908_),
    .Y(_0910_),
    .A1(_1465_),
    .A2(\pwmc[1] ));
 sg13g2_xor2_1 _2794_ (.B(\pwmc[0] ),
    .A(\pwmbuf[0] ),
    .X(_0911_));
 sg13g2_xor2_1 _2795_ (.B(\pwmc[5] ),
    .A(\pwmbuf[5] ),
    .X(_0912_));
 sg13g2_xor2_1 _2796_ (.B(\pwmc[6] ),
    .A(\pwmbuf[6] ),
    .X(_0913_));
 sg13g2_nor4_1 _2797_ (.A(_0910_),
    .B(_0911_),
    .C(_0912_),
    .D(_0913_),
    .Y(_0914_));
 sg13g2_nand4_1 _2798_ (.B(_0906_),
    .C(_0907_),
    .A(_0905_),
    .Y(_0915_),
    .D(_0909_));
 sg13g2_a221oi_1 _2799_ (.B2(_1464_),
    .C1(_0915_),
    .B1(\pwmc[4] ),
    .A1(_1465_),
    .Y(_0916_),
    .A2(\pwmc[1] ));
 sg13g2_a22oi_1 _2800_ (.Y(_0271_),
    .B1(_0914_),
    .B2(_0916_),
    .A2(_0900_),
    .A1(_1463_));
 sg13g2_nand4_1 _2801_ (.B(\pwmc[3] ),
    .C(\pwmc[2] ),
    .A(\pwmc[1] ),
    .Y(_0917_),
    .D(\pwmc[5] ));
 sg13g2_nand2_1 _2802_ (.Y(_0918_),
    .A(\pwmc[4] ),
    .B(\pwmc[6] ));
 sg13g2_nand2_1 _2803_ (.Y(_0919_),
    .A(\pwmc[7] ),
    .B(net936));
 sg13g2_nor3_2 _2804_ (.A(_0917_),
    .B(_0918_),
    .C(_0919_),
    .Y(_0920_));
 sg13g2_mux2_1 _2805_ (.A0(\pwmbuf[7] ),
    .A1(\pwmhold[7] ),
    .S(_0920_),
    .X(_0270_));
 sg13g2_mux2_1 _2806_ (.A0(\pwmbuf[6] ),
    .A1(\pwmhold[6] ),
    .S(_0920_),
    .X(_0269_));
 sg13g2_mux2_1 _2807_ (.A0(\pwmbuf[5] ),
    .A1(\pwmhold[5] ),
    .S(_0920_),
    .X(_0268_));
 sg13g2_mux2_1 _2808_ (.A0(\pwmbuf[4] ),
    .A1(\pwmhold[4] ),
    .S(_0920_),
    .X(_0267_));
 sg13g2_mux2_1 _2809_ (.A0(\pwmbuf[3] ),
    .A1(\pwmhold[3] ),
    .S(_0920_),
    .X(_0266_));
 sg13g2_mux2_1 _2810_ (.A0(\pwmbuf[2] ),
    .A1(\pwmhold[2] ),
    .S(_0920_),
    .X(_0265_));
 sg13g2_mux2_1 _2811_ (.A0(\pwmbuf[1] ),
    .A1(\pwmhold[1] ),
    .S(_0920_),
    .X(_0264_));
 sg13g2_mux2_1 _2812_ (.A0(\pwmbuf[0] ),
    .A1(\pwmhold[0] ),
    .S(_0920_),
    .X(_0263_));
 sg13g2_and2_1 _2813_ (.A(_0180_),
    .B(_0880_),
    .X(_0921_));
 sg13g2_a21o_1 _2814_ (.A2(net718),
    .A1(_0579_),
    .B1(_0921_),
    .X(_0261_));
 sg13g2_nor2_1 _2815_ (.A(_0179_),
    .B(net868),
    .Y(_0922_));
 sg13g2_a21oi_1 _2816_ (.A1(\uart0.txsh[8] ),
    .A2(net868),
    .Y(_0923_),
    .B1(_0922_));
 sg13g2_nor2_1 _2817_ (.A(net718),
    .B(_0923_),
    .Y(_0924_));
 sg13g2_a21oi_1 _2818_ (.A1(_0551_),
    .A2(net718),
    .Y(_0260_),
    .B1(_0924_));
 sg13g2_nor3_1 _2819_ (.A(\uart0.txsh[7] ),
    .B(_0874_),
    .C(net719),
    .Y(_0925_));
 sg13g2_a22oi_1 _2820_ (.Y(_0926_),
    .B1(_0880_),
    .B2(_0178_),
    .A2(net718),
    .A1(_0624_));
 sg13g2_nand2b_1 _2821_ (.Y(_0259_),
    .B(_0926_),
    .A_N(_0925_));
 sg13g2_nor2_1 _2822_ (.A(_0177_),
    .B(net868),
    .Y(_0927_));
 sg13g2_a21oi_1 _2823_ (.A1(\uart0.txsh[6] ),
    .A2(net868),
    .Y(_0928_),
    .B1(_0927_));
 sg13g2_mux2_1 _2824_ (.A0(_0605_),
    .A1(_0928_),
    .S(_0878_),
    .X(_0258_));
 sg13g2_nor2_1 _2825_ (.A(_0176_),
    .B(net869),
    .Y(_0929_));
 sg13g2_a21oi_1 _2826_ (.A1(\uart0.txsh[5] ),
    .A2(net868),
    .Y(_0930_),
    .B1(_0929_));
 sg13g2_nor2_1 _2827_ (.A(net718),
    .B(_0930_),
    .Y(_0931_));
 sg13g2_a21oi_1 _2828_ (.A1(_0521_),
    .A2(net718),
    .Y(_0257_),
    .B1(_0931_));
 sg13g2_nor2_1 _2829_ (.A(_0175_),
    .B(net868),
    .Y(_0932_));
 sg13g2_a21oi_1 _2830_ (.A1(\uart0.txsh[4] ),
    .A2(net868),
    .Y(_0933_),
    .B1(_0932_));
 sg13g2_mux2_1 _2831_ (.A0(_0497_),
    .A1(_0933_),
    .S(_0878_),
    .X(_0256_));
 sg13g2_nor3_1 _2832_ (.A(\uart0.txsh[3] ),
    .B(_0874_),
    .C(net718),
    .Y(_0934_));
 sg13g2_a22oi_1 _2833_ (.Y(_0935_),
    .B1(_0880_),
    .B2(_0174_),
    .A2(net719),
    .A1(_0439_));
 sg13g2_nand2b_1 _2834_ (.Y(_0255_),
    .B(_0935_),
    .A_N(_0934_));
 sg13g2_nor2_1 _2835_ (.A(_0173_),
    .B(net869),
    .Y(_0936_));
 sg13g2_a21oi_1 _2836_ (.A1(\uart0.txsh[2] ),
    .A2(net869),
    .Y(_0937_),
    .B1(_0936_));
 sg13g2_nor2_1 _2837_ (.A(net719),
    .B(_0937_),
    .Y(_0938_));
 sg13g2_a21oi_1 _2838_ (.A1(_0463_),
    .A2(net719),
    .Y(_0254_),
    .B1(_0938_));
 sg13g2_nand2_1 _2839_ (.Y(_0939_),
    .A(\uart0.txsh[1] ),
    .B(net869));
 sg13g2_o21ai_1 _2840_ (.B1(_0939_),
    .Y(_0940_),
    .A1(_0172_),
    .A2(net869));
 sg13g2_nand2_1 _2841_ (.Y(_0253_),
    .A(_0878_),
    .B(_0940_));
 sg13g2_nor2b_1 _2842_ (.A(net230),
    .B_N(net935),
    .Y(xlah));
 sg13g2_nor2_1 _2843_ (.A(_0845_),
    .B(_0851_),
    .Y(_0941_));
 sg13g2_nor2_2 _2844_ (.A(_0851_),
    .B(_0857_),
    .Y(_0942_));
 sg13g2_nor3_1 _2845_ (.A(_0845_),
    .B(_0851_),
    .C(net736),
    .Y(_0943_));
 sg13g2_inv_1 _2846_ (.Y(_0944_),
    .A(net732));
 sg13g2_nor4_2 _2847_ (.A(_0767_),
    .B(_0828_),
    .C(_0836_),
    .Y(_0945_),
    .D(_0944_));
 sg13g2_nand2_1 _2848_ (.Y(_0946_),
    .A(\GUScpu0.PC0[15] ),
    .B(_0945_));
 sg13g2_nor3_2 _2849_ (.A(_0767_),
    .B(_0828_),
    .C(_0835_),
    .Y(_0947_));
 sg13g2_o21ai_1 _2850_ (.B1(net755),
    .Y(_0948_),
    .A1(_0528_),
    .A2(_0762_));
 sg13g2_a21oi_1 _2851_ (.A1(net766),
    .A2(_0525_),
    .Y(_0949_),
    .B1(_0948_));
 sg13g2_a21oi_1 _2852_ (.A1(_0476_),
    .A2(_0501_),
    .Y(_0950_),
    .B1(_0500_));
 sg13g2_o21ai_1 _2853_ (.B1(net758),
    .Y(_0951_),
    .A1(_0527_),
    .A2(_0950_));
 sg13g2_a21oi_1 _2854_ (.A1(_0527_),
    .A2(_0950_),
    .Y(_0952_),
    .B1(_0951_));
 sg13g2_nor2_2 _2855_ (.A(_0949_),
    .B(_0952_),
    .Y(_0953_));
 sg13g2_mux2_2 _2856_ (.A0(_0511_),
    .A1(_0953_),
    .S(net857),
    .X(_0954_));
 sg13g2_inv_1 _2857_ (.Y(_0955_),
    .A(_0954_));
 sg13g2_xnor2_1 _2858_ (.Y(_0956_),
    .A(_0531_),
    .B(_0609_));
 sg13g2_a22oi_1 _2859_ (.Y(_0957_),
    .B1(_0609_),
    .B2(net753),
    .A2(_0608_),
    .A1(net768));
 sg13g2_o21ai_1 _2860_ (.B1(_0957_),
    .Y(_0958_),
    .A1(net755),
    .A2(_0956_));
 sg13g2_nor2_1 _2861_ (.A(net860),
    .B(_0958_),
    .Y(_0959_));
 sg13g2_or2_1 _2862_ (.X(_0960_),
    .B(_0596_),
    .A(net859));
 sg13g2_nor2b_1 _2863_ (.A(_0959_),
    .B_N(_0960_),
    .Y(_0961_));
 sg13g2_o21ai_1 _2864_ (.B1(_0960_),
    .Y(_0962_),
    .A1(net860),
    .A2(_0958_));
 sg13g2_nor2_2 _2865_ (.A(_0955_),
    .B(net730),
    .Y(_0963_));
 sg13g2_nand2_2 _2866_ (.Y(_0964_),
    .A(_0954_),
    .B(_0962_));
 sg13g2_nor2_1 _2867_ (.A(_0954_),
    .B(net729),
    .Y(_0965_));
 sg13g2_nand2_1 _2868_ (.Y(_0966_),
    .A(_0859_),
    .B(_0965_));
 sg13g2_o21ai_1 _2869_ (.B1(_0966_),
    .Y(_0967_),
    .A1(_0944_),
    .A2(_0964_));
 sg13g2_and2_1 _2870_ (.A(_0844_),
    .B(_0967_),
    .X(_0968_));
 sg13g2_a22oi_1 _2871_ (.Y(_0969_),
    .B1(net721),
    .B2(_0968_),
    .A2(net724),
    .A1(net16));
 sg13g2_nand2_2 _2872_ (.Y(\GUScpu0.cdi[15] ),
    .A(_0946_),
    .B(_0969_));
 sg13g2_nor2_2 _2873_ (.A(net935),
    .B(\ckd[1] ),
    .Y(xlal));
 sg13g2_nand2_2 _2874_ (.Y(_0970_),
    .A(_0845_),
    .B(net735));
 sg13g2_a21oi_1 _2875_ (.A1(_0844_),
    .A2(_0858_),
    .Y(_0971_),
    .B1(net735));
 sg13g2_nand2_1 _2876_ (.Y(_0972_),
    .A(_0845_),
    .B(_0857_));
 sg13g2_inv_1 _2877_ (.Y(_0973_),
    .A(_0972_));
 sg13g2_xnor2_1 _2878_ (.Y(_0974_),
    .A(_0844_),
    .B(net736));
 sg13g2_and2_1 _2879_ (.A(_0851_),
    .B(_0974_),
    .X(_0975_));
 sg13g2_nand2_1 _2880_ (.Y(_0976_),
    .A(_0851_),
    .B(_0974_));
 sg13g2_nand2_1 _2881_ (.Y(_0977_),
    .A(_0970_),
    .B(_0976_));
 sg13g2_nor2_2 _2882_ (.A(_0942_),
    .B(_0977_),
    .Y(_0978_));
 sg13g2_nor2_2 _2883_ (.A(net736),
    .B(_0970_),
    .Y(_0979_));
 sg13g2_a22oi_1 _2884_ (.Y(_0980_),
    .B1(_0979_),
    .B2(\GUScpu0.flag0[0] ),
    .A2(net733),
    .A1(\uart0.q[0] ));
 sg13g2_nor2_1 _2885_ (.A(_0851_),
    .B(_0972_),
    .Y(_0981_));
 sg13g2_a22oi_1 _2886_ (.Y(_0982_),
    .B1(net727),
    .B2(gpo),
    .A2(net731),
    .A1(\GUScpu0.PC0[0] ));
 sg13g2_a22oi_1 _2887_ (.Y(_0983_),
    .B1(_0978_),
    .B2(\irqen[0] ),
    .A2(_0902_),
    .A1(_1497_));
 sg13g2_nand4_1 _2888_ (.B(_0980_),
    .C(_0982_),
    .A(net722),
    .Y(_0984_),
    .D(_0983_));
 sg13g2_nand2_1 _2889_ (.Y(_0985_),
    .A(net730),
    .B(_0970_));
 sg13g2_a22oi_1 _2890_ (.Y(_0986_),
    .B1(net728),
    .B2(_0962_),
    .A2(_0971_),
    .A1(net726));
 sg13g2_nand2_1 _2891_ (.Y(_0987_),
    .A(_0985_),
    .B(_0986_));
 sg13g2_nand2_1 _2892_ (.Y(_0988_),
    .A(net721),
    .B(_0987_));
 sg13g2_nand2b_1 _2893_ (.Y(_0989_),
    .B(_0829_),
    .A_N(\xdi[0] ));
 sg13g2_and3_2 _2894_ (.X(\GUScpu0.cdi[0] ),
    .A(_0984_),
    .B(_0988_),
    .C(_0989_));
 sg13g2_a22oi_1 _2895_ (.Y(_0990_),
    .B1(net727),
    .B2(net1),
    .A2(_0979_),
    .A1(\GUScpu0.cv[0][1] ));
 sg13g2_a22oi_1 _2896_ (.Y(_0991_),
    .B1(net731),
    .B2(\GUScpu0.PC0[1] ),
    .A2(net733),
    .A1(\uart0.q[1] ));
 sg13g2_a22oi_1 _2897_ (.Y(_0992_),
    .B1(_0978_),
    .B2(\irqen[1] ),
    .A2(_0902_),
    .A1(_0863_));
 sg13g2_nand4_1 _2898_ (.B(_0990_),
    .C(_0991_),
    .A(net722),
    .Y(_0993_),
    .D(_0992_));
 sg13g2_o21ai_1 _2899_ (.B1(_0963_),
    .Y(_0994_),
    .A1(_0902_),
    .A2(net731));
 sg13g2_nor2b_2 _2900_ (.A(_0901_),
    .B_N(_0970_),
    .Y(_0995_));
 sg13g2_nand3_1 _2901_ (.B(net726),
    .C(_0995_),
    .A(net736),
    .Y(_0996_));
 sg13g2_nor2_1 _2902_ (.A(net735),
    .B(_0972_),
    .Y(_0997_));
 sg13g2_o21ai_1 _2903_ (.B1(net729),
    .Y(_0998_),
    .A1(_0941_),
    .A2(_0997_));
 sg13g2_inv_1 _2904_ (.Y(_0999_),
    .A(_0998_));
 sg13g2_nand4_1 _2905_ (.B(_0994_),
    .C(_0996_),
    .A(net721),
    .Y(_1000_),
    .D(_0998_));
 sg13g2_nand2_1 _2906_ (.Y(_1001_),
    .A(_1499_),
    .B(net724));
 sg13g2_and3_1 _2907_ (.X(\GUScpu0.cdi[1] ),
    .A(_0993_),
    .B(_1000_),
    .C(_1001_));
 sg13g2_a21oi_1 _2908_ (.A1(_0858_),
    .A2(_0901_),
    .Y(_1002_),
    .B1(_0985_));
 sg13g2_nor3_1 _2909_ (.A(_0859_),
    .B(_0954_),
    .C(net729),
    .Y(_1003_));
 sg13g2_nor2_1 _2910_ (.A(_1002_),
    .B(_1003_),
    .Y(_1004_));
 sg13g2_o21ai_1 _2911_ (.B1(_1004_),
    .Y(_1005_),
    .A1(_0901_),
    .A2(_0964_));
 sg13g2_a22oi_1 _2912_ (.Y(_1006_),
    .B1(net727),
    .B2(net2),
    .A2(net734),
    .A1(\uart0.q[2] ));
 sg13g2_a22oi_1 _2913_ (.Y(_1007_),
    .B1(_0979_),
    .B2(\GUScpu0.flag0[2] ),
    .A2(net731),
    .A1(\GUScpu0.PC0[2] ));
 sg13g2_a22oi_1 _2914_ (.Y(_1008_),
    .B1(_0978_),
    .B2(\irqen[2] ),
    .A2(_0902_),
    .A1(\uart0.rxoverr ));
 sg13g2_and4_1 _2915_ (.A(net722),
    .B(_1006_),
    .C(_1007_),
    .D(_1008_),
    .X(_1009_));
 sg13g2_a221oi_1 _2916_ (.B2(_1005_),
    .C1(_1009_),
    .B1(net721),
    .A1(_1500_),
    .Y(\GUScpu0.cdi[2] ),
    .A2(net725));
 sg13g2_a22oi_1 _2917_ (.Y(_1010_),
    .B1(net731),
    .B2(\GUScpu0.PC0[3] ),
    .A2(net734),
    .A1(\uart0.q[3] ));
 sg13g2_a22oi_1 _2918_ (.Y(_1011_),
    .B1(net727),
    .B2(net3),
    .A2(_0979_),
    .A1(\GUScpu0.cv[0][0] ));
 sg13g2_nand2b_1 _2919_ (.Y(_1012_),
    .B(_0902_),
    .A_N(\uart0.urxbuffer[8] ));
 sg13g2_nand3_1 _2920_ (.B(_1011_),
    .C(_1012_),
    .A(_1010_),
    .Y(_1013_));
 sg13g2_a21oi_1 _2921_ (.A1(\irqen[3] ),
    .A2(_0978_),
    .Y(_1014_),
    .B1(_1013_));
 sg13g2_a21oi_1 _2922_ (.A1(_0941_),
    .A2(_0964_),
    .Y(_1015_),
    .B1(_0967_));
 sg13g2_nor2b_1 _2923_ (.A(\xdi[3] ),
    .B_N(net725),
    .Y(_1016_));
 sg13g2_a221oi_1 _2924_ (.B2(net720),
    .C1(_1016_),
    .B1(_1015_),
    .A1(net722),
    .Y(\GUScpu0.cdi[3] ),
    .A2(_1014_));
 sg13g2_nand2_1 _2925_ (.Y(_1017_),
    .A(\uart0.q[4] ),
    .B(net734));
 sg13g2_a22oi_1 _2926_ (.Y(_1018_),
    .B1(net727),
    .B2(net5),
    .A2(net731),
    .A1(\GUScpu0.PC0[4] ));
 sg13g2_a22oi_1 _2927_ (.Y(_1019_),
    .B1(_0978_),
    .B2(\irqen[4] ),
    .A2(_0902_),
    .A1(pwmirq));
 sg13g2_nand3_1 _2928_ (.B(_1018_),
    .C(_1019_),
    .A(_1017_),
    .Y(_1020_));
 sg13g2_a22oi_1 _2929_ (.Y(_1021_),
    .B1(_1020_),
    .B2(net723),
    .A2(_0999_),
    .A1(net720));
 sg13g2_a22oi_1 _2930_ (.Y(_1022_),
    .B1(net721),
    .B2(_0968_),
    .A2(_0829_),
    .A1(\xdi[4] ));
 sg13g2_nand2_2 _2931_ (.Y(\GUScpu0.cdi[4] ),
    .A(_1021_),
    .B(_1022_));
 sg13g2_a21oi_1 _2932_ (.A1(net732),
    .A2(_0963_),
    .Y(_1023_),
    .B1(_1002_));
 sg13g2_o21ai_1 _2933_ (.B1(net726),
    .Y(_1024_),
    .A1(_0901_),
    .A2(_0973_));
 sg13g2_and3_1 _2934_ (.X(_1025_),
    .A(net720),
    .B(_1023_),
    .C(_1024_));
 sg13g2_a22oi_1 _2935_ (.Y(_1026_),
    .B1(_0902_),
    .B2(sdty),
    .A2(net734),
    .A1(\uart0.q[5] ));
 sg13g2_a22oi_1 _2936_ (.Y(_1027_),
    .B1(net727),
    .B2(net6),
    .A2(net731),
    .A1(\GUScpu0.PC0[5] ));
 sg13g2_and2_1 _2937_ (.A(_1026_),
    .B(_1027_),
    .X(_1028_));
 sg13g2_a221oi_1 _2938_ (.B2(_1028_),
    .C1(_1025_),
    .B1(net723),
    .A1(_1502_),
    .Y(\GUScpu0.cdi[5] ),
    .A2(net725));
 sg13g2_nor4_1 _2939_ (.A(\uart0.q[7] ),
    .B(\uart0.q[6] ),
    .C(\uart0.q[5] ),
    .D(\uart0.q[4] ),
    .Y(_1029_));
 sg13g2_nor2_1 _2940_ (.A(\uart0.q[3] ),
    .B(\uart0.q[2] ),
    .Y(_1030_));
 sg13g2_nand4_1 _2941_ (.B(\uart0.q[0] ),
    .C(_1029_),
    .A(\uart0.q[1] ),
    .Y(_1031_),
    .D(_1030_));
 sg13g2_nor3_1 _2942_ (.A(_0077_),
    .B(_0903_),
    .C(_1031_),
    .Y(_1032_));
 sg13g2_a21o_1 _2943_ (.A2(net727),
    .A1(net7),
    .B1(_1032_),
    .X(_1033_));
 sg13g2_a221oi_1 _2944_ (.B2(\GUScpu0.PC0[6] ),
    .C1(_1033_),
    .B1(net731),
    .A1(\uart0.q[6] ),
    .Y(_1034_),
    .A2(net733));
 sg13g2_or2_1 _2945_ (.X(_1035_),
    .B(_0997_),
    .A(_0942_));
 sg13g2_nor2_1 _2946_ (.A(_0941_),
    .B(_1035_),
    .Y(_1036_));
 sg13g2_nor3_1 _2947_ (.A(_0851_),
    .B(_0964_),
    .C(_0974_),
    .Y(_1037_));
 sg13g2_a221oi_1 _2948_ (.B2(net726),
    .C1(_1037_),
    .B1(_1036_),
    .A1(net729),
    .Y(_1038_),
    .A2(_0970_));
 sg13g2_nor2b_1 _2949_ (.A(\xdi[6] ),
    .B_N(net724),
    .Y(_1039_));
 sg13g2_a221oi_1 _2950_ (.B2(net720),
    .C1(_1039_),
    .B1(_1038_),
    .A1(net723),
    .Y(\GUScpu0.cdi[6] ),
    .A2(_1034_));
 sg13g2_nand2_1 _2951_ (.Y(_1040_),
    .A(net8),
    .B(net727));
 sg13g2_a22oi_1 _2952_ (.Y(_1041_),
    .B1(net732),
    .B2(\GUScpu0.PC0[7] ),
    .A2(net734),
    .A1(\uart0.q[7] ));
 sg13g2_nand2_1 _2953_ (.Y(_1042_),
    .A(_1040_),
    .B(_1041_));
 sg13g2_nand2_1 _2954_ (.Y(_1043_),
    .A(\xdi[7] ),
    .B(net724));
 sg13g2_o21ai_1 _2955_ (.B1(net726),
    .Y(_1044_),
    .A1(_0901_),
    .A2(net728));
 sg13g2_nand2_1 _2956_ (.Y(_1045_),
    .A(_1023_),
    .B(_1044_));
 sg13g2_a22oi_1 _2957_ (.Y(_1046_),
    .B1(_1045_),
    .B2(net721),
    .A2(_1042_),
    .A1(net723));
 sg13g2_nand2_2 _2958_ (.Y(\GUScpu0.cdi[7] ),
    .A(_1043_),
    .B(_1046_));
 sg13g2_nor4_2 _2959_ (.A(net735),
    .B(_0954_),
    .C(net729),
    .Y(_1047_),
    .D(_0974_));
 sg13g2_a221oi_1 _2960_ (.B2(_1035_),
    .C1(_1047_),
    .B1(_0963_),
    .A1(_0859_),
    .Y(_1048_),
    .A2(net729));
 sg13g2_nand2b_1 _2961_ (.Y(_1049_),
    .B(net720),
    .A_N(_1048_));
 sg13g2_a22oi_1 _2962_ (.Y(_1050_),
    .B1(_0945_),
    .B2(\GUScpu0.PC0[8] ),
    .A2(net725),
    .A1(net9));
 sg13g2_nand2_2 _2963_ (.Y(\GUScpu0.cdi[8] ),
    .A(_1049_),
    .B(_1050_));
 sg13g2_nand2_1 _2964_ (.Y(_1051_),
    .A(net735),
    .B(_0860_));
 sg13g2_nand3_1 _2965_ (.B(_0976_),
    .C(_1051_),
    .A(net726),
    .Y(_1052_));
 sg13g2_o21ai_1 _2966_ (.B1(_1052_),
    .Y(_1053_),
    .A1(_0964_),
    .A2(_1036_));
 sg13g2_nand2_1 _2967_ (.Y(_1054_),
    .A(net10),
    .B(net724));
 sg13g2_a22oi_1 _2968_ (.Y(_1055_),
    .B1(net720),
    .B2(_1053_),
    .A2(_0945_),
    .A1(\GUScpu0.PC0[9] ));
 sg13g2_nand2_2 _2969_ (.Y(\GUScpu0.cdi[9] ),
    .A(_1054_),
    .B(_1055_));
 sg13g2_and3_1 _2970_ (.X(_1056_),
    .A(_0858_),
    .B(_0963_),
    .C(_0995_));
 sg13g2_o21ai_1 _2971_ (.B1(net720),
    .Y(_1057_),
    .A1(_1047_),
    .A2(_1056_));
 sg13g2_a22oi_1 _2972_ (.Y(_1058_),
    .B1(_0945_),
    .B2(\GUScpu0.PC0[10] ),
    .A2(net724),
    .A1(net11));
 sg13g2_nand2_2 _2973_ (.Y(\GUScpu0.cdi[10] ),
    .A(_1057_),
    .B(_1058_));
 sg13g2_nor2_1 _2974_ (.A(_0942_),
    .B(_0964_),
    .Y(_1059_));
 sg13g2_nand2_1 _2975_ (.Y(_1060_),
    .A(_0970_),
    .B(_1003_));
 sg13g2_a22oi_1 _2976_ (.Y(_1061_),
    .B1(_1059_),
    .B2(_0844_),
    .A2(_0975_),
    .A1(net729));
 sg13g2_nand3_1 _2977_ (.B(_1060_),
    .C(_1061_),
    .A(net720),
    .Y(_1062_));
 sg13g2_a22oi_1 _2978_ (.Y(_1063_),
    .B1(_0945_),
    .B2(\GUScpu0.PC0[11] ),
    .A2(net724),
    .A1(net12));
 sg13g2_nand2_2 _2979_ (.Y(\GUScpu0.cdi[11] ),
    .A(_1062_),
    .B(_1063_));
 sg13g2_nand2_1 _2980_ (.Y(_1064_),
    .A(net13),
    .B(net724));
 sg13g2_a22oi_1 _2981_ (.Y(_1065_),
    .B1(_1059_),
    .B2(_0845_),
    .A2(_0977_),
    .A1(_0964_));
 sg13g2_a22oi_1 _2982_ (.Y(_1066_),
    .B1(_0947_),
    .B2(_1065_),
    .A2(_0945_),
    .A1(\GUScpu0.PC0[12] ));
 sg13g2_nand2_2 _2983_ (.Y(\GUScpu0.cdi[12] ),
    .A(_1064_),
    .B(_1066_));
 sg13g2_nand2_1 _2984_ (.Y(_1067_),
    .A(\GUScpu0.PC0[13] ),
    .B(net732));
 sg13g2_nor3_1 _2985_ (.A(_0942_),
    .B(_0964_),
    .C(_0995_),
    .Y(_1068_));
 sg13g2_nand2_1 _2986_ (.Y(_1069_),
    .A(_0903_),
    .B(_1051_));
 sg13g2_a221oi_1 _2987_ (.B2(net726),
    .C1(_1068_),
    .B1(_1069_),
    .A1(net729),
    .Y(_1070_),
    .A2(_0975_));
 sg13g2_and2_1 _2988_ (.A(net721),
    .B(_1070_),
    .X(_1071_));
 sg13g2_a221oi_1 _2989_ (.B2(_1067_),
    .C1(_1071_),
    .B1(net723),
    .A1(_1503_),
    .Y(\GUScpu0.cdi[13] ),
    .A2(net725));
 sg13g2_nand2_1 _2990_ (.Y(_1072_),
    .A(\GUScpu0.PC0[14] ),
    .B(net732));
 sg13g2_o21ai_1 _2991_ (.B1(net726),
    .Y(_1073_),
    .A1(net736),
    .A2(_0995_));
 sg13g2_nand2_1 _2992_ (.Y(_1074_),
    .A(_0985_),
    .B(_1073_));
 sg13g2_nor4_1 _2993_ (.A(net725),
    .B(_0835_),
    .C(_1068_),
    .D(_1074_),
    .Y(_1075_));
 sg13g2_a221oi_1 _2994_ (.B2(_1072_),
    .C1(_1075_),
    .B1(net723),
    .A1(_1504_),
    .Y(\GUScpu0.cdi[14] ),
    .A2(net725));
 sg13g2_nor3_2 _2995_ (.A(_0078_),
    .B(_0917_),
    .C(_0918_),
    .Y(_1076_));
 sg13g2_nor2_1 _2996_ (.A(\pwmc[0] ),
    .B(_1076_),
    .Y(_0000_));
 sg13g2_and2_1 _2997_ (.A(\pwmc[0] ),
    .B(\pwmc[1] ),
    .X(_1077_));
 sg13g2_nor3_1 _2998_ (.A(_0899_),
    .B(_1076_),
    .C(_1077_),
    .Y(_0001_));
 sg13g2_xnor2_1 _2999_ (.Y(_1078_),
    .A(\pwmc[2] ),
    .B(_1077_));
 sg13g2_nor2_1 _3000_ (.A(_1076_),
    .B(_1078_),
    .Y(_0002_));
 sg13g2_a21oi_1 _3001_ (.A1(\pwmc[2] ),
    .A2(_1077_),
    .Y(_1079_),
    .B1(\pwmc[3] ));
 sg13g2_and3_1 _3002_ (.X(_1080_),
    .A(\pwmc[3] ),
    .B(\pwmc[2] ),
    .C(_1077_));
 sg13g2_nor3_1 _3003_ (.A(_1076_),
    .B(_1079_),
    .C(_1080_),
    .Y(_0003_));
 sg13g2_nor2_1 _3004_ (.A(\pwmc[4] ),
    .B(_1080_),
    .Y(_1081_));
 sg13g2_and2_1 _3005_ (.A(\pwmc[4] ),
    .B(_1080_),
    .X(_1082_));
 sg13g2_nor3_1 _3006_ (.A(_1076_),
    .B(_1081_),
    .C(_1082_),
    .Y(_0004_));
 sg13g2_xnor2_1 _3007_ (.Y(_1083_),
    .A(\pwmc[5] ),
    .B(_1082_));
 sg13g2_nor2_1 _3008_ (.A(_1076_),
    .B(_1083_),
    .Y(_0005_));
 sg13g2_a21oi_1 _3009_ (.A1(\pwmc[5] ),
    .A2(_1082_),
    .Y(_1084_),
    .B1(\pwmc[6] ));
 sg13g2_nand3_1 _3010_ (.B(\pwmc[6] ),
    .C(_1082_),
    .A(\pwmc[5] ),
    .Y(_1085_));
 sg13g2_nand2b_1 _3011_ (.Y(_1086_),
    .B(_1085_),
    .A_N(_1084_));
 sg13g2_nor2_1 _3012_ (.A(_1076_),
    .B(_1086_),
    .Y(_0006_));
 sg13g2_a21oi_1 _3013_ (.A1(_0078_),
    .A2(_1085_),
    .Y(_0007_),
    .B1(_1076_));
 sg13g2_nor2_1 _3014_ (.A(_0083_),
    .B(_1521_),
    .Y(_1087_));
 sg13g2_nor4_1 _3015_ (.A(_0083_),
    .B(_0101_),
    .C(_1521_),
    .D(_1530_),
    .Y(_1088_));
 sg13g2_nand2_1 _3016_ (.Y(_1089_),
    .A(net884),
    .B(_1088_));
 sg13g2_nand3_1 _3017_ (.B(\GUScpu0.IR[0] ),
    .C(_1088_),
    .A(\GUScpu0.IR[1] ),
    .Y(_1090_));
 sg13g2_nor4_1 _3018_ (.A(_0083_),
    .B(_0101_),
    .C(_1521_),
    .D(_1530_),
    .Y(_1091_));
 sg13g2_nand2_1 _3019_ (.Y(_1092_),
    .A(net871),
    .B(_1090_));
 sg13g2_mux2_1 _3020_ (.A0(\GUScpu0.flag0[0] ),
    .A1(\GUScpu0.zn[1][1] ),
    .S(net870),
    .X(_1093_));
 sg13g2_mux2_1 _3021_ (.A0(_1093_),
    .A1(_0472_),
    .S(\GUScpu0.IR[13] ),
    .X(_1094_));
 sg13g2_a21oi_1 _3022_ (.A1(_0079_),
    .A2(_1094_),
    .Y(_1095_),
    .B1(\GUScpu0.IR[14] ));
 sg13g2_o21ai_1 _3023_ (.B1(_1095_),
    .Y(_1096_),
    .A1(_0079_),
    .A2(_1094_));
 sg13g2_nor2_1 _3024_ (.A(_1472_),
    .B(\GUScpu0.zn[1][0] ),
    .Y(_1097_));
 sg13g2_nor2_1 _3025_ (.A(net870),
    .B(\GUScpu0.flag0[2] ),
    .Y(_1098_));
 sg13g2_nor3_1 _3026_ (.A(\GUScpu0.IR[13] ),
    .B(_1097_),
    .C(_1098_),
    .Y(_1099_));
 sg13g2_nor2_1 _3027_ (.A(_1472_),
    .B(\GUScpu0.cv[1][0] ),
    .Y(_1100_));
 sg13g2_o21ai_1 _3028_ (.B1(\GUScpu0.IR[13] ),
    .Y(_1101_),
    .A1(net870),
    .A2(\GUScpu0.cv[0][0] ));
 sg13g2_o21ai_1 _3029_ (.B1(_0079_),
    .Y(_1102_),
    .A1(_1100_),
    .A2(_1101_));
 sg13g2_nand2b_1 _3030_ (.Y(_1103_),
    .B(_1102_),
    .A_N(_1099_));
 sg13g2_nand2_1 _3031_ (.Y(_1104_),
    .A(_0079_),
    .B(_1099_));
 sg13g2_nand3_1 _3032_ (.B(_1103_),
    .C(_1104_),
    .A(\GUScpu0.IR[14] ),
    .Y(_1105_));
 sg13g2_nand4_1 _3033_ (.B(\GUScpu0.opval ),
    .C(_1096_),
    .A(\GUScpu0.IR[15] ),
    .Y(_1106_),
    .D(_1105_));
 sg13g2_nand3_1 _3034_ (.B(_1089_),
    .C(_1106_),
    .A(net848),
    .Y(_1107_));
 sg13g2_nor2b_1 _3035_ (.A(net871),
    .B_N(\GUScpu0.irqq0 ),
    .Y(_1108_));
 sg13g2_and2_1 _3036_ (.A(_1529_),
    .B(_1091_),
    .X(_1109_));
 sg13g2_nor2b_1 _3037_ (.A(_1109_),
    .B_N(_1108_),
    .Y(_1110_));
 sg13g2_nor2_1 _3038_ (.A(net857),
    .B(_1110_),
    .Y(_1111_));
 sg13g2_nor2_1 _3039_ (.A(_0843_),
    .B(_1110_),
    .Y(_1112_));
 sg13g2_nand2_1 _3040_ (.Y(_1113_),
    .A(_0428_),
    .B(_1112_));
 sg13g2_nand3_1 _3041_ (.B(_0489_),
    .C(_1112_),
    .A(_0428_),
    .Y(_1114_));
 sg13g2_nand2_1 _3042_ (.Y(_1115_),
    .A(_0488_),
    .B(_1113_));
 sg13g2_a21oi_1 _3043_ (.A1(_1114_),
    .A2(_1115_),
    .Y(_1116_),
    .B1(net759));
 sg13g2_and2_2 _3044_ (.A(_0101_),
    .B(_1087_),
    .X(_1117_));
 sg13g2_nand2_1 _3045_ (.Y(_1118_),
    .A(_0134_),
    .B(_1117_));
 sg13g2_nand2b_1 _3046_ (.Y(_1119_),
    .B(_1527_),
    .A_N(_1117_));
 sg13g2_nand2_1 _3047_ (.Y(_1120_),
    .A(_1118_),
    .B(_1119_));
 sg13g2_and2_1 _3048_ (.A(_1118_),
    .B(_1119_),
    .X(_1121_));
 sg13g2_nand2_1 _3049_ (.Y(_1122_),
    .A(\GUScpu0.IR[1] ),
    .B(_1117_));
 sg13g2_nand2_1 _3050_ (.Y(_1123_),
    .A(\GUScpu0.IR[5] ),
    .B(_1117_));
 sg13g2_and2_1 _3051_ (.A(_1480_),
    .B(_1117_),
    .X(_1124_));
 sg13g2_nand2_1 _3052_ (.Y(_1125_),
    .A(_1480_),
    .B(_1117_));
 sg13g2_nand2_1 _3053_ (.Y(_1126_),
    .A(_0791_),
    .B(net809));
 sg13g2_o21ai_1 _3054_ (.B1(_1126_),
    .Y(_1127_),
    .A1(_0770_),
    .A2(net808));
 sg13g2_nand2_1 _3055_ (.Y(_1128_),
    .A(_0848_),
    .B(net809));
 sg13g2_o21ai_1 _3056_ (.B1(_1128_),
    .Y(_1129_),
    .A1(_0803_),
    .A2(net808));
 sg13g2_mux2_1 _3057_ (.A0(_1127_),
    .A1(_1129_),
    .S(net813),
    .X(_1130_));
 sg13g2_nand2_1 _3058_ (.Y(_1131_),
    .A(net814),
    .B(_1130_));
 sg13g2_nand2_1 _3059_ (.Y(_1132_),
    .A(_1527_),
    .B(_0841_));
 sg13g2_a221oi_1 _3060_ (.B2(_0760_),
    .C1(_0765_),
    .B1(net758),
    .A1(_1522_),
    .Y(_1133_),
    .A2(_1524_));
 sg13g2_o21ai_1 _3061_ (.B1(_1526_),
    .Y(_1134_),
    .A1(net884),
    .A2(_0472_));
 sg13g2_o21ai_1 _3062_ (.B1(_1132_),
    .Y(_1135_),
    .A1(_1133_),
    .A2(_1134_));
 sg13g2_mux4_1 _3063_ (.S0(net810),
    .A0(_0797_),
    .A1(_1135_),
    .A2(_0958_),
    .A3(_0782_),
    .S1(net813),
    .X(_1136_));
 sg13g2_o21ai_1 _3064_ (.B1(_1131_),
    .Y(_1137_),
    .A1(net818),
    .A2(_1136_));
 sg13g2_nand2_1 _3065_ (.Y(_1138_),
    .A(net771),
    .B(_1137_));
 sg13g2_or2_1 _3066_ (.X(_1139_),
    .B(_1109_),
    .A(_1516_));
 sg13g2_nor2_1 _3067_ (.A(_0834_),
    .B(net810),
    .Y(_1140_));
 sg13g2_a21oi_1 _3068_ (.A1(_0816_),
    .A2(net810),
    .Y(_1141_),
    .B1(_1140_));
 sg13g2_nand2_1 _3069_ (.Y(_1142_),
    .A(_0808_),
    .B(net808));
 sg13g2_o21ai_1 _3070_ (.B1(_1142_),
    .Y(_1143_),
    .A1(_0855_),
    .A2(net808));
 sg13g2_mux2_1 _3071_ (.A0(_1143_),
    .A1(_1141_),
    .S(net812),
    .X(_1144_));
 sg13g2_nor2_1 _3072_ (.A(net815),
    .B(_1144_),
    .Y(_1145_));
 sg13g2_mux2_1 _3073_ (.A0(_0777_),
    .A1(_0953_),
    .S(net808),
    .X(_1146_));
 sg13g2_mux2_1 _3074_ (.A0(_0766_),
    .A1(_0823_),
    .S(net808),
    .X(_1147_));
 sg13g2_mux2_1 _3075_ (.A0(_1147_),
    .A1(_1146_),
    .S(net812),
    .X(_1148_));
 sg13g2_a21oi_1 _3076_ (.A1(net815),
    .A2(_1148_),
    .Y(_1149_),
    .B1(_1145_));
 sg13g2_a21oi_1 _3077_ (.A1(net769),
    .A2(_1149_),
    .Y(_1150_),
    .B1(net803));
 sg13g2_a22oi_1 _3078_ (.Y(_1151_),
    .B1(_1150_),
    .B2(_1138_),
    .A2(net807),
    .A1(\GUScpu0.cdi[2] ));
 sg13g2_a21oi_1 _3079_ (.A1(net759),
    .A2(_1151_),
    .Y(_1152_),
    .B1(_1116_));
 sg13g2_a22oi_1 _3080_ (.Y(_1153_),
    .B1(_0863_),
    .B2(\irqen[1] ),
    .A2(\irqen[3] ),
    .A1(pwmirq));
 sg13g2_a21oi_2 _3081_ (.B1(_1153_),
    .Y(_1154_),
    .A2(\irqen[0] ),
    .A1(\uart0.rxvalid ));
 sg13g2_mux2_1 _3082_ (.A0(_1152_),
    .A1(_1154_),
    .S(net819),
    .X(_0008_));
 sg13g2_nand2b_1 _3083_ (.Y(_1155_),
    .B(_0511_),
    .A_N(_1114_));
 sg13g2_xnor2_1 _3084_ (.Y(_1156_),
    .A(_0511_),
    .B(_1114_));
 sg13g2_nand2_1 _3085_ (.Y(_1157_),
    .A(_0848_),
    .B(net811));
 sg13g2_o21ai_1 _3086_ (.B1(_1157_),
    .Y(_1158_),
    .A1(_0803_),
    .A2(net810));
 sg13g2_mux2_1 _3087_ (.A0(_1158_),
    .A1(_1127_),
    .S(net813),
    .X(_1159_));
 sg13g2_nor2_1 _3088_ (.A(net814),
    .B(_1159_),
    .Y(_1160_));
 sg13g2_a21oi_1 _3089_ (.A1(net818),
    .A2(_1136_),
    .Y(_1161_),
    .B1(_1160_));
 sg13g2_nand2_1 _3090_ (.Y(_1162_),
    .A(net769),
    .B(_1161_));
 sg13g2_a21oi_1 _3091_ (.A1(net771),
    .A2(_1149_),
    .Y(_1163_),
    .B1(net802));
 sg13g2_a22oi_1 _3092_ (.Y(_1164_),
    .B1(_1162_),
    .B2(_1163_),
    .A2(net807),
    .A1(\GUScpu0.cdi[3] ));
 sg13g2_nand2_1 _3093_ (.Y(_1165_),
    .A(net759),
    .B(_1164_));
 sg13g2_o21ai_1 _3094_ (.B1(_1165_),
    .Y(_1166_),
    .A1(net759),
    .A2(_1156_));
 sg13g2_a22oi_1 _3095_ (.Y(_1167_),
    .B1(\irqen[1] ),
    .B2(_0863_),
    .A2(\irqen[0] ),
    .A1(\uart0.rxvalid ));
 sg13g2_nand4_1 _3096_ (.B(\irqen[3] ),
    .C(net819),
    .A(pwmirq),
    .Y(_1168_),
    .D(_1167_));
 sg13g2_o21ai_1 _3097_ (.B1(_1168_),
    .Y(_0009_),
    .A1(net821),
    .A2(_1166_));
 sg13g2_nor2b_1 _3098_ (.A(_1155_),
    .B_N(_0596_),
    .Y(_1169_));
 sg13g2_xnor2_1 _3099_ (.Y(_1170_),
    .A(_0596_),
    .B(_1155_));
 sg13g2_nand2_1 _3100_ (.Y(_1171_),
    .A(net771),
    .B(_1161_));
 sg13g2_mux2_1 _3101_ (.A0(_0777_),
    .A1(_0953_),
    .S(net810),
    .X(_1172_));
 sg13g2_mux2_1 _3102_ (.A0(_1172_),
    .A1(_1147_),
    .S(net812),
    .X(_1173_));
 sg13g2_nand2_1 _3103_ (.Y(_1174_),
    .A(net815),
    .B(_1144_));
 sg13g2_o21ai_1 _3104_ (.B1(_1174_),
    .Y(_1175_),
    .A1(net815),
    .A2(_1173_));
 sg13g2_a21oi_1 _3105_ (.A1(net769),
    .A2(_1175_),
    .Y(_1176_),
    .B1(net802));
 sg13g2_a22oi_1 _3106_ (.Y(_1177_),
    .B1(_1171_),
    .B2(_1176_),
    .A2(net807),
    .A1(\GUScpu0.cdi[4] ));
 sg13g2_nand2_1 _3107_ (.Y(_1178_),
    .A(net759),
    .B(_1177_));
 sg13g2_o21ai_1 _3108_ (.B1(_1178_),
    .Y(_1179_),
    .A1(net759),
    .A2(_1170_));
 sg13g2_o21ai_1 _3109_ (.B1(_1167_),
    .Y(_1180_),
    .A1(_1462_),
    .A2(_1501_));
 sg13g2_nand2b_1 _3110_ (.Y(_1181_),
    .B(net819),
    .A_N(_1180_));
 sg13g2_o21ai_1 _3111_ (.B1(_1181_),
    .Y(_0010_),
    .A1(net819),
    .A2(_1179_));
 sg13g2_nor2_1 _3112_ (.A(\uart0.txdiv[0] ),
    .B(_0881_),
    .Y(_0019_));
 sg13g2_nor2_1 _3113_ (.A(\uart0.txdiv[0] ),
    .B(\uart0.txdiv[1] ),
    .Y(_1182_));
 sg13g2_nor3_1 _3114_ (.A(_0871_),
    .B(net718),
    .C(_1182_),
    .Y(_0020_));
 sg13g2_and2_1 _3115_ (.A(\uart0.txdiv[2] ),
    .B(_0871_),
    .X(_1183_));
 sg13g2_o21ai_1 _3116_ (.B1(_0880_),
    .Y(_1184_),
    .A1(\uart0.txdiv[2] ),
    .A2(_0871_));
 sg13g2_nor2_1 _3117_ (.A(_1183_),
    .B(_1184_),
    .Y(_0021_));
 sg13g2_and2_1 _3118_ (.A(\uart0.txdiv[3] ),
    .B(_1183_),
    .X(_1185_));
 sg13g2_nor2_1 _3119_ (.A(\uart0.txdiv[3] ),
    .B(_1183_),
    .Y(_1186_));
 sg13g2_nor3_1 _3120_ (.A(_0881_),
    .B(_1185_),
    .C(_1186_),
    .Y(_0022_));
 sg13g2_or2_1 _3121_ (.X(_1187_),
    .B(_1185_),
    .A(\uart0.txdiv[4] ));
 sg13g2_nand2_1 _3122_ (.Y(_1188_),
    .A(\uart0.txdiv[4] ),
    .B(_1185_));
 sg13g2_and3_1 _3123_ (.X(_0023_),
    .A(_0880_),
    .B(_1187_),
    .C(_1188_));
 sg13g2_xor2_1 _3124_ (.B(_1188_),
    .A(\uart0.txdiv[5] ),
    .X(_1189_));
 sg13g2_nor2_1 _3125_ (.A(_0881_),
    .B(_1189_),
    .Y(_0024_));
 sg13g2_xnor2_1 _3126_ (.Y(_1190_),
    .A(\uart0.rxreg[0] ),
    .B(\uart0.rxreg[1] ));
 sg13g2_nand2_1 _3127_ (.Y(_1191_),
    .A(\uart0.rxdiv[1] ),
    .B(\uart0.rxdiv[0] ));
 sg13g2_nor2_1 _3128_ (.A(\uart0.rxdiv[2] ),
    .B(\uart0.rxdiv[3] ),
    .Y(_1192_));
 sg13g2_nand3_1 _3129_ (.B(\uart0.rxdiv[4] ),
    .C(_1192_),
    .A(\uart0.rxdiv[5] ),
    .Y(_1193_));
 sg13g2_o21ai_1 _3130_ (.B1(_1190_),
    .Y(_1194_),
    .A1(_1191_),
    .A2(_1193_));
 sg13g2_inv_1 _3131_ (.Y(_1195_),
    .A(_1194_));
 sg13g2_nor2_1 _3132_ (.A(\uart0.rxdiv[0] ),
    .B(_1194_),
    .Y(_0013_));
 sg13g2_or2_1 _3133_ (.X(_1196_),
    .B(\uart0.rxdiv[0] ),
    .A(\uart0.rxdiv[1] ));
 sg13g2_and3_1 _3134_ (.X(_0014_),
    .A(_1190_),
    .B(_1191_),
    .C(_1196_));
 sg13g2_a21oi_1 _3135_ (.A1(\uart0.rxdiv[1] ),
    .A2(\uart0.rxdiv[0] ),
    .Y(_1197_),
    .B1(\uart0.rxdiv[2] ));
 sg13g2_and3_1 _3136_ (.X(_1198_),
    .A(\uart0.rxdiv[1] ),
    .B(\uart0.rxdiv[0] ),
    .C(\uart0.rxdiv[2] ));
 sg13g2_nor3_1 _3137_ (.A(_1194_),
    .B(_1197_),
    .C(_1198_),
    .Y(_0015_));
 sg13g2_nor2_1 _3138_ (.A(\uart0.rxdiv[3] ),
    .B(_1198_),
    .Y(_1199_));
 sg13g2_and2_1 _3139_ (.A(\uart0.rxdiv[3] ),
    .B(_1198_),
    .X(_1200_));
 sg13g2_nor3_1 _3140_ (.A(_1194_),
    .B(_1199_),
    .C(_1200_),
    .Y(_0016_));
 sg13g2_nand2_1 _3141_ (.Y(_1201_),
    .A(\uart0.rxdiv[4] ),
    .B(_1200_));
 sg13g2_o21ai_1 _3142_ (.B1(_1195_),
    .Y(_1202_),
    .A1(\uart0.rxdiv[4] ),
    .A2(_1200_));
 sg13g2_nor2b_1 _3143_ (.A(_1202_),
    .B_N(_1201_),
    .Y(_0017_));
 sg13g2_xor2_1 _3144_ (.B(_1201_),
    .A(\uart0.rxdiv[5] ),
    .X(_1203_));
 sg13g2_nor2_1 _3145_ (.A(_1194_),
    .B(_1203_),
    .Y(_0018_));
 sg13g2_nand2b_1 _3146_ (.Y(_1204_),
    .B(net923),
    .A_N(_0799_));
 sg13g2_o21ai_1 _3147_ (.B1(\ckd[0] ),
    .Y(_1205_),
    .A1(_1468_),
    .A2(_0659_));
 sg13g2_nor2_1 _3148_ (.A(net935),
    .B(_1468_),
    .Y(_1206_));
 sg13g2_nand2b_2 _3149_ (.Y(_1207_),
    .B(net231),
    .A_N(net935));
 sg13g2_o21ai_1 _3150_ (.B1(_1205_),
    .Y(_1208_),
    .A1(_0463_),
    .A2(net922));
 sg13g2_nand2_2 _3151_ (.Y(_1209_),
    .A(net935),
    .B(\ckd[1] ));
 sg13g2_a22oi_1 _3152_ (.Y(uio_out[0]),
    .B1(_1204_),
    .B2(_1208_),
    .A2(xlal),
    .A1(_0845_));
 sg13g2_nor2_1 _3153_ (.A(_0439_),
    .B(net922),
    .Y(_1210_));
 sg13g2_a221oi_1 _3154_ (.B2(_0858_),
    .C1(_1210_),
    .B1(xlal),
    .A1(_0810_),
    .Y(_1211_),
    .A2(net923));
 sg13g2_o21ai_1 _3155_ (.B1(_1211_),
    .Y(uio_out[1]),
    .A1(_0686_),
    .A2(_1209_));
 sg13g2_nor2_1 _3156_ (.A(_0497_),
    .B(net922),
    .Y(_1212_));
 sg13g2_a221oi_1 _3157_ (.B2(_0852_),
    .C1(_1212_),
    .B1(xlal),
    .A1(_0804_),
    .Y(_1213_),
    .A2(net923));
 sg13g2_o21ai_1 _3158_ (.B1(_1213_),
    .Y(uio_out[2]),
    .A1(_0741_),
    .A2(_1209_));
 sg13g2_o21ai_1 _3159_ (.B1(net923),
    .Y(_1214_),
    .A1(_0778_),
    .A2(_0779_));
 sg13g2_o21ai_1 _3160_ (.B1(net935),
    .Y(_1215_),
    .A1(_1468_),
    .A2(_0714_));
 sg13g2_o21ai_1 _3161_ (.B1(_1215_),
    .Y(_1216_),
    .A1(_0521_),
    .A2(net922));
 sg13g2_a22oi_1 _3162_ (.Y(uio_out[3]),
    .B1(_1214_),
    .B2(_1216_),
    .A2(xlal),
    .A1(_0955_));
 sg13g2_nor2_1 _3163_ (.A(_0605_),
    .B(net922),
    .Y(_1217_));
 sg13g2_a221oi_1 _3164_ (.B2(xlal),
    .C1(_1217_),
    .B1(net730),
    .A1(_0783_),
    .Y(_1218_),
    .A2(net923));
 sg13g2_o21ai_1 _3165_ (.B1(_1218_),
    .Y(uio_out[4]),
    .A1(_1703_),
    .A2(_1209_));
 sg13g2_mux4_1 _3166_ (.S0(net935),
    .A0(_0836_),
    .A1(_0818_),
    .A2(_0624_),
    .A3(_1678_),
    .S1(\ckd[1] ),
    .X(_1219_));
 sg13g2_inv_2 _3167_ (.Y(uio_out[5]),
    .A(_1219_));
 sg13g2_nor2b_1 _3168_ (.A(_0772_),
    .B_N(net923),
    .Y(_1220_));
 sg13g2_a221oi_1 _3169_ (.B2(_0551_),
    .C1(_1220_),
    .B1(net885),
    .A1(_0794_),
    .Y(_1221_),
    .A2(xlal));
 sg13g2_o21ai_1 _3170_ (.B1(_1221_),
    .Y(uio_out[6]),
    .A1(_1651_),
    .A2(_1209_));
 sg13g2_a221oi_1 _3171_ (.B2(net885),
    .C1(net923),
    .B1(_0579_),
    .A1(net935),
    .Y(_1222_),
    .A2(_1623_));
 sg13g2_a21oi_1 _3172_ (.A1(_0767_),
    .A2(net923),
    .Y(_1223_),
    .B1(_1222_));
 sg13g2_a21oi_2 _3173_ (.B1(_1223_),
    .Y(uio_out[7]),
    .A2(xlal),
    .A1(_0826_));
 sg13g2_or2_2 _3174_ (.X(xoeb),
    .B(net867),
    .A(net934));
 sg13g2_nor4_1 _3175_ (.A(net866),
    .B(net760),
    .C(_1108_),
    .D(net807),
    .Y(\GUScpu0.opvali ));
 sg13g2_nand3b_1 _3176_ (.B(net867),
    .C(\ckd[1] ),
    .Y(xweb),
    .A_N(clknet_1_0__leaf_clk));
 sg13g2_or2_2 _3177_ (.X(\GUScpu0.clk ),
    .B(_0867_),
    .A(net927));
 sg13g2_nand2b_1 _3178_ (.Y(_1224_),
    .B(_1090_),
    .A_N(_0082_));
 sg13g2_a21oi_1 _3179_ (.A1(_1472_),
    .A2(\irqen[4] ),
    .Y(_1225_),
    .B1(_1180_));
 sg13g2_o21ai_1 _3180_ (.B1(_1224_),
    .Y(_0011_),
    .A1(_0867_),
    .A2(_1225_));
 sg13g2_nor2b_1 _3181_ (.A(_0082_),
    .B_N(_0011_),
    .Y(_0012_));
 sg13g2_nand2b_1 _3182_ (.Y(_0171_),
    .B(net922),
    .A_N(xlah));
 sg13g2_nor3_2 _3183_ (.A(_1528_),
    .B(_1586_),
    .C(_1590_),
    .Y(_1226_));
 sg13g2_nor2_1 _3184_ (.A(_1515_),
    .B(_1593_),
    .Y(_1227_));
 sg13g2_a21oi_2 _3185_ (.B1(_0083_),
    .Y(_1228_),
    .A2(_1227_),
    .A1(_1226_));
 sg13g2_nand2_1 _3186_ (.Y(_1229_),
    .A(net870),
    .B(_1228_));
 sg13g2_mux4_1 _3187_ (.S0(net813),
    .A0(_0782_),
    .A1(_0797_),
    .A2(_0958_),
    .A3(_1135_),
    .S1(net809),
    .X(_1230_));
 sg13g2_nor2_1 _3188_ (.A(net816),
    .B(_1130_),
    .Y(_1231_));
 sg13g2_a21oi_1 _3189_ (.A1(net816),
    .A2(_1230_),
    .Y(_1232_),
    .B1(_1231_));
 sg13g2_nand2_1 _3190_ (.Y(_1233_),
    .A(net769),
    .B(_1232_));
 sg13g2_nand2_1 _3191_ (.Y(_1234_),
    .A(_0808_),
    .B(net810));
 sg13g2_o21ai_1 _3192_ (.B1(_1234_),
    .Y(_1235_),
    .A1(_0855_),
    .A2(net810));
 sg13g2_mux2_1 _3193_ (.A0(_1141_),
    .A1(_1235_),
    .S(net812),
    .X(_1236_));
 sg13g2_nor2_1 _3194_ (.A(net814),
    .B(_1236_),
    .Y(_1237_));
 sg13g2_mux2_1 _3195_ (.A0(_0766_),
    .A1(_0823_),
    .S(net810),
    .X(_1238_));
 sg13g2_mux2_1 _3196_ (.A0(_1146_),
    .A1(_1238_),
    .S(net812),
    .X(_1239_));
 sg13g2_a21oi_1 _3197_ (.A1(net814),
    .A2(_1239_),
    .Y(_1240_),
    .B1(_1237_));
 sg13g2_a21oi_1 _3198_ (.A1(net772),
    .A2(_1240_),
    .Y(_1241_),
    .B1(net802));
 sg13g2_a22oi_1 _3199_ (.Y(_1242_),
    .B1(_1233_),
    .B2(_1241_),
    .A2(net803),
    .A1(\GUScpu0.cdi[15] ));
 sg13g2_inv_1 _3200_ (.Y(_1243_),
    .A(_1242_));
 sg13g2_nand2_1 _3201_ (.Y(_1244_),
    .A(\GUScpu0.zn[1][0] ),
    .B(_1229_));
 sg13g2_o21ai_1 _3202_ (.B1(_1244_),
    .Y(_0192_),
    .A1(_1229_),
    .A2(_1242_));
 sg13g2_nand2_1 _3203_ (.Y(_1245_),
    .A(_0791_),
    .B(net811));
 sg13g2_o21ai_1 _3204_ (.B1(_1245_),
    .Y(_1246_),
    .A1(_0770_),
    .A2(net811));
 sg13g2_mux2_1 _3205_ (.A0(_1129_),
    .A1(_1246_),
    .S(net813),
    .X(_1247_));
 sg13g2_nand2_1 _3206_ (.Y(_1248_),
    .A(net817),
    .B(_1247_));
 sg13g2_o21ai_1 _3207_ (.B1(_1248_),
    .Y(_1249_),
    .A1(net817),
    .A2(_1230_));
 sg13g2_nand2_1 _3208_ (.Y(_1250_),
    .A(net770),
    .B(_1249_));
 sg13g2_nor2_1 _3209_ (.A(_0834_),
    .B(net808),
    .Y(_1251_));
 sg13g2_a21oi_1 _3210_ (.A1(_0816_),
    .A2(net808),
    .Y(_1252_),
    .B1(_1251_));
 sg13g2_mux2_1 _3211_ (.A0(_1235_),
    .A1(_1252_),
    .S(net812),
    .X(_1253_));
 sg13g2_nand2_1 _3212_ (.Y(_1254_),
    .A(net814),
    .B(_1253_));
 sg13g2_o21ai_1 _3213_ (.B1(_1254_),
    .Y(_1255_),
    .A1(net816),
    .A2(_1239_));
 sg13g2_a21oi_1 _3214_ (.A1(net772),
    .A2(_1255_),
    .Y(_1256_),
    .B1(net804));
 sg13g2_a22oi_1 _3215_ (.Y(_1257_),
    .B1(_1250_),
    .B2(_1256_),
    .A2(net805),
    .A1(\GUScpu0.cdi[13] ));
 sg13g2_mux4_1 _3216_ (.S0(net813),
    .A0(_0797_),
    .A1(_0958_),
    .A2(_1135_),
    .A3(_0782_),
    .S1(net809),
    .X(_1258_));
 sg13g2_nor2_1 _3217_ (.A(net817),
    .B(_1247_),
    .Y(_1259_));
 sg13g2_a21oi_1 _3218_ (.A1(net817),
    .A2(_1258_),
    .Y(_1260_),
    .B1(_1259_));
 sg13g2_nand2_1 _3219_ (.Y(_1261_),
    .A(net772),
    .B(_1260_));
 sg13g2_a21oi_1 _3220_ (.A1(net770),
    .A2(_1255_),
    .Y(_1262_),
    .B1(net804));
 sg13g2_a22oi_1 _3221_ (.Y(_1263_),
    .B1(_1261_),
    .B2(_1262_),
    .A2(net805),
    .A1(\GUScpu0.cdi[12] ));
 sg13g2_mux4_1 _3222_ (.S0(net813),
    .A0(_0782_),
    .A1(_0797_),
    .A2(_0958_),
    .A3(_1135_),
    .S1(net811),
    .X(_1264_));
 sg13g2_mux2_1 _3223_ (.A0(_1246_),
    .A1(_1158_),
    .S(net813),
    .X(_1265_));
 sg13g2_nor2_1 _3224_ (.A(net817),
    .B(_1265_),
    .Y(_1266_));
 sg13g2_a21oi_1 _3225_ (.A1(net816),
    .A2(_1264_),
    .Y(_1267_),
    .B1(_1266_));
 sg13g2_nand2_1 _3226_ (.Y(_1268_),
    .A(net772),
    .B(_1267_));
 sg13g2_mux2_1 _3227_ (.A0(_1238_),
    .A1(_1172_),
    .S(net812),
    .X(_1269_));
 sg13g2_mux2_1 _3228_ (.A0(_1252_),
    .A1(_1143_),
    .S(net812),
    .X(_1270_));
 sg13g2_nand2_1 _3229_ (.Y(_1271_),
    .A(net814),
    .B(_1270_));
 sg13g2_o21ai_1 _3230_ (.B1(_1271_),
    .Y(_1272_),
    .A1(net816),
    .A2(_1269_));
 sg13g2_a21oi_1 _3231_ (.A1(net770),
    .A2(_1272_),
    .Y(_1273_),
    .B1(net804));
 sg13g2_a22oi_1 _3232_ (.Y(_1274_),
    .B1(_1268_),
    .B2(_1273_),
    .A2(net804),
    .A1(\GUScpu0.cdi[8] ));
 sg13g2_nand2_1 _3233_ (.Y(_1275_),
    .A(net772),
    .B(_1249_));
 sg13g2_a21oi_1 _3234_ (.A1(net770),
    .A2(_1240_),
    .Y(_1276_),
    .B1(net804));
 sg13g2_a22oi_1 _3235_ (.Y(_1277_),
    .B1(_1275_),
    .B2(_1276_),
    .A2(net804),
    .A1(\GUScpu0.cdi[14] ));
 sg13g2_nand4_1 _3236_ (.B(_1263_),
    .C(_1274_),
    .A(_1257_),
    .Y(_1278_),
    .D(_1277_));
 sg13g2_nand4_1 _3237_ (.B(_1164_),
    .C(_1177_),
    .A(_1151_),
    .Y(_1279_),
    .D(_1242_));
 sg13g2_nand2_1 _3238_ (.Y(_1280_),
    .A(net771),
    .B(_1232_));
 sg13g2_nand2_1 _3239_ (.Y(_1281_),
    .A(net815),
    .B(_1236_));
 sg13g2_o21ai_1 _3240_ (.B1(_1281_),
    .Y(_1282_),
    .A1(net815),
    .A2(_1148_));
 sg13g2_a21oi_1 _3241_ (.A1(net769),
    .A2(_1282_),
    .Y(_1283_),
    .B1(net802));
 sg13g2_a22oi_1 _3242_ (.Y(_1284_),
    .B1(_1280_),
    .B2(_1283_),
    .A2(net803),
    .A1(\GUScpu0.cdi[0] ));
 sg13g2_nand2_1 _3243_ (.Y(_1285_),
    .A(net816),
    .B(_1159_));
 sg13g2_o21ai_1 _3244_ (.B1(_1285_),
    .Y(_1286_),
    .A1(net814),
    .A2(_1264_));
 sg13g2_nand2_1 _3245_ (.Y(_1287_),
    .A(net769),
    .B(_1286_));
 sg13g2_a21oi_1 _3246_ (.A1(net771),
    .A2(_1175_),
    .Y(_1288_),
    .B1(net802));
 sg13g2_a22oi_1 _3247_ (.Y(_1289_),
    .B1(_1287_),
    .B2(_1288_),
    .A2(net802),
    .A1(\GUScpu0.cdi[5] ));
 sg13g2_nand2_1 _3248_ (.Y(_1290_),
    .A(net771),
    .B(_1286_));
 sg13g2_nor2_1 _3249_ (.A(net814),
    .B(_1270_),
    .Y(_1291_));
 sg13g2_a21oi_1 _3250_ (.A1(net815),
    .A2(_1173_),
    .Y(_1292_),
    .B1(_1291_));
 sg13g2_a21oi_1 _3251_ (.A1(net769),
    .A2(_1292_),
    .Y(_1293_),
    .B1(net802));
 sg13g2_a22oi_1 _3252_ (.Y(_1294_),
    .B1(_1290_),
    .B2(_1293_),
    .A2(net803),
    .A1(\GUScpu0.cdi[6] ));
 sg13g2_nand2_1 _3253_ (.Y(_1295_),
    .A(net769),
    .B(_1137_));
 sg13g2_a21oi_1 _3254_ (.A1(net771),
    .A2(_1282_),
    .Y(_1296_),
    .B1(net803));
 sg13g2_a22oi_1 _3255_ (.Y(_1297_),
    .B1(_1295_),
    .B2(_1296_),
    .A2(net803),
    .A1(\GUScpu0.cdi[1] ));
 sg13g2_nand4_1 _3256_ (.B(_1289_),
    .C(_1294_),
    .A(_1284_),
    .Y(_1298_),
    .D(_1297_));
 sg13g2_nand2_1 _3257_ (.Y(_1299_),
    .A(net817),
    .B(_1265_));
 sg13g2_o21ai_1 _3258_ (.B1(_1299_),
    .Y(_1300_),
    .A1(net817),
    .A2(_1258_));
 sg13g2_nand2_1 _3259_ (.Y(_1301_),
    .A(net772),
    .B(_1300_));
 sg13g2_nor2_1 _3260_ (.A(net816),
    .B(_1253_),
    .Y(_1302_));
 sg13g2_a21oi_1 _3261_ (.A1(net816),
    .A2(_1269_),
    .Y(_1303_),
    .B1(_1302_));
 sg13g2_a21oi_1 _3262_ (.A1(net770),
    .A2(_1303_),
    .Y(_1304_),
    .B1(net805));
 sg13g2_a22oi_1 _3263_ (.Y(_1305_),
    .B1(_1301_),
    .B2(_1304_),
    .A2(net805),
    .A1(\GUScpu0.cdi[10] ));
 sg13g2_nand2_1 _3264_ (.Y(_1306_),
    .A(net770),
    .B(_1267_));
 sg13g2_a21oi_1 _3265_ (.A1(net771),
    .A2(_1292_),
    .Y(_1307_),
    .B1(net802));
 sg13g2_a22oi_1 _3266_ (.Y(_1308_),
    .B1(_1306_),
    .B2(_1307_),
    .A2(net804),
    .A1(\GUScpu0.cdi[7] ));
 sg13g2_nand2_1 _3267_ (.Y(_1309_),
    .A(net770),
    .B(_1260_));
 sg13g2_a21oi_1 _3268_ (.A1(net772),
    .A2(_1303_),
    .Y(_1310_),
    .B1(net805));
 sg13g2_a22oi_1 _3269_ (.Y(_1311_),
    .B1(_1309_),
    .B2(_1310_),
    .A2(net805),
    .A1(\GUScpu0.cdi[11] ));
 sg13g2_nand2_1 _3270_ (.Y(_1312_),
    .A(net770),
    .B(_1300_));
 sg13g2_a21oi_1 _3271_ (.A1(net772),
    .A2(_1272_),
    .Y(_1313_),
    .B1(net804));
 sg13g2_a22oi_1 _3272_ (.Y(_1314_),
    .B1(_1312_),
    .B2(_1313_),
    .A2(net805),
    .A1(\GUScpu0.cdi[9] ));
 sg13g2_nand4_1 _3273_ (.B(_1308_),
    .C(_1311_),
    .A(_1305_),
    .Y(_1315_),
    .D(_1314_));
 sg13g2_nor4_2 _3274_ (.A(_1278_),
    .B(_1279_),
    .C(_1298_),
    .Y(_1316_),
    .D(_1315_));
 sg13g2_mux2_1 _3275_ (.A0(_1316_),
    .A1(\GUScpu0.zn[1][1] ),
    .S(_1229_),
    .X(_0193_));
 sg13g2_mux2_1 _3276_ (.A0(net225),
    .A1(net9),
    .S(_1206_),
    .X(_0194_));
 sg13g2_nor2_1 _3277_ (.A(net10),
    .B(net922),
    .Y(_1317_));
 sg13g2_a21oi_1 _3278_ (.A1(_1499_),
    .A2(_1207_),
    .Y(_0195_),
    .B1(_1317_));
 sg13g2_nor2_1 _3279_ (.A(net11),
    .B(_1207_),
    .Y(_1318_));
 sg13g2_a21oi_1 _3280_ (.A1(_1500_),
    .A2(net922),
    .Y(_0196_),
    .B1(_1318_));
 sg13g2_mux2_1 _3281_ (.A0(net224),
    .A1(net12),
    .S(net885),
    .X(_0197_));
 sg13g2_mux2_1 _3282_ (.A0(net223),
    .A1(net13),
    .S(net885),
    .X(_0198_));
 sg13g2_nor2_1 _3283_ (.A(net228),
    .B(net885),
    .Y(_1319_));
 sg13g2_a21oi_1 _3284_ (.A1(_1503_),
    .A2(net885),
    .Y(_0199_),
    .B1(_1319_));
 sg13g2_nor2_1 _3285_ (.A(net229),
    .B(net885),
    .Y(_1320_));
 sg13g2_a21oi_1 _3286_ (.A1(_1504_),
    .A2(net885),
    .Y(_0200_),
    .B1(_1320_));
 sg13g2_mux2_1 _3287_ (.A0(net16),
    .A1(net227),
    .S(_1207_),
    .X(_0201_));
 sg13g2_nand3b_1 _3288_ (.B(_1558_),
    .C(_1592_),
    .Y(_1321_),
    .A_N(_1515_));
 sg13g2_nor3_1 _3289_ (.A(_1532_),
    .B(_1545_),
    .C(_1321_),
    .Y(_1322_));
 sg13g2_a21oi_2 _3290_ (.B1(_1471_),
    .Y(_1323_),
    .A2(_1322_),
    .A1(_1226_));
 sg13g2_and2_1 _3291_ (.A(\GUScpu0.IR[8] ),
    .B(_1323_),
    .X(_1324_));
 sg13g2_nand2_1 _3292_ (.Y(_1325_),
    .A(_0089_),
    .B(net849));
 sg13g2_nor2_1 _3293_ (.A(net883),
    .B(_1325_),
    .Y(_1326_));
 sg13g2_nand2_1 _3294_ (.Y(_1327_),
    .A(_1324_),
    .B(_1326_));
 sg13g2_nor2_1 _3295_ (.A(net848),
    .B(_0454_),
    .Y(_1328_));
 sg13g2_a21oi_2 _3296_ (.B1(_1328_),
    .Y(_1329_),
    .A2(_1284_),
    .A1(net848));
 sg13g2_mux2_1 _3297_ (.A0(_1329_),
    .A1(\GUScpu0.regs[5][0] ),
    .S(net747),
    .X(_0202_));
 sg13g2_nor2_1 _3298_ (.A(net848),
    .B(_0428_),
    .Y(_1330_));
 sg13g2_a21oi_2 _3299_ (.B1(_1330_),
    .Y(_1331_),
    .A2(_1297_),
    .A1(net848));
 sg13g2_mux2_1 _3300_ (.A0(_1331_),
    .A1(\GUScpu0.regs[5][1] ),
    .S(net747),
    .X(_0203_));
 sg13g2_nor2_1 _3301_ (.A(net850),
    .B(_0489_),
    .Y(_1332_));
 sg13g2_a21oi_2 _3302_ (.B1(_1332_),
    .Y(_1333_),
    .A2(_1151_),
    .A1(net850));
 sg13g2_mux2_1 _3303_ (.A0(_1333_),
    .A1(\GUScpu0.regs[5][2] ),
    .S(net747),
    .X(_0204_));
 sg13g2_nor2_1 _3304_ (.A(net848),
    .B(_0511_),
    .Y(_1334_));
 sg13g2_a21oi_2 _3305_ (.B1(_1334_),
    .Y(_1335_),
    .A2(_1164_),
    .A1(net848));
 sg13g2_mux2_1 _3306_ (.A0(_1335_),
    .A1(\GUScpu0.regs[5][3] ),
    .S(net747),
    .X(_0205_));
 sg13g2_nor2_1 _3307_ (.A(net849),
    .B(_0596_),
    .Y(_1336_));
 sg13g2_a21oi_2 _3308_ (.B1(_1336_),
    .Y(_1337_),
    .A2(_1177_),
    .A1(net849));
 sg13g2_mux2_1 _3309_ (.A0(_1337_),
    .A1(\GUScpu0.regs[5][4] ),
    .S(net747),
    .X(_0206_));
 sg13g2_nor2_1 _3310_ (.A(net851),
    .B(_0615_),
    .Y(_1338_));
 sg13g2_a21oi_2 _3311_ (.B1(_1338_),
    .Y(_1339_),
    .A2(_1289_),
    .A1(net851));
 sg13g2_mux2_1 _3312_ (.A0(_1339_),
    .A1(\GUScpu0.regs[5][5] ),
    .S(net747),
    .X(_0207_));
 sg13g2_nor2_1 _3313_ (.A(net850),
    .B(_0542_),
    .Y(_1340_));
 sg13g2_a21oi_2 _3314_ (.B1(_1340_),
    .Y(_1341_),
    .A2(_1294_),
    .A1(net850));
 sg13g2_mux2_1 _3315_ (.A0(_1341_),
    .A1(\GUScpu0.regs[5][6] ),
    .S(net748),
    .X(_0208_));
 sg13g2_nor2_1 _3316_ (.A(net851),
    .B(_0569_),
    .Y(_1342_));
 sg13g2_a21oi_2 _3317_ (.B1(_1342_),
    .Y(_1343_),
    .A2(_1308_),
    .A1(net851));
 sg13g2_mux2_1 _3318_ (.A0(_1343_),
    .A1(\GUScpu0.regs[5][7] ),
    .S(net747),
    .X(_0209_));
 sg13g2_nor2_1 _3319_ (.A(net854),
    .B(_0648_),
    .Y(_1344_));
 sg13g2_a21oi_2 _3320_ (.B1(_1344_),
    .Y(_1345_),
    .A2(_1274_),
    .A1(net854));
 sg13g2_mux2_1 _3321_ (.A0(_1345_),
    .A1(\GUScpu0.regs[5][8] ),
    .S(net748),
    .X(_0210_));
 sg13g2_nor2_1 _3322_ (.A(net852),
    .B(_0677_),
    .Y(_1346_));
 sg13g2_a21oi_2 _3323_ (.B1(_1346_),
    .Y(_1347_),
    .A2(_1314_),
    .A1(net852));
 sg13g2_mux2_1 _3324_ (.A0(_1347_),
    .A1(\GUScpu0.regs[5][9] ),
    .S(net748),
    .X(_0211_));
 sg13g2_nor2_1 _3325_ (.A(net853),
    .B(_0731_),
    .Y(_1348_));
 sg13g2_a21oi_2 _3326_ (.B1(_1348_),
    .Y(_1349_),
    .A2(_1305_),
    .A1(net853));
 sg13g2_mux2_1 _3327_ (.A0(_1349_),
    .A1(\GUScpu0.regs[5][10] ),
    .S(net748),
    .X(_0212_));
 sg13g2_nor2_1 _3328_ (.A(net852),
    .B(_0705_),
    .Y(_1350_));
 sg13g2_a21oi_2 _3329_ (.B1(_1350_),
    .Y(_1351_),
    .A2(_1311_),
    .A1(net854));
 sg13g2_mux2_1 _3330_ (.A0(_1351_),
    .A1(\GUScpu0.regs[5][11] ),
    .S(net748),
    .X(_0213_));
 sg13g2_nor2_1 _3331_ (.A(net853),
    .B(_1693_),
    .Y(_1352_));
 sg13g2_a21oi_2 _3332_ (.B1(_1352_),
    .Y(_1353_),
    .A2(_1263_),
    .A1(net852));
 sg13g2_mux2_1 _3333_ (.A0(_1353_),
    .A1(\GUScpu0.regs[5][12] ),
    .S(net748),
    .X(_0214_));
 sg13g2_nor2_1 _3334_ (.A(net852),
    .B(_1668_),
    .Y(_1354_));
 sg13g2_a21oi_2 _3335_ (.B1(_1354_),
    .Y(_1355_),
    .A2(_1257_),
    .A1(net852));
 sg13g2_mux2_1 _3336_ (.A0(_1355_),
    .A1(\GUScpu0.regs[5][13] ),
    .S(net748),
    .X(_0215_));
 sg13g2_nor2_1 _3337_ (.A(net852),
    .B(_1642_),
    .Y(_1356_));
 sg13g2_a21oi_2 _3338_ (.B1(_1356_),
    .Y(_1357_),
    .A2(_1277_),
    .A1(net852));
 sg13g2_mux2_1 _3339_ (.A0(_1357_),
    .A1(\GUScpu0.regs[5][14] ),
    .S(net748),
    .X(_0216_));
 sg13g2_nor2_1 _3340_ (.A(_1597_),
    .B(net850),
    .Y(_1358_));
 sg13g2_a21oi_2 _3341_ (.B1(_1358_),
    .Y(_1359_),
    .A2(_1242_),
    .A1(net850));
 sg13g2_mux2_1 _3342_ (.A0(_1359_),
    .A1(\GUScpu0.regs[5][15] ),
    .S(net747),
    .X(_0217_));
 sg13g2_nand2_1 _3343_ (.Y(_1360_),
    .A(net883),
    .B(net849));
 sg13g2_o21ai_1 _3344_ (.B1(net849),
    .Y(_1361_),
    .A1(_0089_),
    .A2(net883));
 sg13g2_nand2_1 _3345_ (.Y(_1362_),
    .A(\GUScpu0.IR[8] ),
    .B(net849));
 sg13g2_nand3_1 _3346_ (.B(_1361_),
    .C(_1362_),
    .A(_1323_),
    .Y(_1363_));
 sg13g2_mux2_1 _3347_ (.A0(_1329_),
    .A1(\GUScpu0.regs[6][0] ),
    .S(net751),
    .X(_0218_));
 sg13g2_mux2_1 _3348_ (.A0(_1331_),
    .A1(\GUScpu0.regs[6][1] ),
    .S(net751),
    .X(_0219_));
 sg13g2_mux2_1 _3349_ (.A0(_1333_),
    .A1(\GUScpu0.regs[6][2] ),
    .S(net751),
    .X(_0220_));
 sg13g2_mux2_1 _3350_ (.A0(_1335_),
    .A1(\GUScpu0.regs[6][3] ),
    .S(net751),
    .X(_0221_));
 sg13g2_mux2_1 _3351_ (.A0(_1337_),
    .A1(\GUScpu0.regs[6][4] ),
    .S(net751),
    .X(_0222_));
 sg13g2_mux2_1 _3352_ (.A0(_1339_),
    .A1(\GUScpu0.regs[6][5] ),
    .S(net751),
    .X(_0223_));
 sg13g2_mux2_1 _3353_ (.A0(_1341_),
    .A1(\GUScpu0.regs[6][6] ),
    .S(net751),
    .X(_0224_));
 sg13g2_mux2_1 _3354_ (.A0(_1343_),
    .A1(\GUScpu0.regs[6][7] ),
    .S(net751),
    .X(_0225_));
 sg13g2_mux2_1 _3355_ (.A0(_1345_),
    .A1(\GUScpu0.regs[6][8] ),
    .S(_1363_),
    .X(_0226_));
 sg13g2_mux2_1 _3356_ (.A0(_1347_),
    .A1(\GUScpu0.regs[6][9] ),
    .S(net752),
    .X(_0227_));
 sg13g2_mux2_1 _3357_ (.A0(_1349_),
    .A1(\GUScpu0.regs[6][10] ),
    .S(net752),
    .X(_0228_));
 sg13g2_mux2_1 _3358_ (.A0(_1351_),
    .A1(\GUScpu0.regs[6][11] ),
    .S(net752),
    .X(_0229_));
 sg13g2_mux2_1 _3359_ (.A0(_1353_),
    .A1(\GUScpu0.regs[6][12] ),
    .S(net752),
    .X(_0230_));
 sg13g2_mux2_1 _3360_ (.A0(_1355_),
    .A1(\GUScpu0.regs[6][13] ),
    .S(net752),
    .X(_0231_));
 sg13g2_mux2_1 _3361_ (.A0(_1357_),
    .A1(\GUScpu0.regs[6][14] ),
    .S(net752),
    .X(_0232_));
 sg13g2_mux2_1 _3362_ (.A0(_1359_),
    .A1(\GUScpu0.regs[6][15] ),
    .S(net752),
    .X(_0233_));
 sg13g2_nand2b_2 _3363_ (.Y(_1364_),
    .B(_1323_),
    .A_N(\GUScpu0.IR[8] ));
 sg13g2_nor3_2 _3364_ (.A(_1475_),
    .B(_1360_),
    .C(_1364_),
    .Y(_1365_));
 sg13g2_mux2_1 _3365_ (.A0(\GUScpu0.regs[0][0] ),
    .A1(_1329_),
    .S(net745),
    .X(_0234_));
 sg13g2_mux2_1 _3366_ (.A0(\GUScpu0.regs[0][1] ),
    .A1(_1331_),
    .S(net745),
    .X(_0235_));
 sg13g2_mux2_1 _3367_ (.A0(\GUScpu0.regs[0][2] ),
    .A1(_1333_),
    .S(net745),
    .X(_0236_));
 sg13g2_mux2_1 _3368_ (.A0(\GUScpu0.regs[0][3] ),
    .A1(_1335_),
    .S(net745),
    .X(_0237_));
 sg13g2_mux2_1 _3369_ (.A0(\GUScpu0.regs[0][4] ),
    .A1(_1337_),
    .S(net745),
    .X(_0238_));
 sg13g2_mux2_1 _3370_ (.A0(\GUScpu0.regs[0][5] ),
    .A1(_1339_),
    .S(net745),
    .X(_0239_));
 sg13g2_mux2_1 _3371_ (.A0(\GUScpu0.regs[0][6] ),
    .A1(_1341_),
    .S(net745),
    .X(_0240_));
 sg13g2_mux2_1 _3372_ (.A0(\GUScpu0.regs[0][7] ),
    .A1(_1343_),
    .S(net746),
    .X(_0241_));
 sg13g2_mux2_1 _3373_ (.A0(\GUScpu0.regs[0][8] ),
    .A1(_1345_),
    .S(_1365_),
    .X(_0242_));
 sg13g2_mux2_1 _3374_ (.A0(\GUScpu0.regs[0][9] ),
    .A1(_1347_),
    .S(net746),
    .X(_0243_));
 sg13g2_mux2_1 _3375_ (.A0(\GUScpu0.regs[0][10] ),
    .A1(_1349_),
    .S(net746),
    .X(_0244_));
 sg13g2_mux2_1 _3376_ (.A0(\GUScpu0.regs[0][11] ),
    .A1(_1351_),
    .S(net746),
    .X(_0245_));
 sg13g2_mux2_1 _3377_ (.A0(\GUScpu0.regs[0][12] ),
    .A1(_1353_),
    .S(net746),
    .X(_0246_));
 sg13g2_mux2_1 _3378_ (.A0(\GUScpu0.regs[0][13] ),
    .A1(_1355_),
    .S(net746),
    .X(_0247_));
 sg13g2_mux2_1 _3379_ (.A0(\GUScpu0.regs[0][14] ),
    .A1(_1357_),
    .S(net746),
    .X(_0248_));
 sg13g2_mux2_1 _3380_ (.A0(\GUScpu0.regs[0][15] ),
    .A1(_1359_),
    .S(net745),
    .X(_0249_));
 sg13g2_a21oi_1 _3381_ (.A1(net880),
    .A2(_1538_),
    .Y(_1366_),
    .B1(_1600_));
 sg13g2_and4_1 _3382_ (.A(_1527_),
    .B(_1587_),
    .C(_0469_),
    .D(_1366_),
    .X(_1367_));
 sg13g2_a21oi_1 _3383_ (.A1(_1591_),
    .A2(_1367_),
    .Y(_1368_),
    .B1(_0083_));
 sg13g2_and2_1 _3384_ (.A(_0081_),
    .B(_1368_),
    .X(_1369_));
 sg13g2_nand3_1 _3385_ (.B(_1629_),
    .C(_0759_),
    .A(net758),
    .Y(_1370_));
 sg13g2_o21ai_1 _3386_ (.B1(_1370_),
    .Y(_1371_),
    .A1(_1627_),
    .A2(_0766_));
 sg13g2_mux2_1 _3387_ (.A0(\GUScpu0.cv[0][0] ),
    .A1(_1371_),
    .S(_1369_),
    .X(_0250_));
 sg13g2_nor2_1 _3388_ (.A(net755),
    .B(_1629_),
    .Y(_1372_));
 sg13g2_o21ai_1 _3389_ (.B1(_1372_),
    .Y(_1373_),
    .A1(_1626_),
    .A2(_0759_));
 sg13g2_o21ai_1 _3390_ (.B1(_1373_),
    .Y(_1374_),
    .A1(_1527_),
    .A2(_0464_));
 sg13g2_mux2_1 _3391_ (.A0(\GUScpu0.cv[0][1] ),
    .A1(_1374_),
    .S(_1369_),
    .X(_0251_));
 sg13g2_a22oi_1 _3392_ (.Y(_1375_),
    .B1(_0865_),
    .B2(sdty),
    .A2(_0864_),
    .A1(net733));
 sg13g2_inv_1 _3393_ (.Y(_0252_),
    .A(_1375_));
 sg13g2_nand2_1 _3394_ (.Y(_1376_),
    .A(_0864_),
    .B(net728));
 sg13g2_mux2_1 _3395_ (.A0(_0463_),
    .A1(gpo),
    .S(_1376_),
    .X(_0262_));
 sg13g2_mux2_1 _3396_ (.A0(\pwmhold[0] ),
    .A1(_0463_),
    .S(net716),
    .X(_0273_));
 sg13g2_nor2_1 _3397_ (.A(\pwmhold[1] ),
    .B(net717),
    .Y(_1377_));
 sg13g2_a21oi_1 _3398_ (.A1(_0439_),
    .A2(net717),
    .Y(_0274_),
    .B1(_1377_));
 sg13g2_nor2_1 _3399_ (.A(\pwmhold[2] ),
    .B(net716),
    .Y(_1378_));
 sg13g2_a21oi_1 _3400_ (.A1(_0497_),
    .A2(net716),
    .Y(_0275_),
    .B1(_1378_));
 sg13g2_nor2_1 _3401_ (.A(\pwmhold[3] ),
    .B(net716),
    .Y(_1379_));
 sg13g2_a21oi_1 _3402_ (.A1(_0520_),
    .A2(net716),
    .Y(_0276_),
    .B1(_1379_));
 sg13g2_nor2_1 _3403_ (.A(\pwmhold[4] ),
    .B(net717),
    .Y(_1380_));
 sg13g2_a21oi_1 _3404_ (.A1(_0605_),
    .A2(net716),
    .Y(_0277_),
    .B1(_1380_));
 sg13g2_nor2_1 _3405_ (.A(\pwmhold[5] ),
    .B(net716),
    .Y(_1381_));
 sg13g2_a21oi_1 _3406_ (.A1(_0624_),
    .A2(net716),
    .Y(_0278_),
    .B1(_1381_));
 sg13g2_mux2_1 _3407_ (.A0(\pwmhold[6] ),
    .A1(_0551_),
    .S(net717),
    .X(_0279_));
 sg13g2_nor2_1 _3408_ (.A(\pwmhold[7] ),
    .B(net717),
    .Y(_1382_));
 sg13g2_a21oi_1 _3409_ (.A1(_0579_),
    .A2(net717),
    .Y(_0280_),
    .B1(_1382_));
 sg13g2_nand2_1 _3410_ (.Y(_1383_),
    .A(_0864_),
    .B(_0997_));
 sg13g2_mux2_1 _3411_ (.A0(_0463_),
    .A1(\irqen[0] ),
    .S(net715),
    .X(_0281_));
 sg13g2_nand2_1 _3412_ (.Y(_1384_),
    .A(\irqen[1] ),
    .B(net715));
 sg13g2_o21ai_1 _3413_ (.B1(_1384_),
    .Y(_0282_),
    .A1(_0439_),
    .A2(net715));
 sg13g2_nand2_1 _3414_ (.Y(_1385_),
    .A(\irqen[2] ),
    .B(_1383_));
 sg13g2_o21ai_1 _3415_ (.B1(_1385_),
    .Y(_0283_),
    .A1(_0497_),
    .A2(net715));
 sg13g2_nor2_1 _3416_ (.A(_0521_),
    .B(net715),
    .Y(_1386_));
 sg13g2_a21oi_1 _3417_ (.A1(_1501_),
    .A2(net715),
    .Y(_0284_),
    .B1(_1386_));
 sg13g2_nand2_1 _3418_ (.Y(_1387_),
    .A(\irqen[4] ),
    .B(net715));
 sg13g2_o21ai_1 _3419_ (.B1(_1387_),
    .Y(_0285_),
    .A1(_0605_),
    .A2(net715));
 sg13g2_nand2_1 _3420_ (.Y(_1388_),
    .A(net760),
    .B(_1284_));
 sg13g2_xor2_1 _3421_ (.B(_1111_),
    .A(_0454_),
    .X(_1389_));
 sg13g2_o21ai_1 _3422_ (.B1(_1388_),
    .Y(_1390_),
    .A1(net760),
    .A2(_1389_));
 sg13g2_nor2_1 _3423_ (.A(net819),
    .B(_1390_),
    .Y(_0286_));
 sg13g2_o21ai_1 _3424_ (.B1(_0429_),
    .Y(_1391_),
    .A1(_0843_),
    .A2(_1110_));
 sg13g2_a21oi_1 _3425_ (.A1(_1113_),
    .A2(_1391_),
    .Y(_1392_),
    .B1(net760));
 sg13g2_a21oi_1 _3426_ (.A1(net760),
    .A2(_1297_),
    .Y(_1393_),
    .B1(_1392_));
 sg13g2_nor2b_1 _3427_ (.A(net819),
    .B_N(_1393_),
    .Y(_0287_));
 sg13g2_and2_1 _3428_ (.A(_0615_),
    .B(_1169_),
    .X(_1394_));
 sg13g2_xor2_1 _3429_ (.B(_1169_),
    .A(_0615_),
    .X(_1395_));
 sg13g2_nand2_1 _3430_ (.Y(_1396_),
    .A(net759),
    .B(_1289_));
 sg13g2_o21ai_1 _3431_ (.B1(_1396_),
    .Y(_1397_),
    .A1(net759),
    .A2(_1395_));
 sg13g2_nor2_1 _3432_ (.A(net819),
    .B(_1397_),
    .Y(_0288_));
 sg13g2_nand2_1 _3433_ (.Y(_1398_),
    .A(net760),
    .B(_1294_));
 sg13g2_xnor2_1 _3434_ (.Y(_1399_),
    .A(_0543_),
    .B(_1394_));
 sg13g2_o21ai_1 _3435_ (.B1(_1398_),
    .Y(_1400_),
    .A1(net760),
    .A2(_1399_));
 sg13g2_nor2_1 _3436_ (.A(net819),
    .B(_1400_),
    .Y(_0289_));
 sg13g2_nand2_1 _3437_ (.Y(_1401_),
    .A(net763),
    .B(_1308_));
 sg13g2_nand3_1 _3438_ (.B(_0569_),
    .C(_1394_),
    .A(_0542_),
    .Y(_1402_));
 sg13g2_a21o_1 _3439_ (.A2(_1394_),
    .A1(_0542_),
    .B1(_0569_),
    .X(_1403_));
 sg13g2_and2_1 _3440_ (.A(_1402_),
    .B(_1403_),
    .X(_1404_));
 sg13g2_o21ai_1 _3441_ (.B1(_1401_),
    .Y(_1405_),
    .A1(net763),
    .A2(_1404_));
 sg13g2_nor2_1 _3442_ (.A(net820),
    .B(_1405_),
    .Y(_0290_));
 sg13g2_nor2b_2 _3443_ (.A(_1402_),
    .B_N(_0648_),
    .Y(_1406_));
 sg13g2_xnor2_1 _3444_ (.Y(_1407_),
    .A(_0648_),
    .B(_1402_));
 sg13g2_nand2_1 _3445_ (.Y(_1408_),
    .A(net763),
    .B(_1274_));
 sg13g2_o21ai_1 _3446_ (.B1(_1408_),
    .Y(_1409_),
    .A1(net763),
    .A2(_1407_));
 sg13g2_nand2b_1 _3447_ (.Y(_0291_),
    .B(_1409_),
    .A_N(net820));
 sg13g2_nand2_1 _3448_ (.Y(_1410_),
    .A(net763),
    .B(_1314_));
 sg13g2_nand2_1 _3449_ (.Y(_1411_),
    .A(_0677_),
    .B(_1406_));
 sg13g2_xor2_1 _3450_ (.B(_1406_),
    .A(_0677_),
    .X(_1412_));
 sg13g2_o21ai_1 _3451_ (.B1(_1410_),
    .Y(_1413_),
    .A1(net762),
    .A2(_1412_));
 sg13g2_nor2_1 _3452_ (.A(net820),
    .B(_1413_),
    .Y(_0292_));
 sg13g2_nor3_2 _3453_ (.A(net883),
    .B(_1325_),
    .C(_1364_),
    .Y(_1414_));
 sg13g2_mux2_1 _3454_ (.A0(\GUScpu0.regs[4][0] ),
    .A1(_1329_),
    .S(net743),
    .X(_0293_));
 sg13g2_mux2_1 _3455_ (.A0(\GUScpu0.regs[4][1] ),
    .A1(_1331_),
    .S(net743),
    .X(_0294_));
 sg13g2_mux2_1 _3456_ (.A0(\GUScpu0.regs[4][2] ),
    .A1(_1333_),
    .S(net743),
    .X(_0295_));
 sg13g2_mux2_1 _3457_ (.A0(\GUScpu0.regs[4][3] ),
    .A1(_1335_),
    .S(net743),
    .X(_0296_));
 sg13g2_mux2_1 _3458_ (.A0(\GUScpu0.regs[4][4] ),
    .A1(_1337_),
    .S(net743),
    .X(_0297_));
 sg13g2_mux2_1 _3459_ (.A0(\GUScpu0.regs[4][5] ),
    .A1(_1339_),
    .S(net743),
    .X(_0298_));
 sg13g2_mux2_1 _3460_ (.A0(\GUScpu0.regs[4][6] ),
    .A1(_1341_),
    .S(net744),
    .X(_0299_));
 sg13g2_mux2_1 _3461_ (.A0(\GUScpu0.regs[4][7] ),
    .A1(_1343_),
    .S(net743),
    .X(_0300_));
 sg13g2_mux2_1 _3462_ (.A0(\GUScpu0.regs[4][8] ),
    .A1(_1345_),
    .S(net744),
    .X(_0301_));
 sg13g2_mux2_1 _3463_ (.A0(\GUScpu0.regs[4][9] ),
    .A1(_1347_),
    .S(net744),
    .X(_0302_));
 sg13g2_mux2_1 _3464_ (.A0(\GUScpu0.regs[4][10] ),
    .A1(_1349_),
    .S(net744),
    .X(_0303_));
 sg13g2_mux2_1 _3465_ (.A0(\GUScpu0.regs[4][11] ),
    .A1(_1351_),
    .S(net744),
    .X(_0304_));
 sg13g2_mux2_1 _3466_ (.A0(\GUScpu0.regs[4][12] ),
    .A1(_1353_),
    .S(net744),
    .X(_0305_));
 sg13g2_mux2_1 _3467_ (.A0(\GUScpu0.regs[4][13] ),
    .A1(_1355_),
    .S(net744),
    .X(_0306_));
 sg13g2_mux2_1 _3468_ (.A0(\GUScpu0.regs[4][14] ),
    .A1(_1357_),
    .S(net744),
    .X(_0307_));
 sg13g2_mux2_1 _3469_ (.A0(\GUScpu0.regs[4][15] ),
    .A1(_1359_),
    .S(net743),
    .X(_0308_));
 sg13g2_and2_1 _3470_ (.A(net870),
    .B(_1368_),
    .X(_1415_));
 sg13g2_mux2_1 _3471_ (.A0(\GUScpu0.cv[1][0] ),
    .A1(_1371_),
    .S(_1415_),
    .X(_0309_));
 sg13g2_mux2_1 _3472_ (.A0(\GUScpu0.cv[1][1] ),
    .A1(_1374_),
    .S(_1415_),
    .X(_0310_));
 sg13g2_nor2_1 _3473_ (.A(_0089_),
    .B(_1360_),
    .Y(_1416_));
 sg13g2_nand2_2 _3474_ (.Y(_1417_),
    .A(_1324_),
    .B(_1416_));
 sg13g2_mux2_1 _3475_ (.A0(_1329_),
    .A1(\GUScpu0.regs[3][0] ),
    .S(net741),
    .X(_0311_));
 sg13g2_mux2_1 _3476_ (.A0(_1331_),
    .A1(\GUScpu0.regs[3][1] ),
    .S(net741),
    .X(_0312_));
 sg13g2_mux2_1 _3477_ (.A0(_1333_),
    .A1(\GUScpu0.regs[3][2] ),
    .S(net741),
    .X(_0313_));
 sg13g2_mux2_1 _3478_ (.A0(_1335_),
    .A1(\GUScpu0.regs[3][3] ),
    .S(net741),
    .X(_0314_));
 sg13g2_mux2_1 _3479_ (.A0(_1337_),
    .A1(\GUScpu0.regs[3][4] ),
    .S(net741),
    .X(_0315_));
 sg13g2_mux2_1 _3480_ (.A0(_1339_),
    .A1(\GUScpu0.regs[3][5] ),
    .S(net741),
    .X(_0316_));
 sg13g2_mux2_1 _3481_ (.A0(_1341_),
    .A1(\GUScpu0.regs[3][6] ),
    .S(net741),
    .X(_0317_));
 sg13g2_mux2_1 _3482_ (.A0(_1343_),
    .A1(\GUScpu0.regs[3][7] ),
    .S(net742),
    .X(_0318_));
 sg13g2_mux2_1 _3483_ (.A0(_1345_),
    .A1(\GUScpu0.regs[3][8] ),
    .S(_1417_),
    .X(_0319_));
 sg13g2_mux2_1 _3484_ (.A0(_1347_),
    .A1(\GUScpu0.regs[3][9] ),
    .S(net742),
    .X(_0320_));
 sg13g2_mux2_1 _3485_ (.A0(_1349_),
    .A1(\GUScpu0.regs[3][10] ),
    .S(net742),
    .X(_0321_));
 sg13g2_mux2_1 _3486_ (.A0(_1351_),
    .A1(\GUScpu0.regs[3][11] ),
    .S(net742),
    .X(_0322_));
 sg13g2_mux2_1 _3487_ (.A0(_1353_),
    .A1(\GUScpu0.regs[3][12] ),
    .S(net742),
    .X(_0323_));
 sg13g2_mux2_1 _3488_ (.A0(_1355_),
    .A1(\GUScpu0.regs[3][13] ),
    .S(net742),
    .X(_0324_));
 sg13g2_mux2_1 _3489_ (.A0(_1357_),
    .A1(\GUScpu0.regs[3][14] ),
    .S(net742),
    .X(_0325_));
 sg13g2_mux2_1 _3490_ (.A0(_1359_),
    .A1(\GUScpu0.regs[3][15] ),
    .S(net741),
    .X(_0326_));
 sg13g2_nor2b_2 _3491_ (.A(_1364_),
    .B_N(_1416_),
    .Y(_1418_));
 sg13g2_mux2_1 _3492_ (.A0(\GUScpu0.regs[2][0] ),
    .A1(_1329_),
    .S(net739),
    .X(_0327_));
 sg13g2_mux2_1 _3493_ (.A0(\GUScpu0.regs[2][1] ),
    .A1(_1331_),
    .S(net740),
    .X(_0328_));
 sg13g2_mux2_1 _3494_ (.A0(\GUScpu0.regs[2][2] ),
    .A1(_1333_),
    .S(net739),
    .X(_0329_));
 sg13g2_mux2_1 _3495_ (.A0(\GUScpu0.regs[2][3] ),
    .A1(_1335_),
    .S(net739),
    .X(_0330_));
 sg13g2_mux2_1 _3496_ (.A0(\GUScpu0.regs[2][4] ),
    .A1(_1337_),
    .S(net739),
    .X(_0331_));
 sg13g2_mux2_1 _3497_ (.A0(\GUScpu0.regs[2][5] ),
    .A1(_1339_),
    .S(net739),
    .X(_0332_));
 sg13g2_mux2_1 _3498_ (.A0(\GUScpu0.regs[2][6] ),
    .A1(_1341_),
    .S(net739),
    .X(_0333_));
 sg13g2_mux2_1 _3499_ (.A0(\GUScpu0.regs[2][7] ),
    .A1(_1343_),
    .S(net739),
    .X(_0334_));
 sg13g2_mux2_1 _3500_ (.A0(\GUScpu0.regs[2][8] ),
    .A1(_1345_),
    .S(_1418_),
    .X(_0335_));
 sg13g2_mux2_1 _3501_ (.A0(\GUScpu0.regs[2][9] ),
    .A1(_1347_),
    .S(net740),
    .X(_0336_));
 sg13g2_mux2_1 _3502_ (.A0(\GUScpu0.regs[2][10] ),
    .A1(_1349_),
    .S(net740),
    .X(_0337_));
 sg13g2_mux2_1 _3503_ (.A0(\GUScpu0.regs[2][11] ),
    .A1(_1351_),
    .S(net740),
    .X(_0338_));
 sg13g2_mux2_1 _3504_ (.A0(\GUScpu0.regs[2][12] ),
    .A1(_1353_),
    .S(net740),
    .X(_0339_));
 sg13g2_mux2_1 _3505_ (.A0(\GUScpu0.regs[2][13] ),
    .A1(_1355_),
    .S(net740),
    .X(_0340_));
 sg13g2_mux2_1 _3506_ (.A0(\GUScpu0.regs[2][14] ),
    .A1(_1357_),
    .S(net740),
    .X(_0341_));
 sg13g2_mux2_1 _3507_ (.A0(\GUScpu0.regs[2][15] ),
    .A1(_1359_),
    .S(net739),
    .X(_0342_));
 sg13g2_nand3_1 _3508_ (.B(_0731_),
    .C(_1406_),
    .A(_0677_),
    .Y(_1419_));
 sg13g2_xnor2_1 _3509_ (.Y(_1420_),
    .A(_0731_),
    .B(_1411_));
 sg13g2_nand2_1 _3510_ (.Y(_1421_),
    .A(net761),
    .B(_1305_));
 sg13g2_o21ai_1 _3511_ (.B1(_1421_),
    .Y(_1422_),
    .A1(net761),
    .A2(_1420_));
 sg13g2_nor2_1 _3512_ (.A(net821),
    .B(_1422_),
    .Y(_0343_));
 sg13g2_nand2_1 _3513_ (.Y(_1423_),
    .A(net762),
    .B(_1311_));
 sg13g2_nor2b_1 _3514_ (.A(_1419_),
    .B_N(_0705_),
    .Y(_1424_));
 sg13g2_xnor2_1 _3515_ (.Y(_1425_),
    .A(_0705_),
    .B(_1419_));
 sg13g2_o21ai_1 _3516_ (.B1(_1423_),
    .Y(_1426_),
    .A1(net761),
    .A2(_1425_));
 sg13g2_nor2_1 _3517_ (.A(net820),
    .B(_1426_),
    .Y(_0344_));
 sg13g2_and2_1 _3518_ (.A(_1693_),
    .B(_1424_),
    .X(_1427_));
 sg13g2_xor2_1 _3519_ (.B(_1424_),
    .A(_1693_),
    .X(_1428_));
 sg13g2_nand2_1 _3520_ (.Y(_1429_),
    .A(net761),
    .B(_1263_));
 sg13g2_o21ai_1 _3521_ (.B1(_1429_),
    .Y(_1430_),
    .A1(net761),
    .A2(_1428_));
 sg13g2_nor2_1 _3522_ (.A(net820),
    .B(_1430_),
    .Y(_0345_));
 sg13g2_nand2_1 _3523_ (.Y(_1431_),
    .A(net762),
    .B(_1257_));
 sg13g2_nand2_1 _3524_ (.Y(_1432_),
    .A(_1668_),
    .B(_1427_));
 sg13g2_xor2_1 _3525_ (.B(_1427_),
    .A(_1668_),
    .X(_1433_));
 sg13g2_o21ai_1 _3526_ (.B1(_1431_),
    .Y(_1434_),
    .A1(net761),
    .A2(_1433_));
 sg13g2_nor2_1 _3527_ (.A(net820),
    .B(_1434_),
    .Y(_0346_));
 sg13g2_nand2_1 _3528_ (.Y(_1435_),
    .A(net761),
    .B(_1277_));
 sg13g2_nor2b_1 _3529_ (.A(_1432_),
    .B_N(_1642_),
    .Y(_1436_));
 sg13g2_xnor2_1 _3530_ (.Y(_1437_),
    .A(_1642_),
    .B(_1432_));
 sg13g2_o21ai_1 _3531_ (.B1(_1435_),
    .Y(_1438_),
    .A1(net761),
    .A2(_1437_));
 sg13g2_nor2_1 _3532_ (.A(net820),
    .B(_1438_),
    .Y(_0347_));
 sg13g2_xnor2_1 _3533_ (.Y(_1439_),
    .A(_1597_),
    .B(_1436_));
 sg13g2_nor2_1 _3534_ (.A(net763),
    .B(_1439_),
    .Y(_1440_));
 sg13g2_a21oi_1 _3535_ (.A1(net763),
    .A2(_1243_),
    .Y(_1441_),
    .B1(_1440_));
 sg13g2_nor2_1 _3536_ (.A(net820),
    .B(_1441_),
    .Y(_0348_));
 sg13g2_nand2_1 _3537_ (.Y(_1442_),
    .A(_0081_),
    .B(_1228_));
 sg13g2_nand2_1 _3538_ (.Y(_1443_),
    .A(\GUScpu0.flag0[2] ),
    .B(_1442_));
 sg13g2_o21ai_1 _3539_ (.B1(_1443_),
    .Y(_0349_),
    .A1(_1242_),
    .A2(_1442_));
 sg13g2_mux2_1 _3540_ (.A0(_1316_),
    .A1(\GUScpu0.flag0[0] ),
    .S(_1442_),
    .X(_0350_));
 sg13g2_nand4_1 _3541_ (.B(net849),
    .C(_1323_),
    .A(\GUScpu0.IR[8] ),
    .Y(_1444_),
    .D(_1361_));
 sg13g2_mux2_1 _3542_ (.A0(_1329_),
    .A1(\GUScpu0.regs[7][0] ),
    .S(net749),
    .X(_0351_));
 sg13g2_mux2_1 _3543_ (.A0(_1331_),
    .A1(\GUScpu0.regs[7][1] ),
    .S(net749),
    .X(_0352_));
 sg13g2_mux2_1 _3544_ (.A0(_1333_),
    .A1(\GUScpu0.regs[7][2] ),
    .S(net749),
    .X(_0353_));
 sg13g2_mux2_1 _3545_ (.A0(_1335_),
    .A1(\GUScpu0.regs[7][3] ),
    .S(net749),
    .X(_0354_));
 sg13g2_mux2_1 _3546_ (.A0(_1337_),
    .A1(\GUScpu0.regs[7][4] ),
    .S(net749),
    .X(_0355_));
 sg13g2_mux2_1 _3547_ (.A0(_1339_),
    .A1(\GUScpu0.regs[7][5] ),
    .S(net749),
    .X(_0356_));
 sg13g2_mux2_1 _3548_ (.A0(_1341_),
    .A1(\GUScpu0.regs[7][6] ),
    .S(net749),
    .X(_0357_));
 sg13g2_mux2_1 _3549_ (.A0(_1343_),
    .A1(\GUScpu0.regs[7][7] ),
    .S(net749),
    .X(_0358_));
 sg13g2_mux2_1 _3550_ (.A0(_1345_),
    .A1(\GUScpu0.regs[7][8] ),
    .S(_1444_),
    .X(_0359_));
 sg13g2_mux2_1 _3551_ (.A0(_1347_),
    .A1(\GUScpu0.regs[7][9] ),
    .S(net750),
    .X(_0360_));
 sg13g2_mux2_1 _3552_ (.A0(_1349_),
    .A1(\GUScpu0.regs[7][10] ),
    .S(net750),
    .X(_0361_));
 sg13g2_mux2_1 _3553_ (.A0(_1351_),
    .A1(\GUScpu0.regs[7][11] ),
    .S(net750),
    .X(_0362_));
 sg13g2_mux2_1 _3554_ (.A0(_1353_),
    .A1(\GUScpu0.regs[7][12] ),
    .S(net750),
    .X(_0363_));
 sg13g2_mux2_1 _3555_ (.A0(_1355_),
    .A1(\GUScpu0.regs[7][13] ),
    .S(net750),
    .X(_0364_));
 sg13g2_mux2_1 _3556_ (.A0(_1357_),
    .A1(\GUScpu0.regs[7][14] ),
    .S(net750),
    .X(_0365_));
 sg13g2_mux2_1 _3557_ (.A0(_1359_),
    .A1(\GUScpu0.regs[7][15] ),
    .S(net750),
    .X(_0366_));
 sg13g2_nand2_1 _3558_ (.Y(_1445_),
    .A(net871),
    .B(\GUScpu0.PC0[0] ));
 sg13g2_o21ai_1 _3559_ (.B1(_1445_),
    .Y(_0391_),
    .A1(net871),
    .A2(_1390_));
 sg13g2_mux2_1 _3560_ (.A0(\GUScpu0.PC0[1] ),
    .A1(_1393_),
    .S(_1472_),
    .X(_0392_));
 sg13g2_mux2_1 _3561_ (.A0(\GUScpu0.PC0[2] ),
    .A1(_1152_),
    .S(_1472_),
    .X(_0393_));
 sg13g2_nand2_1 _3562_ (.Y(_1446_),
    .A(net874),
    .B(\GUScpu0.PC0[3] ));
 sg13g2_o21ai_1 _3563_ (.B1(_1446_),
    .Y(_0394_),
    .A1(net874),
    .A2(_1166_));
 sg13g2_nand2_1 _3564_ (.Y(_1447_),
    .A(net872),
    .B(\GUScpu0.PC0[4] ));
 sg13g2_o21ai_1 _3565_ (.B1(_1447_),
    .Y(_0395_),
    .A1(net872),
    .A2(_1179_));
 sg13g2_nand2_1 _3566_ (.Y(_1448_),
    .A(\GUScpu0.PC0[5] ),
    .B(net872));
 sg13g2_o21ai_1 _3567_ (.B1(_1448_),
    .Y(_0396_),
    .A1(net872),
    .A2(_1397_));
 sg13g2_nand2_1 _3568_ (.Y(_1449_),
    .A(net874),
    .B(\GUScpu0.PC0[6] ));
 sg13g2_o21ai_1 _3569_ (.B1(_1449_),
    .Y(_0397_),
    .A1(net874),
    .A2(_1400_));
 sg13g2_nand2_1 _3570_ (.Y(_1450_),
    .A(net874),
    .B(\GUScpu0.PC0[7] ));
 sg13g2_o21ai_1 _3571_ (.B1(_1450_),
    .Y(_0398_),
    .A1(net874),
    .A2(_1405_));
 sg13g2_nand2_1 _3572_ (.Y(_1451_),
    .A(net875),
    .B(\GUScpu0.PC0[8] ));
 sg13g2_o21ai_1 _3573_ (.B1(_1451_),
    .Y(_0399_),
    .A1(net875),
    .A2(_1409_));
 sg13g2_nand2_1 _3574_ (.Y(_1452_),
    .A(net878),
    .B(\GUScpu0.PC0[9] ));
 sg13g2_o21ai_1 _3575_ (.B1(_1452_),
    .Y(_0400_),
    .A1(net878),
    .A2(_1413_));
 sg13g2_nand2_1 _3576_ (.Y(_1453_),
    .A(net877),
    .B(\GUScpu0.PC0[10] ));
 sg13g2_o21ai_1 _3577_ (.B1(_1453_),
    .Y(_0401_),
    .A1(net877),
    .A2(_1422_));
 sg13g2_nand2_1 _3578_ (.Y(_1454_),
    .A(net877),
    .B(\GUScpu0.PC0[11] ));
 sg13g2_o21ai_1 _3579_ (.B1(_1454_),
    .Y(_0402_),
    .A1(net877),
    .A2(_1426_));
 sg13g2_nand2_1 _3580_ (.Y(_1455_),
    .A(net876),
    .B(\GUScpu0.PC0[12] ));
 sg13g2_o21ai_1 _3581_ (.B1(_1455_),
    .Y(_0403_),
    .A1(net876),
    .A2(_1430_));
 sg13g2_nand2_1 _3582_ (.Y(_1456_),
    .A(net876),
    .B(\GUScpu0.PC0[13] ));
 sg13g2_o21ai_1 _3583_ (.B1(_1456_),
    .Y(_0404_),
    .A1(net877),
    .A2(_1434_));
 sg13g2_nand2_1 _3584_ (.Y(_1457_),
    .A(net876),
    .B(\GUScpu0.PC0[14] ));
 sg13g2_o21ai_1 _3585_ (.B1(_1457_),
    .Y(_0405_),
    .A1(net876),
    .A2(_1438_));
 sg13g2_nand2_1 _3586_ (.Y(_1458_),
    .A(net875),
    .B(\GUScpu0.PC0[15] ));
 sg13g2_o21ai_1 _3587_ (.B1(_1458_),
    .Y(_0406_),
    .A1(net875),
    .A2(_1441_));
 sg13g2_nand4_1 _3588_ (.B(net883),
    .C(net849),
    .A(_0089_),
    .Y(_1459_),
    .D(_1324_));
 sg13g2_mux2_1 _3589_ (.A0(_1329_),
    .A1(\GUScpu0.regs[1][0] ),
    .S(net737),
    .X(_0407_));
 sg13g2_mux2_1 _3590_ (.A0(_1331_),
    .A1(\GUScpu0.regs[1][1] ),
    .S(net738),
    .X(_0408_));
 sg13g2_mux2_1 _3591_ (.A0(_1333_),
    .A1(\GUScpu0.regs[1][2] ),
    .S(net737),
    .X(_0409_));
 sg13g2_mux2_1 _3592_ (.A0(_1335_),
    .A1(\GUScpu0.regs[1][3] ),
    .S(net737),
    .X(_0410_));
 sg13g2_mux2_1 _3593_ (.A0(_1337_),
    .A1(\GUScpu0.regs[1][4] ),
    .S(net737),
    .X(_0411_));
 sg13g2_mux2_1 _3594_ (.A0(_1339_),
    .A1(\GUScpu0.regs[1][5] ),
    .S(net737),
    .X(_0412_));
 sg13g2_mux2_1 _3595_ (.A0(_1341_),
    .A1(\GUScpu0.regs[1][6] ),
    .S(net737),
    .X(_0413_));
 sg13g2_mux2_1 _3596_ (.A0(_1343_),
    .A1(\GUScpu0.regs[1][7] ),
    .S(net737),
    .X(_0414_));
 sg13g2_mux2_1 _3597_ (.A0(_1345_),
    .A1(\GUScpu0.regs[1][8] ),
    .S(_1459_),
    .X(_0415_));
 sg13g2_mux2_1 _3598_ (.A0(_1347_),
    .A1(\GUScpu0.regs[1][9] ),
    .S(net738),
    .X(_0416_));
 sg13g2_mux2_1 _3599_ (.A0(_1349_),
    .A1(\GUScpu0.regs[1][10] ),
    .S(net738),
    .X(_0417_));
 sg13g2_mux2_1 _3600_ (.A0(_1351_),
    .A1(\GUScpu0.regs[1][11] ),
    .S(net738),
    .X(_0418_));
 sg13g2_mux2_1 _3601_ (.A0(_1353_),
    .A1(\GUScpu0.regs[1][12] ),
    .S(net738),
    .X(_0419_));
 sg13g2_mux2_1 _3602_ (.A0(_1355_),
    .A1(\GUScpu0.regs[1][13] ),
    .S(net738),
    .X(_0420_));
 sg13g2_mux2_1 _3603_ (.A0(_1357_),
    .A1(\GUScpu0.regs[1][14] ),
    .S(net738),
    .X(_0421_));
 sg13g2_mux2_1 _3604_ (.A0(_1359_),
    .A1(\GUScpu0.regs[1][15] ),
    .S(net737),
    .X(_0422_));
 sg13g2_dfrbp_1 _3605_ (.CLK(net902),
    .RESET_B(net45),
    .D(_0192_),
    .Q_N(_1815_),
    .Q(\GUScpu0.zn[1][0] ));
 sg13g2_dfrbp_1 _3606_ (.CLK(net903),
    .RESET_B(net105),
    .D(_0193_),
    .Q_N(_1814_),
    .Q(\GUScpu0.zn[1][1] ));
 sg13g2_dfrbp_1 _3607_ (.CLK(clknet_1_0__leaf_clk_regs),
    .RESET_B(net104),
    .D(_0194_),
    .Q_N(_1813_),
    .Q(\xdi[0] ));
 sg13g2_dfrbp_1 _3608_ (.CLK(clknet_1_1__leaf_clk_regs),
    .RESET_B(net103),
    .D(net222),
    .Q_N(_1812_),
    .Q(\xdi[1] ));
 sg13g2_dfrbp_1 _3609_ (.CLK(clknet_1_1__leaf_clk_regs),
    .RESET_B(net102),
    .D(_0196_),
    .Q_N(_1811_),
    .Q(\xdi[2] ));
 sg13g2_dfrbp_1 _3610_ (.CLK(clknet_1_0__leaf_clk_regs),
    .RESET_B(net101),
    .D(_0197_),
    .Q_N(_1810_),
    .Q(\xdi[3] ));
 sg13g2_dfrbp_1 _3611_ (.CLK(clknet_1_0__leaf_clk_regs),
    .RESET_B(net100),
    .D(_0198_),
    .Q_N(_1809_),
    .Q(\xdi[4] ));
 sg13g2_dfrbp_1 _3612_ (.CLK(clknet_1_1__leaf_clk_regs),
    .RESET_B(net99),
    .D(_0199_),
    .Q_N(_1808_),
    .Q(\xdi[5] ));
 sg13g2_dfrbp_1 _3613_ (.CLK(clknet_1_1__leaf_clk_regs),
    .RESET_B(net98),
    .D(_0200_),
    .Q_N(_1807_),
    .Q(\xdi[6] ));
 sg13g2_dfrbp_1 _3614_ (.CLK(clknet_1_1__leaf_clk_regs),
    .RESET_B(net97),
    .D(_0201_),
    .Q_N(_1806_),
    .Q(\xdi[7] ));
 sg13g2_dfrbp_1 _3615_ (.CLK(net898),
    .RESET_B(net96),
    .D(_0202_),
    .Q_N(_0140_),
    .Q(\GUScpu0.regs[5][0] ));
 sg13g2_dfrbp_1 _3616_ (.CLK(net895),
    .RESET_B(net95),
    .D(_0203_),
    .Q_N(_0131_),
    .Q(\GUScpu0.regs[5][1] ));
 sg13g2_dfrbp_1 _3617_ (.CLK(net899),
    .RESET_B(net94),
    .D(_0204_),
    .Q_N(_0123_),
    .Q(\GUScpu0.regs[5][2] ));
 sg13g2_dfrbp_1 _3618_ (.CLK(net892),
    .RESET_B(net93),
    .D(_0205_),
    .Q_N(_0115_),
    .Q(\GUScpu0.regs[5][3] ));
 sg13g2_dfrbp_1 _3619_ (.CLK(net892),
    .RESET_B(net92),
    .D(_0206_),
    .Q_N(_0107_),
    .Q(\GUScpu0.regs[5][4] ));
 sg13g2_dfrbp_1 _3620_ (.CLK(net889),
    .RESET_B(net91),
    .D(_0207_),
    .Q_N(_0096_),
    .Q(\GUScpu0.regs[5][5] ));
 sg13g2_dfrbp_1 _3621_ (.CLK(net908),
    .RESET_B(net90),
    .D(_0208_),
    .Q_N(_0148_),
    .Q(\GUScpu0.regs[5][6] ));
 sg13g2_dfrbp_1 _3622_ (.CLK(net893),
    .RESET_B(net89),
    .D(_0209_),
    .Q_N(_0156_),
    .Q(\GUScpu0.regs[5][7] ));
 sg13g2_dfrbp_1 _3623_ (.CLK(net907),
    .RESET_B(net88),
    .D(_0210_),
    .Q_N(_0164_),
    .Q(\GUScpu0.regs[5][8] ));
 sg13g2_dfrbp_1 _3624_ (.CLK(net906),
    .RESET_B(net87),
    .D(_0211_),
    .Q_N(_0026_),
    .Q(\GUScpu0.regs[5][9] ));
 sg13g2_dfrbp_1 _3625_ (.CLK(net909),
    .RESET_B(net86),
    .D(_0212_),
    .Q_N(_0034_),
    .Q(\GUScpu0.regs[5][10] ));
 sg13g2_dfrbp_1 _3626_ (.CLK(net906),
    .RESET_B(net85),
    .D(_0213_),
    .Q_N(_0042_),
    .Q(\GUScpu0.regs[5][11] ));
 sg13g2_dfrbp_1 _3627_ (.CLK(net909),
    .RESET_B(net84),
    .D(_0214_),
    .Q_N(_0050_),
    .Q(\GUScpu0.regs[5][12] ));
 sg13g2_dfrbp_1 _3628_ (.CLK(net913),
    .RESET_B(net83),
    .D(_0215_),
    .Q_N(_0058_),
    .Q(\GUScpu0.regs[5][13] ));
 sg13g2_dfrbp_1 _3629_ (.CLK(net913),
    .RESET_B(net82),
    .D(_0216_),
    .Q_N(_0066_),
    .Q(\GUScpu0.regs[5][14] ));
 sg13g2_dfrbp_1 _3630_ (.CLK(net894),
    .RESET_B(net81),
    .D(_0217_),
    .Q_N(_0074_),
    .Q(\GUScpu0.regs[5][15] ));
 sg13g2_dfrbp_1 _3631_ (.CLK(net889),
    .RESET_B(net80),
    .D(_0218_),
    .Q_N(_0141_),
    .Q(\GUScpu0.regs[6][0] ));
 sg13g2_dfrbp_1 _3632_ (.CLK(net895),
    .RESET_B(net79),
    .D(_0219_),
    .Q_N(_0132_),
    .Q(\GUScpu0.regs[6][1] ));
 sg13g2_dfrbp_1 _3633_ (.CLK(net899),
    .RESET_B(net78),
    .D(_0220_),
    .Q_N(_0124_),
    .Q(\GUScpu0.regs[6][2] ));
 sg13g2_dfrbp_1 _3634_ (.CLK(net892),
    .RESET_B(net77),
    .D(_0221_),
    .Q_N(_0116_),
    .Q(\GUScpu0.regs[6][3] ));
 sg13g2_dfrbp_1 _3635_ (.CLK(net890),
    .RESET_B(net76),
    .D(_0222_),
    .Q_N(_0108_),
    .Q(\GUScpu0.regs[6][4] ));
 sg13g2_dfrbp_1 _3636_ (.CLK(net888),
    .RESET_B(net75),
    .D(_0223_),
    .Q_N(_0097_),
    .Q(\GUScpu0.regs[6][5] ));
 sg13g2_dfrbp_1 _3637_ (.CLK(net896),
    .RESET_B(net74),
    .D(_0224_),
    .Q_N(_0149_),
    .Q(\GUScpu0.regs[6][6] ));
 sg13g2_dfrbp_1 _3638_ (.CLK(net893),
    .RESET_B(net53),
    .D(_0225_),
    .Q_N(_0157_),
    .Q(\GUScpu0.regs[6][7] ));
 sg13g2_dfrbp_1 _3639_ (.CLK(net907),
    .RESET_B(net52),
    .D(_0226_),
    .Q_N(_0165_),
    .Q(\GUScpu0.regs[6][8] ));
 sg13g2_dfrbp_1 _3640_ (.CLK(net912),
    .RESET_B(net51),
    .D(_0227_),
    .Q_N(_0027_),
    .Q(\GUScpu0.regs[6][9] ));
 sg13g2_dfrbp_1 _3641_ (.CLK(net912),
    .RESET_B(net50),
    .D(_0228_),
    .Q_N(_0035_),
    .Q(\GUScpu0.regs[6][10] ));
 sg13g2_dfrbp_1 _3642_ (.CLK(net908),
    .RESET_B(net49),
    .D(_0229_),
    .Q_N(_0043_),
    .Q(\GUScpu0.regs[6][11] ));
 sg13g2_dfrbp_1 _3643_ (.CLK(net911),
    .RESET_B(net48),
    .D(_0230_),
    .Q_N(_0051_),
    .Q(\GUScpu0.regs[6][12] ));
 sg13g2_dfrbp_1 _3644_ (.CLK(net914),
    .RESET_B(net47),
    .D(_0231_),
    .Q_N(_0059_),
    .Q(\GUScpu0.regs[6][13] ));
 sg13g2_dfrbp_1 _3645_ (.CLK(net913),
    .RESET_B(net46),
    .D(_0232_),
    .Q_N(_0067_),
    .Q(\GUScpu0.regs[6][14] ));
 sg13g2_dfrbp_1 _3646_ (.CLK(net894),
    .RESET_B(net44),
    .D(_0233_),
    .Q_N(_0075_),
    .Q(\GUScpu0.regs[6][15] ));
 sg13g2_dfrbp_1 _3647_ (.CLK(net888),
    .RESET_B(net43),
    .D(_0234_),
    .Q_N(_0135_),
    .Q(\GUScpu0.regs[0][0] ));
 sg13g2_dfrbp_1 _3648_ (.CLK(net895),
    .RESET_B(net42),
    .D(_0235_),
    .Q_N(_0126_),
    .Q(\GUScpu0.regs[0][1] ));
 sg13g2_dfrbp_1 _3649_ (.CLK(net899),
    .RESET_B(net41),
    .D(_0236_),
    .Q_N(_0118_),
    .Q(\GUScpu0.regs[0][2] ));
 sg13g2_dfrbp_1 _3650_ (.CLK(net891),
    .RESET_B(net40),
    .D(_0237_),
    .Q_N(_0110_),
    .Q(\GUScpu0.regs[0][3] ));
 sg13g2_dfrbp_1 _3651_ (.CLK(net890),
    .RESET_B(net39),
    .D(_0238_),
    .Q_N(_0102_),
    .Q(\GUScpu0.regs[0][4] ));
 sg13g2_dfrbp_1 _3652_ (.CLK(net889),
    .RESET_B(net38),
    .D(_0239_),
    .Q_N(_0085_),
    .Q(\GUScpu0.regs[0][5] ));
 sg13g2_dfrbp_1 _3653_ (.CLK(net896),
    .RESET_B(net37),
    .D(_0240_),
    .Q_N(_0143_),
    .Q(\GUScpu0.regs[0][6] ));
 sg13g2_dfrbp_1 _3654_ (.CLK(net893),
    .RESET_B(net36),
    .D(_0241_),
    .Q_N(_0151_),
    .Q(\GUScpu0.regs[0][7] ));
 sg13g2_dfrbp_1 _3655_ (.CLK(net907),
    .RESET_B(net35),
    .D(_0242_),
    .Q_N(_0159_),
    .Q(\GUScpu0.regs[0][8] ));
 sg13g2_dfrbp_1 _3656_ (.CLK(net909),
    .RESET_B(net34),
    .D(_0243_),
    .Q_N(_0167_),
    .Q(\GUScpu0.regs[0][9] ));
 sg13g2_dfrbp_1 _3657_ (.CLK(net910),
    .RESET_B(net33),
    .D(_0244_),
    .Q_N(_0029_),
    .Q(\GUScpu0.regs[0][10] ));
 sg13g2_dfrbp_1 _3658_ (.CLK(net906),
    .RESET_B(net32),
    .D(_0245_),
    .Q_N(_0037_),
    .Q(\GUScpu0.regs[0][11] ));
 sg13g2_dfrbp_1 _3659_ (.CLK(net910),
    .RESET_B(net31),
    .D(_0246_),
    .Q_N(_0045_),
    .Q(\GUScpu0.regs[0][12] ));
 sg13g2_dfrbp_1 _3660_ (.CLK(net911),
    .RESET_B(net30),
    .D(_0247_),
    .Q_N(_0053_),
    .Q(\GUScpu0.regs[0][13] ));
 sg13g2_dfrbp_1 _3661_ (.CLK(net914),
    .RESET_B(net29),
    .D(_0248_),
    .Q_N(_0061_),
    .Q(\GUScpu0.regs[0][14] ));
 sg13g2_dfrbp_1 _3662_ (.CLK(net894),
    .RESET_B(net28),
    .D(_0249_),
    .Q_N(_0069_),
    .Q(\GUScpu0.regs[0][15] ));
 sg13g2_dfrbp_1 _3663_ (.CLK(net902),
    .RESET_B(net27),
    .D(_0250_),
    .Q_N(_1805_),
    .Q(\GUScpu0.cv[0][0] ));
 sg13g2_dfrbp_1 _3664_ (.CLK(net902),
    .RESET_B(net26),
    .D(_0251_),
    .Q_N(_1804_),
    .Q(\GUScpu0.cv[0][1] ));
 sg13g2_dfrbp_1 _3665_ (.CLK(net920),
    .RESET_B(net25),
    .D(_0252_),
    .Q_N(_1803_),
    .Q(sdty));
 sg13g2_dfrbp_1 _3666_ (.CLK(net930),
    .RESET_B(net944),
    .D(_0253_),
    .Q_N(txd),
    .Q(_0172_));
 sg13g2_dfrbp_1 _3667_ (.CLK(net929),
    .RESET_B(net940),
    .D(_0254_),
    .Q_N(\uart0.txsh[1] ),
    .Q(_0173_));
 sg13g2_dfrbp_1 _3668_ (.CLK(net926),
    .RESET_B(net938),
    .D(_0255_),
    .Q_N(\uart0.txsh[2] ),
    .Q(_0174_));
 sg13g2_dfrbp_1 _3669_ (.CLK(net926),
    .RESET_B(net938),
    .D(_0256_),
    .Q_N(\uart0.txsh[3] ),
    .Q(_0175_));
 sg13g2_dfrbp_1 _3670_ (.CLK(net927),
    .RESET_B(net939),
    .D(_0257_),
    .Q_N(\uart0.txsh[4] ),
    .Q(_0176_));
 sg13g2_dfrbp_1 _3671_ (.CLK(net927),
    .RESET_B(net938),
    .D(_0258_),
    .Q_N(\uart0.txsh[5] ),
    .Q(_0177_));
 sg13g2_dfrbp_1 _3672_ (.CLK(net927),
    .RESET_B(net938),
    .D(_0259_),
    .Q_N(\uart0.txsh[6] ),
    .Q(_0178_));
 sg13g2_dfrbp_1 _3673_ (.CLK(net927),
    .RESET_B(net939),
    .D(_0260_),
    .Q_N(\uart0.txsh[7] ),
    .Q(_0179_));
 sg13g2_dfrbp_1 _3674_ (.CLK(net927),
    .RESET_B(net939),
    .D(_0261_),
    .Q_N(\uart0.txsh[8] ),
    .Q(_0180_));
 sg13g2_dfrbp_1 _3675_ (.CLK(net924),
    .RESET_B(net936),
    .D(_0000_),
    .Q_N(_1802_),
    .Q(\pwmc[0] ));
 sg13g2_dfrbp_1 _3676_ (.CLK(net925),
    .RESET_B(net936),
    .D(_0001_),
    .Q_N(_1801_),
    .Q(\pwmc[1] ));
 sg13g2_dfrbp_1 _3677_ (.CLK(net924),
    .RESET_B(net937),
    .D(_0002_),
    .Q_N(_1800_),
    .Q(\pwmc[2] ));
 sg13g2_dfrbp_1 _3678_ (.CLK(net924),
    .RESET_B(net936),
    .D(_0003_),
    .Q_N(_1799_),
    .Q(\pwmc[3] ));
 sg13g2_dfrbp_1 _3679_ (.CLK(net925),
    .RESET_B(net936),
    .D(_0004_),
    .Q_N(_1798_),
    .Q(\pwmc[4] ));
 sg13g2_dfrbp_1 _3680_ (.CLK(net925),
    .RESET_B(net936),
    .D(_0005_),
    .Q_N(_1797_),
    .Q(\pwmc[5] ));
 sg13g2_dfrbp_1 _3681_ (.CLK(net925),
    .RESET_B(net936),
    .D(_0006_),
    .Q_N(_1796_),
    .Q(\pwmc[6] ));
 sg13g2_dfrbp_1 _3682_ (.CLK(net925),
    .RESET_B(net936),
    .D(_0007_),
    .Q_N(_0078_),
    .Q(\pwmc[7] ));
 sg13g2_dfrbp_1 _3683_ (.CLK(net920),
    .RESET_B(net212),
    .D(_0262_),
    .Q_N(_1795_),
    .Q(gpo));
 sg13g2_dfrbp_1 _3684_ (.CLK(net924),
    .RESET_B(net211),
    .D(_0263_),
    .Q_N(_1794_),
    .Q(\pwmbuf[0] ));
 sg13g2_dfrbp_1 _3685_ (.CLK(net925),
    .RESET_B(net209),
    .D(_0264_),
    .Q_N(_1793_),
    .Q(\pwmbuf[1] ));
 sg13g2_dfrbp_1 _3686_ (.CLK(net924),
    .RESET_B(net207),
    .D(_0265_),
    .Q_N(_1792_),
    .Q(\pwmbuf[2] ));
 sg13g2_dfrbp_1 _3687_ (.CLK(net924),
    .RESET_B(net205),
    .D(_0266_),
    .Q_N(_1791_),
    .Q(\pwmbuf[3] ));
 sg13g2_dfrbp_1 _3688_ (.CLK(net924),
    .RESET_B(net203),
    .D(_0267_),
    .Q_N(_1790_),
    .Q(\pwmbuf[4] ));
 sg13g2_dfrbp_1 _3689_ (.CLK(net924),
    .RESET_B(net201),
    .D(_0268_),
    .Q_N(_1789_),
    .Q(\pwmbuf[5] ));
 sg13g2_dfrbp_1 _3690_ (.CLK(net925),
    .RESET_B(net199),
    .D(_0269_),
    .Q_N(_1788_),
    .Q(\pwmbuf[6] ));
 sg13g2_dfrbp_1 _3691_ (.CLK(net928),
    .RESET_B(net197),
    .D(_0270_),
    .Q_N(_1787_),
    .Q(\pwmbuf[7] ));
 sg13g2_dfrbp_1 _3692_ (.CLK(net928),
    .RESET_B(net937),
    .D(_0271_),
    .Q_N(_1786_),
    .Q(pwmout));
 sg13g2_dfrbp_1 _3693_ (.CLK(net930),
    .RESET_B(net939),
    .D(_0272_),
    .Q_N(_1785_),
    .Q(pwmirq));
 sg13g2_dfrbp_1 _3694_ (.CLK(net905),
    .RESET_B(net194),
    .D(_0273_),
    .Q_N(_1784_),
    .Q(\pwmhold[0] ));
 sg13g2_dfrbp_1 _3695_ (.CLK(net903),
    .RESET_B(net193),
    .D(_0274_),
    .Q_N(_1783_),
    .Q(\pwmhold[1] ));
 sg13g2_dfrbp_1 _3696_ (.CLK(net904),
    .RESET_B(net192),
    .D(_0275_),
    .Q_N(_1782_),
    .Q(\pwmhold[2] ));
 sg13g2_dfrbp_1 _3697_ (.CLK(net902),
    .RESET_B(net191),
    .D(_0276_),
    .Q_N(_1781_),
    .Q(\pwmhold[3] ));
 sg13g2_dfrbp_1 _3698_ (.CLK(net904),
    .RESET_B(net190),
    .D(_0277_),
    .Q_N(_1780_),
    .Q(\pwmhold[4] ));
 sg13g2_dfrbp_1 _3699_ (.CLK(net902),
    .RESET_B(net189),
    .D(_0278_),
    .Q_N(_1779_),
    .Q(\pwmhold[5] ));
 sg13g2_dfrbp_1 _3700_ (.CLK(net904),
    .RESET_B(net188),
    .D(_0279_),
    .Q_N(_1778_),
    .Q(\pwmhold[6] ));
 sg13g2_dfrbp_1 _3701_ (.CLK(net904),
    .RESET_B(net187),
    .D(_0280_),
    .Q_N(_1777_),
    .Q(\pwmhold[7] ));
 sg13g2_dfrbp_1 _3702_ (.CLK(net920),
    .RESET_B(net943),
    .D(_0281_),
    .Q_N(_1776_),
    .Q(\irqen[0] ));
 sg13g2_dfrbp_1 _3703_ (.CLK(net920),
    .RESET_B(net943),
    .D(_0282_),
    .Q_N(_1775_),
    .Q(\irqen[1] ));
 sg13g2_dfrbp_1 _3704_ (.CLK(net920),
    .RESET_B(net943),
    .D(_0283_),
    .Q_N(_1774_),
    .Q(\irqen[2] ));
 sg13g2_dfrbp_1 _3705_ (.CLK(net917),
    .RESET_B(net943),
    .D(_0284_),
    .Q_N(_1773_),
    .Q(\irqen[3] ));
 sg13g2_dfrbp_1 _3706_ (.CLK(net916),
    .RESET_B(net943),
    .D(_0285_),
    .Q_N(_1816_),
    .Q(\irqen[4] ));
 sg13g2_dfrbp_1 _3707_ (.CLK(clknet_1_0__leaf_clk_regs),
    .RESET_B(net942),
    .D(net220),
    .Q_N(_1712_),
    .Q(\ckd[0] ));
 sg13g2_dfrbp_1 _3708_ (.CLK(clknet_1_0__leaf_clk_regs),
    .RESET_B(net942),
    .D(_0171_),
    .Q_N(_0080_),
    .Q(\ckd[1] ));
 sg13g2_dfrbp_1 _3709_ (.CLK(net929),
    .RESET_B(net943),
    .D(_0191_),
    .Q_N(\uart0.urxsh[0] ),
    .Q(_0181_));
 sg13g2_dfrbp_1 _3710_ (.CLK(net903),
    .RESET_B(net186),
    .D(_0286_),
    .Q_N(_1772_),
    .Q(\GUScpu0.PC1[0] ));
 sg13g2_dfrbp_1 _3711_ (.CLK(net915),
    .RESET_B(net185),
    .D(_0287_),
    .Q_N(_1771_),
    .Q(\GUScpu0.PC1[1] ));
 sg13g2_dfrbp_1 _3712_ (.CLK(net915),
    .RESET_B(net184),
    .D(_0288_),
    .Q_N(_1770_),
    .Q(\GUScpu0.PC1[5] ));
 sg13g2_dfrbp_1 _3713_ (.CLK(net917),
    .RESET_B(net183),
    .D(_0289_),
    .Q_N(_1769_),
    .Q(\GUScpu0.PC1[6] ));
 sg13g2_dfrbp_1 _3714_ (.CLK(net916),
    .RESET_B(net182),
    .D(_0290_),
    .Q_N(_1768_),
    .Q(\GUScpu0.PC1[7] ));
 sg13g2_dfrbp_1 _3715_ (.CLK(net917),
    .RESET_B(net181),
    .D(_0291_),
    .Q_N(_1767_),
    .Q(\GUScpu0.PC1[8] ));
 sg13g2_dfrbp_1 _3716_ (.CLK(net919),
    .RESET_B(net54),
    .D(_0292_),
    .Q_N(_1817_),
    .Q(\GUScpu0.PC1[9] ));
 sg13g2_dfrbp_1 _3717_ (.CLK(net915),
    .RESET_B(net55),
    .D(_0008_),
    .Q_N(_1818_),
    .Q(\GUScpu0.PC1[2] ));
 sg13g2_dfrbp_1 _3718_ (.CLK(net916),
    .RESET_B(net56),
    .D(_0009_),
    .Q_N(_1819_),
    .Q(\GUScpu0.PC1[3] ));
 sg13g2_dfrbp_1 _3719_ (.CLK(net915),
    .RESET_B(net57),
    .D(_0010_),
    .Q_N(_1820_),
    .Q(\GUScpu0.PC1[4] ));
 sg13g2_dfrbp_1 _3720_ (.CLK(net900),
    .RESET_B(net58),
    .D(\GUScpu0.cdi[0] ),
    .Q_N(_0134_),
    .Q(\GUScpu0.IR[0] ));
 sg13g2_dfrbp_1 _3721_ (.CLK(net915),
    .RESET_B(net59),
    .D(\GUScpu0.cdi[1] ),
    .Q_N(_1821_),
    .Q(\GUScpu0.IR[1] ));
 sg13g2_dfrbp_1 _3722_ (.CLK(net900),
    .RESET_B(net60),
    .D(\GUScpu0.cdi[2] ),
    .Q_N(_0088_),
    .Q(\GUScpu0.IR[2] ));
 sg13g2_dfrbp_1 _3723_ (.CLK(net900),
    .RESET_B(net61),
    .D(\GUScpu0.cdi[3] ),
    .Q_N(_0090_),
    .Q(\GUScpu0.IR[3] ));
 sg13g2_dfrbp_1 _3724_ (.CLK(net901),
    .RESET_B(net62),
    .D(\GUScpu0.cdi[4] ),
    .Q_N(_0094_),
    .Q(\GUScpu0.IR[4] ));
 sg13g2_dfrbp_1 _3725_ (.CLK(net900),
    .RESET_B(net63),
    .D(\GUScpu0.cdi[5] ),
    .Q_N(_0099_),
    .Q(\GUScpu0.IR[5] ));
 sg13g2_dfrbp_1 _3726_ (.CLK(net900),
    .RESET_B(net64),
    .D(\GUScpu0.cdi[6] ),
    .Q_N(_0100_),
    .Q(\GUScpu0.IR[6] ));
 sg13g2_dfrbp_1 _3727_ (.CLK(net900),
    .RESET_B(net65),
    .D(\GUScpu0.cdi[7] ),
    .Q_N(_0101_),
    .Q(\GUScpu0.IR[7] ));
 sg13g2_dfrbp_1 _3728_ (.CLK(net900),
    .RESET_B(net66),
    .D(\GUScpu0.cdi[8] ),
    .Q_N(_0087_),
    .Q(\GUScpu0.IR[8] ));
 sg13g2_dfrbp_1 _3729_ (.CLK(net908),
    .RESET_B(net67),
    .D(\GUScpu0.cdi[9] ),
    .Q_N(_0089_),
    .Q(\GUScpu0.IR[9] ));
 sg13g2_dfrbp_1 _3730_ (.CLK(net917),
    .RESET_B(net68),
    .D(\GUScpu0.cdi[10] ),
    .Q_N(_0093_),
    .Q(\GUScpu0.IR[10] ));
 sg13g2_dfrbp_1 _3731_ (.CLK(net900),
    .RESET_B(net69),
    .D(\GUScpu0.cdi[11] ),
    .Q_N(_1822_),
    .Q(\GUScpu0.IR[11] ));
 sg13g2_dfrbp_1 _3732_ (.CLK(net901),
    .RESET_B(net70),
    .D(\GUScpu0.cdi[12] ),
    .Q_N(_0079_),
    .Q(\GUScpu0.IR[12] ));
 sg13g2_dfrbp_1 _3733_ (.CLK(net902),
    .RESET_B(net71),
    .D(\GUScpu0.cdi[13] ),
    .Q_N(_1823_),
    .Q(\GUScpu0.IR[13] ));
 sg13g2_dfrbp_1 _3734_ (.CLK(net899),
    .RESET_B(net72),
    .D(\GUScpu0.cdi[14] ),
    .Q_N(_1824_),
    .Q(\GUScpu0.IR[14] ));
 sg13g2_dfrbp_1 _3735_ (.CLK(net901),
    .RESET_B(net73),
    .D(\GUScpu0.cdi[15] ),
    .Q_N(_0084_),
    .Q(\GUScpu0.IR[15] ));
 sg13g2_dfrbp_1 _3736_ (.CLK(net901),
    .RESET_B(net941),
    .D(\GUScpu0.opvali ),
    .Q_N(_0083_),
    .Q(\GUScpu0.opval ));
 sg13g2_dfrbp_1 _3737_ (.CLK(net903),
    .RESET_B(net941),
    .D(_0012_),
    .Q_N(_0081_),
    .Q(\GUScpu0.imode ));
 sg13g2_dfrbp_1 _3738_ (.CLK(net903),
    .RESET_B(net941),
    .D(_0011_),
    .Q_N(_0082_),
    .Q(\GUScpu0.irqq0 ));
 sg13g2_dfrbp_1 _3739_ (.CLK(net889),
    .RESET_B(net180),
    .D(_0293_),
    .Q_N(_0139_),
    .Q(\GUScpu0.regs[4][0] ));
 sg13g2_dfrbp_1 _3740_ (.CLK(net895),
    .RESET_B(net179),
    .D(_0294_),
    .Q_N(_0130_),
    .Q(\GUScpu0.regs[4][1] ));
 sg13g2_dfrbp_1 _3741_ (.CLK(net899),
    .RESET_B(net178),
    .D(_0295_),
    .Q_N(_0122_),
    .Q(\GUScpu0.regs[4][2] ));
 sg13g2_dfrbp_1 _3742_ (.CLK(net890),
    .RESET_B(net177),
    .D(_0296_),
    .Q_N(_0114_),
    .Q(\GUScpu0.regs[4][3] ));
 sg13g2_dfrbp_1 _3743_ (.CLK(net892),
    .RESET_B(net176),
    .D(_0297_),
    .Q_N(_0106_),
    .Q(\GUScpu0.regs[4][4] ));
 sg13g2_dfrbp_1 _3744_ (.CLK(net888),
    .RESET_B(net175),
    .D(_0298_),
    .Q_N(_0095_),
    .Q(\GUScpu0.regs[4][5] ));
 sg13g2_dfrbp_1 _3745_ (.CLK(net908),
    .RESET_B(net174),
    .D(_0299_),
    .Q_N(_0147_),
    .Q(\GUScpu0.regs[4][6] ));
 sg13g2_dfrbp_1 _3746_ (.CLK(net893),
    .RESET_B(net173),
    .D(_0300_),
    .Q_N(_0155_),
    .Q(\GUScpu0.regs[4][7] ));
 sg13g2_dfrbp_1 _3747_ (.CLK(net907),
    .RESET_B(net172),
    .D(_0301_),
    .Q_N(_0163_),
    .Q(\GUScpu0.regs[4][8] ));
 sg13g2_dfrbp_1 _3748_ (.CLK(net906),
    .RESET_B(net171),
    .D(_0302_),
    .Q_N(_0025_),
    .Q(\GUScpu0.regs[4][9] ));
 sg13g2_dfrbp_1 _3749_ (.CLK(net909),
    .RESET_B(net170),
    .D(_0303_),
    .Q_N(_0033_),
    .Q(\GUScpu0.regs[4][10] ));
 sg13g2_dfrbp_1 _3750_ (.CLK(net906),
    .RESET_B(net169),
    .D(_0304_),
    .Q_N(_0041_),
    .Q(\GUScpu0.regs[4][11] ));
 sg13g2_dfrbp_1 _3751_ (.CLK(net909),
    .RESET_B(net168),
    .D(_0305_),
    .Q_N(_0049_),
    .Q(\GUScpu0.regs[4][12] ));
 sg13g2_dfrbp_1 _3752_ (.CLK(net913),
    .RESET_B(net167),
    .D(_0306_),
    .Q_N(_0057_),
    .Q(\GUScpu0.regs[4][13] ));
 sg13g2_dfrbp_1 _3753_ (.CLK(net913),
    .RESET_B(net166),
    .D(_0307_),
    .Q_N(_0065_),
    .Q(\GUScpu0.regs[4][14] ));
 sg13g2_dfrbp_1 _3754_ (.CLK(net894),
    .RESET_B(net165),
    .D(_0308_),
    .Q_N(_0073_),
    .Q(\GUScpu0.regs[4][15] ));
 sg13g2_dfrbp_1 _3755_ (.CLK(net902),
    .RESET_B(net164),
    .D(_0309_),
    .Q_N(_1766_),
    .Q(\GUScpu0.cv[1][0] ));
 sg13g2_dfrbp_1 _3756_ (.CLK(net902),
    .RESET_B(net163),
    .D(_0310_),
    .Q_N(_1765_),
    .Q(\GUScpu0.cv[1][1] ));
 sg13g2_dfrbp_1 _3757_ (.CLK(net888),
    .RESET_B(net162),
    .D(_0311_),
    .Q_N(_0138_),
    .Q(\GUScpu0.regs[3][0] ));
 sg13g2_dfrbp_1 _3758_ (.CLK(net895),
    .RESET_B(net161),
    .D(_0312_),
    .Q_N(_0129_),
    .Q(\GUScpu0.regs[3][1] ));
 sg13g2_dfrbp_1 _3759_ (.CLK(net899),
    .RESET_B(net160),
    .D(_0313_),
    .Q_N(_0121_),
    .Q(\GUScpu0.regs[3][2] ));
 sg13g2_dfrbp_1 _3760_ (.CLK(net891),
    .RESET_B(net159),
    .D(_0314_),
    .Q_N(_0113_),
    .Q(\GUScpu0.regs[3][3] ));
 sg13g2_dfrbp_1 _3761_ (.CLK(net890),
    .RESET_B(net158),
    .D(_0315_),
    .Q_N(_0105_),
    .Q(\GUScpu0.regs[3][4] ));
 sg13g2_dfrbp_1 _3762_ (.CLK(net889),
    .RESET_B(net157),
    .D(_0316_),
    .Q_N(_0092_),
    .Q(\GUScpu0.regs[3][5] ));
 sg13g2_dfrbp_1 _3763_ (.CLK(net896),
    .RESET_B(net156),
    .D(_0317_),
    .Q_N(_0146_),
    .Q(\GUScpu0.regs[3][6] ));
 sg13g2_dfrbp_1 _3764_ (.CLK(net893),
    .RESET_B(net155),
    .D(_0318_),
    .Q_N(_0154_),
    .Q(\GUScpu0.regs[3][7] ));
 sg13g2_dfrbp_1 _3765_ (.CLK(net907),
    .RESET_B(net154),
    .D(_0319_),
    .Q_N(_0162_),
    .Q(\GUScpu0.regs[3][8] ));
 sg13g2_dfrbp_1 _3766_ (.CLK(net909),
    .RESET_B(net153),
    .D(_0320_),
    .Q_N(_0170_),
    .Q(\GUScpu0.regs[3][9] ));
 sg13g2_dfrbp_1 _3767_ (.CLK(net910),
    .RESET_B(net152),
    .D(_0321_),
    .Q_N(_0032_),
    .Q(\GUScpu0.regs[3][10] ));
 sg13g2_dfrbp_1 _3768_ (.CLK(net906),
    .RESET_B(net151),
    .D(_0322_),
    .Q_N(_0040_),
    .Q(\GUScpu0.regs[3][11] ));
 sg13g2_dfrbp_1 _3769_ (.CLK(net911),
    .RESET_B(net150),
    .D(_0323_),
    .Q_N(_0048_),
    .Q(\GUScpu0.regs[3][12] ));
 sg13g2_dfrbp_1 _3770_ (.CLK(net911),
    .RESET_B(net149),
    .D(_0324_),
    .Q_N(_0056_),
    .Q(\GUScpu0.regs[3][13] ));
 sg13g2_dfrbp_1 _3771_ (.CLK(net913),
    .RESET_B(net148),
    .D(_0325_),
    .Q_N(_0064_),
    .Q(\GUScpu0.regs[3][14] ));
 sg13g2_dfrbp_1 _3772_ (.CLK(net894),
    .RESET_B(net147),
    .D(_0326_),
    .Q_N(_0072_),
    .Q(\GUScpu0.regs[3][15] ));
 sg13g2_dfrbp_1 _3773_ (.CLK(net888),
    .RESET_B(net146),
    .D(_0327_),
    .Q_N(_0137_),
    .Q(\GUScpu0.regs[2][0] ));
 sg13g2_dfrbp_1 _3774_ (.CLK(net895),
    .RESET_B(net145),
    .D(_0328_),
    .Q_N(_0128_),
    .Q(\GUScpu0.regs[2][1] ));
 sg13g2_dfrbp_1 _3775_ (.CLK(net899),
    .RESET_B(net144),
    .D(_0329_),
    .Q_N(_0120_),
    .Q(\GUScpu0.regs[2][2] ));
 sg13g2_dfrbp_1 _3776_ (.CLK(net890),
    .RESET_B(net143),
    .D(_0330_),
    .Q_N(_0112_),
    .Q(\GUScpu0.regs[2][3] ));
 sg13g2_dfrbp_1 _3777_ (.CLK(net890),
    .RESET_B(net142),
    .D(_0331_),
    .Q_N(_0104_),
    .Q(\GUScpu0.regs[2][4] ));
 sg13g2_dfrbp_1 _3778_ (.CLK(net889),
    .RESET_B(net141),
    .D(_0332_),
    .Q_N(_0091_),
    .Q(\GUScpu0.regs[2][5] ));
 sg13g2_dfrbp_1 _3779_ (.CLK(net896),
    .RESET_B(net140),
    .D(_0333_),
    .Q_N(_0145_),
    .Q(\GUScpu0.regs[2][6] ));
 sg13g2_dfrbp_1 _3780_ (.CLK(net893),
    .RESET_B(net139),
    .D(_0334_),
    .Q_N(_0153_),
    .Q(\GUScpu0.regs[2][7] ));
 sg13g2_dfrbp_1 _3781_ (.CLK(net907),
    .RESET_B(net138),
    .D(_0335_),
    .Q_N(_0161_),
    .Q(\GUScpu0.regs[2][8] ));
 sg13g2_dfrbp_1 _3782_ (.CLK(net909),
    .RESET_B(net137),
    .D(_0336_),
    .Q_N(_0169_),
    .Q(\GUScpu0.regs[2][9] ));
 sg13g2_dfrbp_1 _3783_ (.CLK(net910),
    .RESET_B(net136),
    .D(_0337_),
    .Q_N(_0031_),
    .Q(\GUScpu0.regs[2][10] ));
 sg13g2_dfrbp_1 _3784_ (.CLK(net906),
    .RESET_B(net135),
    .D(_0338_),
    .Q_N(_0039_),
    .Q(\GUScpu0.regs[2][11] ));
 sg13g2_dfrbp_1 _3785_ (.CLK(net910),
    .RESET_B(net134),
    .D(_0339_),
    .Q_N(_0047_),
    .Q(\GUScpu0.regs[2][12] ));
 sg13g2_dfrbp_1 _3786_ (.CLK(net911),
    .RESET_B(net133),
    .D(_0340_),
    .Q_N(_0055_),
    .Q(\GUScpu0.regs[2][13] ));
 sg13g2_dfrbp_1 _3787_ (.CLK(net913),
    .RESET_B(net132),
    .D(_0341_),
    .Q_N(_0063_),
    .Q(\GUScpu0.regs[2][14] ));
 sg13g2_dfrbp_1 _3788_ (.CLK(net894),
    .RESET_B(net131),
    .D(_0342_),
    .Q_N(_0071_),
    .Q(\GUScpu0.regs[2][15] ));
 sg13g2_dfrbp_1 _3789_ (.CLK(net918),
    .RESET_B(net130),
    .D(_0343_),
    .Q_N(_1764_),
    .Q(\GUScpu0.PC1[10] ));
 sg13g2_dfrbp_1 _3790_ (.CLK(net918),
    .RESET_B(net129),
    .D(_0344_),
    .Q_N(_1763_),
    .Q(\GUScpu0.PC1[11] ));
 sg13g2_dfrbp_1 _3791_ (.CLK(net918),
    .RESET_B(net128),
    .D(_0345_),
    .Q_N(_1762_),
    .Q(\GUScpu0.PC1[12] ));
 sg13g2_dfrbp_1 _3792_ (.CLK(net918),
    .RESET_B(net127),
    .D(_0346_),
    .Q_N(_1761_),
    .Q(\GUScpu0.PC1[13] ));
 sg13g2_dfrbp_1 _3793_ (.CLK(net918),
    .RESET_B(net126),
    .D(_0347_),
    .Q_N(_1760_),
    .Q(\GUScpu0.PC1[14] ));
 sg13g2_dfrbp_1 _3794_ (.CLK(net917),
    .RESET_B(net125),
    .D(_0348_),
    .Q_N(_1759_),
    .Q(\GUScpu0.PC1[15] ));
 sg13g2_dfrbp_1 _3795_ (.CLK(net903),
    .RESET_B(net124),
    .D(_0349_),
    .Q_N(_1758_),
    .Q(\GUScpu0.flag0[2] ));
 sg13g2_dfrbp_1 _3796_ (.CLK(net903),
    .RESET_B(net123),
    .D(_0350_),
    .Q_N(_1757_),
    .Q(\GUScpu0.flag0[0] ));
 sg13g2_dfrbp_1 _3797_ (.CLK(net888),
    .RESET_B(net122),
    .D(_0351_),
    .Q_N(_0142_),
    .Q(\GUScpu0.regs[7][0] ));
 sg13g2_dfrbp_1 _3798_ (.CLK(net895),
    .RESET_B(net121),
    .D(_0352_),
    .Q_N(_0133_),
    .Q(\GUScpu0.regs[7][1] ));
 sg13g2_dfrbp_1 _3799_ (.CLK(net899),
    .RESET_B(net120),
    .D(_0353_),
    .Q_N(_0125_),
    .Q(\GUScpu0.regs[7][2] ));
 sg13g2_dfrbp_1 _3800_ (.CLK(net892),
    .RESET_B(net119),
    .D(_0354_),
    .Q_N(_0117_),
    .Q(\GUScpu0.regs[7][3] ));
 sg13g2_dfrbp_1 _3801_ (.CLK(net890),
    .RESET_B(net118),
    .D(_0355_),
    .Q_N(_0109_),
    .Q(\GUScpu0.regs[7][4] ));
 sg13g2_dfrbp_1 _3802_ (.CLK(net888),
    .RESET_B(net117),
    .D(_0356_),
    .Q_N(_0098_),
    .Q(\GUScpu0.regs[7][5] ));
 sg13g2_dfrbp_1 _3803_ (.CLK(net896),
    .RESET_B(net116),
    .D(_0357_),
    .Q_N(_0150_),
    .Q(\GUScpu0.regs[7][6] ));
 sg13g2_dfrbp_1 _3804_ (.CLK(net893),
    .RESET_B(net115),
    .D(_0358_),
    .Q_N(_0158_),
    .Q(\GUScpu0.regs[7][7] ));
 sg13g2_dfrbp_1 _3805_ (.CLK(net907),
    .RESET_B(net114),
    .D(_0359_),
    .Q_N(_0166_),
    .Q(\GUScpu0.regs[7][8] ));
 sg13g2_dfrbp_1 _3806_ (.CLK(net908),
    .RESET_B(net113),
    .D(_0360_),
    .Q_N(_0028_),
    .Q(\GUScpu0.regs[7][9] ));
 sg13g2_dfrbp_1 _3807_ (.CLK(net910),
    .RESET_B(net112),
    .D(_0361_),
    .Q_N(_0036_),
    .Q(\GUScpu0.regs[7][10] ));
 sg13g2_dfrbp_1 _3808_ (.CLK(net908),
    .RESET_B(net111),
    .D(_0362_),
    .Q_N(_0044_),
    .Q(\GUScpu0.regs[7][11] ));
 sg13g2_dfrbp_1 _3809_ (.CLK(net911),
    .RESET_B(net110),
    .D(_0363_),
    .Q_N(_0052_),
    .Q(\GUScpu0.regs[7][12] ));
 sg13g2_dfrbp_1 _3810_ (.CLK(net912),
    .RESET_B(net109),
    .D(_0364_),
    .Q_N(_0060_),
    .Q(\GUScpu0.regs[7][13] ));
 sg13g2_dfrbp_1 _3811_ (.CLK(net914),
    .RESET_B(net108),
    .D(_0365_),
    .Q_N(_0068_),
    .Q(\GUScpu0.regs[7][14] ));
 sg13g2_dfrbp_1 _3812_ (.CLK(net894),
    .RESET_B(net107),
    .D(_0366_),
    .Q_N(_0076_),
    .Q(\GUScpu0.regs[7][15] ));
 sg13g2_dfrbp_1 _3813_ (.CLK(net932),
    .RESET_B(net944),
    .D(_0367_),
    .Q_N(\uart0.urxsh[1] ),
    .Q(_0182_));
 sg13g2_dfrbp_1 _3814_ (.CLK(net932),
    .RESET_B(net944),
    .D(_0368_),
    .Q_N(\uart0.urxsh[2] ),
    .Q(_0183_));
 sg13g2_dfrbp_1 _3815_ (.CLK(net932),
    .RESET_B(net946),
    .D(_0369_),
    .Q_N(\uart0.urxsh[3] ),
    .Q(_0184_));
 sg13g2_dfrbp_1 _3816_ (.CLK(net932),
    .RESET_B(net946),
    .D(_0370_),
    .Q_N(\uart0.urxsh[4] ),
    .Q(_0185_));
 sg13g2_dfrbp_1 _3817_ (.CLK(net932),
    .RESET_B(net946),
    .D(_0371_),
    .Q_N(\uart0.urxsh[5] ),
    .Q(_0186_));
 sg13g2_dfrbp_1 _3818_ (.CLK(net931),
    .RESET_B(net945),
    .D(_0372_),
    .Q_N(\uart0.urxsh[6] ),
    .Q(_0187_));
 sg13g2_dfrbp_1 _3819_ (.CLK(net931),
    .RESET_B(net945),
    .D(_0373_),
    .Q_N(\uart0.urxsh[7] ),
    .Q(_0188_));
 sg13g2_dfrbp_1 _3820_ (.CLK(net931),
    .RESET_B(net945),
    .D(_0374_),
    .Q_N(\uart0.urxsh[8] ),
    .Q(_0189_));
 sg13g2_dfrbp_1 _3821_ (.CLK(net931),
    .RESET_B(net945),
    .D(_0375_),
    .Q_N(\uart0.urxsh[9] ),
    .Q(_0190_));
 sg13g2_dfrbp_1 _3822_ (.CLK(net933),
    .RESET_B(net945),
    .D(_0013_),
    .Q_N(_1756_),
    .Q(\uart0.rxdiv[0] ));
 sg13g2_dfrbp_1 _3823_ (.CLK(net931),
    .RESET_B(net946),
    .D(_0014_),
    .Q_N(_1755_),
    .Q(\uart0.rxdiv[1] ));
 sg13g2_dfrbp_1 _3824_ (.CLK(net933),
    .RESET_B(net945),
    .D(_0015_),
    .Q_N(_1754_),
    .Q(\uart0.rxdiv[2] ));
 sg13g2_dfrbp_1 _3825_ (.CLK(net933),
    .RESET_B(net946),
    .D(_0016_),
    .Q_N(_1753_),
    .Q(\uart0.rxdiv[3] ));
 sg13g2_dfrbp_1 _3826_ (.CLK(net932),
    .RESET_B(net946),
    .D(_0017_),
    .Q_N(_1752_),
    .Q(\uart0.rxdiv[4] ));
 sg13g2_dfrbp_1 _3827_ (.CLK(net931),
    .RESET_B(net946),
    .D(_0018_),
    .Q_N(_1751_),
    .Q(\uart0.rxdiv[5] ));
 sg13g2_dfrbp_1 _3828_ (.CLK(net929),
    .RESET_B(net944),
    .D(_0376_),
    .Q_N(_1750_),
    .Q(\uart0.txbitcnt[0] ));
 sg13g2_dfrbp_1 _3829_ (.CLK(net929),
    .RESET_B(net944),
    .D(_0377_),
    .Q_N(_1749_),
    .Q(\uart0.txbitcnt[1] ));
 sg13g2_dfrbp_1 _3830_ (.CLK(net929),
    .RESET_B(net944),
    .D(_0378_),
    .Q_N(_1748_),
    .Q(\uart0.txbitcnt[2] ));
 sg13g2_dfrbp_1 _3831_ (.CLK(net929),
    .RESET_B(net944),
    .D(_0379_),
    .Q_N(_1747_),
    .Q(\uart0.txbitcnt[3] ));
 sg13g2_dfrbp_1 _3832_ (.CLK(net930),
    .RESET_B(net18),
    .D(_0380_),
    .Q_N(_1746_),
    .Q(\uart0.q[0] ));
 sg13g2_dfrbp_1 _3833_ (.CLK(net930),
    .RESET_B(net219),
    .D(_0381_),
    .Q_N(_1745_),
    .Q(\uart0.q[1] ));
 sg13g2_dfrbp_1 _3834_ (.CLK(net929),
    .RESET_B(net217),
    .D(_0382_),
    .Q_N(_1744_),
    .Q(\uart0.q[2] ));
 sg13g2_dfrbp_1 _3835_ (.CLK(net929),
    .RESET_B(net215),
    .D(_0383_),
    .Q_N(_1743_),
    .Q(\uart0.q[3] ));
 sg13g2_dfrbp_1 _3836_ (.CLK(net932),
    .RESET_B(net213),
    .D(_0384_),
    .Q_N(_1742_),
    .Q(\uart0.q[4] ));
 sg13g2_dfrbp_1 _3837_ (.CLK(net933),
    .RESET_B(net208),
    .D(_0385_),
    .Q_N(_1741_),
    .Q(\uart0.q[5] ));
 sg13g2_dfrbp_1 _3838_ (.CLK(net933),
    .RESET_B(net204),
    .D(_0386_),
    .Q_N(_1740_),
    .Q(\uart0.q[6] ));
 sg13g2_dfrbp_1 _3839_ (.CLK(net933),
    .RESET_B(net200),
    .D(_0387_),
    .Q_N(_1739_),
    .Q(\uart0.q[7] ));
 sg13g2_dfrbp_1 _3840_ (.CLK(net933),
    .RESET_B(net196),
    .D(_0388_),
    .Q_N(_1738_),
    .Q(\uart0.urxbuffer[8] ));
 sg13g2_dfrbp_1 _3841_ (.CLK(net931),
    .RESET_B(net945),
    .D(net4),
    .Q_N(_1737_),
    .Q(\uart0.rxreg[0] ));
 sg13g2_dfrbp_1 _3842_ (.CLK(net931),
    .RESET_B(net945),
    .D(\uart0.rxreg[0] ),
    .Q_N(_1736_),
    .Q(\uart0.rxreg[1] ));
 sg13g2_dfrbp_1 _3843_ (.CLK(net930),
    .RESET_B(net943),
    .D(_0389_),
    .Q_N(_0077_),
    .Q(\uart0.rxvalid ));
 sg13g2_dfrbp_1 _3844_ (.CLK(net930),
    .RESET_B(net943),
    .D(_0390_),
    .Q_N(_1735_),
    .Q(\uart0.rxoverr ));
 sg13g2_dfrbp_1 _3845_ (.CLK(net903),
    .RESET_B(net941),
    .D(_0391_),
    .Q_N(_1734_),
    .Q(\GUScpu0.PC0[0] ));
 sg13g2_dfrbp_1 _3846_ (.CLK(net916),
    .RESET_B(net937),
    .D(_0392_),
    .Q_N(_1733_),
    .Q(\GUScpu0.PC0[1] ));
 sg13g2_dfrbp_1 _3847_ (.CLK(net915),
    .RESET_B(net939),
    .D(_0393_),
    .Q_N(_1732_),
    .Q(\GUScpu0.PC0[2] ));
 sg13g2_dfrbp_1 _3848_ (.CLK(net916),
    .RESET_B(net939),
    .D(_0394_),
    .Q_N(_1731_),
    .Q(\GUScpu0.PC0[3] ));
 sg13g2_dfrbp_1 _3849_ (.CLK(net915),
    .RESET_B(net939),
    .D(_0395_),
    .Q_N(_1730_),
    .Q(\GUScpu0.PC0[4] ));
 sg13g2_dfrbp_1 _3850_ (.CLK(net915),
    .RESET_B(net941),
    .D(_0396_),
    .Q_N(_1729_),
    .Q(\GUScpu0.PC0[5] ));
 sg13g2_dfrbp_1 _3851_ (.CLK(net916),
    .RESET_B(net941),
    .D(_0397_),
    .Q_N(_1728_),
    .Q(\GUScpu0.PC0[6] ));
 sg13g2_dfrbp_1 _3852_ (.CLK(net916),
    .RESET_B(net942),
    .D(_0398_),
    .Q_N(_1727_),
    .Q(\GUScpu0.PC0[7] ));
 sg13g2_dfrbp_1 _3853_ (.CLK(net917),
    .RESET_B(net942),
    .D(_0399_),
    .Q_N(_1726_),
    .Q(\GUScpu0.PC0[8] ));
 sg13g2_dfrbp_1 _3854_ (.CLK(net919),
    .RESET_B(net942),
    .D(_0400_),
    .Q_N(_1725_),
    .Q(\GUScpu0.PC0[9] ));
 sg13g2_dfrbp_1 _3855_ (.CLK(net918),
    .RESET_B(net947),
    .D(_0401_),
    .Q_N(_1724_),
    .Q(\GUScpu0.PC0[10] ));
 sg13g2_dfrbp_1 _3856_ (.CLK(net918),
    .RESET_B(net947),
    .D(_0402_),
    .Q_N(_1723_),
    .Q(\GUScpu0.PC0[11] ));
 sg13g2_dfrbp_1 _3857_ (.CLK(net919),
    .RESET_B(net947),
    .D(_0403_),
    .Q_N(_1722_),
    .Q(\GUScpu0.PC0[12] ));
 sg13g2_dfrbp_1 _3858_ (.CLK(net918),
    .RESET_B(net942),
    .D(_0404_),
    .Q_N(_1721_),
    .Q(\GUScpu0.PC0[13] ));
 sg13g2_dfrbp_1 _3859_ (.CLK(net919),
    .RESET_B(net942),
    .D(_0405_),
    .Q_N(_1720_),
    .Q(\GUScpu0.PC0[14] ));
 sg13g2_dfrbp_1 _3860_ (.CLK(net919),
    .RESET_B(net942),
    .D(_0406_),
    .Q_N(_1719_),
    .Q(\GUScpu0.PC0[15] ));
 sg13g2_dfrbp_1 _3861_ (.CLK(net926),
    .RESET_B(net940),
    .D(_0019_),
    .Q_N(_1718_),
    .Q(\uart0.txdiv[0] ));
 sg13g2_dfrbp_1 _3862_ (.CLK(net926),
    .RESET_B(net938),
    .D(_0020_),
    .Q_N(_1717_),
    .Q(\uart0.txdiv[1] ));
 sg13g2_dfrbp_1 _3863_ (.CLK(net926),
    .RESET_B(net938),
    .D(_0021_),
    .Q_N(_1716_),
    .Q(\uart0.txdiv[2] ));
 sg13g2_dfrbp_1 _3864_ (.CLK(net926),
    .RESET_B(net938),
    .D(_0022_),
    .Q_N(_1715_),
    .Q(\uart0.txdiv[3] ));
 sg13g2_dfrbp_1 _3865_ (.CLK(net926),
    .RESET_B(net938),
    .D(_0023_),
    .Q_N(_1714_),
    .Q(\uart0.txdiv[4] ));
 sg13g2_dfrbp_1 _3866_ (.CLK(net926),
    .RESET_B(net940),
    .D(_0024_),
    .Q_N(_1713_),
    .Q(\uart0.txdiv[5] ));
 sg13g2_dfrbp_1 _3867_ (.CLK(net888),
    .RESET_B(net24),
    .D(_0407_),
    .Q_N(_0136_),
    .Q(\GUScpu0.regs[1][0] ));
 sg13g2_dfrbp_1 _3868_ (.CLK(net895),
    .RESET_B(net23),
    .D(_0408_),
    .Q_N(_0127_),
    .Q(\GUScpu0.regs[1][1] ));
 sg13g2_dfrbp_1 _3869_ (.CLK(net891),
    .RESET_B(net22),
    .D(_0409_),
    .Q_N(_0119_),
    .Q(\GUScpu0.regs[1][2] ));
 sg13g2_dfrbp_1 _3870_ (.CLK(net891),
    .RESET_B(net21),
    .D(_0410_),
    .Q_N(_0111_),
    .Q(\GUScpu0.regs[1][3] ));
 sg13g2_dfrbp_1 _3871_ (.CLK(net890),
    .RESET_B(net20),
    .D(_0411_),
    .Q_N(_0103_),
    .Q(\GUScpu0.regs[1][4] ));
 sg13g2_dfrbp_1 _3872_ (.CLK(net889),
    .RESET_B(net19),
    .D(_0412_),
    .Q_N(_0086_),
    .Q(\GUScpu0.regs[1][5] ));
 sg13g2_dfrbp_1 _3873_ (.CLK(net896),
    .RESET_B(net17),
    .D(_0413_),
    .Q_N(_0144_),
    .Q(\GUScpu0.regs[1][6] ));
 sg13g2_dfrbp_1 _3874_ (.CLK(net893),
    .RESET_B(net218),
    .D(_0414_),
    .Q_N(_0152_),
    .Q(\GUScpu0.regs[1][7] ));
 sg13g2_dfrbp_1 _3875_ (.CLK(net907),
    .RESET_B(net216),
    .D(_0415_),
    .Q_N(_0160_),
    .Q(\GUScpu0.regs[1][8] ));
 sg13g2_dfrbp_1 _3876_ (.CLK(net909),
    .RESET_B(net214),
    .D(_0416_),
    .Q_N(_0168_),
    .Q(\GUScpu0.regs[1][9] ));
 sg13g2_dfrbp_1 _3877_ (.CLK(net910),
    .RESET_B(net210),
    .D(_0417_),
    .Q_N(_0030_),
    .Q(\GUScpu0.regs[1][10] ));
 sg13g2_dfrbp_1 _3878_ (.CLK(net906),
    .RESET_B(net206),
    .D(_0418_),
    .Q_N(_0038_),
    .Q(\GUScpu0.regs[1][11] ));
 sg13g2_dfrbp_1 _3879_ (.CLK(net910),
    .RESET_B(net202),
    .D(_0419_),
    .Q_N(_0046_),
    .Q(\GUScpu0.regs[1][12] ));
 sg13g2_dfrbp_1 _3880_ (.CLK(net911),
    .RESET_B(net198),
    .D(_0420_),
    .Q_N(_0054_),
    .Q(\GUScpu0.regs[1][13] ));
 sg13g2_dfrbp_1 _3881_ (.CLK(net913),
    .RESET_B(net195),
    .D(_0421_),
    .Q_N(_0062_),
    .Q(\GUScpu0.regs[1][14] ));
 sg13g2_dfrbp_1 _3882_ (.CLK(net894),
    .RESET_B(net106),
    .D(_0422_),
    .Q_N(_0070_),
    .Q(\GUScpu0.regs[1][15] ));
 sg13g2_tiehi _3832__18 (.L_HI(net18));
 sg13g2_tiehi _3872__19 (.L_HI(net19));
 sg13g2_tiehi _3871__20 (.L_HI(net20));
 sg13g2_tiehi _3870__21 (.L_HI(net21));
 sg13g2_tiehi _3869__22 (.L_HI(net22));
 sg13g2_tiehi _3868__23 (.L_HI(net23));
 sg13g2_tiehi _3867__24 (.L_HI(net24));
 sg13g2_tiehi _3665__25 (.L_HI(net25));
 sg13g2_tiehi _3664__26 (.L_HI(net26));
 sg13g2_tiehi _3663__27 (.L_HI(net27));
 sg13g2_tiehi _3662__28 (.L_HI(net28));
 sg13g2_tiehi _3661__29 (.L_HI(net29));
 sg13g2_tiehi _3660__30 (.L_HI(net30));
 sg13g2_tiehi _3659__31 (.L_HI(net31));
 sg13g2_tiehi _3658__32 (.L_HI(net32));
 sg13g2_tiehi _3657__33 (.L_HI(net33));
 sg13g2_tiehi _3656__34 (.L_HI(net34));
 sg13g2_tiehi _3655__35 (.L_HI(net35));
 sg13g2_tiehi _3654__36 (.L_HI(net36));
 sg13g2_tiehi _3653__37 (.L_HI(net37));
 sg13g2_tiehi _3652__38 (.L_HI(net38));
 sg13g2_tiehi _3651__39 (.L_HI(net39));
 sg13g2_tiehi _3650__40 (.L_HI(net40));
 sg13g2_tiehi _3649__41 (.L_HI(net41));
 sg13g2_tiehi _3648__42 (.L_HI(net42));
 sg13g2_tiehi _3647__43 (.L_HI(net43));
 sg13g2_tiehi _3646__44 (.L_HI(net44));
 sg13g2_tiehi _3605__45 (.L_HI(net45));
 sg13g2_tiehi _3645__46 (.L_HI(net46));
 sg13g2_tiehi _3644__47 (.L_HI(net47));
 sg13g2_tiehi _3643__48 (.L_HI(net48));
 sg13g2_tiehi _3642__49 (.L_HI(net49));
 sg13g2_tiehi _3641__50 (.L_HI(net50));
 sg13g2_tiehi _3640__51 (.L_HI(net51));
 sg13g2_tiehi _3639__52 (.L_HI(net52));
 sg13g2_tiehi _3638__53 (.L_HI(net53));
 sg13g2_tiehi _3716__54 (.L_HI(net54));
 sg13g2_tiehi _3717__55 (.L_HI(net55));
 sg13g2_tiehi _3718__56 (.L_HI(net56));
 sg13g2_tiehi _3719__57 (.L_HI(net57));
 sg13g2_tiehi _3720__58 (.L_HI(net58));
 sg13g2_tiehi _3721__59 (.L_HI(net59));
 sg13g2_tiehi _3722__60 (.L_HI(net60));
 sg13g2_tiehi _3723__61 (.L_HI(net61));
 sg13g2_tiehi _3724__62 (.L_HI(net62));
 sg13g2_tiehi _3725__63 (.L_HI(net63));
 sg13g2_tiehi _3726__64 (.L_HI(net64));
 sg13g2_tiehi _3727__65 (.L_HI(net65));
 sg13g2_tiehi _3728__66 (.L_HI(net66));
 sg13g2_tiehi _3729__67 (.L_HI(net67));
 sg13g2_tiehi _3730__68 (.L_HI(net68));
 sg13g2_tiehi _3731__69 (.L_HI(net69));
 sg13g2_tiehi _3732__70 (.L_HI(net70));
 sg13g2_tiehi _3733__71 (.L_HI(net71));
 sg13g2_tiehi _3734__72 (.L_HI(net72));
 sg13g2_tiehi _3735__73 (.L_HI(net73));
 sg13g2_tiehi _3637__74 (.L_HI(net74));
 sg13g2_tiehi _3636__75 (.L_HI(net75));
 sg13g2_tiehi _3635__76 (.L_HI(net76));
 sg13g2_tiehi _3634__77 (.L_HI(net77));
 sg13g2_tiehi _3633__78 (.L_HI(net78));
 sg13g2_tiehi _3632__79 (.L_HI(net79));
 sg13g2_tiehi _3631__80 (.L_HI(net80));
 sg13g2_tiehi _3630__81 (.L_HI(net81));
 sg13g2_tiehi _3629__82 (.L_HI(net82));
 sg13g2_tiehi _3628__83 (.L_HI(net83));
 sg13g2_tiehi _3627__84 (.L_HI(net84));
 sg13g2_tiehi _3626__85 (.L_HI(net85));
 sg13g2_tiehi _3625__86 (.L_HI(net86));
 sg13g2_tiehi _3624__87 (.L_HI(net87));
 sg13g2_tiehi _3623__88 (.L_HI(net88));
 sg13g2_tiehi _3622__89 (.L_HI(net89));
 sg13g2_tiehi _3621__90 (.L_HI(net90));
 sg13g2_tiehi _3620__91 (.L_HI(net91));
 sg13g2_tiehi _3619__92 (.L_HI(net92));
 sg13g2_tiehi _3618__93 (.L_HI(net93));
 sg13g2_tiehi _3617__94 (.L_HI(net94));
 sg13g2_tiehi _3616__95 (.L_HI(net95));
 sg13g2_tiehi _3615__96 (.L_HI(net96));
 sg13g2_tiehi _3614__97 (.L_HI(net97));
 sg13g2_tiehi _3613__98 (.L_HI(net98));
 sg13g2_tiehi _3612__99 (.L_HI(net99));
 sg13g2_tiehi _3611__100 (.L_HI(net100));
 sg13g2_tiehi _3610__101 (.L_HI(net101));
 sg13g2_tiehi _3609__102 (.L_HI(net102));
 sg13g2_tiehi _3608__103 (.L_HI(net103));
 sg13g2_tiehi _3607__104 (.L_HI(net104));
 sg13g2_tiehi _3606__105 (.L_HI(net105));
 sg13g2_tiehi _3882__106 (.L_HI(net106));
 sg13g2_tiehi _3812__107 (.L_HI(net107));
 sg13g2_tiehi _3811__108 (.L_HI(net108));
 sg13g2_tiehi _3810__109 (.L_HI(net109));
 sg13g2_tiehi _3809__110 (.L_HI(net110));
 sg13g2_tiehi _3808__111 (.L_HI(net111));
 sg13g2_tiehi _3807__112 (.L_HI(net112));
 sg13g2_tiehi _3806__113 (.L_HI(net113));
 sg13g2_tiehi _3805__114 (.L_HI(net114));
 sg13g2_tiehi _3804__115 (.L_HI(net115));
 sg13g2_tiehi _3803__116 (.L_HI(net116));
 sg13g2_tiehi _3802__117 (.L_HI(net117));
 sg13g2_tiehi _3801__118 (.L_HI(net118));
 sg13g2_tiehi _3800__119 (.L_HI(net119));
 sg13g2_tiehi _3799__120 (.L_HI(net120));
 sg13g2_tiehi _3798__121 (.L_HI(net121));
 sg13g2_tiehi _3797__122 (.L_HI(net122));
 sg13g2_tiehi _3796__123 (.L_HI(net123));
 sg13g2_tiehi _3795__124 (.L_HI(net124));
 sg13g2_tiehi _3794__125 (.L_HI(net125));
 sg13g2_tiehi _3793__126 (.L_HI(net126));
 sg13g2_tiehi _3792__127 (.L_HI(net127));
 sg13g2_tiehi _3791__128 (.L_HI(net128));
 sg13g2_tiehi _3790__129 (.L_HI(net129));
 sg13g2_tiehi _3789__130 (.L_HI(net130));
 sg13g2_tiehi _3788__131 (.L_HI(net131));
 sg13g2_tiehi _3787__132 (.L_HI(net132));
 sg13g2_tiehi _3786__133 (.L_HI(net133));
 sg13g2_tiehi _3785__134 (.L_HI(net134));
 sg13g2_tiehi _3784__135 (.L_HI(net135));
 sg13g2_tiehi _3783__136 (.L_HI(net136));
 sg13g2_tiehi _3782__137 (.L_HI(net137));
 sg13g2_tiehi _3781__138 (.L_HI(net138));
 sg13g2_tiehi _3780__139 (.L_HI(net139));
 sg13g2_tiehi _3779__140 (.L_HI(net140));
 sg13g2_tiehi _3778__141 (.L_HI(net141));
 sg13g2_tiehi _3777__142 (.L_HI(net142));
 sg13g2_tiehi _3776__143 (.L_HI(net143));
 sg13g2_tiehi _3775__144 (.L_HI(net144));
 sg13g2_tiehi _3774__145 (.L_HI(net145));
 sg13g2_tiehi _3773__146 (.L_HI(net146));
 sg13g2_tiehi _3772__147 (.L_HI(net147));
 sg13g2_tiehi _3771__148 (.L_HI(net148));
 sg13g2_tiehi _3770__149 (.L_HI(net149));
 sg13g2_tiehi _3769__150 (.L_HI(net150));
 sg13g2_tiehi _3768__151 (.L_HI(net151));
 sg13g2_tiehi _3767__152 (.L_HI(net152));
 sg13g2_tiehi _3766__153 (.L_HI(net153));
 sg13g2_tiehi _3765__154 (.L_HI(net154));
 sg13g2_tiehi _3764__155 (.L_HI(net155));
 sg13g2_tiehi _3763__156 (.L_HI(net156));
 sg13g2_tiehi _3762__157 (.L_HI(net157));
 sg13g2_tiehi _3761__158 (.L_HI(net158));
 sg13g2_tiehi _3760__159 (.L_HI(net159));
 sg13g2_tiehi _3759__160 (.L_HI(net160));
 sg13g2_tiehi _3758__161 (.L_HI(net161));
 sg13g2_tiehi _3757__162 (.L_HI(net162));
 sg13g2_tiehi _3756__163 (.L_HI(net163));
 sg13g2_tiehi _3755__164 (.L_HI(net164));
 sg13g2_tiehi _3754__165 (.L_HI(net165));
 sg13g2_tiehi _3753__166 (.L_HI(net166));
 sg13g2_tiehi _3752__167 (.L_HI(net167));
 sg13g2_tiehi _3751__168 (.L_HI(net168));
 sg13g2_tiehi _3750__169 (.L_HI(net169));
 sg13g2_tiehi _3749__170 (.L_HI(net170));
 sg13g2_tiehi _3748__171 (.L_HI(net171));
 sg13g2_tiehi _3747__172 (.L_HI(net172));
 sg13g2_tiehi _3746__173 (.L_HI(net173));
 sg13g2_tiehi _3745__174 (.L_HI(net174));
 sg13g2_tiehi _3744__175 (.L_HI(net175));
 sg13g2_tiehi _3743__176 (.L_HI(net176));
 sg13g2_tiehi _3742__177 (.L_HI(net177));
 sg13g2_tiehi _3741__178 (.L_HI(net178));
 sg13g2_tiehi _3740__179 (.L_HI(net179));
 sg13g2_tiehi _3739__180 (.L_HI(net180));
 sg13g2_tiehi _3715__181 (.L_HI(net181));
 sg13g2_tiehi _3714__182 (.L_HI(net182));
 sg13g2_tiehi _3713__183 (.L_HI(net183));
 sg13g2_tiehi _3712__184 (.L_HI(net184));
 sg13g2_tiehi _3711__185 (.L_HI(net185));
 sg13g2_tiehi _3710__186 (.L_HI(net186));
 sg13g2_tiehi _3701__187 (.L_HI(net187));
 sg13g2_tiehi _3700__188 (.L_HI(net188));
 sg13g2_tiehi _3699__189 (.L_HI(net189));
 sg13g2_tiehi _3698__190 (.L_HI(net190));
 sg13g2_tiehi _3697__191 (.L_HI(net191));
 sg13g2_tiehi _3696__192 (.L_HI(net192));
 sg13g2_tiehi _3695__193 (.L_HI(net193));
 sg13g2_tiehi _3694__194 (.L_HI(net194));
 sg13g2_tiehi _3881__195 (.L_HI(net195));
 sg13g2_tiehi _3840__196 (.L_HI(net196));
 sg13g2_tiehi _3691__197 (.L_HI(net197));
 sg13g2_tiehi _3880__198 (.L_HI(net198));
 sg13g2_tiehi _3690__199 (.L_HI(net199));
 sg13g2_tiehi _3839__200 (.L_HI(net200));
 sg13g2_tiehi _3689__201 (.L_HI(net201));
 sg13g2_tiehi _3879__202 (.L_HI(net202));
 sg13g2_tiehi _3688__203 (.L_HI(net203));
 sg13g2_tiehi _3838__204 (.L_HI(net204));
 sg13g2_tiehi _3687__205 (.L_HI(net205));
 sg13g2_tiehi _3878__206 (.L_HI(net206));
 sg13g2_tiehi _3686__207 (.L_HI(net207));
 sg13g2_tiehi _3837__208 (.L_HI(net208));
 sg13g2_tiehi _3685__209 (.L_HI(net209));
 sg13g2_tiehi _3877__210 (.L_HI(net210));
 sg13g2_tiehi _3684__211 (.L_HI(net211));
 sg13g2_tiehi _3683__212 (.L_HI(net212));
 sg13g2_tiehi _3836__213 (.L_HI(net213));
 sg13g2_tiehi _3876__214 (.L_HI(net214));
 sg13g2_tiehi _3835__215 (.L_HI(net215));
 sg13g2_tiehi _3875__216 (.L_HI(net216));
 sg13g2_tiehi _3834__217 (.L_HI(net217));
 sg13g2_tiehi _3874__218 (.L_HI(net218));
 sg13g2_tiehi _3833__219 (.L_HI(net219));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_buf_1 _4086_ (.A(xoeb),
    .X(uio_oe[0]));
 sg13g2_buf_1 _4087_ (.A(xoeb),
    .X(uio_oe[1]));
 sg13g2_buf_1 _4088_ (.A(xoeb),
    .X(uio_oe[2]));
 sg13g2_buf_2 _4089_ (.A(xoeb),
    .X(uio_oe[3]));
 sg13g2_buf_2 _4090_ (.A(xoeb),
    .X(uio_oe[4]));
 sg13g2_buf_2 _4091_ (.A(xoeb),
    .X(uio_oe[5]));
 sg13g2_buf_2 _4092_ (.A(xoeb),
    .X(uio_oe[6]));
 sg13g2_buf_2 _4093_ (.A(xoeb),
    .X(uio_oe[7]));
 sg13g2_buf_1 _4094_ (.A(\ckd[0] ),
    .X(uo_out[0]));
 sg13g2_buf_1 _4095_ (.A(xlal),
    .X(uo_out[1]));
 sg13g2_buf_1 _4096_ (.A(xlah),
    .X(uo_out[2]));
 sg13g2_buf_2 _4097_ (.A(pwmout),
    .X(uo_out[3]));
 sg13g2_buf_2 _4098_ (.A(txd),
    .X(uo_out[4]));
 sg13g2_buf_2 _4099_ (.A(gpo),
    .X(uo_out[5]));
 sg13g2_buf_1 _4100_ (.A(xoeb),
    .X(uo_out[6]));
 sg13g2_buf_1 _4101_ (.A(xweb),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout715 (.A(_1383_),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(net717),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(_0904_),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(net719),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(_0877_),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(net721),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(_0947_),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(_0837_),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_0837_),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(net725),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(_0829_),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(_0965_),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(net728),
    .X(net727));
 sg13g2_buf_1 fanout728 (.A(_0981_),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(net730),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(_0961_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(net732),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(_0943_),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(_0861_),
    .X(net733));
 sg13g2_buf_1 fanout734 (.A(_0861_),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(_0852_),
    .X(net735));
 sg13g2_buf_4 fanout736 (.X(net736),
    .A(_0857_));
 sg13g2_buf_4 fanout737 (.X(net737),
    .A(net738));
 sg13g2_buf_8 fanout738 (.A(_1459_),
    .X(net738));
 sg13g2_buf_4 fanout739 (.X(net739),
    .A(net740));
 sg13g2_buf_8 fanout740 (.A(_1418_),
    .X(net740));
 sg13g2_buf_4 fanout741 (.X(net741),
    .A(net742));
 sg13g2_buf_8 fanout742 (.A(_1417_),
    .X(net742));
 sg13g2_buf_4 fanout743 (.X(net743),
    .A(_1414_));
 sg13g2_buf_4 fanout744 (.X(net744),
    .A(_1414_));
 sg13g2_buf_4 fanout745 (.X(net745),
    .A(net746));
 sg13g2_buf_4 fanout746 (.X(net746),
    .A(_1365_));
 sg13g2_buf_4 fanout747 (.X(net747),
    .A(_1327_));
 sg13g2_buf_4 fanout748 (.X(net748),
    .A(_1327_));
 sg13g2_buf_4 fanout749 (.X(net749),
    .A(net750));
 sg13g2_buf_4 fanout750 (.X(net750),
    .A(_1444_));
 sg13g2_buf_4 fanout751 (.X(net751),
    .A(net752));
 sg13g2_buf_8 fanout752 (.A(_1363_),
    .X(net752));
 sg13g2_buf_4 fanout753 (.X(net753),
    .A(_0763_));
 sg13g2_buf_4 fanout754 (.X(net754),
    .A(_0763_));
 sg13g2_buf_4 fanout755 (.X(net755),
    .A(_1556_));
 sg13g2_buf_2 fanout756 (.A(_1556_),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(_1596_),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(_1555_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(net760),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_1107_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(net762),
    .X(net761));
 sg13g2_buf_1 fanout762 (.A(net763),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(_1107_),
    .X(net763));
 sg13g2_buf_4 fanout764 (.X(net764),
    .A(net765));
 sg13g2_buf_4 fanout765 (.X(net765),
    .A(_1574_));
 sg13g2_buf_2 fanout766 (.A(net768),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(net768),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(_1551_),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(_1121_),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(_1121_),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(_1120_),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(_1120_),
    .X(net772));
 sg13g2_buf_4 fanout773 (.X(net773),
    .A(net774));
 sg13g2_buf_4 fanout774 (.X(net774),
    .A(_1602_));
 sg13g2_buf_4 fanout775 (.X(net775),
    .A(_1573_));
 sg13g2_buf_2 fanout776 (.A(_1573_),
    .X(net776));
 sg13g2_buf_4 fanout777 (.X(net777),
    .A(net780));
 sg13g2_buf_4 fanout778 (.X(net778),
    .A(net780));
 sg13g2_buf_2 fanout779 (.A(net780),
    .X(net779));
 sg13g2_buf_4 fanout780 (.X(net780),
    .A(_1570_));
 sg13g2_buf_2 fanout781 (.A(net782),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(net783),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_1569_),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(net785),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(net786),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(_1569_),
    .X(net786));
 sg13g2_buf_4 fanout787 (.X(net787),
    .A(net788));
 sg13g2_buf_4 fanout788 (.X(net788),
    .A(net789));
 sg13g2_buf_4 fanout789 (.X(net789),
    .A(net797));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(net791));
 sg13g2_buf_2 fanout791 (.A(net797),
    .X(net791));
 sg13g2_buf_4 fanout792 (.X(net792),
    .A(net797));
 sg13g2_buf_2 fanout793 (.A(net795),
    .X(net793));
 sg13g2_buf_1 fanout794 (.A(net795),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(net796),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(net797),
    .X(net796));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(_1568_));
 sg13g2_buf_4 fanout798 (.X(net798),
    .A(_1567_));
 sg13g2_buf_2 fanout799 (.A(_1567_),
    .X(net799));
 sg13g2_buf_4 fanout800 (.X(net800),
    .A(net801));
 sg13g2_buf_2 fanout801 (.A(_1567_),
    .X(net801));
 sg13g2_buf_2 fanout802 (.A(net806),
    .X(net802));
 sg13g2_buf_2 fanout803 (.A(net806),
    .X(net803));
 sg13g2_buf_2 fanout804 (.A(net806),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(net806),
    .X(net805));
 sg13g2_buf_1 fanout806 (.A(net807),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(_1139_),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(_1125_),
    .X(net808));
 sg13g2_buf_1 fanout809 (.A(_1125_),
    .X(net809));
 sg13g2_buf_4 fanout810 (.X(net810),
    .A(_1124_));
 sg13g2_buf_1 fanout811 (.A(_1124_),
    .X(net811));
 sg13g2_buf_4 fanout812 (.X(net812),
    .A(_1123_));
 sg13g2_buf_4 fanout813 (.X(net813),
    .A(_1123_));
 sg13g2_buf_2 fanout814 (.A(net815),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(net818),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(net818),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(net818),
    .X(net817));
 sg13g2_buf_1 fanout818 (.A(_1122_),
    .X(net818));
 sg13g2_buf_4 fanout819 (.X(net819),
    .A(net821));
 sg13g2_buf_4 fanout820 (.X(net820),
    .A(net821));
 sg13g2_buf_4 fanout821 (.X(net821),
    .A(_1092_));
 sg13g2_buf_4 fanout822 (.X(net822),
    .A(net823));
 sg13g2_buf_2 fanout823 (.A(_1618_),
    .X(net823));
 sg13g2_buf_2 fanout824 (.A(net825),
    .X(net824));
 sg13g2_buf_4 fanout825 (.X(net825),
    .A(_1618_));
 sg13g2_buf_4 fanout826 (.X(net826),
    .A(_1610_));
 sg13g2_buf_4 fanout827 (.X(net827),
    .A(_1610_));
 sg13g2_buf_4 fanout828 (.X(net828),
    .A(_1608_));
 sg13g2_buf_2 fanout829 (.A(_1608_),
    .X(net829));
 sg13g2_buf_4 fanout830 (.X(net830),
    .A(_1564_));
 sg13g2_buf_2 fanout831 (.A(_1564_),
    .X(net831));
 sg13g2_buf_4 fanout832 (.X(net832),
    .A(_1563_));
 sg13g2_buf_2 fanout833 (.A(_0889_),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(_0887_),
    .X(net834));
 sg13g2_buf_4 fanout835 (.X(net835),
    .A(net837));
 sg13g2_buf_2 fanout836 (.A(net837),
    .X(net836));
 sg13g2_buf_4 fanout837 (.X(net837),
    .A(_1611_));
 sg13g2_buf_4 fanout838 (.X(net838),
    .A(net839));
 sg13g2_buf_4 fanout839 (.X(net839),
    .A(_1611_));
 sg13g2_buf_4 fanout840 (.X(net840),
    .A(net841));
 sg13g2_buf_4 fanout841 (.X(net841),
    .A(net842));
 sg13g2_buf_4 fanout842 (.X(net842),
    .A(net844));
 sg13g2_buf_4 fanout843 (.X(net843),
    .A(net844));
 sg13g2_buf_2 fanout844 (.A(_1607_),
    .X(net844));
 sg13g2_buf_4 fanout845 (.X(net845),
    .A(net846));
 sg13g2_buf_4 fanout846 (.X(net846),
    .A(net847));
 sg13g2_buf_4 fanout847 (.X(net847),
    .A(_1607_));
 sg13g2_buf_2 fanout848 (.A(net850),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(net850),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(_1603_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_1603_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(net853),
    .X(net852));
 sg13g2_buf_1 fanout853 (.A(net854),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_1603_),
    .X(net854));
 sg13g2_buf_4 fanout855 (.X(net855),
    .A(_1559_));
 sg13g2_buf_4 fanout856 (.X(net856),
    .A(_1559_));
 sg13g2_buf_4 fanout857 (.X(net857),
    .A(_1518_));
 sg13g2_buf_2 fanout858 (.A(net859),
    .X(net858));
 sg13g2_buf_1 fanout859 (.A(_1518_),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(net861),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_1517_),
    .X(net861));
 sg13g2_buf_4 fanout862 (.X(net862),
    .A(net863));
 sg13g2_buf_4 fanout863 (.X(net863),
    .A(net864));
 sg13g2_buf_4 fanout864 (.X(net864),
    .A(_1560_));
 sg13g2_buf_2 fanout865 (.A(net866),
    .X(net865));
 sg13g2_buf_1 fanout866 (.A(net867),
    .X(net866));
 sg13g2_buf_4 fanout867 (.X(net867),
    .A(_1510_));
 sg13g2_buf_2 fanout868 (.A(net869),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(_0873_),
    .X(net869));
 sg13g2_buf_4 fanout870 (.X(net870),
    .A(net873));
 sg13g2_buf_1 fanout871 (.A(net873),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(net873),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(\GUScpu0.imode ),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(net875),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(\GUScpu0.imode ),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(net878),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(net878),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(\GUScpu0.imode ),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(\GUScpu0.IR[13] ),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(net881),
    .X(net880));
 sg13g2_buf_1 fanout881 (.A(\GUScpu0.IR[12] ),
    .X(net881));
 sg13g2_buf_4 fanout882 (.X(net882),
    .A(\GUScpu0.IR[11] ));
 sg13g2_buf_4 fanout883 (.X(net883),
    .A(_0093_));
 sg13g2_buf_4 fanout884 (.X(net884),
    .A(\GUScpu0.IR[1] ));
 sg13g2_buf_4 fanout885 (.X(net885),
    .A(_1206_));
 sg13g2_buf_4 fanout886 (.X(net886),
    .A(\uart0.urxsh[0] ));
 sg13g2_buf_2 fanout887 (.A(\uart0.urxsh[0] ),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(net889),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(net898),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(net892),
    .X(net890));
 sg13g2_buf_1 fanout891 (.A(net892),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(net898),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(net897),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(net897),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(net897),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(net897),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(net898),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(\GUScpu0.clk ),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(net905),
    .X(net899));
 sg13g2_buf_4 fanout900 (.X(net900),
    .A(net901));
 sg13g2_buf_2 fanout901 (.A(net905),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(net904),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(net904),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(net905),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(\GUScpu0.clk ),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(net908),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(net908),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(net921),
    .X(net908));
 sg13g2_buf_2 fanout909 (.A(net912),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(net911),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(net912),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(net914),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(net914),
    .X(net913));
 sg13g2_buf_2 fanout914 (.A(net921),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(net916),
    .X(net915));
 sg13g2_buf_4 fanout916 (.X(net916),
    .A(net917));
 sg13g2_buf_2 fanout917 (.A(net921),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(net919),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(net920),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(net921),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(\GUScpu0.clk ),
    .X(net921));
 sg13g2_buf_4 fanout922 (.X(net922),
    .A(_1207_));
 sg13g2_buf_2 fanout923 (.A(xlah),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(net925),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(net928),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(net927),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(net928),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(net934),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(net930),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(net934),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(net932),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(net933),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(net934),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(_0080_),
    .X(net934));
 sg13g2_buf_4 fanout935 (.X(net935),
    .A(\ckd[0] ));
 sg13g2_buf_4 fanout936 (.X(net936),
    .A(net937));
 sg13g2_buf_2 fanout937 (.A(net940),
    .X(net937));
 sg13g2_buf_4 fanout938 (.X(net938),
    .A(net939));
 sg13g2_buf_4 fanout939 (.X(net939),
    .A(net940));
 sg13g2_buf_2 fanout940 (.A(net941),
    .X(net940));
 sg13g2_buf_4 fanout941 (.X(net941),
    .A(rst_n));
 sg13g2_buf_4 fanout942 (.X(net942),
    .A(net947));
 sg13g2_buf_4 fanout943 (.X(net943),
    .A(net947));
 sg13g2_buf_4 fanout944 (.X(net944),
    .A(net947));
 sg13g2_buf_4 fanout945 (.X(net945),
    .A(net946));
 sg13g2_buf_4 fanout946 (.X(net946),
    .A(net947));
 sg13g2_buf_4 fanout947 (.X(net947),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_tiehi _3873__17 (.L_HI(net17));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_1_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_1_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_1_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_1_1__leaf_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(_1712_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold2 (.A(\xdi[1] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0195_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold4 (.A(\xdi[4] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold5 (.A(\xdi[3] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold6 (.A(\xdi[0] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold7 (.A(\xdi[2] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold8 (.A(\xdi[7] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold9 (.A(\xdi[5] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold10 (.A(\xdi[6] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold11 (.A(\ckd[1] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold12 (.A(\ckd[1] ),
    .X(net231));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_108 ();
 sg13g2_decap_4 FILLER_0_115 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_fill_1 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_165 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_4 FILLER_1_70 ();
 sg13g2_fill_2 FILLER_1_74 ();
 sg13g2_decap_4 FILLER_1_112 ();
 sg13g2_fill_2 FILLER_1_116 ();
 sg13g2_decap_8 FILLER_1_144 ();
 sg13g2_decap_8 FILLER_1_191 ();
 sg13g2_decap_8 FILLER_1_198 ();
 sg13g2_decap_8 FILLER_1_205 ();
 sg13g2_decap_8 FILLER_1_212 ();
 sg13g2_decap_8 FILLER_1_219 ();
 sg13g2_decap_8 FILLER_1_226 ();
 sg13g2_decap_8 FILLER_1_233 ();
 sg13g2_decap_8 FILLER_1_240 ();
 sg13g2_decap_8 FILLER_1_247 ();
 sg13g2_decap_8 FILLER_1_254 ();
 sg13g2_decap_8 FILLER_1_261 ();
 sg13g2_decap_8 FILLER_1_268 ();
 sg13g2_decap_8 FILLER_1_275 ();
 sg13g2_decap_8 FILLER_1_282 ();
 sg13g2_decap_8 FILLER_1_289 ();
 sg13g2_decap_8 FILLER_1_296 ();
 sg13g2_decap_8 FILLER_1_303 ();
 sg13g2_decap_8 FILLER_1_310 ();
 sg13g2_decap_8 FILLER_1_317 ();
 sg13g2_decap_8 FILLER_1_324 ();
 sg13g2_decap_8 FILLER_1_331 ();
 sg13g2_decap_8 FILLER_1_338 ();
 sg13g2_decap_8 FILLER_1_345 ();
 sg13g2_decap_8 FILLER_1_352 ();
 sg13g2_decap_8 FILLER_1_359 ();
 sg13g2_decap_8 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_373 ();
 sg13g2_decap_8 FILLER_1_380 ();
 sg13g2_decap_8 FILLER_1_387 ();
 sg13g2_decap_8 FILLER_1_394 ();
 sg13g2_decap_8 FILLER_1_401 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_4 FILLER_2_70 ();
 sg13g2_fill_1 FILLER_2_74 ();
 sg13g2_fill_2 FILLER_2_85 ();
 sg13g2_fill_1 FILLER_2_87 ();
 sg13g2_fill_2 FILLER_2_114 ();
 sg13g2_fill_1 FILLER_2_116 ();
 sg13g2_decap_8 FILLER_2_195 ();
 sg13g2_decap_8 FILLER_2_202 ();
 sg13g2_decap_8 FILLER_2_209 ();
 sg13g2_decap_8 FILLER_2_216 ();
 sg13g2_decap_8 FILLER_2_223 ();
 sg13g2_decap_8 FILLER_2_230 ();
 sg13g2_decap_8 FILLER_2_237 ();
 sg13g2_decap_8 FILLER_2_244 ();
 sg13g2_decap_8 FILLER_2_251 ();
 sg13g2_decap_8 FILLER_2_258 ();
 sg13g2_decap_8 FILLER_2_265 ();
 sg13g2_decap_8 FILLER_2_272 ();
 sg13g2_decap_8 FILLER_2_279 ();
 sg13g2_decap_8 FILLER_2_286 ();
 sg13g2_decap_8 FILLER_2_293 ();
 sg13g2_decap_8 FILLER_2_300 ();
 sg13g2_decap_8 FILLER_2_307 ();
 sg13g2_decap_8 FILLER_2_314 ();
 sg13g2_decap_8 FILLER_2_321 ();
 sg13g2_decap_8 FILLER_2_328 ();
 sg13g2_decap_8 FILLER_2_335 ();
 sg13g2_decap_8 FILLER_2_342 ();
 sg13g2_decap_8 FILLER_2_349 ();
 sg13g2_decap_8 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_4 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_4 FILLER_3_70 ();
 sg13g2_fill_2 FILLER_3_114 ();
 sg13g2_fill_1 FILLER_3_140 ();
 sg13g2_fill_2 FILLER_3_167 ();
 sg13g2_fill_1 FILLER_3_169 ();
 sg13g2_fill_1 FILLER_3_184 ();
 sg13g2_decap_8 FILLER_3_211 ();
 sg13g2_decap_8 FILLER_3_218 ();
 sg13g2_decap_8 FILLER_3_225 ();
 sg13g2_decap_8 FILLER_3_232 ();
 sg13g2_decap_8 FILLER_3_239 ();
 sg13g2_decap_8 FILLER_3_246 ();
 sg13g2_decap_8 FILLER_3_253 ();
 sg13g2_decap_8 FILLER_3_260 ();
 sg13g2_decap_8 FILLER_3_267 ();
 sg13g2_decap_8 FILLER_3_274 ();
 sg13g2_decap_8 FILLER_3_281 ();
 sg13g2_decap_8 FILLER_3_288 ();
 sg13g2_decap_8 FILLER_3_295 ();
 sg13g2_decap_8 FILLER_3_302 ();
 sg13g2_decap_8 FILLER_3_309 ();
 sg13g2_decap_8 FILLER_3_316 ();
 sg13g2_decap_8 FILLER_3_323 ();
 sg13g2_decap_8 FILLER_3_330 ();
 sg13g2_decap_8 FILLER_3_337 ();
 sg13g2_decap_8 FILLER_3_344 ();
 sg13g2_decap_8 FILLER_3_351 ();
 sg13g2_decap_8 FILLER_3_358 ();
 sg13g2_decap_8 FILLER_3_365 ();
 sg13g2_decap_8 FILLER_3_372 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_3_386 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_decap_8 FILLER_3_400 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_fill_2 FILLER_4_63 ();
 sg13g2_decap_4 FILLER_4_95 ();
 sg13g2_decap_8 FILLER_4_103 ();
 sg13g2_decap_4 FILLER_4_110 ();
 sg13g2_fill_1 FILLER_4_114 ();
 sg13g2_decap_8 FILLER_4_141 ();
 sg13g2_decap_4 FILLER_4_148 ();
 sg13g2_fill_2 FILLER_4_152 ();
 sg13g2_decap_8 FILLER_4_162 ();
 sg13g2_decap_4 FILLER_4_169 ();
 sg13g2_fill_1 FILLER_4_173 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_4 FILLER_5_49 ();
 sg13g2_fill_1 FILLER_5_53 ();
 sg13g2_fill_1 FILLER_5_88 ();
 sg13g2_decap_8 FILLER_5_103 ();
 sg13g2_decap_4 FILLER_5_110 ();
 sg13g2_fill_2 FILLER_5_114 ();
 sg13g2_decap_8 FILLER_5_130 ();
 sg13g2_decap_8 FILLER_5_137 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_decap_4 FILLER_5_155 ();
 sg13g2_decap_8 FILLER_5_169 ();
 sg13g2_decap_4 FILLER_5_176 ();
 sg13g2_decap_4 FILLER_5_190 ();
 sg13g2_decap_8 FILLER_5_202 ();
 sg13g2_decap_8 FILLER_5_209 ();
 sg13g2_decap_8 FILLER_5_216 ();
 sg13g2_decap_8 FILLER_5_223 ();
 sg13g2_decap_8 FILLER_5_230 ();
 sg13g2_decap_8 FILLER_5_237 ();
 sg13g2_decap_8 FILLER_5_244 ();
 sg13g2_decap_8 FILLER_5_251 ();
 sg13g2_decap_8 FILLER_5_258 ();
 sg13g2_decap_8 FILLER_5_265 ();
 sg13g2_decap_8 FILLER_5_272 ();
 sg13g2_decap_8 FILLER_5_279 ();
 sg13g2_decap_8 FILLER_5_286 ();
 sg13g2_decap_8 FILLER_5_293 ();
 sg13g2_decap_8 FILLER_5_300 ();
 sg13g2_decap_8 FILLER_5_307 ();
 sg13g2_decap_8 FILLER_5_314 ();
 sg13g2_decap_8 FILLER_5_321 ();
 sg13g2_decap_8 FILLER_5_328 ();
 sg13g2_decap_8 FILLER_5_335 ();
 sg13g2_decap_8 FILLER_5_342 ();
 sg13g2_decap_8 FILLER_5_349 ();
 sg13g2_decap_8 FILLER_5_356 ();
 sg13g2_decap_8 FILLER_5_363 ();
 sg13g2_decap_8 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_decap_8 FILLER_5_384 ();
 sg13g2_decap_8 FILLER_5_391 ();
 sg13g2_decap_8 FILLER_5_398 ();
 sg13g2_decap_4 FILLER_5_405 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_4 FILLER_6_63 ();
 sg13g2_fill_1 FILLER_6_67 ();
 sg13g2_decap_4 FILLER_6_78 ();
 sg13g2_fill_1 FILLER_6_82 ();
 sg13g2_decap_4 FILLER_6_109 ();
 sg13g2_fill_1 FILLER_6_113 ();
 sg13g2_decap_4 FILLER_6_140 ();
 sg13g2_fill_2 FILLER_6_144 ();
 sg13g2_decap_8 FILLER_6_176 ();
 sg13g2_decap_8 FILLER_6_183 ();
 sg13g2_fill_2 FILLER_6_190 ();
 sg13g2_fill_1 FILLER_6_192 ();
 sg13g2_decap_8 FILLER_6_197 ();
 sg13g2_decap_8 FILLER_6_204 ();
 sg13g2_decap_8 FILLER_6_211 ();
 sg13g2_decap_8 FILLER_6_218 ();
 sg13g2_decap_8 FILLER_6_225 ();
 sg13g2_decap_8 FILLER_6_232 ();
 sg13g2_decap_8 FILLER_6_239 ();
 sg13g2_decap_8 FILLER_6_246 ();
 sg13g2_decap_8 FILLER_6_253 ();
 sg13g2_decap_8 FILLER_6_260 ();
 sg13g2_decap_8 FILLER_6_267 ();
 sg13g2_decap_8 FILLER_6_274 ();
 sg13g2_decap_8 FILLER_6_281 ();
 sg13g2_decap_8 FILLER_6_288 ();
 sg13g2_decap_8 FILLER_6_295 ();
 sg13g2_decap_8 FILLER_6_302 ();
 sg13g2_decap_8 FILLER_6_309 ();
 sg13g2_decap_8 FILLER_6_316 ();
 sg13g2_decap_8 FILLER_6_323 ();
 sg13g2_decap_8 FILLER_6_330 ();
 sg13g2_decap_8 FILLER_6_337 ();
 sg13g2_decap_8 FILLER_6_344 ();
 sg13g2_decap_8 FILLER_6_351 ();
 sg13g2_decap_8 FILLER_6_358 ();
 sg13g2_decap_8 FILLER_6_365 ();
 sg13g2_decap_8 FILLER_6_372 ();
 sg13g2_decap_8 FILLER_6_379 ();
 sg13g2_decap_8 FILLER_6_386 ();
 sg13g2_decap_8 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_400 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_fill_2 FILLER_7_45 ();
 sg13g2_decap_8 FILLER_7_51 ();
 sg13g2_decap_8 FILLER_7_58 ();
 sg13g2_fill_2 FILLER_7_65 ();
 sg13g2_fill_1 FILLER_7_67 ();
 sg13g2_fill_2 FILLER_7_72 ();
 sg13g2_fill_1 FILLER_7_74 ();
 sg13g2_decap_8 FILLER_7_80 ();
 sg13g2_decap_8 FILLER_7_87 ();
 sg13g2_decap_4 FILLER_7_120 ();
 sg13g2_fill_1 FILLER_7_124 ();
 sg13g2_fill_2 FILLER_7_184 ();
 sg13g2_fill_1 FILLER_7_186 ();
 sg13g2_decap_8 FILLER_7_208 ();
 sg13g2_decap_8 FILLER_7_215 ();
 sg13g2_decap_8 FILLER_7_222 ();
 sg13g2_decap_8 FILLER_7_229 ();
 sg13g2_decap_8 FILLER_7_236 ();
 sg13g2_decap_8 FILLER_7_243 ();
 sg13g2_decap_8 FILLER_7_250 ();
 sg13g2_decap_8 FILLER_7_257 ();
 sg13g2_decap_8 FILLER_7_264 ();
 sg13g2_decap_8 FILLER_7_271 ();
 sg13g2_decap_8 FILLER_7_278 ();
 sg13g2_decap_8 FILLER_7_285 ();
 sg13g2_decap_8 FILLER_7_292 ();
 sg13g2_decap_8 FILLER_7_299 ();
 sg13g2_decap_8 FILLER_7_306 ();
 sg13g2_decap_8 FILLER_7_313 ();
 sg13g2_decap_8 FILLER_7_320 ();
 sg13g2_decap_8 FILLER_7_327 ();
 sg13g2_decap_8 FILLER_7_334 ();
 sg13g2_decap_8 FILLER_7_341 ();
 sg13g2_decap_8 FILLER_7_348 ();
 sg13g2_decap_8 FILLER_7_355 ();
 sg13g2_decap_8 FILLER_7_362 ();
 sg13g2_decap_8 FILLER_7_369 ();
 sg13g2_decap_8 FILLER_7_376 ();
 sg13g2_decap_8 FILLER_7_383 ();
 sg13g2_decap_8 FILLER_7_390 ();
 sg13g2_decap_8 FILLER_7_397 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_4 FILLER_8_28 ();
 sg13g2_fill_1 FILLER_8_94 ();
 sg13g2_decap_8 FILLER_8_124 ();
 sg13g2_fill_1 FILLER_8_131 ();
 sg13g2_fill_2 FILLER_8_155 ();
 sg13g2_decap_8 FILLER_8_213 ();
 sg13g2_decap_8 FILLER_8_220 ();
 sg13g2_decap_8 FILLER_8_227 ();
 sg13g2_decap_8 FILLER_8_234 ();
 sg13g2_decap_8 FILLER_8_241 ();
 sg13g2_decap_8 FILLER_8_248 ();
 sg13g2_decap_8 FILLER_8_255 ();
 sg13g2_decap_8 FILLER_8_262 ();
 sg13g2_decap_8 FILLER_8_269 ();
 sg13g2_decap_8 FILLER_8_276 ();
 sg13g2_decap_8 FILLER_8_283 ();
 sg13g2_decap_8 FILLER_8_290 ();
 sg13g2_decap_8 FILLER_8_297 ();
 sg13g2_decap_8 FILLER_8_304 ();
 sg13g2_decap_8 FILLER_8_311 ();
 sg13g2_decap_8 FILLER_8_318 ();
 sg13g2_decap_8 FILLER_8_325 ();
 sg13g2_decap_8 FILLER_8_332 ();
 sg13g2_decap_8 FILLER_8_339 ();
 sg13g2_decap_8 FILLER_8_346 ();
 sg13g2_decap_8 FILLER_8_353 ();
 sg13g2_decap_8 FILLER_8_360 ();
 sg13g2_decap_8 FILLER_8_367 ();
 sg13g2_decap_8 FILLER_8_374 ();
 sg13g2_decap_8 FILLER_8_381 ();
 sg13g2_decap_8 FILLER_8_388 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_fill_1 FILLER_9_105 ();
 sg13g2_fill_2 FILLER_9_111 ();
 sg13g2_fill_1 FILLER_9_113 ();
 sg13g2_decap_4 FILLER_9_136 ();
 sg13g2_fill_2 FILLER_9_159 ();
 sg13g2_fill_1 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_fill_1 FILLER_10_35 ();
 sg13g2_fill_1 FILLER_10_80 ();
 sg13g2_decap_8 FILLER_10_107 ();
 sg13g2_decap_4 FILLER_10_114 ();
 sg13g2_fill_1 FILLER_10_118 ();
 sg13g2_decap_4 FILLER_10_145 ();
 sg13g2_fill_2 FILLER_10_149 ();
 sg13g2_decap_8 FILLER_10_177 ();
 sg13g2_decap_8 FILLER_10_184 ();
 sg13g2_fill_2 FILLER_10_191 ();
 sg13g2_decap_8 FILLER_10_198 ();
 sg13g2_decap_8 FILLER_10_205 ();
 sg13g2_decap_8 FILLER_10_212 ();
 sg13g2_decap_8 FILLER_10_219 ();
 sg13g2_decap_8 FILLER_10_226 ();
 sg13g2_decap_8 FILLER_10_233 ();
 sg13g2_decap_8 FILLER_10_240 ();
 sg13g2_decap_8 FILLER_10_247 ();
 sg13g2_decap_8 FILLER_10_254 ();
 sg13g2_decap_8 FILLER_10_261 ();
 sg13g2_decap_8 FILLER_10_268 ();
 sg13g2_decap_8 FILLER_10_275 ();
 sg13g2_decap_8 FILLER_10_282 ();
 sg13g2_decap_8 FILLER_10_289 ();
 sg13g2_decap_8 FILLER_10_296 ();
 sg13g2_decap_8 FILLER_10_303 ();
 sg13g2_decap_8 FILLER_10_310 ();
 sg13g2_decap_8 FILLER_10_317 ();
 sg13g2_decap_8 FILLER_10_324 ();
 sg13g2_decap_8 FILLER_10_331 ();
 sg13g2_decap_8 FILLER_10_338 ();
 sg13g2_decap_8 FILLER_10_345 ();
 sg13g2_decap_8 FILLER_10_352 ();
 sg13g2_decap_8 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_366 ();
 sg13g2_decap_8 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_8 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_fill_2 FILLER_11_42 ();
 sg13g2_fill_1 FILLER_11_44 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_fill_2 FILLER_11_56 ();
 sg13g2_fill_1 FILLER_11_58 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_fill_1 FILLER_11_82 ();
 sg13g2_decap_4 FILLER_11_87 ();
 sg13g2_fill_1 FILLER_11_91 ();
 sg13g2_decap_4 FILLER_11_96 ();
 sg13g2_decap_8 FILLER_11_113 ();
 sg13g2_decap_8 FILLER_11_149 ();
 sg13g2_decap_4 FILLER_11_156 ();
 sg13g2_fill_1 FILLER_11_160 ();
 sg13g2_decap_8 FILLER_11_165 ();
 sg13g2_decap_4 FILLER_11_172 ();
 sg13g2_fill_1 FILLER_11_176 ();
 sg13g2_decap_8 FILLER_11_185 ();
 sg13g2_fill_2 FILLER_11_192 ();
 sg13g2_decap_8 FILLER_11_198 ();
 sg13g2_decap_8 FILLER_11_205 ();
 sg13g2_decap_8 FILLER_11_212 ();
 sg13g2_decap_8 FILLER_11_219 ();
 sg13g2_decap_8 FILLER_11_226 ();
 sg13g2_decap_8 FILLER_11_233 ();
 sg13g2_decap_8 FILLER_11_240 ();
 sg13g2_decap_8 FILLER_11_247 ();
 sg13g2_decap_8 FILLER_11_254 ();
 sg13g2_decap_8 FILLER_11_261 ();
 sg13g2_decap_8 FILLER_11_268 ();
 sg13g2_decap_8 FILLER_11_275 ();
 sg13g2_decap_8 FILLER_11_282 ();
 sg13g2_decap_8 FILLER_11_289 ();
 sg13g2_decap_8 FILLER_11_296 ();
 sg13g2_decap_8 FILLER_11_303 ();
 sg13g2_decap_8 FILLER_11_310 ();
 sg13g2_decap_8 FILLER_11_317 ();
 sg13g2_decap_8 FILLER_11_324 ();
 sg13g2_decap_8 FILLER_11_331 ();
 sg13g2_decap_8 FILLER_11_338 ();
 sg13g2_decap_8 FILLER_11_345 ();
 sg13g2_decap_8 FILLER_11_352 ();
 sg13g2_decap_8 FILLER_11_359 ();
 sg13g2_decap_8 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_4 FILLER_12_42 ();
 sg13g2_fill_1 FILLER_12_46 ();
 sg13g2_decap_8 FILLER_12_51 ();
 sg13g2_fill_2 FILLER_12_58 ();
 sg13g2_fill_1 FILLER_12_60 ();
 sg13g2_fill_2 FILLER_12_82 ();
 sg13g2_fill_2 FILLER_12_97 ();
 sg13g2_decap_4 FILLER_12_119 ();
 sg13g2_decap_4 FILLER_12_137 ();
 sg13g2_fill_1 FILLER_12_141 ();
 sg13g2_decap_4 FILLER_12_160 ();
 sg13g2_fill_2 FILLER_12_183 ();
 sg13g2_decap_8 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_256 ();
 sg13g2_decap_8 FILLER_12_263 ();
 sg13g2_decap_8 FILLER_12_270 ();
 sg13g2_decap_8 FILLER_12_277 ();
 sg13g2_decap_8 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_fill_1 FILLER_13_35 ();
 sg13g2_fill_2 FILLER_13_99 ();
 sg13g2_fill_2 FILLER_13_113 ();
 sg13g2_decap_4 FILLER_13_120 ();
 sg13g2_fill_1 FILLER_13_134 ();
 sg13g2_fill_1 FILLER_13_155 ();
 sg13g2_fill_1 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_221 ();
 sg13g2_decap_8 FILLER_13_228 ();
 sg13g2_decap_8 FILLER_13_235 ();
 sg13g2_decap_8 FILLER_13_242 ();
 sg13g2_decap_8 FILLER_13_249 ();
 sg13g2_decap_8 FILLER_13_256 ();
 sg13g2_decap_8 FILLER_13_263 ();
 sg13g2_decap_8 FILLER_13_270 ();
 sg13g2_decap_8 FILLER_13_277 ();
 sg13g2_decap_8 FILLER_13_284 ();
 sg13g2_decap_8 FILLER_13_291 ();
 sg13g2_decap_8 FILLER_13_298 ();
 sg13g2_decap_8 FILLER_13_305 ();
 sg13g2_decap_8 FILLER_13_312 ();
 sg13g2_decap_8 FILLER_13_319 ();
 sg13g2_decap_8 FILLER_13_326 ();
 sg13g2_decap_8 FILLER_13_333 ();
 sg13g2_decap_8 FILLER_13_340 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_361 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_4 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_fill_1 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_49 ();
 sg13g2_fill_1 FILLER_14_116 ();
 sg13g2_fill_2 FILLER_14_186 ();
 sg13g2_decap_8 FILLER_14_213 ();
 sg13g2_decap_8 FILLER_14_220 ();
 sg13g2_decap_8 FILLER_14_227 ();
 sg13g2_decap_8 FILLER_14_234 ();
 sg13g2_decap_8 FILLER_14_241 ();
 sg13g2_decap_8 FILLER_14_248 ();
 sg13g2_decap_8 FILLER_14_255 ();
 sg13g2_decap_8 FILLER_14_262 ();
 sg13g2_decap_8 FILLER_14_269 ();
 sg13g2_decap_8 FILLER_14_276 ();
 sg13g2_decap_8 FILLER_14_283 ();
 sg13g2_decap_8 FILLER_14_290 ();
 sg13g2_decap_8 FILLER_14_297 ();
 sg13g2_decap_8 FILLER_14_304 ();
 sg13g2_decap_8 FILLER_14_311 ();
 sg13g2_decap_8 FILLER_14_318 ();
 sg13g2_decap_8 FILLER_14_325 ();
 sg13g2_decap_8 FILLER_14_332 ();
 sg13g2_decap_8 FILLER_14_339 ();
 sg13g2_decap_8 FILLER_14_346 ();
 sg13g2_decap_8 FILLER_14_353 ();
 sg13g2_decap_8 FILLER_14_360 ();
 sg13g2_decap_8 FILLER_14_367 ();
 sg13g2_decap_8 FILLER_14_374 ();
 sg13g2_decap_8 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_14_388 ();
 sg13g2_decap_8 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_4 FILLER_15_28 ();
 sg13g2_fill_1 FILLER_15_32 ();
 sg13g2_decap_8 FILLER_15_73 ();
 sg13g2_fill_1 FILLER_15_80 ();
 sg13g2_fill_1 FILLER_15_96 ();
 sg13g2_fill_2 FILLER_15_101 ();
 sg13g2_fill_1 FILLER_15_103 ();
 sg13g2_decap_4 FILLER_15_144 ();
 sg13g2_fill_1 FILLER_15_148 ();
 sg13g2_decap_8 FILLER_15_157 ();
 sg13g2_decap_4 FILLER_15_164 ();
 sg13g2_fill_2 FILLER_15_168 ();
 sg13g2_decap_4 FILLER_15_183 ();
 sg13g2_fill_2 FILLER_15_187 ();
 sg13g2_decap_8 FILLER_15_205 ();
 sg13g2_decap_8 FILLER_15_212 ();
 sg13g2_decap_8 FILLER_15_219 ();
 sg13g2_decap_8 FILLER_15_226 ();
 sg13g2_decap_8 FILLER_15_233 ();
 sg13g2_decap_8 FILLER_15_240 ();
 sg13g2_decap_8 FILLER_15_247 ();
 sg13g2_decap_8 FILLER_15_254 ();
 sg13g2_decap_8 FILLER_15_261 ();
 sg13g2_decap_8 FILLER_15_268 ();
 sg13g2_decap_8 FILLER_15_275 ();
 sg13g2_decap_8 FILLER_15_282 ();
 sg13g2_decap_8 FILLER_15_289 ();
 sg13g2_decap_8 FILLER_15_296 ();
 sg13g2_decap_8 FILLER_15_303 ();
 sg13g2_decap_8 FILLER_15_310 ();
 sg13g2_decap_8 FILLER_15_317 ();
 sg13g2_decap_8 FILLER_15_324 ();
 sg13g2_decap_8 FILLER_15_331 ();
 sg13g2_decap_8 FILLER_15_338 ();
 sg13g2_decap_8 FILLER_15_345 ();
 sg13g2_decap_8 FILLER_15_352 ();
 sg13g2_decap_8 FILLER_15_359 ();
 sg13g2_decap_8 FILLER_15_366 ();
 sg13g2_decap_8 FILLER_15_373 ();
 sg13g2_decap_8 FILLER_15_380 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_fill_2 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_48 ();
 sg13g2_decap_8 FILLER_16_55 ();
 sg13g2_decap_8 FILLER_16_62 ();
 sg13g2_decap_8 FILLER_16_69 ();
 sg13g2_decap_8 FILLER_16_76 ();
 sg13g2_decap_4 FILLER_16_83 ();
 sg13g2_fill_1 FILLER_16_113 ();
 sg13g2_decap_4 FILLER_16_122 ();
 sg13g2_fill_2 FILLER_16_152 ();
 sg13g2_fill_1 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_165 ();
 sg13g2_decap_4 FILLER_16_185 ();
 sg13g2_fill_1 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_205 ();
 sg13g2_decap_8 FILLER_16_212 ();
 sg13g2_decap_8 FILLER_16_219 ();
 sg13g2_decap_8 FILLER_16_226 ();
 sg13g2_decap_8 FILLER_16_233 ();
 sg13g2_decap_8 FILLER_16_240 ();
 sg13g2_decap_8 FILLER_16_247 ();
 sg13g2_decap_8 FILLER_16_254 ();
 sg13g2_decap_8 FILLER_16_261 ();
 sg13g2_decap_8 FILLER_16_268 ();
 sg13g2_decap_8 FILLER_16_275 ();
 sg13g2_decap_8 FILLER_16_282 ();
 sg13g2_decap_8 FILLER_16_289 ();
 sg13g2_decap_8 FILLER_16_296 ();
 sg13g2_decap_8 FILLER_16_303 ();
 sg13g2_decap_8 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_317 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_decap_8 FILLER_16_331 ();
 sg13g2_decap_8 FILLER_16_338 ();
 sg13g2_decap_8 FILLER_16_345 ();
 sg13g2_decap_8 FILLER_16_352 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_fill_2 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_40 ();
 sg13g2_decap_8 FILLER_17_47 ();
 sg13g2_fill_2 FILLER_17_54 ();
 sg13g2_decap_8 FILLER_17_82 ();
 sg13g2_decap_8 FILLER_17_89 ();
 sg13g2_decap_8 FILLER_17_96 ();
 sg13g2_decap_8 FILLER_17_103 ();
 sg13g2_decap_8 FILLER_17_110 ();
 sg13g2_decap_8 FILLER_17_117 ();
 sg13g2_decap_8 FILLER_17_124 ();
 sg13g2_fill_1 FILLER_17_136 ();
 sg13g2_decap_8 FILLER_17_141 ();
 sg13g2_decap_4 FILLER_17_148 ();
 sg13g2_decap_8 FILLER_17_214 ();
 sg13g2_decap_4 FILLER_17_221 ();
 sg13g2_decap_8 FILLER_17_240 ();
 sg13g2_decap_8 FILLER_17_247 ();
 sg13g2_decap_8 FILLER_17_254 ();
 sg13g2_decap_8 FILLER_17_261 ();
 sg13g2_decap_8 FILLER_17_268 ();
 sg13g2_decap_8 FILLER_17_275 ();
 sg13g2_decap_8 FILLER_17_282 ();
 sg13g2_decap_8 FILLER_17_289 ();
 sg13g2_decap_8 FILLER_17_296 ();
 sg13g2_decap_8 FILLER_17_303 ();
 sg13g2_decap_8 FILLER_17_310 ();
 sg13g2_decap_8 FILLER_17_317 ();
 sg13g2_decap_8 FILLER_17_324 ();
 sg13g2_decap_8 FILLER_17_331 ();
 sg13g2_decap_8 FILLER_17_338 ();
 sg13g2_decap_8 FILLER_17_345 ();
 sg13g2_decap_8 FILLER_17_352 ();
 sg13g2_decap_8 FILLER_17_359 ();
 sg13g2_decap_8 FILLER_17_366 ();
 sg13g2_decap_8 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_23 ();
 sg13g2_fill_1 FILLER_18_54 ();
 sg13g2_decap_8 FILLER_18_94 ();
 sg13g2_fill_1 FILLER_18_101 ();
 sg13g2_decap_4 FILLER_18_110 ();
 sg13g2_decap_8 FILLER_18_127 ();
 sg13g2_decap_8 FILLER_18_134 ();
 sg13g2_decap_8 FILLER_18_141 ();
 sg13g2_fill_2 FILLER_18_148 ();
 sg13g2_fill_1 FILLER_18_150 ();
 sg13g2_fill_2 FILLER_18_191 ();
 sg13g2_fill_2 FILLER_18_197 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_fill_2 FILLER_18_217 ();
 sg13g2_fill_2 FILLER_18_229 ();
 sg13g2_fill_1 FILLER_18_231 ();
 sg13g2_fill_2 FILLER_18_243 ();
 sg13g2_fill_1 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_250 ();
 sg13g2_decap_8 FILLER_18_257 ();
 sg13g2_decap_8 FILLER_18_264 ();
 sg13g2_decap_8 FILLER_18_271 ();
 sg13g2_decap_8 FILLER_18_278 ();
 sg13g2_decap_8 FILLER_18_285 ();
 sg13g2_decap_8 FILLER_18_292 ();
 sg13g2_decap_8 FILLER_18_299 ();
 sg13g2_decap_8 FILLER_18_306 ();
 sg13g2_decap_8 FILLER_18_313 ();
 sg13g2_decap_8 FILLER_18_320 ();
 sg13g2_decap_8 FILLER_18_327 ();
 sg13g2_decap_8 FILLER_18_334 ();
 sg13g2_decap_8 FILLER_18_341 ();
 sg13g2_decap_8 FILLER_18_348 ();
 sg13g2_decap_8 FILLER_18_355 ();
 sg13g2_decap_8 FILLER_18_362 ();
 sg13g2_decap_8 FILLER_18_369 ();
 sg13g2_decap_8 FILLER_18_376 ();
 sg13g2_decap_8 FILLER_18_383 ();
 sg13g2_decap_8 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_397 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_4 FILLER_19_14 ();
 sg13g2_fill_2 FILLER_19_78 ();
 sg13g2_decap_4 FILLER_19_151 ();
 sg13g2_fill_2 FILLER_19_155 ();
 sg13g2_fill_1 FILLER_19_171 ();
 sg13g2_fill_2 FILLER_19_229 ();
 sg13g2_fill_2 FILLER_19_237 ();
 sg13g2_decap_8 FILLER_19_260 ();
 sg13g2_decap_8 FILLER_19_267 ();
 sg13g2_decap_8 FILLER_19_274 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_decap_8 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_decap_8 FILLER_19_302 ();
 sg13g2_decap_8 FILLER_19_309 ();
 sg13g2_decap_8 FILLER_19_316 ();
 sg13g2_decap_8 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_330 ();
 sg13g2_decap_8 FILLER_19_337 ();
 sg13g2_decap_8 FILLER_19_344 ();
 sg13g2_decap_8 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_fill_2 FILLER_20_21 ();
 sg13g2_fill_1 FILLER_20_23 ();
 sg13g2_decap_8 FILLER_20_50 ();
 sg13g2_decap_8 FILLER_20_57 ();
 sg13g2_fill_2 FILLER_20_64 ();
 sg13g2_fill_1 FILLER_20_66 ();
 sg13g2_fill_2 FILLER_20_71 ();
 sg13g2_fill_1 FILLER_20_79 ();
 sg13g2_fill_2 FILLER_20_105 ();
 sg13g2_fill_2 FILLER_20_126 ();
 sg13g2_decap_4 FILLER_20_164 ();
 sg13g2_fill_1 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_194 ();
 sg13g2_fill_1 FILLER_20_201 ();
 sg13g2_fill_1 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_269 ();
 sg13g2_decap_8 FILLER_20_276 ();
 sg13g2_decap_8 FILLER_20_283 ();
 sg13g2_decap_8 FILLER_20_290 ();
 sg13g2_decap_8 FILLER_20_297 ();
 sg13g2_decap_8 FILLER_20_304 ();
 sg13g2_decap_8 FILLER_20_311 ();
 sg13g2_decap_8 FILLER_20_318 ();
 sg13g2_decap_8 FILLER_20_325 ();
 sg13g2_decap_8 FILLER_20_332 ();
 sg13g2_decap_8 FILLER_20_339 ();
 sg13g2_decap_8 FILLER_20_346 ();
 sg13g2_decap_8 FILLER_20_353 ();
 sg13g2_decap_8 FILLER_20_360 ();
 sg13g2_decap_8 FILLER_20_367 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_decap_8 FILLER_20_381 ();
 sg13g2_decap_8 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_43 ();
 sg13g2_fill_2 FILLER_21_50 ();
 sg13g2_fill_2 FILLER_21_62 ();
 sg13g2_fill_1 FILLER_21_85 ();
 sg13g2_fill_1 FILLER_21_125 ();
 sg13g2_fill_2 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_4 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_204 ();
 sg13g2_decap_8 FILLER_21_258 ();
 sg13g2_fill_1 FILLER_21_265 ();
 sg13g2_decap_8 FILLER_21_292 ();
 sg13g2_decap_8 FILLER_21_299 ();
 sg13g2_decap_8 FILLER_21_306 ();
 sg13g2_decap_8 FILLER_21_313 ();
 sg13g2_decap_8 FILLER_21_320 ();
 sg13g2_decap_8 FILLER_21_327 ();
 sg13g2_decap_8 FILLER_21_334 ();
 sg13g2_decap_8 FILLER_21_341 ();
 sg13g2_decap_8 FILLER_21_348 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_21_383 ();
 sg13g2_decap_8 FILLER_21_390 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_4 FILLER_22_42 ();
 sg13g2_fill_2 FILLER_22_46 ();
 sg13g2_fill_2 FILLER_22_89 ();
 sg13g2_decap_4 FILLER_22_107 ();
 sg13g2_fill_2 FILLER_22_111 ();
 sg13g2_decap_4 FILLER_22_137 ();
 sg13g2_fill_2 FILLER_22_141 ();
 sg13g2_fill_1 FILLER_22_153 ();
 sg13g2_decap_8 FILLER_22_162 ();
 sg13g2_fill_2 FILLER_22_169 ();
 sg13g2_fill_1 FILLER_22_171 ();
 sg13g2_decap_8 FILLER_22_180 ();
 sg13g2_decap_8 FILLER_22_187 ();
 sg13g2_fill_1 FILLER_22_194 ();
 sg13g2_decap_8 FILLER_22_200 ();
 sg13g2_decap_8 FILLER_22_207 ();
 sg13g2_decap_4 FILLER_22_214 ();
 sg13g2_fill_2 FILLER_22_218 ();
 sg13g2_fill_2 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_fill_2 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_291 ();
 sg13g2_decap_8 FILLER_22_298 ();
 sg13g2_decap_8 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_312 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_decap_8 FILLER_22_326 ();
 sg13g2_decap_8 FILLER_22_333 ();
 sg13g2_decap_8 FILLER_22_340 ();
 sg13g2_decap_8 FILLER_22_347 ();
 sg13g2_decap_8 FILLER_22_354 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_fill_2 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_30 ();
 sg13g2_decap_4 FILLER_23_65 ();
 sg13g2_fill_1 FILLER_23_69 ();
 sg13g2_fill_2 FILLER_23_88 ();
 sg13g2_fill_1 FILLER_23_90 ();
 sg13g2_decap_4 FILLER_23_134 ();
 sg13g2_fill_2 FILLER_23_138 ();
 sg13g2_fill_2 FILLER_23_150 ();
 sg13g2_fill_2 FILLER_23_156 ();
 sg13g2_decap_4 FILLER_23_163 ();
 sg13g2_fill_1 FILLER_23_167 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_fill_2 FILLER_23_201 ();
 sg13g2_fill_1 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_225 ();
 sg13g2_fill_1 FILLER_23_231 ();
 sg13g2_decap_4 FILLER_23_236 ();
 sg13g2_fill_1 FILLER_23_240 ();
 sg13g2_decap_4 FILLER_23_254 ();
 sg13g2_fill_2 FILLER_23_258 ();
 sg13g2_fill_2 FILLER_23_284 ();
 sg13g2_decap_8 FILLER_23_312 ();
 sg13g2_decap_8 FILLER_23_319 ();
 sg13g2_decap_8 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_347 ();
 sg13g2_decap_8 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_62 ();
 sg13g2_decap_8 FILLER_24_69 ();
 sg13g2_decap_8 FILLER_24_76 ();
 sg13g2_decap_8 FILLER_24_83 ();
 sg13g2_decap_4 FILLER_24_90 ();
 sg13g2_fill_2 FILLER_24_94 ();
 sg13g2_decap_8 FILLER_24_101 ();
 sg13g2_fill_2 FILLER_24_108 ();
 sg13g2_fill_2 FILLER_24_114 ();
 sg13g2_fill_1 FILLER_24_121 ();
 sg13g2_fill_2 FILLER_24_201 ();
 sg13g2_fill_1 FILLER_24_203 ();
 sg13g2_decap_4 FILLER_24_257 ();
 sg13g2_fill_2 FILLER_24_261 ();
 sg13g2_fill_1 FILLER_24_273 ();
 sg13g2_fill_1 FILLER_24_284 ();
 sg13g2_decap_8 FILLER_24_311 ();
 sg13g2_decap_8 FILLER_24_318 ();
 sg13g2_decap_8 FILLER_24_325 ();
 sg13g2_decap_8 FILLER_24_332 ();
 sg13g2_decap_8 FILLER_24_339 ();
 sg13g2_decap_8 FILLER_24_346 ();
 sg13g2_decap_8 FILLER_24_353 ();
 sg13g2_decap_8 FILLER_24_360 ();
 sg13g2_decap_8 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_388 ();
 sg13g2_decap_8 FILLER_24_395 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_4 FILLER_25_21 ();
 sg13g2_fill_1 FILLER_25_25 ();
 sg13g2_decap_4 FILLER_25_58 ();
 sg13g2_fill_1 FILLER_25_62 ();
 sg13g2_fill_2 FILLER_25_89 ();
 sg13g2_fill_1 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_97 ();
 sg13g2_decap_8 FILLER_25_104 ();
 sg13g2_decap_8 FILLER_25_111 ();
 sg13g2_decap_8 FILLER_25_136 ();
 sg13g2_decap_4 FILLER_25_147 ();
 sg13g2_fill_1 FILLER_25_151 ();
 sg13g2_fill_2 FILLER_25_168 ();
 sg13g2_fill_1 FILLER_25_198 ();
 sg13g2_fill_1 FILLER_25_211 ();
 sg13g2_fill_1 FILLER_25_241 ();
 sg13g2_fill_2 FILLER_25_250 ();
 sg13g2_fill_1 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_fill_2 FILLER_25_273 ();
 sg13g2_fill_1 FILLER_25_295 ();
 sg13g2_decap_8 FILLER_25_304 ();
 sg13g2_decap_8 FILLER_25_311 ();
 sg13g2_decap_8 FILLER_25_318 ();
 sg13g2_decap_8 FILLER_25_325 ();
 sg13g2_decap_8 FILLER_25_332 ();
 sg13g2_decap_8 FILLER_25_339 ();
 sg13g2_decap_8 FILLER_25_346 ();
 sg13g2_decap_8 FILLER_25_353 ();
 sg13g2_decap_8 FILLER_25_360 ();
 sg13g2_decap_8 FILLER_25_367 ();
 sg13g2_decap_8 FILLER_25_374 ();
 sg13g2_decap_8 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_4 FILLER_26_28 ();
 sg13g2_fill_2 FILLER_26_32 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_fill_2 FILLER_26_71 ();
 sg13g2_decap_4 FILLER_26_120 ();
 sg13g2_fill_1 FILLER_26_124 ();
 sg13g2_fill_2 FILLER_26_135 ();
 sg13g2_fill_1 FILLER_26_137 ();
 sg13g2_decap_8 FILLER_26_143 ();
 sg13g2_decap_8 FILLER_26_150 ();
 sg13g2_fill_1 FILLER_26_187 ();
 sg13g2_decap_8 FILLER_26_201 ();
 sg13g2_decap_8 FILLER_26_208 ();
 sg13g2_fill_2 FILLER_26_215 ();
 sg13g2_decap_4 FILLER_26_266 ();
 sg13g2_fill_2 FILLER_26_270 ();
 sg13g2_decap_4 FILLER_26_276 ();
 sg13g2_fill_2 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_286 ();
 sg13g2_decap_8 FILLER_26_293 ();
 sg13g2_decap_8 FILLER_26_300 ();
 sg13g2_decap_8 FILLER_26_307 ();
 sg13g2_decap_8 FILLER_26_314 ();
 sg13g2_decap_8 FILLER_26_326 ();
 sg13g2_decap_8 FILLER_26_333 ();
 sg13g2_decap_8 FILLER_26_340 ();
 sg13g2_decap_8 FILLER_26_347 ();
 sg13g2_decap_8 FILLER_26_354 ();
 sg13g2_decap_8 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_39 ();
 sg13g2_fill_1 FILLER_27_46 ();
 sg13g2_fill_1 FILLER_27_112 ();
 sg13g2_decap_4 FILLER_27_139 ();
 sg13g2_decap_4 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_decap_8 FILLER_27_193 ();
 sg13g2_decap_8 FILLER_27_200 ();
 sg13g2_fill_1 FILLER_27_207 ();
 sg13g2_fill_1 FILLER_27_216 ();
 sg13g2_decap_8 FILLER_27_236 ();
 sg13g2_decap_8 FILLER_27_243 ();
 sg13g2_fill_2 FILLER_27_250 ();
 sg13g2_fill_2 FILLER_27_293 ();
 sg13g2_fill_1 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_307 ();
 sg13g2_fill_2 FILLER_27_314 ();
 sg13g2_fill_1 FILLER_27_326 ();
 sg13g2_decap_8 FILLER_27_353 ();
 sg13g2_decap_8 FILLER_27_360 ();
 sg13g2_decap_8 FILLER_27_367 ();
 sg13g2_decap_8 FILLER_27_374 ();
 sg13g2_decap_8 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_decap_8 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_4 FILLER_28_54 ();
 sg13g2_fill_2 FILLER_28_68 ();
 sg13g2_fill_2 FILLER_28_80 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_fill_2 FILLER_28_168 ();
 sg13g2_fill_1 FILLER_28_175 ();
 sg13g2_fill_2 FILLER_28_191 ();
 sg13g2_fill_1 FILLER_28_198 ();
 sg13g2_fill_2 FILLER_28_224 ();
 sg13g2_fill_1 FILLER_28_238 ();
 sg13g2_fill_2 FILLER_28_251 ();
 sg13g2_fill_2 FILLER_28_256 ();
 sg13g2_fill_1 FILLER_28_258 ();
 sg13g2_fill_2 FILLER_28_273 ();
 sg13g2_fill_2 FILLER_28_285 ();
 sg13g2_fill_1 FILLER_28_287 ();
 sg13g2_decap_8 FILLER_28_354 ();
 sg13g2_decap_8 FILLER_28_361 ();
 sg13g2_decap_8 FILLER_28_368 ();
 sg13g2_decap_8 FILLER_28_375 ();
 sg13g2_decap_8 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_4 ();
 sg13g2_decap_4 FILLER_29_65 ();
 sg13g2_fill_2 FILLER_29_69 ();
 sg13g2_decap_8 FILLER_29_81 ();
 sg13g2_fill_2 FILLER_29_88 ();
 sg13g2_fill_1 FILLER_29_90 ();
 sg13g2_fill_2 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_142 ();
 sg13g2_fill_1 FILLER_29_148 ();
 sg13g2_decap_8 FILLER_29_158 ();
 sg13g2_decap_8 FILLER_29_165 ();
 sg13g2_decap_4 FILLER_29_172 ();
 sg13g2_fill_2 FILLER_29_176 ();
 sg13g2_fill_2 FILLER_29_195 ();
 sg13g2_decap_4 FILLER_29_202 ();
 sg13g2_fill_1 FILLER_29_232 ();
 sg13g2_decap_4 FILLER_29_307 ();
 sg13g2_fill_2 FILLER_29_311 ();
 sg13g2_fill_2 FILLER_29_347 ();
 sg13g2_fill_1 FILLER_29_349 ();
 sg13g2_decap_8 FILLER_29_376 ();
 sg13g2_decap_8 FILLER_29_383 ();
 sg13g2_decap_8 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_4 FILLER_30_14 ();
 sg13g2_fill_1 FILLER_30_18 ();
 sg13g2_fill_1 FILLER_30_27 ();
 sg13g2_fill_2 FILLER_30_38 ();
 sg13g2_fill_2 FILLER_30_97 ();
 sg13g2_fill_1 FILLER_30_99 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_4 FILLER_30_119 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_decap_8 FILLER_30_128 ();
 sg13g2_decap_8 FILLER_30_135 ();
 sg13g2_fill_2 FILLER_30_142 ();
 sg13g2_fill_1 FILLER_30_144 ();
 sg13g2_decap_8 FILLER_30_148 ();
 sg13g2_decap_4 FILLER_30_155 ();
 sg13g2_fill_1 FILLER_30_159 ();
 sg13g2_fill_1 FILLER_30_173 ();
 sg13g2_fill_2 FILLER_30_202 ();
 sg13g2_decap_4 FILLER_30_208 ();
 sg13g2_fill_1 FILLER_30_212 ();
 sg13g2_decap_8 FILLER_30_218 ();
 sg13g2_fill_1 FILLER_30_235 ();
 sg13g2_fill_1 FILLER_30_249 ();
 sg13g2_fill_2 FILLER_30_254 ();
 sg13g2_fill_2 FILLER_30_260 ();
 sg13g2_fill_1 FILLER_30_262 ();
 sg13g2_decap_8 FILLER_30_269 ();
 sg13g2_decap_4 FILLER_30_276 ();
 sg13g2_fill_2 FILLER_30_280 ();
 sg13g2_decap_4 FILLER_30_286 ();
 sg13g2_fill_2 FILLER_30_290 ();
 sg13g2_decap_8 FILLER_30_302 ();
 sg13g2_decap_8 FILLER_30_309 ();
 sg13g2_decap_4 FILLER_30_316 ();
 sg13g2_fill_2 FILLER_30_320 ();
 sg13g2_fill_2 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_30_377 ();
 sg13g2_decap_8 FILLER_30_384 ();
 sg13g2_decap_8 FILLER_30_391 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_4 FILLER_31_42 ();
 sg13g2_fill_2 FILLER_31_46 ();
 sg13g2_decap_8 FILLER_31_62 ();
 sg13g2_decap_8 FILLER_31_69 ();
 sg13g2_decap_8 FILLER_31_80 ();
 sg13g2_fill_1 FILLER_31_87 ();
 sg13g2_decap_8 FILLER_31_99 ();
 sg13g2_decap_8 FILLER_31_106 ();
 sg13g2_fill_1 FILLER_31_113 ();
 sg13g2_fill_2 FILLER_31_119 ();
 sg13g2_fill_1 FILLER_31_121 ();
 sg13g2_decap_4 FILLER_31_127 ();
 sg13g2_fill_2 FILLER_31_131 ();
 sg13g2_fill_1 FILLER_31_150 ();
 sg13g2_fill_1 FILLER_31_186 ();
 sg13g2_fill_2 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_219 ();
 sg13g2_fill_2 FILLER_31_226 ();
 sg13g2_fill_1 FILLER_31_233 ();
 sg13g2_decap_8 FILLER_31_237 ();
 sg13g2_fill_1 FILLER_31_244 ();
 sg13g2_decap_8 FILLER_31_271 ();
 sg13g2_fill_2 FILLER_31_278 ();
 sg13g2_fill_1 FILLER_31_284 ();
 sg13g2_decap_4 FILLER_31_325 ();
 sg13g2_fill_2 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_335 ();
 sg13g2_fill_1 FILLER_31_342 ();
 sg13g2_fill_1 FILLER_31_353 ();
 sg13g2_decap_8 FILLER_31_380 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_41 ();
 sg13g2_decap_8 FILLER_32_48 ();
 sg13g2_decap_4 FILLER_32_55 ();
 sg13g2_decap_8 FILLER_32_69 ();
 sg13g2_fill_2 FILLER_32_95 ();
 sg13g2_decap_4 FILLER_32_106 ();
 sg13g2_fill_1 FILLER_32_110 ();
 sg13g2_fill_2 FILLER_32_124 ();
 sg13g2_fill_1 FILLER_32_150 ();
 sg13g2_decap_8 FILLER_32_198 ();
 sg13g2_decap_8 FILLER_32_213 ();
 sg13g2_decap_4 FILLER_32_220 ();
 sg13g2_fill_1 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_fill_2 FILLER_32_272 ();
 sg13g2_fill_1 FILLER_32_274 ();
 sg13g2_decap_8 FILLER_32_341 ();
 sg13g2_fill_1 FILLER_32_348 ();
 sg13g2_decap_8 FILLER_32_367 ();
 sg13g2_decap_8 FILLER_32_374 ();
 sg13g2_decap_8 FILLER_32_381 ();
 sg13g2_decap_8 FILLER_32_388 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_4 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_18 ();
 sg13g2_decap_4 FILLER_33_160 ();
 sg13g2_fill_1 FILLER_33_169 ();
 sg13g2_fill_1 FILLER_33_178 ();
 sg13g2_decap_8 FILLER_33_188 ();
 sg13g2_decap_8 FILLER_33_195 ();
 sg13g2_fill_2 FILLER_33_202 ();
 sg13g2_fill_1 FILLER_33_209 ();
 sg13g2_decap_8 FILLER_33_236 ();
 sg13g2_decap_8 FILLER_33_243 ();
 sg13g2_decap_8 FILLER_33_276 ();
 sg13g2_decap_4 FILLER_33_283 ();
 sg13g2_fill_2 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_303 ();
 sg13g2_fill_2 FILLER_33_312 ();
 sg13g2_fill_1 FILLER_33_314 ();
 sg13g2_fill_2 FILLER_33_320 ();
 sg13g2_fill_2 FILLER_33_348 ();
 sg13g2_fill_1 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_377 ();
 sg13g2_decap_8 FILLER_33_384 ();
 sg13g2_decap_8 FILLER_33_391 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_4 FILLER_34_14 ();
 sg13g2_fill_2 FILLER_34_18 ();
 sg13g2_fill_1 FILLER_34_48 ();
 sg13g2_fill_2 FILLER_34_75 ();
 sg13g2_fill_1 FILLER_34_131 ();
 sg13g2_decap_8 FILLER_34_137 ();
 sg13g2_fill_1 FILLER_34_165 ();
 sg13g2_decap_4 FILLER_34_171 ();
 sg13g2_fill_1 FILLER_34_175 ();
 sg13g2_fill_2 FILLER_34_180 ();
 sg13g2_decap_4 FILLER_34_186 ();
 sg13g2_fill_2 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_202 ();
 sg13g2_decap_4 FILLER_34_212 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_decap_8 FILLER_34_247 ();
 sg13g2_fill_2 FILLER_34_254 ();
 sg13g2_fill_1 FILLER_34_256 ();
 sg13g2_decap_8 FILLER_34_261 ();
 sg13g2_fill_1 FILLER_34_268 ();
 sg13g2_decap_8 FILLER_34_295 ();
 sg13g2_decap_8 FILLER_34_302 ();
 sg13g2_decap_8 FILLER_34_309 ();
 sg13g2_decap_4 FILLER_34_316 ();
 sg13g2_fill_1 FILLER_34_346 ();
 sg13g2_decap_8 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_384 ();
 sg13g2_decap_8 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_45 ();
 sg13g2_fill_2 FILLER_35_52 ();
 sg13g2_fill_2 FILLER_35_72 ();
 sg13g2_fill_1 FILLER_35_74 ();
 sg13g2_decap_8 FILLER_35_115 ();
 sg13g2_decap_8 FILLER_35_122 ();
 sg13g2_fill_1 FILLER_35_129 ();
 sg13g2_decap_8 FILLER_35_142 ();
 sg13g2_decap_4 FILLER_35_149 ();
 sg13g2_fill_1 FILLER_35_153 ();
 sg13g2_decap_8 FILLER_35_159 ();
 sg13g2_decap_4 FILLER_35_166 ();
 sg13g2_fill_1 FILLER_35_170 ();
 sg13g2_fill_2 FILLER_35_181 ();
 sg13g2_fill_1 FILLER_35_183 ();
 sg13g2_fill_1 FILLER_35_191 ();
 sg13g2_fill_1 FILLER_35_202 ();
 sg13g2_fill_1 FILLER_35_215 ();
 sg13g2_fill_2 FILLER_35_225 ();
 sg13g2_fill_1 FILLER_35_244 ();
 sg13g2_decap_8 FILLER_35_270 ();
 sg13g2_decap_8 FILLER_35_277 ();
 sg13g2_decap_4 FILLER_35_284 ();
 sg13g2_fill_2 FILLER_35_292 ();
 sg13g2_fill_1 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_299 ();
 sg13g2_decap_8 FILLER_35_306 ();
 sg13g2_decap_8 FILLER_35_313 ();
 sg13g2_decap_4 FILLER_35_320 ();
 sg13g2_fill_1 FILLER_35_324 ();
 sg13g2_fill_1 FILLER_35_367 ();
 sg13g2_decap_8 FILLER_35_394 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_4 FILLER_36_28 ();
 sg13g2_fill_1 FILLER_36_32 ();
 sg13g2_decap_4 FILLER_36_41 ();
 sg13g2_fill_2 FILLER_36_57 ();
 sg13g2_fill_1 FILLER_36_59 ();
 sg13g2_decap_8 FILLER_36_65 ();
 sg13g2_decap_8 FILLER_36_80 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_145 ();
 sg13g2_fill_2 FILLER_36_156 ();
 sg13g2_fill_1 FILLER_36_158 ();
 sg13g2_decap_8 FILLER_36_169 ();
 sg13g2_decap_4 FILLER_36_176 ();
 sg13g2_fill_1 FILLER_36_180 ();
 sg13g2_fill_2 FILLER_36_194 ();
 sg13g2_fill_1 FILLER_36_233 ();
 sg13g2_fill_2 FILLER_36_250 ();
 sg13g2_fill_2 FILLER_36_283 ();
 sg13g2_fill_1 FILLER_36_285 ();
 sg13g2_fill_1 FILLER_36_294 ();
 sg13g2_fill_2 FILLER_36_321 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_fill_1 FILLER_36_329 ();
 sg13g2_fill_2 FILLER_36_334 ();
 sg13g2_fill_1 FILLER_36_336 ();
 sg13g2_decap_8 FILLER_36_347 ();
 sg13g2_decap_8 FILLER_36_354 ();
 sg13g2_fill_2 FILLER_36_361 ();
 sg13g2_fill_1 FILLER_36_375 ();
 sg13g2_fill_2 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_4 FILLER_37_28 ();
 sg13g2_fill_1 FILLER_37_32 ();
 sg13g2_fill_2 FILLER_37_44 ();
 sg13g2_fill_1 FILLER_37_46 ();
 sg13g2_fill_1 FILLER_37_66 ();
 sg13g2_decap_8 FILLER_37_80 ();
 sg13g2_decap_8 FILLER_37_87 ();
 sg13g2_decap_8 FILLER_37_94 ();
 sg13g2_decap_4 FILLER_37_101 ();
 sg13g2_fill_2 FILLER_37_140 ();
 sg13g2_fill_2 FILLER_37_166 ();
 sg13g2_fill_1 FILLER_37_178 ();
 sg13g2_decap_8 FILLER_37_193 ();
 sg13g2_fill_2 FILLER_37_200 ();
 sg13g2_fill_2 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_216 ();
 sg13g2_decap_8 FILLER_37_223 ();
 sg13g2_fill_1 FILLER_37_230 ();
 sg13g2_fill_2 FILLER_37_259 ();
 sg13g2_fill_1 FILLER_37_261 ();
 sg13g2_fill_2 FILLER_37_348 ();
 sg13g2_fill_1 FILLER_37_350 ();
 sg13g2_decap_4 FILLER_37_356 ();
 sg13g2_decap_4 FILLER_37_363 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_4 FILLER_38_21 ();
 sg13g2_fill_2 FILLER_38_25 ();
 sg13g2_fill_2 FILLER_38_57 ();
 sg13g2_fill_1 FILLER_38_59 ();
 sg13g2_fill_2 FILLER_38_102 ();
 sg13g2_fill_1 FILLER_38_104 ();
 sg13g2_fill_2 FILLER_38_113 ();
 sg13g2_fill_2 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_fill_2 FILLER_38_207 ();
 sg13g2_decap_4 FILLER_38_214 ();
 sg13g2_fill_1 FILLER_38_233 ();
 sg13g2_fill_2 FILLER_38_239 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_fill_1 FILLER_38_252 ();
 sg13g2_fill_1 FILLER_38_270 ();
 sg13g2_fill_1 FILLER_38_290 ();
 sg13g2_decap_8 FILLER_38_316 ();
 sg13g2_fill_2 FILLER_38_323 ();
 sg13g2_fill_1 FILLER_38_325 ();
 sg13g2_decap_8 FILLER_38_330 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_fill_1 FILLER_39_21 ();
 sg13g2_fill_2 FILLER_39_41 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_fill_2 FILLER_39_105 ();
 sg13g2_fill_1 FILLER_39_115 ();
 sg13g2_fill_1 FILLER_39_162 ();
 sg13g2_decap_8 FILLER_39_181 ();
 sg13g2_fill_2 FILLER_39_188 ();
 sg13g2_fill_1 FILLER_39_190 ();
 sg13g2_fill_1 FILLER_39_225 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_decap_8 FILLER_39_272 ();
 sg13g2_decap_4 FILLER_39_295 ();
 sg13g2_fill_1 FILLER_39_299 ();
 sg13g2_decap_8 FILLER_39_310 ();
 sg13g2_decap_8 FILLER_39_317 ();
 sg13g2_decap_4 FILLER_39_324 ();
 sg13g2_decap_4 FILLER_39_342 ();
 sg13g2_fill_2 FILLER_39_346 ();
 sg13g2_fill_2 FILLER_39_352 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_fill_1 FILLER_40_14 ();
 sg13g2_fill_1 FILLER_40_41 ();
 sg13g2_fill_2 FILLER_40_54 ();
 sg13g2_fill_1 FILLER_40_56 ();
 sg13g2_fill_2 FILLER_40_62 ();
 sg13g2_decap_4 FILLER_40_74 ();
 sg13g2_fill_1 FILLER_40_78 ();
 sg13g2_decap_4 FILLER_40_87 ();
 sg13g2_fill_2 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_4 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_121 ();
 sg13g2_decap_4 FILLER_40_128 ();
 sg13g2_fill_2 FILLER_40_144 ();
 sg13g2_decap_4 FILLER_40_150 ();
 sg13g2_fill_2 FILLER_40_154 ();
 sg13g2_fill_1 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_166 ();
 sg13g2_fill_1 FILLER_40_173 ();
 sg13g2_decap_8 FILLER_40_187 ();
 sg13g2_fill_2 FILLER_40_194 ();
 sg13g2_fill_2 FILLER_40_201 ();
 sg13g2_decap_4 FILLER_40_227 ();
 sg13g2_fill_1 FILLER_40_231 ();
 sg13g2_decap_8 FILLER_40_240 ();
 sg13g2_decap_8 FILLER_40_247 ();
 sg13g2_fill_1 FILLER_40_254 ();
 sg13g2_decap_8 FILLER_40_277 ();
 sg13g2_decap_4 FILLER_40_284 ();
 sg13g2_fill_2 FILLER_40_288 ();
 sg13g2_fill_2 FILLER_40_294 ();
 sg13g2_decap_8 FILLER_40_353 ();
 sg13g2_fill_1 FILLER_40_360 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_fill_2 FILLER_40_406 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_fill_2 FILLER_41_21 ();
 sg13g2_fill_1 FILLER_41_23 ();
 sg13g2_decap_4 FILLER_41_38 ();
 sg13g2_fill_1 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_4 FILLER_41_84 ();
 sg13g2_fill_2 FILLER_41_88 ();
 sg13g2_fill_2 FILLER_41_115 ();
 sg13g2_fill_1 FILLER_41_117 ();
 sg13g2_decap_4 FILLER_41_123 ();
 sg13g2_fill_1 FILLER_41_127 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_fill_2 FILLER_41_140 ();
 sg13g2_fill_1 FILLER_41_169 ();
 sg13g2_decap_8 FILLER_41_182 ();
 sg13g2_decap_4 FILLER_41_189 ();
 sg13g2_fill_1 FILLER_41_193 ();
 sg13g2_decap_8 FILLER_41_202 ();
 sg13g2_fill_2 FILLER_41_209 ();
 sg13g2_decap_4 FILLER_41_219 ();
 sg13g2_fill_1 FILLER_41_223 ();
 sg13g2_decap_8 FILLER_41_244 ();
 sg13g2_decap_8 FILLER_41_251 ();
 sg13g2_decap_8 FILLER_41_258 ();
 sg13g2_fill_2 FILLER_41_265 ();
 sg13g2_fill_1 FILLER_41_267 ();
 sg13g2_fill_2 FILLER_41_277 ();
 sg13g2_fill_2 FILLER_41_305 ();
 sg13g2_fill_1 FILLER_41_307 ();
 sg13g2_decap_4 FILLER_41_334 ();
 sg13g2_fill_1 FILLER_41_338 ();
 sg13g2_decap_8 FILLER_41_373 ();
 sg13g2_fill_2 FILLER_41_380 ();
 sg13g2_fill_1 FILLER_41_382 ();
 sg13g2_fill_1 FILLER_41_387 ();
 sg13g2_decap_8 FILLER_41_397 ();
 sg13g2_decap_4 FILLER_41_404 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_4 FILLER_42_39 ();
 sg13g2_decap_8 FILLER_42_69 ();
 sg13g2_fill_2 FILLER_42_76 ();
 sg13g2_fill_1 FILLER_42_78 ();
 sg13g2_decap_8 FILLER_42_134 ();
 sg13g2_fill_2 FILLER_42_157 ();
 sg13g2_fill_2 FILLER_42_187 ();
 sg13g2_decap_8 FILLER_42_204 ();
 sg13g2_decap_8 FILLER_42_211 ();
 sg13g2_decap_8 FILLER_42_218 ();
 sg13g2_fill_1 FILLER_42_229 ();
 sg13g2_decap_4 FILLER_42_240 ();
 sg13g2_fill_1 FILLER_42_268 ();
 sg13g2_fill_2 FILLER_42_277 ();
 sg13g2_fill_2 FILLER_42_283 ();
 sg13g2_fill_1 FILLER_42_285 ();
 sg13g2_fill_2 FILLER_42_291 ();
 sg13g2_fill_1 FILLER_42_293 ();
 sg13g2_decap_8 FILLER_42_325 ();
 sg13g2_decap_8 FILLER_42_332 ();
 sg13g2_fill_2 FILLER_42_339 ();
 sg13g2_decap_4 FILLER_42_355 ();
 sg13g2_fill_2 FILLER_42_359 ();
 sg13g2_decap_4 FILLER_42_364 ();
 sg13g2_fill_1 FILLER_42_368 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_fill_2 FILLER_43_14 ();
 sg13g2_fill_1 FILLER_43_16 ();
 sg13g2_decap_4 FILLER_43_43 ();
 sg13g2_fill_2 FILLER_43_123 ();
 sg13g2_fill_2 FILLER_43_187 ();
 sg13g2_fill_1 FILLER_43_189 ();
 sg13g2_fill_2 FILLER_43_200 ();
 sg13g2_fill_1 FILLER_43_202 ();
 sg13g2_decap_8 FILLER_43_221 ();
 sg13g2_decap_4 FILLER_43_228 ();
 sg13g2_fill_1 FILLER_43_232 ();
 sg13g2_fill_1 FILLER_43_254 ();
 sg13g2_fill_2 FILLER_43_258 ();
 sg13g2_fill_1 FILLER_43_264 ();
 sg13g2_decap_8 FILLER_43_309 ();
 sg13g2_decap_8 FILLER_43_316 ();
 sg13g2_decap_4 FILLER_43_323 ();
 sg13g2_fill_1 FILLER_43_327 ();
 sg13g2_fill_2 FILLER_43_337 ();
 sg13g2_fill_2 FILLER_43_380 ();
 sg13g2_fill_1 FILLER_43_382 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_32 ();
 sg13g2_fill_1 FILLER_44_93 ();
 sg13g2_fill_2 FILLER_44_114 ();
 sg13g2_fill_1 FILLER_44_116 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_fill_2 FILLER_44_168 ();
 sg13g2_fill_1 FILLER_44_200 ();
 sg13g2_decap_8 FILLER_44_221 ();
 sg13g2_fill_1 FILLER_44_228 ();
 sg13g2_fill_2 FILLER_44_238 ();
 sg13g2_fill_1 FILLER_44_240 ();
 sg13g2_fill_2 FILLER_44_257 ();
 sg13g2_fill_2 FILLER_44_267 ();
 sg13g2_fill_1 FILLER_44_269 ();
 sg13g2_decap_8 FILLER_44_300 ();
 sg13g2_decap_4 FILLER_44_307 ();
 sg13g2_fill_2 FILLER_44_311 ();
 sg13g2_fill_2 FILLER_44_317 ();
 sg13g2_fill_2 FILLER_44_381 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_4 FILLER_45_14 ();
 sg13g2_fill_2 FILLER_45_18 ();
 sg13g2_decap_8 FILLER_45_46 ();
 sg13g2_decap_8 FILLER_45_53 ();
 sg13g2_decap_4 FILLER_45_60 ();
 sg13g2_fill_1 FILLER_45_64 ();
 sg13g2_fill_2 FILLER_45_80 ();
 sg13g2_fill_1 FILLER_45_87 ();
 sg13g2_fill_2 FILLER_45_93 ();
 sg13g2_decap_8 FILLER_45_115 ();
 sg13g2_decap_4 FILLER_45_122 ();
 sg13g2_fill_1 FILLER_45_126 ();
 sg13g2_fill_1 FILLER_45_146 ();
 sg13g2_fill_2 FILLER_45_159 ();
 sg13g2_fill_1 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_169 ();
 sg13g2_decap_4 FILLER_45_176 ();
 sg13g2_fill_1 FILLER_45_180 ();
 sg13g2_fill_2 FILLER_45_185 ();
 sg13g2_decap_8 FILLER_45_220 ();
 sg13g2_fill_1 FILLER_45_227 ();
 sg13g2_fill_1 FILLER_45_237 ();
 sg13g2_fill_2 FILLER_45_261 ();
 sg13g2_fill_1 FILLER_45_288 ();
 sg13g2_fill_2 FILLER_45_294 ();
 sg13g2_fill_1 FILLER_45_296 ();
 sg13g2_fill_1 FILLER_45_333 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_fill_1 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_58 ();
 sg13g2_decap_8 FILLER_46_65 ();
 sg13g2_fill_1 FILLER_46_72 ();
 sg13g2_decap_8 FILLER_46_83 ();
 sg13g2_fill_2 FILLER_46_90 ();
 sg13g2_fill_1 FILLER_46_92 ();
 sg13g2_decap_8 FILLER_46_96 ();
 sg13g2_decap_8 FILLER_46_108 ();
 sg13g2_decap_8 FILLER_46_115 ();
 sg13g2_decap_4 FILLER_46_122 ();
 sg13g2_fill_1 FILLER_46_126 ();
 sg13g2_fill_2 FILLER_46_135 ();
 sg13g2_fill_1 FILLER_46_137 ();
 sg13g2_fill_1 FILLER_46_175 ();
 sg13g2_fill_2 FILLER_46_179 ();
 sg13g2_fill_2 FILLER_46_229 ();
 sg13g2_decap_4 FILLER_46_262 ();
 sg13g2_fill_1 FILLER_46_266 ();
 sg13g2_decap_8 FILLER_46_276 ();
 sg13g2_decap_4 FILLER_46_283 ();
 sg13g2_fill_1 FILLER_46_287 ();
 sg13g2_decap_8 FILLER_46_326 ();
 sg13g2_decap_8 FILLER_46_333 ();
 sg13g2_decap_8 FILLER_46_340 ();
 sg13g2_fill_2 FILLER_46_347 ();
 sg13g2_fill_1 FILLER_46_349 ();
 sg13g2_decap_8 FILLER_46_354 ();
 sg13g2_decap_8 FILLER_46_361 ();
 sg13g2_fill_2 FILLER_46_368 ();
 sg13g2_decap_4 FILLER_46_374 ();
 sg13g2_fill_1 FILLER_46_378 ();
 sg13g2_decap_8 FILLER_46_397 ();
 sg13g2_decap_4 FILLER_46_404 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_4 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_43 ();
 sg13g2_fill_2 FILLER_47_50 ();
 sg13g2_fill_1 FILLER_47_62 ();
 sg13g2_decap_4 FILLER_47_67 ();
 sg13g2_fill_1 FILLER_47_71 ();
 sg13g2_decap_8 FILLER_47_82 ();
 sg13g2_fill_2 FILLER_47_89 ();
 sg13g2_fill_1 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_100 ();
 sg13g2_decap_4 FILLER_47_107 ();
 sg13g2_decap_8 FILLER_47_127 ();
 sg13g2_fill_2 FILLER_47_196 ();
 sg13g2_fill_1 FILLER_47_207 ();
 sg13g2_fill_2 FILLER_47_218 ();
 sg13g2_fill_1 FILLER_47_220 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_fill_2 FILLER_47_280 ();
 sg13g2_fill_1 FILLER_47_282 ();
 sg13g2_fill_2 FILLER_47_301 ();
 sg13g2_decap_8 FILLER_47_342 ();
 sg13g2_decap_8 FILLER_47_349 ();
 sg13g2_decap_8 FILLER_47_356 ();
 sg13g2_decap_8 FILLER_47_363 ();
 sg13g2_decap_8 FILLER_47_370 ();
 sg13g2_decap_8 FILLER_47_377 ();
 sg13g2_decap_8 FILLER_47_384 ();
 sg13g2_decap_8 FILLER_47_391 ();
 sg13g2_decap_8 FILLER_47_398 ();
 sg13g2_decap_4 FILLER_47_405 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_4 FILLER_48_35 ();
 sg13g2_fill_1 FILLER_48_39 ();
 sg13g2_fill_2 FILLER_48_50 ();
 sg13g2_decap_4 FILLER_48_87 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_fill_2 FILLER_48_112 ();
 sg13g2_fill_2 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_fill_2 FILLER_48_182 ();
 sg13g2_fill_1 FILLER_48_184 ();
 sg13g2_decap_8 FILLER_48_198 ();
 sg13g2_decap_8 FILLER_48_205 ();
 sg13g2_decap_8 FILLER_48_212 ();
 sg13g2_fill_2 FILLER_48_219 ();
 sg13g2_fill_1 FILLER_48_238 ();
 sg13g2_fill_2 FILLER_48_254 ();
 sg13g2_decap_8 FILLER_48_359 ();
 sg13g2_fill_2 FILLER_48_366 ();
 sg13g2_fill_1 FILLER_48_368 ();
 sg13g2_decap_8 FILLER_48_374 ();
 sg13g2_decap_8 FILLER_48_381 ();
 sg13g2_decap_8 FILLER_48_388 ();
 sg13g2_decap_8 FILLER_48_395 ();
 sg13g2_decap_8 FILLER_48_402 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_4 FILLER_49_28 ();
 sg13g2_decap_4 FILLER_49_114 ();
 sg13g2_fill_1 FILLER_49_118 ();
 sg13g2_decap_8 FILLER_49_128 ();
 sg13g2_decap_8 FILLER_49_135 ();
 sg13g2_decap_8 FILLER_49_142 ();
 sg13g2_fill_2 FILLER_49_149 ();
 sg13g2_decap_8 FILLER_49_156 ();
 sg13g2_decap_8 FILLER_49_163 ();
 sg13g2_decap_8 FILLER_49_170 ();
 sg13g2_decap_8 FILLER_49_177 ();
 sg13g2_decap_4 FILLER_49_184 ();
 sg13g2_fill_1 FILLER_49_188 ();
 sg13g2_fill_2 FILLER_49_205 ();
 sg13g2_fill_2 FILLER_49_227 ();
 sg13g2_fill_2 FILLER_49_239 ();
 sg13g2_fill_1 FILLER_49_241 ();
 sg13g2_fill_2 FILLER_49_251 ();
 sg13g2_decap_4 FILLER_49_263 ();
 sg13g2_fill_1 FILLER_49_267 ();
 sg13g2_fill_2 FILLER_49_280 ();
 sg13g2_fill_1 FILLER_49_282 ();
 sg13g2_fill_2 FILLER_49_329 ();
 sg13g2_decap_8 FILLER_49_365 ();
 sg13g2_decap_8 FILLER_49_372 ();
 sg13g2_decap_8 FILLER_49_379 ();
 sg13g2_decap_8 FILLER_49_386 ();
 sg13g2_decap_8 FILLER_49_393 ();
 sg13g2_decap_8 FILLER_49_400 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_fill_2 FILLER_50_28 ();
 sg13g2_fill_1 FILLER_50_30 ();
 sg13g2_decap_4 FILLER_50_129 ();
 sg13g2_fill_1 FILLER_50_133 ();
 sg13g2_decap_4 FILLER_50_147 ();
 sg13g2_fill_1 FILLER_50_156 ();
 sg13g2_fill_1 FILLER_50_161 ();
 sg13g2_decap_8 FILLER_50_167 ();
 sg13g2_decap_8 FILLER_50_174 ();
 sg13g2_fill_2 FILLER_50_181 ();
 sg13g2_fill_2 FILLER_50_214 ();
 sg13g2_fill_1 FILLER_50_216 ();
 sg13g2_decap_8 FILLER_50_246 ();
 sg13g2_decap_8 FILLER_50_253 ();
 sg13g2_decap_8 FILLER_50_260 ();
 sg13g2_decap_8 FILLER_50_267 ();
 sg13g2_fill_1 FILLER_50_274 ();
 sg13g2_decap_8 FILLER_50_301 ();
 sg13g2_decap_8 FILLER_50_308 ();
 sg13g2_decap_8 FILLER_50_315 ();
 sg13g2_decap_4 FILLER_50_322 ();
 sg13g2_fill_1 FILLER_50_326 ();
 sg13g2_fill_1 FILLER_50_339 ();
 sg13g2_fill_2 FILLER_50_348 ();
 sg13g2_fill_1 FILLER_50_350 ();
 sg13g2_fill_2 FILLER_50_356 ();
 sg13g2_decap_8 FILLER_50_395 ();
 sg13g2_decap_8 FILLER_50_402 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_4 FILLER_51_28 ();
 sg13g2_fill_2 FILLER_51_32 ();
 sg13g2_fill_1 FILLER_51_48 ();
 sg13g2_decap_8 FILLER_51_53 ();
 sg13g2_decap_8 FILLER_51_60 ();
 sg13g2_decap_4 FILLER_51_67 ();
 sg13g2_fill_1 FILLER_51_81 ();
 sg13g2_fill_1 FILLER_51_87 ();
 sg13g2_fill_2 FILLER_51_107 ();
 sg13g2_fill_2 FILLER_51_119 ();
 sg13g2_fill_2 FILLER_51_131 ();
 sg13g2_fill_1 FILLER_51_146 ();
 sg13g2_decap_4 FILLER_51_167 ();
 sg13g2_fill_2 FILLER_51_201 ();
 sg13g2_fill_1 FILLER_51_203 ();
 sg13g2_fill_1 FILLER_51_219 ();
 sg13g2_fill_2 FILLER_51_235 ();
 sg13g2_fill_1 FILLER_51_237 ();
 sg13g2_decap_4 FILLER_51_253 ();
 sg13g2_decap_8 FILLER_51_261 ();
 sg13g2_fill_1 FILLER_51_268 ();
 sg13g2_decap_4 FILLER_51_273 ();
 sg13g2_fill_2 FILLER_51_277 ();
 sg13g2_fill_2 FILLER_51_284 ();
 sg13g2_decap_8 FILLER_51_321 ();
 sg13g2_decap_4 FILLER_51_328 ();
 sg13g2_fill_1 FILLER_51_332 ();
 sg13g2_fill_2 FILLER_51_338 ();
 sg13g2_decap_8 FILLER_51_397 ();
 sg13g2_decap_4 FILLER_51_404 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_fill_2 FILLER_52_28 ();
 sg13g2_fill_1 FILLER_52_30 ();
 sg13g2_decap_8 FILLER_52_57 ();
 sg13g2_fill_2 FILLER_52_64 ();
 sg13g2_fill_1 FILLER_52_66 ();
 sg13g2_decap_4 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_86 ();
 sg13g2_decap_8 FILLER_52_93 ();
 sg13g2_decap_4 FILLER_52_103 ();
 sg13g2_fill_1 FILLER_52_133 ();
 sg13g2_fill_1 FILLER_52_151 ();
 sg13g2_fill_2 FILLER_52_185 ();
 sg13g2_fill_1 FILLER_52_202 ();
 sg13g2_fill_2 FILLER_52_217 ();
 sg13g2_fill_1 FILLER_52_219 ();
 sg13g2_fill_1 FILLER_52_228 ();
 sg13g2_fill_2 FILLER_52_244 ();
 sg13g2_decap_4 FILLER_52_302 ();
 sg13g2_fill_2 FILLER_52_306 ();
 sg13g2_fill_1 FILLER_52_313 ();
 sg13g2_decap_8 FILLER_52_322 ();
 sg13g2_decap_8 FILLER_52_329 ();
 sg13g2_decap_8 FILLER_52_336 ();
 sg13g2_decap_8 FILLER_52_343 ();
 sg13g2_fill_1 FILLER_52_350 ();
 sg13g2_fill_2 FILLER_52_381 ();
 sg13g2_decap_8 FILLER_52_392 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_fill_2 FILLER_52_406 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_4 FILLER_53_21 ();
 sg13g2_fill_2 FILLER_53_39 ();
 sg13g2_fill_2 FILLER_53_93 ();
 sg13g2_fill_2 FILLER_53_135 ();
 sg13g2_fill_2 FILLER_53_162 ();
 sg13g2_fill_1 FILLER_53_180 ();
 sg13g2_fill_1 FILLER_53_202 ();
 sg13g2_fill_2 FILLER_53_213 ();
 sg13g2_fill_1 FILLER_53_215 ();
 sg13g2_decap_4 FILLER_53_224 ();
 sg13g2_fill_1 FILLER_53_228 ();
 sg13g2_fill_2 FILLER_53_233 ();
 sg13g2_decap_8 FILLER_53_239 ();
 sg13g2_decap_4 FILLER_53_246 ();
 sg13g2_fill_2 FILLER_53_298 ();
 sg13g2_fill_1 FILLER_53_300 ();
 sg13g2_fill_2 FILLER_53_313 ();
 sg13g2_decap_8 FILLER_53_341 ();
 sg13g2_decap_8 FILLER_53_348 ();
 sg13g2_fill_2 FILLER_53_355 ();
 sg13g2_fill_1 FILLER_53_357 ();
 sg13g2_decap_4 FILLER_53_363 ();
 sg13g2_decap_8 FILLER_53_393 ();
 sg13g2_decap_8 FILLER_53_400 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_4 FILLER_54_28 ();
 sg13g2_fill_2 FILLER_54_32 ();
 sg13g2_fill_1 FILLER_54_44 ();
 sg13g2_fill_1 FILLER_54_55 ();
 sg13g2_decap_8 FILLER_54_60 ();
 sg13g2_decap_8 FILLER_54_67 ();
 sg13g2_decap_4 FILLER_54_74 ();
 sg13g2_decap_8 FILLER_54_82 ();
 sg13g2_decap_4 FILLER_54_89 ();
 sg13g2_decap_8 FILLER_54_133 ();
 sg13g2_fill_1 FILLER_54_145 ();
 sg13g2_decap_4 FILLER_54_151 ();
 sg13g2_decap_8 FILLER_54_159 ();
 sg13g2_decap_8 FILLER_54_169 ();
 sg13g2_decap_4 FILLER_54_176 ();
 sg13g2_fill_2 FILLER_54_180 ();
 sg13g2_decap_4 FILLER_54_203 ();
 sg13g2_fill_1 FILLER_54_207 ();
 sg13g2_fill_2 FILLER_54_238 ();
 sg13g2_fill_2 FILLER_54_256 ();
 sg13g2_decap_4 FILLER_54_263 ();
 sg13g2_fill_2 FILLER_54_267 ();
 sg13g2_fill_1 FILLER_54_278 ();
 sg13g2_decap_8 FILLER_54_290 ();
 sg13g2_fill_2 FILLER_54_297 ();
 sg13g2_decap_4 FILLER_54_328 ();
 sg13g2_fill_1 FILLER_54_332 ();
 sg13g2_decap_8 FILLER_54_363 ();
 sg13g2_fill_1 FILLER_54_370 ();
 sg13g2_fill_2 FILLER_54_379 ();
 sg13g2_decap_8 FILLER_54_398 ();
 sg13g2_decap_4 FILLER_54_405 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_4 FILLER_55_14 ();
 sg13g2_fill_2 FILLER_55_18 ();
 sg13g2_decap_8 FILLER_55_46 ();
 sg13g2_decap_8 FILLER_55_53 ();
 sg13g2_decap_8 FILLER_55_60 ();
 sg13g2_fill_2 FILLER_55_86 ();
 sg13g2_decap_8 FILLER_55_97 ();
 sg13g2_decap_8 FILLER_55_108 ();
 sg13g2_fill_2 FILLER_55_115 ();
 sg13g2_decap_8 FILLER_55_125 ();
 sg13g2_decap_8 FILLER_55_132 ();
 sg13g2_fill_2 FILLER_55_139 ();
 sg13g2_decap_8 FILLER_55_149 ();
 sg13g2_decap_4 FILLER_55_156 ();
 sg13g2_fill_1 FILLER_55_160 ();
 sg13g2_decap_8 FILLER_55_179 ();
 sg13g2_decap_4 FILLER_55_186 ();
 sg13g2_decap_8 FILLER_55_194 ();
 sg13g2_decap_8 FILLER_55_201 ();
 sg13g2_decap_8 FILLER_55_208 ();
 sg13g2_fill_1 FILLER_55_215 ();
 sg13g2_decap_8 FILLER_55_265 ();
 sg13g2_decap_8 FILLER_55_272 ();
 sg13g2_fill_1 FILLER_55_279 ();
 sg13g2_decap_4 FILLER_55_284 ();
 sg13g2_fill_1 FILLER_55_288 ();
 sg13g2_decap_4 FILLER_55_369 ();
 sg13g2_fill_2 FILLER_55_373 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_fill_2 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_fill_1 FILLER_56_56 ();
 sg13g2_fill_1 FILLER_56_88 ();
 sg13g2_fill_2 FILLER_56_103 ();
 sg13g2_fill_2 FILLER_56_115 ();
 sg13g2_fill_1 FILLER_56_117 ();
 sg13g2_fill_2 FILLER_56_123 ();
 sg13g2_decap_8 FILLER_56_130 ();
 sg13g2_fill_1 FILLER_56_137 ();
 sg13g2_fill_1 FILLER_56_172 ();
 sg13g2_fill_2 FILLER_56_192 ();
 sg13g2_fill_2 FILLER_56_203 ();
 sg13g2_decap_4 FILLER_56_218 ();
 sg13g2_fill_2 FILLER_56_235 ();
 sg13g2_decap_8 FILLER_56_256 ();
 sg13g2_decap_8 FILLER_56_263 ();
 sg13g2_fill_2 FILLER_56_270 ();
 sg13g2_fill_2 FILLER_56_277 ();
 sg13g2_fill_1 FILLER_56_279 ();
 sg13g2_fill_1 FILLER_56_288 ();
 sg13g2_fill_2 FILLER_56_297 ();
 sg13g2_fill_1 FILLER_56_299 ();
 sg13g2_decap_8 FILLER_56_313 ();
 sg13g2_decap_8 FILLER_56_320 ();
 sg13g2_decap_4 FILLER_56_327 ();
 sg13g2_fill_2 FILLER_56_355 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_7 ();
 sg13g2_fill_1 FILLER_57_9 ();
 sg13g2_fill_2 FILLER_57_101 ();
 sg13g2_fill_2 FILLER_57_134 ();
 sg13g2_fill_2 FILLER_57_189 ();
 sg13g2_fill_1 FILLER_57_191 ();
 sg13g2_decap_8 FILLER_57_223 ();
 sg13g2_decap_8 FILLER_57_230 ();
 sg13g2_decap_8 FILLER_57_241 ();
 sg13g2_fill_2 FILLER_57_248 ();
 sg13g2_fill_1 FILLER_57_250 ();
 sg13g2_fill_1 FILLER_57_268 ();
 sg13g2_decap_8 FILLER_57_295 ();
 sg13g2_decap_8 FILLER_57_302 ();
 sg13g2_decap_8 FILLER_57_309 ();
 sg13g2_decap_8 FILLER_57_316 ();
 sg13g2_decap_4 FILLER_57_323 ();
 sg13g2_fill_2 FILLER_57_327 ();
 sg13g2_decap_4 FILLER_57_334 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_4 FILLER_58_14 ();
 sg13g2_fill_1 FILLER_58_18 ();
 sg13g2_fill_2 FILLER_58_43 ();
 sg13g2_fill_1 FILLER_58_59 ();
 sg13g2_fill_1 FILLER_58_156 ();
 sg13g2_decap_4 FILLER_58_201 ();
 sg13g2_fill_2 FILLER_58_210 ();
 sg13g2_decap_8 FILLER_58_216 ();
 sg13g2_fill_2 FILLER_58_223 ();
 sg13g2_fill_1 FILLER_58_225 ();
 sg13g2_decap_8 FILLER_58_230 ();
 sg13g2_fill_2 FILLER_58_237 ();
 sg13g2_decap_4 FILLER_58_343 ();
 sg13g2_fill_1 FILLER_58_347 ();
 sg13g2_decap_8 FILLER_58_396 ();
 sg13g2_decap_4 FILLER_58_403 ();
 sg13g2_fill_2 FILLER_58_407 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_4 FILLER_59_28 ();
 sg13g2_fill_2 FILLER_59_32 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_54 ();
 sg13g2_decap_8 FILLER_59_61 ();
 sg13g2_decap_8 FILLER_59_68 ();
 sg13g2_fill_2 FILLER_59_85 ();
 sg13g2_fill_1 FILLER_59_87 ();
 sg13g2_decap_8 FILLER_59_96 ();
 sg13g2_decap_8 FILLER_59_103 ();
 sg13g2_decap_4 FILLER_59_110 ();
 sg13g2_fill_2 FILLER_59_114 ();
 sg13g2_fill_1 FILLER_59_140 ();
 sg13g2_decap_8 FILLER_59_169 ();
 sg13g2_fill_2 FILLER_59_176 ();
 sg13g2_fill_1 FILLER_59_178 ();
 sg13g2_fill_2 FILLER_59_184 ();
 sg13g2_fill_1 FILLER_59_196 ();
 sg13g2_decap_4 FILLER_59_205 ();
 sg13g2_fill_1 FILLER_59_209 ();
 sg13g2_fill_2 FILLER_59_227 ();
 sg13g2_fill_1 FILLER_59_229 ();
 sg13g2_decap_4 FILLER_59_241 ();
 sg13g2_fill_2 FILLER_59_281 ();
 sg13g2_fill_1 FILLER_59_283 ();
 sg13g2_fill_2 FILLER_59_295 ();
 sg13g2_decap_8 FILLER_59_333 ();
 sg13g2_decap_8 FILLER_59_340 ();
 sg13g2_decap_4 FILLER_59_347 ();
 sg13g2_decap_8 FILLER_59_355 ();
 sg13g2_fill_1 FILLER_59_362 ();
 sg13g2_decap_8 FILLER_59_372 ();
 sg13g2_decap_4 FILLER_59_379 ();
 sg13g2_decap_8 FILLER_59_387 ();
 sg13g2_decap_8 FILLER_59_394 ();
 sg13g2_decap_8 FILLER_59_401 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_38 ();
 sg13g2_decap_8 FILLER_60_45 ();
 sg13g2_decap_8 FILLER_60_52 ();
 sg13g2_decap_8 FILLER_60_59 ();
 sg13g2_fill_2 FILLER_60_66 ();
 sg13g2_fill_1 FILLER_60_68 ();
 sg13g2_decap_8 FILLER_60_79 ();
 sg13g2_fill_2 FILLER_60_86 ();
 sg13g2_decap_8 FILLER_60_93 ();
 sg13g2_fill_2 FILLER_60_100 ();
 sg13g2_fill_1 FILLER_60_102 ();
 sg13g2_decap_8 FILLER_60_108 ();
 sg13g2_decap_8 FILLER_60_115 ();
 sg13g2_decap_8 FILLER_60_122 ();
 sg13g2_fill_2 FILLER_60_129 ();
 sg13g2_decap_8 FILLER_60_136 ();
 sg13g2_decap_8 FILLER_60_143 ();
 sg13g2_fill_1 FILLER_60_158 ();
 sg13g2_decap_8 FILLER_60_162 ();
 sg13g2_decap_4 FILLER_60_169 ();
 sg13g2_fill_2 FILLER_60_173 ();
 sg13g2_fill_2 FILLER_60_212 ();
 sg13g2_fill_1 FILLER_60_214 ();
 sg13g2_fill_2 FILLER_60_249 ();
 sg13g2_fill_1 FILLER_60_251 ();
 sg13g2_fill_2 FILLER_60_256 ();
 sg13g2_fill_1 FILLER_60_258 ();
 sg13g2_decap_4 FILLER_60_279 ();
 sg13g2_fill_1 FILLER_60_283 ();
 sg13g2_fill_1 FILLER_60_315 ();
 sg13g2_decap_8 FILLER_60_330 ();
 sg13g2_fill_2 FILLER_60_337 ();
 sg13g2_fill_2 FILLER_60_370 ();
 sg13g2_fill_1 FILLER_60_372 ();
 sg13g2_fill_2 FILLER_60_383 ();
 sg13g2_fill_1 FILLER_60_385 ();
 sg13g2_decap_8 FILLER_60_391 ();
 sg13g2_decap_8 FILLER_60_398 ();
 sg13g2_decap_4 FILLER_60_405 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_4 FILLER_61_7 ();
 sg13g2_fill_2 FILLER_61_63 ();
 sg13g2_fill_1 FILLER_61_79 ();
 sg13g2_fill_2 FILLER_61_108 ();
 sg13g2_fill_1 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_139 ();
 sg13g2_decap_8 FILLER_61_146 ();
 sg13g2_decap_8 FILLER_61_153 ();
 sg13g2_decap_4 FILLER_61_160 ();
 sg13g2_fill_1 FILLER_61_164 ();
 sg13g2_fill_1 FILLER_61_183 ();
 sg13g2_fill_2 FILLER_61_210 ();
 sg13g2_fill_1 FILLER_61_212 ();
 sg13g2_decap_4 FILLER_61_246 ();
 sg13g2_fill_1 FILLER_61_250 ();
 sg13g2_decap_8 FILLER_61_257 ();
 sg13g2_decap_8 FILLER_61_264 ();
 sg13g2_decap_8 FILLER_61_271 ();
 sg13g2_decap_8 FILLER_61_278 ();
 sg13g2_decap_8 FILLER_61_285 ();
 sg13g2_decap_8 FILLER_61_301 ();
 sg13g2_decap_4 FILLER_61_308 ();
 sg13g2_fill_2 FILLER_61_312 ();
 sg13g2_decap_8 FILLER_61_320 ();
 sg13g2_decap_4 FILLER_61_327 ();
 sg13g2_fill_1 FILLER_61_331 ();
 sg13g2_decap_4 FILLER_61_353 ();
 sg13g2_decap_4 FILLER_61_404 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_4 FILLER_62_7 ();
 sg13g2_fill_2 FILLER_62_11 ();
 sg13g2_fill_1 FILLER_62_43 ();
 sg13g2_fill_1 FILLER_62_54 ();
 sg13g2_fill_1 FILLER_62_81 ();
 sg13g2_fill_2 FILLER_62_122 ();
 sg13g2_fill_2 FILLER_62_154 ();
 sg13g2_fill_1 FILLER_62_156 ();
 sg13g2_decap_4 FILLER_62_165 ();
 sg13g2_fill_1 FILLER_62_169 ();
 sg13g2_fill_1 FILLER_62_188 ();
 sg13g2_fill_2 FILLER_62_199 ();
 sg13g2_fill_1 FILLER_62_201 ();
 sg13g2_fill_1 FILLER_62_208 ();
 sg13g2_decap_8 FILLER_62_213 ();
 sg13g2_fill_1 FILLER_62_220 ();
 sg13g2_fill_2 FILLER_62_226 ();
 sg13g2_fill_2 FILLER_62_232 ();
 sg13g2_fill_2 FILLER_62_238 ();
 sg13g2_fill_2 FILLER_62_246 ();
 sg13g2_fill_1 FILLER_62_253 ();
 sg13g2_decap_8 FILLER_62_262 ();
 sg13g2_fill_1 FILLER_62_287 ();
 sg13g2_decap_8 FILLER_62_292 ();
 sg13g2_fill_2 FILLER_62_299 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_fill_2 FILLER_63_21 ();
 sg13g2_fill_1 FILLER_63_37 ();
 sg13g2_fill_2 FILLER_63_74 ();
 sg13g2_fill_1 FILLER_63_76 ();
 sg13g2_fill_2 FILLER_63_142 ();
 sg13g2_fill_1 FILLER_63_188 ();
 sg13g2_fill_2 FILLER_63_197 ();
 sg13g2_decap_8 FILLER_63_224 ();
 sg13g2_decap_8 FILLER_63_231 ();
 sg13g2_decap_8 FILLER_63_238 ();
 sg13g2_fill_2 FILLER_63_250 ();
 sg13g2_decap_4 FILLER_63_256 ();
 sg13g2_fill_1 FILLER_63_260 ();
 sg13g2_fill_2 FILLER_63_269 ();
 sg13g2_fill_1 FILLER_63_271 ();
 sg13g2_decap_4 FILLER_63_286 ();
 sg13g2_fill_1 FILLER_63_290 ();
 sg13g2_fill_1 FILLER_63_313 ();
 sg13g2_fill_1 FILLER_63_349 ();
 sg13g2_decap_4 FILLER_63_362 ();
 sg13g2_fill_2 FILLER_63_366 ();
 sg13g2_fill_2 FILLER_63_373 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_4 FILLER_64_35 ();
 sg13g2_fill_2 FILLER_64_39 ();
 sg13g2_decap_8 FILLER_64_59 ();
 sg13g2_fill_2 FILLER_64_66 ();
 sg13g2_fill_2 FILLER_64_83 ();
 sg13g2_fill_1 FILLER_64_85 ();
 sg13g2_fill_1 FILLER_64_91 ();
 sg13g2_fill_1 FILLER_64_127 ();
 sg13g2_decap_4 FILLER_64_142 ();
 sg13g2_fill_1 FILLER_64_146 ();
 sg13g2_decap_8 FILLER_64_167 ();
 sg13g2_fill_2 FILLER_64_174 ();
 sg13g2_fill_2 FILLER_64_206 ();
 sg13g2_decap_8 FILLER_64_214 ();
 sg13g2_fill_1 FILLER_64_221 ();
 sg13g2_fill_2 FILLER_64_234 ();
 sg13g2_fill_1 FILLER_64_236 ();
 sg13g2_fill_1 FILLER_64_259 ();
 sg13g2_fill_2 FILLER_64_275 ();
 sg13g2_fill_1 FILLER_64_277 ();
 sg13g2_decap_8 FILLER_64_339 ();
 sg13g2_decap_8 FILLER_64_346 ();
 sg13g2_decap_8 FILLER_64_353 ();
 sg13g2_decap_8 FILLER_64_360 ();
 sg13g2_decap_8 FILLER_64_367 ();
 sg13g2_fill_1 FILLER_64_379 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_4 FILLER_65_21 ();
 sg13g2_fill_1 FILLER_65_25 ();
 sg13g2_decap_4 FILLER_65_52 ();
 sg13g2_fill_2 FILLER_65_56 ();
 sg13g2_fill_2 FILLER_65_72 ();
 sg13g2_fill_1 FILLER_65_79 ();
 sg13g2_decap_4 FILLER_65_92 ();
 sg13g2_fill_1 FILLER_65_96 ();
 sg13g2_fill_2 FILLER_65_100 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_fill_2 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_132 ();
 sg13g2_decap_8 FILLER_65_139 ();
 sg13g2_decap_8 FILLER_65_146 ();
 sg13g2_decap_8 FILLER_65_153 ();
 sg13g2_decap_4 FILLER_65_160 ();
 sg13g2_fill_1 FILLER_65_164 ();
 sg13g2_fill_2 FILLER_65_173 ();
 sg13g2_fill_1 FILLER_65_175 ();
 sg13g2_decap_8 FILLER_65_180 ();
 sg13g2_fill_2 FILLER_65_187 ();
 sg13g2_fill_2 FILLER_65_201 ();
 sg13g2_fill_2 FILLER_65_214 ();
 sg13g2_fill_1 FILLER_65_227 ();
 sg13g2_decap_8 FILLER_65_330 ();
 sg13g2_decap_8 FILLER_65_337 ();
 sg13g2_decap_4 FILLER_65_344 ();
 sg13g2_fill_2 FILLER_65_348 ();
 sg13g2_fill_1 FILLER_65_360 ();
 sg13g2_decap_8 FILLER_65_365 ();
 sg13g2_decap_8 FILLER_65_372 ();
 sg13g2_decap_4 FILLER_65_379 ();
 sg13g2_decap_4 FILLER_65_405 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_fill_1 FILLER_66_57 ();
 sg13g2_fill_2 FILLER_66_79 ();
 sg13g2_fill_1 FILLER_66_86 ();
 sg13g2_fill_1 FILLER_66_100 ();
 sg13g2_decap_8 FILLER_66_104 ();
 sg13g2_decap_8 FILLER_66_111 ();
 sg13g2_decap_4 FILLER_66_118 ();
 sg13g2_fill_1 FILLER_66_122 ();
 sg13g2_decap_8 FILLER_66_136 ();
 sg13g2_decap_4 FILLER_66_143 ();
 sg13g2_fill_1 FILLER_66_147 ();
 sg13g2_fill_2 FILLER_66_165 ();
 sg13g2_decap_8 FILLER_66_185 ();
 sg13g2_decap_4 FILLER_66_202 ();
 sg13g2_fill_2 FILLER_66_214 ();
 sg13g2_fill_2 FILLER_66_241 ();
 sg13g2_fill_1 FILLER_66_243 ();
 sg13g2_fill_2 FILLER_66_260 ();
 sg13g2_decap_8 FILLER_66_294 ();
 sg13g2_fill_1 FILLER_66_301 ();
 sg13g2_decap_8 FILLER_66_323 ();
 sg13g2_decap_8 FILLER_66_382 ();
 sg13g2_decap_8 FILLER_66_389 ();
 sg13g2_decap_8 FILLER_66_396 ();
 sg13g2_decap_4 FILLER_66_403 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_fill_2 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_48 ();
 sg13g2_decap_8 FILLER_67_55 ();
 sg13g2_decap_4 FILLER_67_62 ();
 sg13g2_fill_1 FILLER_67_66 ();
 sg13g2_fill_1 FILLER_67_88 ();
 sg13g2_decap_4 FILLER_67_110 ();
 sg13g2_fill_2 FILLER_67_145 ();
 sg13g2_fill_2 FILLER_67_171 ();
 sg13g2_decap_4 FILLER_67_190 ();
 sg13g2_fill_2 FILLER_67_194 ();
 sg13g2_decap_8 FILLER_67_222 ();
 sg13g2_decap_4 FILLER_67_240 ();
 sg13g2_fill_1 FILLER_67_244 ();
 sg13g2_fill_1 FILLER_67_259 ();
 sg13g2_fill_1 FILLER_67_276 ();
 sg13g2_fill_1 FILLER_67_289 ();
 sg13g2_fill_2 FILLER_67_295 ();
 sg13g2_fill_1 FILLER_67_297 ();
 sg13g2_decap_8 FILLER_67_320 ();
 sg13g2_fill_1 FILLER_67_327 ();
 sg13g2_fill_2 FILLER_67_338 ();
 sg13g2_fill_1 FILLER_67_340 ();
 sg13g2_decap_8 FILLER_67_345 ();
 sg13g2_fill_1 FILLER_67_352 ();
 sg13g2_decap_4 FILLER_67_405 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_4 FILLER_68_35 ();
 sg13g2_fill_1 FILLER_68_39 ();
 sg13g2_fill_2 FILLER_68_66 ();
 sg13g2_fill_1 FILLER_68_68 ();
 sg13g2_decap_8 FILLER_68_82 ();
 sg13g2_decap_8 FILLER_68_89 ();
 sg13g2_decap_4 FILLER_68_96 ();
 sg13g2_fill_2 FILLER_68_146 ();
 sg13g2_fill_1 FILLER_68_148 ();
 sg13g2_fill_2 FILLER_68_214 ();
 sg13g2_fill_1 FILLER_68_243 ();
 sg13g2_fill_1 FILLER_68_248 ();
 sg13g2_fill_2 FILLER_68_257 ();
 sg13g2_fill_2 FILLER_68_282 ();
 sg13g2_fill_1 FILLER_68_288 ();
 sg13g2_fill_1 FILLER_68_293 ();
 sg13g2_fill_2 FILLER_68_406 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_4 FILLER_69_35 ();
 sg13g2_fill_1 FILLER_69_39 ();
 sg13g2_fill_1 FILLER_69_50 ();
 sg13g2_fill_2 FILLER_69_81 ();
 sg13g2_fill_1 FILLER_69_83 ();
 sg13g2_decap_4 FILLER_69_144 ();
 sg13g2_fill_1 FILLER_69_148 ();
 sg13g2_decap_8 FILLER_69_176 ();
 sg13g2_decap_8 FILLER_69_183 ();
 sg13g2_decap_8 FILLER_69_190 ();
 sg13g2_fill_2 FILLER_69_197 ();
 sg13g2_fill_1 FILLER_69_208 ();
 sg13g2_fill_2 FILLER_69_250 ();
 sg13g2_fill_1 FILLER_69_252 ();
 sg13g2_fill_2 FILLER_69_267 ();
 sg13g2_fill_2 FILLER_69_280 ();
 sg13g2_decap_4 FILLER_69_287 ();
 sg13g2_fill_2 FILLER_69_291 ();
 sg13g2_decap_4 FILLER_69_306 ();
 sg13g2_fill_1 FILLER_69_310 ();
 sg13g2_decap_8 FILLER_69_345 ();
 sg13g2_fill_2 FILLER_69_361 ();
 sg13g2_fill_1 FILLER_69_363 ();
 sg13g2_fill_2 FILLER_69_388 ();
 sg13g2_decap_8 FILLER_69_394 ();
 sg13g2_decap_8 FILLER_69_401 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_4 FILLER_70_28 ();
 sg13g2_fill_2 FILLER_70_32 ();
 sg13g2_fill_2 FILLER_70_60 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_fill_1 FILLER_70_119 ();
 sg13g2_decap_4 FILLER_70_124 ();
 sg13g2_fill_2 FILLER_70_128 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_decap_4 FILLER_70_154 ();
 sg13g2_fill_2 FILLER_70_158 ();
 sg13g2_decap_4 FILLER_70_169 ();
 sg13g2_fill_2 FILLER_70_173 ();
 sg13g2_decap_8 FILLER_70_179 ();
 sg13g2_fill_1 FILLER_70_186 ();
 sg13g2_fill_2 FILLER_70_198 ();
 sg13g2_fill_1 FILLER_70_200 ();
 sg13g2_decap_8 FILLER_70_210 ();
 sg13g2_fill_2 FILLER_70_217 ();
 sg13g2_decap_4 FILLER_70_223 ();
 sg13g2_fill_1 FILLER_70_227 ();
 sg13g2_decap_4 FILLER_70_233 ();
 sg13g2_fill_1 FILLER_70_242 ();
 sg13g2_fill_1 FILLER_70_260 ();
 sg13g2_decap_8 FILLER_70_287 ();
 sg13g2_fill_1 FILLER_70_294 ();
 sg13g2_decap_4 FILLER_70_316 ();
 sg13g2_fill_2 FILLER_70_320 ();
 sg13g2_decap_8 FILLER_70_326 ();
 sg13g2_decap_4 FILLER_70_333 ();
 sg13g2_fill_2 FILLER_70_337 ();
 sg13g2_decap_8 FILLER_70_347 ();
 sg13g2_decap_8 FILLER_70_354 ();
 sg13g2_decap_4 FILLER_70_361 ();
 sg13g2_decap_8 FILLER_70_374 ();
 sg13g2_decap_8 FILLER_70_381 ();
 sg13g2_fill_2 FILLER_70_388 ();
 sg13g2_decap_8 FILLER_70_402 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_4 FILLER_71_28 ();
 sg13g2_fill_2 FILLER_71_32 ();
 sg13g2_fill_1 FILLER_71_44 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_fill_1 FILLER_71_63 ();
 sg13g2_fill_2 FILLER_71_73 ();
 sg13g2_fill_1 FILLER_71_75 ();
 sg13g2_decap_4 FILLER_71_90 ();
 sg13g2_fill_1 FILLER_71_94 ();
 sg13g2_decap_8 FILLER_71_100 ();
 sg13g2_decap_8 FILLER_71_107 ();
 sg13g2_decap_4 FILLER_71_114 ();
 sg13g2_fill_2 FILLER_71_118 ();
 sg13g2_decap_8 FILLER_71_146 ();
 sg13g2_decap_8 FILLER_71_157 ();
 sg13g2_decap_8 FILLER_71_207 ();
 sg13g2_decap_8 FILLER_71_214 ();
 sg13g2_fill_2 FILLER_71_221 ();
 sg13g2_fill_1 FILLER_71_223 ();
 sg13g2_fill_2 FILLER_71_248 ();
 sg13g2_fill_2 FILLER_71_258 ();
 sg13g2_fill_1 FILLER_71_260 ();
 sg13g2_fill_1 FILLER_71_283 ();
 sg13g2_fill_1 FILLER_71_295 ();
 sg13g2_decap_8 FILLER_71_317 ();
 sg13g2_decap_8 FILLER_71_324 ();
 sg13g2_decap_8 FILLER_71_331 ();
 sg13g2_decap_8 FILLER_71_343 ();
 sg13g2_fill_2 FILLER_71_350 ();
 sg13g2_fill_1 FILLER_71_352 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_4 FILLER_72_68 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_fill_2 FILLER_72_105 ();
 sg13g2_fill_2 FILLER_72_116 ();
 sg13g2_fill_1 FILLER_72_191 ();
 sg13g2_fill_2 FILLER_72_218 ();
 sg13g2_fill_2 FILLER_72_242 ();
 sg13g2_fill_2 FILLER_72_255 ();
 sg13g2_fill_2 FILLER_72_267 ();
 sg13g2_fill_2 FILLER_72_298 ();
 sg13g2_fill_2 FILLER_72_317 ();
 sg13g2_fill_1 FILLER_72_319 ();
 sg13g2_decap_4 FILLER_72_334 ();
 sg13g2_fill_2 FILLER_72_338 ();
 sg13g2_fill_2 FILLER_72_375 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_4 FILLER_73_42 ();
 sg13g2_fill_1 FILLER_73_46 ();
 sg13g2_decap_4 FILLER_73_73 ();
 sg13g2_fill_1 FILLER_73_77 ();
 sg13g2_fill_2 FILLER_73_128 ();
 sg13g2_fill_1 FILLER_73_144 ();
 sg13g2_fill_1 FILLER_73_182 ();
 sg13g2_fill_1 FILLER_73_209 ();
 sg13g2_fill_1 FILLER_73_253 ();
 sg13g2_decap_4 FILLER_73_262 ();
 sg13g2_decap_4 FILLER_73_272 ();
 sg13g2_fill_1 FILLER_73_276 ();
 sg13g2_decap_4 FILLER_73_280 ();
 sg13g2_fill_2 FILLER_73_310 ();
 sg13g2_fill_1 FILLER_73_312 ();
 sg13g2_fill_1 FILLER_73_380 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_4 FILLER_74_42 ();
 sg13g2_fill_2 FILLER_74_46 ();
 sg13g2_decap_4 FILLER_74_66 ();
 sg13g2_fill_1 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_123 ();
 sg13g2_fill_1 FILLER_74_130 ();
 sg13g2_decap_8 FILLER_74_135 ();
 sg13g2_decap_8 FILLER_74_142 ();
 sg13g2_decap_4 FILLER_74_149 ();
 sg13g2_decap_4 FILLER_74_165 ();
 sg13g2_fill_1 FILLER_74_178 ();
 sg13g2_decap_4 FILLER_74_210 ();
 sg13g2_fill_2 FILLER_74_219 ();
 sg13g2_fill_1 FILLER_74_221 ();
 sg13g2_fill_1 FILLER_74_226 ();
 sg13g2_fill_2 FILLER_74_245 ();
 sg13g2_fill_1 FILLER_74_289 ();
 sg13g2_fill_1 FILLER_74_293 ();
 sg13g2_decap_4 FILLER_74_302 ();
 sg13g2_fill_2 FILLER_74_306 ();
 sg13g2_decap_4 FILLER_74_334 ();
 sg13g2_fill_2 FILLER_74_348 ();
 sg13g2_decap_4 FILLER_74_376 ();
 sg13g2_fill_1 FILLER_74_380 ();
 sg13g2_decap_4 FILLER_74_403 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_4 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_fill_2 FILLER_75_80 ();
 sg13g2_fill_1 FILLER_75_82 ();
 sg13g2_decap_8 FILLER_75_87 ();
 sg13g2_decap_8 FILLER_75_94 ();
 sg13g2_decap_4 FILLER_75_101 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_4 FILLER_75_147 ();
 sg13g2_fill_2 FILLER_75_151 ();
 sg13g2_decap_8 FILLER_75_157 ();
 sg13g2_decap_8 FILLER_75_164 ();
 sg13g2_fill_1 FILLER_75_176 ();
 sg13g2_decap_8 FILLER_75_187 ();
 sg13g2_decap_8 FILLER_75_194 ();
 sg13g2_fill_1 FILLER_75_201 ();
 sg13g2_decap_8 FILLER_75_206 ();
 sg13g2_fill_2 FILLER_75_213 ();
 sg13g2_fill_1 FILLER_75_215 ();
 sg13g2_fill_2 FILLER_75_225 ();
 sg13g2_fill_2 FILLER_75_280 ();
 sg13g2_decap_8 FILLER_75_291 ();
 sg13g2_decap_8 FILLER_75_298 ();
 sg13g2_decap_8 FILLER_75_305 ();
 sg13g2_fill_2 FILLER_75_312 ();
 sg13g2_decap_4 FILLER_75_328 ();
 sg13g2_fill_1 FILLER_75_332 ();
 sg13g2_decap_8 FILLER_75_355 ();
 sg13g2_fill_2 FILLER_75_362 ();
 sg13g2_decap_8 FILLER_75_368 ();
 sg13g2_decap_8 FILLER_75_375 ();
 sg13g2_fill_2 FILLER_75_386 ();
 sg13g2_fill_1 FILLER_75_393 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_fill_1 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_66 ();
 sg13g2_decap_4 FILLER_76_73 ();
 sg13g2_fill_2 FILLER_76_77 ();
 sg13g2_fill_2 FILLER_76_83 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_4 FILLER_76_112 ();
 sg13g2_fill_2 FILLER_76_116 ();
 sg13g2_fill_2 FILLER_76_128 ();
 sg13g2_decap_8 FILLER_76_134 ();
 sg13g2_fill_2 FILLER_76_141 ();
 sg13g2_fill_2 FILLER_76_192 ();
 sg13g2_decap_8 FILLER_76_283 ();
 sg13g2_decap_8 FILLER_76_290 ();
 sg13g2_fill_2 FILLER_76_297 ();
 sg13g2_decap_8 FILLER_76_314 ();
 sg13g2_decap_4 FILLER_76_321 ();
 sg13g2_fill_1 FILLER_76_325 ();
 sg13g2_fill_2 FILLER_76_331 ();
 sg13g2_decap_8 FILLER_76_352 ();
 sg13g2_decap_4 FILLER_76_359 ();
 sg13g2_decap_8 FILLER_76_368 ();
 sg13g2_fill_1 FILLER_76_375 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_4 FILLER_77_42 ();
 sg13g2_fill_2 FILLER_77_66 ();
 sg13g2_fill_1 FILLER_77_98 ();
 sg13g2_decap_4 FILLER_77_145 ();
 sg13g2_fill_2 FILLER_77_157 ();
 sg13g2_fill_1 FILLER_77_235 ();
 sg13g2_fill_2 FILLER_77_267 ();
 sg13g2_fill_1 FILLER_77_291 ();
 sg13g2_fill_1 FILLER_77_344 ();
 sg13g2_fill_1 FILLER_77_371 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_fill_1 FILLER_78_42 ();
 sg13g2_decap_4 FILLER_78_147 ();
 sg13g2_fill_2 FILLER_78_177 ();
 sg13g2_fill_1 FILLER_78_210 ();
 sg13g2_fill_1 FILLER_78_242 ();
 sg13g2_fill_1 FILLER_78_283 ();
 sg13g2_fill_2 FILLER_78_289 ();
 sg13g2_fill_1 FILLER_78_291 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_fill_2 FILLER_79_49 ();
 sg13g2_decap_4 FILLER_79_103 ();
 sg13g2_fill_1 FILLER_79_107 ();
 sg13g2_fill_1 FILLER_79_170 ();
 sg13g2_decap_8 FILLER_79_208 ();
 sg13g2_fill_1 FILLER_79_215 ();
 sg13g2_fill_1 FILLER_79_230 ();
 sg13g2_fill_2 FILLER_79_302 ();
 sg13g2_fill_2 FILLER_79_314 ();
 sg13g2_fill_1 FILLER_79_316 ();
 sg13g2_fill_2 FILLER_79_343 ();
 sg13g2_fill_1 FILLER_79_345 ();
 sg13g2_fill_2 FILLER_79_380 ();
 sg13g2_fill_1 FILLER_79_382 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_fill_2 FILLER_80_63 ();
 sg13g2_fill_1 FILLER_80_65 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_decap_8 FILLER_80_77 ();
 sg13g2_fill_2 FILLER_80_84 ();
 sg13g2_fill_1 FILLER_80_86 ();
 sg13g2_fill_1 FILLER_80_91 ();
 sg13g2_decap_8 FILLER_80_102 ();
 sg13g2_decap_8 FILLER_80_109 ();
 sg13g2_fill_2 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_126 ();
 sg13g2_fill_2 FILLER_80_130 ();
 sg13g2_decap_8 FILLER_80_136 ();
 sg13g2_decap_8 FILLER_80_143 ();
 sg13g2_decap_4 FILLER_80_150 ();
 sg13g2_fill_1 FILLER_80_154 ();
 sg13g2_fill_2 FILLER_80_159 ();
 sg13g2_fill_1 FILLER_80_161 ();
 sg13g2_decap_8 FILLER_80_166 ();
 sg13g2_fill_1 FILLER_80_178 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_fill_2 FILLER_80_226 ();
 sg13g2_fill_1 FILLER_80_228 ();
 sg13g2_decap_4 FILLER_80_238 ();
 sg13g2_fill_2 FILLER_80_246 ();
 sg13g2_fill_2 FILLER_80_252 ();
 sg13g2_fill_2 FILLER_80_267 ();
 sg13g2_fill_2 FILLER_80_277 ();
 sg13g2_fill_1 FILLER_80_279 ();
 sg13g2_fill_1 FILLER_80_293 ();
 sg13g2_fill_2 FILLER_80_323 ();
 sg13g2_fill_1 FILLER_80_325 ();
 sg13g2_decap_8 FILLER_80_395 ();
 sg13g2_decap_8 FILLER_80_402 ();
endmodule

module tt_um_faramire_rotary_ring_wrapper (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire clknet_0_clk;
 wire \ctr1.intensity_out[0] ;
 wire \ctr1.intensity_out[1] ;
 wire \ctr1.intensity_out[3] ;
 wire \ctr1.intensity_out[5] ;
 wire \ctr1.inverted ;
 wire \ctr1.led_binary[0] ;
 wire \ctr1.led_binary[1] ;
 wire \ctr1.led_binary[2] ;
 wire \ctr1.led_binary[3] ;
 wire \ctr1.led_mask_i[0] ;
 wire \ctr1.led_mask_i[10] ;
 wire \ctr1.led_mask_i[11] ;
 wire \ctr1.led_mask_i[1] ;
 wire \ctr1.led_mask_i[2] ;
 wire \ctr1.led_mask_i[3] ;
 wire \ctr1.led_mask_i[4] ;
 wire \ctr1.led_mask_i[5] ;
 wire \ctr1.led_mask_i[6] ;
 wire \ctr1.led_mask_i[7] ;
 wire \ctr1.led_mask_i[8] ;
 wire \ctr1.led_mask_i[9] ;
 wire \ctr1.rot_dn ;
 wire \ctr1.rot_up ;
 wire \leddriv1.byte_pos[0] ;
 wire \leddriv1.byte_pos[1] ;
 wire \leddriv1.byte_pos[2] ;
 wire \leddriv1.grb_pos[0] ;
 wire \leddriv1.grb_pos[1] ;
 wire \leddriv1.led_dout ;
 wire \leddriv1.led_pos[0] ;
 wire \leddriv1.led_pos[1] ;
 wire \leddriv1.led_pos[2] ;
 wire \leddriv1.led_pos[3] ;
 wire \leddriv1.reg_colour[0] ;
 wire \leddriv1.reg_colour[1] ;
 wire \leddriv1.reg_colour[2] ;
 wire \leddriv1.reg_intensity[0] ;
 wire \leddriv1.reg_intensity[1] ;
 wire \leddriv1.reg_intensity[3] ;
 wire \leddriv1.reg_intensity[5] ;
 wire \leddriv1.reg_led_mask[0] ;
 wire \leddriv1.reg_led_mask[10] ;
 wire \leddriv1.reg_led_mask[11] ;
 wire \leddriv1.reg_led_mask[1] ;
 wire \leddriv1.reg_led_mask[2] ;
 wire \leddriv1.reg_led_mask[3] ;
 wire \leddriv1.reg_led_mask[4] ;
 wire \leddriv1.reg_led_mask[5] ;
 wire \leddriv1.reg_led_mask[6] ;
 wire \leddriv1.reg_led_mask[7] ;
 wire \leddriv1.reg_led_mask[8] ;
 wire \leddriv1.reg_led_mask[9] ;
 wire \leddriv1.rs_counter[0] ;
 wire \leddriv1.rs_counter[10] ;
 wire \leddriv1.rs_counter[1] ;
 wire \leddriv1.rs_counter[2] ;
 wire \leddriv1.rs_counter[3] ;
 wire \leddriv1.rs_counter[4] ;
 wire \leddriv1.rs_counter[5] ;
 wire \leddriv1.rs_counter[6] ;
 wire \leddriv1.rs_counter[7] ;
 wire \leddriv1.rs_counter[8] ;
 wire \leddriv1.rs_counter[9] ;
 wire \leddriv1.skip_calc ;
 wire \leddriv1.state[0] ;
 wire \leddriv1.state[1] ;
 wire \leddriv1.state[2] ;
 wire \leddriv1.state[3] ;
 wire \leddriv1.th_counter[0] ;
 wire \leddriv1.th_counter[1] ;
 wire \leddriv1.th_counter[2] ;
 wire \leddriv1.th_counter[3] ;
 wire \leddriv1.th_counter[4] ;
 wire \leddriv1.th_counter[5] ;
 wire \leddriv1.tl_counter[0] ;
 wire \leddriv1.tl_counter[1] ;
 wire \leddriv1.tl_counter[2] ;
 wire \leddriv1.tl_counter[3] ;
 wire \leddriv1.tl_counter[4] ;
 wire \leddriv1.tl_counter[5] ;
 wire \leddriv1.tl_max[1] ;
 wire \rdec1.dn_detected ;
 wire \rdec1.pause_counter[0] ;
 wire \rdec1.pause_counter[10] ;
 wire \rdec1.pause_counter[11] ;
 wire \rdec1.pause_counter[12] ;
 wire \rdec1.pause_counter[13] ;
 wire \rdec1.pause_counter[14] ;
 wire \rdec1.pause_counter[1] ;
 wire \rdec1.pause_counter[2] ;
 wire \rdec1.pause_counter[3] ;
 wire \rdec1.pause_counter[4] ;
 wire \rdec1.pause_counter[5] ;
 wire \rdec1.pause_counter[6] ;
 wire \rdec1.pause_counter[7] ;
 wire \rdec1.pause_counter[8] ;
 wire \rdec1.pause_counter[9] ;
 wire \rdec1.state[0] ;
 wire \rdec1.state[1] ;
 wire \rdec1.state[2] ;
 wire \rdec1.state[3] ;
 wire \rdec1.up_detected ;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;

 sg13g2_inv_1 _0644_ (.Y(_0118_),
    .A(\leddriv1.state[1] ));
 sg13g2_inv_1 _0645_ (.Y(_0119_),
    .A(net230));
 sg13g2_inv_1 _0646_ (.Y(_0120_),
    .A(\ctr1.rot_up ));
 sg13g2_inv_1 _0647_ (.Y(_0121_),
    .A(net172));
 sg13g2_inv_1 _0648_ (.Y(_0122_),
    .A(net248));
 sg13g2_inv_1 _0649_ (.Y(_0123_),
    .A(net222));
 sg13g2_inv_1 _0650_ (.Y(_0124_),
    .A(net232));
 sg13g2_inv_1 _0651_ (.Y(_0125_),
    .A(net215));
 sg13g2_inv_1 _0652_ (.Y(_0126_),
    .A(net307));
 sg13g2_inv_1 _0653_ (.Y(_0127_),
    .A(\leddriv1.led_pos[3] ));
 sg13g2_inv_1 _0654_ (.Y(_0128_),
    .A(net275));
 sg13g2_inv_1 _0655_ (.Y(_0129_),
    .A(\leddriv1.byte_pos[0] ));
 sg13g2_inv_1 _0656_ (.Y(_0130_),
    .A(\leddriv1.tl_counter[0] ));
 sg13g2_inv_1 _0657_ (.Y(_0131_),
    .A(net266));
 sg13g2_inv_1 _0658_ (.Y(_0132_),
    .A(net309));
 sg13g2_inv_1 _0659_ (.Y(_0133_),
    .A(net330));
 sg13g2_inv_1 _0660_ (.Y(_0134_),
    .A(net177));
 sg13g2_inv_1 _0661_ (.Y(_0135_),
    .A(\leddriv1.th_counter[3] ));
 sg13g2_inv_1 _0662_ (.Y(_0136_),
    .A(net204));
 sg13g2_inv_1 _0663_ (.Y(_0137_),
    .A(net249));
 sg13g2_inv_1 _0664_ (.Y(_0138_),
    .A(net306));
 sg13g2_inv_1 _0665_ (.Y(_0139_),
    .A(net251));
 sg13g2_inv_1 _0666_ (.Y(_0140_),
    .A(net256));
 sg13g2_inv_1 _0667_ (.Y(_0141_),
    .A(net319));
 sg13g2_inv_1 _0668_ (.Y(_0142_),
    .A(net246));
 sg13g2_inv_1 _0669_ (.Y(_0143_),
    .A(net210));
 sg13g2_inv_1 _0670_ (.Y(_0144_),
    .A(net218));
 sg13g2_inv_1 _0671_ (.Y(_0145_),
    .A(net315));
 sg13g2_inv_1 _0672_ (.Y(_0146_),
    .A(\rdec1.pause_counter[14] ));
 sg13g2_inv_1 _0673_ (.Y(_0147_),
    .A(net2));
 sg13g2_nand2_1 _0674_ (.Y(_0148_),
    .A(net115),
    .B(\leddriv1.state[0] ));
 sg13g2_nor2b_1 _0675_ (.A(\leddriv1.tl_counter[1] ),
    .B_N(\leddriv1.tl_max[1] ),
    .Y(_0149_));
 sg13g2_nand4_1 _0676_ (.B(_0132_),
    .C(_0133_),
    .A(_0131_),
    .Y(_0150_),
    .D(_0149_));
 sg13g2_nand3_1 _0677_ (.B(net233),
    .C(_0150_),
    .A(net116),
    .Y(_0151_));
 sg13g2_or3_1 _0678_ (.A(\leddriv1.th_counter[3] ),
    .B(\leddriv1.th_counter[2] ),
    .C(\leddriv1.th_counter[1] ),
    .X(_0152_));
 sg13g2_a21oi_1 _0679_ (.A1(net177),
    .A2(_0152_),
    .Y(_0153_),
    .B1(net176));
 sg13g2_nand2b_1 _0680_ (.Y(_0154_),
    .B(\leddriv1.state[1] ),
    .A_N(_0153_));
 sg13g2_nor2_1 _0681_ (.A(_0151_),
    .B(_0154_),
    .Y(_0155_));
 sg13g2_or2_1 _0682_ (.X(_0156_),
    .B(net297),
    .A(_0151_));
 sg13g2_o21ai_1 _0683_ (.B1(net100),
    .Y(_0003_),
    .A1(net262),
    .A2(_0156_));
 sg13g2_nand4_1 _0684_ (.B(net251),
    .C(net228),
    .A(\leddriv1.rs_counter[7] ),
    .Y(_0157_),
    .D(net258));
 sg13g2_o21ai_1 _0685_ (.B1(net256),
    .Y(_0158_),
    .A1(\leddriv1.rs_counter[5] ),
    .A2(\leddriv1.rs_counter[4] ));
 sg13g2_nor2_2 _0686_ (.A(_0157_),
    .B(_0158_),
    .Y(_0159_));
 sg13g2_nand2_1 _0687_ (.Y(_0160_),
    .A(net281),
    .B(net116));
 sg13g2_nor2_2 _0688_ (.A(_0159_),
    .B(_0160_),
    .Y(_0161_));
 sg13g2_a21o_1 _0689_ (.A2(_0155_),
    .A1(net262),
    .B1(_0161_),
    .X(_0004_));
 sg13g2_nand2_1 _0690_ (.Y(_0162_),
    .A(net281),
    .B(_0159_));
 sg13g2_nand2_1 _0691_ (.Y(_0001_),
    .A(net116),
    .B(net282));
 sg13g2_nand2_1 _0692_ (.Y(_0163_),
    .A(\rdec1.pause_counter[0] ),
    .B(net238));
 sg13g2_nor2_1 _0693_ (.A(_0141_),
    .B(_0163_),
    .Y(_0164_));
 sg13g2_and4_1 _0694_ (.A(\rdec1.pause_counter[0] ),
    .B(net238),
    .C(net192),
    .D(\rdec1.pause_counter[2] ),
    .X(_0165_));
 sg13g2_nand2_1 _0695_ (.Y(_0166_),
    .A(net268),
    .B(_0165_));
 sg13g2_nand4_1 _0696_ (.B(_0142_),
    .C(\rdec1.pause_counter[4] ),
    .A(net107),
    .Y(_0167_),
    .D(_0165_));
 sg13g2_nor4_1 _0697_ (.A(_0145_),
    .B(\rdec1.pause_counter[13] ),
    .C(\rdec1.pause_counter[12] ),
    .D(_0146_),
    .Y(_0168_));
 sg13g2_and2_1 _0698_ (.A(\rdec1.pause_counter[10] ),
    .B(\rdec1.pause_counter[11] ),
    .X(_0169_));
 sg13g2_nand2_1 _0699_ (.Y(_0170_),
    .A(\rdec1.pause_counter[10] ),
    .B(\rdec1.pause_counter[11] ));
 sg13g2_nand2b_1 _0700_ (.Y(_0171_),
    .B(net115),
    .A_N(\rdec1.pause_counter[7] ));
 sg13g2_nor4_1 _0701_ (.A(net226),
    .B(net218),
    .C(_0170_),
    .D(_0171_),
    .Y(_0172_));
 sg13g2_nand3b_1 _0702_ (.B(_0168_),
    .C(_0172_),
    .Y(_0173_),
    .A_N(_0167_));
 sg13g2_nand2_1 _0703_ (.Y(_0174_),
    .A(net115),
    .B(_0173_));
 sg13g2_and3_2 _0704_ (.X(_0175_),
    .A(net108),
    .B(net115),
    .C(_0173_));
 sg13g2_nand3_1 _0705_ (.B(net115),
    .C(_0173_),
    .A(net107),
    .Y(_0176_));
 sg13g2_a21o_1 _0706_ (.A2(net301),
    .A1(net115),
    .B1(_0175_),
    .X(_0006_));
 sg13g2_nand2_1 _0707_ (.Y(_0177_),
    .A(net3),
    .B(net2));
 sg13g2_nand3_1 _0708_ (.B(net260),
    .C(_0177_),
    .A(net1),
    .Y(_0178_));
 sg13g2_nand2_1 _0709_ (.Y(_0007_),
    .A(_0173_),
    .B(_0178_));
 sg13g2_a21oi_1 _0710_ (.A1(net233),
    .A2(_0150_),
    .Y(_0179_),
    .B1(_0118_));
 sg13g2_and2_1 _0711_ (.A(net114),
    .B(_0179_),
    .X(_0180_));
 sg13g2_nand2_1 _0712_ (.Y(_0181_),
    .A(net114),
    .B(_0179_));
 sg13g2_nand2_1 _0713_ (.Y(_0182_),
    .A(\leddriv1.state[1] ),
    .B(_0153_));
 sg13g2_nor2_2 _0714_ (.A(_0151_),
    .B(_0182_),
    .Y(_0183_));
 sg13g2_nand2_1 _0715_ (.Y(_0184_),
    .A(net106),
    .B(net116));
 sg13g2_nor2_1 _0716_ (.A(_0180_),
    .B(_0183_),
    .Y(_0185_));
 sg13g2_nand2_1 _0717_ (.Y(_0002_),
    .A(_0184_),
    .B(_0185_));
 sg13g2_a21oi_1 _0718_ (.A1(net3),
    .A2(net260),
    .Y(_0186_),
    .B1(net274));
 sg13g2_o21ai_1 _0719_ (.B1(net117),
    .Y(_0005_),
    .A1(_0147_),
    .A2(_0186_));
 sg13g2_nand3_1 _0720_ (.B(_0147_),
    .C(net274),
    .A(net117),
    .Y(_0187_));
 sg13g2_inv_1 _0721_ (.Y(_0000_),
    .A(_0187_));
 sg13g2_nor2_1 _0722_ (.A(\ctr1.led_mask_i[5] ),
    .B(\ctr1.led_mask_i[4] ),
    .Y(_0188_));
 sg13g2_nor3_2 _0723_ (.A(\ctr1.led_mask_i[7] ),
    .B(\ctr1.led_mask_i[5] ),
    .C(\ctr1.led_mask_i[4] ),
    .Y(_0189_));
 sg13g2_nor2_1 _0724_ (.A(\ctr1.led_mask_i[6] ),
    .B(\ctr1.led_mask_i[2] ),
    .Y(_0190_));
 sg13g2_nor2_1 _0725_ (.A(\ctr1.led_mask_i[1] ),
    .B(\ctr1.led_mask_i[0] ),
    .Y(_0191_));
 sg13g2_nor2b_1 _0726_ (.A(net298),
    .B_N(_0189_),
    .Y(_0192_));
 sg13g2_nand2b_1 _0727_ (.Y(_0193_),
    .B(_0189_),
    .A_N(\ctr1.led_mask_i[6] ));
 sg13g2_nand4_1 _0728_ (.B(_0189_),
    .C(_0190_),
    .A(\ctr1.led_mask_i[3] ),
    .Y(_0194_),
    .D(_0191_));
 sg13g2_nor3_2 _0729_ (.A(\ctr1.led_mask_i[3] ),
    .B(\ctr1.led_mask_i[1] ),
    .C(\ctr1.led_mask_i[0] ),
    .Y(_0195_));
 sg13g2_nand2_1 _0730_ (.Y(_0196_),
    .A(_0190_),
    .B(_0195_));
 sg13g2_nand4_1 _0731_ (.B(_0188_),
    .C(_0190_),
    .A(\ctr1.led_mask_i[7] ),
    .Y(_0197_),
    .D(_0195_));
 sg13g2_xor2_1 _0732_ (.B(\ctr1.led_mask_i[2] ),
    .A(\ctr1.led_mask_i[6] ),
    .X(_0198_));
 sg13g2_nand3_1 _0733_ (.B(_0195_),
    .C(_0198_),
    .A(_0189_),
    .Y(_0199_));
 sg13g2_nor2_1 _0734_ (.A(\ctr1.led_mask_i[11] ),
    .B(\ctr1.led_mask_i[10] ),
    .Y(_0200_));
 sg13g2_nand4_1 _0735_ (.B(_0197_),
    .C(_0199_),
    .A(_0194_),
    .Y(_0201_),
    .D(_0200_));
 sg13g2_or2_1 _0736_ (.X(_0202_),
    .B(\ctr1.led_mask_i[8] ),
    .A(\ctr1.led_mask_i[9] ));
 sg13g2_a21oi_1 _0737_ (.A1(\ctr1.led_mask_i[11] ),
    .A2(\ctr1.led_mask_i[10] ),
    .Y(_0203_),
    .B1(_0202_));
 sg13g2_nand3_1 _0738_ (.B(_0190_),
    .C(_0195_),
    .A(_0189_),
    .Y(_0204_));
 sg13g2_nand2b_1 _0739_ (.Y(_0205_),
    .B(_0204_),
    .A_N(_0200_));
 sg13g2_nand3_1 _0740_ (.B(_0203_),
    .C(_0205_),
    .A(_0201_),
    .Y(_0206_));
 sg13g2_or3_2 _0741_ (.A(\ctr1.led_mask_i[11] ),
    .B(\ctr1.led_mask_i[10] ),
    .C(_0202_),
    .X(_0207_));
 sg13g2_inv_1 _0742_ (.Y(_0208_),
    .A(_0207_));
 sg13g2_nand2b_1 _0743_ (.Y(_0209_),
    .B(\ctr1.led_mask_i[5] ),
    .A_N(\ctr1.led_mask_i[4] ));
 sg13g2_xnor2_1 _0744_ (.Y(_0210_),
    .A(\ctr1.led_mask_i[5] ),
    .B(\ctr1.led_mask_i[4] ));
 sg13g2_or4_1 _0745_ (.A(\ctr1.led_mask_i[7] ),
    .B(_0196_),
    .C(_0207_),
    .D(_0210_),
    .X(_0211_));
 sg13g2_nand2_1 _0746_ (.Y(_0212_),
    .A(\ctr1.led_mask_i[1] ),
    .B(\ctr1.led_mask_i[0] ));
 sg13g2_nor2_1 _0747_ (.A(\ctr1.led_mask_i[3] ),
    .B(\ctr1.led_mask_i[2] ),
    .Y(_0213_));
 sg13g2_nand2_1 _0748_ (.Y(_0214_),
    .A(\ctr1.led_mask_i[9] ),
    .B(\ctr1.led_mask_i[8] ));
 sg13g2_nand3_1 _0749_ (.B(_0202_),
    .C(_0214_),
    .A(_0200_),
    .Y(_0215_));
 sg13g2_nor2_1 _0750_ (.A(_0204_),
    .B(_0215_),
    .Y(_0216_));
 sg13g2_nand2_1 _0751_ (.Y(_0217_),
    .A(_0212_),
    .B(_0213_));
 sg13g2_nor4_1 _0752_ (.A(_0191_),
    .B(_0193_),
    .C(_0207_),
    .D(_0217_),
    .Y(_0218_));
 sg13g2_nor2_1 _0753_ (.A(_0216_),
    .B(_0218_),
    .Y(_0219_));
 sg13g2_nand3_1 _0754_ (.B(_0211_),
    .C(_0219_),
    .A(_0206_),
    .Y(_0220_));
 sg13g2_o21ai_1 _0755_ (.B1(net112),
    .Y(_0221_),
    .A1(net196),
    .A2(_0220_));
 sg13g2_nand2_1 _0756_ (.Y(_0222_),
    .A(\ctr1.led_mask_i[1] ),
    .B(_0213_));
 sg13g2_nor4_1 _0757_ (.A(\ctr1.led_mask_i[0] ),
    .B(_0193_),
    .C(_0207_),
    .D(_0222_),
    .Y(_0223_));
 sg13g2_a21oi_1 _0758_ (.A1(_0194_),
    .A2(_0197_),
    .Y(_0224_),
    .B1(_0207_));
 sg13g2_nor4_1 _0759_ (.A(\ctr1.led_mask_i[7] ),
    .B(_0196_),
    .C(_0207_),
    .D(_0209_),
    .Y(_0225_));
 sg13g2_xnor2_1 _0760_ (.Y(_0226_),
    .A(\ctr1.led_mask_i[11] ),
    .B(\ctr1.led_mask_i[9] ));
 sg13g2_nor4_1 _0761_ (.A(\ctr1.led_mask_i[10] ),
    .B(\ctr1.led_mask_i[8] ),
    .C(_0204_),
    .D(_0226_),
    .Y(_0227_));
 sg13g2_nor4_1 _0762_ (.A(_0223_),
    .B(_0224_),
    .C(_0225_),
    .D(_0227_),
    .Y(_0228_));
 sg13g2_a21oi_1 _0763_ (.A1(_0220_),
    .A2(_0228_),
    .Y(_0019_),
    .B1(_0221_));
 sg13g2_o21ai_1 _0764_ (.B1(_0206_),
    .Y(_0229_),
    .A1(_0122_),
    .A2(_0220_));
 sg13g2_and2_1 _0765_ (.A(net112),
    .B(_0229_),
    .X(_0020_));
 sg13g2_o21ai_1 _0766_ (.B1(net112),
    .Y(_0230_),
    .A1(net214),
    .A2(_0220_));
 sg13g2_a21oi_1 _0767_ (.A1(_0192_),
    .A2(_0220_),
    .Y(_0021_),
    .B1(_0230_));
 sg13g2_o21ai_1 _0768_ (.B1(net112),
    .Y(_0231_),
    .A1(net179),
    .A2(_0220_));
 sg13g2_a21oi_1 _0769_ (.A1(_0208_),
    .A2(_0220_),
    .Y(_0022_),
    .B1(_0231_));
 sg13g2_or2_1 _0770_ (.X(_0232_),
    .B(\ctr1.rot_dn ),
    .A(\ctr1.rot_up ));
 sg13g2_nand2_1 _0771_ (.Y(_0233_),
    .A(net102),
    .B(\ctr1.led_mask_i[1] ));
 sg13g2_nand3b_1 _0772_ (.B(net93),
    .C(_0233_),
    .Y(_0234_),
    .A_N(\ctr1.led_mask_i[11] ));
 sg13g2_o21ai_1 _0773_ (.B1(_0234_),
    .Y(_0235_),
    .A1(net341),
    .A2(net93));
 sg13g2_nand2_1 _0774_ (.Y(_0023_),
    .A(net114),
    .B(net342));
 sg13g2_nand2_2 _0775_ (.Y(_0236_),
    .A(net102),
    .B(\ctr1.rot_dn ));
 sg13g2_nor2_1 _0776_ (.A(net333),
    .B(net92),
    .Y(_0237_));
 sg13g2_o21ai_1 _0777_ (.B1(net114),
    .Y(_0238_),
    .A1(net102),
    .A2(\ctr1.led_mask_i[0] ));
 sg13g2_nor2_1 _0778_ (.A(\ctr1.led_mask_i[1] ),
    .B(net93),
    .Y(_0239_));
 sg13g2_nor3_1 _0779_ (.A(_0237_),
    .B(_0238_),
    .C(_0239_),
    .Y(_0024_));
 sg13g2_nor2_1 _0780_ (.A(net335),
    .B(_0236_),
    .Y(_0240_));
 sg13g2_o21ai_1 _0781_ (.B1(net111),
    .Y(_0241_),
    .A1(net103),
    .A2(\ctr1.led_mask_i[1] ));
 sg13g2_nor2_1 _0782_ (.A(net333),
    .B(net94),
    .Y(_0242_));
 sg13g2_nor3_1 _0783_ (.A(net336),
    .B(_0241_),
    .C(_0242_),
    .Y(_0025_));
 sg13g2_nor2_1 _0784_ (.A(net338),
    .B(_0236_),
    .Y(_0243_));
 sg13g2_o21ai_1 _0785_ (.B1(net111),
    .Y(_0244_),
    .A1(net103),
    .A2(net333));
 sg13g2_nor2_1 _0786_ (.A(net335),
    .B(net93),
    .Y(_0245_));
 sg13g2_nor3_1 _0787_ (.A(net339),
    .B(_0244_),
    .C(_0245_),
    .Y(_0026_));
 sg13g2_nor2_1 _0788_ (.A(net340),
    .B(net92),
    .Y(_0246_));
 sg13g2_o21ai_1 _0789_ (.B1(net111),
    .Y(_0247_),
    .A1(net103),
    .A2(net335));
 sg13g2_nor2_1 _0790_ (.A(net338),
    .B(net93),
    .Y(_0248_));
 sg13g2_nor3_1 _0791_ (.A(_0246_),
    .B(_0247_),
    .C(_0248_),
    .Y(_0027_));
 sg13g2_nor2_1 _0792_ (.A(net298),
    .B(net92),
    .Y(_0249_));
 sg13g2_o21ai_1 _0793_ (.B1(net111),
    .Y(_0250_),
    .A1(net103),
    .A2(net338));
 sg13g2_nor2_1 _0794_ (.A(net340),
    .B(net94),
    .Y(_0251_));
 sg13g2_nor3_1 _0795_ (.A(_0249_),
    .B(_0250_),
    .C(_0251_),
    .Y(_0028_));
 sg13g2_nor2_1 _0796_ (.A(net325),
    .B(net92),
    .Y(_0252_));
 sg13g2_o21ai_1 _0797_ (.B1(net111),
    .Y(_0253_),
    .A1(net103),
    .A2(net340));
 sg13g2_nor2_1 _0798_ (.A(net298),
    .B(net94),
    .Y(_0254_));
 sg13g2_nor3_1 _0799_ (.A(_0252_),
    .B(_0253_),
    .C(_0254_),
    .Y(_0029_));
 sg13g2_nor2_1 _0800_ (.A(net299),
    .B(_0236_),
    .Y(_0255_));
 sg13g2_o21ai_1 _0801_ (.B1(net111),
    .Y(_0256_),
    .A1(net102),
    .A2(net298));
 sg13g2_nor2_1 _0802_ (.A(net325),
    .B(net94),
    .Y(_0257_));
 sg13g2_nor3_1 _0803_ (.A(_0255_),
    .B(_0256_),
    .C(_0257_),
    .Y(_0030_));
 sg13g2_nor2_1 _0804_ (.A(net323),
    .B(net92),
    .Y(_0258_));
 sg13g2_o21ai_1 _0805_ (.B1(net111),
    .Y(_0259_),
    .A1(net102),
    .A2(\ctr1.led_mask_i[7] ));
 sg13g2_nor2_1 _0806_ (.A(net299),
    .B(net93),
    .Y(_0260_));
 sg13g2_nor3_1 _0807_ (.A(_0258_),
    .B(_0259_),
    .C(_0260_),
    .Y(_0031_));
 sg13g2_nor2_1 _0808_ (.A(net305),
    .B(net92),
    .Y(_0261_));
 sg13g2_o21ai_1 _0809_ (.B1(net114),
    .Y(_0262_),
    .A1(net102),
    .A2(net299));
 sg13g2_nor2_1 _0810_ (.A(net323),
    .B(net93),
    .Y(_0263_));
 sg13g2_nor3_1 _0811_ (.A(_0261_),
    .B(_0262_),
    .C(_0263_),
    .Y(_0032_));
 sg13g2_or2_1 _0812_ (.X(_0264_),
    .B(net93),
    .A(net305));
 sg13g2_o21ai_1 _0813_ (.B1(net114),
    .Y(_0265_),
    .A1(net102),
    .A2(net323));
 sg13g2_o21ai_1 _0814_ (.B1(_0264_),
    .Y(_0266_),
    .A1(net332),
    .A2(net92));
 sg13g2_nor2_1 _0815_ (.A(_0265_),
    .B(_0266_),
    .Y(_0033_));
 sg13g2_o21ai_1 _0816_ (.B1(net92),
    .Y(_0267_),
    .A1(net208),
    .A2(net332));
 sg13g2_o21ai_1 _0817_ (.B1(net114),
    .Y(_0268_),
    .A1(net102),
    .A2(net305));
 sg13g2_nor2_1 _0818_ (.A(_0267_),
    .B(_0268_),
    .Y(_0034_));
 sg13g2_nand2b_1 _0819_ (.Y(_0035_),
    .B(net113),
    .A_N(net196));
 sg13g2_nand2_1 _0820_ (.Y(_0036_),
    .A(_0122_),
    .B(net113));
 sg13g2_nand2b_1 _0821_ (.Y(_0037_),
    .B(net112),
    .A_N(net214));
 sg13g2_nand2b_1 _0822_ (.Y(_0038_),
    .B(net112),
    .A_N(net179));
 sg13g2_nand2b_1 _0823_ (.Y(_0039_),
    .B(net111),
    .A_N(net110));
 sg13g2_o21ai_1 _0824_ (.B1(net117),
    .Y(_0269_),
    .A1(net110),
    .A2(net4));
 sg13g2_a21oi_1 _0825_ (.A1(_0121_),
    .A2(net4),
    .Y(_0040_),
    .B1(_0269_));
 sg13g2_mux2_1 _0826_ (.A0(net3),
    .A1(net220),
    .S(_0187_),
    .X(_0041_));
 sg13g2_nand2_1 _0827_ (.Y(_0270_),
    .A(net201),
    .B(_0187_));
 sg13g2_o21ai_1 _0828_ (.B1(net202),
    .Y(_0042_),
    .A1(net3),
    .A2(_0187_));
 sg13g2_nor2_2 _0829_ (.A(net108),
    .B(\rdec1.state[2] ),
    .Y(_0271_));
 sg13g2_nor2_2 _0830_ (.A(_0174_),
    .B(_0271_),
    .Y(_0272_));
 sg13g2_nand3b_1 _0831_ (.B(net115),
    .C(_0173_),
    .Y(_0273_),
    .A_N(_0271_));
 sg13g2_a22oi_1 _0832_ (.Y(_0274_),
    .B1(net91),
    .B2(\rdec1.pause_counter[0] ),
    .A2(_0175_),
    .A1(net170));
 sg13g2_inv_1 _0833_ (.Y(_0043_),
    .A(net171));
 sg13g2_a21oi_1 _0834_ (.A1(\rdec1.pause_counter[0] ),
    .A2(_0272_),
    .Y(_0275_),
    .B1(net238));
 sg13g2_nor2b_1 _0835_ (.A(net108),
    .B_N(\rdec1.state[2] ),
    .Y(_0276_));
 sg13g2_nor2_1 _0836_ (.A(net107),
    .B(net90),
    .Y(_0277_));
 sg13g2_a21oi_1 _0837_ (.A1(net108),
    .A2(_0163_),
    .Y(_0278_),
    .B1(net91));
 sg13g2_nor2_1 _0838_ (.A(net239),
    .B(_0278_),
    .Y(_0044_));
 sg13g2_nor2b_1 _0839_ (.A(_0164_),
    .B_N(net107),
    .Y(_0279_));
 sg13g2_nor2_1 _0840_ (.A(net91),
    .B(_0279_),
    .Y(_0280_));
 sg13g2_o21ai_1 _0841_ (.B1(_0141_),
    .Y(_0281_),
    .A1(_0163_),
    .A2(net91));
 sg13g2_nor2b_1 _0842_ (.A(_0280_),
    .B_N(net320),
    .Y(_0045_));
 sg13g2_a21oi_1 _0843_ (.A1(_0164_),
    .A2(_0175_),
    .Y(_0282_),
    .B1(net192));
 sg13g2_a21oi_1 _0844_ (.A1(net192),
    .A2(_0280_),
    .Y(_0046_),
    .B1(_0282_));
 sg13g2_a21oi_1 _0845_ (.A1(_0165_),
    .A2(_0272_),
    .Y(_0283_),
    .B1(net268));
 sg13g2_a21oi_1 _0846_ (.A1(net107),
    .A2(_0166_),
    .Y(_0284_),
    .B1(net90));
 sg13g2_nor2_1 _0847_ (.A(net269),
    .B(_0284_),
    .Y(_0047_));
 sg13g2_nand2b_1 _0848_ (.Y(_0285_),
    .B(net246),
    .A_N(_0284_));
 sg13g2_o21ai_1 _0849_ (.B1(_0285_),
    .Y(_0048_),
    .A1(_0167_),
    .A2(net90));
 sg13g2_nor2_1 _0850_ (.A(_0142_),
    .B(_0166_),
    .Y(_0286_));
 sg13g2_nand4_1 _0851_ (.B(net268),
    .C(net226),
    .A(net246),
    .Y(_0287_),
    .D(_0165_));
 sg13g2_nor2_1 _0852_ (.A(_0176_),
    .B(_0287_),
    .Y(_0288_));
 sg13g2_or2_1 _0853_ (.X(_0289_),
    .B(_0288_),
    .A(_0277_));
 sg13g2_a21oi_1 _0854_ (.A1(_0272_),
    .A2(_0286_),
    .Y(_0290_),
    .B1(net226));
 sg13g2_nor2_1 _0855_ (.A(_0289_),
    .B(net227),
    .Y(_0049_));
 sg13g2_nor2_1 _0856_ (.A(net210),
    .B(_0288_),
    .Y(_0291_));
 sg13g2_a21oi_1 _0857_ (.A1(net210),
    .A2(_0289_),
    .Y(_0050_),
    .B1(_0291_));
 sg13g2_nor2_1 _0858_ (.A(_0143_),
    .B(_0287_),
    .Y(_0292_));
 sg13g2_nor3_2 _0859_ (.A(_0143_),
    .B(_0144_),
    .C(_0287_),
    .Y(_0293_));
 sg13g2_nor2b_1 _0860_ (.A(_0293_),
    .B_N(net107),
    .Y(_0294_));
 sg13g2_nor2_1 _0861_ (.A(net90),
    .B(_0294_),
    .Y(_0295_));
 sg13g2_a21oi_1 _0862_ (.A1(_0272_),
    .A2(_0292_),
    .Y(_0296_),
    .B1(net218));
 sg13g2_nor2_1 _0863_ (.A(_0295_),
    .B(net219),
    .Y(_0051_));
 sg13g2_nand3_1 _0864_ (.B(_0175_),
    .C(_0293_),
    .A(_0145_),
    .Y(_0297_));
 sg13g2_o21ai_1 _0865_ (.B1(_0297_),
    .Y(_0052_),
    .A1(_0145_),
    .A2(_0295_));
 sg13g2_nand2_1 _0866_ (.Y(_0298_),
    .A(\rdec1.pause_counter[9] ),
    .B(_0293_));
 sg13g2_nand3_1 _0867_ (.B(net293),
    .C(_0293_),
    .A(\rdec1.pause_counter[9] ),
    .Y(_0299_));
 sg13g2_a21oi_1 _0868_ (.A1(net107),
    .A2(_0299_),
    .Y(_0300_),
    .B1(net90));
 sg13g2_nor2_1 _0869_ (.A(net90),
    .B(_0298_),
    .Y(_0301_));
 sg13g2_nor2_1 _0870_ (.A(net293),
    .B(_0301_),
    .Y(_0302_));
 sg13g2_nor2_1 _0871_ (.A(_0300_),
    .B(net294),
    .Y(_0053_));
 sg13g2_nor3_1 _0872_ (.A(net291),
    .B(_0176_),
    .C(_0299_),
    .Y(_0303_));
 sg13g2_nand2b_1 _0873_ (.Y(_0304_),
    .B(net291),
    .A_N(_0300_));
 sg13g2_nand2b_1 _0874_ (.Y(_0054_),
    .B(_0304_),
    .A_N(_0303_));
 sg13g2_nand4_1 _0875_ (.B(net271),
    .C(_0169_),
    .A(\rdec1.pause_counter[9] ),
    .Y(_0305_),
    .D(_0293_));
 sg13g2_a21oi_1 _0876_ (.A1(net107),
    .A2(_0305_),
    .Y(_0306_),
    .B1(net90));
 sg13g2_a21oi_1 _0877_ (.A1(_0169_),
    .A2(_0301_),
    .Y(_0307_),
    .B1(net271));
 sg13g2_nor2_1 _0878_ (.A(_0306_),
    .B(net272),
    .Y(_0055_));
 sg13g2_nor3_1 _0879_ (.A(net286),
    .B(_0176_),
    .C(_0305_),
    .Y(_0308_));
 sg13g2_nand2b_1 _0880_ (.Y(_0309_),
    .B(net286),
    .A_N(_0306_));
 sg13g2_nand2b_1 _0881_ (.Y(_0056_),
    .B(_0309_),
    .A_N(_0308_));
 sg13g2_nand2_1 _0882_ (.Y(_0310_),
    .A(net286),
    .B(net271));
 sg13g2_nor4_1 _0883_ (.A(_0170_),
    .B(net90),
    .C(_0298_),
    .D(_0310_),
    .Y(_0311_));
 sg13g2_xnor2_1 _0884_ (.Y(_0312_),
    .A(net288),
    .B(_0311_));
 sg13g2_nor2_1 _0885_ (.A(_0277_),
    .B(net289),
    .Y(_0057_));
 sg13g2_a22oi_1 _0886_ (.Y(_0313_),
    .B1(_0276_),
    .B2(net220),
    .A2(_0271_),
    .A1(\ctr1.rot_dn ));
 sg13g2_nor2b_1 _0887_ (.A(net221),
    .B_N(net116),
    .Y(_0058_));
 sg13g2_a22oi_1 _0888_ (.Y(_0314_),
    .B1(_0276_),
    .B2(net201),
    .A2(_0271_),
    .A1(net208));
 sg13g2_nor2b_1 _0889_ (.A(net209),
    .B_N(net115),
    .Y(_0059_));
 sg13g2_mux2_1 _0890_ (.A0(net180),
    .A1(\leddriv1.reg_intensity[0] ),
    .S(net101),
    .X(_0060_));
 sg13g2_mux2_1 _0891_ (.A0(net190),
    .A1(\leddriv1.reg_intensity[1] ),
    .S(net101),
    .X(_0061_));
 sg13g2_mux2_1 _0892_ (.A0(net216),
    .A1(\leddriv1.reg_intensity[3] ),
    .S(net100),
    .X(_0062_));
 sg13g2_mux2_1 _0893_ (.A0(net186),
    .A1(\leddriv1.reg_intensity[5] ),
    .S(net100),
    .X(_0063_));
 sg13g2_a21oi_1 _0894_ (.A1(\leddriv1.led_pos[0] ),
    .A2(\leddriv1.reg_led_mask[5] ),
    .Y(_0315_),
    .B1(\leddriv1.led_pos[1] ));
 sg13g2_o21ai_1 _0895_ (.B1(_0315_),
    .Y(_0316_),
    .A1(net104),
    .A2(_0123_));
 sg13g2_nor2b_1 _0896_ (.A(net104),
    .B_N(\leddriv1.led_pos[1] ),
    .Y(_0317_));
 sg13g2_and2_1 _0897_ (.A(net104),
    .B(\leddriv1.led_pos[1] ),
    .X(_0318_));
 sg13g2_nand2_1 _0898_ (.Y(_0319_),
    .A(net104),
    .B(net311));
 sg13g2_a221oi_1 _0899_ (.B2(_0125_),
    .C1(\leddriv1.led_pos[3] ),
    .B1(_0318_),
    .A1(_0124_),
    .Y(_0320_),
    .A2(_0317_));
 sg13g2_a21oi_2 _0900_ (.B1(_0126_),
    .Y(_0321_),
    .A2(_0320_),
    .A1(_0316_));
 sg13g2_mux4_1 _0901_ (.S0(net104),
    .A0(\leddriv1.reg_led_mask[0] ),
    .A1(\leddriv1.reg_led_mask[1] ),
    .A2(\leddriv1.reg_led_mask[2] ),
    .A3(\leddriv1.reg_led_mask[3] ),
    .S1(\leddriv1.led_pos[1] ),
    .X(_0322_));
 sg13g2_or3_1 _0902_ (.A(\leddriv1.led_pos[2] ),
    .B(\leddriv1.led_pos[3] ),
    .C(_0322_),
    .X(_0323_));
 sg13g2_mux4_1 _0903_ (.S0(net104),
    .A0(\leddriv1.reg_led_mask[8] ),
    .A1(\leddriv1.reg_led_mask[9] ),
    .A2(\leddriv1.reg_led_mask[10] ),
    .A3(\leddriv1.reg_led_mask[11] ),
    .S1(\leddriv1.led_pos[1] ),
    .X(_0324_));
 sg13g2_o21ai_1 _0904_ (.B1(_0323_),
    .Y(_0325_),
    .A1(_0127_),
    .A2(_0324_));
 sg13g2_or3_2 _0905_ (.A(_0184_),
    .B(_0321_),
    .C(_0325_),
    .X(_0326_));
 sg13g2_or2_1 _0906_ (.X(_0327_),
    .B(net100),
    .A(net106));
 sg13g2_nor3_2 _0907_ (.A(_0009_),
    .B(_0321_),
    .C(_0325_),
    .Y(_0328_));
 sg13g2_nand2_1 _0908_ (.Y(_0329_),
    .A(\leddriv1.byte_pos[0] ),
    .B(net241));
 sg13g2_nor2_2 _0909_ (.A(_0010_),
    .B(_0329_),
    .Y(_0330_));
 sg13g2_nand2_1 _0910_ (.Y(_0331_),
    .A(\leddriv1.grb_pos[1] ),
    .B(_0330_));
 sg13g2_nand2_1 _0911_ (.Y(_0332_),
    .A(_0126_),
    .B(_0319_));
 sg13g2_nand4_1 _0912_ (.B(\leddriv1.grb_pos[1] ),
    .C(_0330_),
    .A(\leddriv1.led_pos[3] ),
    .Y(_0333_),
    .D(_0332_));
 sg13g2_nor4_2 _0913_ (.A(_0009_),
    .B(_0321_),
    .C(_0325_),
    .Y(_0334_),
    .D(_0333_));
 sg13g2_a21oi_2 _0914_ (.B1(_0334_),
    .Y(_0335_),
    .A2(_0327_),
    .A1(_0326_));
 sg13g2_nor2b_1 _0915_ (.A(_0330_),
    .B_N(\leddriv1.state[2] ),
    .Y(_0336_));
 sg13g2_nand3_1 _0916_ (.B(_0335_),
    .C(_0336_),
    .A(net165),
    .Y(_0337_));
 sg13g2_o21ai_1 _0917_ (.B1(net166),
    .Y(_0064_),
    .A1(_0129_),
    .A2(_0335_));
 sg13g2_a21oi_1 _0918_ (.A1(\leddriv1.byte_pos[0] ),
    .A2(_0335_),
    .Y(_0338_),
    .B1(net241));
 sg13g2_nand2_1 _0919_ (.Y(_0339_),
    .A(net106),
    .B(_0329_));
 sg13g2_a21oi_1 _0920_ (.A1(_0335_),
    .A2(_0339_),
    .Y(_0065_),
    .B1(net242));
 sg13g2_nand2_1 _0921_ (.Y(_0340_),
    .A(_0010_),
    .B(_0329_));
 sg13g2_nand3_1 _0922_ (.B(_0336_),
    .C(_0340_),
    .A(_0335_),
    .Y(_0341_));
 sg13g2_o21ai_1 _0923_ (.B1(_0341_),
    .Y(_0066_),
    .A1(_0128_),
    .A2(_0335_));
 sg13g2_nand2b_1 _0924_ (.Y(_0342_),
    .B(_0328_),
    .A_N(_0330_));
 sg13g2_nand2_1 _0925_ (.Y(_0343_),
    .A(_0335_),
    .B(_0342_));
 sg13g2_nor2_1 _0926_ (.A(_0009_),
    .B(net321),
    .Y(_0344_));
 sg13g2_and2_1 _0927_ (.A(net283),
    .B(_0344_),
    .X(_0345_));
 sg13g2_mux2_1 _0928_ (.A0(net284),
    .A1(\leddriv1.grb_pos[0] ),
    .S(_0343_),
    .X(_0067_));
 sg13g2_and2_1 _0929_ (.A(\leddriv1.grb_pos[0] ),
    .B(_0344_),
    .X(_0346_));
 sg13g2_mux2_1 _0930_ (.A0(_0346_),
    .A1(net321),
    .S(_0343_),
    .X(_0068_));
 sg13g2_a221oi_1 _0931_ (.B2(_0331_),
    .C1(_0334_),
    .B1(_0328_),
    .A1(_0326_),
    .Y(_0347_),
    .A2(_0327_));
 sg13g2_and2_1 _0932_ (.A(net106),
    .B(net313),
    .X(_0348_));
 sg13g2_mux2_1 _0933_ (.A0(net104),
    .A1(_0348_),
    .S(_0347_),
    .X(_0069_));
 sg13g2_a21oi_1 _0934_ (.A1(net104),
    .A2(_0347_),
    .Y(_0349_),
    .B1(net311));
 sg13g2_nand2_1 _0935_ (.Y(_0350_),
    .A(net106),
    .B(_0319_));
 sg13g2_a21oi_1 _0936_ (.A1(_0347_),
    .A2(_0350_),
    .Y(_0070_),
    .B1(net312));
 sg13g2_nand2_1 _0937_ (.Y(_0351_),
    .A(net307),
    .B(_0318_));
 sg13g2_nand4_1 _0938_ (.B(_0332_),
    .C(_0347_),
    .A(net106),
    .Y(_0352_),
    .D(_0351_));
 sg13g2_o21ai_1 _0939_ (.B1(_0352_),
    .Y(_0071_),
    .A1(_0126_),
    .A2(_0347_));
 sg13g2_nand3_1 _0940_ (.B(_0318_),
    .C(_0347_),
    .A(net307),
    .Y(_0353_));
 sg13g2_o21ai_1 _0941_ (.B1(net106),
    .Y(_0354_),
    .A1(_0127_),
    .A2(_0351_));
 sg13g2_a22oi_1 _0942_ (.Y(_0072_),
    .B1(_0354_),
    .B2(_0347_),
    .A2(_0353_),
    .A1(_0127_));
 sg13g2_mux2_1 _0943_ (.A0(\leddriv1.th_counter[0] ),
    .A1(net174),
    .S(_0183_),
    .X(_0073_));
 sg13g2_nand3_1 _0944_ (.B(net327),
    .C(_0183_),
    .A(\leddriv1.th_counter[0] ),
    .Y(_0355_));
 sg13g2_a21o_1 _0945_ (.A2(_0183_),
    .A1(\leddriv1.th_counter[0] ),
    .B1(net327),
    .X(_0356_));
 sg13g2_and2_1 _0946_ (.A(_0355_),
    .B(net328),
    .X(_0074_));
 sg13g2_nand4_1 _0947_ (.B(net236),
    .C(\leddriv1.th_counter[1] ),
    .A(\leddriv1.th_counter[0] ),
    .Y(_0357_),
    .D(_0183_));
 sg13g2_xnor2_1 _0948_ (.Y(_0075_),
    .A(net236),
    .B(_0355_));
 sg13g2_xnor2_1 _0949_ (.Y(_0076_),
    .A(net244),
    .B(_0357_));
 sg13g2_o21ai_1 _0950_ (.B1(_0134_),
    .Y(_0077_),
    .A1(_0135_),
    .A2(_0357_));
 sg13g2_o21ai_1 _0951_ (.B1(net116),
    .Y(_0358_),
    .A1(\leddriv1.state[3] ),
    .A2(\leddriv1.state[0] ));
 sg13g2_a21oi_2 _0952_ (.B1(_0358_),
    .Y(_0359_),
    .A2(_0159_),
    .A1(net105));
 sg13g2_a21o_2 _0953_ (.A2(_0159_),
    .A1(net105),
    .B1(_0358_),
    .X(_0360_));
 sg13g2_a22oi_1 _0954_ (.Y(_0361_),
    .B1(_0360_),
    .B2(\leddriv1.rs_counter[0] ),
    .A2(_0161_),
    .A1(net168));
 sg13g2_inv_1 _0955_ (.Y(_0079_),
    .A(net169));
 sg13g2_nand3_1 _0956_ (.B(net316),
    .C(_0359_),
    .A(\leddriv1.rs_counter[0] ),
    .Y(_0362_));
 sg13g2_nor2_1 _0957_ (.A(net105),
    .B(net100),
    .Y(_0363_));
 sg13g2_a21oi_1 _0958_ (.A1(\leddriv1.rs_counter[0] ),
    .A2(_0359_),
    .Y(_0364_),
    .B1(net316));
 sg13g2_nor2_1 _0959_ (.A(_0363_),
    .B(net317),
    .Y(_0365_));
 sg13g2_and2_1 _0960_ (.A(_0362_),
    .B(_0365_),
    .X(_0080_));
 sg13g2_and3_1 _0961_ (.X(_0366_),
    .A(\leddriv1.rs_counter[0] ),
    .B(\leddriv1.rs_counter[1] ),
    .C(net204));
 sg13g2_nor2b_1 _0962_ (.A(_0366_),
    .B_N(net105),
    .Y(_0367_));
 sg13g2_nor2_1 _0963_ (.A(_0360_),
    .B(_0367_),
    .Y(_0368_));
 sg13g2_a21oi_1 _0964_ (.A1(_0136_),
    .A2(_0362_),
    .Y(_0081_),
    .B1(_0368_));
 sg13g2_nand2_1 _0965_ (.Y(_0369_),
    .A(_0161_),
    .B(_0366_));
 sg13g2_nand2b_1 _0966_ (.Y(_0370_),
    .B(net253),
    .A_N(_0368_));
 sg13g2_o21ai_1 _0967_ (.B1(_0370_),
    .Y(_0082_),
    .A1(net253),
    .A2(_0369_));
 sg13g2_and3_1 _0968_ (.X(_0371_),
    .A(net253),
    .B(net249),
    .C(_0366_));
 sg13g2_inv_1 _0969_ (.Y(_0372_),
    .A(_0371_));
 sg13g2_a21oi_1 _0970_ (.A1(net105),
    .A2(_0372_),
    .Y(_0373_),
    .B1(_0360_));
 sg13g2_nand3_1 _0971_ (.B(_0359_),
    .C(_0366_),
    .A(\leddriv1.rs_counter[3] ),
    .Y(_0374_));
 sg13g2_a21oi_1 _0972_ (.A1(_0137_),
    .A2(_0374_),
    .Y(_0083_),
    .B1(_0373_));
 sg13g2_a21oi_1 _0973_ (.A1(_0161_),
    .A2(_0371_),
    .Y(_0375_),
    .B1(net264));
 sg13g2_a21oi_1 _0974_ (.A1(net264),
    .A2(_0373_),
    .Y(_0084_),
    .B1(_0375_));
 sg13g2_nand3_1 _0975_ (.B(net251),
    .C(_0371_),
    .A(net264),
    .Y(_0376_));
 sg13g2_a21oi_1 _0976_ (.A1(net105),
    .A2(_0376_),
    .Y(_0377_),
    .B1(_0360_));
 sg13g2_nand3_1 _0977_ (.B(_0359_),
    .C(_0371_),
    .A(\leddriv1.rs_counter[5] ),
    .Y(_0378_));
 sg13g2_a21oi_1 _0978_ (.A1(_0139_),
    .A2(_0378_),
    .Y(_0085_),
    .B1(_0377_));
 sg13g2_nand3b_1 _0979_ (.B(_0138_),
    .C(_0161_),
    .Y(_0379_),
    .A_N(_0376_));
 sg13g2_o21ai_1 _0980_ (.B1(_0379_),
    .Y(_0086_),
    .A1(_0138_),
    .A2(_0377_));
 sg13g2_nor2_1 _0981_ (.A(_0138_),
    .B(_0376_),
    .Y(_0380_));
 sg13g2_and2_1 _0982_ (.A(\leddriv1.rs_counter[8] ),
    .B(_0380_),
    .X(_0381_));
 sg13g2_nand2_1 _0983_ (.Y(_0382_),
    .A(net258),
    .B(_0380_));
 sg13g2_a21oi_1 _0984_ (.A1(net105),
    .A2(_0382_),
    .Y(_0383_),
    .B1(_0360_));
 sg13g2_a21oi_1 _0985_ (.A1(_0359_),
    .A2(_0380_),
    .Y(_0384_),
    .B1(net258));
 sg13g2_nor2_1 _0986_ (.A(_0383_),
    .B(net259),
    .Y(_0087_));
 sg13g2_a21oi_1 _0987_ (.A1(_0161_),
    .A2(_0381_),
    .Y(_0385_),
    .B1(net228));
 sg13g2_a21oi_1 _0988_ (.A1(net228),
    .A2(_0383_),
    .Y(_0088_),
    .B1(_0385_));
 sg13g2_nand3_1 _0989_ (.B(_0161_),
    .C(_0381_),
    .A(net228),
    .Y(_0386_));
 sg13g2_o21ai_1 _0990_ (.B1(_0386_),
    .Y(_0089_),
    .A1(_0140_),
    .A2(_0363_));
 sg13g2_mux2_1 _0991_ (.A0(net5),
    .A1(net255),
    .S(net100),
    .X(_0090_));
 sg13g2_mux2_1 _0992_ (.A0(net6),
    .A1(net277),
    .S(net100),
    .X(_0091_));
 sg13g2_mux2_1 _0993_ (.A0(net7),
    .A1(net278),
    .S(net100),
    .X(_0092_));
 sg13g2_xnor2_1 _0994_ (.Y(_0387_),
    .A(net109),
    .B(\ctr1.led_mask_i[0] ));
 sg13g2_nand2_1 _0995_ (.Y(_0388_),
    .A(net197),
    .B(net95));
 sg13g2_o21ai_1 _0996_ (.B1(_0388_),
    .Y(_0093_),
    .A1(net95),
    .A2(_0387_));
 sg13g2_xnor2_1 _0997_ (.Y(_0389_),
    .A(net109),
    .B(\ctr1.led_mask_i[1] ));
 sg13g2_nand2_1 _0998_ (.Y(_0390_),
    .A(net182),
    .B(net95));
 sg13g2_o21ai_1 _0999_ (.B1(_0390_),
    .Y(_0094_),
    .A1(net95),
    .A2(_0389_));
 sg13g2_xnor2_1 _1000_ (.Y(_0391_),
    .A(net109),
    .B(\ctr1.led_mask_i[2] ));
 sg13g2_nand2_1 _1001_ (.Y(_0392_),
    .A(net188),
    .B(net97));
 sg13g2_o21ai_1 _1002_ (.B1(_0392_),
    .Y(_0095_),
    .A1(net97),
    .A2(_0391_));
 sg13g2_xnor2_1 _1003_ (.Y(_0393_),
    .A(net109),
    .B(\ctr1.led_mask_i[3] ));
 sg13g2_nand2_1 _1004_ (.Y(_0394_),
    .A(net206),
    .B(net97));
 sg13g2_o21ai_1 _1005_ (.B1(_0394_),
    .Y(_0096_),
    .A1(net97),
    .A2(_0393_));
 sg13g2_xor2_1 _1006_ (.B(\ctr1.led_mask_i[4] ),
    .A(net110),
    .X(_0395_));
 sg13g2_nor2_1 _1007_ (.A(net98),
    .B(_0395_),
    .Y(_0396_));
 sg13g2_a21oi_1 _1008_ (.A1(_0123_),
    .A2(net97),
    .Y(_0097_),
    .B1(_0396_));
 sg13g2_xnor2_1 _1009_ (.Y(_0397_),
    .A(net110),
    .B(\ctr1.led_mask_i[5] ));
 sg13g2_nand2_1 _1010_ (.Y(_0398_),
    .A(net184),
    .B(net97));
 sg13g2_o21ai_1 _1011_ (.B1(_0398_),
    .Y(_0098_),
    .A1(net97),
    .A2(_0397_));
 sg13g2_xor2_1 _1012_ (.B(net344),
    .A(net110),
    .X(_0399_));
 sg13g2_nor2_1 _1013_ (.A(net98),
    .B(_0399_),
    .Y(_0400_));
 sg13g2_a21oi_1 _1014_ (.A1(_0124_),
    .A2(net98),
    .Y(_0099_),
    .B1(_0400_));
 sg13g2_xor2_1 _1015_ (.B(net345),
    .A(net110),
    .X(_0401_));
 sg13g2_nor2_1 _1016_ (.A(net97),
    .B(_0401_),
    .Y(_0402_));
 sg13g2_a21oi_1 _1017_ (.A1(_0125_),
    .A2(net98),
    .Y(_0100_),
    .B1(_0402_));
 sg13g2_xnor2_1 _1018_ (.Y(_0403_),
    .A(net109),
    .B(\ctr1.led_mask_i[8] ));
 sg13g2_nand2_1 _1019_ (.Y(_0404_),
    .A(net224),
    .B(net95));
 sg13g2_o21ai_1 _1020_ (.B1(_0404_),
    .Y(_0101_),
    .A1(net95),
    .A2(_0403_));
 sg13g2_xnor2_1 _1021_ (.Y(_0405_),
    .A(net109),
    .B(\ctr1.led_mask_i[9] ));
 sg13g2_nand2_1 _1022_ (.Y(_0406_),
    .A(net194),
    .B(net95));
 sg13g2_o21ai_1 _1023_ (.B1(_0406_),
    .Y(_0102_),
    .A1(net95),
    .A2(_0405_));
 sg13g2_xnor2_1 _1024_ (.Y(_0407_),
    .A(net109),
    .B(\ctr1.led_mask_i[10] ));
 sg13g2_nand2_1 _1025_ (.Y(_0408_),
    .A(net212),
    .B(net96));
 sg13g2_o21ai_1 _1026_ (.B1(_0408_),
    .Y(_0103_),
    .A1(net96),
    .A2(_0407_));
 sg13g2_xnor2_1 _1027_ (.Y(_0409_),
    .A(net109),
    .B(\ctr1.led_mask_i[11] ));
 sg13g2_nand2_1 _1028_ (.Y(_0410_),
    .A(net199),
    .B(net96));
 sg13g2_o21ai_1 _1029_ (.B1(_0410_),
    .Y(_0104_),
    .A1(net96),
    .A2(_0409_));
 sg13g2_a22oi_1 _1030_ (.Y(_0411_),
    .B1(_0328_),
    .B2(_0333_),
    .A2(_0327_),
    .A1(_0326_));
 sg13g2_mux2_1 _1031_ (.A0(net262),
    .A1(net106),
    .S(_0411_),
    .X(_0105_));
 sg13g2_nand2b_1 _1032_ (.Y(_0412_),
    .B(\leddriv1.byte_pos[0] ),
    .A_N(\leddriv1.reg_intensity[1] ));
 sg13g2_o21ai_1 _1033_ (.B1(_0412_),
    .Y(_0413_),
    .A1(\leddriv1.byte_pos[0] ),
    .A2(\leddriv1.reg_intensity[0] ));
 sg13g2_nand3_1 _1034_ (.B(\leddriv1.byte_pos[1] ),
    .C(\leddriv1.reg_intensity[3] ),
    .A(\leddriv1.byte_pos[0] ),
    .Y(_0414_));
 sg13g2_o21ai_1 _1035_ (.B1(_0414_),
    .Y(_0415_),
    .A1(\leddriv1.byte_pos[1] ),
    .A2(_0413_));
 sg13g2_nand3_1 _1036_ (.B(\leddriv1.reg_intensity[5] ),
    .C(_0011_),
    .A(\leddriv1.byte_pos[0] ),
    .Y(_0416_));
 sg13g2_mux2_1 _1037_ (.A0(\leddriv1.reg_colour[0] ),
    .A1(\leddriv1.reg_colour[1] ),
    .S(\leddriv1.grb_pos[0] ),
    .X(_0417_));
 sg13g2_nand2b_1 _1038_ (.Y(_0418_),
    .B(_0417_),
    .A_N(\leddriv1.grb_pos[1] ));
 sg13g2_nand3b_1 _1039_ (.B(\leddriv1.reg_colour[2] ),
    .C(\leddriv1.grb_pos[1] ),
    .Y(_0419_),
    .A_N(\leddriv1.grb_pos[0] ));
 sg13g2_a22oi_1 _1040_ (.Y(_0420_),
    .B1(_0418_),
    .B2(_0419_),
    .A2(_0416_),
    .A1(net275));
 sg13g2_o21ai_1 _1041_ (.B1(_0420_),
    .Y(_0421_),
    .A1(net275),
    .A2(_0415_));
 sg13g2_mux2_1 _1042_ (.A0(_0421_),
    .A1(net300),
    .S(_0326_),
    .X(_0106_));
 sg13g2_nand2b_1 _1043_ (.Y(_0422_),
    .B(net116),
    .A_N(_0179_));
 sg13g2_a221oi_1 _1044_ (.B2(_0119_),
    .C1(_0422_),
    .B1(_0182_),
    .A1(net105),
    .Y(_0107_),
    .A2(_0154_));
 sg13g2_nor2_1 _1045_ (.A(net296),
    .B(net99),
    .Y(_0423_));
 sg13g2_or2_2 _1046_ (.X(_0424_),
    .B(_0423_),
    .A(_0180_));
 sg13g2_nand2_1 _1047_ (.Y(_0425_),
    .A(net163),
    .B(_0180_));
 sg13g2_o21ai_1 _1048_ (.B1(_0425_),
    .Y(_0108_),
    .A1(_0130_),
    .A2(_0424_));
 sg13g2_a21oi_1 _1049_ (.A1(\leddriv1.tl_counter[0] ),
    .A2(_0424_),
    .Y(_0426_),
    .B1(net302));
 sg13g2_and3_1 _1050_ (.X(_0427_),
    .A(\leddriv1.tl_counter[0] ),
    .B(net302),
    .C(_0424_));
 sg13g2_nand3_1 _1051_ (.B(net302),
    .C(_0424_),
    .A(\leddriv1.tl_counter[0] ),
    .Y(_0428_));
 sg13g2_nor3_1 _1052_ (.A(_0423_),
    .B(net303),
    .C(_0427_),
    .Y(_0109_));
 sg13g2_and3_1 _1053_ (.X(_0429_),
    .A(\leddriv1.tl_counter[0] ),
    .B(\leddriv1.tl_counter[2] ),
    .C(\leddriv1.tl_counter[1] ));
 sg13g2_nand3_1 _1054_ (.B(net309),
    .C(net302),
    .A(\leddriv1.tl_counter[0] ),
    .Y(_0430_));
 sg13g2_nand2_1 _1055_ (.Y(_0431_),
    .A(net296),
    .B(_0430_));
 sg13g2_a22oi_1 _1056_ (.Y(_0110_),
    .B1(_0431_),
    .B2(_0424_),
    .A2(_0428_),
    .A1(_0132_));
 sg13g2_nor3_1 _1057_ (.A(net330),
    .B(_0181_),
    .C(_0430_),
    .Y(_0432_));
 sg13g2_a21oi_1 _1058_ (.A1(_0424_),
    .A2(_0431_),
    .Y(_0433_),
    .B1(_0133_));
 sg13g2_or2_1 _1059_ (.X(_0111_),
    .B(_0433_),
    .A(net331));
 sg13g2_nand3_1 _1060_ (.B(\leddriv1.tl_counter[3] ),
    .C(_0429_),
    .A(net266),
    .Y(_0434_));
 sg13g2_nand2_1 _1061_ (.Y(_0435_),
    .A(\leddriv1.state[1] ),
    .B(_0434_));
 sg13g2_o21ai_1 _1062_ (.B1(_0435_),
    .Y(_0436_),
    .A1(_0180_),
    .A2(_0423_));
 sg13g2_nand3_1 _1063_ (.B(_0424_),
    .C(_0429_),
    .A(\leddriv1.tl_counter[3] ),
    .Y(_0437_));
 sg13g2_a22oi_1 _1064_ (.Y(_0112_),
    .B1(_0437_),
    .B2(_0131_),
    .A2(_0435_),
    .A1(_0424_));
 sg13g2_nand2_1 _1065_ (.Y(_0438_),
    .A(net233),
    .B(_0436_));
 sg13g2_o21ai_1 _1066_ (.B1(net234),
    .Y(_0113_),
    .A1(_0181_),
    .A2(_0434_));
 sg13g2_nand2_1 _1067_ (.Y(_0439_),
    .A(net117),
    .B(net9));
 sg13g2_nand2_1 _1068_ (.Y(_0440_),
    .A(net117),
    .B(net8));
 sg13g2_and3_1 _1069_ (.X(_0114_),
    .A(net117),
    .B(net9),
    .C(net8));
 sg13g2_nor2_1 _1070_ (.A(net8),
    .B(_0439_),
    .Y(_0115_));
 sg13g2_nor2_1 _1071_ (.A(net9),
    .B(_0440_),
    .Y(_0116_));
 sg13g2_o21ai_1 _1072_ (.B1(net117),
    .Y(_0117_),
    .A1(net9),
    .A2(net8));
 sg13g2_buf_1 _1073_ (.A(net176),
    .X(_0078_));
 sg13g2_dfrbp_1 _1074_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net73),
    .D(_0019_),
    .Q_N(_0529_),
    .Q(\ctr1.led_binary[0] ));
 sg13g2_dfrbp_1 _1075_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net43),
    .D(_0020_),
    .Q_N(_0528_),
    .Q(\ctr1.led_binary[1] ));
 sg13g2_dfrbp_1 _1076_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net41),
    .D(_0021_),
    .Q_N(_0527_),
    .Q(\ctr1.led_binary[2] ));
 sg13g2_dfrbp_1 _1077_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net39),
    .D(_0022_),
    .Q_N(_0526_),
    .Q(\ctr1.led_binary[3] ));
 sg13g2_dfrbp_1 _1078_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net37),
    .D(_0023_),
    .Q_N(_0525_),
    .Q(\ctr1.led_mask_i[0] ));
 sg13g2_dfrbp_1 _1079_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net35),
    .D(net334),
    .Q_N(_0524_),
    .Q(\ctr1.led_mask_i[1] ));
 sg13g2_dfrbp_1 _1080_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net33),
    .D(net337),
    .Q_N(_0523_),
    .Q(\ctr1.led_mask_i[2] ));
 sg13g2_dfrbp_1 _1081_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net31),
    .D(_0026_),
    .Q_N(_0522_),
    .Q(\ctr1.led_mask_i[3] ));
 sg13g2_dfrbp_1 _1082_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net29),
    .D(_0027_),
    .Q_N(_0521_),
    .Q(\ctr1.led_mask_i[4] ));
 sg13g2_dfrbp_1 _1083_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net162),
    .D(_0028_),
    .Q_N(_0520_),
    .Q(\ctr1.led_mask_i[5] ));
 sg13g2_dfrbp_1 _1084_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net160),
    .D(_0029_),
    .Q_N(_0519_),
    .Q(\ctr1.led_mask_i[6] ));
 sg13g2_dfrbp_1 _1085_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net158),
    .D(net326),
    .Q_N(_0518_),
    .Q(\ctr1.led_mask_i[7] ));
 sg13g2_dfrbp_1 _1086_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net156),
    .D(net324),
    .Q_N(_0517_),
    .Q(\ctr1.led_mask_i[8] ));
 sg13g2_dfrbp_1 _1087_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net154),
    .D(_0032_),
    .Q_N(_0516_),
    .Q(\ctr1.led_mask_i[9] ));
 sg13g2_dfrbp_1 _1088_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net152),
    .D(_0033_),
    .Q_N(_0515_),
    .Q(\ctr1.led_mask_i[10] ));
 sg13g2_dfrbp_1 _1089_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net150),
    .D(_0034_),
    .Q_N(_0514_),
    .Q(\ctr1.led_mask_i[11] ));
 sg13g2_dfrbp_1 _1090_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net148),
    .D(_0035_),
    .Q_N(_0513_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1091_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net147),
    .D(_0036_),
    .Q_N(_0512_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1092_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net146),
    .D(_0037_),
    .Q_N(_0511_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _1093_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net145),
    .D(_0038_),
    .Q_N(_0510_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _1094_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net144),
    .D(_0039_),
    .Q_N(_0509_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1095_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net143),
    .D(net173),
    .Q_N(_0008_),
    .Q(\ctr1.inverted ));
 sg13g2_dfrbp_1 _1096_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net141),
    .D(_0041_),
    .Q_N(_0508_),
    .Q(\rdec1.dn_detected ));
 sg13g2_dfrbp_1 _1097_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net140),
    .D(net203),
    .Q_N(_0507_),
    .Q(\rdec1.up_detected ));
 sg13g2_dfrbp_1 _1098_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net139),
    .D(_0043_),
    .Q_N(_0018_),
    .Q(\rdec1.pause_counter[0] ));
 sg13g2_dfrbp_1 _1099_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net137),
    .D(net240),
    .Q_N(_0506_),
    .Q(\rdec1.pause_counter[1] ));
 sg13g2_dfrbp_1 _1100_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net135),
    .D(_0045_),
    .Q_N(_0505_),
    .Q(\rdec1.pause_counter[2] ));
 sg13g2_dfrbp_1 _1101_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net133),
    .D(net193),
    .Q_N(_0504_),
    .Q(\rdec1.pause_counter[3] ));
 sg13g2_dfrbp_1 _1102_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net131),
    .D(net270),
    .Q_N(_0503_),
    .Q(\rdec1.pause_counter[4] ));
 sg13g2_dfrbp_1 _1103_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net129),
    .D(net247),
    .Q_N(_0502_),
    .Q(\rdec1.pause_counter[5] ));
 sg13g2_dfrbp_1 _1104_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net127),
    .D(_0049_),
    .Q_N(_0501_),
    .Q(\rdec1.pause_counter[6] ));
 sg13g2_dfrbp_1 _1105_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net125),
    .D(net211),
    .Q_N(_0500_),
    .Q(\rdec1.pause_counter[7] ));
 sg13g2_dfrbp_1 _1106_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net123),
    .D(_0051_),
    .Q_N(_0499_),
    .Q(\rdec1.pause_counter[8] ));
 sg13g2_dfrbp_1 _1107_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net121),
    .D(_0052_),
    .Q_N(_0498_),
    .Q(\rdec1.pause_counter[9] ));
 sg13g2_dfrbp_1 _1108_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net119),
    .D(net295),
    .Q_N(_0497_),
    .Q(\rdec1.pause_counter[10] ));
 sg13g2_dfrbp_1 _1109_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net89),
    .D(net292),
    .Q_N(_0496_),
    .Q(\rdec1.pause_counter[11] ));
 sg13g2_dfrbp_1 _1110_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net87),
    .D(net273),
    .Q_N(_0495_),
    .Q(\rdec1.pause_counter[12] ));
 sg13g2_dfrbp_1 _1111_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net85),
    .D(net287),
    .Q_N(_0494_),
    .Q(\rdec1.pause_counter[13] ));
 sg13g2_dfrbp_1 _1112_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net83),
    .D(net290),
    .Q_N(_0493_),
    .Q(\rdec1.pause_counter[14] ));
 sg13g2_dfrbp_1 _1113_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net81),
    .D(_0058_),
    .Q_N(_0492_),
    .Q(\ctr1.rot_dn ));
 sg13g2_dfrbp_1 _1114_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net71),
    .D(_0059_),
    .Q_N(_0491_),
    .Q(\ctr1.rot_up ));
 sg13g2_dfrbp_1 _1115_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net69),
    .D(net181),
    .Q_N(_0490_),
    .Q(\leddriv1.reg_intensity[0] ));
 sg13g2_dfrbp_1 _1116_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net68),
    .D(net191),
    .Q_N(_0489_),
    .Q(\leddriv1.reg_intensity[1] ));
 sg13g2_dfrbp_1 _1117_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net67),
    .D(net217),
    .Q_N(_0488_),
    .Q(\leddriv1.reg_intensity[3] ));
 sg13g2_dfrbp_1 _1118_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net74),
    .D(net187),
    .Q_N(_0530_),
    .Q(\leddriv1.reg_intensity[5] ));
 sg13g2_dfrbp_1 _1119_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net75),
    .D(_0005_),
    .Q_N(_0531_),
    .Q(\rdec1.state[0] ));
 sg13g2_dfrbp_1 _1120_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net76),
    .D(_0006_),
    .Q_N(_0532_),
    .Q(\rdec1.state[1] ));
 sg13g2_dfrbp_1 _1121_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net77),
    .D(_0000_),
    .Q_N(_0533_),
    .Q(\rdec1.state[2] ));
 sg13g2_dfrbp_1 _1122_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net78),
    .D(net261),
    .Q_N(_0534_),
    .Q(\rdec1.state[3] ));
 sg13g2_dfrbp_1 _1123_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net79),
    .D(_0001_),
    .Q_N(_0535_),
    .Q(\leddriv1.state[0] ));
 sg13g2_dfrbp_1 _1124_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net80),
    .D(_0002_),
    .Q_N(_0536_),
    .Q(\leddriv1.state[1] ));
 sg13g2_dfrbp_1 _1125_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net28),
    .D(_0003_),
    .Q_N(_0009_),
    .Q(\leddriv1.state[2] ));
 sg13g2_dfrbp_1 _1126_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net66),
    .D(net263),
    .Q_N(_0487_),
    .Q(\leddriv1.state[3] ));
 sg13g2_dfrbp_1 _1127_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net65),
    .D(net167),
    .Q_N(_0017_),
    .Q(\leddriv1.byte_pos[0] ));
 sg13g2_dfrbp_1 _1128_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net63),
    .D(net243),
    .Q_N(_0011_),
    .Q(\leddriv1.byte_pos[1] ));
 sg13g2_dfrbp_1 _1129_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net61),
    .D(net276),
    .Q_N(_0010_),
    .Q(\leddriv1.byte_pos[2] ));
 sg13g2_dfrbp_1 _1130_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net59),
    .D(net285),
    .Q_N(_0016_),
    .Q(\leddriv1.grb_pos[0] ));
 sg13g2_dfrbp_1 _1131_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net57),
    .D(net322),
    .Q_N(_0486_),
    .Q(\leddriv1.grb_pos[1] ));
 sg13g2_dfrbp_1 _1132_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net55),
    .D(net314),
    .Q_N(_0015_),
    .Q(\leddriv1.led_pos[0] ));
 sg13g2_dfrbp_1 _1133_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net53),
    .D(_0070_),
    .Q_N(_0485_),
    .Q(\leddriv1.led_pos[1] ));
 sg13g2_dfrbp_1 _1134_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net51),
    .D(_0071_),
    .Q_N(_0484_),
    .Q(\leddriv1.led_pos[2] ));
 sg13g2_dfrbp_1 _1135_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net49),
    .D(net308),
    .Q_N(_0483_),
    .Q(\leddriv1.led_pos[3] ));
 sg13g2_dfrbp_1 _1136_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net47),
    .D(net175),
    .Q_N(_0014_),
    .Q(\leddriv1.th_counter[0] ));
 sg13g2_dfrbp_1 _1137_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net46),
    .D(net329),
    .Q_N(_0482_),
    .Q(\leddriv1.th_counter[1] ));
 sg13g2_dfrbp_1 _1138_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net45),
    .D(net237),
    .Q_N(_0481_),
    .Q(\leddriv1.th_counter[2] ));
 sg13g2_dfrbp_1 _1139_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net44),
    .D(net245),
    .Q_N(_0480_),
    .Q(\leddriv1.th_counter[3] ));
 sg13g2_dfrbp_1 _1140_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net42),
    .D(net178),
    .Q_N(_0479_),
    .Q(\leddriv1.th_counter[4] ));
 sg13g2_dfrbp_1 _1141_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net40),
    .D(_0078_),
    .Q_N(_0478_),
    .Q(\leddriv1.th_counter[5] ));
 sg13g2_dfrbp_1 _1142_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net38),
    .D(_0079_),
    .Q_N(_0013_),
    .Q(\leddriv1.rs_counter[0] ));
 sg13g2_dfrbp_1 _1143_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net34),
    .D(net318),
    .Q_N(_0477_),
    .Q(\leddriv1.rs_counter[1] ));
 sg13g2_dfrbp_1 _1144_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net30),
    .D(net205),
    .Q_N(_0476_),
    .Q(\leddriv1.rs_counter[2] ));
 sg13g2_dfrbp_1 _1145_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net161),
    .D(net254),
    .Q_N(_0475_),
    .Q(\leddriv1.rs_counter[3] ));
 sg13g2_dfrbp_1 _1146_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net157),
    .D(net250),
    .Q_N(_0474_),
    .Q(\leddriv1.rs_counter[4] ));
 sg13g2_dfrbp_1 _1147_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net153),
    .D(net265),
    .Q_N(_0473_),
    .Q(\leddriv1.rs_counter[5] ));
 sg13g2_dfrbp_1 _1148_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net149),
    .D(net252),
    .Q_N(_0472_),
    .Q(\leddriv1.rs_counter[6] ));
 sg13g2_dfrbp_1 _1149_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net138),
    .D(_0086_),
    .Q_N(_0471_),
    .Q(\leddriv1.rs_counter[7] ));
 sg13g2_dfrbp_1 _1150_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net134),
    .D(_0087_),
    .Q_N(_0470_),
    .Q(\leddriv1.rs_counter[8] ));
 sg13g2_dfrbp_1 _1151_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net130),
    .D(net229),
    .Q_N(_0469_),
    .Q(\leddriv1.rs_counter[9] ));
 sg13g2_dfrbp_1 _1152_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net126),
    .D(net257),
    .Q_N(_0468_),
    .Q(\leddriv1.rs_counter[10] ));
 sg13g2_dfrbp_1 _1153_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net122),
    .D(_0090_),
    .Q_N(_0467_),
    .Q(\leddriv1.reg_colour[0] ));
 sg13g2_dfrbp_1 _1154_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net120),
    .D(_0091_),
    .Q_N(_0466_),
    .Q(\leddriv1.reg_colour[1] ));
 sg13g2_dfrbp_1 _1155_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net118),
    .D(_0092_),
    .Q_N(_0465_),
    .Q(\leddriv1.reg_colour[2] ));
 sg13g2_dfrbp_1 _1156_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net88),
    .D(net198),
    .Q_N(_0464_),
    .Q(\leddriv1.reg_led_mask[0] ));
 sg13g2_dfrbp_1 _1157_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net86),
    .D(net183),
    .Q_N(_0463_),
    .Q(\leddriv1.reg_led_mask[1] ));
 sg13g2_dfrbp_1 _1158_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net84),
    .D(net189),
    .Q_N(_0462_),
    .Q(\leddriv1.reg_led_mask[2] ));
 sg13g2_dfrbp_1 _1159_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net82),
    .D(net207),
    .Q_N(_0461_),
    .Q(\leddriv1.reg_led_mask[3] ));
 sg13g2_dfrbp_1 _1160_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net72),
    .D(net223),
    .Q_N(_0460_),
    .Q(\leddriv1.reg_led_mask[4] ));
 sg13g2_dfrbp_1 _1161_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net70),
    .D(net185),
    .Q_N(_0459_),
    .Q(\leddriv1.reg_led_mask[5] ));
 sg13g2_dfrbp_1 _1162_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net64),
    .D(_0099_),
    .Q_N(_0458_),
    .Q(\leddriv1.reg_led_mask[6] ));
 sg13g2_dfrbp_1 _1163_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net62),
    .D(_0100_),
    .Q_N(_0457_),
    .Q(\leddriv1.reg_led_mask[7] ));
 sg13g2_dfrbp_1 _1164_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net60),
    .D(net225),
    .Q_N(_0456_),
    .Q(\leddriv1.reg_led_mask[8] ));
 sg13g2_dfrbp_1 _1165_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net58),
    .D(net195),
    .Q_N(_0455_),
    .Q(\leddriv1.reg_led_mask[9] ));
 sg13g2_dfrbp_1 _1166_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net56),
    .D(net213),
    .Q_N(_0454_),
    .Q(\leddriv1.reg_led_mask[10] ));
 sg13g2_dfrbp_1 _1167_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net54),
    .D(net200),
    .Q_N(_0453_),
    .Q(\leddriv1.reg_led_mask[11] ));
 sg13g2_dfrbp_1 _1168_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net52),
    .D(net280),
    .Q_N(_0452_),
    .Q(\leddriv1.skip_calc ));
 sg13g2_dfrbp_1 _1169_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net50),
    .D(_0106_),
    .Q_N(_0451_),
    .Q(\leddriv1.tl_max[1] ));
 sg13g2_dfrbp_1 _1170_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net48),
    .D(net231),
    .Q_N(_0450_),
    .Q(\leddriv1.led_dout ));
 sg13g2_dfrbp_1 _1171_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net32),
    .D(net164),
    .Q_N(_0012_),
    .Q(\leddriv1.tl_counter[0] ));
 sg13g2_dfrbp_1 _1172_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net159),
    .D(net304),
    .Q_N(_0449_),
    .Q(\leddriv1.tl_counter[1] ));
 sg13g2_dfrbp_1 _1173_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net151),
    .D(net310),
    .Q_N(_0448_),
    .Q(\leddriv1.tl_counter[2] ));
 sg13g2_dfrbp_1 _1174_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net136),
    .D(_0111_),
    .Q_N(_0447_),
    .Q(\leddriv1.tl_counter[3] ));
 sg13g2_dfrbp_1 _1175_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net128),
    .D(net267),
    .Q_N(_0446_),
    .Q(\leddriv1.tl_counter[4] ));
 sg13g2_dfrbp_1 _1176_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net36),
    .D(net235),
    .Q_N(_0445_),
    .Q(\leddriv1.tl_counter[5] ));
 sg13g2_dfrbp_1 _1177_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net155),
    .D(_0114_),
    .Q_N(_0444_),
    .Q(\ctr1.intensity_out[5] ));
 sg13g2_dfrbp_1 _1178_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net142),
    .D(_0115_),
    .Q_N(_0443_),
    .Q(\ctr1.intensity_out[3] ));
 sg13g2_dfrbp_1 _1179_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net132),
    .D(_0116_),
    .Q_N(_0442_),
    .Q(\ctr1.intensity_out[1] ));
 sg13g2_dfrbp_1 _1180_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net124),
    .D(_0117_),
    .Q_N(_0441_),
    .Q(\ctr1.intensity_out[0] ));
 sg13g2_tiehi _1082__29 (.L_HI(net29));
 sg13g2_tiehi _1144__30 (.L_HI(net30));
 sg13g2_tiehi _1081__31 (.L_HI(net31));
 sg13g2_tiehi _1171__32 (.L_HI(net32));
 sg13g2_tiehi _1080__33 (.L_HI(net33));
 sg13g2_tiehi _1143__34 (.L_HI(net34));
 sg13g2_tiehi _1079__35 (.L_HI(net35));
 sg13g2_tiehi _1176__36 (.L_HI(net36));
 sg13g2_tiehi _1078__37 (.L_HI(net37));
 sg13g2_tiehi _1142__38 (.L_HI(net38));
 sg13g2_tiehi _1077__39 (.L_HI(net39));
 sg13g2_tiehi _1141__40 (.L_HI(net40));
 sg13g2_tiehi _1076__41 (.L_HI(net41));
 sg13g2_tiehi _1140__42 (.L_HI(net42));
 sg13g2_tiehi _1075__43 (.L_HI(net43));
 sg13g2_tiehi _1139__44 (.L_HI(net44));
 sg13g2_tiehi _1138__45 (.L_HI(net45));
 sg13g2_tiehi _1137__46 (.L_HI(net46));
 sg13g2_tiehi _1136__47 (.L_HI(net47));
 sg13g2_tiehi _1170__48 (.L_HI(net48));
 sg13g2_tiehi _1135__49 (.L_HI(net49));
 sg13g2_tiehi _1169__50 (.L_HI(net50));
 sg13g2_tiehi _1134__51 (.L_HI(net51));
 sg13g2_tiehi _1168__52 (.L_HI(net52));
 sg13g2_tiehi _1133__53 (.L_HI(net53));
 sg13g2_tiehi _1167__54 (.L_HI(net54));
 sg13g2_tiehi _1132__55 (.L_HI(net55));
 sg13g2_tiehi _1166__56 (.L_HI(net56));
 sg13g2_tiehi _1131__57 (.L_HI(net57));
 sg13g2_tiehi _1165__58 (.L_HI(net58));
 sg13g2_tiehi _1130__59 (.L_HI(net59));
 sg13g2_tiehi _1164__60 (.L_HI(net60));
 sg13g2_tiehi _1129__61 (.L_HI(net61));
 sg13g2_tiehi _1163__62 (.L_HI(net62));
 sg13g2_tiehi _1128__63 (.L_HI(net63));
 sg13g2_tiehi _1162__64 (.L_HI(net64));
 sg13g2_tiehi _1127__65 (.L_HI(net65));
 sg13g2_tiehi _1126__66 (.L_HI(net66));
 sg13g2_tiehi _1117__67 (.L_HI(net67));
 sg13g2_tiehi _1116__68 (.L_HI(net68));
 sg13g2_tiehi _1115__69 (.L_HI(net69));
 sg13g2_tiehi _1161__70 (.L_HI(net70));
 sg13g2_tiehi _1114__71 (.L_HI(net71));
 sg13g2_tiehi _1160__72 (.L_HI(net72));
 sg13g2_tiehi _1074__73 (.L_HI(net73));
 sg13g2_tiehi _1118__74 (.L_HI(net74));
 sg13g2_tiehi _1119__75 (.L_HI(net75));
 sg13g2_tiehi _1120__76 (.L_HI(net76));
 sg13g2_tiehi _1121__77 (.L_HI(net77));
 sg13g2_tiehi _1122__78 (.L_HI(net78));
 sg13g2_tiehi _1123__79 (.L_HI(net79));
 sg13g2_tiehi _1124__80 (.L_HI(net80));
 sg13g2_tiehi _1113__81 (.L_HI(net81));
 sg13g2_tiehi _1159__82 (.L_HI(net82));
 sg13g2_tiehi _1112__83 (.L_HI(net83));
 sg13g2_tiehi _1158__84 (.L_HI(net84));
 sg13g2_tiehi _1111__85 (.L_HI(net85));
 sg13g2_tiehi _1157__86 (.L_HI(net86));
 sg13g2_tiehi _1110__87 (.L_HI(net87));
 sg13g2_tiehi _1156__88 (.L_HI(net88));
 sg13g2_tiehi _1109__89 (.L_HI(net89));
 sg13g2_tiehi _1155__90 (.L_HI(net118));
 sg13g2_tiehi _1108__91 (.L_HI(net119));
 sg13g2_tiehi _1154__92 (.L_HI(net120));
 sg13g2_tiehi _1107__93 (.L_HI(net121));
 sg13g2_tiehi _1153__94 (.L_HI(net122));
 sg13g2_tiehi _1106__95 (.L_HI(net123));
 sg13g2_tiehi _1180__96 (.L_HI(net124));
 sg13g2_tiehi _1105__97 (.L_HI(net125));
 sg13g2_tiehi _1152__98 (.L_HI(net126));
 sg13g2_tiehi _1104__99 (.L_HI(net127));
 sg13g2_tiehi _1175__100 (.L_HI(net128));
 sg13g2_tiehi _1103__101 (.L_HI(net129));
 sg13g2_tiehi _1151__102 (.L_HI(net130));
 sg13g2_tiehi _1102__103 (.L_HI(net131));
 sg13g2_tiehi _1179__104 (.L_HI(net132));
 sg13g2_tiehi _1101__105 (.L_HI(net133));
 sg13g2_tiehi _1150__106 (.L_HI(net134));
 sg13g2_tiehi _1100__107 (.L_HI(net135));
 sg13g2_tiehi _1174__108 (.L_HI(net136));
 sg13g2_tiehi _1099__109 (.L_HI(net137));
 sg13g2_tiehi _1149__110 (.L_HI(net138));
 sg13g2_tiehi _1098__111 (.L_HI(net139));
 sg13g2_tiehi _1097__112 (.L_HI(net140));
 sg13g2_tiehi _1096__113 (.L_HI(net141));
 sg13g2_tiehi _1178__114 (.L_HI(net142));
 sg13g2_tiehi _1095__115 (.L_HI(net143));
 sg13g2_tiehi _1094__116 (.L_HI(net144));
 sg13g2_tiehi _1093__117 (.L_HI(net145));
 sg13g2_tiehi _1092__118 (.L_HI(net146));
 sg13g2_tiehi _1091__119 (.L_HI(net147));
 sg13g2_tiehi _1090__120 (.L_HI(net148));
 sg13g2_tiehi _1148__121 (.L_HI(net149));
 sg13g2_tiehi _1089__122 (.L_HI(net150));
 sg13g2_tiehi _1173__123 (.L_HI(net151));
 sg13g2_tiehi _1088__124 (.L_HI(net152));
 sg13g2_tiehi _1147__125 (.L_HI(net153));
 sg13g2_tiehi _1087__126 (.L_HI(net154));
 sg13g2_tiehi _1177__127 (.L_HI(net155));
 sg13g2_tiehi _1086__128 (.L_HI(net156));
 sg13g2_tiehi _1146__129 (.L_HI(net157));
 sg13g2_tiehi _1085__130 (.L_HI(net158));
 sg13g2_tiehi _1172__131 (.L_HI(net159));
 sg13g2_tiehi _1084__132 (.L_HI(net160));
 sg13g2_tiehi _1145__133 (.L_HI(net161));
 sg13g2_tiehi _1083__134 (.L_HI(net162));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_11 (.L_LO(net11));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_12 (.L_LO(net12));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_13 (.L_LO(net13));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_14 (.L_LO(net14));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_15 (.L_LO(net15));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_16 (.L_LO(net16));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_17 (.L_LO(net17));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_18 (.L_LO(net18));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_19 (.L_LO(net19));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_20 (.L_LO(net20));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_21 (.L_LO(net21));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_22 (.L_LO(net22));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_23 (.L_LO(net23));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_24 (.L_LO(net24));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_25 (.L_LO(net25));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_26 (.L_LO(net26));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_27 (.L_LO(net27));
 sg13g2_tiehi _1125__28 (.L_HI(net28));
 sg13g2_buf_1 _1306_ (.A(\leddriv1.led_dout ),
    .X(uo_out[0]));
 sg13g2_buf_2 fanout90 (.A(_0273_),
    .X(net90));
 sg13g2_buf_1 fanout91 (.A(_0273_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0236_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_0232_),
    .X(net93));
 sg13g2_buf_1 fanout94 (.A(_0232_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(net99),
    .X(net95));
 sg13g2_buf_1 fanout96 (.A(net99),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(net98),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(net99),
    .X(net98));
 sg13g2_buf_1 fanout99 (.A(net101),
    .X(net99));
 sg13g2_buf_4 fanout100 (.X(net100),
    .A(net101));
 sg13g2_buf_2 fanout101 (.A(_0148_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_0120_),
    .X(net102));
 sg13g2_buf_1 fanout103 (.A(_0120_),
    .X(net103));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(\leddriv1.led_pos[0] ));
 sg13g2_buf_2 fanout105 (.A(net346),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(net279),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(\rdec1.state[1] ),
    .X(net107));
 sg13g2_buf_1 fanout108 (.A(\rdec1.state[1] ),
    .X(net108));
 sg13g2_buf_4 fanout109 (.X(net109),
    .A(\ctr1.inverted ));
 sg13g2_buf_2 fanout110 (.A(net343),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(net113),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(net113),
    .X(net112));
 sg13g2_buf_1 fanout113 (.A(net114),
    .X(net113));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(net1));
 sg13g2_buf_2 fanout115 (.A(net116),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(net117),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(net1),
    .X(net117));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_tielo tt_um_faramire_rotary_ring_wrapper_10 (.L_LO(net10));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0012_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0108_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0017_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0337_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0064_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0013_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0361_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0018_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0274_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0008_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0040_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0014_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0073_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold14 (.A(\leddriv1.th_counter[5] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold15 (.A(\leddriv1.th_counter[4] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0077_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold17 (.A(\ctr1.led_binary[3] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold18 (.A(\ctr1.intensity_out[0] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0060_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold20 (.A(\leddriv1.reg_led_mask[1] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0094_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold22 (.A(\leddriv1.reg_led_mask[5] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0098_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold24 (.A(\ctr1.intensity_out[5] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0063_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold26 (.A(\leddriv1.reg_led_mask[2] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0095_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold28 (.A(\ctr1.intensity_out[1] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0061_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold30 (.A(\rdec1.pause_counter[3] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0046_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold32 (.A(\leddriv1.reg_led_mask[9] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0102_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold34 (.A(\ctr1.led_binary[0] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold35 (.A(\leddriv1.reg_led_mask[0] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0093_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold37 (.A(\leddriv1.reg_led_mask[11] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0104_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold39 (.A(\rdec1.up_detected ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0270_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0042_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold42 (.A(\leddriv1.rs_counter[2] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0081_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold44 (.A(\leddriv1.reg_led_mask[3] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0096_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold46 (.A(\ctr1.rot_up ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0314_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold48 (.A(\rdec1.pause_counter[7] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0050_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold50 (.A(\leddriv1.reg_led_mask[10] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0103_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold52 (.A(\ctr1.led_binary[2] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold53 (.A(\leddriv1.reg_led_mask[7] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold54 (.A(\ctr1.intensity_out[3] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0062_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold56 (.A(\rdec1.pause_counter[8] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0296_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold58 (.A(\rdec1.dn_detected ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0313_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold60 (.A(\leddriv1.reg_led_mask[4] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0097_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold62 (.A(\leddriv1.reg_led_mask[8] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0101_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold64 (.A(\rdec1.pause_counter[6] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0290_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold66 (.A(\leddriv1.rs_counter[9] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0088_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold68 (.A(\leddriv1.led_dout ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0107_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold70 (.A(\leddriv1.reg_led_mask[6] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold71 (.A(\leddriv1.tl_counter[5] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0438_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0113_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold74 (.A(\leddriv1.th_counter[2] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0075_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold76 (.A(\rdec1.pause_counter[1] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0275_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0044_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold79 (.A(\leddriv1.byte_pos[1] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0338_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0065_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold82 (.A(\leddriv1.th_counter[3] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0076_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold84 (.A(\rdec1.pause_counter[5] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0048_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold86 (.A(\ctr1.led_binary[1] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold87 (.A(\leddriv1.rs_counter[4] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0083_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold89 (.A(\leddriv1.rs_counter[6] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0085_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold91 (.A(\leddriv1.rs_counter[3] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0082_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold93 (.A(\leddriv1.reg_colour[0] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold94 (.A(\leddriv1.rs_counter[10] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0089_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold96 (.A(\leddriv1.rs_counter[8] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0384_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold98 (.A(\rdec1.state[3] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0007_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold100 (.A(\leddriv1.skip_calc ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0004_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold102 (.A(\leddriv1.rs_counter[5] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0084_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold104 (.A(\leddriv1.tl_counter[4] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0112_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold106 (.A(\rdec1.pause_counter[4] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0283_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0047_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold109 (.A(\rdec1.pause_counter[12] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0307_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0055_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold112 (.A(\rdec1.state[0] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold113 (.A(\leddriv1.byte_pos[2] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0066_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold115 (.A(\leddriv1.reg_colour[1] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold116 (.A(\leddriv1.reg_colour[2] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold117 (.A(\leddriv1.state[2] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0105_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold119 (.A(\leddriv1.state[3] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0162_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0016_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0345_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0067_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold124 (.A(\rdec1.pause_counter[13] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0056_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold126 (.A(\rdec1.pause_counter[14] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0312_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0057_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold129 (.A(\rdec1.pause_counter[11] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0054_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold131 (.A(\rdec1.pause_counter[10] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0302_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0053_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold134 (.A(\leddriv1.state[1] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0154_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold136 (.A(\ctr1.led_mask_i[6] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold137 (.A(\ctr1.led_mask_i[8] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold138 (.A(\leddriv1.tl_max[1] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold139 (.A(\rdec1.state[2] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold140 (.A(\leddriv1.tl_counter[1] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0426_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0109_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold143 (.A(\ctr1.led_mask_i[10] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold144 (.A(\leddriv1.rs_counter[7] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold145 (.A(\leddriv1.led_pos[2] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0072_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold147 (.A(\leddriv1.tl_counter[2] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0110_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold149 (.A(\leddriv1.led_pos[1] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0349_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0015_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0069_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold153 (.A(\rdec1.pause_counter[9] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold154 (.A(\leddriv1.rs_counter[1] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0364_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0080_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold157 (.A(\rdec1.pause_counter[2] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0281_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold159 (.A(\leddriv1.grb_pos[1] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0068_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold161 (.A(\ctr1.led_mask_i[9] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0031_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold163 (.A(\ctr1.led_mask_i[7] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0030_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold165 (.A(\leddriv1.th_counter[1] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0356_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0074_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold168 (.A(\leddriv1.tl_counter[3] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0432_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold170 (.A(\ctr1.led_mask_i[11] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold171 (.A(\ctr1.led_mask_i[2] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0024_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold173 (.A(\ctr1.led_mask_i[3] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0240_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0025_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold176 (.A(\ctr1.led_mask_i[4] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0243_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold178 (.A(\ctr1.led_mask_i[5] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold179 (.A(\ctr1.led_mask_i[0] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0235_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold181 (.A(\ctr1.inverted ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold182 (.A(\ctr1.led_mask_i[6] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold183 (.A(\ctr1.led_mask_i[7] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold184 (.A(\leddriv1.state[3] ),
    .X(net346));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_fill_2 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_278 ();
 sg13g2_decap_8 FILLER_13_285 ();
 sg13g2_decap_8 FILLER_13_292 ();
 sg13g2_decap_8 FILLER_13_299 ();
 sg13g2_decap_8 FILLER_13_306 ();
 sg13g2_decap_8 FILLER_13_313 ();
 sg13g2_decap_8 FILLER_13_320 ();
 sg13g2_decap_8 FILLER_13_327 ();
 sg13g2_decap_8 FILLER_13_334 ();
 sg13g2_decap_8 FILLER_13_341 ();
 sg13g2_decap_8 FILLER_13_348 ();
 sg13g2_decap_8 FILLER_13_355 ();
 sg13g2_decap_8 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_13_369 ();
 sg13g2_decap_8 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_fill_1 FILLER_14_231 ();
 sg13g2_fill_2 FILLER_14_245 ();
 sg13g2_decap_4 FILLER_14_260 ();
 sg13g2_fill_1 FILLER_14_273 ();
 sg13g2_fill_2 FILLER_14_288 ();
 sg13g2_decap_8 FILLER_14_304 ();
 sg13g2_decap_8 FILLER_14_311 ();
 sg13g2_decap_8 FILLER_14_318 ();
 sg13g2_decap_8 FILLER_14_325 ();
 sg13g2_decap_8 FILLER_14_332 ();
 sg13g2_decap_8 FILLER_14_339 ();
 sg13g2_fill_2 FILLER_14_346 ();
 sg13g2_fill_2 FILLER_14_356 ();
 sg13g2_fill_1 FILLER_14_363 ();
 sg13g2_fill_2 FILLER_14_381 ();
 sg13g2_fill_1 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_388 ();
 sg13g2_decap_8 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_fill_2 FILLER_15_217 ();
 sg13g2_fill_2 FILLER_15_223 ();
 sg13g2_fill_1 FILLER_15_225 ();
 sg13g2_decap_8 FILLER_15_312 ();
 sg13g2_decap_8 FILLER_15_319 ();
 sg13g2_decap_8 FILLER_15_326 ();
 sg13g2_decap_4 FILLER_15_333 ();
 sg13g2_fill_2 FILLER_15_337 ();
 sg13g2_fill_2 FILLER_15_365 ();
 sg13g2_fill_1 FILLER_15_367 ();
 sg13g2_fill_1 FILLER_15_382 ();
 sg13g2_fill_2 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_4 FILLER_16_203 ();
 sg13g2_fill_1 FILLER_16_207 ();
 sg13g2_fill_1 FILLER_16_273 ();
 sg13g2_fill_2 FILLER_16_283 ();
 sg13g2_fill_2 FILLER_16_294 ();
 sg13g2_fill_2 FILLER_16_343 ();
 sg13g2_fill_2 FILLER_16_359 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_4 FILLER_17_196 ();
 sg13g2_fill_2 FILLER_17_200 ();
 sg13g2_fill_1 FILLER_17_277 ();
 sg13g2_fill_2 FILLER_17_321 ();
 sg13g2_fill_1 FILLER_17_323 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_fill_2 FILLER_18_144 ();
 sg13g2_decap_8 FILLER_18_151 ();
 sg13g2_decap_8 FILLER_18_158 ();
 sg13g2_decap_8 FILLER_18_165 ();
 sg13g2_decap_8 FILLER_18_172 ();
 sg13g2_decap_8 FILLER_18_179 ();
 sg13g2_decap_8 FILLER_18_186 ();
 sg13g2_decap_8 FILLER_18_193 ();
 sg13g2_decap_8 FILLER_18_200 ();
 sg13g2_decap_4 FILLER_18_207 ();
 sg13g2_fill_2 FILLER_18_211 ();
 sg13g2_fill_2 FILLER_18_217 ();
 sg13g2_fill_2 FILLER_18_228 ();
 sg13g2_fill_1 FILLER_18_270 ();
 sg13g2_fill_1 FILLER_18_327 ();
 sg13g2_fill_1 FILLER_18_350 ();
 sg13g2_fill_2 FILLER_18_361 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_fill_2 FILLER_19_145 ();
 sg13g2_fill_1 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_157 ();
 sg13g2_fill_1 FILLER_19_164 ();
 sg13g2_fill_1 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_187 ();
 sg13g2_decap_8 FILLER_19_194 ();
 sg13g2_fill_2 FILLER_19_201 ();
 sg13g2_fill_1 FILLER_19_203 ();
 sg13g2_fill_1 FILLER_19_273 ();
 sg13g2_fill_1 FILLER_19_322 ();
 sg13g2_fill_1 FILLER_19_372 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_fill_2 FILLER_20_112 ();
 sg13g2_fill_1 FILLER_20_118 ();
 sg13g2_decap_4 FILLER_20_202 ();
 sg13g2_fill_2 FILLER_20_206 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_fill_1 FILLER_20_269 ();
 sg13g2_fill_2 FILLER_20_279 ();
 sg13g2_decap_4 FILLER_20_324 ();
 sg13g2_fill_1 FILLER_20_328 ();
 sg13g2_fill_2 FILLER_20_387 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_4 FILLER_21_98 ();
 sg13g2_fill_1 FILLER_21_102 ();
 sg13g2_fill_1 FILLER_21_138 ();
 sg13g2_decap_4 FILLER_21_165 ();
 sg13g2_decap_4 FILLER_21_182 ();
 sg13g2_fill_1 FILLER_21_186 ();
 sg13g2_fill_1 FILLER_21_223 ();
 sg13g2_fill_1 FILLER_21_237 ();
 sg13g2_fill_1 FILLER_21_256 ();
 sg13g2_fill_1 FILLER_21_333 ();
 sg13g2_fill_1 FILLER_21_353 ();
 sg13g2_fill_2 FILLER_21_364 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_fill_2 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_107 ();
 sg13g2_fill_1 FILLER_22_128 ();
 sg13g2_fill_2 FILLER_22_137 ();
 sg13g2_fill_1 FILLER_22_139 ();
 sg13g2_fill_2 FILLER_22_212 ();
 sg13g2_fill_1 FILLER_22_253 ();
 sg13g2_fill_2 FILLER_22_312 ();
 sg13g2_fill_1 FILLER_22_314 ();
 sg13g2_fill_2 FILLER_22_372 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_4 FILLER_23_105 ();
 sg13g2_fill_2 FILLER_23_154 ();
 sg13g2_fill_1 FILLER_23_156 ();
 sg13g2_fill_2 FILLER_23_170 ();
 sg13g2_fill_2 FILLER_23_198 ();
 sg13g2_fill_1 FILLER_23_216 ();
 sg13g2_fill_1 FILLER_23_238 ();
 sg13g2_fill_1 FILLER_23_264 ();
 sg13g2_fill_1 FILLER_23_279 ();
 sg13g2_decap_4 FILLER_23_321 ();
 sg13g2_fill_2 FILLER_23_325 ();
 sg13g2_fill_1 FILLER_23_360 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_4 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_102 ();
 sg13g2_fill_2 FILLER_24_112 ();
 sg13g2_fill_1 FILLER_24_114 ();
 sg13g2_fill_1 FILLER_24_132 ();
 sg13g2_fill_1 FILLER_24_319 ();
 sg13g2_fill_2 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_4 FILLER_25_49 ();
 sg13g2_fill_2 FILLER_25_53 ();
 sg13g2_decap_8 FILLER_25_81 ();
 sg13g2_fill_2 FILLER_25_92 ();
 sg13g2_fill_1 FILLER_25_94 ();
 sg13g2_fill_1 FILLER_25_157 ();
 sg13g2_fill_2 FILLER_25_176 ();
 sg13g2_fill_1 FILLER_25_212 ();
 sg13g2_fill_2 FILLER_25_224 ();
 sg13g2_fill_1 FILLER_25_261 ();
 sg13g2_fill_1 FILLER_25_319 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_4 FILLER_26_35 ();
 sg13g2_fill_1 FILLER_26_39 ();
 sg13g2_decap_4 FILLER_26_44 ();
 sg13g2_fill_2 FILLER_26_48 ();
 sg13g2_fill_2 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_65 ();
 sg13g2_fill_2 FILLER_26_70 ();
 sg13g2_fill_1 FILLER_26_72 ();
 sg13g2_fill_2 FILLER_26_134 ();
 sg13g2_fill_2 FILLER_26_184 ();
 sg13g2_fill_1 FILLER_26_186 ();
 sg13g2_fill_1 FILLER_26_226 ();
 sg13g2_fill_2 FILLER_26_287 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_fill_1 FILLER_26_303 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_fill_2 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_56 ();
 sg13g2_fill_1 FILLER_27_58 ();
 sg13g2_fill_2 FILLER_27_64 ();
 sg13g2_decap_8 FILLER_27_85 ();
 sg13g2_fill_2 FILLER_27_117 ();
 sg13g2_fill_1 FILLER_27_133 ();
 sg13g2_fill_2 FILLER_27_142 ();
 sg13g2_fill_1 FILLER_27_144 ();
 sg13g2_fill_1 FILLER_27_163 ();
 sg13g2_decap_4 FILLER_27_190 ();
 sg13g2_fill_2 FILLER_27_194 ();
 sg13g2_fill_1 FILLER_27_235 ();
 sg13g2_decap_8 FILLER_27_302 ();
 sg13g2_fill_2 FILLER_27_354 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_4 FILLER_28_21 ();
 sg13g2_fill_1 FILLER_28_25 ();
 sg13g2_fill_2 FILLER_28_81 ();
 sg13g2_fill_1 FILLER_28_83 ();
 sg13g2_fill_2 FILLER_28_119 ();
 sg13g2_decap_4 FILLER_28_181 ();
 sg13g2_fill_2 FILLER_28_185 ();
 sg13g2_fill_1 FILLER_28_247 ();
 sg13g2_fill_2 FILLER_28_271 ();
 sg13g2_fill_1 FILLER_28_283 ();
 sg13g2_decap_4 FILLER_28_297 ();
 sg13g2_fill_2 FILLER_28_314 ();
 sg13g2_fill_2 FILLER_28_328 ();
 sg13g2_fill_1 FILLER_28_380 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_fill_1 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_48 ();
 sg13g2_fill_1 FILLER_29_73 ();
 sg13g2_fill_2 FILLER_29_89 ();
 sg13g2_fill_1 FILLER_29_91 ();
 sg13g2_fill_2 FILLER_29_121 ();
 sg13g2_fill_2 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_142 ();
 sg13g2_fill_2 FILLER_29_199 ();
 sg13g2_fill_1 FILLER_29_201 ();
 sg13g2_fill_1 FILLER_29_246 ();
 sg13g2_fill_1 FILLER_29_277 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_47 ();
 sg13g2_fill_1 FILLER_30_75 ();
 sg13g2_decap_4 FILLER_30_90 ();
 sg13g2_fill_2 FILLER_30_135 ();
 sg13g2_fill_1 FILLER_30_151 ();
 sg13g2_fill_1 FILLER_30_243 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_277 ();
 sg13g2_fill_2 FILLER_30_287 ();
 sg13g2_fill_1 FILLER_30_293 ();
 sg13g2_fill_2 FILLER_30_303 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_fill_1 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_4 FILLER_31_14 ();
 sg13g2_fill_1 FILLER_31_18 ();
 sg13g2_fill_2 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_51 ();
 sg13g2_fill_2 FILLER_31_76 ();
 sg13g2_fill_1 FILLER_31_86 ();
 sg13g2_fill_2 FILLER_31_115 ();
 sg13g2_fill_1 FILLER_31_117 ();
 sg13g2_fill_1 FILLER_31_123 ();
 sg13g2_fill_2 FILLER_31_171 ();
 sg13g2_fill_1 FILLER_31_173 ();
 sg13g2_fill_1 FILLER_31_197 ();
 sg13g2_decap_4 FILLER_31_202 ();
 sg13g2_decap_4 FILLER_31_209 ();
 sg13g2_fill_2 FILLER_31_213 ();
 sg13g2_fill_1 FILLER_31_260 ();
 sg13g2_fill_1 FILLER_31_317 ();
 sg13g2_fill_1 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_fill_2 FILLER_32_61 ();
 sg13g2_fill_1 FILLER_32_63 ();
 sg13g2_fill_2 FILLER_32_78 ();
 sg13g2_fill_1 FILLER_32_80 ();
 sg13g2_fill_2 FILLER_32_114 ();
 sg13g2_fill_2 FILLER_32_128 ();
 sg13g2_fill_1 FILLER_32_130 ();
 sg13g2_fill_1 FILLER_32_145 ();
 sg13g2_fill_2 FILLER_32_172 ();
 sg13g2_fill_1 FILLER_32_174 ();
 sg13g2_fill_2 FILLER_32_222 ();
 sg13g2_fill_1 FILLER_32_254 ();
 sg13g2_fill_2 FILLER_32_261 ();
 sg13g2_fill_1 FILLER_32_344 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_16 ();
 sg13g2_fill_1 FILLER_33_47 ();
 sg13g2_fill_1 FILLER_33_80 ();
 sg13g2_fill_2 FILLER_33_119 ();
 sg13g2_fill_1 FILLER_33_121 ();
 sg13g2_fill_2 FILLER_33_132 ();
 sg13g2_fill_2 FILLER_33_155 ();
 sg13g2_fill_1 FILLER_33_157 ();
 sg13g2_fill_2 FILLER_33_162 ();
 sg13g2_fill_2 FILLER_33_173 ();
 sg13g2_fill_1 FILLER_33_175 ();
 sg13g2_fill_1 FILLER_33_232 ();
 sg13g2_fill_2 FILLER_33_236 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_fill_2 FILLER_33_276 ();
 sg13g2_fill_1 FILLER_33_350 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_4 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_25 ();
 sg13g2_fill_2 FILLER_34_53 ();
 sg13g2_fill_1 FILLER_34_55 ();
 sg13g2_fill_2 FILLER_34_66 ();
 sg13g2_fill_2 FILLER_34_82 ();
 sg13g2_fill_1 FILLER_34_84 ();
 sg13g2_fill_1 FILLER_34_94 ();
 sg13g2_fill_1 FILLER_34_113 ();
 sg13g2_fill_2 FILLER_34_141 ();
 sg13g2_fill_2 FILLER_34_155 ();
 sg13g2_fill_2 FILLER_34_185 ();
 sg13g2_fill_1 FILLER_34_195 ();
 sg13g2_fill_2 FILLER_34_228 ();
 sg13g2_fill_2 FILLER_34_284 ();
 sg13g2_fill_1 FILLER_34_309 ();
 sg13g2_fill_1 FILLER_34_333 ();
 sg13g2_fill_2 FILLER_34_343 ();
 sg13g2_fill_1 FILLER_34_345 ();
 sg13g2_fill_2 FILLER_34_358 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_4 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_32 ();
 sg13g2_fill_2 FILLER_35_60 ();
 sg13g2_fill_1 FILLER_35_76 ();
 sg13g2_fill_2 FILLER_35_174 ();
 sg13g2_fill_1 FILLER_35_176 ();
 sg13g2_fill_1 FILLER_35_187 ();
 sg13g2_fill_1 FILLER_35_249 ();
 sg13g2_fill_1 FILLER_35_254 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_fill_2 FILLER_36_42 ();
 sg13g2_decap_4 FILLER_36_48 ();
 sg13g2_fill_1 FILLER_36_56 ();
 sg13g2_fill_1 FILLER_36_93 ();
 sg13g2_fill_2 FILLER_36_156 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_fill_1 FILLER_36_254 ();
 sg13g2_fill_2 FILLER_36_298 ();
 sg13g2_fill_2 FILLER_36_310 ();
 sg13g2_fill_1 FILLER_36_347 ();
 sg13g2_fill_1 FILLER_36_378 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_fill_2 FILLER_37_64 ();
 sg13g2_fill_1 FILLER_37_66 ();
 sg13g2_fill_2 FILLER_37_135 ();
 sg13g2_fill_1 FILLER_37_137 ();
 sg13g2_fill_2 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_231 ();
 sg13g2_fill_1 FILLER_37_233 ();
 sg13g2_fill_1 FILLER_37_280 ();
 sg13g2_fill_2 FILLER_37_291 ();
 sg13g2_fill_1 FILLER_37_303 ();
 sg13g2_fill_2 FILLER_37_340 ();
 sg13g2_fill_1 FILLER_37_350 ();
 sg13g2_fill_2 FILLER_37_380 ();
 sg13g2_fill_1 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_fill_2 FILLER_38_68 ();
 sg13g2_fill_2 FILLER_38_154 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_fill_2 FILLER_38_187 ();
 sg13g2_fill_1 FILLER_38_215 ();
 sg13g2_fill_2 FILLER_38_254 ();
 sg13g2_fill_1 FILLER_38_256 ();
 sg13g2_fill_1 FILLER_38_269 ();
 sg13g2_fill_2 FILLER_38_283 ();
 sg13g2_fill_1 FILLER_38_285 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net10;
 assign uio_oe[1] = net11;
 assign uio_oe[2] = net12;
 assign uio_oe[3] = net13;
 assign uio_oe[4] = net14;
 assign uio_oe[5] = net15;
 assign uio_oe[6] = net16;
 assign uio_oe[7] = net17;
 assign uio_out[0] = net18;
 assign uio_out[1] = net19;
 assign uio_out[2] = net20;
 assign uio_out[3] = net21;
 assign uio_out[4] = net22;
 assign uio_out[5] = net23;
 assign uio_out[6] = net24;
 assign uio_out[7] = net25;
 assign uo_out[6] = net26;
 assign uo_out[7] = net27;
endmodule

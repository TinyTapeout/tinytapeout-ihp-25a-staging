module tt_um_asheldon44_dsm_decimation_filter (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \CIC.dec_clk ;
 wire \CIC.inc_out[0] ;
 wire \CIC.inc_out[10] ;
 wire \CIC.inc_out[11] ;
 wire \CIC.inc_out[12] ;
 wire \CIC.inc_out[13] ;
 wire \CIC.inc_out[14] ;
 wire \CIC.inc_out[15] ;
 wire \CIC.inc_out[16] ;
 wire \CIC.inc_out[17] ;
 wire \CIC.inc_out[18] ;
 wire \CIC.inc_out[19] ;
 wire \CIC.inc_out[1] ;
 wire \CIC.inc_out[20] ;
 wire \CIC.inc_out[21] ;
 wire \CIC.inc_out[22] ;
 wire \CIC.inc_out[23] ;
 wire \CIC.inc_out[2] ;
 wire \CIC.inc_out[3] ;
 wire \CIC.inc_out[4] ;
 wire \CIC.inc_out[5] ;
 wire \CIC.inc_out[6] ;
 wire \CIC.inc_out[7] ;
 wire \CIC.inc_out[8] ;
 wire \CIC.inc_out[9] ;
 wire \CIC.int_1_out[0] ;
 wire \CIC.int_1_out[10] ;
 wire \CIC.int_1_out[11] ;
 wire \CIC.int_1_out[12] ;
 wire \CIC.int_1_out[13] ;
 wire \CIC.int_1_out[14] ;
 wire \CIC.int_1_out[15] ;
 wire \CIC.int_1_out[16] ;
 wire \CIC.int_1_out[17] ;
 wire \CIC.int_1_out[18] ;
 wire \CIC.int_1_out[19] ;
 wire \CIC.int_1_out[1] ;
 wire \CIC.int_1_out[20] ;
 wire \CIC.int_1_out[21] ;
 wire \CIC.int_1_out[22] ;
 wire \CIC.int_1_out[23] ;
 wire \CIC.int_1_out[2] ;
 wire \CIC.int_1_out[3] ;
 wire \CIC.int_1_out[4] ;
 wire \CIC.int_1_out[5] ;
 wire \CIC.int_1_out[6] ;
 wire \CIC.int_1_out[7] ;
 wire \CIC.int_1_out[8] ;
 wire \CIC.int_1_out[9] ;
 wire \CIC.int_2_out[0] ;
 wire \CIC.int_2_out[10] ;
 wire \CIC.int_2_out[11] ;
 wire \CIC.int_2_out[12] ;
 wire \CIC.int_2_out[13] ;
 wire \CIC.int_2_out[14] ;
 wire \CIC.int_2_out[15] ;
 wire \CIC.int_2_out[16] ;
 wire \CIC.int_2_out[17] ;
 wire \CIC.int_2_out[18] ;
 wire \CIC.int_2_out[19] ;
 wire \CIC.int_2_out[1] ;
 wire \CIC.int_2_out[20] ;
 wire \CIC.int_2_out[21] ;
 wire \CIC.int_2_out[22] ;
 wire \CIC.int_2_out[23] ;
 wire \CIC.int_2_out[2] ;
 wire \CIC.int_2_out[3] ;
 wire \CIC.int_2_out[4] ;
 wire \CIC.int_2_out[5] ;
 wire \CIC.int_2_out[6] ;
 wire \CIC.int_2_out[7] ;
 wire \CIC.int_2_out[8] ;
 wire \CIC.int_2_out[9] ;
 wire \CIC.out[0] ;
 wire \CIC.out[10] ;
 wire \CIC.out[11] ;
 wire \CIC.out[12] ;
 wire \CIC.out[13] ;
 wire \CIC.out[14] ;
 wire \CIC.out[15] ;
 wire \CIC.out[16] ;
 wire \CIC.out[17] ;
 wire \CIC.out[18] ;
 wire \CIC.out[19] ;
 wire \CIC.out[1] ;
 wire \CIC.out[20] ;
 wire \CIC.out[21] ;
 wire \CIC.out[22] ;
 wire \CIC.out[23] ;
 wire \CIC.out[2] ;
 wire \CIC.out[3] ;
 wire \CIC.out[4] ;
 wire \CIC.out[5] ;
 wire \CIC.out[6] ;
 wire \CIC.out[7] ;
 wire \CIC.out[8] ;
 wire \CIC.out[9] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[0] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[10] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[11] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[12] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[13] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[14] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[15] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[16] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[17] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[18] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[19] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[1] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[20] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[21] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[22] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[23] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[2] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[3] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[4] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[5] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[6] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[7] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[8] ;
 wire \CIC.u_differentiator.a_mux4to1.d1[9] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[0] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[10] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[11] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[12] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[13] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[14] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[15] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[16] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[17] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[18] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[19] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[1] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[20] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[21] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[22] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[23] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[2] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[3] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[4] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[5] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[6] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[7] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[8] ;
 wire \CIC.u_differentiator.a_mux4to1.d2[9] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[0] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[10] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[11] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[12] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[13] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[14] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[15] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[16] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[17] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[18] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[19] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[1] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[20] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[21] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[22] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[23] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[2] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[3] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[4] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[5] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[6] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[7] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[8] ;
 wire \CIC.u_differentiator.a_mux4to1.d3[9] ;
 wire \CIC.u_differentiator.a_mux4to1.sel[0] ;
 wire \CIC.u_differentiator.a_mux4to1.sel[1] ;
 wire \CIC.u_differentiator.count[2] ;
 wire \CIC.u_differentiator.prev_lr_clk ;
 wire \CIC.u_differentiator.temp[0] ;
 wire \CIC.u_differentiator.temp[10] ;
 wire \CIC.u_differentiator.temp[11] ;
 wire \CIC.u_differentiator.temp[12] ;
 wire \CIC.u_differentiator.temp[13] ;
 wire \CIC.u_differentiator.temp[14] ;
 wire \CIC.u_differentiator.temp[15] ;
 wire \CIC.u_differentiator.temp[16] ;
 wire \CIC.u_differentiator.temp[17] ;
 wire \CIC.u_differentiator.temp[18] ;
 wire \CIC.u_differentiator.temp[19] ;
 wire \CIC.u_differentiator.temp[1] ;
 wire \CIC.u_differentiator.temp[20] ;
 wire \CIC.u_differentiator.temp[21] ;
 wire \CIC.u_differentiator.temp[22] ;
 wire \CIC.u_differentiator.temp[23] ;
 wire \CIC.u_differentiator.temp[2] ;
 wire \CIC.u_differentiator.temp[3] ;
 wire \CIC.u_differentiator.temp[4] ;
 wire \CIC.u_differentiator.temp[5] ;
 wire \CIC.u_differentiator.temp[6] ;
 wire \CIC.u_differentiator.temp[7] ;
 wire \CIC.u_differentiator.temp[8] ;
 wire \CIC.u_differentiator.temp[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire div_clk8x;
 wire \divideby64.clkOutDiv1 ;
 wire \divideby64.clkOutDiv2 ;
 wire \divideby64.clkOutDiv4 ;
 wire \divideby64.clkOutDiv5 ;
 wire \outmux.count[0] ;
 wire \outmux.count[1] ;
 wire \outmux.count[2] ;
 wire net39;
 wire net3;
 wire clknet_0_clk;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net1;
 wire net2;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;

 sg13g2_inv_1 _1104_ (.Y(_0448_),
    .A(net375));
 sg13g2_inv_2 _1105_ (.Y(_0449_),
    .A(net379));
 sg13g2_inv_1 _1106_ (.Y(_0450_),
    .A(\CIC.u_differentiator.a_mux4to1.d3[0] ));
 sg13g2_inv_1 _1107_ (.Y(_0451_),
    .A(\CIC.u_differentiator.a_mux4to1.d2[0] ));
 sg13g2_inv_1 _1108_ (.Y(_0452_),
    .A(\CIC.u_differentiator.a_mux4to1.d3[4] ));
 sg13g2_inv_1 _1109_ (.Y(_0453_),
    .A(\CIC.u_differentiator.a_mux4to1.d2[4] ));
 sg13g2_inv_1 _1110_ (.Y(_0454_),
    .A(\CIC.u_differentiator.a_mux4to1.d3[6] ));
 sg13g2_inv_1 _1111_ (.Y(_0455_),
    .A(\CIC.u_differentiator.a_mux4to1.d2[6] ));
 sg13g2_inv_1 _1112_ (.Y(_0456_),
    .A(\CIC.u_differentiator.a_mux4to1.d3[7] ));
 sg13g2_inv_1 _1113_ (.Y(_0457_),
    .A(\CIC.u_differentiator.a_mux4to1.d2[7] ));
 sg13g2_inv_1 _1114_ (.Y(_0458_),
    .A(\CIC.u_differentiator.a_mux4to1.d3[12] ));
 sg13g2_inv_1 _1115_ (.Y(_0459_),
    .A(\CIC.u_differentiator.a_mux4to1.d2[12] ));
 sg13g2_inv_1 _1116_ (.Y(_0460_),
    .A(\CIC.u_differentiator.a_mux4to1.d2[20] ));
 sg13g2_inv_1 _1117_ (.Y(_0461_),
    .A(\CIC.u_differentiator.a_mux4to1.d2[22] ));
 sg13g2_inv_1 _1118_ (.Y(_0462_),
    .A(net245));
 sg13g2_inv_1 _1119_ (.Y(_0463_),
    .A(\CIC.inc_out[22] ));
 sg13g2_inv_1 _1120_ (.Y(_0464_),
    .A(net230));
 sg13g2_inv_1 _1121_ (.Y(_0465_),
    .A(\CIC.u_differentiator.temp[7] ));
 sg13g2_inv_1 _1122_ (.Y(_0466_),
    .A(_0006_));
 sg13g2_inv_1 _1123_ (.Y(_0467_),
    .A(\CIC.u_differentiator.temp[11] ));
 sg13g2_inv_1 _1124_ (.Y(_0468_),
    .A(net218));
 sg13g2_inv_1 _1125_ (.Y(_0469_),
    .A(\CIC.u_differentiator.temp[14] ));
 sg13g2_inv_1 _1126_ (.Y(_0470_),
    .A(_0008_));
 sg13g2_inv_1 _1127_ (.Y(_0471_),
    .A(\CIC.u_differentiator.temp[15] ));
 sg13g2_inv_1 _1128_ (.Y(_0472_),
    .A(\CIC.u_differentiator.temp[21] ));
 sg13g2_nand3b_1 _1129_ (.B(\outmux.count[1] ),
    .C(_0010_),
    .Y(_0473_),
    .A_N(\outmux.count[0] ));
 sg13g2_nor2_1 _1130_ (.A(\CIC.out[16] ),
    .B(net349),
    .Y(_0474_));
 sg13g2_nand2_1 _1131_ (.Y(_0475_),
    .A(\outmux.count[0] ),
    .B(\outmux.count[1] ));
 sg13g2_nor2_2 _1132_ (.A(\outmux.count[2] ),
    .B(_0475_),
    .Y(_0476_));
 sg13g2_nor3_2 _1133_ (.A(\outmux.count[0] ),
    .B(\outmux.count[1] ),
    .C(_0010_),
    .Y(_0477_));
 sg13g2_a22oi_1 _1134_ (.Y(_0478_),
    .B1(_0477_),
    .B2(\CIC.out[0] ),
    .A2(_0476_),
    .A1(\CIC.out[8] ));
 sg13g2_a21oi_1 _1135_ (.A1(net349),
    .A2(_0478_),
    .Y(uo_out[0]),
    .B1(_0474_));
 sg13g2_nor2_1 _1136_ (.A(\CIC.out[17] ),
    .B(net349),
    .Y(_0479_));
 sg13g2_a22oi_1 _1137_ (.Y(_0480_),
    .B1(_0477_),
    .B2(\CIC.out[1] ),
    .A2(_0476_),
    .A1(\CIC.out[9] ));
 sg13g2_a21oi_1 _1138_ (.A1(net349),
    .A2(_0480_),
    .Y(uo_out[1]),
    .B1(_0479_));
 sg13g2_nor2_1 _1139_ (.A(\CIC.out[18] ),
    .B(net349),
    .Y(_0481_));
 sg13g2_a22oi_1 _1140_ (.Y(_0482_),
    .B1(_0477_),
    .B2(\CIC.out[2] ),
    .A2(_0476_),
    .A1(\CIC.out[10] ));
 sg13g2_a21oi_1 _1141_ (.A1(net349),
    .A2(_0482_),
    .Y(uo_out[2]),
    .B1(_0481_));
 sg13g2_nor2_1 _1142_ (.A(\CIC.out[19] ),
    .B(net348),
    .Y(_0483_));
 sg13g2_a22oi_1 _1143_ (.Y(_0484_),
    .B1(_0477_),
    .B2(\CIC.out[3] ),
    .A2(_0476_),
    .A1(\CIC.out[11] ));
 sg13g2_a21oi_2 _1144_ (.B1(_0483_),
    .Y(uo_out[3]),
    .A2(_0484_),
    .A1(net349));
 sg13g2_a22oi_1 _1145_ (.Y(_0485_),
    .B1(_0477_),
    .B2(\CIC.out[4] ),
    .A2(_0476_),
    .A1(\CIC.out[12] ));
 sg13g2_nor2_1 _1146_ (.A(\CIC.out[20] ),
    .B(net348),
    .Y(_0486_));
 sg13g2_a21oi_1 _1147_ (.A1(_0473_),
    .A2(_0485_),
    .Y(uo_out[4]),
    .B1(_0486_));
 sg13g2_nor2_1 _1148_ (.A(\CIC.out[21] ),
    .B(net348),
    .Y(_0487_));
 sg13g2_a22oi_1 _1149_ (.Y(_0488_),
    .B1(_0477_),
    .B2(\CIC.out[5] ),
    .A2(_0476_),
    .A1(\CIC.out[13] ));
 sg13g2_a21oi_2 _1150_ (.B1(_0487_),
    .Y(uo_out[5]),
    .A2(_0488_),
    .A1(net348));
 sg13g2_nor2_1 _1151_ (.A(\CIC.out[22] ),
    .B(net348),
    .Y(_0489_));
 sg13g2_a22oi_1 _1152_ (.Y(_0490_),
    .B1(_0477_),
    .B2(\CIC.out[6] ),
    .A2(_0476_),
    .A1(\CIC.out[14] ));
 sg13g2_a21oi_1 _1153_ (.A1(net348),
    .A2(_0490_),
    .Y(uo_out[6]),
    .B1(_0489_));
 sg13g2_nor2_1 _1154_ (.A(\CIC.out[23] ),
    .B(net348),
    .Y(_0491_));
 sg13g2_a22oi_1 _1155_ (.Y(_0492_),
    .B1(_0477_),
    .B2(\CIC.out[7] ),
    .A2(_0476_),
    .A1(\CIC.out[15] ));
 sg13g2_a21oi_2 _1156_ (.B1(_0491_),
    .Y(uo_out[7]),
    .A2(_0492_),
    .A1(net348));
 sg13g2_xor2_1 _1157_ (.B(net1),
    .A(net255),
    .X(_0034_));
 sg13g2_nand3_1 _1158_ (.B(net1),
    .C(net301),
    .A(net255),
    .Y(_0493_));
 sg13g2_a21o_1 _1159_ (.A2(net1),
    .A1(net255),
    .B1(net301),
    .X(_0494_));
 sg13g2_and2_1 _1160_ (.A(_0493_),
    .B(_0494_),
    .X(_0045_));
 sg13g2_and4_2 _1161_ (.A(net442),
    .B(net1),
    .C(\CIC.inc_out[1] ),
    .D(net168),
    .X(_0495_));
 sg13g2_xnor2_1 _1162_ (.Y(_0050_),
    .A(net168),
    .B(_0493_));
 sg13g2_xor2_1 _1163_ (.B(net443),
    .A(net252),
    .X(_0051_));
 sg13g2_and3_1 _1164_ (.X(_0496_),
    .A(\CIC.inc_out[3] ),
    .B(net116),
    .C(_0495_));
 sg13g2_a21oi_1 _1165_ (.A1(\CIC.inc_out[3] ),
    .A2(_0495_),
    .Y(_0497_),
    .B1(net116));
 sg13g2_nor2_1 _1166_ (.A(_0496_),
    .B(net117),
    .Y(_0052_));
 sg13g2_xor2_1 _1167_ (.B(_0496_),
    .A(net187),
    .X(_0053_));
 sg13g2_and3_1 _1168_ (.X(_0498_),
    .A(net187),
    .B(net159),
    .C(_0496_));
 sg13g2_a21oi_1 _1169_ (.A1(\CIC.inc_out[5] ),
    .A2(_0496_),
    .Y(_0499_),
    .B1(net159));
 sg13g2_nor2_1 _1170_ (.A(_0498_),
    .B(net160),
    .Y(_0054_));
 sg13g2_xor2_1 _1171_ (.B(_0498_),
    .A(net238),
    .X(_0055_));
 sg13g2_and3_1 _1172_ (.X(_0500_),
    .A(net238),
    .B(net205),
    .C(_0498_));
 sg13g2_a21oi_1 _1173_ (.A1(\CIC.inc_out[7] ),
    .A2(_0498_),
    .Y(_0501_),
    .B1(net205));
 sg13g2_nor2_1 _1174_ (.A(_0500_),
    .B(net206),
    .Y(_0056_));
 sg13g2_xor2_1 _1175_ (.B(_0500_),
    .A(net253),
    .X(_0057_));
 sg13g2_and3_1 _1176_ (.X(_0502_),
    .A(net436),
    .B(net152),
    .C(_0500_));
 sg13g2_a21oi_1 _1177_ (.A1(\CIC.inc_out[9] ),
    .A2(_0500_),
    .Y(_0503_),
    .B1(net152));
 sg13g2_nor2_1 _1178_ (.A(_0502_),
    .B(net153),
    .Y(_0035_));
 sg13g2_xor2_1 _1179_ (.B(_0502_),
    .A(net261),
    .X(_0036_));
 sg13g2_and3_1 _1180_ (.X(_0504_),
    .A(net444),
    .B(net174),
    .C(_0502_));
 sg13g2_a21oi_1 _1181_ (.A1(\CIC.inc_out[11] ),
    .A2(_0502_),
    .Y(_0505_),
    .B1(net174));
 sg13g2_nor2_1 _1182_ (.A(_0504_),
    .B(net175),
    .Y(_0037_));
 sg13g2_xor2_1 _1183_ (.B(_0504_),
    .A(net254),
    .X(_0038_));
 sg13g2_nand3_1 _1184_ (.B(net269),
    .C(_0504_),
    .A(net254),
    .Y(_0506_));
 sg13g2_a21o_1 _1185_ (.A2(_0504_),
    .A1(net254),
    .B1(net269),
    .X(_0507_));
 sg13g2_and2_1 _1186_ (.A(_0506_),
    .B(_0507_),
    .X(_0039_));
 sg13g2_nor2_1 _1187_ (.A(_0462_),
    .B(_0506_),
    .Y(_0508_));
 sg13g2_xnor2_1 _1188_ (.Y(_0040_),
    .A(net245),
    .B(_0506_));
 sg13g2_and2_1 _1189_ (.A(net247),
    .B(_0508_),
    .X(_0509_));
 sg13g2_xor2_1 _1190_ (.B(_0508_),
    .A(net247),
    .X(_0041_));
 sg13g2_xor2_1 _1191_ (.B(_0509_),
    .A(net258),
    .X(_0042_));
 sg13g2_and3_2 _1192_ (.X(_0510_),
    .A(net445),
    .B(net138),
    .C(_0509_));
 sg13g2_a21oi_1 _1193_ (.A1(\CIC.inc_out[17] ),
    .A2(_0509_),
    .Y(_0511_),
    .B1(net138));
 sg13g2_nor2_1 _1194_ (.A(_0510_),
    .B(net139),
    .Y(_0043_));
 sg13g2_xor2_1 _1195_ (.B(_0510_),
    .A(net263),
    .X(_0044_));
 sg13g2_nand3_1 _1196_ (.B(net287),
    .C(_0510_),
    .A(net263),
    .Y(_0512_));
 sg13g2_a21o_1 _1197_ (.A2(_0510_),
    .A1(net263),
    .B1(net287),
    .X(_0513_));
 sg13g2_and2_1 _1198_ (.A(_0512_),
    .B(_0513_),
    .X(_0046_));
 sg13g2_nand4_1 _1199_ (.B(\CIC.inc_out[20] ),
    .C(\CIC.inc_out[21] ),
    .A(\CIC.inc_out[19] ),
    .Y(_0514_),
    .D(_0510_));
 sg13g2_xnor2_1 _1200_ (.Y(_0047_),
    .A(net256),
    .B(_0512_));
 sg13g2_nor2_1 _1201_ (.A(_0463_),
    .B(_0514_),
    .Y(_0515_));
 sg13g2_xnor2_1 _1202_ (.Y(_0048_),
    .A(net250),
    .B(_0514_));
 sg13g2_xor2_1 _1203_ (.B(_0515_),
    .A(net72),
    .X(_0049_));
 sg13g2_xor2_1 _1204_ (.B(\outmux.count[1] ),
    .A(\outmux.count[0] ),
    .X(_0106_));
 sg13g2_xnor2_1 _1205_ (.Y(_0107_),
    .A(\outmux.count[2] ),
    .B(_0475_));
 sg13g2_nand2_1 _1206_ (.Y(_0516_),
    .A(net93),
    .B(net170));
 sg13g2_nand2_1 _1207_ (.Y(_0517_),
    .A(net259),
    .B(\CIC.int_1_out[1] ));
 sg13g2_nor2_1 _1208_ (.A(\CIC.int_2_out[1] ),
    .B(\CIC.int_1_out[1] ),
    .Y(_0518_));
 sg13g2_xor2_1 _1209_ (.B(\CIC.int_1_out[1] ),
    .A(net259),
    .X(_0519_));
 sg13g2_xnor2_1 _1210_ (.Y(_0093_),
    .A(_0516_),
    .B(net260));
 sg13g2_and2_1 _1211_ (.A(net172),
    .B(\CIC.int_1_out[2] ),
    .X(_0520_));
 sg13g2_xor2_1 _1212_ (.B(net423),
    .A(net172),
    .X(_0521_));
 sg13g2_o21ai_1 _1213_ (.B1(_0517_),
    .Y(_0522_),
    .A1(_0516_),
    .A2(_0518_));
 sg13g2_xor2_1 _1214_ (.B(_0522_),
    .A(_0521_),
    .X(_0098_));
 sg13g2_a21oi_2 _1215_ (.B1(_0520_),
    .Y(_0523_),
    .A2(_0522_),
    .A1(_0521_));
 sg13g2_nand2_1 _1216_ (.Y(_0524_),
    .A(net272),
    .B(net278));
 sg13g2_xnor2_1 _1217_ (.Y(_0525_),
    .A(net272),
    .B(\CIC.int_1_out[3] ));
 sg13g2_xor2_1 _1218_ (.B(net273),
    .A(_0523_),
    .X(_0099_));
 sg13g2_and2_1 _1219_ (.A(net216),
    .B(\CIC.int_1_out[4] ),
    .X(_0526_));
 sg13g2_xor2_1 _1220_ (.B(net298),
    .A(net216),
    .X(_0527_));
 sg13g2_o21ai_1 _1221_ (.B1(_0524_),
    .Y(_0528_),
    .A1(_0523_),
    .A2(_0525_));
 sg13g2_xor2_1 _1222_ (.B(_0528_),
    .A(_0527_),
    .X(_0100_));
 sg13g2_nor2_1 _1223_ (.A(net432),
    .B(\CIC.int_1_out[5] ),
    .Y(_0529_));
 sg13g2_xor2_1 _1224_ (.B(\CIC.int_1_out[5] ),
    .A(net280),
    .X(_0530_));
 sg13g2_a21oi_1 _1225_ (.A1(_0527_),
    .A2(_0528_),
    .Y(_0531_),
    .B1(_0526_));
 sg13g2_xnor2_1 _1226_ (.Y(_0101_),
    .A(net281),
    .B(_0531_));
 sg13g2_and2_1 _1227_ (.A(net140),
    .B(net454),
    .X(_0532_));
 sg13g2_xnor2_1 _1228_ (.Y(_0533_),
    .A(net140),
    .B(\CIC.int_1_out[6] ));
 sg13g2_a221oi_1 _1229_ (.B2(_0528_),
    .C1(_0526_),
    .B1(_0527_),
    .A1(\CIC.int_2_out[5] ),
    .Y(_0534_),
    .A2(\CIC.int_1_out[5] ));
 sg13g2_nor3_2 _1230_ (.A(_0529_),
    .B(_0533_),
    .C(_0534_),
    .Y(_0535_));
 sg13g2_o21ai_1 _1231_ (.B1(_0533_),
    .Y(_0536_),
    .A1(_0529_),
    .A2(_0534_));
 sg13g2_nor2b_1 _1232_ (.A(_0535_),
    .B_N(_0536_),
    .Y(_0102_));
 sg13g2_nor2_1 _1233_ (.A(_0532_),
    .B(_0535_),
    .Y(_0537_));
 sg13g2_nand2_1 _1234_ (.Y(_0538_),
    .A(net285),
    .B(\CIC.int_1_out[7] ));
 sg13g2_xor2_1 _1235_ (.B(net275),
    .A(net199),
    .X(_0539_));
 sg13g2_o21ai_1 _1236_ (.B1(_0539_),
    .Y(_0540_),
    .A1(_0532_),
    .A2(_0535_));
 sg13g2_xnor2_1 _1237_ (.Y(_0103_),
    .A(_0537_),
    .B(_0539_));
 sg13g2_nand2_1 _1238_ (.Y(_0541_),
    .A(net286),
    .B(_0540_));
 sg13g2_nand2_1 _1239_ (.Y(_0542_),
    .A(net197),
    .B(net276));
 sg13g2_xnor2_1 _1240_ (.Y(_0543_),
    .A(net197),
    .B(net276));
 sg13g2_nand2b_1 _1241_ (.Y(_0544_),
    .B(_0541_),
    .A_N(_0543_));
 sg13g2_xnor2_1 _1242_ (.Y(_0104_),
    .A(_0541_),
    .B(_0543_));
 sg13g2_nor2_1 _1243_ (.A(net283),
    .B(\CIC.int_1_out[9] ),
    .Y(_0545_));
 sg13g2_nand2_1 _1244_ (.Y(_0546_),
    .A(net283),
    .B(\CIC.int_1_out[9] ));
 sg13g2_nand2b_1 _1245_ (.Y(_0547_),
    .B(net284),
    .A_N(_0545_));
 sg13g2_nand2_1 _1246_ (.Y(_0548_),
    .A(_0542_),
    .B(_0544_));
 sg13g2_xnor2_1 _1247_ (.Y(_0105_),
    .A(_0547_),
    .B(_0548_));
 sg13g2_nand2_1 _1248_ (.Y(_0549_),
    .A(net185),
    .B(net292));
 sg13g2_xor2_1 _1249_ (.B(net292),
    .A(net185),
    .X(_0550_));
 sg13g2_inv_1 _1250_ (.Y(_0551_),
    .A(_0550_));
 sg13g2_o21ai_1 _1251_ (.B1(_0546_),
    .Y(_0552_),
    .A1(_0542_),
    .A2(_0545_));
 sg13g2_nor2_1 _1252_ (.A(_0543_),
    .B(_0547_),
    .Y(_0553_));
 sg13g2_a21oi_1 _1253_ (.A1(_0541_),
    .A2(_0553_),
    .Y(_0554_),
    .B1(_0552_));
 sg13g2_xnor2_1 _1254_ (.Y(_0083_),
    .A(_0550_),
    .B(_0554_));
 sg13g2_nor2_1 _1255_ (.A(net241),
    .B(\CIC.int_1_out[11] ),
    .Y(_0555_));
 sg13g2_nand2_1 _1256_ (.Y(_0556_),
    .A(net241),
    .B(net293));
 sg13g2_nand2b_1 _1257_ (.Y(_0557_),
    .B(_0556_),
    .A_N(_0555_));
 sg13g2_o21ai_1 _1258_ (.B1(_0549_),
    .Y(_0558_),
    .A1(_0551_),
    .A2(_0554_));
 sg13g2_xnor2_1 _1259_ (.Y(_0084_),
    .A(net294),
    .B(_0558_));
 sg13g2_nand2_1 _1260_ (.Y(_0559_),
    .A(net417),
    .B(net296));
 sg13g2_xor2_1 _1261_ (.B(\CIC.int_1_out[12] ),
    .A(\CIC.int_2_out[12] ),
    .X(_0560_));
 sg13g2_nor2_1 _1262_ (.A(_0551_),
    .B(_0557_),
    .Y(_0561_));
 sg13g2_o21ai_1 _1263_ (.B1(_0556_),
    .Y(_0562_),
    .A1(_0549_),
    .A2(_0555_));
 sg13g2_a21oi_1 _1264_ (.A1(_0552_),
    .A2(_0561_),
    .Y(_0563_),
    .B1(_0562_));
 sg13g2_inv_1 _1265_ (.Y(_0564_),
    .A(_0563_));
 sg13g2_nand2_1 _1266_ (.Y(_0565_),
    .A(_0553_),
    .B(_0561_));
 sg13g2_a21oi_2 _1267_ (.B1(_0565_),
    .Y(_0566_),
    .A2(_0540_),
    .A1(_0538_));
 sg13g2_o21ai_1 _1268_ (.B1(_0560_),
    .Y(_0567_),
    .A1(_0564_),
    .A2(_0566_));
 sg13g2_or3_1 _1269_ (.A(_0560_),
    .B(_0564_),
    .C(_0566_),
    .X(_0568_));
 sg13g2_and2_1 _1270_ (.A(_0567_),
    .B(_0568_),
    .X(_0085_));
 sg13g2_nor2_1 _1271_ (.A(net430),
    .B(\CIC.int_1_out[13] ),
    .Y(_0569_));
 sg13g2_xor2_1 _1272_ (.B(\CIC.int_1_out[13] ),
    .A(\CIC.int_2_out[13] ),
    .X(_0570_));
 sg13g2_nand2_1 _1273_ (.Y(_0571_),
    .A(_0559_),
    .B(_0567_));
 sg13g2_xor2_1 _1274_ (.B(_0571_),
    .A(_0570_),
    .X(_0086_));
 sg13g2_nand2_1 _1275_ (.Y(_0572_),
    .A(net226),
    .B(net305));
 sg13g2_xor2_1 _1276_ (.B(net305),
    .A(net226),
    .X(_0573_));
 sg13g2_a22oi_1 _1277_ (.Y(_0574_),
    .B1(\CIC.int_2_out[13] ),
    .B2(\CIC.int_1_out[13] ),
    .A2(\CIC.int_1_out[12] ),
    .A1(\CIC.int_2_out[12] ));
 sg13g2_a21oi_1 _1278_ (.A1(_0567_),
    .A2(_0574_),
    .Y(_0575_),
    .B1(_0569_));
 sg13g2_nand2_1 _1279_ (.Y(_0576_),
    .A(_0573_),
    .B(_0575_));
 sg13g2_xor2_1 _1280_ (.B(_0575_),
    .A(_0573_),
    .X(_0087_));
 sg13g2_nor2_1 _1281_ (.A(\CIC.int_2_out[15] ),
    .B(\CIC.int_1_out[15] ),
    .Y(_0577_));
 sg13g2_xor2_1 _1282_ (.B(\CIC.int_1_out[15] ),
    .A(net421),
    .X(_0578_));
 sg13g2_nand2_1 _1283_ (.Y(_0579_),
    .A(_0572_),
    .B(_0576_));
 sg13g2_xor2_1 _1284_ (.B(_0579_),
    .A(net422),
    .X(_0088_));
 sg13g2_nand2_1 _1285_ (.Y(_0580_),
    .A(net236),
    .B(net452));
 sg13g2_nor2_1 _1286_ (.A(net236),
    .B(net452),
    .Y(_0581_));
 sg13g2_or2_1 _1287_ (.X(_0582_),
    .B(\CIC.int_1_out[16] ),
    .A(net434));
 sg13g2_and2_1 _1288_ (.A(_0580_),
    .B(_0582_),
    .X(_0583_));
 sg13g2_and2_1 _1289_ (.A(_0573_),
    .B(_0578_),
    .X(_0584_));
 sg13g2_nor2_1 _1290_ (.A(_0569_),
    .B(_0574_),
    .Y(_0585_));
 sg13g2_nor2_1 _1291_ (.A(_0572_),
    .B(_0577_),
    .Y(_0586_));
 sg13g2_a221oi_1 _1292_ (.B2(_0585_),
    .C1(_0586_),
    .B1(_0584_),
    .A1(\CIC.int_2_out[15] ),
    .Y(_0587_),
    .A2(\CIC.int_1_out[15] ));
 sg13g2_nand3_1 _1293_ (.B(_0570_),
    .C(_0584_),
    .A(_0560_),
    .Y(_0588_));
 sg13g2_nand2_1 _1294_ (.Y(_0589_),
    .A(_0587_),
    .B(_0588_));
 sg13g2_nand2_1 _1295_ (.Y(_0590_),
    .A(_0563_),
    .B(_0587_));
 sg13g2_o21ai_1 _1296_ (.B1(_0589_),
    .Y(_0591_),
    .A1(_0566_),
    .A2(_0590_));
 sg13g2_xnor2_1 _1297_ (.Y(_0089_),
    .A(net435),
    .B(_0591_));
 sg13g2_nand2_1 _1298_ (.Y(_0592_),
    .A(\CIC.int_2_out[17] ),
    .B(\CIC.int_1_out[17] ));
 sg13g2_xnor2_1 _1299_ (.Y(_0593_),
    .A(net290),
    .B(\CIC.int_1_out[17] ));
 sg13g2_o21ai_1 _1300_ (.B1(_0580_),
    .Y(_0594_),
    .A1(_0581_),
    .A2(_0591_));
 sg13g2_xnor2_1 _1301_ (.Y(_0090_),
    .A(net291),
    .B(_0594_));
 sg13g2_nand2_1 _1302_ (.Y(_0595_),
    .A(net212),
    .B(net289));
 sg13g2_xnor2_1 _1303_ (.Y(_0596_),
    .A(net212),
    .B(net289));
 sg13g2_nand2_1 _1304_ (.Y(_0597_),
    .A(_0580_),
    .B(_0592_));
 sg13g2_o21ai_1 _1305_ (.B1(_0597_),
    .Y(_0598_),
    .A1(net300),
    .A2(\CIC.int_1_out[17] ));
 sg13g2_nand3b_1 _1306_ (.B(_0582_),
    .C(_0580_),
    .Y(_0599_),
    .A_N(_0593_));
 sg13g2_o21ai_1 _1307_ (.B1(_0598_),
    .Y(_0600_),
    .A1(_0591_),
    .A2(_0599_));
 sg13g2_nand2b_1 _1308_ (.Y(_0601_),
    .B(_0600_),
    .A_N(_0596_));
 sg13g2_xnor2_1 _1309_ (.Y(_0091_),
    .A(_0596_),
    .B(_0600_));
 sg13g2_nor2_1 _1310_ (.A(net150),
    .B(\CIC.int_1_out[19] ),
    .Y(_0602_));
 sg13g2_nand2_1 _1311_ (.Y(_0603_),
    .A(net150),
    .B(\CIC.int_1_out[19] ));
 sg13g2_nor2b_1 _1312_ (.A(_0602_),
    .B_N(_0603_),
    .Y(_0604_));
 sg13g2_and2_1 _1313_ (.A(_0595_),
    .B(_0601_),
    .X(_0605_));
 sg13g2_xnor2_1 _1314_ (.Y(_0092_),
    .A(_0604_),
    .B(_0605_));
 sg13g2_nand2b_1 _1315_ (.Y(_0606_),
    .B(_0604_),
    .A_N(_0596_));
 sg13g2_or2_1 _1316_ (.X(_0607_),
    .B(_0606_),
    .A(_0599_));
 sg13g2_o21ai_1 _1317_ (.B1(_0603_),
    .Y(_0608_),
    .A1(_0595_),
    .A2(_0602_));
 sg13g2_nor2_1 _1318_ (.A(_0598_),
    .B(_0606_),
    .Y(_0609_));
 sg13g2_nor2_1 _1319_ (.A(_0608_),
    .B(_0609_),
    .Y(_0610_));
 sg13g2_o21ai_1 _1320_ (.B1(_0610_),
    .Y(_0611_),
    .A1(_0591_),
    .A2(_0607_));
 sg13g2_and2_1 _1321_ (.A(net243),
    .B(net419),
    .X(_0612_));
 sg13g2_xor2_1 _1322_ (.B(net419),
    .A(net243),
    .X(_0613_));
 sg13g2_xor2_1 _1323_ (.B(_0613_),
    .A(_0611_),
    .X(_0094_));
 sg13g2_or2_1 _1324_ (.X(_0614_),
    .B(\CIC.int_1_out[21] ),
    .A(\CIC.int_2_out[21] ));
 sg13g2_and2_1 _1325_ (.A(net214),
    .B(\CIC.int_1_out[21] ),
    .X(_0615_));
 sg13g2_xor2_1 _1326_ (.B(\CIC.int_1_out[21] ),
    .A(net214),
    .X(_0616_));
 sg13g2_a21oi_1 _1327_ (.A1(_0611_),
    .A2(_0613_),
    .Y(_0617_),
    .B1(_0612_));
 sg13g2_xnor2_1 _1328_ (.Y(_0095_),
    .A(_0616_),
    .B(_0617_));
 sg13g2_nand2_1 _1329_ (.Y(_0618_),
    .A(net234),
    .B(net446));
 sg13g2_nor2_1 _1330_ (.A(net234),
    .B(net451),
    .Y(_0619_));
 sg13g2_xor2_1 _1331_ (.B(net270),
    .A(net234),
    .X(_0620_));
 sg13g2_and2_1 _1332_ (.A(_0613_),
    .B(_0616_),
    .X(_0621_));
 sg13g2_a221oi_1 _1333_ (.B2(_0611_),
    .C1(_0615_),
    .B1(_0621_),
    .A1(_0612_),
    .Y(_0622_),
    .A2(_0614_));
 sg13g2_xnor2_1 _1334_ (.Y(_0096_),
    .A(_0620_),
    .B(_0622_));
 sg13g2_o21ai_1 _1335_ (.B1(_0618_),
    .Y(_0623_),
    .A1(_0619_),
    .A2(_0622_));
 sg13g2_xnor2_1 _1336_ (.Y(_0624_),
    .A(net95),
    .B(net249));
 sg13g2_xnor2_1 _1337_ (.Y(_0097_),
    .A(_0623_),
    .B(_0624_));
 sg13g2_xor2_1 _1338_ (.B(\CIC.int_1_out[0] ),
    .A(net93),
    .X(_0082_));
 sg13g2_nand2_1 _1339_ (.Y(_0625_),
    .A(net255),
    .B(net170));
 sg13g2_nand2_1 _1340_ (.Y(_0626_),
    .A(net301),
    .B(net266));
 sg13g2_nor2_1 _1341_ (.A(\CIC.inc_out[1] ),
    .B(\CIC.int_1_out[1] ),
    .Y(_0627_));
 sg13g2_xor2_1 _1342_ (.B(net266),
    .A(\CIC.inc_out[1] ),
    .X(_0628_));
 sg13g2_xnor2_1 _1343_ (.Y(_0069_),
    .A(_0625_),
    .B(net267));
 sg13g2_and2_1 _1344_ (.A(net168),
    .B(net437),
    .X(_0629_));
 sg13g2_or2_1 _1345_ (.X(_0630_),
    .B(net423),
    .A(net168));
 sg13g2_nand2b_1 _1346_ (.Y(_0631_),
    .B(_0630_),
    .A_N(_0629_));
 sg13g2_o21ai_1 _1347_ (.B1(_0626_),
    .Y(_0632_),
    .A1(_0625_),
    .A2(_0627_));
 sg13g2_xnor2_1 _1348_ (.Y(_0074_),
    .A(_0631_),
    .B(_0632_));
 sg13g2_a21oi_2 _1349_ (.B1(_0629_),
    .Y(_0633_),
    .A2(_0632_),
    .A1(_0630_));
 sg13g2_nand2_1 _1350_ (.Y(_0634_),
    .A(net431),
    .B(net278));
 sg13g2_xnor2_1 _1351_ (.Y(_0635_),
    .A(net252),
    .B(net278));
 sg13g2_xor2_1 _1352_ (.B(_0635_),
    .A(_0633_),
    .X(_0075_));
 sg13g2_nand2_1 _1353_ (.Y(_0636_),
    .A(net116),
    .B(net298));
 sg13g2_xor2_1 _1354_ (.B(net298),
    .A(net116),
    .X(_0637_));
 sg13g2_o21ai_1 _1355_ (.B1(_0634_),
    .Y(_0638_),
    .A1(_0633_),
    .A2(_0635_));
 sg13g2_nand2_1 _1356_ (.Y(_0639_),
    .A(_0637_),
    .B(_0638_));
 sg13g2_xor2_1 _1357_ (.B(_0638_),
    .A(_0637_),
    .X(_0076_));
 sg13g2_nor2_1 _1358_ (.A(net438),
    .B(\CIC.int_1_out[5] ),
    .Y(_0640_));
 sg13g2_nand2_1 _1359_ (.Y(_0641_),
    .A(net187),
    .B(\CIC.int_1_out[5] ));
 sg13g2_nand2b_1 _1360_ (.Y(_0642_),
    .B(_0641_),
    .A_N(_0640_));
 sg13g2_nand2_1 _1361_ (.Y(_0643_),
    .A(_0636_),
    .B(_0639_));
 sg13g2_xnor2_1 _1362_ (.Y(_0077_),
    .A(_0642_),
    .B(_0643_));
 sg13g2_and2_1 _1363_ (.A(net159),
    .B(net295),
    .X(_0644_));
 sg13g2_xnor2_1 _1364_ (.Y(_0645_),
    .A(net159),
    .B(\CIC.int_1_out[6] ));
 sg13g2_nand2_1 _1365_ (.Y(_0646_),
    .A(_0636_),
    .B(_0641_));
 sg13g2_a21oi_1 _1366_ (.A1(_0637_),
    .A2(_0638_),
    .Y(_0647_),
    .B1(_0646_));
 sg13g2_nor3_2 _1367_ (.A(_0640_),
    .B(_0645_),
    .C(_0647_),
    .Y(_0648_));
 sg13g2_o21ai_1 _1368_ (.B1(_0645_),
    .Y(_0649_),
    .A1(_0640_),
    .A2(_0647_));
 sg13g2_nor2b_1 _1369_ (.A(_0648_),
    .B_N(_0649_),
    .Y(_0078_));
 sg13g2_nor2_1 _1370_ (.A(_0644_),
    .B(_0648_),
    .Y(_0650_));
 sg13g2_nand2_1 _1371_ (.Y(_0651_),
    .A(net425),
    .B(\CIC.int_1_out[7] ));
 sg13g2_xor2_1 _1372_ (.B(net275),
    .A(net238),
    .X(_0652_));
 sg13g2_o21ai_1 _1373_ (.B1(_0652_),
    .Y(_0653_),
    .A1(_0644_),
    .A2(_0648_));
 sg13g2_xnor2_1 _1374_ (.Y(_0079_),
    .A(_0650_),
    .B(_0652_));
 sg13g2_nand2_1 _1375_ (.Y(_0654_),
    .A(net426),
    .B(_0653_));
 sg13g2_nand2_1 _1376_ (.Y(_0655_),
    .A(net205),
    .B(net276));
 sg13g2_xnor2_1 _1377_ (.Y(_0656_),
    .A(net205),
    .B(net276));
 sg13g2_nand2b_1 _1378_ (.Y(_0657_),
    .B(_0654_),
    .A_N(_0656_));
 sg13g2_xnor2_1 _1379_ (.Y(_0080_),
    .A(_0654_),
    .B(_0656_));
 sg13g2_nor2_1 _1380_ (.A(\CIC.inc_out[9] ),
    .B(\CIC.int_1_out[9] ),
    .Y(_0658_));
 sg13g2_xnor2_1 _1381_ (.Y(_0659_),
    .A(net253),
    .B(\CIC.int_1_out[9] ));
 sg13g2_nand2_1 _1382_ (.Y(_0660_),
    .A(_0655_),
    .B(_0657_));
 sg13g2_xnor2_1 _1383_ (.Y(_0081_),
    .A(_0659_),
    .B(_0660_));
 sg13g2_and2_1 _1384_ (.A(net152),
    .B(net292),
    .X(_0661_));
 sg13g2_xor2_1 _1385_ (.B(net292),
    .A(net152),
    .X(_0662_));
 sg13g2_a22oi_1 _1386_ (.Y(_0663_),
    .B1(\CIC.int_1_out[9] ),
    .B2(\CIC.inc_out[9] ),
    .A2(\CIC.int_1_out[8] ),
    .A1(net302));
 sg13g2_a21oi_1 _1387_ (.A1(_0657_),
    .A2(net303),
    .Y(_0664_),
    .B1(_0658_));
 sg13g2_xor2_1 _1388_ (.B(net304),
    .A(_0662_),
    .X(_0059_));
 sg13g2_xor2_1 _1389_ (.B(net293),
    .A(net261),
    .X(_0665_));
 sg13g2_a21oi_1 _1390_ (.A1(_0662_),
    .A2(_0664_),
    .Y(_0666_),
    .B1(_0661_));
 sg13g2_xnor2_1 _1391_ (.Y(_0060_),
    .A(_0665_),
    .B(_0666_));
 sg13g2_nand2_1 _1392_ (.Y(_0667_),
    .A(net174),
    .B(net296));
 sg13g2_xnor2_1 _1393_ (.Y(_0668_),
    .A(\CIC.inc_out[12] ),
    .B(\CIC.int_1_out[12] ));
 sg13g2_inv_1 _1394_ (.Y(_0669_),
    .A(_0668_));
 sg13g2_nand2_1 _1395_ (.Y(_0670_),
    .A(_0662_),
    .B(_0665_));
 sg13g2_nor3_1 _1396_ (.A(_0658_),
    .B(_0663_),
    .C(_0670_),
    .Y(_0671_));
 sg13g2_o21ai_1 _1397_ (.B1(_0661_),
    .Y(_0672_),
    .A1(\CIC.inc_out[11] ),
    .A2(\CIC.int_1_out[11] ));
 sg13g2_a21oi_1 _1398_ (.A1(\CIC.inc_out[11] ),
    .A2(\CIC.int_1_out[11] ),
    .Y(_0673_),
    .B1(_0671_));
 sg13g2_nand2_1 _1399_ (.Y(_0674_),
    .A(_0672_),
    .B(_0673_));
 sg13g2_or3_1 _1400_ (.A(_0656_),
    .B(_0659_),
    .C(_0670_),
    .X(_0675_));
 sg13g2_a21oi_2 _1401_ (.B1(_0675_),
    .Y(_0676_),
    .A2(_0653_),
    .A1(_0651_));
 sg13g2_o21ai_1 _1402_ (.B1(_0669_),
    .Y(_0677_),
    .A1(_0674_),
    .A2(_0676_));
 sg13g2_or3_1 _1403_ (.A(_0669_),
    .B(_0674_),
    .C(_0676_),
    .X(_0678_));
 sg13g2_and2_1 _1404_ (.A(_0677_),
    .B(_0678_),
    .X(_0061_));
 sg13g2_nor2_1 _1405_ (.A(net440),
    .B(\CIC.int_1_out[13] ),
    .Y(_0679_));
 sg13g2_xnor2_1 _1406_ (.Y(_0680_),
    .A(net254),
    .B(\CIC.int_1_out[13] ));
 sg13g2_nand2_1 _1407_ (.Y(_0681_),
    .A(_0667_),
    .B(_0677_));
 sg13g2_xnor2_1 _1408_ (.Y(_0062_),
    .A(_0680_),
    .B(_0681_));
 sg13g2_and2_1 _1409_ (.A(net269),
    .B(net305),
    .X(_0682_));
 sg13g2_xor2_1 _1410_ (.B(\CIC.int_1_out[14] ),
    .A(net269),
    .X(_0683_));
 sg13g2_inv_1 _1411_ (.Y(_0684_),
    .A(_0683_));
 sg13g2_a22oi_1 _1412_ (.Y(_0685_),
    .B1(\CIC.int_1_out[13] ),
    .B2(\CIC.inc_out[13] ),
    .A2(\CIC.int_1_out[12] ),
    .A1(\CIC.inc_out[12] ));
 sg13g2_nor2_1 _1413_ (.A(_0679_),
    .B(_0685_),
    .Y(_0686_));
 sg13g2_a21oi_1 _1414_ (.A1(_0677_),
    .A2(_0685_),
    .Y(_0687_),
    .B1(_0679_));
 sg13g2_xnor2_1 _1415_ (.Y(_0063_),
    .A(_0684_),
    .B(_0687_));
 sg13g2_nor2_1 _1416_ (.A(\CIC.inc_out[15] ),
    .B(\CIC.int_1_out[15] ),
    .Y(_0688_));
 sg13g2_xnor2_1 _1417_ (.Y(_0689_),
    .A(\CIC.inc_out[15] ),
    .B(\CIC.int_1_out[15] ));
 sg13g2_a21oi_1 _1418_ (.A1(_0683_),
    .A2(_0687_),
    .Y(_0690_),
    .B1(_0682_));
 sg13g2_xor2_1 _1419_ (.B(net306),
    .A(_0689_),
    .X(_0064_));
 sg13g2_a21oi_1 _1420_ (.A1(\CIC.inc_out[15] ),
    .A2(\CIC.int_1_out[15] ),
    .Y(_0691_),
    .B1(_0682_));
 sg13g2_nor2_1 _1421_ (.A(_0684_),
    .B(_0689_),
    .Y(_0692_));
 sg13g2_nor4_2 _1422_ (.A(_0668_),
    .B(_0680_),
    .C(_0684_),
    .Y(_0693_),
    .D(_0689_));
 sg13g2_a22oi_1 _1423_ (.Y(_0694_),
    .B1(_0693_),
    .B2(_0674_),
    .A2(_0692_),
    .A1(_0686_));
 sg13g2_o21ai_1 _1424_ (.B1(_0694_),
    .Y(_0695_),
    .A1(_0688_),
    .A2(_0691_));
 sg13g2_a21oi_2 _1425_ (.B1(_0695_),
    .Y(_0696_),
    .A2(_0693_),
    .A1(_0676_));
 sg13g2_nand2_1 _1426_ (.Y(_0697_),
    .A(net247),
    .B(net308));
 sg13g2_xor2_1 _1427_ (.B(net308),
    .A(net247),
    .X(_0698_));
 sg13g2_nand2b_1 _1428_ (.Y(_0699_),
    .B(_0698_),
    .A_N(_0696_));
 sg13g2_xnor2_1 _1429_ (.Y(_0065_),
    .A(_0696_),
    .B(_0698_));
 sg13g2_nor2_1 _1430_ (.A(net445),
    .B(\CIC.int_1_out[17] ),
    .Y(_0700_));
 sg13g2_xor2_1 _1431_ (.B(\CIC.int_1_out[17] ),
    .A(net258),
    .X(_0701_));
 sg13g2_nand2_1 _1432_ (.Y(_0702_),
    .A(_0697_),
    .B(_0699_));
 sg13g2_xor2_1 _1433_ (.B(_0702_),
    .A(_0701_),
    .X(_0066_));
 sg13g2_and2_1 _1434_ (.A(net138),
    .B(net289),
    .X(_0703_));
 sg13g2_xor2_1 _1435_ (.B(net448),
    .A(net455),
    .X(_0704_));
 sg13g2_a22oi_1 _1436_ (.Y(_0705_),
    .B1(\CIC.int_1_out[17] ),
    .B2(\CIC.inc_out[17] ),
    .A2(\CIC.int_1_out[16] ),
    .A1(\CIC.inc_out[16] ));
 sg13g2_a21oi_1 _1437_ (.A1(_0699_),
    .A2(_0705_),
    .Y(_0706_),
    .B1(_0700_));
 sg13g2_xor2_1 _1438_ (.B(_0706_),
    .A(net449),
    .X(_0067_));
 sg13g2_nor2_1 _1439_ (.A(\CIC.inc_out[19] ),
    .B(\CIC.int_1_out[19] ),
    .Y(_0707_));
 sg13g2_xor2_1 _1440_ (.B(net415),
    .A(\CIC.inc_out[19] ),
    .X(_0708_));
 sg13g2_a21oi_1 _1441_ (.A1(_0704_),
    .A2(_0706_),
    .Y(_0709_),
    .B1(_0703_));
 sg13g2_xnor2_1 _1442_ (.Y(_0068_),
    .A(net416),
    .B(_0709_));
 sg13g2_nand2_1 _1443_ (.Y(_0710_),
    .A(_0704_),
    .B(_0708_));
 sg13g2_nand4_1 _1444_ (.B(_0701_),
    .C(_0704_),
    .A(_0698_),
    .Y(_0711_),
    .D(_0708_));
 sg13g2_a21oi_1 _1445_ (.A1(\CIC.inc_out[19] ),
    .A2(\CIC.int_1_out[19] ),
    .Y(_0712_),
    .B1(_0703_));
 sg13g2_nor2_1 _1446_ (.A(_0707_),
    .B(_0712_),
    .Y(_0713_));
 sg13g2_nor3_1 _1447_ (.A(_0700_),
    .B(_0705_),
    .C(_0710_),
    .Y(_0714_));
 sg13g2_nor2_1 _1448_ (.A(_0713_),
    .B(_0714_),
    .Y(_0715_));
 sg13g2_o21ai_1 _1449_ (.B1(_0715_),
    .Y(_0716_),
    .A1(_0696_),
    .A2(_0711_));
 sg13g2_and2_1 _1450_ (.A(net287),
    .B(net419),
    .X(_0717_));
 sg13g2_xor2_1 _1451_ (.B(net419),
    .A(net287),
    .X(_0718_));
 sg13g2_xor2_1 _1452_ (.B(_0718_),
    .A(_0716_),
    .X(_0070_));
 sg13g2_xor2_1 _1453_ (.B(net427),
    .A(net256),
    .X(_0719_));
 sg13g2_a21oi_1 _1454_ (.A1(_0716_),
    .A2(_0718_),
    .Y(_0720_),
    .B1(_0717_));
 sg13g2_xnor2_1 _1455_ (.Y(_0071_),
    .A(_0719_),
    .B(_0720_));
 sg13g2_nand2_1 _1456_ (.Y(_0721_),
    .A(net250),
    .B(net446));
 sg13g2_nor2_1 _1457_ (.A(net265),
    .B(\CIC.int_1_out[22] ),
    .Y(_0722_));
 sg13g2_xor2_1 _1458_ (.B(net270),
    .A(net250),
    .X(_0723_));
 sg13g2_and2_1 _1459_ (.A(_0718_),
    .B(_0719_),
    .X(_0724_));
 sg13g2_o21ai_1 _1460_ (.B1(_0717_),
    .Y(_0725_),
    .A1(\CIC.inc_out[21] ),
    .A2(\CIC.int_1_out[21] ));
 sg13g2_inv_1 _1461_ (.Y(_0726_),
    .A(_0725_));
 sg13g2_a221oi_1 _1462_ (.B2(_0724_),
    .C1(_0726_),
    .B1(_0716_),
    .A1(net428),
    .Y(_0727_),
    .A2(\CIC.int_1_out[21] ));
 sg13g2_xnor2_1 _1463_ (.Y(_0072_),
    .A(_0723_),
    .B(net429));
 sg13g2_o21ai_1 _1464_ (.B1(_0721_),
    .Y(_0728_),
    .A1(_0722_),
    .A2(_0727_));
 sg13g2_xnor2_1 _1465_ (.Y(_0729_),
    .A(net72),
    .B(net249));
 sg13g2_xnor2_1 _1466_ (.Y(_0073_),
    .A(net447),
    .B(_0729_));
 sg13g2_xor2_1 _1467_ (.B(net170),
    .A(\CIC.inc_out[0] ),
    .X(_0058_));
 sg13g2_nand2b_2 _1468_ (.Y(_0730_),
    .B(\CIC.dec_clk ),
    .A_N(\CIC.u_differentiator.prev_lr_clk ));
 sg13g2_nor2b_1 _1469_ (.A(net380),
    .B_N(net372),
    .Y(_0731_));
 sg13g2_nand2b_1 _1470_ (.Y(_0732_),
    .B(net372),
    .A_N(net380));
 sg13g2_nor2_1 _1471_ (.A(\CIC.u_differentiator.count[2] ),
    .B(net369),
    .Y(_0733_));
 sg13g2_nand2b_2 _1472_ (.Y(_0734_),
    .B(net370),
    .A_N(\CIC.u_differentiator.count[2] ));
 sg13g2_and2_1 _1473_ (.A(_0730_),
    .B(net360),
    .X(_0735_));
 sg13g2_nor2_1 _1474_ (.A(net119),
    .B(net345),
    .Y(_0736_));
 sg13g2_and2_1 _1475_ (.A(net376),
    .B(net379),
    .X(_0737_));
 sg13g2_nand2_1 _1476_ (.Y(_0738_),
    .A(net372),
    .B(net380));
 sg13g2_nor2_1 _1477_ (.A(net374),
    .B(net380),
    .Y(_0739_));
 sg13g2_or2_1 _1478_ (.X(_0740_),
    .B(net380),
    .A(net372));
 sg13g2_a21oi_1 _1479_ (.A1(net378),
    .A2(\CIC.u_differentiator.a_mux4to1.d1[0] ),
    .Y(_0741_),
    .B1(net376));
 sg13g2_a221oi_1 _1480_ (.B2(_0450_),
    .C1(_0741_),
    .B1(net367),
    .A1(_0451_),
    .Y(_0742_),
    .A2(net370));
 sg13g2_nand2b_1 _1481_ (.Y(_0743_),
    .B(\CIC.u_differentiator.temp[0] ),
    .A_N(_0742_));
 sg13g2_xnor2_1 _1482_ (.Y(_0744_),
    .A(\CIC.u_differentiator.temp[0] ),
    .B(_0742_));
 sg13g2_a21oi_1 _1483_ (.A1(net345),
    .A2(_0744_),
    .Y(_0108_),
    .B1(_0736_));
 sg13g2_nor2_1 _1484_ (.A(net43),
    .B(net345),
    .Y(_0745_));
 sg13g2_xnor2_1 _1485_ (.Y(_0746_),
    .A(net376),
    .B(net378));
 sg13g2_nand2b_1 _1486_ (.Y(_0747_),
    .B(net376),
    .A_N(_0012_));
 sg13g2_nor2b_1 _1487_ (.A(net375),
    .B_N(_0031_),
    .Y(_0748_));
 sg13g2_a221oi_1 _1488_ (.B2(_0449_),
    .C1(_0748_),
    .B1(_0747_),
    .A1(_0011_),
    .Y(_0749_),
    .A2(_0746_));
 sg13g2_nand2b_1 _1489_ (.Y(_0750_),
    .B(_0749_),
    .A_N(\CIC.u_differentiator.temp[1] ));
 sg13g2_inv_1 _1490_ (.Y(_0751_),
    .A(_0750_));
 sg13g2_xnor2_1 _1491_ (.Y(_0752_),
    .A(\CIC.u_differentiator.temp[1] ),
    .B(_0749_));
 sg13g2_and2_1 _1492_ (.A(_0743_),
    .B(_0752_),
    .X(_0753_));
 sg13g2_xnor2_1 _1493_ (.Y(_0754_),
    .A(_0743_),
    .B(_0752_));
 sg13g2_a21oi_1 _1494_ (.A1(net345),
    .A2(_0754_),
    .Y(_0109_),
    .B1(_0745_));
 sg13g2_nor2_1 _1495_ (.A(net110),
    .B(net347),
    .Y(_0755_));
 sg13g2_nor2_1 _1496_ (.A(_0751_),
    .B(_0753_),
    .Y(_0756_));
 sg13g2_nor2_1 _1497_ (.A(\CIC.u_differentiator.a_mux4to1.d3[2] ),
    .B(net365),
    .Y(_0757_));
 sg13g2_a21oi_1 _1498_ (.A1(net378),
    .A2(\CIC.u_differentiator.a_mux4to1.d1[2] ),
    .Y(_0758_),
    .B1(net376));
 sg13g2_nor2_1 _1499_ (.A(\CIC.u_differentiator.a_mux4to1.d2[2] ),
    .B(net369),
    .Y(_0759_));
 sg13g2_nor3_1 _1500_ (.A(_0757_),
    .B(_0758_),
    .C(_0759_),
    .Y(_0760_));
 sg13g2_nor2b_1 _1501_ (.A(\CIC.u_differentiator.temp[2] ),
    .B_N(_0760_),
    .Y(_0761_));
 sg13g2_xnor2_1 _1502_ (.Y(_0762_),
    .A(\CIC.u_differentiator.temp[2] ),
    .B(_0760_));
 sg13g2_o21ai_1 _1503_ (.B1(_0762_),
    .Y(_0763_),
    .A1(_0751_),
    .A2(_0753_));
 sg13g2_xor2_1 _1504_ (.B(_0762_),
    .A(_0756_),
    .X(_0764_));
 sg13g2_a21oi_1 _1505_ (.A1(net347),
    .A2(_0764_),
    .Y(_0110_),
    .B1(_0755_));
 sg13g2_nor2_1 _1506_ (.A(net54),
    .B(net345),
    .Y(_0765_));
 sg13g2_nand2b_1 _1507_ (.Y(_0766_),
    .B(_0763_),
    .A_N(_0761_));
 sg13g2_nand2_1 _1508_ (.Y(_0767_),
    .A(_0013_),
    .B(net367));
 sg13g2_a22oi_1 _1509_ (.Y(_0768_),
    .B1(net370),
    .B2(_0014_),
    .A2(_0032_),
    .A1(_0448_));
 sg13g2_nand3_1 _1510_ (.B(_0767_),
    .C(_0768_),
    .A(net363),
    .Y(_0769_));
 sg13g2_and2_1 _1511_ (.A(\CIC.u_differentiator.temp[3] ),
    .B(_0769_),
    .X(_0770_));
 sg13g2_nor2_1 _1512_ (.A(\CIC.u_differentiator.temp[3] ),
    .B(_0769_),
    .Y(_0771_));
 sg13g2_nor2_1 _1513_ (.A(_0770_),
    .B(_0771_),
    .Y(_0772_));
 sg13g2_xnor2_1 _1514_ (.Y(_0773_),
    .A(_0766_),
    .B(_0772_));
 sg13g2_a21oi_1 _1515_ (.A1(net345),
    .A2(_0773_),
    .Y(_0111_),
    .B1(_0765_));
 sg13g2_nor2_1 _1516_ (.A(net165),
    .B(net344),
    .Y(_0774_));
 sg13g2_a21oi_1 _1517_ (.A1(net378),
    .A2(\CIC.u_differentiator.a_mux4to1.d1[4] ),
    .Y(_0775_),
    .B1(net375));
 sg13g2_a221oi_1 _1518_ (.B2(_0452_),
    .C1(_0775_),
    .B1(net367),
    .A1(_0453_),
    .Y(_0776_),
    .A2(net370));
 sg13g2_nor2b_1 _1519_ (.A(\CIC.u_differentiator.temp[4] ),
    .B_N(_0776_),
    .Y(_0777_));
 sg13g2_xnor2_1 _1520_ (.Y(_0778_),
    .A(\CIC.u_differentiator.temp[4] ),
    .B(_0776_));
 sg13g2_nor2_1 _1521_ (.A(_0761_),
    .B(_0771_),
    .Y(_0779_));
 sg13g2_a21oi_2 _1522_ (.B1(_0770_),
    .Y(_0780_),
    .A2(_0779_),
    .A1(_0763_));
 sg13g2_xnor2_1 _1523_ (.Y(_0781_),
    .A(_0778_),
    .B(_0780_));
 sg13g2_a21oi_1 _1524_ (.A1(net344),
    .A2(_0781_),
    .Y(_0112_),
    .B1(_0774_));
 sg13g2_nand3_1 _1525_ (.B(net378),
    .C(_0015_),
    .A(net375),
    .Y(_0782_));
 sg13g2_nand2b_1 _1526_ (.Y(_0783_),
    .B(_0033_),
    .A_N(net375));
 sg13g2_nand3b_1 _1527_ (.B(_0016_),
    .C(net375),
    .Y(_0784_),
    .A_N(net378));
 sg13g2_and4_1 _1528_ (.A(net363),
    .B(_0782_),
    .C(_0783_),
    .D(_0784_),
    .X(_0785_));
 sg13g2_nand4_1 _1529_ (.B(_0782_),
    .C(_0783_),
    .A(net363),
    .Y(_0786_),
    .D(_0784_));
 sg13g2_xnor2_1 _1530_ (.Y(_0787_),
    .A(\CIC.u_differentiator.temp[5] ),
    .B(_0785_));
 sg13g2_a21oi_1 _1531_ (.A1(_0778_),
    .A2(_0780_),
    .Y(_0788_),
    .B1(_0777_));
 sg13g2_xor2_1 _1532_ (.B(_0788_),
    .A(_0787_),
    .X(_0789_));
 sg13g2_nor2_1 _1533_ (.A(net53),
    .B(net344),
    .Y(_0790_));
 sg13g2_a21oi_1 _1534_ (.A1(net344),
    .A2(_0789_),
    .Y(_0113_),
    .B1(_0790_));
 sg13g2_nor2_1 _1535_ (.A(net122),
    .B(net343),
    .Y(_0791_));
 sg13g2_a21oi_1 _1536_ (.A1(net378),
    .A2(\CIC.u_differentiator.a_mux4to1.d1[6] ),
    .Y(_0792_),
    .B1(net375));
 sg13g2_a221oi_1 _1537_ (.B2(_0454_),
    .C1(_0792_),
    .B1(net367),
    .A1(_0455_),
    .Y(_0793_),
    .A2(net371));
 sg13g2_nand2b_1 _1538_ (.Y(_0794_),
    .B(_0793_),
    .A_N(\CIC.u_differentiator.temp[6] ));
 sg13g2_xnor2_1 _1539_ (.Y(_0795_),
    .A(\CIC.u_differentiator.temp[6] ),
    .B(_0793_));
 sg13g2_nand2_1 _1540_ (.Y(_0796_),
    .A(_0778_),
    .B(_0787_));
 sg13g2_nand2b_1 _1541_ (.Y(_0797_),
    .B(_0780_),
    .A_N(_0796_));
 sg13g2_a21oi_1 _1542_ (.A1(_0464_),
    .A2(_0785_),
    .Y(_0798_),
    .B1(_0777_));
 sg13g2_a21o_1 _1543_ (.A2(_0786_),
    .A1(\CIC.u_differentiator.temp[5] ),
    .B1(_0798_),
    .X(_0799_));
 sg13g2_and2_1 _1544_ (.A(_0797_),
    .B(_0799_),
    .X(_0800_));
 sg13g2_nand2b_1 _1545_ (.Y(_0801_),
    .B(_0795_),
    .A_N(_0800_));
 sg13g2_xor2_1 _1546_ (.B(_0800_),
    .A(_0795_),
    .X(_0802_));
 sg13g2_a21oi_1 _1547_ (.A1(net343),
    .A2(_0802_),
    .Y(_0114_),
    .B1(_0791_));
 sg13g2_nor2_1 _1548_ (.A(net57),
    .B(net343),
    .Y(_0803_));
 sg13g2_a21oi_1 _1549_ (.A1(net378),
    .A2(\CIC.u_differentiator.a_mux4to1.d1[7] ),
    .Y(_0804_),
    .B1(net375));
 sg13g2_a221oi_1 _1550_ (.B2(_0456_),
    .C1(_0804_),
    .B1(net366),
    .A1(_0457_),
    .Y(_0805_),
    .A2(net371));
 sg13g2_inv_1 _1551_ (.Y(_0806_),
    .A(_0805_));
 sg13g2_xnor2_1 _1552_ (.Y(_0807_),
    .A(\CIC.u_differentiator.temp[7] ),
    .B(_0805_));
 sg13g2_nand2_1 _1553_ (.Y(_0808_),
    .A(_0794_),
    .B(_0801_));
 sg13g2_xnor2_1 _1554_ (.Y(_0809_),
    .A(_0807_),
    .B(_0808_));
 sg13g2_a21oi_1 _1555_ (.A1(net343),
    .A2(_0809_),
    .Y(_0115_),
    .B1(_0803_));
 sg13g2_nor2_1 _1556_ (.A(net81),
    .B(net343),
    .Y(_0810_));
 sg13g2_nor2_1 _1557_ (.A(\CIC.u_differentiator.a_mux4to1.d2[8] ),
    .B(net369),
    .Y(_0811_));
 sg13g2_nor2_1 _1558_ (.A(net377),
    .B(\CIC.u_differentiator.a_mux4to1.d1[8] ),
    .Y(_0812_));
 sg13g2_o21ai_1 _1559_ (.B1(net363),
    .Y(_0813_),
    .A1(\CIC.u_differentiator.a_mux4to1.d3[8] ),
    .A2(net365));
 sg13g2_nor3_1 _1560_ (.A(_0811_),
    .B(_0812_),
    .C(_0813_),
    .Y(_0814_));
 sg13g2_nor2b_1 _1561_ (.A(\CIC.u_differentiator.temp[8] ),
    .B_N(_0814_),
    .Y(_0815_));
 sg13g2_xnor2_1 _1562_ (.Y(_0816_),
    .A(\CIC.u_differentiator.temp[8] ),
    .B(_0814_));
 sg13g2_a21oi_1 _1563_ (.A1(\CIC.u_differentiator.temp[7] ),
    .A2(_0806_),
    .Y(_0817_),
    .B1(_0794_));
 sg13g2_a21oi_1 _1564_ (.A1(_0465_),
    .A2(_0805_),
    .Y(_0818_),
    .B1(_0817_));
 sg13g2_nand2_1 _1565_ (.Y(_0819_),
    .A(_0795_),
    .B(_0807_));
 sg13g2_or2_1 _1566_ (.X(_0820_),
    .B(_0819_),
    .A(_0796_));
 sg13g2_a221oi_1 _1567_ (.B2(_0763_),
    .C1(_0820_),
    .B1(_0779_),
    .A1(\CIC.u_differentiator.temp[3] ),
    .Y(_0821_),
    .A2(_0769_));
 sg13g2_o21ai_1 _1568_ (.B1(_0818_),
    .Y(_0822_),
    .A1(_0799_),
    .A2(_0819_));
 sg13g2_nor2_2 _1569_ (.A(_0821_),
    .B(_0822_),
    .Y(_0823_));
 sg13g2_o21ai_1 _1570_ (.B1(_0816_),
    .Y(_0824_),
    .A1(_0821_),
    .A2(_0822_));
 sg13g2_xor2_1 _1571_ (.B(_0823_),
    .A(_0816_),
    .X(_0825_));
 sg13g2_a21oi_1 _1572_ (.A1(net343),
    .A2(_0825_),
    .Y(_0116_),
    .B1(_0810_));
 sg13g2_a21oi_1 _1573_ (.A1(net379),
    .A2(_0466_),
    .Y(_0826_),
    .B1(net377));
 sg13g2_a221oi_1 _1574_ (.B2(_0019_),
    .C1(_0826_),
    .B1(net366),
    .A1(_0020_),
    .Y(_0827_),
    .A2(net371));
 sg13g2_nand2b_1 _1575_ (.Y(_0828_),
    .B(\CIC.u_differentiator.temp[9] ),
    .A_N(_0827_));
 sg13g2_nor2b_1 _1576_ (.A(\CIC.u_differentiator.temp[9] ),
    .B_N(_0827_),
    .Y(_0829_));
 sg13g2_xnor2_1 _1577_ (.Y(_0830_),
    .A(\CIC.u_differentiator.temp[9] ),
    .B(_0827_));
 sg13g2_nand2b_1 _1578_ (.Y(_0831_),
    .B(_0824_),
    .A_N(_0815_));
 sg13g2_xnor2_1 _1579_ (.Y(_0832_),
    .A(_0830_),
    .B(_0831_));
 sg13g2_nor2_1 _1580_ (.A(net41),
    .B(net343),
    .Y(_0833_));
 sg13g2_a21oi_1 _1581_ (.A1(net343),
    .A2(_0832_),
    .Y(_0117_),
    .B1(_0833_));
 sg13g2_nor2_1 _1582_ (.A(net92),
    .B(net346),
    .Y(_0834_));
 sg13g2_nor2_1 _1583_ (.A(\CIC.u_differentiator.a_mux4to1.d2[10] ),
    .B(net369),
    .Y(_0835_));
 sg13g2_nor2_1 _1584_ (.A(net377),
    .B(\CIC.u_differentiator.a_mux4to1.d1[10] ),
    .Y(_0836_));
 sg13g2_o21ai_1 _1585_ (.B1(net363),
    .Y(_0837_),
    .A1(\CIC.u_differentiator.a_mux4to1.d3[10] ),
    .A2(net365));
 sg13g2_nor3_1 _1586_ (.A(_0835_),
    .B(_0836_),
    .C(_0837_),
    .Y(_0838_));
 sg13g2_nor2b_1 _1587_ (.A(\CIC.u_differentiator.temp[10] ),
    .B_N(_0838_),
    .Y(_0839_));
 sg13g2_xnor2_1 _1588_ (.Y(_0840_),
    .A(\CIC.u_differentiator.temp[10] ),
    .B(_0838_));
 sg13g2_nand2_1 _1589_ (.Y(_0841_),
    .A(_0816_),
    .B(_0830_));
 sg13g2_a21oi_1 _1590_ (.A1(_0815_),
    .A2(_0828_),
    .Y(_0842_),
    .B1(_0829_));
 sg13g2_inv_1 _1591_ (.Y(_0843_),
    .A(_0842_));
 sg13g2_o21ai_1 _1592_ (.B1(_0842_),
    .Y(_0844_),
    .A1(_0823_),
    .A2(_0841_));
 sg13g2_xnor2_1 _1593_ (.Y(_0845_),
    .A(_0840_),
    .B(_0844_));
 sg13g2_a21oi_1 _1594_ (.A1(net346),
    .A2(_0845_),
    .Y(_0118_),
    .B1(_0834_));
 sg13g2_nor2_1 _1595_ (.A(net105),
    .B(net341),
    .Y(_0846_));
 sg13g2_nor2_1 _1596_ (.A(\CIC.u_differentiator.a_mux4to1.d2[11] ),
    .B(net368),
    .Y(_0847_));
 sg13g2_nor2_1 _1597_ (.A(net374),
    .B(\CIC.u_differentiator.a_mux4to1.d1[11] ),
    .Y(_0848_));
 sg13g2_o21ai_1 _1598_ (.B1(net362),
    .Y(_0849_),
    .A1(\CIC.u_differentiator.a_mux4to1.d3[11] ),
    .A2(net365));
 sg13g2_nor3_2 _1599_ (.A(_0847_),
    .B(_0848_),
    .C(_0849_),
    .Y(_0850_));
 sg13g2_nor2_1 _1600_ (.A(_0467_),
    .B(_0850_),
    .Y(_0851_));
 sg13g2_xnor2_1 _1601_ (.Y(_0852_),
    .A(\CIC.u_differentiator.temp[11] ),
    .B(_0850_));
 sg13g2_a21oi_1 _1602_ (.A1(_0840_),
    .A2(_0844_),
    .Y(_0853_),
    .B1(_0839_));
 sg13g2_xor2_1 _1603_ (.B(_0853_),
    .A(_0852_),
    .X(_0854_));
 sg13g2_a21oi_1 _1604_ (.A1(net341),
    .A2(_0854_),
    .Y(_0119_),
    .B1(_0846_));
 sg13g2_nor2_1 _1605_ (.A(net86),
    .B(net346),
    .Y(_0855_));
 sg13g2_a21oi_1 _1606_ (.A1(net379),
    .A2(\CIC.u_differentiator.a_mux4to1.d1[12] ),
    .Y(_0856_),
    .B1(net377));
 sg13g2_a221oi_1 _1607_ (.B2(_0458_),
    .C1(_0856_),
    .B1(net366),
    .A1(_0459_),
    .Y(_0857_),
    .A2(net371));
 sg13g2_nor2b_1 _1608_ (.A(\CIC.u_differentiator.temp[12] ),
    .B_N(_0857_),
    .Y(_0858_));
 sg13g2_xnor2_1 _1609_ (.Y(_0859_),
    .A(\CIC.u_differentiator.temp[12] ),
    .B(_0857_));
 sg13g2_nand2_1 _1610_ (.Y(_0860_),
    .A(_0840_),
    .B(_0852_));
 sg13g2_inv_1 _1611_ (.Y(_0861_),
    .A(_0860_));
 sg13g2_a21oi_1 _1612_ (.A1(_0467_),
    .A2(_0850_),
    .Y(_0862_),
    .B1(_0839_));
 sg13g2_nor2_1 _1613_ (.A(_0851_),
    .B(_0862_),
    .Y(_0863_));
 sg13g2_a21oi_2 _1614_ (.B1(_0863_),
    .Y(_0864_),
    .A2(_0861_),
    .A1(_0844_));
 sg13g2_nor2b_1 _1615_ (.A(_0864_),
    .B_N(_0859_),
    .Y(_0865_));
 sg13g2_xor2_1 _1616_ (.B(_0864_),
    .A(_0859_),
    .X(_0866_));
 sg13g2_a21oi_1 _1617_ (.A1(net346),
    .A2(_0866_),
    .Y(_0120_),
    .B1(_0855_));
 sg13g2_nand2_1 _1618_ (.Y(_0867_),
    .A(_0023_),
    .B(net366));
 sg13g2_nand2b_1 _1619_ (.Y(_0868_),
    .B(_0007_),
    .A_N(net374));
 sg13g2_nand2_1 _1620_ (.Y(_0869_),
    .A(_0024_),
    .B(net370));
 sg13g2_and4_1 _1621_ (.A(net363),
    .B(_0867_),
    .C(_0868_),
    .D(_0869_),
    .X(_0870_));
 sg13g2_nand4_1 _1622_ (.B(_0867_),
    .C(_0868_),
    .A(net362),
    .Y(_0871_),
    .D(_0869_));
 sg13g2_xnor2_1 _1623_ (.Y(_0872_),
    .A(\CIC.u_differentiator.temp[13] ),
    .B(_0870_));
 sg13g2_nor2_1 _1624_ (.A(_0858_),
    .B(_0865_),
    .Y(_0873_));
 sg13g2_xor2_1 _1625_ (.B(_0873_),
    .A(_0872_),
    .X(_0874_));
 sg13g2_nor2_1 _1626_ (.A(net42),
    .B(net346),
    .Y(_0875_));
 sg13g2_a21oi_1 _1627_ (.A1(net346),
    .A2(_0874_),
    .Y(_0121_),
    .B1(_0875_));
 sg13g2_nor2_1 _1628_ (.A(net142),
    .B(net341),
    .Y(_0876_));
 sg13g2_nor2_1 _1629_ (.A(\CIC.u_differentiator.a_mux4to1.d2[14] ),
    .B(net368),
    .Y(_0877_));
 sg13g2_nor2_1 _1630_ (.A(net374),
    .B(\CIC.u_differentiator.a_mux4to1.d1[14] ),
    .Y(_0878_));
 sg13g2_o21ai_1 _1631_ (.B1(net363),
    .Y(_0879_),
    .A1(\CIC.u_differentiator.a_mux4to1.d3[14] ),
    .A2(net364));
 sg13g2_nor3_2 _1632_ (.A(_0877_),
    .B(_0878_),
    .C(_0879_),
    .Y(_0880_));
 sg13g2_and2_1 _1633_ (.A(_0469_),
    .B(_0880_),
    .X(_0881_));
 sg13g2_nand2_1 _1634_ (.Y(_0882_),
    .A(_0469_),
    .B(_0880_));
 sg13g2_xnor2_1 _1635_ (.Y(_0883_),
    .A(\CIC.u_differentiator.temp[14] ),
    .B(_0880_));
 sg13g2_nand2_1 _1636_ (.Y(_0884_),
    .A(_0859_),
    .B(_0872_));
 sg13g2_a21oi_1 _1637_ (.A1(_0468_),
    .A2(_0870_),
    .Y(_0885_),
    .B1(_0858_));
 sg13g2_a21o_1 _1638_ (.A2(_0871_),
    .A1(\CIC.u_differentiator.temp[13] ),
    .B1(_0885_),
    .X(_0886_));
 sg13g2_o21ai_1 _1639_ (.B1(_0886_),
    .Y(_0887_),
    .A1(_0864_),
    .A2(_0884_));
 sg13g2_xnor2_1 _1640_ (.Y(_0888_),
    .A(_0883_),
    .B(_0887_));
 sg13g2_a21oi_1 _1641_ (.A1(net341),
    .A2(_0888_),
    .Y(_0122_),
    .B1(_0876_));
 sg13g2_nor2_1 _1642_ (.A(net48),
    .B(net341),
    .Y(_0889_));
 sg13g2_a21oi_1 _1643_ (.A1(net380),
    .A2(_0470_),
    .Y(_0890_),
    .B1(net374));
 sg13g2_a221oi_1 _1644_ (.B2(_0025_),
    .C1(_0890_),
    .B1(net366),
    .A1(_0026_),
    .Y(_0891_),
    .A2(net370));
 sg13g2_nand2_1 _1645_ (.Y(_0892_),
    .A(_0471_),
    .B(_0891_));
 sg13g2_nor2_1 _1646_ (.A(_0471_),
    .B(_0891_),
    .Y(_0893_));
 sg13g2_xnor2_1 _1647_ (.Y(_0894_),
    .A(\CIC.u_differentiator.temp[15] ),
    .B(_0891_));
 sg13g2_a21oi_1 _1648_ (.A1(_0883_),
    .A2(_0887_),
    .Y(_0895_),
    .B1(_0881_));
 sg13g2_xor2_1 _1649_ (.B(_0895_),
    .A(_0894_),
    .X(_0896_));
 sg13g2_a21oi_1 _1650_ (.A1(net341),
    .A2(_0896_),
    .Y(_0123_),
    .B1(_0889_));
 sg13g2_nor2_1 _1651_ (.A(net97),
    .B(net342),
    .Y(_0897_));
 sg13g2_nand2_1 _1652_ (.Y(_0898_),
    .A(_0883_),
    .B(_0894_));
 sg13g2_nor2_1 _1653_ (.A(_0884_),
    .B(_0898_),
    .Y(_0899_));
 sg13g2_nor3_1 _1654_ (.A(_0860_),
    .B(_0884_),
    .C(_0898_),
    .Y(_0900_));
 sg13g2_nand2b_1 _1655_ (.Y(_0901_),
    .B(_0900_),
    .A_N(_0841_));
 sg13g2_a21o_1 _1656_ (.A2(_0892_),
    .A1(_0882_),
    .B1(_0893_),
    .X(_0902_));
 sg13g2_o21ai_1 _1657_ (.B1(_0902_),
    .Y(_0903_),
    .A1(_0886_),
    .A2(_0898_));
 sg13g2_a221oi_1 _1658_ (.B2(_0843_),
    .C1(_0903_),
    .B1(_0900_),
    .A1(_0863_),
    .Y(_0904_),
    .A2(_0899_));
 sg13g2_o21ai_1 _1659_ (.B1(_0904_),
    .Y(_0905_),
    .A1(_0823_),
    .A2(_0901_));
 sg13g2_nor2_1 _1660_ (.A(\CIC.u_differentiator.a_mux4to1.d2[16] ),
    .B(net368),
    .Y(_0906_));
 sg13g2_nor2_1 _1661_ (.A(net373),
    .B(\CIC.u_differentiator.a_mux4to1.d1[16] ),
    .Y(_0907_));
 sg13g2_o21ai_1 _1662_ (.B1(net362),
    .Y(_0908_),
    .A1(\CIC.u_differentiator.a_mux4to1.d3[16] ),
    .A2(net365));
 sg13g2_nor3_1 _1663_ (.A(_0906_),
    .B(_0907_),
    .C(_0908_),
    .Y(_0231_));
 sg13g2_nor2b_1 _1664_ (.A(\CIC.u_differentiator.temp[16] ),
    .B_N(_0231_),
    .Y(_0232_));
 sg13g2_xnor2_1 _1665_ (.Y(_0233_),
    .A(\CIC.u_differentiator.temp[16] ),
    .B(_0231_));
 sg13g2_xnor2_1 _1666_ (.Y(_0234_),
    .A(_0905_),
    .B(_0233_));
 sg13g2_a21oi_1 _1667_ (.A1(net341),
    .A2(_0234_),
    .Y(_0124_),
    .B1(_0897_));
 sg13g2_nor2_1 _1668_ (.A(net156),
    .B(net341),
    .Y(_0235_));
 sg13g2_nor2_1 _1669_ (.A(\CIC.u_differentiator.a_mux4to1.d2[17] ),
    .B(net368),
    .Y(_0236_));
 sg13g2_nor2_1 _1670_ (.A(net372),
    .B(\CIC.u_differentiator.a_mux4to1.d1[17] ),
    .Y(_0237_));
 sg13g2_o21ai_1 _1671_ (.B1(net362),
    .Y(_0238_),
    .A1(\CIC.u_differentiator.a_mux4to1.d3[17] ),
    .A2(net364));
 sg13g2_nor3_1 _1672_ (.A(_0236_),
    .B(_0237_),
    .C(_0238_),
    .Y(_0239_));
 sg13g2_nand2b_1 _1673_ (.Y(_0240_),
    .B(\CIC.u_differentiator.temp[17] ),
    .A_N(_0239_));
 sg13g2_inv_1 _1674_ (.Y(_0241_),
    .A(_0240_));
 sg13g2_nor2b_1 _1675_ (.A(\CIC.u_differentiator.temp[17] ),
    .B_N(_0239_),
    .Y(_0242_));
 sg13g2_nor2_1 _1676_ (.A(_0241_),
    .B(_0242_),
    .Y(_0243_));
 sg13g2_a21oi_1 _1677_ (.A1(_0905_),
    .A2(_0233_),
    .Y(_0244_),
    .B1(_0232_));
 sg13g2_xor2_1 _1678_ (.B(_0244_),
    .A(_0243_),
    .X(_0245_));
 sg13g2_a21oi_1 _1679_ (.A1(net339),
    .A2(_0245_),
    .Y(_0125_),
    .B1(_0235_));
 sg13g2_nor2_1 _1680_ (.A(net80),
    .B(net339),
    .Y(_0246_));
 sg13g2_nor2_1 _1681_ (.A(\CIC.u_differentiator.a_mux4to1.d2[18] ),
    .B(net368),
    .Y(_0247_));
 sg13g2_nor2_1 _1682_ (.A(net372),
    .B(\CIC.u_differentiator.a_mux4to1.d1[18] ),
    .Y(_0248_));
 sg13g2_o21ai_1 _1683_ (.B1(net362),
    .Y(_0249_),
    .A1(\CIC.u_differentiator.a_mux4to1.d3[18] ),
    .A2(net364));
 sg13g2_nor3_1 _1684_ (.A(_0247_),
    .B(_0248_),
    .C(_0249_),
    .Y(_0250_));
 sg13g2_nor2b_1 _1685_ (.A(\CIC.u_differentiator.temp[18] ),
    .B_N(_0250_),
    .Y(_0251_));
 sg13g2_xnor2_1 _1686_ (.Y(_0252_),
    .A(\CIC.u_differentiator.temp[18] ),
    .B(_0250_));
 sg13g2_a21oi_1 _1687_ (.A1(_0232_),
    .A2(_0240_),
    .Y(_0253_),
    .B1(_0242_));
 sg13g2_and2_1 _1688_ (.A(_0233_),
    .B(_0243_),
    .X(_0254_));
 sg13g2_a221oi_1 _1689_ (.B2(_0905_),
    .C1(_0242_),
    .B1(_0254_),
    .A1(_0232_),
    .Y(_0255_),
    .A2(_0240_));
 sg13g2_nor2b_1 _1690_ (.A(_0255_),
    .B_N(_0252_),
    .Y(_0256_));
 sg13g2_xor2_1 _1691_ (.B(_0255_),
    .A(_0252_),
    .X(_0257_));
 sg13g2_a21oi_1 _1692_ (.A1(net339),
    .A2(_0257_),
    .Y(_0126_),
    .B1(_0246_));
 sg13g2_nor2_1 _1693_ (.A(net98),
    .B(net339),
    .Y(_0258_));
 sg13g2_or2_1 _1694_ (.X(_0259_),
    .B(\CIC.u_differentiator.a_mux4to1.d1[19] ),
    .A(net372));
 sg13g2_o21ai_1 _1695_ (.B1(net362),
    .Y(_0260_),
    .A1(\CIC.u_differentiator.a_mux4to1.d3[19] ),
    .A2(net364));
 sg13g2_o21ai_1 _1696_ (.B1(_0259_),
    .Y(_0261_),
    .A1(\CIC.u_differentiator.a_mux4to1.d2[19] ),
    .A2(net368));
 sg13g2_o21ai_1 _1697_ (.B1(\CIC.u_differentiator.temp[19] ),
    .Y(_0262_),
    .A1(_0260_),
    .A2(_0261_));
 sg13g2_or3_1 _1698_ (.A(\CIC.u_differentiator.temp[19] ),
    .B(_0260_),
    .C(_0261_),
    .X(_0263_));
 sg13g2_and2_1 _1699_ (.A(_0262_),
    .B(_0263_),
    .X(_0264_));
 sg13g2_nor2_1 _1700_ (.A(_0251_),
    .B(_0256_),
    .Y(_0265_));
 sg13g2_xor2_1 _1701_ (.B(_0265_),
    .A(_0264_),
    .X(_0266_));
 sg13g2_a21oi_1 _1702_ (.A1(net339),
    .A2(_0266_),
    .Y(_0127_),
    .B1(_0258_));
 sg13g2_nor2_1 _1703_ (.A(net99),
    .B(net340),
    .Y(_0267_));
 sg13g2_nand2_1 _1704_ (.Y(_0268_),
    .A(_0252_),
    .B(_0264_));
 sg13g2_and3_1 _1705_ (.X(_0269_),
    .A(_0252_),
    .B(_0254_),
    .C(_0264_));
 sg13g2_o21ai_1 _1706_ (.B1(_0263_),
    .Y(_0270_),
    .A1(_0253_),
    .A2(_0268_));
 sg13g2_a221oi_1 _1707_ (.B2(_0905_),
    .C1(_0270_),
    .B1(_0269_),
    .A1(_0251_),
    .Y(_0271_),
    .A2(_0262_));
 sg13g2_a21oi_1 _1708_ (.A1(net380),
    .A2(\CIC.u_differentiator.a_mux4to1.d1[20] ),
    .Y(_0272_),
    .B1(net373));
 sg13g2_a21oi_1 _1709_ (.A1(_0460_),
    .A2(net370),
    .Y(_0273_),
    .B1(_0272_));
 sg13g2_o21ai_1 _1710_ (.B1(_0273_),
    .Y(_0274_),
    .A1(\CIC.u_differentiator.a_mux4to1.d3[20] ),
    .A2(net364));
 sg13g2_xor2_1 _1711_ (.B(_0274_),
    .A(\CIC.u_differentiator.temp[20] ),
    .X(_0275_));
 sg13g2_nand2b_1 _1712_ (.Y(_0276_),
    .B(_0275_),
    .A_N(_0271_));
 sg13g2_xor2_1 _1713_ (.B(_0275_),
    .A(_0271_),
    .X(_0277_));
 sg13g2_a21oi_1 _1714_ (.A1(net339),
    .A2(_0277_),
    .Y(_0128_),
    .B1(_0267_));
 sg13g2_nor2_1 _1715_ (.A(net112),
    .B(net340),
    .Y(_0278_));
 sg13g2_nor2_1 _1716_ (.A(\CIC.u_differentiator.a_mux4to1.d2[21] ),
    .B(net368),
    .Y(_0279_));
 sg13g2_nor2_1 _1717_ (.A(net373),
    .B(\CIC.u_differentiator.a_mux4to1.d1[21] ),
    .Y(_0280_));
 sg13g2_o21ai_1 _1718_ (.B1(net362),
    .Y(_0281_),
    .A1(\CIC.u_differentiator.a_mux4to1.d3[21] ),
    .A2(net364));
 sg13g2_nor3_2 _1719_ (.A(_0279_),
    .B(_0280_),
    .C(_0281_),
    .Y(_0282_));
 sg13g2_nor2_1 _1720_ (.A(_0472_),
    .B(_0282_),
    .Y(_0283_));
 sg13g2_xnor2_1 _1721_ (.Y(_0284_),
    .A(\CIC.u_differentiator.temp[21] ),
    .B(_0282_));
 sg13g2_o21ai_1 _1722_ (.B1(_0276_),
    .Y(_0285_),
    .A1(\CIC.u_differentiator.temp[20] ),
    .A2(_0274_));
 sg13g2_xnor2_1 _1723_ (.Y(_0286_),
    .A(_0284_),
    .B(_0285_));
 sg13g2_a21oi_1 _1724_ (.A1(net340),
    .A2(_0286_),
    .Y(_0129_),
    .B1(_0278_));
 sg13g2_nor2_1 _1725_ (.A(net101),
    .B(net339),
    .Y(_0287_));
 sg13g2_nand2_1 _1726_ (.Y(_0288_),
    .A(_0275_),
    .B(_0284_));
 sg13g2_nor3_1 _1727_ (.A(\CIC.u_differentiator.temp[20] ),
    .B(_0274_),
    .C(_0283_),
    .Y(_0289_));
 sg13g2_a21oi_1 _1728_ (.A1(_0472_),
    .A2(_0282_),
    .Y(_0290_),
    .B1(_0289_));
 sg13g2_o21ai_1 _1729_ (.B1(_0290_),
    .Y(_0291_),
    .A1(_0271_),
    .A2(_0288_));
 sg13g2_a21oi_1 _1730_ (.A1(net380),
    .A2(\CIC.u_differentiator.a_mux4to1.d1[22] ),
    .Y(_0292_),
    .B1(net373));
 sg13g2_a21oi_1 _1731_ (.A1(_0461_),
    .A2(net370),
    .Y(_0293_),
    .B1(_0292_));
 sg13g2_o21ai_1 _1732_ (.B1(_0293_),
    .Y(_0294_),
    .A1(\CIC.u_differentiator.a_mux4to1.d3[22] ),
    .A2(net364));
 sg13g2_nor2_1 _1733_ (.A(\CIC.u_differentiator.temp[22] ),
    .B(_0294_),
    .Y(_0295_));
 sg13g2_xor2_1 _1734_ (.B(_0294_),
    .A(\CIC.u_differentiator.temp[22] ),
    .X(_0296_));
 sg13g2_xnor2_1 _1735_ (.Y(_0297_),
    .A(_0291_),
    .B(_0296_));
 sg13g2_a21oi_1 _1736_ (.A1(net339),
    .A2(_0297_),
    .Y(_0130_),
    .B1(_0287_));
 sg13g2_nor2_1 _1737_ (.A(net127),
    .B(net340),
    .Y(_0298_));
 sg13g2_a21oi_1 _1738_ (.A1(_0291_),
    .A2(_0296_),
    .Y(_0299_),
    .B1(_0295_));
 sg13g2_nor2_1 _1739_ (.A(\CIC.u_differentiator.a_mux4to1.d2[23] ),
    .B(net368),
    .Y(_0300_));
 sg13g2_nor2_1 _1740_ (.A(net372),
    .B(\CIC.u_differentiator.a_mux4to1.d1[23] ),
    .Y(_0301_));
 sg13g2_o21ai_1 _1741_ (.B1(net362),
    .Y(_0302_),
    .A1(\CIC.u_differentiator.a_mux4to1.d3[23] ),
    .A2(net364));
 sg13g2_nor3_1 _1742_ (.A(_0300_),
    .B(_0301_),
    .C(_0302_),
    .Y(_0303_));
 sg13g2_xor2_1 _1743_ (.B(_0303_),
    .A(\CIC.u_differentiator.temp[23] ),
    .X(_0304_));
 sg13g2_xnor2_1 _1744_ (.Y(_0305_),
    .A(_0299_),
    .B(_0304_));
 sg13g2_a21oi_1 _1745_ (.A1(net340),
    .A2(_0305_),
    .Y(_0131_),
    .B1(_0298_));
 sg13g2_nand2_1 _1746_ (.Y(_0306_),
    .A(net182),
    .B(_0739_));
 sg13g2_nand3_1 _1747_ (.B(_0730_),
    .C(_0739_),
    .A(_0009_),
    .Y(_0307_));
 sg13g2_nor3_1 _1748_ (.A(net377),
    .B(_0449_),
    .C(\CIC.u_differentiator.count[2] ),
    .Y(_0308_));
 sg13g2_and2_1 _1749_ (.A(_0730_),
    .B(net356),
    .X(_0309_));
 sg13g2_or2_1 _1750_ (.X(_0310_),
    .B(net332),
    .A(net346));
 sg13g2_nor2b_1 _1751_ (.A(_0310_),
    .B_N(net336),
    .Y(_0311_));
 sg13g2_nor2_1 _1752_ (.A(net360),
    .B(net355),
    .Y(_0312_));
 sg13g2_nand2_1 _1753_ (.Y(_0313_),
    .A(net136),
    .B(net358));
 sg13g2_a22oi_1 _1754_ (.Y(_0314_),
    .B1(net353),
    .B2(\CIC.u_differentiator.a_mux4to1.d1[0] ),
    .A2(net361),
    .A1(net119));
 sg13g2_a21oi_1 _1755_ (.A1(_0313_),
    .A2(_0314_),
    .Y(_0315_),
    .B1(net314));
 sg13g2_a21o_1 _1756_ (.A2(net314),
    .A1(net176),
    .B1(_0315_),
    .X(_0132_));
 sg13g2_nand2b_1 _1757_ (.Y(_0316_),
    .B(net357),
    .A_N(_0012_));
 sg13g2_o21ai_1 _1758_ (.B1(_0316_),
    .Y(_0317_),
    .A1(_0011_),
    .A2(_0734_));
 sg13g2_a21oi_1 _1759_ (.A1(\CIC.u_differentiator.a_mux4to1.d1[1] ),
    .A2(net352),
    .Y(_0318_),
    .B1(_0317_));
 sg13g2_nand2_1 _1760_ (.Y(_0319_),
    .A(net103),
    .B(net314));
 sg13g2_o21ai_1 _1761_ (.B1(_0319_),
    .Y(_0133_),
    .A1(net314),
    .A2(_0318_));
 sg13g2_nand2_1 _1762_ (.Y(_0320_),
    .A(\CIC.u_differentiator.a_mux4to1.d1[2] ),
    .B(net352));
 sg13g2_a22oi_1 _1763_ (.Y(_0321_),
    .B1(net357),
    .B2(\CIC.u_differentiator.a_mux4to1.d2[2] ),
    .A2(net361),
    .A1(net110));
 sg13g2_a21oi_1 _1764_ (.A1(_0320_),
    .A2(_0321_),
    .Y(_0322_),
    .B1(net314));
 sg13g2_a21o_1 _1765_ (.A2(net314),
    .A1(net195),
    .B1(_0322_),
    .X(_0134_));
 sg13g2_nand2b_1 _1766_ (.Y(_0323_),
    .B(net357),
    .A_N(_0014_));
 sg13g2_o21ai_1 _1767_ (.B1(_0323_),
    .Y(_0324_),
    .A1(_0013_),
    .A2(_0734_));
 sg13g2_a21oi_1 _1768_ (.A1(net154),
    .A2(net352),
    .Y(_0325_),
    .B1(_0324_));
 sg13g2_nand2_1 _1769_ (.Y(_0326_),
    .A(net162),
    .B(net314));
 sg13g2_o21ai_1 _1770_ (.B1(_0326_),
    .Y(_0135_),
    .A1(net314),
    .A2(_0325_));
 sg13g2_nand2_1 _1771_ (.Y(_0327_),
    .A(net109),
    .B(net357));
 sg13g2_a22oi_1 _1772_ (.Y(_0328_),
    .B1(net352),
    .B2(\CIC.u_differentiator.a_mux4to1.d1[4] ),
    .A2(net361),
    .A1(net165));
 sg13g2_a21oi_1 _1773_ (.A1(_0327_),
    .A2(_0328_),
    .Y(_0329_),
    .B1(net313));
 sg13g2_a21o_1 _1774_ (.A2(net313),
    .A1(net191),
    .B1(_0329_),
    .X(_0136_));
 sg13g2_nand2_1 _1775_ (.Y(_0330_),
    .A(net123),
    .B(net353));
 sg13g2_nor2b_1 _1776_ (.A(_0016_),
    .B_N(net357),
    .Y(_0331_));
 sg13g2_o21ai_1 _1777_ (.B1(_0330_),
    .Y(_0332_),
    .A1(_0015_),
    .A2(net359));
 sg13g2_nor3_1 _1778_ (.A(net313),
    .B(_0331_),
    .C(_0332_),
    .Y(_0333_));
 sg13g2_a21oi_1 _1779_ (.A1(_0464_),
    .A2(net313),
    .Y(_0137_),
    .B1(_0333_));
 sg13g2_nand2_1 _1780_ (.Y(_0334_),
    .A(\CIC.u_differentiator.a_mux4to1.d1[6] ),
    .B(net353));
 sg13g2_a22oi_1 _1781_ (.Y(_0335_),
    .B1(net357),
    .B2(net78),
    .A2(net361),
    .A1(net122));
 sg13g2_a21oi_1 _1782_ (.A1(_0334_),
    .A2(_0335_),
    .Y(_0336_),
    .B1(net313));
 sg13g2_a21o_1 _1783_ (.A2(net313),
    .A1(net189),
    .B1(_0336_),
    .X(_0138_));
 sg13g2_nand2_1 _1784_ (.Y(_0337_),
    .A(\CIC.u_differentiator.a_mux4to1.d1[7] ),
    .B(net353));
 sg13g2_nor2b_1 _1785_ (.A(net147),
    .B_N(net357),
    .Y(_0338_));
 sg13g2_o21ai_1 _1786_ (.B1(_0337_),
    .Y(_0339_),
    .A1(_0017_),
    .A2(net359));
 sg13g2_nor3_1 _1787_ (.A(net313),
    .B(_0338_),
    .C(_0339_),
    .Y(_0340_));
 sg13g2_a21oi_1 _1788_ (.A1(_0465_),
    .A2(net313),
    .Y(_0139_),
    .B1(net148));
 sg13g2_nand2_1 _1789_ (.Y(_0341_),
    .A(\CIC.u_differentiator.a_mux4to1.d1[8] ),
    .B(net352));
 sg13g2_a22oi_1 _1790_ (.Y(_0342_),
    .B1(net357),
    .B2(net106),
    .A2(net361),
    .A1(net81));
 sg13g2_a21oi_1 _1791_ (.A1(_0341_),
    .A2(_0342_),
    .Y(_0343_),
    .B1(net312));
 sg13g2_a21o_1 _1792_ (.A2(net312),
    .A1(net202),
    .B1(_0343_),
    .X(_0140_));
 sg13g2_nand2b_1 _1793_ (.Y(_0344_),
    .B(net358),
    .A_N(_0020_));
 sg13g2_o21ai_1 _1794_ (.B1(_0344_),
    .Y(_0345_),
    .A1(_0019_),
    .A2(net359));
 sg13g2_a21oi_1 _1795_ (.A1(\CIC.u_differentiator.a_mux4to1.d1[9] ),
    .A2(net352),
    .Y(_0346_),
    .B1(_0345_));
 sg13g2_nand2_1 _1796_ (.Y(_0347_),
    .A(net145),
    .B(net312));
 sg13g2_o21ai_1 _1797_ (.B1(_0347_),
    .Y(_0141_),
    .A1(net312),
    .A2(_0346_));
 sg13g2_nand2_1 _1798_ (.Y(_0348_),
    .A(\CIC.u_differentiator.a_mux4to1.d1[10] ),
    .B(net352));
 sg13g2_a22oi_1 _1799_ (.Y(_0349_),
    .B1(net358),
    .B2(net135),
    .A2(_0733_),
    .A1(net92));
 sg13g2_a21oi_1 _1800_ (.A1(_0348_),
    .A2(_0349_),
    .Y(_0350_),
    .B1(net312));
 sg13g2_a21o_1 _1801_ (.A2(net312),
    .A1(net193),
    .B1(_0350_),
    .X(_0142_));
 sg13g2_nand2_1 _1802_ (.Y(_0351_),
    .A(\CIC.u_differentiator.a_mux4to1.d1[11] ),
    .B(net351));
 sg13g2_nor2b_1 _1803_ (.A(net131),
    .B_N(net356),
    .Y(_0352_));
 sg13g2_o21ai_1 _1804_ (.B1(_0351_),
    .Y(_0353_),
    .A1(_0021_),
    .A2(net359));
 sg13g2_nor3_1 _1805_ (.A(net311),
    .B(_0352_),
    .C(_0353_),
    .Y(_0354_));
 sg13g2_a21oi_1 _1806_ (.A1(_0467_),
    .A2(net311),
    .Y(_0143_),
    .B1(net132));
 sg13g2_nand2_1 _1807_ (.Y(_0355_),
    .A(\CIC.u_differentiator.a_mux4to1.d1[12] ),
    .B(net352));
 sg13g2_a22oi_1 _1808_ (.Y(_0356_),
    .B1(net358),
    .B2(net164),
    .A2(net361),
    .A1(net86));
 sg13g2_a21oi_1 _1809_ (.A1(_0355_),
    .A2(_0356_),
    .Y(_0357_),
    .B1(net312));
 sg13g2_a21o_1 _1810_ (.A2(net312),
    .A1(net210),
    .B1(_0357_),
    .X(_0144_));
 sg13g2_nand2_1 _1811_ (.Y(_0358_),
    .A(net166),
    .B(net351));
 sg13g2_nor2b_1 _1812_ (.A(_0024_),
    .B_N(net358),
    .Y(_0359_));
 sg13g2_o21ai_1 _1813_ (.B1(_0358_),
    .Y(_0360_),
    .A1(_0023_),
    .A2(net359));
 sg13g2_nor3_1 _1814_ (.A(net311),
    .B(_0359_),
    .C(_0360_),
    .Y(_0361_));
 sg13g2_a21oi_1 _1815_ (.A1(_0468_),
    .A2(net311),
    .Y(_0145_),
    .B1(_0361_));
 sg13g2_nand2_1 _1816_ (.Y(_0362_),
    .A(\CIC.u_differentiator.a_mux4to1.d1[14] ),
    .B(net351));
 sg13g2_a22oi_1 _1817_ (.Y(_0363_),
    .B1(net356),
    .B2(net91),
    .A2(net361),
    .A1(net142));
 sg13g2_a21oi_1 _1818_ (.A1(_0362_),
    .A2(_0363_),
    .Y(_0364_),
    .B1(net311));
 sg13g2_a21o_1 _1819_ (.A2(net311),
    .A1(net220),
    .B1(_0364_),
    .X(_0146_));
 sg13g2_nand2b_1 _1820_ (.Y(_0365_),
    .B(net356),
    .A_N(_0026_));
 sg13g2_o21ai_1 _1821_ (.B1(_0365_),
    .Y(_0366_),
    .A1(_0025_),
    .A2(net359));
 sg13g2_a21oi_1 _1822_ (.A1(\CIC.u_differentiator.a_mux4to1.d1[15] ),
    .A2(net351),
    .Y(_0367_),
    .B1(_0366_));
 sg13g2_nand2_1 _1823_ (.Y(_0368_),
    .A(net107),
    .B(net311));
 sg13g2_o21ai_1 _1824_ (.B1(_0368_),
    .Y(_0147_),
    .A1(net311),
    .A2(_0367_));
 sg13g2_nand2_1 _1825_ (.Y(_0369_),
    .A(\CIC.u_differentiator.a_mux4to1.d1[16] ),
    .B(net350));
 sg13g2_a22oi_1 _1826_ (.Y(_0370_),
    .B1(net355),
    .B2(net134),
    .A2(net360),
    .A1(net97));
 sg13g2_a21oi_1 _1827_ (.A1(_0369_),
    .A2(_0370_),
    .Y(_0371_),
    .B1(net310));
 sg13g2_a21o_1 _1828_ (.A2(net316),
    .A1(net180),
    .B1(_0371_),
    .X(_0148_));
 sg13g2_nand2_1 _1829_ (.Y(_0372_),
    .A(net88),
    .B(net310));
 sg13g2_nand2b_1 _1830_ (.Y(_0373_),
    .B(net355),
    .A_N(_0028_));
 sg13g2_o21ai_1 _1831_ (.B1(_0373_),
    .Y(_0374_),
    .A1(_0027_),
    .A2(net359));
 sg13g2_a21oi_1 _1832_ (.A1(\CIC.u_differentiator.a_mux4to1.d1[17] ),
    .A2(net350),
    .Y(_0375_),
    .B1(_0374_));
 sg13g2_o21ai_1 _1833_ (.B1(_0372_),
    .Y(_0149_),
    .A1(net310),
    .A2(_0375_));
 sg13g2_nand2_1 _1834_ (.Y(_0376_),
    .A(\CIC.u_differentiator.a_mux4to1.d1[18] ),
    .B(net350));
 sg13g2_a22oi_1 _1835_ (.Y(_0377_),
    .B1(net355),
    .B2(net100),
    .A2(net360),
    .A1(net80));
 sg13g2_a21oi_1 _1836_ (.A1(_0376_),
    .A2(_0377_),
    .Y(_0378_),
    .B1(net310));
 sg13g2_a21o_1 _1837_ (.A2(net310),
    .A1(net222),
    .B1(_0378_),
    .X(_0150_));
 sg13g2_nand2b_1 _1838_ (.Y(_0379_),
    .B(net355),
    .A_N(_0030_));
 sg13g2_o21ai_1 _1839_ (.B1(_0379_),
    .Y(_0380_),
    .A1(_0029_),
    .A2(net359));
 sg13g2_a21oi_1 _1840_ (.A1(\CIC.u_differentiator.a_mux4to1.d1[19] ),
    .A2(net350),
    .Y(_0381_),
    .B1(_0380_));
 sg13g2_nand2_1 _1841_ (.Y(_0382_),
    .A(net84),
    .B(net310));
 sg13g2_o21ai_1 _1842_ (.B1(_0382_),
    .Y(_0151_),
    .A1(net310),
    .A2(_0381_));
 sg13g2_nand2_1 _1843_ (.Y(_0383_),
    .A(\CIC.u_differentiator.a_mux4to1.d1[20] ),
    .B(net350));
 sg13g2_a22oi_1 _1844_ (.Y(_0384_),
    .B1(net355),
    .B2(net128),
    .A2(net360),
    .A1(net99));
 sg13g2_a21oi_1 _1845_ (.A1(_0383_),
    .A2(_0384_),
    .Y(_0385_),
    .B1(net309));
 sg13g2_a21o_1 _1846_ (.A2(net309),
    .A1(net239),
    .B1(_0385_),
    .X(_0152_));
 sg13g2_nand2_1 _1847_ (.Y(_0386_),
    .A(net130),
    .B(net355));
 sg13g2_a22oi_1 _1848_ (.Y(_0387_),
    .B1(net350),
    .B2(\CIC.u_differentiator.a_mux4to1.d1[21] ),
    .A2(net360),
    .A1(net112));
 sg13g2_a21oi_1 _1849_ (.A1(_0386_),
    .A2(_0387_),
    .Y(_0388_),
    .B1(net309));
 sg13g2_a21o_1 _1850_ (.A2(net309),
    .A1(net224),
    .B1(_0388_),
    .X(_0153_));
 sg13g2_nand2_1 _1851_ (.Y(_0389_),
    .A(\CIC.u_differentiator.a_mux4to1.d1[22] ),
    .B(net350));
 sg13g2_a22oi_1 _1852_ (.Y(_0390_),
    .B1(net355),
    .B2(net121),
    .A2(net360),
    .A1(net101));
 sg13g2_a21oi_1 _1853_ (.A1(_0389_),
    .A2(_0390_),
    .Y(_0391_),
    .B1(net309));
 sg13g2_a21o_1 _1854_ (.A2(net309),
    .A1(net208),
    .B1(_0391_),
    .X(_0154_));
 sg13g2_nand2_1 _1855_ (.Y(_0392_),
    .A(net90),
    .B(net356));
 sg13g2_a22oi_1 _1856_ (.Y(_0393_),
    .B1(net350),
    .B2(\CIC.u_differentiator.a_mux4to1.d1[23] ),
    .A2(net360),
    .A1(\CIC.u_differentiator.a_mux4to1.d3[23] ));
 sg13g2_a21oi_1 _1857_ (.A1(_0392_),
    .A2(_0393_),
    .Y(_0394_),
    .B1(net309));
 sg13g2_a21o_1 _1858_ (.A2(net309),
    .A1(net125),
    .B1(_0394_),
    .X(_0155_));
 sg13g2_and4_1 _1859_ (.A(net395),
    .B(net453),
    .C(_0730_),
    .D(net366),
    .X(_0395_));
 sg13g2_nor2_1 _1860_ (.A(net113),
    .B(net323),
    .Y(_0396_));
 sg13g2_a21oi_1 _1861_ (.A1(_0744_),
    .A2(net323),
    .Y(_0156_),
    .B1(_0396_));
 sg13g2_nor2_1 _1862_ (.A(net59),
    .B(net322),
    .Y(_0397_));
 sg13g2_a21oi_1 _1863_ (.A1(_0754_),
    .A2(net323),
    .Y(_0157_),
    .B1(_0397_));
 sg13g2_nor2_1 _1864_ (.A(net102),
    .B(net322),
    .Y(_0398_));
 sg13g2_a21oi_1 _1865_ (.A1(_0764_),
    .A2(net323),
    .Y(_0158_),
    .B1(_0398_));
 sg13g2_nor2_1 _1866_ (.A(net70),
    .B(net321),
    .Y(_0399_));
 sg13g2_a21oi_1 _1867_ (.A1(_0773_),
    .A2(net321),
    .Y(_0159_),
    .B1(_0399_));
 sg13g2_nor2_1 _1868_ (.A(net74),
    .B(net322),
    .Y(_0400_));
 sg13g2_a21oi_1 _1869_ (.A1(_0781_),
    .A2(net324),
    .Y(_0160_),
    .B1(_0400_));
 sg13g2_nor2_1 _1870_ (.A(net82),
    .B(net324),
    .Y(_0401_));
 sg13g2_a21oi_1 _1871_ (.A1(_0789_),
    .A2(net324),
    .Y(_0161_),
    .B1(_0401_));
 sg13g2_nor2_1 _1872_ (.A(net67),
    .B(net319),
    .Y(_0402_));
 sg13g2_a21oi_1 _1873_ (.A1(_0802_),
    .A2(net319),
    .Y(_0162_),
    .B1(_0402_));
 sg13g2_nor2_1 _1874_ (.A(net76),
    .B(net319),
    .Y(_0403_));
 sg13g2_a21oi_1 _1875_ (.A1(_0809_),
    .A2(net319),
    .Y(_0163_),
    .B1(_0403_));
 sg13g2_nor2_1 _1876_ (.A(net58),
    .B(net322),
    .Y(_0404_));
 sg13g2_a21oi_1 _1877_ (.A1(_0825_),
    .A2(net322),
    .Y(_0164_),
    .B1(_0404_));
 sg13g2_nor2_1 _1878_ (.A(net65),
    .B(net322),
    .Y(_0405_));
 sg13g2_a21oi_1 _1879_ (.A1(_0832_),
    .A2(net322),
    .Y(_0165_),
    .B1(_0405_));
 sg13g2_nor2_1 _1880_ (.A(net63),
    .B(net322),
    .Y(_0406_));
 sg13g2_a21oi_1 _1881_ (.A1(_0845_),
    .A2(net325),
    .Y(_0166_),
    .B1(_0406_));
 sg13g2_nor2_1 _1882_ (.A(net56),
    .B(net321),
    .Y(_0407_));
 sg13g2_a21oi_1 _1883_ (.A1(_0854_),
    .A2(net321),
    .Y(_0167_),
    .B1(_0407_));
 sg13g2_nor2_1 _1884_ (.A(net55),
    .B(net321),
    .Y(_0408_));
 sg13g2_a21oi_1 _1885_ (.A1(_0866_),
    .A2(net321),
    .Y(_0168_),
    .B1(_0408_));
 sg13g2_nor2_1 _1886_ (.A(net62),
    .B(net321),
    .Y(_0409_));
 sg13g2_a21oi_1 _1887_ (.A1(_0874_),
    .A2(net321),
    .Y(_0169_),
    .B1(_0409_));
 sg13g2_nor2_1 _1888_ (.A(net68),
    .B(net320),
    .Y(_0410_));
 sg13g2_a21oi_1 _1889_ (.A1(_0888_),
    .A2(net320),
    .Y(_0170_),
    .B1(_0410_));
 sg13g2_nor2_1 _1890_ (.A(net61),
    .B(net319),
    .Y(_0411_));
 sg13g2_a21oi_1 _1891_ (.A1(_0896_),
    .A2(net319),
    .Y(_0171_),
    .B1(_0411_));
 sg13g2_nor2_1 _1892_ (.A(net69),
    .B(net325),
    .Y(_0412_));
 sg13g2_a21oi_1 _1893_ (.A1(_0234_),
    .A2(net325),
    .Y(_0172_),
    .B1(_0412_));
 sg13g2_nor2_1 _1894_ (.A(net83),
    .B(net319),
    .Y(_0413_));
 sg13g2_a21oi_1 _1895_ (.A1(_0245_),
    .A2(net317),
    .Y(_0173_),
    .B1(_0413_));
 sg13g2_nor2_1 _1896_ (.A(net129),
    .B(net319),
    .Y(_0414_));
 sg13g2_a21oi_1 _1897_ (.A1(_0257_),
    .A2(net318),
    .Y(_0174_),
    .B1(_0414_));
 sg13g2_nor2_1 _1898_ (.A(net79),
    .B(net317),
    .Y(_0415_));
 sg13g2_a21oi_1 _1899_ (.A1(_0266_),
    .A2(net317),
    .Y(_0175_),
    .B1(_0415_));
 sg13g2_nor2_1 _1900_ (.A(net111),
    .B(net317),
    .Y(_0416_));
 sg13g2_a21oi_1 _1901_ (.A1(_0277_),
    .A2(net318),
    .Y(_0176_),
    .B1(_0416_));
 sg13g2_nor2_1 _1902_ (.A(net71),
    .B(net317),
    .Y(_0417_));
 sg13g2_a21oi_1 _1903_ (.A1(_0286_),
    .A2(net317),
    .Y(_0177_),
    .B1(_0417_));
 sg13g2_nor2_1 _1904_ (.A(net115),
    .B(net318),
    .Y(_0418_));
 sg13g2_a21oi_1 _1905_ (.A1(_0297_),
    .A2(net318),
    .Y(_0178_),
    .B1(_0418_));
 sg13g2_nor2_1 _1906_ (.A(net87),
    .B(net317),
    .Y(_0419_));
 sg13g2_a21oi_1 _1907_ (.A1(_0305_),
    .A2(net317),
    .Y(_0179_),
    .B1(_0419_));
 sg13g2_nor2_1 _1908_ (.A(net136),
    .B(net331),
    .Y(_0420_));
 sg13g2_a21oi_1 _1909_ (.A1(_0744_),
    .A2(net331),
    .Y(_0180_),
    .B1(_0420_));
 sg13g2_nor2_1 _1910_ (.A(net46),
    .B(net330),
    .Y(_0421_));
 sg13g2_a21oi_1 _1911_ (.A1(_0754_),
    .A2(net330),
    .Y(_0181_),
    .B1(_0421_));
 sg13g2_nor2_1 _1912_ (.A(net201),
    .B(net331),
    .Y(_0422_));
 sg13g2_a21oi_1 _1913_ (.A1(_0764_),
    .A2(net331),
    .Y(_0182_),
    .B1(_0422_));
 sg13g2_nor2_1 _1914_ (.A(net49),
    .B(net330),
    .Y(_0423_));
 sg13g2_a21oi_1 _1915_ (.A1(_0773_),
    .A2(net330),
    .Y(_0183_),
    .B1(_0423_));
 sg13g2_nor2_1 _1916_ (.A(net109),
    .B(net330),
    .Y(_0424_));
 sg13g2_a21oi_1 _1917_ (.A1(_0781_),
    .A2(net329),
    .Y(_0184_),
    .B1(_0424_));
 sg13g2_nor2_1 _1918_ (.A(net50),
    .B(net330),
    .Y(_0425_));
 sg13g2_a21oi_1 _1919_ (.A1(_0789_),
    .A2(net330),
    .Y(_0185_),
    .B1(_0425_));
 sg13g2_nor2_1 _1920_ (.A(net78),
    .B(net329),
    .Y(_0426_));
 sg13g2_a21oi_1 _1921_ (.A1(_0802_),
    .A2(net329),
    .Y(_0186_),
    .B1(_0426_));
 sg13g2_nor2_1 _1922_ (.A(net64),
    .B(net329),
    .Y(_0427_));
 sg13g2_a21oi_1 _1923_ (.A1(_0809_),
    .A2(net329),
    .Y(_0187_),
    .B1(_0427_));
 sg13g2_nor2_1 _1924_ (.A(net106),
    .B(net329),
    .Y(_0428_));
 sg13g2_a21oi_1 _1925_ (.A1(_0825_),
    .A2(net329),
    .Y(_0188_),
    .B1(_0428_));
 sg13g2_nor2_1 _1926_ (.A(net52),
    .B(net329),
    .Y(_0429_));
 sg13g2_a21oi_1 _1927_ (.A1(_0832_),
    .A2(net332),
    .Y(_0189_),
    .B1(_0429_));
 sg13g2_nor2_1 _1928_ (.A(net135),
    .B(net332),
    .Y(_0430_));
 sg13g2_a21oi_1 _1929_ (.A1(_0845_),
    .A2(net332),
    .Y(_0190_),
    .B1(_0430_));
 sg13g2_nor2_1 _1930_ (.A(net75),
    .B(net328),
    .Y(_0431_));
 sg13g2_a21oi_1 _1931_ (.A1(_0854_),
    .A2(net328),
    .Y(_0191_),
    .B1(_0431_));
 sg13g2_nor2_1 _1932_ (.A(net164),
    .B(net332),
    .Y(_0432_));
 sg13g2_a21oi_1 _1933_ (.A1(_0866_),
    .A2(net332),
    .Y(_0192_),
    .B1(_0432_));
 sg13g2_nor2_1 _1934_ (.A(net51),
    .B(net332),
    .Y(_0433_));
 sg13g2_a21oi_1 _1935_ (.A1(_0874_),
    .A2(net332),
    .Y(_0193_),
    .B1(_0433_));
 sg13g2_nor2_1 _1936_ (.A(net91),
    .B(net328),
    .Y(_0434_));
 sg13g2_a21oi_1 _1937_ (.A1(_0888_),
    .A2(net328),
    .Y(_0194_),
    .B1(_0434_));
 sg13g2_nor2_1 _1938_ (.A(net45),
    .B(net328),
    .Y(_0435_));
 sg13g2_a21oi_1 _1939_ (.A1(_0896_),
    .A2(net328),
    .Y(_0195_),
    .B1(_0435_));
 sg13g2_nor2_1 _1940_ (.A(net134),
    .B(net333),
    .Y(_0436_));
 sg13g2_a21oi_1 _1941_ (.A1(_0234_),
    .A2(net333),
    .Y(_0196_),
    .B1(_0436_));
 sg13g2_nor2_1 _1942_ (.A(net66),
    .B(net326),
    .Y(_0437_));
 sg13g2_a21oi_1 _1943_ (.A1(_0245_),
    .A2(net326),
    .Y(_0197_),
    .B1(_0437_));
 sg13g2_nor2_1 _1944_ (.A(net100),
    .B(net326),
    .Y(_0438_));
 sg13g2_a21oi_1 _1945_ (.A1(_0257_),
    .A2(net326),
    .Y(_0198_),
    .B1(_0438_));
 sg13g2_nor2_1 _1946_ (.A(net77),
    .B(net326),
    .Y(_0439_));
 sg13g2_a21oi_1 _1947_ (.A1(_0266_),
    .A2(net326),
    .Y(_0199_),
    .B1(_0439_));
 sg13g2_nor2_1 _1948_ (.A(net128),
    .B(net327),
    .Y(_0440_));
 sg13g2_a21oi_1 _1949_ (.A1(_0277_),
    .A2(net326),
    .Y(_0200_),
    .B1(_0440_));
 sg13g2_nor2_1 _1950_ (.A(net130),
    .B(net327),
    .Y(_0441_));
 sg13g2_a21oi_1 _1951_ (.A1(_0286_),
    .A2(net327),
    .Y(_0201_),
    .B1(_0441_));
 sg13g2_nor2_1 _1952_ (.A(net121),
    .B(net327),
    .Y(_0442_));
 sg13g2_a21oi_1 _1953_ (.A1(_0297_),
    .A2(net326),
    .Y(_0202_),
    .B1(_0442_));
 sg13g2_nor2_1 _1954_ (.A(net90),
    .B(net327),
    .Y(_0443_));
 sg13g2_a21oi_1 _1955_ (.A1(_0305_),
    .A2(net327),
    .Y(_0203_),
    .B1(_0443_));
 sg13g2_nand3_1 _1956_ (.B(_0306_),
    .C(net351),
    .A(_0730_),
    .Y(_0444_));
 sg13g2_a21oi_1 _1957_ (.A1(net182),
    .A2(net366),
    .Y(_0445_),
    .B1(_0444_));
 sg13g2_nor2_1 _1958_ (.A(_0449_),
    .B(_0445_),
    .Y(_0446_));
 sg13g2_a21oi_1 _1959_ (.A1(_0449_),
    .A2(net315),
    .Y(_0204_),
    .B1(_0446_));
 sg13g2_a21o_1 _1960_ (.A2(_0445_),
    .A1(net377),
    .B1(_0310_),
    .X(_0205_));
 sg13g2_a21oi_1 _1961_ (.A1(net182),
    .A2(net366),
    .Y(_0447_),
    .B1(\CIC.u_differentiator.count[2] ));
 sg13g2_nor2_1 _1962_ (.A(_0444_),
    .B(net183),
    .Y(_0206_));
 sg13g2_mux2_1 _1963_ (.A0(net93),
    .A1(net204),
    .S(net337),
    .X(_0207_));
 sg13g2_mux2_1 _1964_ (.A0(\CIC.int_2_out[1] ),
    .A1(net143),
    .S(net336),
    .X(_0208_));
 sg13g2_mux2_1 _1965_ (.A0(net172),
    .A1(\CIC.u_differentiator.a_mux4to1.d1[2] ),
    .S(net336),
    .X(_0209_));
 sg13g2_mux2_1 _1966_ (.A0(\CIC.int_2_out[3] ),
    .A1(net154),
    .S(net336),
    .X(_0210_));
 sg13g2_mux2_1 _1967_ (.A0(net216),
    .A1(\CIC.u_differentiator.a_mux4to1.d1[4] ),
    .S(net337),
    .X(_0211_));
 sg13g2_mux2_1 _1968_ (.A0(\CIC.int_2_out[5] ),
    .A1(net123),
    .S(net337),
    .X(_0212_));
 sg13g2_mux2_1 _1969_ (.A0(net140),
    .A1(\CIC.u_differentiator.a_mux4to1.d1[6] ),
    .S(net337),
    .X(_0213_));
 sg13g2_mux2_1 _1970_ (.A0(net199),
    .A1(\CIC.u_differentiator.a_mux4to1.d1[7] ),
    .S(net337),
    .X(_0214_));
 sg13g2_mux2_1 _1971_ (.A0(net197),
    .A1(\CIC.u_differentiator.a_mux4to1.d1[8] ),
    .S(net336),
    .X(_0215_));
 sg13g2_mux2_1 _1972_ (.A0(\CIC.int_2_out[9] ),
    .A1(net178),
    .S(net336),
    .X(_0216_));
 sg13g2_mux2_1 _1973_ (.A0(net185),
    .A1(\CIC.u_differentiator.a_mux4to1.d1[10] ),
    .S(net336),
    .X(_0217_));
 sg13g2_mux2_1 _1974_ (.A0(net241),
    .A1(\CIC.u_differentiator.a_mux4to1.d1[11] ),
    .S(net336),
    .X(_0218_));
 sg13g2_mux2_1 _1975_ (.A0(\CIC.int_2_out[12] ),
    .A1(net232),
    .S(net335),
    .X(_0219_));
 sg13g2_mux2_1 _1976_ (.A0(\CIC.int_2_out[13] ),
    .A1(net166),
    .S(net335),
    .X(_0220_));
 sg13g2_mux2_1 _1977_ (.A0(net226),
    .A1(\CIC.u_differentiator.a_mux4to1.d1[14] ),
    .S(net335),
    .X(_0221_));
 sg13g2_mux2_1 _1978_ (.A0(\CIC.int_2_out[15] ),
    .A1(net157),
    .S(net335),
    .X(_0222_));
 sg13g2_mux2_1 _1979_ (.A0(net236),
    .A1(\CIC.u_differentiator.a_mux4to1.d1[16] ),
    .S(net334),
    .X(_0223_));
 sg13g2_mux2_1 _1980_ (.A0(\CIC.int_2_out[17] ),
    .A1(net228),
    .S(net334),
    .X(_0224_));
 sg13g2_mux2_1 _1981_ (.A0(net212),
    .A1(\CIC.u_differentiator.a_mux4to1.d1[18] ),
    .S(net334),
    .X(_0225_));
 sg13g2_mux2_1 _1982_ (.A0(net150),
    .A1(\CIC.u_differentiator.a_mux4to1.d1[19] ),
    .S(net334),
    .X(_0226_));
 sg13g2_mux2_1 _1983_ (.A0(net243),
    .A1(\CIC.u_differentiator.a_mux4to1.d1[20] ),
    .S(net334),
    .X(_0227_));
 sg13g2_mux2_1 _1984_ (.A0(net214),
    .A1(\CIC.u_differentiator.a_mux4to1.d1[21] ),
    .S(net334),
    .X(_0228_));
 sg13g2_mux2_1 _1985_ (.A0(net234),
    .A1(\CIC.u_differentiator.a_mux4to1.d1[22] ),
    .S(net334),
    .X(_0229_));
 sg13g2_mux2_1 _1986_ (.A0(net95),
    .A1(\CIC.u_differentiator.a_mux4to1.d1[23] ),
    .S(net334),
    .X(_0230_));
 sg13g2_dfrbp_1 _1987_ (.CLK(\divideby64.clkOutDiv5 ),
    .RESET_B(net393),
    .D(_0005_),
    .Q_N(_0005_),
    .Q(\CIC.dec_clk ));
 sg13g2_dfrbp_1 _1988_ (.CLK(\divideby64.clkOutDiv4 ),
    .RESET_B(net393),
    .D(_0004_),
    .Q_N(_0004_),
    .Q(\divideby64.clkOutDiv5 ));
 sg13g2_dfrbp_1 _1989_ (.CLK(div_clk8x),
    .RESET_B(net392),
    .D(_0003_),
    .Q_N(_0003_),
    .Q(\divideby64.clkOutDiv4 ));
 sg13g2_dfrbp_1 _1990_ (.CLK(\divideby64.clkOutDiv2 ),
    .RESET_B(net392),
    .D(_0002_),
    .Q_N(_0002_),
    .Q(div_clk8x));
 sg13g2_dfrbp_1 _1991_ (.CLK(\divideby64.clkOutDiv1 ),
    .RESET_B(net392),
    .D(_0001_),
    .Q_N(_0001_),
    .Q(\divideby64.clkOutDiv2 ));
 sg13g2_dfrbp_1 _1992_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net392),
    .D(net40),
    .Q_N(_0000_),
    .Q(\divideby64.clkOutDiv1 ));
 sg13g2_dfrbp_1 _1993_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net411),
    .D(net120),
    .Q_N(_1006_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[0] ));
 sg13g2_dfrbp_1 _1994_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net411),
    .D(net44),
    .Q_N(_0011_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[1] ));
 sg13g2_dfrbp_1 _1995_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net407),
    .D(_0110_),
    .Q_N(_1005_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[2] ));
 sg13g2_dfrbp_1 _1996_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net408),
    .D(_0111_),
    .Q_N(_0013_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[3] ));
 sg13g2_dfrbp_1 _1997_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net408),
    .D(_0112_),
    .Q_N(_1004_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[4] ));
 sg13g2_dfrbp_1 _1998_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net408),
    .D(_0113_),
    .Q_N(_0015_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[5] ));
 sg13g2_dfrbp_1 _1999_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net399),
    .D(_0114_),
    .Q_N(_1003_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[6] ));
 sg13g2_dfrbp_1 _2000_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net400),
    .D(_0115_),
    .Q_N(_0017_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[7] ));
 sg13g2_dfrbp_1 _2001_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net407),
    .D(_0116_),
    .Q_N(_1002_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[8] ));
 sg13g2_dfrbp_1 _2002_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net399),
    .D(_0117_),
    .Q_N(_0019_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[9] ));
 sg13g2_dfrbp_1 _2003_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net406),
    .D(_0118_),
    .Q_N(_1001_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[10] ));
 sg13g2_dfrbp_1 _2004_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net395),
    .D(_0119_),
    .Q_N(_0021_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[11] ));
 sg13g2_dfrbp_1 _2005_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net399),
    .D(_0120_),
    .Q_N(_1000_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[12] ));
 sg13g2_dfrbp_1 _2006_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net389),
    .D(_0121_),
    .Q_N(_0023_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[13] ));
 sg13g2_dfrbp_1 _2007_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net394),
    .D(_0122_),
    .Q_N(_0999_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[14] ));
 sg13g2_dfrbp_1 _2008_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net388),
    .D(_0123_),
    .Q_N(_0025_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[15] ));
 sg13g2_dfrbp_1 _2009_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net394),
    .D(_0124_),
    .Q_N(_0998_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[16] ));
 sg13g2_dfrbp_1 _2010_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net383),
    .D(_0125_),
    .Q_N(_0027_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[17] ));
 sg13g2_dfrbp_1 _2011_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net390),
    .D(_0126_),
    .Q_N(_0997_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[18] ));
 sg13g2_dfrbp_1 _2012_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net390),
    .D(_0127_),
    .Q_N(_0029_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[19] ));
 sg13g2_dfrbp_1 _2013_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net393),
    .D(_0128_),
    .Q_N(_0996_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[20] ));
 sg13g2_dfrbp_1 _2014_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net392),
    .D(_0129_),
    .Q_N(_0995_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[21] ));
 sg13g2_dfrbp_1 _2015_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net393),
    .D(_0130_),
    .Q_N(_0994_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[22] ));
 sg13g2_dfrbp_1 _2016_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net391),
    .D(_0131_),
    .Q_N(_1007_),
    .Q(\CIC.u_differentiator.a_mux4to1.d3[23] ));
 sg13g2_dfrbp_1 _2017_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net395),
    .D(\CIC.dec_clk ),
    .Q_N(_0993_),
    .Q(\CIC.u_differentiator.prev_lr_clk ));
 sg13g2_dfrbp_1 _2018_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net411),
    .D(net177),
    .Q_N(_0992_),
    .Q(\CIC.u_differentiator.temp[0] ));
 sg13g2_dfrbp_1 _2019_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net410),
    .D(net104),
    .Q_N(_0991_),
    .Q(\CIC.u_differentiator.temp[1] ));
 sg13g2_dfrbp_1 _2020_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net406),
    .D(net196),
    .Q_N(_0990_),
    .Q(\CIC.u_differentiator.temp[2] ));
 sg13g2_dfrbp_1 _2021_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net409),
    .D(net163),
    .Q_N(_0989_),
    .Q(\CIC.u_differentiator.temp[3] ));
 sg13g2_dfrbp_1 _2022_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net409),
    .D(net192),
    .Q_N(_0988_),
    .Q(\CIC.u_differentiator.temp[4] ));
 sg13g2_dfrbp_1 _2023_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net409),
    .D(net231),
    .Q_N(_0987_),
    .Q(\CIC.u_differentiator.temp[5] ));
 sg13g2_dfrbp_1 _2024_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net403),
    .D(net190),
    .Q_N(_0986_),
    .Q(\CIC.u_differentiator.temp[6] ));
 sg13g2_dfrbp_1 _2025_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net403),
    .D(net149),
    .Q_N(_0985_),
    .Q(\CIC.u_differentiator.temp[7] ));
 sg13g2_dfrbp_1 _2026_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net407),
    .D(net203),
    .Q_N(_0984_),
    .Q(\CIC.u_differentiator.temp[8] ));
 sg13g2_dfrbp_1 _2027_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net400),
    .D(net146),
    .Q_N(_0983_),
    .Q(\CIC.u_differentiator.temp[9] ));
 sg13g2_dfrbp_1 _2028_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net406),
    .D(net194),
    .Q_N(_0982_),
    .Q(\CIC.u_differentiator.temp[10] ));
 sg13g2_dfrbp_1 _2029_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net395),
    .D(net133),
    .Q_N(_0981_),
    .Q(\CIC.u_differentiator.temp[11] ));
 sg13g2_dfrbp_1 _2030_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net394),
    .D(net211),
    .Q_N(_0980_),
    .Q(\CIC.u_differentiator.temp[12] ));
 sg13g2_dfrbp_1 _2031_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net388),
    .D(net219),
    .Q_N(_0979_),
    .Q(\CIC.u_differentiator.temp[13] ));
 sg13g2_dfrbp_1 _2032_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net388),
    .D(net221),
    .Q_N(_0978_),
    .Q(\CIC.u_differentiator.temp[14] ));
 sg13g2_dfrbp_1 _2033_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net389),
    .D(net108),
    .Q_N(_0977_),
    .Q(\CIC.u_differentiator.temp[15] ));
 sg13g2_dfrbp_1 _2034_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net394),
    .D(net181),
    .Q_N(_0976_),
    .Q(\CIC.u_differentiator.temp[16] ));
 sg13g2_dfrbp_1 _2035_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net384),
    .D(net89),
    .Q_N(_0975_),
    .Q(\CIC.u_differentiator.temp[17] ));
 sg13g2_dfrbp_1 _2036_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net390),
    .D(net223),
    .Q_N(_0974_),
    .Q(\CIC.u_differentiator.temp[18] ));
 sg13g2_dfrbp_1 _2037_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net391),
    .D(net85),
    .Q_N(_0973_),
    .Q(\CIC.u_differentiator.temp[19] ));
 sg13g2_dfrbp_1 _2038_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net393),
    .D(net240),
    .Q_N(_0972_),
    .Q(\CIC.u_differentiator.temp[20] ));
 sg13g2_dfrbp_1 _2039_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net392),
    .D(net225),
    .Q_N(_0971_),
    .Q(\CIC.u_differentiator.temp[21] ));
 sg13g2_dfrbp_1 _2040_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net392),
    .D(net209),
    .Q_N(_0970_),
    .Q(\CIC.u_differentiator.temp[22] ));
 sg13g2_dfrbp_1 _2041_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net390),
    .D(net126),
    .Q_N(_0969_),
    .Q(\CIC.u_differentiator.temp[23] ));
 sg13g2_dfrbp_1 _2042_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net37),
    .D(net114),
    .Q_N(_0968_),
    .Q(\CIC.out[0] ));
 sg13g2_dfrbp_1 _2043_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net36),
    .D(net60),
    .Q_N(_0967_),
    .Q(\CIC.out[1] ));
 sg13g2_dfrbp_1 _2044_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net35),
    .D(_0158_),
    .Q_N(_0966_),
    .Q(\CIC.out[2] ));
 sg13g2_dfrbp_1 _2045_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net34),
    .D(_0159_),
    .Q_N(_0965_),
    .Q(\CIC.out[3] ));
 sg13g2_dfrbp_1 _2046_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net33),
    .D(_0160_),
    .Q_N(_0964_),
    .Q(\CIC.out[4] ));
 sg13g2_dfrbp_1 _2047_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net32),
    .D(_0161_),
    .Q_N(_0963_),
    .Q(\CIC.out[5] ));
 sg13g2_dfrbp_1 _2048_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net31),
    .D(_0162_),
    .Q_N(_0962_),
    .Q(\CIC.out[6] ));
 sg13g2_dfrbp_1 _2049_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net30),
    .D(_0163_),
    .Q_N(_0961_),
    .Q(\CIC.out[7] ));
 sg13g2_dfrbp_1 _2050_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net29),
    .D(_0164_),
    .Q_N(_0960_),
    .Q(\CIC.out[8] ));
 sg13g2_dfrbp_1 _2051_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net28),
    .D(_0165_),
    .Q_N(_0959_),
    .Q(\CIC.out[9] ));
 sg13g2_dfrbp_1 _2052_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net27),
    .D(_0166_),
    .Q_N(_0958_),
    .Q(\CIC.out[10] ));
 sg13g2_dfrbp_1 _2053_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net26),
    .D(_0167_),
    .Q_N(_0957_),
    .Q(\CIC.out[11] ));
 sg13g2_dfrbp_1 _2054_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net25),
    .D(_0168_),
    .Q_N(_0956_),
    .Q(\CIC.out[12] ));
 sg13g2_dfrbp_1 _2055_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net24),
    .D(_0169_),
    .Q_N(_0955_),
    .Q(\CIC.out[13] ));
 sg13g2_dfrbp_1 _2056_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net23),
    .D(_0170_),
    .Q_N(_0954_),
    .Q(\CIC.out[14] ));
 sg13g2_dfrbp_1 _2057_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net22),
    .D(_0171_),
    .Q_N(_0953_),
    .Q(\CIC.out[15] ));
 sg13g2_dfrbp_1 _2058_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net21),
    .D(_0172_),
    .Q_N(_0952_),
    .Q(\CIC.out[16] ));
 sg13g2_dfrbp_1 _2059_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net20),
    .D(_0173_),
    .Q_N(_0951_),
    .Q(\CIC.out[17] ));
 sg13g2_dfrbp_1 _2060_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net19),
    .D(_0174_),
    .Q_N(_0950_),
    .Q(\CIC.out[18] ));
 sg13g2_dfrbp_1 _2061_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net18),
    .D(_0175_),
    .Q_N(_0949_),
    .Q(\CIC.out[19] ));
 sg13g2_dfrbp_1 _2062_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net17),
    .D(_0176_),
    .Q_N(_0948_),
    .Q(\CIC.out[20] ));
 sg13g2_dfrbp_1 _2063_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net16),
    .D(_0177_),
    .Q_N(_0947_),
    .Q(\CIC.out[21] ));
 sg13g2_dfrbp_1 _2064_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net15),
    .D(_0178_),
    .Q_N(_0946_),
    .Q(\CIC.out[22] ));
 sg13g2_dfrbp_1 _2065_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net14),
    .D(_0179_),
    .Q_N(_0945_),
    .Q(\CIC.out[23] ));
 sg13g2_dfrbp_1 _2066_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net411),
    .D(net137),
    .Q_N(_0944_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[0] ));
 sg13g2_dfrbp_1 _2067_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net411),
    .D(net47),
    .Q_N(_0012_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[1] ));
 sg13g2_dfrbp_1 _2068_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net407),
    .D(_0182_),
    .Q_N(_0943_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[2] ));
 sg13g2_dfrbp_1 _2069_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net408),
    .D(_0183_),
    .Q_N(_0014_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[3] ));
 sg13g2_dfrbp_1 _2070_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net408),
    .D(_0184_),
    .Q_N(_0942_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[4] ));
 sg13g2_dfrbp_1 _2071_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net408),
    .D(_0185_),
    .Q_N(_0016_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[5] ));
 sg13g2_dfrbp_1 _2072_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net403),
    .D(_0186_),
    .Q_N(_0941_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[6] ));
 sg13g2_dfrbp_1 _2073_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net399),
    .D(_0187_),
    .Q_N(_0018_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[7] ));
 sg13g2_dfrbp_1 _2074_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net406),
    .D(_0188_),
    .Q_N(_0940_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[8] ));
 sg13g2_dfrbp_1 _2075_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net400),
    .D(_0189_),
    .Q_N(_0020_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[9] ));
 sg13g2_dfrbp_1 _2076_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net406),
    .D(_0190_),
    .Q_N(_0939_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[10] ));
 sg13g2_dfrbp_1 _2077_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net394),
    .D(_0191_),
    .Q_N(_0022_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[11] ));
 sg13g2_dfrbp_1 _2078_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net406),
    .D(_0192_),
    .Q_N(_0938_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[12] ));
 sg13g2_dfrbp_1 _2079_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net399),
    .D(_0193_),
    .Q_N(_0024_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[13] ));
 sg13g2_dfrbp_1 _2080_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net394),
    .D(_0194_),
    .Q_N(_0937_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[14] ));
 sg13g2_dfrbp_1 _2081_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net388),
    .D(_0195_),
    .Q_N(_0026_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[15] ));
 sg13g2_dfrbp_1 _2082_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net394),
    .D(_0196_),
    .Q_N(_0936_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[16] ));
 sg13g2_dfrbp_1 _2083_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net391),
    .D(_0197_),
    .Q_N(_0028_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[17] ));
 sg13g2_dfrbp_1 _2084_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net390),
    .D(_0198_),
    .Q_N(_0935_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[18] ));
 sg13g2_dfrbp_1 _2085_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net390),
    .D(_0199_),
    .Q_N(_0030_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[19] ));
 sg13g2_dfrbp_1 _2086_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net393),
    .D(_0200_),
    .Q_N(_0934_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[20] ));
 sg13g2_dfrbp_1 _2087_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net392),
    .D(_0201_),
    .Q_N(_0933_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[21] ));
 sg13g2_dfrbp_1 _2088_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net393),
    .D(_0202_),
    .Q_N(_0932_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[22] ));
 sg13g2_dfrbp_1 _2089_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net390),
    .D(_0203_),
    .Q_N(_0931_),
    .Q(\CIC.u_differentiator.a_mux4to1.d2[23] ));
 sg13g2_dfrbp_1 _2090_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net406),
    .D(_0204_),
    .Q_N(_0930_),
    .Q(\CIC.u_differentiator.a_mux4to1.sel[0] ));
 sg13g2_dfrbp_1 _2091_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net406),
    .D(_0205_),
    .Q_N(_0929_),
    .Q(\CIC.u_differentiator.a_mux4to1.sel[1] ));
 sg13g2_dfrbp_1 _2092_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net394),
    .D(net184),
    .Q_N(_0009_),
    .Q(\CIC.u_differentiator.count[2] ));
 sg13g2_dfrbp_1 _2093_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net410),
    .D(_0207_),
    .Q_N(_0928_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[0] ));
 sg13g2_dfrbp_1 _2094_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net410),
    .D(net144),
    .Q_N(_0031_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[1] ));
 sg13g2_dfrbp_1 _2095_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net409),
    .D(net173),
    .Q_N(_0927_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[2] ));
 sg13g2_dfrbp_1 _2096_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net409),
    .D(net155),
    .Q_N(_0032_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[3] ));
 sg13g2_dfrbp_1 _2097_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net404),
    .D(net217),
    .Q_N(_0926_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[4] ));
 sg13g2_dfrbp_1 _2098_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net404),
    .D(net124),
    .Q_N(_0033_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[5] ));
 sg13g2_dfrbp_1 _2099_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net403),
    .D(net141),
    .Q_N(_0925_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[6] ));
 sg13g2_dfrbp_1 _2100_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net403),
    .D(net200),
    .Q_N(_0924_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[7] ));
 sg13g2_dfrbp_1 _2101_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net400),
    .D(net198),
    .Q_N(_0923_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[8] ));
 sg13g2_dfrbp_1 _2102_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net400),
    .D(net179),
    .Q_N(_0006_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[9] ));
 sg13g2_dfrbp_1 _2103_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net399),
    .D(net186),
    .Q_N(_0922_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[10] ));
 sg13g2_dfrbp_1 _2104_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net399),
    .D(net242),
    .Q_N(_0921_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[11] ));
 sg13g2_dfrbp_1 _2105_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net399),
    .D(net233),
    .Q_N(_0920_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[12] ));
 sg13g2_dfrbp_1 _2106_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net388),
    .D(net167),
    .Q_N(_0007_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[13] ));
 sg13g2_dfrbp_1 _2107_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net388),
    .D(net227),
    .Q_N(_0919_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[14] ));
 sg13g2_dfrbp_1 _2108_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net389),
    .D(net158),
    .Q_N(_0008_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[15] ));
 sg13g2_dfrbp_1 _2109_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net388),
    .D(net237),
    .Q_N(_0918_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[16] ));
 sg13g2_dfrbp_1 _2110_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net384),
    .D(net229),
    .Q_N(_0917_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[17] ));
 sg13g2_dfrbp_1 _2111_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net384),
    .D(net213),
    .Q_N(_0916_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[18] ));
 sg13g2_dfrbp_1 _2112_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net384),
    .D(net151),
    .Q_N(_0915_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[19] ));
 sg13g2_dfrbp_1 _2113_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net384),
    .D(net244),
    .Q_N(_0914_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[20] ));
 sg13g2_dfrbp_1 _2114_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net383),
    .D(net215),
    .Q_N(_0913_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[21] ));
 sg13g2_dfrbp_1 _2115_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net383),
    .D(net235),
    .Q_N(_0912_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[22] ));
 sg13g2_dfrbp_1 _2116_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net390),
    .D(net96),
    .Q_N(_1008_),
    .Q(\CIC.u_differentiator.a_mux4to1.d1[23] ));
 sg13g2_dfrbp_1 _2117_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net411),
    .D(net94),
    .Q_N(_1009_),
    .Q(\CIC.int_2_out[0] ));
 sg13g2_dfrbp_1 _2118_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net410),
    .D(_0093_),
    .Q_N(_1010_),
    .Q(\CIC.int_2_out[1] ));
 sg13g2_dfrbp_1 _2119_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net408),
    .D(net424),
    .Q_N(_1011_),
    .Q(\CIC.int_2_out[2] ));
 sg13g2_dfrbp_1 _2120_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net408),
    .D(net274),
    .Q_N(_1012_),
    .Q(\CIC.int_2_out[3] ));
 sg13g2_dfrbp_1 _2121_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net404),
    .D(_0100_),
    .Q_N(_1013_),
    .Q(\CIC.int_2_out[4] ));
 sg13g2_dfrbp_1 _2122_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net404),
    .D(net282),
    .Q_N(_1014_),
    .Q(\CIC.int_2_out[5] ));
 sg13g2_dfrbp_1 _2123_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net403),
    .D(net433),
    .Q_N(_1015_),
    .Q(\CIC.int_2_out[6] ));
 sg13g2_dfrbp_1 _2124_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net402),
    .D(_0103_),
    .Q_N(_1016_),
    .Q(\CIC.int_2_out[7] ));
 sg13g2_dfrbp_1 _2125_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net398),
    .D(_0104_),
    .Q_N(_1017_),
    .Q(\CIC.int_2_out[8] ));
 sg13g2_dfrbp_1 _2126_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net398),
    .D(_0105_),
    .Q_N(_1018_),
    .Q(\CIC.int_2_out[9] ));
 sg13g2_dfrbp_1 _2127_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net397),
    .D(_0083_),
    .Q_N(_1019_),
    .Q(\CIC.int_2_out[10] ));
 sg13g2_dfrbp_1 _2128_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net397),
    .D(_0084_),
    .Q_N(_1020_),
    .Q(\CIC.int_2_out[11] ));
 sg13g2_dfrbp_1 _2129_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net387),
    .D(_0085_),
    .Q_N(_1021_),
    .Q(\CIC.int_2_out[12] ));
 sg13g2_dfrbp_1 _2130_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net386),
    .D(net418),
    .Q_N(_1022_),
    .Q(\CIC.int_2_out[13] ));
 sg13g2_dfrbp_1 _2131_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net386),
    .D(_0087_),
    .Q_N(_1023_),
    .Q(\CIC.int_2_out[14] ));
 sg13g2_dfrbp_1 _2132_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net387),
    .D(_0088_),
    .Q_N(_1024_),
    .Q(\CIC.int_2_out[15] ));
 sg13g2_dfrbp_1 _2133_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net386),
    .D(_0089_),
    .Q_N(_1025_),
    .Q(\CIC.int_2_out[16] ));
 sg13g2_dfrbp_1 _2134_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net388),
    .D(_0090_),
    .Q_N(_1026_),
    .Q(\CIC.int_2_out[17] ));
 sg13g2_dfrbp_1 _2135_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net384),
    .D(_0091_),
    .Q_N(_1027_),
    .Q(\CIC.int_2_out[18] ));
 sg13g2_dfrbp_1 _2136_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net384),
    .D(_0092_),
    .Q_N(_1028_),
    .Q(\CIC.int_2_out[19] ));
 sg13g2_dfrbp_1 _2137_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net383),
    .D(_0094_),
    .Q_N(_1029_),
    .Q(\CIC.int_2_out[20] ));
 sg13g2_dfrbp_1 _2138_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net383),
    .D(net420),
    .Q_N(_1030_),
    .Q(\CIC.int_2_out[21] ));
 sg13g2_dfrbp_1 _2139_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net383),
    .D(net271),
    .Q_N(_1031_),
    .Q(\CIC.int_2_out[22] ));
 sg13g2_dfrbp_1 _2140_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net383),
    .D(_0097_),
    .Q_N(_1032_),
    .Q(\CIC.int_2_out[23] ));
 sg13g2_dfrbp_1 _2141_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net411),
    .D(net171),
    .Q_N(_1033_),
    .Q(\CIC.int_1_out[0] ));
 sg13g2_dfrbp_1 _2142_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net410),
    .D(_0069_),
    .Q_N(_1034_),
    .Q(\CIC.int_1_out[1] ));
 sg13g2_dfrbp_1 _2143_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net410),
    .D(_0074_),
    .Q_N(_1035_),
    .Q(\CIC.int_1_out[2] ));
 sg13g2_dfrbp_1 _2144_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net403),
    .D(net279),
    .Q_N(_1036_),
    .Q(\CIC.int_1_out[3] ));
 sg13g2_dfrbp_1 _2145_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net404),
    .D(_0076_),
    .Q_N(_1037_),
    .Q(\CIC.int_1_out[4] ));
 sg13g2_dfrbp_1 _2146_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net405),
    .D(net299),
    .Q_N(_1038_),
    .Q(\CIC.int_1_out[5] ));
 sg13g2_dfrbp_1 _2147_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net402),
    .D(net439),
    .Q_N(_1039_),
    .Q(\CIC.int_1_out[6] ));
 sg13g2_dfrbp_1 _2148_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net402),
    .D(_0079_),
    .Q_N(_1040_),
    .Q(\CIC.int_1_out[7] ));
 sg13g2_dfrbp_1 _2149_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net398),
    .D(_0080_),
    .Q_N(_1041_),
    .Q(\CIC.int_1_out[8] ));
 sg13g2_dfrbp_1 _2150_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net398),
    .D(net277),
    .Q_N(_1042_),
    .Q(\CIC.int_1_out[9] ));
 sg13g2_dfrbp_1 _2151_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net397),
    .D(_0059_),
    .Q_N(_1043_),
    .Q(\CIC.int_1_out[10] ));
 sg13g2_dfrbp_1 _2152_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net397),
    .D(_0060_),
    .Q_N(_1044_),
    .Q(\CIC.int_1_out[11] ));
 sg13g2_dfrbp_1 _2153_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net387),
    .D(_0061_),
    .Q_N(_1045_),
    .Q(\CIC.int_1_out[12] ));
 sg13g2_dfrbp_1 _2154_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net387),
    .D(net297),
    .Q_N(_1046_),
    .Q(\CIC.int_1_out[13] ));
 sg13g2_dfrbp_1 _2155_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net386),
    .D(net441),
    .Q_N(_1047_),
    .Q(\CIC.int_1_out[14] ));
 sg13g2_dfrbp_1 _2156_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net387),
    .D(net307),
    .Q_N(_1048_),
    .Q(\CIC.int_1_out[15] ));
 sg13g2_dfrbp_1 _2157_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net386),
    .D(_0065_),
    .Q_N(_1049_),
    .Q(\CIC.int_1_out[16] ));
 sg13g2_dfrbp_1 _2158_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net382),
    .D(net414),
    .Q_N(_1050_),
    .Q(\CIC.int_1_out[17] ));
 sg13g2_dfrbp_1 _2159_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net382),
    .D(net450),
    .Q_N(_1051_),
    .Q(\CIC.int_1_out[18] ));
 sg13g2_dfrbp_1 _2160_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net382),
    .D(_0068_),
    .Q_N(_1052_),
    .Q(\CIC.int_1_out[19] ));
 sg13g2_dfrbp_1 _2161_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net381),
    .D(_0070_),
    .Q_N(_1053_),
    .Q(\CIC.int_1_out[20] ));
 sg13g2_dfrbp_1 _2162_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net381),
    .D(_0071_),
    .Q_N(_1054_),
    .Q(\CIC.int_1_out[21] ));
 sg13g2_dfrbp_1 _2163_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net381),
    .D(_0072_),
    .Q_N(_1055_),
    .Q(\CIC.int_1_out[22] ));
 sg13g2_dfrbp_1 _2164_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net383),
    .D(_0073_),
    .Q_N(_1056_),
    .Q(\CIC.int_1_out[23] ));
 sg13g2_dfrbp_1 _2165_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net412),
    .D(_0034_),
    .Q_N(_1057_),
    .Q(\CIC.inc_out[0] ));
 sg13g2_dfrbp_1 _2166_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net410),
    .D(_0045_),
    .Q_N(_1058_),
    .Q(\CIC.inc_out[1] ));
 sg13g2_dfrbp_1 _2167_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net410),
    .D(net169),
    .Q_N(_1059_),
    .Q(\CIC.inc_out[2] ));
 sg13g2_dfrbp_1 _2168_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net403),
    .D(_0051_),
    .Q_N(_1060_),
    .Q(\CIC.inc_out[3] ));
 sg13g2_dfrbp_1 _2169_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net402),
    .D(net118),
    .Q_N(_1061_),
    .Q(\CIC.inc_out[4] ));
 sg13g2_dfrbp_1 _2170_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net402),
    .D(net188),
    .Q_N(_1062_),
    .Q(\CIC.inc_out[5] ));
 sg13g2_dfrbp_1 _2171_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net402),
    .D(net161),
    .Q_N(_1063_),
    .Q(\CIC.inc_out[6] ));
 sg13g2_dfrbp_1 _2172_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net402),
    .D(_0055_),
    .Q_N(_1064_),
    .Q(\CIC.inc_out[7] ));
 sg13g2_dfrbp_1 _2173_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net402),
    .D(net207),
    .Q_N(_1065_),
    .Q(\CIC.inc_out[8] ));
 sg13g2_dfrbp_1 _2174_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net397),
    .D(_0057_),
    .Q_N(_1066_),
    .Q(\CIC.inc_out[9] ));
 sg13g2_dfrbp_1 _2175_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net397),
    .D(_0035_),
    .Q_N(_1067_),
    .Q(\CIC.inc_out[10] ));
 sg13g2_dfrbp_1 _2176_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net397),
    .D(net262),
    .Q_N(_1068_),
    .Q(\CIC.inc_out[11] ));
 sg13g2_dfrbp_1 _2177_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net397),
    .D(_0037_),
    .Q_N(_1069_),
    .Q(\CIC.inc_out[12] ));
 sg13g2_dfrbp_1 _2178_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net387),
    .D(_0038_),
    .Q_N(_1070_),
    .Q(\CIC.inc_out[13] ));
 sg13g2_dfrbp_1 _2179_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net386),
    .D(_0039_),
    .Q_N(_1071_),
    .Q(\CIC.inc_out[14] ));
 sg13g2_dfrbp_1 _2180_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net386),
    .D(net246),
    .Q_N(_1072_),
    .Q(\CIC.inc_out[15] ));
 sg13g2_dfrbp_1 _2181_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net386),
    .D(net248),
    .Q_N(_1073_),
    .Q(\CIC.inc_out[16] ));
 sg13g2_dfrbp_1 _2182_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net382),
    .D(_0042_),
    .Q_N(_1074_),
    .Q(\CIC.inc_out[17] ));
 sg13g2_dfrbp_1 _2183_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net382),
    .D(_0043_),
    .Q_N(_1075_),
    .Q(\CIC.inc_out[18] ));
 sg13g2_dfrbp_1 _2184_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net381),
    .D(net264),
    .Q_N(_1076_),
    .Q(\CIC.inc_out[19] ));
 sg13g2_dfrbp_1 _2185_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net381),
    .D(_0046_),
    .Q_N(_1077_),
    .Q(\CIC.inc_out[20] ));
 sg13g2_dfrbp_1 _2186_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net381),
    .D(net257),
    .Q_N(_1078_),
    .Q(\CIC.inc_out[21] ));
 sg13g2_dfrbp_1 _2187_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net381),
    .D(net251),
    .Q_N(_1079_),
    .Q(\CIC.inc_out[22] ));
 sg13g2_dfrbp_1 _2188_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net381),
    .D(net73),
    .Q_N(_0911_),
    .Q(\CIC.inc_out[23] ));
 sg13g2_dfrbp_1 _2189_ (.CLK(_0002_),
    .RESET_B(net395),
    .D(_0909_),
    .Q_N(_0909_),
    .Q(\outmux.count[0] ));
 sg13g2_dfrbp_1 _2190_ (.CLK(_0002_),
    .RESET_B(net395),
    .D(_0106_),
    .Q_N(_0910_),
    .Q(\outmux.count[1] ));
 sg13g2_dfrbp_1 _2191_ (.CLK(_0002_),
    .RESET_B(net395),
    .D(_0107_),
    .Q_N(_0010_),
    .Q(\outmux.count[2] ));
 sg13g2_tiehi _2064__15 (.L_HI(net15));
 sg13g2_tiehi _2063__16 (.L_HI(net16));
 sg13g2_tiehi _2062__17 (.L_HI(net17));
 sg13g2_tiehi _2061__18 (.L_HI(net18));
 sg13g2_tiehi _2060__19 (.L_HI(net19));
 sg13g2_tiehi _2059__20 (.L_HI(net20));
 sg13g2_tiehi _2058__21 (.L_HI(net21));
 sg13g2_tiehi _2057__22 (.L_HI(net22));
 sg13g2_tiehi _2056__23 (.L_HI(net23));
 sg13g2_tiehi _2055__24 (.L_HI(net24));
 sg13g2_tiehi _2054__25 (.L_HI(net25));
 sg13g2_tiehi _2053__26 (.L_HI(net26));
 sg13g2_tiehi _2052__27 (.L_HI(net27));
 sg13g2_tiehi _2051__28 (.L_HI(net28));
 sg13g2_tiehi _2050__29 (.L_HI(net29));
 sg13g2_tiehi _2049__30 (.L_HI(net30));
 sg13g2_tiehi _2048__31 (.L_HI(net31));
 sg13g2_tiehi _2047__32 (.L_HI(net32));
 sg13g2_tiehi _2046__33 (.L_HI(net33));
 sg13g2_tiehi _2045__34 (.L_HI(net34));
 sg13g2_tiehi _2044__35 (.L_HI(net35));
 sg13g2_tiehi _2043__36 (.L_HI(net36));
 sg13g2_tiehi _2042__37 (.L_HI(net37));
 sg13g2_tiehi tt_um_asheldon44_dsm_decimation_filter_38 (.L_HI(net38));
 sg13g2_tiehi tt_um_asheldon44_dsm_decimation_filter_39 (.L_HI(net39));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_asheldon44_dsm_decimation_filter_3 (.L_LO(net3));
 sg13g2_tielo tt_um_asheldon44_dsm_decimation_filter_4 (.L_LO(net4));
 sg13g2_tielo tt_um_asheldon44_dsm_decimation_filter_5 (.L_LO(net5));
 sg13g2_tielo tt_um_asheldon44_dsm_decimation_filter_6 (.L_LO(net6));
 sg13g2_tielo tt_um_asheldon44_dsm_decimation_filter_7 (.L_LO(net7));
 sg13g2_tielo tt_um_asheldon44_dsm_decimation_filter_8 (.L_LO(net8));
 sg13g2_tielo tt_um_asheldon44_dsm_decimation_filter_9 (.L_LO(net9));
 sg13g2_tielo tt_um_asheldon44_dsm_decimation_filter_10 (.L_LO(net10));
 sg13g2_tielo tt_um_asheldon44_dsm_decimation_filter_11 (.L_LO(net11));
 sg13g2_tielo tt_um_asheldon44_dsm_decimation_filter_12 (.L_LO(net12));
 sg13g2_tielo tt_um_asheldon44_dsm_decimation_filter_13 (.L_LO(net13));
 sg13g2_tiehi _2065__14 (.L_HI(net14));
 sg13g2_buf_1 _2230_ (.A(div_clk8x),
    .X(uio_out[0]));
 sg13g2_buf_1 _2231_ (.A(\CIC.dec_clk ),
    .X(uio_out[2]));
 sg13g2_buf_2 fanout309 (.A(net310),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(net316),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(net316),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(net315),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(net315),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(net315),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(net316),
    .X(net315));
 sg13g2_buf_1 fanout316 (.A(_0311_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(net320),
    .X(net317));
 sg13g2_buf_1 fanout318 (.A(net320),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(net320),
    .X(net319));
 sg13g2_buf_1 fanout320 (.A(_0395_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(net325),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(net324),
    .X(net322));
 sg13g2_buf_1 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_1 fanout324 (.A(net325),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_0395_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(net328),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(net328),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(net333),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(net330),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(net333),
    .X(net330));
 sg13g2_buf_1 fanout331 (.A(net333),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(net333),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_0309_),
    .X(net333));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(net338));
 sg13g2_buf_2 fanout335 (.A(net338),
    .X(net335));
 sg13g2_buf_4 fanout336 (.X(net336),
    .A(net338));
 sg13g2_buf_4 fanout337 (.X(net337),
    .A(net338));
 sg13g2_buf_2 fanout338 (.A(_0307_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(net342),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(net342),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(net342),
    .X(net341));
 sg13g2_buf_1 fanout342 (.A(net347),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(net345),
    .X(net343));
 sg13g2_buf_1 fanout344 (.A(net345),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(net346),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(net347),
    .X(net346));
 sg13g2_buf_1 fanout347 (.A(_0735_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(net349),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_0473_),
    .X(net349));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(net354));
 sg13g2_buf_2 fanout351 (.A(net354),
    .X(net351));
 sg13g2_buf_4 fanout352 (.X(net352),
    .A(net354));
 sg13g2_buf_2 fanout353 (.A(net354),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_0312_),
    .X(net354));
 sg13g2_buf_4 fanout355 (.X(net355),
    .A(net356));
 sg13g2_buf_2 fanout356 (.A(_0308_),
    .X(net356));
 sg13g2_buf_4 fanout357 (.X(net357),
    .A(net358));
 sg13g2_buf_2 fanout358 (.A(_0308_),
    .X(net358));
 sg13g2_buf_4 fanout359 (.X(net359),
    .A(_0734_));
 sg13g2_buf_2 fanout360 (.A(net361),
    .X(net360));
 sg13g2_buf_4 fanout361 (.X(net361),
    .A(_0733_));
 sg13g2_buf_4 fanout362 (.X(net362),
    .A(net363));
 sg13g2_buf_4 fanout363 (.X(net363),
    .A(_0740_));
 sg13g2_buf_4 fanout364 (.X(net364),
    .A(net365));
 sg13g2_buf_2 fanout365 (.A(_0738_),
    .X(net365));
 sg13g2_buf_4 fanout366 (.X(net366),
    .A(_0737_));
 sg13g2_buf_2 fanout367 (.A(_0737_),
    .X(net367));
 sg13g2_buf_4 fanout368 (.X(net368),
    .A(_0732_));
 sg13g2_buf_2 fanout369 (.A(_0732_),
    .X(net369));
 sg13g2_buf_4 fanout370 (.X(net370),
    .A(_0731_));
 sg13g2_buf_1 fanout371 (.A(_0731_),
    .X(net371));
 sg13g2_buf_4 fanout372 (.X(net372),
    .A(net374));
 sg13g2_buf_1 fanout373 (.A(net374),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(\CIC.u_differentiator.a_mux4to1.sel[1] ),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(net377),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(net377),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(net288),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(net379),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(net268),
    .X(net379));
 sg13g2_buf_4 fanout380 (.X(net380),
    .A(\CIC.u_differentiator.a_mux4to1.sel[0] ));
 sg13g2_buf_4 fanout381 (.X(net381),
    .A(net385));
 sg13g2_buf_4 fanout382 (.X(net382),
    .A(net385));
 sg13g2_buf_4 fanout383 (.X(net383),
    .A(net385));
 sg13g2_buf_4 fanout384 (.X(net384),
    .A(net385));
 sg13g2_buf_2 fanout385 (.A(net396),
    .X(net385));
 sg13g2_buf_4 fanout386 (.X(net386),
    .A(net389));
 sg13g2_buf_4 fanout387 (.X(net387),
    .A(net389));
 sg13g2_buf_4 fanout388 (.X(net388),
    .A(net389));
 sg13g2_buf_2 fanout389 (.A(net396),
    .X(net389));
 sg13g2_buf_4 fanout390 (.X(net390),
    .A(net391));
 sg13g2_buf_2 fanout391 (.A(net396),
    .X(net391));
 sg13g2_buf_4 fanout392 (.X(net392),
    .A(net393));
 sg13g2_buf_4 fanout393 (.X(net393),
    .A(net396));
 sg13g2_buf_4 fanout394 (.X(net394),
    .A(net395));
 sg13g2_buf_4 fanout395 (.X(net395),
    .A(net396));
 sg13g2_buf_2 fanout396 (.A(rst_n),
    .X(net396));
 sg13g2_buf_4 fanout397 (.X(net397),
    .A(net401));
 sg13g2_buf_2 fanout398 (.A(net401),
    .X(net398));
 sg13g2_buf_4 fanout399 (.X(net399),
    .A(net401));
 sg13g2_buf_4 fanout400 (.X(net400),
    .A(net401));
 sg13g2_buf_2 fanout401 (.A(net413),
    .X(net401));
 sg13g2_buf_4 fanout402 (.X(net402),
    .A(net405));
 sg13g2_buf_4 fanout403 (.X(net403),
    .A(net405));
 sg13g2_buf_2 fanout404 (.A(net405),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(net413),
    .X(net405));
 sg13g2_buf_4 fanout406 (.X(net406),
    .A(net407));
 sg13g2_buf_2 fanout407 (.A(net413),
    .X(net407));
 sg13g2_buf_4 fanout408 (.X(net408),
    .A(net412));
 sg13g2_buf_2 fanout409 (.A(net412),
    .X(net409));
 sg13g2_buf_4 fanout410 (.X(net410),
    .A(net411));
 sg13g2_buf_4 fanout411 (.X(net411),
    .A(net412));
 sg13g2_buf_2 fanout412 (.A(net413),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(rst_n),
    .X(net413));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_tielo tt_um_asheldon44_dsm_decimation_filter_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_25__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0000_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold2 (.A(\CIC.u_differentiator.a_mux4to1.d3[9] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold3 (.A(\CIC.u_differentiator.a_mux4to1.d3[13] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold4 (.A(\CIC.u_differentiator.a_mux4to1.d3[1] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0109_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold6 (.A(\CIC.u_differentiator.a_mux4to1.d2[15] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold7 (.A(\CIC.u_differentiator.a_mux4to1.d2[1] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0181_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold9 (.A(\CIC.u_differentiator.a_mux4to1.d3[15] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold10 (.A(\CIC.u_differentiator.a_mux4to1.d2[3] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold11 (.A(\CIC.u_differentiator.a_mux4to1.d2[5] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold12 (.A(\CIC.u_differentiator.a_mux4to1.d2[13] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold13 (.A(\CIC.u_differentiator.a_mux4to1.d2[9] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold14 (.A(\CIC.u_differentiator.a_mux4to1.d3[5] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold15 (.A(\CIC.u_differentiator.a_mux4to1.d3[3] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold16 (.A(\CIC.out[12] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold17 (.A(\CIC.out[11] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold18 (.A(\CIC.u_differentiator.a_mux4to1.d3[7] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold19 (.A(\CIC.out[8] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold20 (.A(\CIC.out[1] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0157_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold22 (.A(\CIC.out[15] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold23 (.A(\CIC.out[13] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold24 (.A(\CIC.out[10] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold25 (.A(\CIC.u_differentiator.a_mux4to1.d2[7] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold26 (.A(\CIC.out[9] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold27 (.A(\CIC.u_differentiator.a_mux4to1.d2[17] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold28 (.A(\CIC.out[6] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold29 (.A(\CIC.out[14] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold30 (.A(\CIC.out[16] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold31 (.A(\CIC.out[3] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold32 (.A(\CIC.out[21] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold33 (.A(\CIC.inc_out[23] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0049_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold35 (.A(\CIC.out[4] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold36 (.A(\CIC.u_differentiator.a_mux4to1.d2[11] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold37 (.A(\CIC.out[7] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold38 (.A(\CIC.u_differentiator.a_mux4to1.d2[19] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold39 (.A(\CIC.u_differentiator.a_mux4to1.d2[6] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold40 (.A(\CIC.out[19] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold41 (.A(\CIC.u_differentiator.a_mux4to1.d3[18] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold42 (.A(\CIC.u_differentiator.a_mux4to1.d3[8] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold43 (.A(\CIC.out[5] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold44 (.A(\CIC.out[17] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold45 (.A(\CIC.u_differentiator.temp[19] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0151_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold47 (.A(\CIC.u_differentiator.a_mux4to1.d3[12] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold48 (.A(\CIC.out[23] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold49 (.A(\CIC.u_differentiator.temp[17] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0149_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold51 (.A(\CIC.u_differentiator.a_mux4to1.d2[23] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold52 (.A(\CIC.u_differentiator.a_mux4to1.d2[14] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold53 (.A(\CIC.u_differentiator.a_mux4to1.d3[10] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold54 (.A(\CIC.int_2_out[0] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0082_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold56 (.A(\CIC.int_2_out[23] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0230_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold58 (.A(\CIC.u_differentiator.a_mux4to1.d3[16] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold59 (.A(\CIC.u_differentiator.a_mux4to1.d3[19] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold60 (.A(\CIC.u_differentiator.a_mux4to1.d3[20] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold61 (.A(\CIC.u_differentiator.a_mux4to1.d2[18] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold62 (.A(\CIC.u_differentiator.a_mux4to1.d3[22] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold63 (.A(\CIC.out[2] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold64 (.A(\CIC.u_differentiator.temp[1] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0133_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold66 (.A(\CIC.u_differentiator.a_mux4to1.d3[11] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold67 (.A(\CIC.u_differentiator.a_mux4to1.d2[8] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold68 (.A(\CIC.u_differentiator.temp[15] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0147_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold70 (.A(\CIC.u_differentiator.a_mux4to1.d2[4] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold71 (.A(\CIC.u_differentiator.a_mux4to1.d3[2] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold72 (.A(\CIC.out[20] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold73 (.A(\CIC.u_differentiator.a_mux4to1.d3[21] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold74 (.A(\CIC.out[0] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0156_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold76 (.A(\CIC.out[22] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold77 (.A(\CIC.inc_out[4] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0497_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0052_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold80 (.A(\CIC.u_differentiator.a_mux4to1.d3[0] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0108_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold82 (.A(\CIC.u_differentiator.a_mux4to1.d2[22] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold83 (.A(\CIC.u_differentiator.a_mux4to1.d3[6] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold84 (.A(\CIC.u_differentiator.a_mux4to1.d1[5] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0212_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold86 (.A(\CIC.u_differentiator.temp[23] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0155_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold88 (.A(\CIC.u_differentiator.a_mux4to1.d3[23] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold89 (.A(\CIC.u_differentiator.a_mux4to1.d2[20] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold90 (.A(\CIC.out[18] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold91 (.A(\CIC.u_differentiator.a_mux4to1.d2[21] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0022_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0354_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0143_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold95 (.A(\CIC.u_differentiator.a_mux4to1.d2[16] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold96 (.A(\CIC.u_differentiator.a_mux4to1.d2[10] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold97 (.A(\CIC.u_differentiator.a_mux4to1.d2[0] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0180_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold99 (.A(\CIC.inc_out[18] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0511_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold101 (.A(\CIC.int_2_out[6] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0213_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold103 (.A(\CIC.u_differentiator.a_mux4to1.d3[14] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold104 (.A(\CIC.u_differentiator.a_mux4to1.d1[1] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0208_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold106 (.A(\CIC.u_differentiator.temp[9] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0141_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0018_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0340_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0139_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold111 (.A(\CIC.int_2_out[19] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0226_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold113 (.A(\CIC.inc_out[10] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0503_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold115 (.A(\CIC.u_differentiator.a_mux4to1.d1[3] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0210_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold117 (.A(\CIC.u_differentiator.a_mux4to1.d3[17] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold118 (.A(\CIC.u_differentiator.a_mux4to1.d1[15] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0222_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold120 (.A(\CIC.inc_out[6] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0499_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0054_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold123 (.A(\CIC.u_differentiator.temp[3] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0135_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold125 (.A(\CIC.u_differentiator.a_mux4to1.d2[12] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold126 (.A(\CIC.u_differentiator.a_mux4to1.d3[4] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold127 (.A(\CIC.u_differentiator.a_mux4to1.d1[13] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0220_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold129 (.A(\CIC.inc_out[2] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0050_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold131 (.A(\CIC.int_1_out[0] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0058_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold133 (.A(\CIC.int_2_out[2] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0209_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold135 (.A(\CIC.inc_out[12] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0505_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold137 (.A(\CIC.u_differentiator.temp[0] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0132_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold139 (.A(\CIC.u_differentiator.a_mux4to1.d1[9] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0216_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold141 (.A(\CIC.u_differentiator.temp[16] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0148_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0009_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0447_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0206_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold146 (.A(\CIC.int_2_out[10] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0217_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold148 (.A(\CIC.inc_out[5] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0053_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold150 (.A(\CIC.u_differentiator.temp[6] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0138_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold152 (.A(\CIC.u_differentiator.temp[4] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0136_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold154 (.A(\CIC.u_differentiator.temp[10] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0142_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold156 (.A(\CIC.u_differentiator.temp[2] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0134_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold158 (.A(\CIC.int_2_out[8] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0215_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold160 (.A(\CIC.int_2_out[7] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0214_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold162 (.A(\CIC.u_differentiator.a_mux4to1.d2[2] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold163 (.A(\CIC.u_differentiator.temp[8] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0140_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold165 (.A(\CIC.u_differentiator.a_mux4to1.d1[0] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold166 (.A(\CIC.inc_out[8] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0501_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0056_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold169 (.A(\CIC.u_differentiator.temp[22] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0154_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold171 (.A(\CIC.u_differentiator.temp[12] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0144_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold173 (.A(\CIC.int_2_out[18] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0225_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold175 (.A(\CIC.int_2_out[21] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0228_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold177 (.A(\CIC.int_2_out[4] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0211_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold179 (.A(\CIC.u_differentiator.temp[13] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0145_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold181 (.A(\CIC.u_differentiator.temp[14] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0146_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold183 (.A(\CIC.u_differentiator.temp[18] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0150_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold185 (.A(\CIC.u_differentiator.temp[21] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0153_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold187 (.A(\CIC.int_2_out[14] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0221_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold189 (.A(\CIC.u_differentiator.a_mux4to1.d1[17] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0224_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold191 (.A(\CIC.u_differentiator.temp[5] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0137_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold193 (.A(\CIC.u_differentiator.a_mux4to1.d1[12] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0219_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold195 (.A(\CIC.int_2_out[22] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0229_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold197 (.A(\CIC.int_2_out[16] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0223_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold199 (.A(\CIC.inc_out[7] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold200 (.A(\CIC.u_differentiator.temp[20] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0152_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold202 (.A(\CIC.int_2_out[11] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0218_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold204 (.A(\CIC.int_2_out[20] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0227_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold206 (.A(\CIC.inc_out[15] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0040_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold208 (.A(\CIC.inc_out[16] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0041_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold210 (.A(\CIC.int_1_out[23] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold211 (.A(\CIC.inc_out[22] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0048_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold213 (.A(\CIC.inc_out[3] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold214 (.A(\CIC.inc_out[9] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold215 (.A(\CIC.inc_out[13] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold216 (.A(\CIC.inc_out[0] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold217 (.A(\CIC.inc_out[21] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0047_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold219 (.A(\CIC.inc_out[17] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold220 (.A(\CIC.int_2_out[1] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0519_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold222 (.A(\CIC.inc_out[11] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0036_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold224 (.A(\CIC.inc_out[19] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0044_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold226 (.A(\CIC.inc_out[22] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold227 (.A(\CIC.int_1_out[1] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0628_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold229 (.A(\CIC.u_differentiator.a_mux4to1.sel[0] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold230 (.A(\CIC.inc_out[14] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold231 (.A(\CIC.int_1_out[22] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0096_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold233 (.A(\CIC.int_2_out[3] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0525_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0099_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold236 (.A(\CIC.int_1_out[7] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold237 (.A(\CIC.int_1_out[8] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0081_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold239 (.A(\CIC.int_1_out[3] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0075_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold241 (.A(\CIC.int_2_out[5] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0530_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0101_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold244 (.A(\CIC.int_2_out[9] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0546_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold246 (.A(\CIC.int_2_out[7] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0538_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold248 (.A(\CIC.inc_out[20] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold249 (.A(\CIC.u_differentiator.a_mux4to1.sel[1] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold250 (.A(\CIC.int_1_out[18] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold251 (.A(\CIC.int_2_out[17] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0593_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold253 (.A(\CIC.int_1_out[10] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold254 (.A(\CIC.int_1_out[11] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0557_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold256 (.A(\CIC.int_1_out[6] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold257 (.A(\CIC.int_1_out[12] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0062_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold259 (.A(\CIC.int_1_out[4] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0077_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold261 (.A(\CIC.int_2_out[17] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold262 (.A(\CIC.inc_out[1] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold263 (.A(\CIC.inc_out[8] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0663_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0664_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold266 (.A(\CIC.int_1_out[14] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0690_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0064_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold269 (.A(\CIC.int_1_out[16] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0066_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold271 (.A(\CIC.int_1_out[19] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0708_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold273 (.A(\CIC.int_2_out[12] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0086_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold275 (.A(\CIC.int_1_out[20] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0095_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold277 (.A(\CIC.int_2_out[15] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0578_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold279 (.A(\CIC.int_1_out[2] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0098_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold281 (.A(\CIC.inc_out[7] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0651_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold283 (.A(\CIC.int_1_out[21] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold284 (.A(\CIC.inc_out[21] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0727_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold286 (.A(\CIC.int_2_out[13] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold287 (.A(\CIC.inc_out[3] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold288 (.A(\CIC.int_2_out[5] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0102_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold290 (.A(\CIC.int_2_out[16] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0583_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold292 (.A(\CIC.inc_out[9] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold293 (.A(\CIC.int_1_out[2] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold294 (.A(\CIC.inc_out[5] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0078_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold296 (.A(\CIC.inc_out[13] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0063_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold298 (.A(\CIC.inc_out[0] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0495_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold300 (.A(\CIC.inc_out[11] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold301 (.A(\CIC.inc_out[17] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold302 (.A(\CIC.int_1_out[22] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0728_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold304 (.A(\CIC.int_1_out[18] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0704_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0067_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold307 (.A(\CIC.int_1_out[22] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold308 (.A(\CIC.int_1_out[16] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0009_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold310 (.A(\CIC.int_1_out[6] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold311 (.A(\CIC.inc_out[18] ),
    .X(net455));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_4 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_163 ();
 sg13g2_decap_8 FILLER_0_170 ();
 sg13g2_decap_8 FILLER_0_177 ();
 sg13g2_decap_8 FILLER_0_184 ();
 sg13g2_decap_8 FILLER_0_191 ();
 sg13g2_decap_8 FILLER_0_198 ();
 sg13g2_decap_8 FILLER_0_205 ();
 sg13g2_decap_8 FILLER_0_212 ();
 sg13g2_decap_8 FILLER_0_219 ();
 sg13g2_decap_8 FILLER_0_226 ();
 sg13g2_decap_8 FILLER_0_233 ();
 sg13g2_decap_8 FILLER_0_240 ();
 sg13g2_decap_8 FILLER_0_247 ();
 sg13g2_decap_8 FILLER_0_254 ();
 sg13g2_decap_8 FILLER_0_261 ();
 sg13g2_decap_8 FILLER_0_268 ();
 sg13g2_decap_8 FILLER_0_275 ();
 sg13g2_decap_8 FILLER_0_282 ();
 sg13g2_decap_8 FILLER_0_289 ();
 sg13g2_decap_8 FILLER_0_296 ();
 sg13g2_decap_8 FILLER_0_303 ();
 sg13g2_decap_8 FILLER_0_310 ();
 sg13g2_decap_8 FILLER_0_317 ();
 sg13g2_decap_8 FILLER_0_324 ();
 sg13g2_decap_8 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_338 ();
 sg13g2_decap_8 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_fill_1 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_12 ();
 sg13g2_decap_8 FILLER_1_19 ();
 sg13g2_decap_8 FILLER_1_26 ();
 sg13g2_decap_8 FILLER_1_33 ();
 sg13g2_decap_8 FILLER_1_40 ();
 sg13g2_decap_8 FILLER_1_47 ();
 sg13g2_decap_8 FILLER_1_54 ();
 sg13g2_decap_8 FILLER_1_61 ();
 sg13g2_decap_8 FILLER_1_72 ();
 sg13g2_decap_4 FILLER_1_79 ();
 sg13g2_fill_1 FILLER_1_83 ();
 sg13g2_fill_2 FILLER_1_88 ();
 sg13g2_fill_1 FILLER_1_90 ();
 sg13g2_decap_4 FILLER_1_95 ();
 sg13g2_decap_8 FILLER_1_103 ();
 sg13g2_decap_4 FILLER_1_110 ();
 sg13g2_fill_1 FILLER_1_114 ();
 sg13g2_decap_8 FILLER_1_128 ();
 sg13g2_decap_4 FILLER_1_135 ();
 sg13g2_fill_2 FILLER_1_139 ();
 sg13g2_fill_1 FILLER_1_145 ();
 sg13g2_decap_8 FILLER_1_179 ();
 sg13g2_decap_4 FILLER_1_186 ();
 sg13g2_decap_8 FILLER_1_194 ();
 sg13g2_fill_2 FILLER_1_201 ();
 sg13g2_decap_8 FILLER_1_207 ();
 sg13g2_decap_8 FILLER_1_214 ();
 sg13g2_decap_8 FILLER_1_221 ();
 sg13g2_decap_8 FILLER_1_228 ();
 sg13g2_decap_8 FILLER_1_235 ();
 sg13g2_decap_8 FILLER_1_242 ();
 sg13g2_decap_8 FILLER_1_249 ();
 sg13g2_fill_1 FILLER_1_256 ();
 sg13g2_decap_8 FILLER_1_261 ();
 sg13g2_decap_8 FILLER_1_268 ();
 sg13g2_fill_2 FILLER_1_275 ();
 sg13g2_decap_8 FILLER_1_282 ();
 sg13g2_decap_8 FILLER_1_289 ();
 sg13g2_fill_1 FILLER_1_296 ();
 sg13g2_fill_2 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_307 ();
 sg13g2_decap_8 FILLER_1_314 ();
 sg13g2_decap_8 FILLER_1_321 ();
 sg13g2_decap_8 FILLER_1_328 ();
 sg13g2_decap_8 FILLER_1_335 ();
 sg13g2_decap_8 FILLER_1_342 ();
 sg13g2_decap_4 FILLER_1_349 ();
 sg13g2_fill_2 FILLER_1_353 ();
 sg13g2_decap_8 FILLER_1_359 ();
 sg13g2_decap_8 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_373 ();
 sg13g2_decap_8 FILLER_1_380 ();
 sg13g2_decap_8 FILLER_1_387 ();
 sg13g2_decap_8 FILLER_1_394 ();
 sg13g2_decap_8 FILLER_1_401 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_30 ();
 sg13g2_decap_4 FILLER_2_55 ();
 sg13g2_fill_1 FILLER_2_59 ();
 sg13g2_fill_2 FILLER_2_84 ();
 sg13g2_fill_1 FILLER_2_91 ();
 sg13g2_fill_1 FILLER_2_139 ();
 sg13g2_decap_8 FILLER_2_242 ();
 sg13g2_fill_2 FILLER_2_284 ();
 sg13g2_fill_2 FILLER_2_306 ();
 sg13g2_fill_1 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_316 ();
 sg13g2_decap_8 FILLER_2_323 ();
 sg13g2_decap_8 FILLER_2_330 ();
 sg13g2_decap_4 FILLER_2_337 ();
 sg13g2_fill_1 FILLER_2_341 ();
 sg13g2_fill_2 FILLER_2_347 ();
 sg13g2_fill_1 FILLER_2_349 ();
 sg13g2_fill_2 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_372 ();
 sg13g2_decap_8 FILLER_2_379 ();
 sg13g2_decap_8 FILLER_2_386 ();
 sg13g2_decap_8 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_400 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_fill_2 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_42 ();
 sg13g2_fill_1 FILLER_3_57 ();
 sg13g2_fill_1 FILLER_3_72 ();
 sg13g2_fill_1 FILLER_3_158 ();
 sg13g2_fill_1 FILLER_3_164 ();
 sg13g2_fill_1 FILLER_3_190 ();
 sg13g2_fill_2 FILLER_3_209 ();
 sg13g2_fill_2 FILLER_3_267 ();
 sg13g2_fill_2 FILLER_3_316 ();
 sg13g2_fill_1 FILLER_3_318 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_4 FILLER_3_403 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_fill_2 FILLER_4_103 ();
 sg13g2_fill_1 FILLER_4_105 ();
 sg13g2_fill_2 FILLER_4_132 ();
 sg13g2_fill_1 FILLER_4_169 ();
 sg13g2_fill_1 FILLER_4_197 ();
 sg13g2_fill_2 FILLER_4_204 ();
 sg13g2_fill_1 FILLER_4_218 ();
 sg13g2_fill_2 FILLER_4_228 ();
 sg13g2_fill_1 FILLER_4_230 ();
 sg13g2_fill_2 FILLER_4_249 ();
 sg13g2_fill_2 FILLER_4_260 ();
 sg13g2_fill_1 FILLER_4_302 ();
 sg13g2_fill_2 FILLER_4_355 ();
 sg13g2_decap_4 FILLER_4_405 ();
 sg13g2_fill_1 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_18 ();
 sg13g2_fill_2 FILLER_5_37 ();
 sg13g2_fill_1 FILLER_5_141 ();
 sg13g2_fill_2 FILLER_5_151 ();
 sg13g2_fill_1 FILLER_5_199 ();
 sg13g2_fill_1 FILLER_5_205 ();
 sg13g2_fill_1 FILLER_5_227 ();
 sg13g2_fill_2 FILLER_5_250 ();
 sg13g2_fill_1 FILLER_5_265 ();
 sg13g2_fill_1 FILLER_5_320 ();
 sg13g2_fill_2 FILLER_5_348 ();
 sg13g2_fill_1 FILLER_5_364 ();
 sg13g2_fill_2 FILLER_5_396 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_fill_1 FILLER_6_8 ();
 sg13g2_fill_1 FILLER_6_89 ();
 sg13g2_fill_2 FILLER_6_117 ();
 sg13g2_fill_1 FILLER_6_119 ();
 sg13g2_fill_2 FILLER_6_192 ();
 sg13g2_fill_2 FILLER_6_240 ();
 sg13g2_fill_1 FILLER_6_250 ();
 sg13g2_fill_1 FILLER_6_264 ();
 sg13g2_fill_1 FILLER_6_355 ();
 sg13g2_fill_2 FILLER_7_108 ();
 sg13g2_fill_2 FILLER_7_153 ();
 sg13g2_fill_2 FILLER_7_189 ();
 sg13g2_fill_2 FILLER_7_228 ();
 sg13g2_fill_2 FILLER_7_247 ();
 sg13g2_fill_1 FILLER_7_286 ();
 sg13g2_fill_1 FILLER_7_316 ();
 sg13g2_fill_2 FILLER_7_339 ();
 sg13g2_fill_1 FILLER_7_363 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_fill_1 FILLER_8_40 ();
 sg13g2_fill_1 FILLER_8_57 ();
 sg13g2_fill_1 FILLER_8_72 ();
 sg13g2_fill_1 FILLER_8_156 ();
 sg13g2_fill_2 FILLER_8_178 ();
 sg13g2_fill_1 FILLER_8_193 ();
 sg13g2_fill_1 FILLER_8_214 ();
 sg13g2_fill_1 FILLER_8_281 ();
 sg13g2_fill_2 FILLER_8_290 ();
 sg13g2_fill_2 FILLER_8_323 ();
 sg13g2_fill_2 FILLER_8_368 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_71 ();
 sg13g2_fill_1 FILLER_9_80 ();
 sg13g2_fill_2 FILLER_9_95 ();
 sg13g2_fill_1 FILLER_9_121 ();
 sg13g2_fill_1 FILLER_9_145 ();
 sg13g2_fill_1 FILLER_9_208 ();
 sg13g2_fill_1 FILLER_9_222 ();
 sg13g2_decap_4 FILLER_9_228 ();
 sg13g2_fill_1 FILLER_9_232 ();
 sg13g2_fill_2 FILLER_9_247 ();
 sg13g2_fill_1 FILLER_9_249 ();
 sg13g2_fill_2 FILLER_9_269 ();
 sg13g2_fill_1 FILLER_9_271 ();
 sg13g2_fill_1 FILLER_9_277 ();
 sg13g2_fill_2 FILLER_9_347 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_71 ();
 sg13g2_fill_1 FILLER_10_82 ();
 sg13g2_fill_1 FILLER_10_156 ();
 sg13g2_fill_1 FILLER_10_183 ();
 sg13g2_fill_1 FILLER_10_193 ();
 sg13g2_fill_2 FILLER_10_222 ();
 sg13g2_fill_1 FILLER_10_233 ();
 sg13g2_decap_4 FILLER_10_254 ();
 sg13g2_fill_2 FILLER_10_258 ();
 sg13g2_fill_2 FILLER_10_280 ();
 sg13g2_fill_2 FILLER_10_304 ();
 sg13g2_fill_1 FILLER_10_306 ();
 sg13g2_fill_1 FILLER_11_35 ();
 sg13g2_fill_2 FILLER_11_62 ();
 sg13g2_fill_2 FILLER_11_80 ();
 sg13g2_fill_2 FILLER_11_92 ();
 sg13g2_fill_1 FILLER_11_104 ();
 sg13g2_fill_1 FILLER_11_156 ();
 sg13g2_fill_1 FILLER_11_192 ();
 sg13g2_decap_8 FILLER_11_248 ();
 sg13g2_fill_2 FILLER_11_255 ();
 sg13g2_fill_1 FILLER_11_257 ();
 sg13g2_fill_1 FILLER_11_266 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_35 ();
 sg13g2_fill_1 FILLER_12_53 ();
 sg13g2_fill_1 FILLER_12_92 ();
 sg13g2_fill_2 FILLER_12_177 ();
 sg13g2_fill_1 FILLER_12_179 ();
 sg13g2_fill_2 FILLER_12_212 ();
 sg13g2_fill_1 FILLER_12_214 ();
 sg13g2_fill_2 FILLER_12_283 ();
 sg13g2_fill_2 FILLER_12_294 ();
 sg13g2_fill_1 FILLER_12_296 ();
 sg13g2_fill_2 FILLER_12_337 ();
 sg13g2_fill_1 FILLER_12_373 ();
 sg13g2_fill_2 FILLER_13_30 ();
 sg13g2_fill_1 FILLER_13_32 ();
 sg13g2_fill_2 FILLER_13_42 ();
 sg13g2_fill_1 FILLER_13_44 ();
 sg13g2_fill_1 FILLER_13_83 ();
 sg13g2_fill_1 FILLER_13_129 ();
 sg13g2_fill_1 FILLER_13_135 ();
 sg13g2_fill_2 FILLER_13_140 ();
 sg13g2_fill_1 FILLER_13_182 ();
 sg13g2_fill_1 FILLER_13_198 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_fill_2 FILLER_13_259 ();
 sg13g2_fill_2 FILLER_13_346 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_43 ();
 sg13g2_fill_2 FILLER_14_109 ();
 sg13g2_fill_2 FILLER_14_192 ();
 sg13g2_fill_1 FILLER_14_194 ();
 sg13g2_fill_2 FILLER_14_218 ();
 sg13g2_fill_1 FILLER_14_220 ();
 sg13g2_decap_4 FILLER_14_247 ();
 sg13g2_fill_2 FILLER_14_251 ();
 sg13g2_fill_1 FILLER_14_307 ();
 sg13g2_fill_2 FILLER_15_83 ();
 sg13g2_fill_2 FILLER_15_109 ();
 sg13g2_fill_2 FILLER_15_128 ();
 sg13g2_fill_1 FILLER_15_130 ();
 sg13g2_fill_2 FILLER_15_184 ();
 sg13g2_fill_2 FILLER_15_212 ();
 sg13g2_fill_2 FILLER_15_251 ();
 sg13g2_fill_1 FILLER_15_253 ();
 sg13g2_fill_1 FILLER_15_310 ();
 sg13g2_fill_1 FILLER_15_341 ();
 sg13g2_fill_2 FILLER_15_383 ();
 sg13g2_fill_1 FILLER_15_399 ();
 sg13g2_fill_1 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_18 ();
 sg13g2_fill_1 FILLER_16_20 ();
 sg13g2_fill_2 FILLER_16_54 ();
 sg13g2_fill_2 FILLER_16_119 ();
 sg13g2_fill_1 FILLER_16_121 ();
 sg13g2_fill_1 FILLER_16_155 ();
 sg13g2_fill_2 FILLER_16_165 ();
 sg13g2_fill_2 FILLER_16_205 ();
 sg13g2_fill_2 FILLER_16_269 ();
 sg13g2_fill_1 FILLER_16_271 ();
 sg13g2_fill_2 FILLER_16_291 ();
 sg13g2_fill_2 FILLER_16_302 ();
 sg13g2_fill_1 FILLER_16_361 ();
 sg13g2_fill_2 FILLER_17_30 ();
 sg13g2_fill_2 FILLER_17_136 ();
 sg13g2_fill_1 FILLER_17_138 ();
 sg13g2_fill_1 FILLER_17_144 ();
 sg13g2_fill_1 FILLER_17_217 ();
 sg13g2_fill_2 FILLER_17_278 ();
 sg13g2_fill_2 FILLER_17_325 ();
 sg13g2_fill_1 FILLER_17_341 ();
 sg13g2_fill_1 FILLER_17_356 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_2 ();
 sg13g2_fill_1 FILLER_18_20 ();
 sg13g2_decap_4 FILLER_18_40 ();
 sg13g2_fill_2 FILLER_18_58 ();
 sg13g2_fill_1 FILLER_18_60 ();
 sg13g2_fill_2 FILLER_18_110 ();
 sg13g2_fill_1 FILLER_18_112 ();
 sg13g2_fill_2 FILLER_18_173 ();
 sg13g2_fill_2 FILLER_18_204 ();
 sg13g2_fill_1 FILLER_18_206 ();
 sg13g2_decap_4 FILLER_18_216 ();
 sg13g2_fill_1 FILLER_18_220 ();
 sg13g2_fill_2 FILLER_18_226 ();
 sg13g2_decap_4 FILLER_18_232 ();
 sg13g2_fill_1 FILLER_18_236 ();
 sg13g2_fill_2 FILLER_18_256 ();
 sg13g2_fill_2 FILLER_18_313 ();
 sg13g2_fill_2 FILLER_18_328 ();
 sg13g2_fill_2 FILLER_18_340 ();
 sg13g2_fill_2 FILLER_19_26 ();
 sg13g2_fill_1 FILLER_19_28 ();
 sg13g2_decap_4 FILLER_19_77 ();
 sg13g2_decap_4 FILLER_19_115 ();
 sg13g2_fill_2 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_232 ();
 sg13g2_fill_2 FILLER_19_240 ();
 sg13g2_fill_1 FILLER_19_293 ();
 sg13g2_fill_2 FILLER_19_303 ();
 sg13g2_fill_1 FILLER_19_332 ();
 sg13g2_fill_1 FILLER_19_358 ();
 sg13g2_fill_2 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_33 ();
 sg13g2_fill_1 FILLER_20_59 ();
 sg13g2_fill_2 FILLER_20_63 ();
 sg13g2_fill_2 FILLER_20_91 ();
 sg13g2_fill_1 FILLER_20_93 ();
 sg13g2_fill_2 FILLER_20_103 ();
 sg13g2_fill_2 FILLER_20_131 ();
 sg13g2_fill_2 FILLER_20_142 ();
 sg13g2_fill_1 FILLER_20_144 ();
 sg13g2_fill_1 FILLER_20_162 ();
 sg13g2_decap_4 FILLER_20_177 ();
 sg13g2_fill_2 FILLER_20_181 ();
 sg13g2_decap_8 FILLER_20_193 ();
 sg13g2_decap_4 FILLER_20_200 ();
 sg13g2_fill_1 FILLER_20_222 ();
 sg13g2_fill_2 FILLER_20_230 ();
 sg13g2_fill_1 FILLER_20_232 ();
 sg13g2_fill_1 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_251 ();
 sg13g2_decap_4 FILLER_20_258 ();
 sg13g2_fill_2 FILLER_20_271 ();
 sg13g2_fill_1 FILLER_20_273 ();
 sg13g2_fill_1 FILLER_20_367 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_4 ();
 sg13g2_fill_2 FILLER_21_32 ();
 sg13g2_fill_2 FILLER_21_43 ();
 sg13g2_decap_4 FILLER_21_81 ();
 sg13g2_fill_1 FILLER_21_94 ();
 sg13g2_decap_8 FILLER_21_113 ();
 sg13g2_decap_4 FILLER_21_120 ();
 sg13g2_fill_1 FILLER_21_138 ();
 sg13g2_decap_8 FILLER_21_149 ();
 sg13g2_decap_4 FILLER_21_156 ();
 sg13g2_decap_4 FILLER_21_176 ();
 sg13g2_decap_8 FILLER_21_239 ();
 sg13g2_fill_1 FILLER_21_246 ();
 sg13g2_decap_4 FILLER_21_252 ();
 sg13g2_fill_2 FILLER_21_256 ();
 sg13g2_fill_2 FILLER_21_293 ();
 sg13g2_fill_2 FILLER_21_309 ();
 sg13g2_fill_1 FILLER_21_311 ();
 sg13g2_fill_1 FILLER_21_321 ();
 sg13g2_fill_1 FILLER_21_377 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_4 ();
 sg13g2_fill_2 FILLER_22_31 ();
 sg13g2_fill_1 FILLER_22_33 ();
 sg13g2_fill_2 FILLER_22_78 ();
 sg13g2_fill_1 FILLER_22_80 ();
 sg13g2_decap_4 FILLER_22_86 ();
 sg13g2_fill_1 FILLER_22_90 ();
 sg13g2_fill_1 FILLER_22_103 ();
 sg13g2_decap_8 FILLER_22_113 ();
 sg13g2_fill_1 FILLER_22_120 ();
 sg13g2_fill_2 FILLER_22_164 ();
 sg13g2_decap_8 FILLER_22_174 ();
 sg13g2_fill_1 FILLER_22_202 ();
 sg13g2_decap_8 FILLER_22_208 ();
 sg13g2_decap_4 FILLER_22_215 ();
 sg13g2_fill_2 FILLER_22_272 ();
 sg13g2_fill_2 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_11 ();
 sg13g2_decap_4 FILLER_23_91 ();
 sg13g2_fill_1 FILLER_23_95 ();
 sg13g2_fill_1 FILLER_23_104 ();
 sg13g2_fill_2 FILLER_23_123 ();
 sg13g2_fill_1 FILLER_23_155 ();
 sg13g2_fill_1 FILLER_23_197 ();
 sg13g2_fill_2 FILLER_23_292 ();
 sg13g2_fill_1 FILLER_23_351 ();
 sg13g2_fill_2 FILLER_23_361 ();
 sg13g2_fill_2 FILLER_23_381 ();
 sg13g2_fill_2 FILLER_24_26 ();
 sg13g2_fill_2 FILLER_24_37 ();
 sg13g2_fill_1 FILLER_24_39 ();
 sg13g2_fill_1 FILLER_24_68 ();
 sg13g2_fill_2 FILLER_24_83 ();
 sg13g2_decap_4 FILLER_24_101 ();
 sg13g2_fill_1 FILLER_24_125 ();
 sg13g2_fill_1 FILLER_24_173 ();
 sg13g2_fill_1 FILLER_24_185 ();
 sg13g2_decap_4 FILLER_24_194 ();
 sg13g2_fill_1 FILLER_24_198 ();
 sg13g2_fill_1 FILLER_24_207 ();
 sg13g2_decap_4 FILLER_24_217 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_fill_1 FILLER_24_231 ();
 sg13g2_fill_2 FILLER_24_258 ();
 sg13g2_fill_1 FILLER_24_274 ();
 sg13g2_fill_2 FILLER_24_321 ();
 sg13g2_fill_1 FILLER_24_328 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_fill_1 FILLER_25_43 ();
 sg13g2_fill_2 FILLER_25_54 ();
 sg13g2_fill_1 FILLER_25_56 ();
 sg13g2_fill_1 FILLER_25_83 ();
 sg13g2_fill_2 FILLER_25_184 ();
 sg13g2_fill_1 FILLER_25_186 ();
 sg13g2_fill_2 FILLER_25_200 ();
 sg13g2_fill_1 FILLER_25_253 ();
 sg13g2_fill_2 FILLER_25_317 ();
 sg13g2_fill_1 FILLER_25_319 ();
 sg13g2_fill_1 FILLER_25_336 ();
 sg13g2_fill_2 FILLER_25_345 ();
 sg13g2_fill_1 FILLER_25_367 ();
 sg13g2_fill_1 FILLER_25_373 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_69 ();
 sg13g2_fill_1 FILLER_26_71 ();
 sg13g2_decap_8 FILLER_26_86 ();
 sg13g2_fill_2 FILLER_26_107 ();
 sg13g2_fill_2 FILLER_26_127 ();
 sg13g2_fill_1 FILLER_26_129 ();
 sg13g2_fill_2 FILLER_26_142 ();
 sg13g2_fill_1 FILLER_26_144 ();
 sg13g2_fill_1 FILLER_26_154 ();
 sg13g2_fill_1 FILLER_26_169 ();
 sg13g2_decap_4 FILLER_26_193 ();
 sg13g2_fill_1 FILLER_26_197 ();
 sg13g2_fill_1 FILLER_26_224 ();
 sg13g2_fill_1 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_266 ();
 sg13g2_fill_1 FILLER_26_268 ();
 sg13g2_fill_2 FILLER_26_273 ();
 sg13g2_fill_1 FILLER_26_318 ();
 sg13g2_fill_1 FILLER_26_339 ();
 sg13g2_fill_2 FILLER_26_345 ();
 sg13g2_fill_1 FILLER_26_373 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_fill_1 FILLER_27_49 ();
 sg13g2_fill_2 FILLER_27_65 ();
 sg13g2_fill_1 FILLER_27_67 ();
 sg13g2_fill_2 FILLER_27_83 ();
 sg13g2_fill_2 FILLER_27_117 ();
 sg13g2_fill_1 FILLER_27_119 ();
 sg13g2_fill_2 FILLER_27_128 ();
 sg13g2_decap_8 FILLER_27_205 ();
 sg13g2_fill_2 FILLER_27_217 ();
 sg13g2_fill_1 FILLER_27_238 ();
 sg13g2_fill_2 FILLER_27_247 ();
 sg13g2_fill_2 FILLER_27_254 ();
 sg13g2_fill_1 FILLER_27_256 ();
 sg13g2_fill_1 FILLER_27_290 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_52 ();
 sg13g2_fill_1 FILLER_28_67 ();
 sg13g2_fill_2 FILLER_28_73 ();
 sg13g2_fill_1 FILLER_28_75 ();
 sg13g2_decap_4 FILLER_28_88 ();
 sg13g2_fill_2 FILLER_28_92 ();
 sg13g2_decap_8 FILLER_28_99 ();
 sg13g2_fill_2 FILLER_28_146 ();
 sg13g2_fill_2 FILLER_28_176 ();
 sg13g2_fill_2 FILLER_28_201 ();
 sg13g2_fill_1 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_209 ();
 sg13g2_fill_2 FILLER_28_216 ();
 sg13g2_fill_2 FILLER_28_248 ();
 sg13g2_fill_2 FILLER_28_272 ();
 sg13g2_fill_1 FILLER_28_278 ();
 sg13g2_fill_2 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_56 ();
 sg13g2_fill_1 FILLER_29_67 ();
 sg13g2_decap_8 FILLER_29_82 ();
 sg13g2_fill_1 FILLER_29_98 ();
 sg13g2_fill_1 FILLER_29_116 ();
 sg13g2_fill_2 FILLER_29_131 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_fill_1 FILLER_29_158 ();
 sg13g2_fill_1 FILLER_29_196 ();
 sg13g2_fill_1 FILLER_29_202 ();
 sg13g2_fill_2 FILLER_29_229 ();
 sg13g2_fill_1 FILLER_29_231 ();
 sg13g2_fill_2 FILLER_29_272 ();
 sg13g2_fill_1 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_280 ();
 sg13g2_fill_2 FILLER_29_350 ();
 sg13g2_fill_1 FILLER_29_352 ();
 sg13g2_fill_1 FILLER_29_362 ();
 sg13g2_fill_2 FILLER_29_380 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_4 ();
 sg13g2_fill_2 FILLER_30_23 ();
 sg13g2_fill_2 FILLER_30_59 ();
 sg13g2_decap_4 FILLER_30_103 ();
 sg13g2_fill_1 FILLER_30_107 ();
 sg13g2_fill_1 FILLER_30_139 ();
 sg13g2_fill_2 FILLER_30_166 ();
 sg13g2_fill_2 FILLER_30_194 ();
 sg13g2_fill_1 FILLER_30_209 ();
 sg13g2_fill_1 FILLER_30_219 ();
 sg13g2_fill_2 FILLER_30_242 ();
 sg13g2_fill_2 FILLER_30_335 ();
 sg13g2_fill_2 FILLER_30_342 ();
 sg13g2_fill_1 FILLER_30_344 ();
 sg13g2_fill_2 FILLER_30_362 ();
 sg13g2_fill_1 FILLER_31_26 ();
 sg13g2_fill_2 FILLER_31_90 ();
 sg13g2_fill_1 FILLER_31_92 ();
 sg13g2_decap_8 FILLER_31_132 ();
 sg13g2_fill_1 FILLER_31_139 ();
 sg13g2_fill_1 FILLER_31_148 ();
 sg13g2_fill_2 FILLER_31_171 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_fill_2 FILLER_31_262 ();
 sg13g2_fill_1 FILLER_31_264 ();
 sg13g2_fill_1 FILLER_31_270 ();
 sg13g2_fill_1 FILLER_31_280 ();
 sg13g2_fill_1 FILLER_31_323 ();
 sg13g2_fill_2 FILLER_32_26 ();
 sg13g2_fill_2 FILLER_32_62 ();
 sg13g2_fill_1 FILLER_32_77 ();
 sg13g2_decap_4 FILLER_32_104 ();
 sg13g2_fill_1 FILLER_32_108 ();
 sg13g2_fill_2 FILLER_32_113 ();
 sg13g2_fill_1 FILLER_32_115 ();
 sg13g2_fill_2 FILLER_32_121 ();
 sg13g2_fill_2 FILLER_32_136 ();
 sg13g2_fill_1 FILLER_32_138 ();
 sg13g2_fill_1 FILLER_32_155 ();
 sg13g2_fill_2 FILLER_32_165 ();
 sg13g2_fill_1 FILLER_32_167 ();
 sg13g2_fill_1 FILLER_32_219 ();
 sg13g2_fill_2 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_234 ();
 sg13g2_fill_2 FILLER_32_356 ();
 sg13g2_fill_1 FILLER_32_399 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_90 ();
 sg13g2_decap_8 FILLER_33_100 ();
 sg13g2_decap_4 FILLER_33_107 ();
 sg13g2_fill_1 FILLER_33_142 ();
 sg13g2_fill_2 FILLER_33_173 ();
 sg13g2_fill_1 FILLER_33_175 ();
 sg13g2_fill_2 FILLER_33_185 ();
 sg13g2_fill_1 FILLER_33_204 ();
 sg13g2_fill_1 FILLER_33_209 ();
 sg13g2_fill_1 FILLER_33_215 ();
 sg13g2_fill_1 FILLER_33_220 ();
 sg13g2_fill_1 FILLER_33_243 ();
 sg13g2_fill_1 FILLER_33_265 ();
 sg13g2_fill_1 FILLER_33_347 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_fill_2 FILLER_34_35 ();
 sg13g2_fill_2 FILLER_34_59 ();
 sg13g2_fill_1 FILLER_34_61 ();
 sg13g2_fill_2 FILLER_34_81 ();
 sg13g2_fill_1 FILLER_34_163 ();
 sg13g2_fill_2 FILLER_34_184 ();
 sg13g2_fill_1 FILLER_34_186 ();
 sg13g2_fill_2 FILLER_34_204 ();
 sg13g2_fill_2 FILLER_34_232 ();
 sg13g2_fill_1 FILLER_34_234 ();
 sg13g2_fill_1 FILLER_34_341 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_fill_2 FILLER_35_26 ();
 sg13g2_fill_2 FILLER_35_106 ();
 sg13g2_fill_1 FILLER_35_108 ();
 sg13g2_fill_1 FILLER_35_127 ();
 sg13g2_fill_2 FILLER_35_208 ();
 sg13g2_fill_2 FILLER_35_222 ();
 sg13g2_fill_1 FILLER_35_224 ();
 sg13g2_fill_2 FILLER_35_231 ();
 sg13g2_fill_1 FILLER_35_233 ();
 sg13g2_fill_2 FILLER_35_260 ();
 sg13g2_fill_1 FILLER_35_262 ();
 sg13g2_fill_1 FILLER_35_289 ();
 sg13g2_fill_2 FILLER_35_334 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_56 ();
 sg13g2_fill_1 FILLER_36_58 ();
 sg13g2_fill_1 FILLER_36_90 ();
 sg13g2_fill_2 FILLER_36_116 ();
 sg13g2_fill_2 FILLER_36_126 ();
 sg13g2_fill_2 FILLER_36_190 ();
 sg13g2_fill_2 FILLER_36_201 ();
 sg13g2_fill_2 FILLER_36_248 ();
 sg13g2_fill_1 FILLER_36_250 ();
 sg13g2_fill_2 FILLER_36_262 ();
 sg13g2_fill_1 FILLER_36_278 ();
 sg13g2_fill_1 FILLER_36_384 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_24 ();
 sg13g2_decap_4 FILLER_37_31 ();
 sg13g2_fill_2 FILLER_37_39 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_fill_2 FILLER_37_337 ();
 sg13g2_fill_1 FILLER_37_339 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_49 ();
 sg13g2_fill_2 FILLER_38_54 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_fill_2 FILLER_38_76 ();
 sg13g2_fill_1 FILLER_38_78 ();
 sg13g2_fill_2 FILLER_38_178 ();
 sg13g2_fill_2 FILLER_38_184 ();
 sg13g2_fill_1 FILLER_38_198 ();
 sg13g2_fill_2 FILLER_38_229 ();
 sg13g2_fill_2 FILLER_38_248 ();
 sg13g2_fill_1 FILLER_38_265 ();
 sg13g2_fill_1 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_fill_1 FILLER_38_372 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net38;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net39;
 assign uio_oe[3] = net3;
 assign uio_oe[4] = net4;
 assign uio_oe[5] = net5;
 assign uio_oe[6] = net6;
 assign uio_oe[7] = net7;
 assign uio_out[1] = net8;
 assign uio_out[3] = net9;
 assign uio_out[4] = net10;
 assign uio_out[5] = net11;
 assign uio_out[6] = net12;
 assign uio_out[7] = net13;
endmodule

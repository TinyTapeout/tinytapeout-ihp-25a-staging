module tt_um_16_mic_beamformer_arghunter (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire out;
 wire \u_top_module.u_cic.inc_out[10] ;
 wire \u_top_module.u_cic.inc_out[11] ;
 wire \u_top_module.u_cic.inc_out[12] ;
 wire \u_top_module.u_cic.inc_out[13] ;
 wire \u_top_module.u_cic.inc_out[14] ;
 wire \u_top_module.u_cic.inc_out[15] ;
 wire \u_top_module.u_cic.inc_out[16] ;
 wire \u_top_module.u_cic.inc_out[17] ;
 wire \u_top_module.u_cic.inc_out[18] ;
 wire \u_top_module.u_cic.inc_out[19] ;
 wire \u_top_module.u_cic.inc_out[1] ;
 wire \u_top_module.u_cic.inc_out[20] ;
 wire \u_top_module.u_cic.inc_out[21] ;
 wire \u_top_module.u_cic.inc_out[22] ;
 wire \u_top_module.u_cic.inc_out[23] ;
 wire \u_top_module.u_cic.inc_out[2] ;
 wire \u_top_module.u_cic.inc_out[3] ;
 wire \u_top_module.u_cic.inc_out[4] ;
 wire \u_top_module.u_cic.inc_out[5] ;
 wire \u_top_module.u_cic.inc_out[6] ;
 wire \u_top_module.u_cic.inc_out[7] ;
 wire \u_top_module.u_cic.inc_out[8] ;
 wire \u_top_module.u_cic.inc_out[9] ;
 wire \u_top_module.u_cic.int_1_out[10] ;
 wire \u_top_module.u_cic.int_1_out[11] ;
 wire \u_top_module.u_cic.int_1_out[12] ;
 wire \u_top_module.u_cic.int_1_out[13] ;
 wire \u_top_module.u_cic.int_1_out[14] ;
 wire \u_top_module.u_cic.int_1_out[15] ;
 wire \u_top_module.u_cic.int_1_out[16] ;
 wire \u_top_module.u_cic.int_1_out[17] ;
 wire \u_top_module.u_cic.int_1_out[18] ;
 wire \u_top_module.u_cic.int_1_out[19] ;
 wire \u_top_module.u_cic.int_1_out[1] ;
 wire \u_top_module.u_cic.int_1_out[20] ;
 wire \u_top_module.u_cic.int_1_out[21] ;
 wire \u_top_module.u_cic.int_1_out[22] ;
 wire \u_top_module.u_cic.int_1_out[23] ;
 wire \u_top_module.u_cic.int_1_out[2] ;
 wire \u_top_module.u_cic.int_1_out[3] ;
 wire \u_top_module.u_cic.int_1_out[4] ;
 wire \u_top_module.u_cic.int_1_out[5] ;
 wire \u_top_module.u_cic.int_1_out[6] ;
 wire \u_top_module.u_cic.int_1_out[7] ;
 wire \u_top_module.u_cic.int_1_out[8] ;
 wire \u_top_module.u_cic.int_1_out[9] ;
 wire \u_top_module.u_cic.int_2_out[10] ;
 wire \u_top_module.u_cic.int_2_out[11] ;
 wire \u_top_module.u_cic.int_2_out[12] ;
 wire \u_top_module.u_cic.int_2_out[13] ;
 wire \u_top_module.u_cic.int_2_out[14] ;
 wire \u_top_module.u_cic.int_2_out[15] ;
 wire \u_top_module.u_cic.int_2_out[16] ;
 wire \u_top_module.u_cic.int_2_out[17] ;
 wire \u_top_module.u_cic.int_2_out[18] ;
 wire \u_top_module.u_cic.int_2_out[19] ;
 wire \u_top_module.u_cic.int_2_out[1] ;
 wire \u_top_module.u_cic.int_2_out[20] ;
 wire \u_top_module.u_cic.int_2_out[21] ;
 wire \u_top_module.u_cic.int_2_out[22] ;
 wire \u_top_module.u_cic.int_2_out[23] ;
 wire \u_top_module.u_cic.int_2_out[2] ;
 wire \u_top_module.u_cic.int_2_out[3] ;
 wire \u_top_module.u_cic.int_2_out[4] ;
 wire \u_top_module.u_cic.int_2_out[5] ;
 wire \u_top_module.u_cic.int_2_out[6] ;
 wire \u_top_module.u_cic.int_2_out[7] ;
 wire \u_top_module.u_cic.int_2_out[8] ;
 wire \u_top_module.u_cic.int_2_out[9] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[10] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[11] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[12] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[13] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[14] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[15] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[16] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[17] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[18] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[19] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[1] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[20] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[21] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[22] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[23] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[2] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[3] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[4] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[5] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[6] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[7] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[8] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d1[9] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[0] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[10] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[11] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[12] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[13] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[14] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[15] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[16] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[17] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[18] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[19] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[1] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[20] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[21] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[22] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[23] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[2] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[3] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[4] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[5] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[6] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[7] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[8] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d2[9] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[0] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[10] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[11] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[12] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[13] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[14] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[15] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[16] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[17] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[18] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[19] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[1] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[20] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[21] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[22] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[23] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[2] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[3] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[4] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[5] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[6] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[7] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[8] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.d3[9] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.sel[0] ;
 wire \u_top_module.u_cic.u_differentiator.a_mux4to1.sel[1] ;
 wire \u_top_module.u_cic.u_differentiator.count[2] ;
 wire \u_top_module.u_cic.u_differentiator.prev_lr_clk ;
 wire \u_top_module.u_cic.u_differentiator.temp[0] ;
 wire \u_top_module.u_cic.u_differentiator.temp[10] ;
 wire \u_top_module.u_cic.u_differentiator.temp[11] ;
 wire \u_top_module.u_cic.u_differentiator.temp[12] ;
 wire \u_top_module.u_cic.u_differentiator.temp[13] ;
 wire \u_top_module.u_cic.u_differentiator.temp[14] ;
 wire \u_top_module.u_cic.u_differentiator.temp[15] ;
 wire \u_top_module.u_cic.u_differentiator.temp[16] ;
 wire \u_top_module.u_cic.u_differentiator.temp[17] ;
 wire \u_top_module.u_cic.u_differentiator.temp[18] ;
 wire \u_top_module.u_cic.u_differentiator.temp[19] ;
 wire \u_top_module.u_cic.u_differentiator.temp[1] ;
 wire \u_top_module.u_cic.u_differentiator.temp[20] ;
 wire \u_top_module.u_cic.u_differentiator.temp[21] ;
 wire \u_top_module.u_cic.u_differentiator.temp[22] ;
 wire \u_top_module.u_cic.u_differentiator.temp[23] ;
 wire \u_top_module.u_cic.u_differentiator.temp[2] ;
 wire \u_top_module.u_cic.u_differentiator.temp[3] ;
 wire \u_top_module.u_cic.u_differentiator.temp[4] ;
 wire \u_top_module.u_cic.u_differentiator.temp[5] ;
 wire \u_top_module.u_cic.u_differentiator.temp[6] ;
 wire \u_top_module.u_cic.u_differentiator.temp[7] ;
 wire \u_top_module.u_cic.u_differentiator.temp[8] ;
 wire \u_top_module.u_cic.u_differentiator.temp[9] ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.prev_lr_clk ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.out ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[9].u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ;
 wire \u_top_module.u_i2s_bus.u_mux_shift.data ;
 wire \u_top_module.u_i2s_bus.u_mux_shift.sum_res ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.ddr_data_falling ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.ddr_data_rising ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.sdr_data_0 ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.sdr_data_1 ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[1].u_ddr_to_sdr.ddr_data_falling ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[1].u_ddr_to_sdr.ddr_data_rising ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[1].u_ddr_to_sdr.sdr_data_0 ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[1].u_ddr_to_sdr.sdr_data_1 ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[2].u_ddr_to_sdr.ddr_data_falling ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[2].u_ddr_to_sdr.ddr_data_rising ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[2].u_ddr_to_sdr.sdr_data_0 ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[2].u_ddr_to_sdr.sdr_data_1 ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[3].u_ddr_to_sdr.ddr_data_falling ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[3].u_ddr_to_sdr.ddr_data_rising ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[3].u_ddr_to_sdr.sdr_data_0 ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[3].u_ddr_to_sdr.sdr_data_1 ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[4].u_ddr_to_sdr.ddr_data_falling ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[4].u_ddr_to_sdr.ddr_data_rising ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[4].u_ddr_to_sdr.sdr_data_0 ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[4].u_ddr_to_sdr.sdr_data_1 ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.ddr_data_falling ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.ddr_data_rising ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.sdr_data_0 ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.sdr_data_1 ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[6].u_ddr_to_sdr.ddr_data_falling ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[6].u_ddr_to_sdr.ddr_data_rising ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[6].u_ddr_to_sdr.sdr_data_0 ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[6].u_ddr_to_sdr.sdr_data_1 ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[7].u_ddr_to_sdr.ddr_data_falling ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[7].u_ddr_to_sdr.ddr_data_rising ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[7].u_ddr_to_sdr.sdr_data_0 ;
 wire \u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[7].u_ddr_to_sdr.sdr_data_1 ;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;

 sg13g2_inv_1 _1431_ (.Y(_0699_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[1] ));
 sg13g2_inv_1 _1432_ (.Y(_0700_),
    .A(_0037_));
 sg13g2_inv_1 _1433_ (.Y(_0701_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[2] ));
 sg13g2_inv_1 _1434_ (.Y(_0702_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[3] ));
 sg13g2_inv_1 _1435_ (.Y(_0703_),
    .A(_0039_));
 sg13g2_inv_1 _1436_ (.Y(_0704_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[4] ));
 sg13g2_inv_1 _1437_ (.Y(_0705_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[5] ));
 sg13g2_inv_1 _1438_ (.Y(_0706_),
    .A(_0041_));
 sg13g2_inv_1 _1439_ (.Y(_0707_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[6] ));
 sg13g2_inv_1 _1440_ (.Y(_0708_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[7] ));
 sg13g2_inv_1 _1441_ (.Y(_0709_),
    .A(_0043_));
 sg13g2_inv_1 _1442_ (.Y(_0710_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[8] ));
 sg13g2_inv_1 _1443_ (.Y(_0711_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[9] ));
 sg13g2_inv_1 _1444_ (.Y(_0712_),
    .A(_0045_));
 sg13g2_inv_1 _1445_ (.Y(_0713_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[10] ));
 sg13g2_inv_1 _1446_ (.Y(_0714_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[11] ));
 sg13g2_inv_1 _1447_ (.Y(_0715_),
    .A(_0047_));
 sg13g2_inv_1 _1448_ (.Y(_0716_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[12] ));
 sg13g2_inv_1 _1449_ (.Y(_0717_),
    .A(_0049_));
 sg13g2_inv_1 _1450_ (.Y(_0718_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[14] ));
 sg13g2_inv_1 _1451_ (.Y(_0719_),
    .A(_0051_));
 sg13g2_inv_1 _1452_ (.Y(_0720_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[16] ));
 sg13g2_inv_1 _1453_ (.Y(_0721_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[17] ));
 sg13g2_inv_1 _1454_ (.Y(_0722_),
    .A(_0053_));
 sg13g2_inv_1 _1455_ (.Y(_0723_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[18] ));
 sg13g2_inv_1 _1456_ (.Y(_0724_),
    .A(_0055_));
 sg13g2_inv_1 _1457_ (.Y(_0725_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[20] ));
 sg13g2_inv_1 _1458_ (.Y(_0726_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[21] ));
 sg13g2_inv_1 _1459_ (.Y(_0727_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[22] ));
 sg13g2_inv_1 _1460_ (.Y(_0728_),
    .A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[23] ));
 sg13g2_inv_1 _1461_ (.Y(_0729_),
    .A(\u_top_module.u_cic.inc_out[6] ));
 sg13g2_inv_1 _1462_ (.Y(_0730_),
    .A(\u_top_module.u_cic.inc_out[8] ));
 sg13g2_inv_1 _1463_ (.Y(_0731_),
    .A(\u_top_module.u_cic.inc_out[12] ));
 sg13g2_inv_1 _1464_ (.Y(_0732_),
    .A(\u_top_module.u_cic.inc_out[13] ));
 sg13g2_inv_1 _1465_ (.Y(_0733_),
    .A(\u_top_module.u_cic.int_1_out[13] ));
 sg13g2_inv_1 _1466_ (.Y(_0734_),
    .A(\u_top_module.u_cic.u_differentiator.temp[9] ));
 sg13g2_inv_1 _1467_ (.Y(_0735_),
    .A(\u_top_module.u_cic.u_differentiator.temp[17] ));
 sg13g2_inv_1 _1468_ (.Y(_0736_),
    .A(_0032_));
 sg13g2_inv_1 _1469_ (.Y(_0737_),
    .A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.sdr_data_0 ));
 sg13g2_inv_1 _1470_ (.Y(_0125_),
    .A(net134));
 sg13g2_and2_1 _1471_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.out ),
    .B(net171),
    .X(_0170_));
 sg13g2_nor2b_1 _1472_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.prev_lr_clk ),
    .B_N(net11),
    .Y(_0738_));
 sg13g2_nand2b_1 _1473_ (.Y(_0739_),
    .B(net11),
    .A_N(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.prev_lr_clk ));
 sg13g2_mux2_1 _1474_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .S(net80),
    .X(_0010_));
 sg13g2_mux2_1 _1475_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .S(net80),
    .X(_0021_));
 sg13g2_mux2_1 _1476_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .S(net80),
    .X(_0024_));
 sg13g2_mux2_1 _1477_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .S(net80),
    .X(_0025_));
 sg13g2_mux2_1 _1478_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .S(net80),
    .X(_0026_));
 sg13g2_mux2_1 _1479_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .S(net79),
    .X(_0027_));
 sg13g2_mux2_1 _1480_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .S(net79),
    .X(_0028_));
 sg13g2_mux2_1 _1481_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .S(net79),
    .X(_0029_));
 sg13g2_mux2_1 _1482_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .S(net79),
    .X(_0030_));
 sg13g2_mux2_1 _1483_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .S(net79),
    .X(_0000_));
 sg13g2_mux2_1 _1484_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .S(net79),
    .X(_0001_));
 sg13g2_mux2_1 _1485_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .S(net81),
    .X(_0002_));
 sg13g2_mux2_1 _1486_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .S(net81),
    .X(_0003_));
 sg13g2_mux2_1 _1487_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .S(net81),
    .X(_0004_));
 sg13g2_mux2_1 _1488_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .S(net78),
    .X(_0005_));
 sg13g2_mux2_1 _1489_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .S(net78),
    .X(_0006_));
 sg13g2_mux2_1 _1490_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .S(net78),
    .X(_0007_));
 sg13g2_mux2_1 _1491_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .S(net78),
    .X(_0008_));
 sg13g2_mux2_1 _1492_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.sum_res ),
    .S(net78),
    .X(_0009_));
 sg13g2_mux2_1 _1493_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.sum_res ),
    .S(net78),
    .X(_0011_));
 sg13g2_mux2_1 _1494_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.sum_res ),
    .S(net78),
    .X(_0012_));
 sg13g2_mux2_2 _1495_ (.A0(\u_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.out ),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.sum_res ),
    .S(net78),
    .X(_0013_));
 sg13g2_and2_2 _1496_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.sum_res ),
    .B(net79),
    .X(_0740_));
 sg13g2_a21o_1 _1497_ (.A2(net77),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.out ),
    .B1(net70),
    .X(_0014_));
 sg13g2_a21o_1 _1498_ (.A2(net77),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.out ),
    .B1(net70),
    .X(_0015_));
 sg13g2_a21o_1 _1499_ (.A2(net77),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.out ),
    .B1(net70),
    .X(_0016_));
 sg13g2_a21o_1 _1500_ (.A2(net77),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.out ),
    .B1(net70),
    .X(_0017_));
 sg13g2_a21o_1 _1501_ (.A2(_0739_),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.out ),
    .B1(_0740_),
    .X(_0018_));
 sg13g2_a21o_1 _1502_ (.A2(net77),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.out ),
    .B1(net70),
    .X(_0019_));
 sg13g2_a21o_1 _1503_ (.A2(net77),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.out ),
    .B1(net70),
    .X(_0020_));
 sg13g2_a21o_1 _1504_ (.A2(net77),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.out ),
    .B1(net70),
    .X(_0022_));
 sg13g2_a21o_1 _1505_ (.A2(net77),
    .A1(\u_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.out ),
    .B1(net70),
    .X(_0023_));
 sg13g2_and2_1 _1506_ (.A(\u_top_module.u_cic.inc_out[1] ),
    .B(\u_top_module.u_cic.int_1_out[1] ),
    .X(_0741_));
 sg13g2_xor2_1 _1507_ (.B(\u_top_module.u_cic.int_1_out[1] ),
    .A(\u_top_module.u_cic.inc_out[1] ),
    .X(_0056_));
 sg13g2_and2_1 _1508_ (.A(\u_top_module.u_cic.inc_out[2] ),
    .B(\u_top_module.u_cic.int_1_out[2] ),
    .X(_0742_));
 sg13g2_xor2_1 _1509_ (.B(\u_top_module.u_cic.int_1_out[2] ),
    .A(\u_top_module.u_cic.inc_out[2] ),
    .X(_0743_));
 sg13g2_xor2_1 _1510_ (.B(_0743_),
    .A(_0741_),
    .X(_0071_));
 sg13g2_a21oi_1 _1511_ (.A1(_0741_),
    .A2(_0743_),
    .Y(_0744_),
    .B1(_0742_));
 sg13g2_nand2_1 _1512_ (.Y(_0745_),
    .A(\u_top_module.u_cic.inc_out[3] ),
    .B(\u_top_module.u_cic.int_1_out[3] ));
 sg13g2_xnor2_1 _1513_ (.Y(_0746_),
    .A(\u_top_module.u_cic.inc_out[3] ),
    .B(\u_top_module.u_cic.int_1_out[3] ));
 sg13g2_xor2_1 _1514_ (.B(_0746_),
    .A(_0744_),
    .X(_0072_));
 sg13g2_and2_1 _1515_ (.A(\u_top_module.u_cic.inc_out[4] ),
    .B(\u_top_module.u_cic.int_1_out[4] ),
    .X(_0747_));
 sg13g2_xor2_1 _1516_ (.B(\u_top_module.u_cic.int_1_out[4] ),
    .A(\u_top_module.u_cic.inc_out[4] ),
    .X(_0748_));
 sg13g2_o21ai_1 _1517_ (.B1(_0745_),
    .Y(_0749_),
    .A1(_0744_),
    .A2(_0746_));
 sg13g2_xor2_1 _1518_ (.B(_0749_),
    .A(_0748_),
    .X(_0073_));
 sg13g2_a21oi_1 _1519_ (.A1(_0748_),
    .A2(_0749_),
    .Y(_0750_),
    .B1(_0747_));
 sg13g2_nor2_1 _1520_ (.A(\u_top_module.u_cic.inc_out[5] ),
    .B(\u_top_module.u_cic.int_1_out[5] ),
    .Y(_0751_));
 sg13g2_xor2_1 _1521_ (.B(\u_top_module.u_cic.int_1_out[5] ),
    .A(\u_top_module.u_cic.inc_out[5] ),
    .X(_0752_));
 sg13g2_xnor2_1 _1522_ (.Y(_0074_),
    .A(_0750_),
    .B(_0752_));
 sg13g2_nand2_1 _1523_ (.Y(_0753_),
    .A(\u_top_module.u_cic.inc_out[6] ),
    .B(\u_top_module.u_cic.int_1_out[6] ));
 sg13g2_xnor2_1 _1524_ (.Y(_0754_),
    .A(\u_top_module.u_cic.inc_out[6] ),
    .B(\u_top_module.u_cic.int_1_out[6] ));
 sg13g2_a221oi_1 _1525_ (.B2(_0749_),
    .C1(_0747_),
    .B1(_0748_),
    .A1(\u_top_module.u_cic.inc_out[5] ),
    .Y(_0755_),
    .A2(\u_top_module.u_cic.int_1_out[5] ));
 sg13g2_or3_1 _1526_ (.A(_0751_),
    .B(_0754_),
    .C(_0755_),
    .X(_0756_));
 sg13g2_o21ai_1 _1527_ (.B1(_0754_),
    .Y(_0757_),
    .A1(_0751_),
    .A2(_0755_));
 sg13g2_and2_1 _1528_ (.A(_0756_),
    .B(_0757_),
    .X(_0075_));
 sg13g2_and2_1 _1529_ (.A(\u_top_module.u_cic.inc_out[7] ),
    .B(\u_top_module.u_cic.int_1_out[7] ),
    .X(_0758_));
 sg13g2_xor2_1 _1530_ (.B(\u_top_module.u_cic.int_1_out[7] ),
    .A(\u_top_module.u_cic.inc_out[7] ),
    .X(_0759_));
 sg13g2_inv_1 _1531_ (.Y(_0760_),
    .A(_0759_));
 sg13g2_a21oi_2 _1532_ (.B1(_0760_),
    .Y(_0761_),
    .A2(_0756_),
    .A1(_0753_));
 sg13g2_nand3_1 _1533_ (.B(_0756_),
    .C(_0760_),
    .A(_0753_),
    .Y(_0762_));
 sg13g2_nor2b_1 _1534_ (.A(_0761_),
    .B_N(_0762_),
    .Y(_0076_));
 sg13g2_nand2_1 _1535_ (.Y(_0763_),
    .A(\u_top_module.u_cic.inc_out[8] ),
    .B(\u_top_module.u_cic.int_1_out[8] ));
 sg13g2_xor2_1 _1536_ (.B(\u_top_module.u_cic.int_1_out[8] ),
    .A(\u_top_module.u_cic.inc_out[8] ),
    .X(_0764_));
 sg13g2_o21ai_1 _1537_ (.B1(_0764_),
    .Y(_0765_),
    .A1(_0758_),
    .A2(_0761_));
 sg13g2_or3_1 _1538_ (.A(_0758_),
    .B(_0761_),
    .C(_0764_),
    .X(_0766_));
 sg13g2_and2_1 _1539_ (.A(_0765_),
    .B(_0766_),
    .X(_0077_));
 sg13g2_and2_1 _1540_ (.A(_0763_),
    .B(_0765_),
    .X(_0767_));
 sg13g2_nor2_1 _1541_ (.A(\u_top_module.u_cic.inc_out[9] ),
    .B(\u_top_module.u_cic.int_1_out[9] ),
    .Y(_0768_));
 sg13g2_and2_1 _1542_ (.A(\u_top_module.u_cic.inc_out[9] ),
    .B(\u_top_module.u_cic.int_1_out[9] ),
    .X(_0769_));
 sg13g2_nor2_1 _1543_ (.A(_0768_),
    .B(_0769_),
    .Y(_0770_));
 sg13g2_xnor2_1 _1544_ (.Y(_0078_),
    .A(_0767_),
    .B(_0770_));
 sg13g2_nand2_1 _1545_ (.Y(_0771_),
    .A(\u_top_module.u_cic.inc_out[10] ),
    .B(\u_top_module.u_cic.int_1_out[10] ));
 sg13g2_xor2_1 _1546_ (.B(\u_top_module.u_cic.int_1_out[10] ),
    .A(\u_top_module.u_cic.inc_out[10] ),
    .X(_0772_));
 sg13g2_a21oi_1 _1547_ (.A1(_0763_),
    .A2(_0765_),
    .Y(_0773_),
    .B1(_0768_));
 sg13g2_nor2_1 _1548_ (.A(_0769_),
    .B(_0773_),
    .Y(_0774_));
 sg13g2_o21ai_1 _1549_ (.B1(_0772_),
    .Y(_0775_),
    .A1(_0769_),
    .A2(_0773_));
 sg13g2_xnor2_1 _1550_ (.Y(_0057_),
    .A(_0772_),
    .B(_0774_));
 sg13g2_nand2_1 _1551_ (.Y(_0776_),
    .A(_0771_),
    .B(_0775_));
 sg13g2_nor2_1 _1552_ (.A(\u_top_module.u_cic.inc_out[11] ),
    .B(\u_top_module.u_cic.int_1_out[11] ),
    .Y(_0777_));
 sg13g2_and2_1 _1553_ (.A(\u_top_module.u_cic.inc_out[11] ),
    .B(\u_top_module.u_cic.int_1_out[11] ),
    .X(_0778_));
 sg13g2_nor2_1 _1554_ (.A(_0777_),
    .B(_0778_),
    .Y(_0779_));
 sg13g2_xor2_1 _1555_ (.B(_0779_),
    .A(_0776_),
    .X(_0058_));
 sg13g2_nand2_1 _1556_ (.Y(_0780_),
    .A(\u_top_module.u_cic.inc_out[12] ),
    .B(\u_top_module.u_cic.int_1_out[12] ));
 sg13g2_xor2_1 _1557_ (.B(\u_top_module.u_cic.int_1_out[12] ),
    .A(\u_top_module.u_cic.inc_out[12] ),
    .X(_0781_));
 sg13g2_a21oi_1 _1558_ (.A1(_0771_),
    .A2(_0775_),
    .Y(_0782_),
    .B1(_0777_));
 sg13g2_o21ai_1 _1559_ (.B1(_0781_),
    .Y(_0783_),
    .A1(_0778_),
    .A2(_0782_));
 sg13g2_or3_1 _1560_ (.A(_0778_),
    .B(_0781_),
    .C(_0782_),
    .X(_0784_));
 sg13g2_and2_1 _1561_ (.A(_0783_),
    .B(_0784_),
    .X(_0059_));
 sg13g2_nand2_1 _1562_ (.Y(_0785_),
    .A(_0780_),
    .B(_0783_));
 sg13g2_nor2_1 _1563_ (.A(_0732_),
    .B(_0733_),
    .Y(_0786_));
 sg13g2_xnor2_1 _1564_ (.Y(_0787_),
    .A(\u_top_module.u_cic.inc_out[13] ),
    .B(\u_top_module.u_cic.int_1_out[13] ));
 sg13g2_xnor2_1 _1565_ (.Y(_0060_),
    .A(_0785_),
    .B(_0787_));
 sg13g2_nand2_1 _1566_ (.Y(_0788_),
    .A(\u_top_module.u_cic.inc_out[14] ),
    .B(\u_top_module.u_cic.int_1_out[14] ));
 sg13g2_xor2_1 _1567_ (.B(\u_top_module.u_cic.int_1_out[14] ),
    .A(\u_top_module.u_cic.inc_out[14] ),
    .X(_0789_));
 sg13g2_a22oi_1 _1568_ (.Y(_0790_),
    .B1(_0780_),
    .B2(_0783_),
    .A2(_0733_),
    .A1(_0732_));
 sg13g2_o21ai_1 _1569_ (.B1(_0789_),
    .Y(_0791_),
    .A1(_0786_),
    .A2(_0790_));
 sg13g2_or3_1 _1570_ (.A(_0786_),
    .B(_0789_),
    .C(_0790_),
    .X(_0792_));
 sg13g2_and2_1 _1571_ (.A(_0791_),
    .B(_0792_),
    .X(_0061_));
 sg13g2_nand2_1 _1572_ (.Y(_0793_),
    .A(_0788_),
    .B(_0791_));
 sg13g2_nor2_1 _1573_ (.A(\u_top_module.u_cic.inc_out[15] ),
    .B(\u_top_module.u_cic.int_1_out[15] ),
    .Y(_0794_));
 sg13g2_and2_1 _1574_ (.A(\u_top_module.u_cic.inc_out[15] ),
    .B(\u_top_module.u_cic.int_1_out[15] ),
    .X(_0795_));
 sg13g2_or2_1 _1575_ (.X(_0796_),
    .B(_0795_),
    .A(_0794_));
 sg13g2_xnor2_1 _1576_ (.Y(_0062_),
    .A(_0793_),
    .B(_0796_));
 sg13g2_nand2_1 _1577_ (.Y(_0797_),
    .A(\u_top_module.u_cic.inc_out[16] ),
    .B(\u_top_module.u_cic.int_1_out[16] ));
 sg13g2_xor2_1 _1578_ (.B(\u_top_module.u_cic.int_1_out[16] ),
    .A(\u_top_module.u_cic.inc_out[16] ),
    .X(_0798_));
 sg13g2_a21oi_1 _1579_ (.A1(_0788_),
    .A2(_0791_),
    .Y(_0799_),
    .B1(_0794_));
 sg13g2_o21ai_1 _1580_ (.B1(_0798_),
    .Y(_0800_),
    .A1(_0795_),
    .A2(_0799_));
 sg13g2_or3_1 _1581_ (.A(_0795_),
    .B(_0798_),
    .C(_0799_),
    .X(_0801_));
 sg13g2_and2_1 _1582_ (.A(_0800_),
    .B(_0801_),
    .X(_0063_));
 sg13g2_nand2_1 _1583_ (.Y(_0802_),
    .A(_0797_),
    .B(_0800_));
 sg13g2_nor2_1 _1584_ (.A(\u_top_module.u_cic.inc_out[17] ),
    .B(\u_top_module.u_cic.int_1_out[17] ),
    .Y(_0803_));
 sg13g2_and2_1 _1585_ (.A(\u_top_module.u_cic.inc_out[17] ),
    .B(\u_top_module.u_cic.int_1_out[17] ),
    .X(_0804_));
 sg13g2_nor2_1 _1586_ (.A(_0803_),
    .B(_0804_),
    .Y(_0805_));
 sg13g2_xor2_1 _1587_ (.B(_0805_),
    .A(_0802_),
    .X(_0064_));
 sg13g2_nand2_1 _1588_ (.Y(_0806_),
    .A(\u_top_module.u_cic.inc_out[18] ),
    .B(\u_top_module.u_cic.int_1_out[18] ));
 sg13g2_xor2_1 _1589_ (.B(\u_top_module.u_cic.int_1_out[18] ),
    .A(\u_top_module.u_cic.inc_out[18] ),
    .X(_0807_));
 sg13g2_inv_1 _1590_ (.Y(_0808_),
    .A(_0807_));
 sg13g2_a21oi_1 _1591_ (.A1(_0797_),
    .A2(_0800_),
    .Y(_0809_),
    .B1(_0803_));
 sg13g2_o21ai_1 _1592_ (.B1(_0807_),
    .Y(_0810_),
    .A1(_0804_),
    .A2(_0809_));
 sg13g2_nor3_1 _1593_ (.A(_0804_),
    .B(_0808_),
    .C(_0809_),
    .Y(_0811_));
 sg13g2_o21ai_1 _1594_ (.B1(_0808_),
    .Y(_0812_),
    .A1(_0804_),
    .A2(_0809_));
 sg13g2_nand2b_1 _1595_ (.Y(_0065_),
    .B(_0812_),
    .A_N(_0811_));
 sg13g2_nor2_1 _1596_ (.A(\u_top_module.u_cic.inc_out[19] ),
    .B(\u_top_module.u_cic.int_1_out[19] ),
    .Y(_0813_));
 sg13g2_xnor2_1 _1597_ (.Y(_0814_),
    .A(\u_top_module.u_cic.inc_out[19] ),
    .B(\u_top_module.u_cic.int_1_out[19] ));
 sg13g2_nand2_1 _1598_ (.Y(_0815_),
    .A(_0806_),
    .B(_0810_));
 sg13g2_xnor2_1 _1599_ (.Y(_0066_),
    .A(_0814_),
    .B(_0815_));
 sg13g2_xnor2_1 _1600_ (.Y(_0816_),
    .A(\u_top_module.u_cic.inc_out[20] ),
    .B(\u_top_module.u_cic.int_1_out[20] ));
 sg13g2_a22oi_1 _1601_ (.Y(_0817_),
    .B1(\u_top_module.u_cic.inc_out[19] ),
    .B2(\u_top_module.u_cic.int_1_out[19] ),
    .A2(\u_top_module.u_cic.int_1_out[18] ),
    .A1(\u_top_module.u_cic.inc_out[18] ));
 sg13g2_a21o_1 _1602_ (.A2(_0817_),
    .A1(_0810_),
    .B1(_0813_),
    .X(_0818_));
 sg13g2_nor2_1 _1603_ (.A(_0816_),
    .B(_0818_),
    .Y(_0819_));
 sg13g2_xor2_1 _1604_ (.B(_0818_),
    .A(_0816_),
    .X(_0067_));
 sg13g2_a21oi_1 _1605_ (.A1(\u_top_module.u_cic.inc_out[20] ),
    .A2(\u_top_module.u_cic.int_1_out[20] ),
    .Y(_0820_),
    .B1(_0819_));
 sg13g2_nor2_1 _1606_ (.A(\u_top_module.u_cic.inc_out[21] ),
    .B(\u_top_module.u_cic.int_1_out[21] ),
    .Y(_0821_));
 sg13g2_nand2_1 _1607_ (.Y(_0822_),
    .A(\u_top_module.u_cic.inc_out[21] ),
    .B(\u_top_module.u_cic.int_1_out[21] ));
 sg13g2_nor2b_1 _1608_ (.A(_0821_),
    .B_N(_0822_),
    .Y(_0823_));
 sg13g2_xnor2_1 _1609_ (.Y(_0068_),
    .A(_0820_),
    .B(_0823_));
 sg13g2_or2_1 _1610_ (.X(_0824_),
    .B(\u_top_module.u_cic.int_1_out[22] ),
    .A(\u_top_module.u_cic.inc_out[22] ));
 sg13g2_and2_1 _1611_ (.A(\u_top_module.u_cic.inc_out[22] ),
    .B(\u_top_module.u_cic.int_1_out[22] ),
    .X(_0825_));
 sg13g2_xnor2_1 _1612_ (.Y(_0826_),
    .A(\u_top_module.u_cic.inc_out[22] ),
    .B(\u_top_module.u_cic.int_1_out[22] ));
 sg13g2_o21ai_1 _1613_ (.B1(_0822_),
    .Y(_0827_),
    .A1(_0820_),
    .A2(_0821_));
 sg13g2_xnor2_1 _1614_ (.Y(_0069_),
    .A(_0826_),
    .B(_0827_));
 sg13g2_a21oi_1 _1615_ (.A1(_0824_),
    .A2(_0827_),
    .Y(_0828_),
    .B1(_0825_));
 sg13g2_xor2_1 _1616_ (.B(\u_top_module.u_cic.int_1_out[23] ),
    .A(\u_top_module.u_cic.inc_out[23] ),
    .X(_0829_));
 sg13g2_xnor2_1 _1617_ (.Y(_0070_),
    .A(_0828_),
    .B(_0829_));
 sg13g2_and2_1 _1618_ (.A(\u_top_module.u_cic.int_1_out[1] ),
    .B(\u_top_module.u_cic.int_2_out[1] ),
    .X(_0830_));
 sg13g2_xor2_1 _1619_ (.B(\u_top_module.u_cic.int_2_out[1] ),
    .A(\u_top_module.u_cic.int_1_out[1] ),
    .X(_0112_));
 sg13g2_and2_1 _1620_ (.A(\u_top_module.u_cic.int_1_out[2] ),
    .B(\u_top_module.u_cic.int_2_out[2] ),
    .X(_0831_));
 sg13g2_xor2_1 _1621_ (.B(\u_top_module.u_cic.int_2_out[2] ),
    .A(\u_top_module.u_cic.int_1_out[2] ),
    .X(_0832_));
 sg13g2_xor2_1 _1622_ (.B(_0832_),
    .A(_0830_),
    .X(_0117_));
 sg13g2_a21oi_2 _1623_ (.B1(_0831_),
    .Y(_0833_),
    .A2(_0832_),
    .A1(_0830_));
 sg13g2_nand2_1 _1624_ (.Y(_0834_),
    .A(\u_top_module.u_cic.int_1_out[3] ),
    .B(\u_top_module.u_cic.int_2_out[3] ));
 sg13g2_xnor2_1 _1625_ (.Y(_0835_),
    .A(\u_top_module.u_cic.int_1_out[3] ),
    .B(\u_top_module.u_cic.int_2_out[3] ));
 sg13g2_xor2_1 _1626_ (.B(_0835_),
    .A(_0833_),
    .X(_0118_));
 sg13g2_and2_1 _1627_ (.A(\u_top_module.u_cic.int_1_out[4] ),
    .B(\u_top_module.u_cic.int_2_out[4] ),
    .X(_0836_));
 sg13g2_xor2_1 _1628_ (.B(\u_top_module.u_cic.int_2_out[4] ),
    .A(\u_top_module.u_cic.int_1_out[4] ),
    .X(_0837_));
 sg13g2_o21ai_1 _1629_ (.B1(_0834_),
    .Y(_0838_),
    .A1(_0833_),
    .A2(_0835_));
 sg13g2_xor2_1 _1630_ (.B(_0838_),
    .A(_0837_),
    .X(_0119_));
 sg13g2_a21oi_1 _1631_ (.A1(_0837_),
    .A2(_0838_),
    .Y(_0839_),
    .B1(_0836_));
 sg13g2_nor2_1 _1632_ (.A(\u_top_module.u_cic.int_1_out[5] ),
    .B(\u_top_module.u_cic.int_2_out[5] ),
    .Y(_0840_));
 sg13g2_xor2_1 _1633_ (.B(\u_top_module.u_cic.int_2_out[5] ),
    .A(\u_top_module.u_cic.int_1_out[5] ),
    .X(_0841_));
 sg13g2_xnor2_1 _1634_ (.Y(_0120_),
    .A(_0839_),
    .B(_0841_));
 sg13g2_nand2_1 _1635_ (.Y(_0842_),
    .A(\u_top_module.u_cic.int_1_out[6] ),
    .B(\u_top_module.u_cic.int_2_out[6] ));
 sg13g2_xnor2_1 _1636_ (.Y(_0843_),
    .A(\u_top_module.u_cic.int_1_out[6] ),
    .B(\u_top_module.u_cic.int_2_out[6] ));
 sg13g2_a221oi_1 _1637_ (.B2(_0838_),
    .C1(_0836_),
    .B1(_0837_),
    .A1(\u_top_module.u_cic.int_1_out[5] ),
    .Y(_0844_),
    .A2(\u_top_module.u_cic.int_2_out[5] ));
 sg13g2_or3_1 _1638_ (.A(_0840_),
    .B(_0843_),
    .C(_0844_),
    .X(_0845_));
 sg13g2_o21ai_1 _1639_ (.B1(_0843_),
    .Y(_0846_),
    .A1(_0840_),
    .A2(_0844_));
 sg13g2_and2_1 _1640_ (.A(_0845_),
    .B(_0846_),
    .X(_0121_));
 sg13g2_and2_1 _1641_ (.A(\u_top_module.u_cic.int_1_out[7] ),
    .B(\u_top_module.u_cic.int_2_out[7] ),
    .X(_0847_));
 sg13g2_xor2_1 _1642_ (.B(\u_top_module.u_cic.int_2_out[7] ),
    .A(\u_top_module.u_cic.int_1_out[7] ),
    .X(_0848_));
 sg13g2_inv_1 _1643_ (.Y(_0849_),
    .A(_0848_));
 sg13g2_a21oi_2 _1644_ (.B1(_0849_),
    .Y(_0850_),
    .A2(_0845_),
    .A1(_0842_));
 sg13g2_nand3_1 _1645_ (.B(_0845_),
    .C(_0849_),
    .A(_0842_),
    .Y(_0851_));
 sg13g2_nor2b_1 _1646_ (.A(_0850_),
    .B_N(_0851_),
    .Y(_0122_));
 sg13g2_nand2_1 _1647_ (.Y(_0852_),
    .A(\u_top_module.u_cic.int_1_out[8] ),
    .B(\u_top_module.u_cic.int_2_out[8] ));
 sg13g2_xor2_1 _1648_ (.B(\u_top_module.u_cic.int_2_out[8] ),
    .A(\u_top_module.u_cic.int_1_out[8] ),
    .X(_0853_));
 sg13g2_o21ai_1 _1649_ (.B1(_0853_),
    .Y(_0854_),
    .A1(_0847_),
    .A2(_0850_));
 sg13g2_or3_1 _1650_ (.A(_0847_),
    .B(_0850_),
    .C(_0853_),
    .X(_0855_));
 sg13g2_and2_1 _1651_ (.A(_0854_),
    .B(_0855_),
    .X(_0123_));
 sg13g2_and2_1 _1652_ (.A(_0852_),
    .B(_0854_),
    .X(_0856_));
 sg13g2_nor2_1 _1653_ (.A(\u_top_module.u_cic.int_1_out[9] ),
    .B(\u_top_module.u_cic.int_2_out[9] ),
    .Y(_0857_));
 sg13g2_and2_1 _1654_ (.A(\u_top_module.u_cic.int_1_out[9] ),
    .B(\u_top_module.u_cic.int_2_out[9] ),
    .X(_0858_));
 sg13g2_nor2_1 _1655_ (.A(_0857_),
    .B(_0858_),
    .Y(_0859_));
 sg13g2_xnor2_1 _1656_ (.Y(_0124_),
    .A(_0856_),
    .B(_0859_));
 sg13g2_nand2_1 _1657_ (.Y(_0860_),
    .A(\u_top_module.u_cic.int_1_out[10] ),
    .B(\u_top_module.u_cic.int_2_out[10] ));
 sg13g2_xor2_1 _1658_ (.B(\u_top_module.u_cic.int_2_out[10] ),
    .A(\u_top_module.u_cic.int_1_out[10] ),
    .X(_0861_));
 sg13g2_a21oi_1 _1659_ (.A1(_0852_),
    .A2(_0854_),
    .Y(_0862_),
    .B1(_0857_));
 sg13g2_nor2_1 _1660_ (.A(_0858_),
    .B(_0862_),
    .Y(_0863_));
 sg13g2_o21ai_1 _1661_ (.B1(_0861_),
    .Y(_0864_),
    .A1(_0858_),
    .A2(_0862_));
 sg13g2_xnor2_1 _1662_ (.Y(_0102_),
    .A(_0861_),
    .B(_0863_));
 sg13g2_nand2_1 _1663_ (.Y(_0865_),
    .A(_0860_),
    .B(_0864_));
 sg13g2_nor2_1 _1664_ (.A(\u_top_module.u_cic.int_1_out[11] ),
    .B(\u_top_module.u_cic.int_2_out[11] ),
    .Y(_0866_));
 sg13g2_and2_1 _1665_ (.A(\u_top_module.u_cic.int_1_out[11] ),
    .B(\u_top_module.u_cic.int_2_out[11] ),
    .X(_0867_));
 sg13g2_or2_1 _1666_ (.X(_0868_),
    .B(_0867_),
    .A(_0866_));
 sg13g2_xnor2_1 _1667_ (.Y(_0103_),
    .A(_0865_),
    .B(_0868_));
 sg13g2_nand2_1 _1668_ (.Y(_0869_),
    .A(\u_top_module.u_cic.int_1_out[12] ),
    .B(\u_top_module.u_cic.int_2_out[12] ));
 sg13g2_xor2_1 _1669_ (.B(\u_top_module.u_cic.int_2_out[12] ),
    .A(\u_top_module.u_cic.int_1_out[12] ),
    .X(_0870_));
 sg13g2_a21oi_1 _1670_ (.A1(_0860_),
    .A2(_0864_),
    .Y(_0871_),
    .B1(_0866_));
 sg13g2_o21ai_1 _1671_ (.B1(_0870_),
    .Y(_0872_),
    .A1(_0867_),
    .A2(_0871_));
 sg13g2_or3_1 _1672_ (.A(_0867_),
    .B(_0870_),
    .C(_0871_),
    .X(_0873_));
 sg13g2_and2_1 _1673_ (.A(_0872_),
    .B(_0873_),
    .X(_0104_));
 sg13g2_nand2_1 _1674_ (.Y(_0874_),
    .A(_0869_),
    .B(_0872_));
 sg13g2_nor2_1 _1675_ (.A(\u_top_module.u_cic.int_1_out[13] ),
    .B(\u_top_module.u_cic.int_2_out[13] ),
    .Y(_0875_));
 sg13g2_and2_1 _1676_ (.A(\u_top_module.u_cic.int_1_out[13] ),
    .B(\u_top_module.u_cic.int_2_out[13] ),
    .X(_0876_));
 sg13g2_nor2_1 _1677_ (.A(_0875_),
    .B(_0876_),
    .Y(_0877_));
 sg13g2_xor2_1 _1678_ (.B(_0877_),
    .A(_0874_),
    .X(_0105_));
 sg13g2_nand2_1 _1679_ (.Y(_0878_),
    .A(\u_top_module.u_cic.int_1_out[14] ),
    .B(\u_top_module.u_cic.int_2_out[14] ));
 sg13g2_xor2_1 _1680_ (.B(\u_top_module.u_cic.int_2_out[14] ),
    .A(\u_top_module.u_cic.int_1_out[14] ),
    .X(_0879_));
 sg13g2_a21oi_1 _1681_ (.A1(_0869_),
    .A2(_0872_),
    .Y(_0880_),
    .B1(_0875_));
 sg13g2_o21ai_1 _1682_ (.B1(_0879_),
    .Y(_0881_),
    .A1(_0876_),
    .A2(_0880_));
 sg13g2_or3_1 _1683_ (.A(_0876_),
    .B(_0879_),
    .C(_0880_),
    .X(_0882_));
 sg13g2_and2_1 _1684_ (.A(_0881_),
    .B(_0882_),
    .X(_0106_));
 sg13g2_nand2_1 _1685_ (.Y(_0883_),
    .A(_0878_),
    .B(_0881_));
 sg13g2_nor2_1 _1686_ (.A(\u_top_module.u_cic.int_1_out[15] ),
    .B(\u_top_module.u_cic.int_2_out[15] ),
    .Y(_0884_));
 sg13g2_and2_1 _1687_ (.A(\u_top_module.u_cic.int_1_out[15] ),
    .B(\u_top_module.u_cic.int_2_out[15] ),
    .X(_0885_));
 sg13g2_or2_1 _1688_ (.X(_0886_),
    .B(_0885_),
    .A(_0884_));
 sg13g2_xnor2_1 _1689_ (.Y(_0107_),
    .A(_0883_),
    .B(_0886_));
 sg13g2_nand2_1 _1690_ (.Y(_0887_),
    .A(\u_top_module.u_cic.int_1_out[16] ),
    .B(\u_top_module.u_cic.int_2_out[16] ));
 sg13g2_xor2_1 _1691_ (.B(\u_top_module.u_cic.int_2_out[16] ),
    .A(\u_top_module.u_cic.int_1_out[16] ),
    .X(_0888_));
 sg13g2_a21oi_1 _1692_ (.A1(_0878_),
    .A2(_0881_),
    .Y(_0889_),
    .B1(_0884_));
 sg13g2_o21ai_1 _1693_ (.B1(_0888_),
    .Y(_0890_),
    .A1(_0885_),
    .A2(_0889_));
 sg13g2_or3_1 _1694_ (.A(_0885_),
    .B(_0888_),
    .C(_0889_),
    .X(_0891_));
 sg13g2_and2_1 _1695_ (.A(_0890_),
    .B(_0891_),
    .X(_0108_));
 sg13g2_nand2_1 _1696_ (.Y(_0892_),
    .A(_0887_),
    .B(_0890_));
 sg13g2_nor2_1 _1697_ (.A(\u_top_module.u_cic.int_1_out[17] ),
    .B(\u_top_module.u_cic.int_2_out[17] ),
    .Y(_0893_));
 sg13g2_and2_1 _1698_ (.A(\u_top_module.u_cic.int_1_out[17] ),
    .B(\u_top_module.u_cic.int_2_out[17] ),
    .X(_0894_));
 sg13g2_nor2_1 _1699_ (.A(_0893_),
    .B(_0894_),
    .Y(_0895_));
 sg13g2_xor2_1 _1700_ (.B(_0895_),
    .A(_0892_),
    .X(_0109_));
 sg13g2_nand2_1 _1701_ (.Y(_0896_),
    .A(\u_top_module.u_cic.int_1_out[18] ),
    .B(\u_top_module.u_cic.int_2_out[18] ));
 sg13g2_xor2_1 _1702_ (.B(\u_top_module.u_cic.int_2_out[18] ),
    .A(\u_top_module.u_cic.int_1_out[18] ),
    .X(_0897_));
 sg13g2_inv_1 _1703_ (.Y(_0898_),
    .A(_0897_));
 sg13g2_a21oi_2 _1704_ (.B1(_0893_),
    .Y(_0899_),
    .A2(_0890_),
    .A1(_0887_));
 sg13g2_o21ai_1 _1705_ (.B1(_0897_),
    .Y(_0900_),
    .A1(_0894_),
    .A2(_0899_));
 sg13g2_nor3_1 _1706_ (.A(_0894_),
    .B(_0898_),
    .C(_0899_),
    .Y(_0901_));
 sg13g2_o21ai_1 _1707_ (.B1(_0898_),
    .Y(_0902_),
    .A1(_0894_),
    .A2(_0899_));
 sg13g2_nand2b_1 _1708_ (.Y(_0110_),
    .B(_0902_),
    .A_N(_0901_));
 sg13g2_nor2_1 _1709_ (.A(\u_top_module.u_cic.int_1_out[19] ),
    .B(\u_top_module.u_cic.int_2_out[19] ),
    .Y(_0903_));
 sg13g2_xnor2_1 _1710_ (.Y(_0904_),
    .A(\u_top_module.u_cic.int_1_out[19] ),
    .B(\u_top_module.u_cic.int_2_out[19] ));
 sg13g2_nand2_1 _1711_ (.Y(_0905_),
    .A(_0896_),
    .B(_0900_));
 sg13g2_xnor2_1 _1712_ (.Y(_0111_),
    .A(_0904_),
    .B(_0905_));
 sg13g2_xnor2_1 _1713_ (.Y(_0906_),
    .A(\u_top_module.u_cic.int_1_out[20] ),
    .B(\u_top_module.u_cic.int_2_out[20] ));
 sg13g2_a22oi_1 _1714_ (.Y(_0907_),
    .B1(\u_top_module.u_cic.int_2_out[19] ),
    .B2(\u_top_module.u_cic.int_1_out[19] ),
    .A2(\u_top_module.u_cic.int_2_out[18] ),
    .A1(\u_top_module.u_cic.int_1_out[18] ));
 sg13g2_a21o_1 _1715_ (.A2(_0907_),
    .A1(_0900_),
    .B1(_0903_),
    .X(_0908_));
 sg13g2_nor2_1 _1716_ (.A(_0906_),
    .B(_0908_),
    .Y(_0909_));
 sg13g2_xor2_1 _1717_ (.B(_0908_),
    .A(_0906_),
    .X(_0113_));
 sg13g2_a21oi_1 _1718_ (.A1(\u_top_module.u_cic.int_1_out[20] ),
    .A2(\u_top_module.u_cic.int_2_out[20] ),
    .Y(_0910_),
    .B1(_0909_));
 sg13g2_nor2_1 _1719_ (.A(\u_top_module.u_cic.int_1_out[21] ),
    .B(\u_top_module.u_cic.int_2_out[21] ),
    .Y(_0911_));
 sg13g2_nand2_1 _1720_ (.Y(_0912_),
    .A(\u_top_module.u_cic.int_1_out[21] ),
    .B(\u_top_module.u_cic.int_2_out[21] ));
 sg13g2_nor2b_1 _1721_ (.A(_0911_),
    .B_N(_0912_),
    .Y(_0913_));
 sg13g2_xnor2_1 _1722_ (.Y(_0114_),
    .A(_0910_),
    .B(_0913_));
 sg13g2_or2_1 _1723_ (.X(_0914_),
    .B(\u_top_module.u_cic.int_2_out[22] ),
    .A(\u_top_module.u_cic.int_1_out[22] ));
 sg13g2_and2_1 _1724_ (.A(\u_top_module.u_cic.int_1_out[22] ),
    .B(\u_top_module.u_cic.int_2_out[22] ),
    .X(_0915_));
 sg13g2_xnor2_1 _1725_ (.Y(_0916_),
    .A(\u_top_module.u_cic.int_1_out[22] ),
    .B(\u_top_module.u_cic.int_2_out[22] ));
 sg13g2_o21ai_1 _1726_ (.B1(_0912_),
    .Y(_0917_),
    .A1(_0910_),
    .A2(_0911_));
 sg13g2_xnor2_1 _1727_ (.Y(_0115_),
    .A(_0916_),
    .B(_0917_));
 sg13g2_a21oi_1 _1728_ (.A1(_0914_),
    .A2(_0917_),
    .Y(_0918_),
    .B1(_0915_));
 sg13g2_xor2_1 _1729_ (.B(\u_top_module.u_cic.int_2_out[23] ),
    .A(\u_top_module.u_cic.int_1_out[23] ),
    .X(_0919_));
 sg13g2_xnor2_1 _1730_ (.Y(_0116_),
    .A(_0918_),
    .B(_0919_));
 sg13g2_nor2_1 _1731_ (.A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[3].u_ddr_to_sdr.sdr_data_0 ),
    .B(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[2].u_ddr_to_sdr.sdr_data_1 ),
    .Y(_0920_));
 sg13g2_xor2_1 _1732_ (.B(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[2].u_ddr_to_sdr.sdr_data_1 ),
    .A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[3].u_ddr_to_sdr.sdr_data_0 ),
    .X(_0921_));
 sg13g2_xnor2_1 _1733_ (.Y(_0922_),
    .A(_0033_),
    .B(_0921_));
 sg13g2_nand2_1 _1734_ (.Y(_0923_),
    .A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[1].u_ddr_to_sdr.sdr_data_1 ),
    .B(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[1].u_ddr_to_sdr.sdr_data_0 ));
 sg13g2_nor2_1 _1735_ (.A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[1].u_ddr_to_sdr.sdr_data_1 ),
    .B(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[1].u_ddr_to_sdr.sdr_data_0 ),
    .Y(_0924_));
 sg13g2_xor2_1 _1736_ (.B(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[1].u_ddr_to_sdr.sdr_data_0 ),
    .A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[1].u_ddr_to_sdr.sdr_data_1 ),
    .X(_0925_));
 sg13g2_xnor2_1 _1737_ (.Y(_0926_),
    .A(_0032_),
    .B(_0925_));
 sg13g2_nand3_1 _1738_ (.B(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.sdr_data_0 ),
    .C(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.sdr_data_1 ),
    .A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[7].u_ddr_to_sdr.sdr_data_1 ),
    .Y(_0927_));
 sg13g2_nor2_1 _1739_ (.A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[7].u_ddr_to_sdr.sdr_data_1 ),
    .B(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.sdr_data_0 ),
    .Y(_0928_));
 sg13g2_nor3_2 _1740_ (.A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[7].u_ddr_to_sdr.sdr_data_1 ),
    .B(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.sdr_data_0 ),
    .C(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.sdr_data_1 ),
    .Y(_0929_));
 sg13g2_a21oi_1 _1741_ (.A1(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[7].u_ddr_to_sdr.sdr_data_1 ),
    .A2(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.sdr_data_0 ),
    .Y(_0930_),
    .B1(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.sdr_data_1 ));
 sg13g2_nor2_1 _1742_ (.A(_0928_),
    .B(_0930_),
    .Y(_0931_));
 sg13g2_o21ai_1 _1743_ (.B1(_0927_),
    .Y(_0932_),
    .A1(_0929_),
    .A2(_0931_));
 sg13g2_xor2_1 _1744_ (.B(_0932_),
    .A(_0926_),
    .X(_0933_));
 sg13g2_nand2b_1 _1745_ (.Y(_0934_),
    .B(_0933_),
    .A_N(_0922_));
 sg13g2_xnor2_1 _1746_ (.Y(_0935_),
    .A(_0922_),
    .B(_0933_));
 sg13g2_nor2_1 _1747_ (.A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[6].u_ddr_to_sdr.sdr_data_0 ),
    .B(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.sdr_data_1 ),
    .Y(_0936_));
 sg13g2_xor2_1 _1748_ (.B(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.sdr_data_1 ),
    .A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[6].u_ddr_to_sdr.sdr_data_0 ),
    .X(_0937_));
 sg13g2_xnor2_1 _1749_ (.Y(_0938_),
    .A(_0034_),
    .B(_0937_));
 sg13g2_inv_1 _1750_ (.Y(_0939_),
    .A(_0938_));
 sg13g2_nand2_1 _1751_ (.Y(_0940_),
    .A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[4].u_ddr_to_sdr.sdr_data_1 ),
    .B(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[4].u_ddr_to_sdr.sdr_data_0 ));
 sg13g2_nand3_1 _1752_ (.B(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[4].u_ddr_to_sdr.sdr_data_0 ),
    .C(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.sdr_data_0 ),
    .A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[4].u_ddr_to_sdr.sdr_data_1 ),
    .Y(_0941_));
 sg13g2_nor2_2 _1753_ (.A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[4].u_ddr_to_sdr.sdr_data_1 ),
    .B(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[4].u_ddr_to_sdr.sdr_data_0 ),
    .Y(_0942_));
 sg13g2_nand2_1 _1754_ (.Y(_0943_),
    .A(_0737_),
    .B(_0942_));
 sg13g2_o21ai_1 _1755_ (.B1(_0940_),
    .Y(_0944_),
    .A1(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.sdr_data_0 ),
    .A2(_0942_));
 sg13g2_a21oi_1 _1756_ (.A1(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.sdr_data_0 ),
    .A2(_0942_),
    .Y(_0945_),
    .B1(_0944_));
 sg13g2_nor2_1 _1757_ (.A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.sdr_data_0 ),
    .B(_0940_),
    .Y(_0946_));
 sg13g2_nor2_1 _1758_ (.A(_0945_),
    .B(_0946_),
    .Y(_0947_));
 sg13g2_xnor2_1 _1759_ (.Y(_0948_),
    .A(_0939_),
    .B(_0947_));
 sg13g2_nand2_1 _1760_ (.Y(_0949_),
    .A(_0935_),
    .B(_0948_));
 sg13g2_xor2_1 _1761_ (.B(_0948_),
    .A(_0935_),
    .X(_0950_));
 sg13g2_nand2_1 _1762_ (.Y(_0951_),
    .A(_0031_),
    .B(_0950_));
 sg13g2_xnor2_1 _1763_ (.Y(_0952_),
    .A(_0031_),
    .B(_0950_));
 sg13g2_inv_1 _1764_ (.Y(_0953_),
    .A(_0952_));
 sg13g2_nand2_1 _1765_ (.Y(_0954_),
    .A(\u_top_module.u_cic.inc_out[1] ),
    .B(_0953_));
 sg13g2_xnor2_1 _1766_ (.Y(_0079_),
    .A(\u_top_module.u_cic.inc_out[1] ),
    .B(_0952_));
 sg13g2_a21oi_1 _1767_ (.A1(_0034_),
    .A2(_0937_),
    .Y(_0955_),
    .B1(_0936_));
 sg13g2_nor2b_2 _1768_ (.A(_0031_),
    .B_N(_0955_),
    .Y(_0956_));
 sg13g2_xnor2_1 _1769_ (.Y(_0957_),
    .A(_0031_),
    .B(_0955_));
 sg13g2_nor2_2 _1770_ (.A(_0938_),
    .B(_0943_),
    .Y(_0958_));
 sg13g2_nand2_1 _1771_ (.Y(_0959_),
    .A(_0941_),
    .B(_0943_));
 sg13g2_xnor2_1 _1772_ (.Y(_0960_),
    .A(_0938_),
    .B(_0959_));
 sg13g2_o21ai_1 _1773_ (.B1(_0960_),
    .Y(_0961_),
    .A1(_0938_),
    .A2(_0947_));
 sg13g2_nor2b_1 _1774_ (.A(_0958_),
    .B_N(_0961_),
    .Y(_0962_));
 sg13g2_a21oi_2 _1775_ (.B1(_0920_),
    .Y(_0963_),
    .A2(_0921_),
    .A1(_0033_));
 sg13g2_inv_1 _1776_ (.Y(_0964_),
    .A(_0963_));
 sg13g2_a21oi_2 _1777_ (.B1(_0924_),
    .Y(_0965_),
    .A2(_0923_),
    .A1(_0032_));
 sg13g2_nor2_1 _1778_ (.A(_0922_),
    .B(_0965_),
    .Y(_0966_));
 sg13g2_nand2_1 _1779_ (.Y(_0967_),
    .A(_0922_),
    .B(_0965_));
 sg13g2_xor2_1 _1780_ (.B(_0965_),
    .A(_0922_),
    .X(_0968_));
 sg13g2_xnor2_1 _1781_ (.Y(_0969_),
    .A(_0963_),
    .B(_0968_));
 sg13g2_nor2_1 _1782_ (.A(_0926_),
    .B(_0931_),
    .Y(_0970_));
 sg13g2_nor2b_1 _1783_ (.A(_0927_),
    .B_N(_0926_),
    .Y(_0971_));
 sg13g2_nor3_1 _1784_ (.A(_0929_),
    .B(_0970_),
    .C(_0971_),
    .Y(_0972_));
 sg13g2_xnor2_1 _1785_ (.Y(_0973_),
    .A(_0969_),
    .B(_0972_));
 sg13g2_nor2_1 _1786_ (.A(_0934_),
    .B(_0973_),
    .Y(_0974_));
 sg13g2_nand2_1 _1787_ (.Y(_0975_),
    .A(_0934_),
    .B(_0973_));
 sg13g2_xnor2_1 _1788_ (.Y(_0976_),
    .A(_0934_),
    .B(_0973_));
 sg13g2_xor2_1 _1789_ (.B(_0976_),
    .A(_0962_),
    .X(_0977_));
 sg13g2_nor2_1 _1790_ (.A(_0949_),
    .B(_0977_),
    .Y(_0978_));
 sg13g2_xor2_1 _1791_ (.B(_0977_),
    .A(_0949_),
    .X(_0979_));
 sg13g2_xnor2_1 _1792_ (.Y(_0980_),
    .A(_0957_),
    .B(_0979_));
 sg13g2_nor2_1 _1793_ (.A(_0951_),
    .B(_0980_),
    .Y(_0981_));
 sg13g2_or2_1 _1794_ (.X(_0982_),
    .B(_0980_),
    .A(_0951_));
 sg13g2_xor2_1 _1795_ (.B(_0980_),
    .A(_0951_),
    .X(_0983_));
 sg13g2_nand2_1 _1796_ (.Y(_0984_),
    .A(\u_top_module.u_cic.inc_out[2] ),
    .B(_0983_));
 sg13g2_xnor2_1 _1797_ (.Y(_0985_),
    .A(\u_top_module.u_cic.inc_out[2] ),
    .B(_0983_));
 sg13g2_xor2_1 _1798_ (.B(_0985_),
    .A(_0954_),
    .X(_0094_));
 sg13g2_o21ai_1 _1799_ (.B1(_0984_),
    .Y(_0986_),
    .A1(_0954_),
    .A2(_0985_));
 sg13g2_a21oi_2 _1800_ (.B1(_0978_),
    .Y(_0987_),
    .A2(_0979_),
    .A1(_0957_));
 sg13g2_a21o_1 _1801_ (.A2(_0979_),
    .A1(_0957_),
    .B1(_0978_),
    .X(_0988_));
 sg13g2_a21oi_1 _1802_ (.A1(_0962_),
    .A2(_0975_),
    .Y(_0989_),
    .B1(_0974_));
 sg13g2_a22oi_1 _1803_ (.Y(_0990_),
    .B1(_0942_),
    .B2(_0737_),
    .A2(_0941_),
    .A1(_0939_));
 sg13g2_a21oi_2 _1804_ (.B1(_0966_),
    .Y(_0991_),
    .A2(_0967_),
    .A1(_0964_));
 sg13g2_xor2_1 _1805_ (.B(_0991_),
    .A(_0960_),
    .X(_0992_));
 sg13g2_nand2b_1 _1806_ (.Y(_0993_),
    .B(_0992_),
    .A_N(_0990_));
 sg13g2_xnor2_1 _1807_ (.Y(_0994_),
    .A(_0990_),
    .B(_0992_));
 sg13g2_nor2b_2 _1808_ (.A(_0926_),
    .B_N(_0929_),
    .Y(_0995_));
 sg13g2_a21oi_1 _1809_ (.A1(_0969_),
    .A2(_0972_),
    .Y(_0996_),
    .B1(_0995_));
 sg13g2_nor2_1 _1810_ (.A(_0971_),
    .B(_0995_),
    .Y(_0997_));
 sg13g2_xor2_1 _1811_ (.B(_0997_),
    .A(_0969_),
    .X(_0998_));
 sg13g2_xnor2_1 _1812_ (.Y(_0999_),
    .A(_0996_),
    .B(_0998_));
 sg13g2_xnor2_1 _1813_ (.Y(_1000_),
    .A(_0994_),
    .B(_0999_));
 sg13g2_nor2_1 _1814_ (.A(_0989_),
    .B(_1000_),
    .Y(_1001_));
 sg13g2_xor2_1 _1815_ (.B(_1000_),
    .A(_0989_),
    .X(_1002_));
 sg13g2_nor2b_1 _1816_ (.A(_0956_),
    .B_N(_0958_),
    .Y(_1003_));
 sg13g2_nand2b_1 _1817_ (.Y(_1004_),
    .B(_0958_),
    .A_N(_0956_));
 sg13g2_xnor2_1 _1818_ (.Y(_1005_),
    .A(_0956_),
    .B(_0958_));
 sg13g2_xnor2_1 _1819_ (.Y(_1006_),
    .A(_1002_),
    .B(_1005_));
 sg13g2_nor2_1 _1820_ (.A(_0987_),
    .B(_1006_),
    .Y(_1007_));
 sg13g2_and2_1 _1821_ (.A(_0987_),
    .B(_1006_),
    .X(_1008_));
 sg13g2_xnor2_1 _1822_ (.Y(_1009_),
    .A(_0988_),
    .B(_1006_));
 sg13g2_xnor2_1 _1823_ (.Y(_1010_),
    .A(_0982_),
    .B(_1009_));
 sg13g2_xnor2_1 _1824_ (.Y(_1011_),
    .A(\u_top_module.u_cic.inc_out[3] ),
    .B(_1010_));
 sg13g2_nor2b_1 _1825_ (.A(_1011_),
    .B_N(_0986_),
    .Y(_1012_));
 sg13g2_xnor2_1 _1826_ (.Y(_0095_),
    .A(_0986_),
    .B(_1011_));
 sg13g2_nand3b_1 _1827_ (.B(_1004_),
    .C(_0988_),
    .Y(_1013_),
    .A_N(_1006_));
 sg13g2_o21ai_1 _1828_ (.B1(_1003_),
    .Y(_1014_),
    .A1(_0987_),
    .A2(_1006_));
 sg13g2_o21ai_1 _1829_ (.B1(_1004_),
    .Y(_1015_),
    .A1(_0987_),
    .A2(_1006_));
 sg13g2_nand3_1 _1830_ (.B(_1002_),
    .C(_1003_),
    .A(_0988_),
    .Y(_1016_));
 sg13g2_a22oi_1 _1831_ (.Y(_1017_),
    .B1(_1013_),
    .B2(_1014_),
    .A2(_1009_),
    .A1(_0981_));
 sg13g2_nor4_2 _1832_ (.A(_0982_),
    .B(_1003_),
    .C(_1007_),
    .Y(_1018_),
    .D(_1008_));
 sg13g2_a22oi_1 _1833_ (.Y(_1019_),
    .B1(_1015_),
    .B2(_1016_),
    .A2(_1009_),
    .A1(_0981_));
 sg13g2_nor4_2 _1834_ (.A(_0982_),
    .B(_1004_),
    .C(_1007_),
    .Y(_1020_),
    .D(_1008_));
 sg13g2_a22oi_1 _1835_ (.Y(_1021_),
    .B1(_0999_),
    .B2(_0994_),
    .A2(_0995_),
    .A1(_0969_));
 sg13g2_a21oi_1 _1836_ (.A1(_0969_),
    .A2(_0997_),
    .Y(_1022_),
    .B1(_0995_));
 sg13g2_xor2_1 _1837_ (.B(_0956_),
    .A(_0034_),
    .X(_1023_));
 sg13g2_xnor2_1 _1838_ (.Y(_1024_),
    .A(_1022_),
    .B(_1023_));
 sg13g2_xnor2_1 _1839_ (.Y(_1025_),
    .A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[3].u_ddr_to_sdr.sdr_data_1 ),
    .B(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.sdr_data_0 ));
 sg13g2_xnor2_1 _1840_ (.Y(_1026_),
    .A(_0937_),
    .B(_1025_));
 sg13g2_xnor2_1 _1841_ (.Y(_1027_),
    .A(_0944_),
    .B(_1026_));
 sg13g2_a21oi_1 _1842_ (.A1(_0926_),
    .A2(_0927_),
    .Y(_1028_),
    .B1(_0929_));
 sg13g2_xnor2_1 _1843_ (.Y(_1029_),
    .A(_1027_),
    .B(_1028_));
 sg13g2_a21oi_1 _1844_ (.A1(_0736_),
    .A2(_0923_),
    .Y(_1030_),
    .B1(_0924_));
 sg13g2_xor2_1 _1845_ (.B(_0921_),
    .A(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[2].u_ddr_to_sdr.sdr_data_0 ),
    .X(_1031_));
 sg13g2_xor2_1 _1846_ (.B(_1030_),
    .A(_0990_),
    .X(_1032_));
 sg13g2_xnor2_1 _1847_ (.Y(_1033_),
    .A(_1029_),
    .B(_1032_));
 sg13g2_xnor2_1 _1848_ (.Y(_1034_),
    .A(_0963_),
    .B(_1031_));
 sg13g2_xnor2_1 _1849_ (.Y(_1035_),
    .A(_0991_),
    .B(_1034_));
 sg13g2_xnor2_1 _1850_ (.Y(_1036_),
    .A(_1033_),
    .B(_1035_));
 sg13g2_xnor2_1 _1851_ (.Y(_1037_),
    .A(_1024_),
    .B(_1036_));
 sg13g2_xnor2_1 _1852_ (.Y(_1038_),
    .A(_1021_),
    .B(_1037_));
 sg13g2_a21oi_1 _1853_ (.A1(_1002_),
    .A2(_1005_),
    .Y(_1039_),
    .B1(_1001_));
 sg13g2_o21ai_1 _1854_ (.B1(_0993_),
    .Y(_1040_),
    .A1(_0960_),
    .A2(_0991_));
 sg13g2_xnor2_1 _1855_ (.Y(_1041_),
    .A(_1038_),
    .B(_1040_));
 sg13g2_xnor2_1 _1856_ (.Y(_1042_),
    .A(_1039_),
    .B(_1041_));
 sg13g2_xor2_1 _1857_ (.B(_1041_),
    .A(_1039_),
    .X(_1043_));
 sg13g2_nor3_2 _1858_ (.A(_1019_),
    .B(_1020_),
    .C(_1043_),
    .Y(_1044_));
 sg13g2_o21ai_1 _1859_ (.B1(_1042_),
    .Y(_1045_),
    .A1(_1017_),
    .A2(_1018_));
 sg13g2_nor3_2 _1860_ (.A(_1017_),
    .B(_1018_),
    .C(_1042_),
    .Y(_1046_));
 sg13g2_o21ai_1 _1861_ (.B1(_1043_),
    .Y(_1047_),
    .A1(_1019_),
    .A2(_1020_));
 sg13g2_nand2_1 _1862_ (.Y(_1048_),
    .A(_1045_),
    .B(_1047_));
 sg13g2_nor2_2 _1863_ (.A(_1044_),
    .B(_1046_),
    .Y(_1049_));
 sg13g2_nand2_1 _1864_ (.Y(_1050_),
    .A(\u_top_module.u_cic.inc_out[4] ),
    .B(net17));
 sg13g2_xnor2_1 _1865_ (.Y(_1051_),
    .A(\u_top_module.u_cic.inc_out[4] ),
    .B(net16));
 sg13g2_a21oi_2 _1866_ (.B1(_1012_),
    .Y(_1052_),
    .A2(_1010_),
    .A1(\u_top_module.u_cic.inc_out[3] ));
 sg13g2_xor2_1 _1867_ (.B(_1052_),
    .A(_1051_),
    .X(_0096_));
 sg13g2_xnor2_1 _1868_ (.Y(_1053_),
    .A(\u_top_module.u_cic.inc_out[5] ),
    .B(net17));
 sg13g2_o21ai_1 _1869_ (.B1(_1050_),
    .Y(_1054_),
    .A1(_1051_),
    .A2(_1052_));
 sg13g2_xnor2_1 _1870_ (.Y(_0097_),
    .A(_1053_),
    .B(_1054_));
 sg13g2_nand3_1 _1871_ (.B(_1045_),
    .C(_1047_),
    .A(_0729_),
    .Y(_1055_));
 sg13g2_nor2_1 _1872_ (.A(_0729_),
    .B(_1049_),
    .Y(_1056_));
 sg13g2_o21ai_1 _1873_ (.B1(\u_top_module.u_cic.inc_out[6] ),
    .Y(_1057_),
    .A1(_1044_),
    .A2(_1046_));
 sg13g2_nand2_1 _1874_ (.Y(_1058_),
    .A(_1055_),
    .B(_1057_));
 sg13g2_nor3_1 _1875_ (.A(_1051_),
    .B(_1052_),
    .C(_1053_),
    .Y(_1059_));
 sg13g2_o21ai_1 _1876_ (.B1(net17),
    .Y(_1060_),
    .A1(\u_top_module.u_cic.inc_out[4] ),
    .A2(\u_top_module.u_cic.inc_out[5] ));
 sg13g2_nand2b_1 _1877_ (.Y(_1061_),
    .B(_1060_),
    .A_N(_1059_));
 sg13g2_xnor2_1 _1878_ (.Y(_0098_),
    .A(_1058_),
    .B(_1061_));
 sg13g2_o21ai_1 _1879_ (.B1(\u_top_module.u_cic.inc_out[7] ),
    .Y(_1062_),
    .A1(_1044_),
    .A2(_1046_));
 sg13g2_nand3b_1 _1880_ (.B(_1045_),
    .C(_1047_),
    .Y(_1063_),
    .A_N(\u_top_module.u_cic.inc_out[7] ));
 sg13g2_nand2_1 _1881_ (.Y(_1064_),
    .A(_1062_),
    .B(_1063_));
 sg13g2_a21oi_1 _1882_ (.A1(_1055_),
    .A2(_1061_),
    .Y(_1065_),
    .B1(_1056_));
 sg13g2_xor2_1 _1883_ (.B(_1065_),
    .A(_1064_),
    .X(_0099_));
 sg13g2_nor2_1 _1884_ (.A(_1058_),
    .B(_1064_),
    .Y(_1066_));
 sg13g2_nand4_1 _1885_ (.B(_1057_),
    .C(_1062_),
    .A(_1055_),
    .Y(_1067_),
    .D(_1063_));
 sg13g2_and2_1 _1886_ (.A(_1057_),
    .B(_1062_),
    .X(_1068_));
 sg13g2_o21ai_1 _1887_ (.B1(_1068_),
    .Y(_1069_),
    .A1(_1060_),
    .A2(_1067_));
 sg13g2_a21o_2 _1888_ (.A2(_1066_),
    .A1(_1059_),
    .B1(_1069_),
    .X(_1070_));
 sg13g2_xnor2_1 _1889_ (.Y(_1071_),
    .A(\u_top_module.u_cic.inc_out[8] ),
    .B(net16));
 sg13g2_nand2b_1 _1890_ (.Y(_1072_),
    .B(_1070_),
    .A_N(_1071_));
 sg13g2_xnor2_1 _1891_ (.Y(_0100_),
    .A(_1070_),
    .B(_1071_));
 sg13g2_xnor2_1 _1892_ (.Y(_1073_),
    .A(\u_top_module.u_cic.inc_out[9] ),
    .B(net16));
 sg13g2_o21ai_1 _1893_ (.B1(_1072_),
    .Y(_1074_),
    .A1(_0730_),
    .A2(_1049_));
 sg13g2_xnor2_1 _1894_ (.Y(_0101_),
    .A(_1073_),
    .B(_1074_));
 sg13g2_xnor2_1 _1895_ (.Y(_1075_),
    .A(\u_top_module.u_cic.inc_out[10] ),
    .B(net16));
 sg13g2_o21ai_1 _1896_ (.B1(net16),
    .Y(_0290_),
    .A1(\u_top_module.u_cic.inc_out[8] ),
    .A2(\u_top_module.u_cic.inc_out[9] ));
 sg13g2_inv_1 _1897_ (.Y(_0291_),
    .A(_0290_));
 sg13g2_o21ai_1 _1898_ (.B1(_0290_),
    .Y(_0292_),
    .A1(_1072_),
    .A2(_1073_));
 sg13g2_nor2b_1 _1899_ (.A(_1075_),
    .B_N(_0292_),
    .Y(_0293_));
 sg13g2_xnor2_1 _1900_ (.Y(_0080_),
    .A(_1075_),
    .B(_0292_));
 sg13g2_xnor2_1 _1901_ (.Y(_0294_),
    .A(\u_top_module.u_cic.inc_out[11] ),
    .B(net16));
 sg13g2_a21oi_1 _1902_ (.A1(\u_top_module.u_cic.inc_out[10] ),
    .A2(net16),
    .Y(_0295_),
    .B1(_0293_));
 sg13g2_xor2_1 _1903_ (.B(_0295_),
    .A(_0294_),
    .X(_0081_));
 sg13g2_nor2_1 _1904_ (.A(_1075_),
    .B(_0294_),
    .Y(_0296_));
 sg13g2_nor4_1 _1905_ (.A(_1071_),
    .B(_1073_),
    .C(_1075_),
    .D(_0294_),
    .Y(_0297_));
 sg13g2_o21ai_1 _1906_ (.B1(net16),
    .Y(_0298_),
    .A1(\u_top_module.u_cic.inc_out[10] ),
    .A2(\u_top_module.u_cic.inc_out[11] ));
 sg13g2_inv_1 _1907_ (.Y(_0299_),
    .A(_0298_));
 sg13g2_a221oi_1 _1908_ (.B2(_1070_),
    .C1(_0299_),
    .B1(_0297_),
    .A1(_0291_),
    .Y(_0300_),
    .A2(_0296_));
 sg13g2_xnor2_1 _1909_ (.Y(_0301_),
    .A(\u_top_module.u_cic.inc_out[12] ),
    .B(net15));
 sg13g2_or2_1 _1910_ (.X(_0302_),
    .B(_0301_),
    .A(_0300_));
 sg13g2_xor2_1 _1911_ (.B(_0301_),
    .A(_0300_),
    .X(_0082_));
 sg13g2_xnor2_1 _1912_ (.Y(_0303_),
    .A(\u_top_module.u_cic.inc_out[13] ),
    .B(net14));
 sg13g2_o21ai_1 _1913_ (.B1(_0302_),
    .Y(_0304_),
    .A1(_0731_),
    .A2(_1049_));
 sg13g2_xnor2_1 _1914_ (.Y(_0083_),
    .A(_0303_),
    .B(_0304_));
 sg13g2_xnor2_1 _1915_ (.Y(_0305_),
    .A(\u_top_module.u_cic.inc_out[14] ),
    .B(net14));
 sg13g2_o21ai_1 _1916_ (.B1(net14),
    .Y(_0306_),
    .A1(\u_top_module.u_cic.inc_out[12] ),
    .A2(\u_top_module.u_cic.inc_out[13] ));
 sg13g2_a22oi_1 _1917_ (.Y(_0307_),
    .B1(_0302_),
    .B2(_0306_),
    .A2(_1049_),
    .A1(_0732_));
 sg13g2_nor2b_1 _1918_ (.A(_0305_),
    .B_N(_0307_),
    .Y(_0308_));
 sg13g2_xnor2_1 _1919_ (.Y(_0084_),
    .A(_0305_),
    .B(_0307_));
 sg13g2_xnor2_1 _1920_ (.Y(_0309_),
    .A(\u_top_module.u_cic.inc_out[15] ),
    .B(net14));
 sg13g2_a21oi_1 _1921_ (.A1(\u_top_module.u_cic.inc_out[14] ),
    .A2(net14),
    .Y(_0310_),
    .B1(_0308_));
 sg13g2_xor2_1 _1922_ (.B(_0310_),
    .A(_0309_),
    .X(_0085_));
 sg13g2_or4_1 _1923_ (.A(_0301_),
    .B(_0303_),
    .C(_0305_),
    .D(_0309_),
    .X(_0311_));
 sg13g2_o21ai_1 _1924_ (.B1(net14),
    .Y(_0312_),
    .A1(\u_top_module.u_cic.inc_out[14] ),
    .A2(\u_top_module.u_cic.inc_out[15] ));
 sg13g2_nor3_1 _1925_ (.A(_0305_),
    .B(_0306_),
    .C(_0309_),
    .Y(_0313_));
 sg13g2_nor2b_1 _1926_ (.A(_0313_),
    .B_N(_0312_),
    .Y(_0314_));
 sg13g2_o21ai_1 _1927_ (.B1(_0314_),
    .Y(_0315_),
    .A1(_0300_),
    .A2(_0311_));
 sg13g2_xnor2_1 _1928_ (.Y(_0316_),
    .A(\u_top_module.u_cic.inc_out[16] ),
    .B(net14));
 sg13g2_nor2b_1 _1929_ (.A(_0316_),
    .B_N(_0315_),
    .Y(_0317_));
 sg13g2_xnor2_1 _1930_ (.Y(_0086_),
    .A(_0315_),
    .B(_0316_));
 sg13g2_a21o_1 _1931_ (.A2(net12),
    .A1(\u_top_module.u_cic.inc_out[16] ),
    .B1(_0317_),
    .X(_0318_));
 sg13g2_xnor2_1 _1932_ (.Y(_0319_),
    .A(_0035_),
    .B(net14));
 sg13g2_inv_1 _1933_ (.Y(_0320_),
    .A(_0319_));
 sg13g2_xnor2_1 _1934_ (.Y(_0087_),
    .A(_0318_),
    .B(_0320_));
 sg13g2_nand2_1 _1935_ (.Y(_0321_),
    .A(\u_top_module.u_cic.inc_out[18] ),
    .B(net13));
 sg13g2_xnor2_1 _1936_ (.Y(_0322_),
    .A(\u_top_module.u_cic.inc_out[18] ),
    .B(net13));
 sg13g2_a21oi_1 _1937_ (.A1(\u_top_module.u_cic.inc_out[16] ),
    .A2(_0035_),
    .Y(_0323_),
    .B1(\u_top_module.u_cic.inc_out[17] ));
 sg13g2_nor2_1 _1938_ (.A(_1049_),
    .B(_0323_),
    .Y(_0324_));
 sg13g2_a21oi_1 _1939_ (.A1(_0317_),
    .A2(_0319_),
    .Y(_0325_),
    .B1(_0324_));
 sg13g2_xor2_1 _1940_ (.B(_0325_),
    .A(_0322_),
    .X(_0088_));
 sg13g2_o21ai_1 _1941_ (.B1(_0321_),
    .Y(_0326_),
    .A1(_0322_),
    .A2(_0325_));
 sg13g2_xnor2_1 _1942_ (.Y(_0327_),
    .A(\u_top_module.u_cic.inc_out[19] ),
    .B(net13));
 sg13g2_xnor2_1 _1943_ (.Y(_0089_),
    .A(_0326_),
    .B(_0327_));
 sg13g2_nor4_1 _1944_ (.A(_0316_),
    .B(_0320_),
    .C(_0322_),
    .D(_0327_),
    .Y(_0328_));
 sg13g2_o21ai_1 _1945_ (.B1(net13),
    .Y(_0329_),
    .A1(\u_top_module.u_cic.inc_out[18] ),
    .A2(\u_top_module.u_cic.inc_out[19] ));
 sg13g2_nand2b_1 _1946_ (.Y(_0330_),
    .B(_0329_),
    .A_N(_0324_));
 sg13g2_a21oi_2 _1947_ (.B1(_0330_),
    .Y(_0331_),
    .A2(_0328_),
    .A1(_0315_));
 sg13g2_nand2_1 _1948_ (.Y(_0332_),
    .A(\u_top_module.u_cic.inc_out[20] ),
    .B(net12));
 sg13g2_xnor2_1 _1949_ (.Y(_0333_),
    .A(\u_top_module.u_cic.inc_out[20] ),
    .B(net12));
 sg13g2_xor2_1 _1950_ (.B(_0333_),
    .A(_0331_),
    .X(_0090_));
 sg13g2_nand2b_1 _1951_ (.Y(_0334_),
    .B(_1049_),
    .A_N(\u_top_module.u_cic.inc_out[21] ));
 sg13g2_and2_1 _1952_ (.A(\u_top_module.u_cic.inc_out[21] ),
    .B(net12),
    .X(_0335_));
 sg13g2_xnor2_1 _1953_ (.Y(_0336_),
    .A(\u_top_module.u_cic.inc_out[21] ),
    .B(net12));
 sg13g2_o21ai_1 _1954_ (.B1(_0332_),
    .Y(_0337_),
    .A1(_0331_),
    .A2(_0333_));
 sg13g2_xnor2_1 _1955_ (.Y(_0091_),
    .A(_0336_),
    .B(_0337_));
 sg13g2_nand2_1 _1956_ (.Y(_0338_),
    .A(\u_top_module.u_cic.inc_out[22] ),
    .B(net12));
 sg13g2_xnor2_1 _1957_ (.Y(_0339_),
    .A(\u_top_module.u_cic.inc_out[22] ),
    .B(net12));
 sg13g2_a21oi_1 _1958_ (.A1(_0334_),
    .A2(_0337_),
    .Y(_0340_),
    .B1(_0335_));
 sg13g2_xor2_1 _1959_ (.B(_0340_),
    .A(_0339_),
    .X(_0092_));
 sg13g2_o21ai_1 _1960_ (.B1(_0338_),
    .Y(_0341_),
    .A1(_0339_),
    .A2(_0340_));
 sg13g2_xnor2_1 _1961_ (.Y(_0342_),
    .A(\u_top_module.u_cic.inc_out[23] ),
    .B(net12));
 sg13g2_xnor2_1 _1962_ (.Y(_0093_),
    .A(_0341_),
    .B(_0342_));
 sg13g2_and2_1 _1963_ (.A(\u_top_module.u_i2s_bus.u_mux_shift.sum_res ),
    .B(net79),
    .X(_0166_));
 sg13g2_nor2b_2 _1964_ (.A(\u_top_module.u_cic.u_differentiator.prev_lr_clk ),
    .B_N(net11),
    .Y(_0343_));
 sg13g2_or2_2 _1965_ (.X(_0344_),
    .B(_0343_),
    .A(\u_top_module.u_cic.u_differentiator.count[2] ));
 sg13g2_nand3b_1 _1966_ (.B(\u_top_module.u_cic.u_differentiator.count[2] ),
    .C(net92),
    .Y(_0345_),
    .A_N(_0343_));
 sg13g2_o21ai_1 _1967_ (.B1(_0345_),
    .Y(_0167_),
    .A1(net92),
    .A2(_0344_));
 sg13g2_nand2_1 _1968_ (.Y(_0346_),
    .A(net84),
    .B(\u_top_module.u_cic.u_differentiator.count[2] ));
 sg13g2_nor2b_2 _1969_ (.A(net82),
    .B_N(net88),
    .Y(_0347_));
 sg13g2_nor2b_2 _1970_ (.A(net94),
    .B_N(net85),
    .Y(_0348_));
 sg13g2_nand2b_2 _1971_ (.Y(_0349_),
    .B(net83),
    .A_N(net90));
 sg13g2_xnor2_1 _1972_ (.Y(_0350_),
    .A(net89),
    .B(net83));
 sg13g2_nand2b_2 _1973_ (.Y(_0351_),
    .B(_0349_),
    .A_N(net76));
 sg13g2_nor2b_1 _1974_ (.A(\u_top_module.u_cic.u_differentiator.count[2] ),
    .B_N(net76),
    .Y(_0352_));
 sg13g2_nor2_2 _1975_ (.A(\u_top_module.u_cic.u_differentiator.count[2] ),
    .B(_0349_),
    .Y(_0353_));
 sg13g2_nand2b_2 _1976_ (.Y(_0354_),
    .B(_0348_),
    .A_N(\u_top_module.u_cic.u_differentiator.count[2] ));
 sg13g2_nor2_1 _1977_ (.A(\u_top_module.u_cic.u_differentiator.count[2] ),
    .B(net72),
    .Y(_0355_));
 sg13g2_nor2_2 _1978_ (.A(net69),
    .B(net66),
    .Y(_0356_));
 sg13g2_nor2b_2 _1979_ (.A(_0343_),
    .B_N(net68),
    .Y(_0357_));
 sg13g2_nor2_2 _1980_ (.A(_0344_),
    .B(_0349_),
    .Y(_0358_));
 sg13g2_a21oi_1 _1981_ (.A1(_0346_),
    .A2(net59),
    .Y(_0168_),
    .B1(_0343_));
 sg13g2_and2_1 _1982_ (.A(net92),
    .B(net84),
    .X(_0359_));
 sg13g2_nor2_1 _1983_ (.A(\u_top_module.u_cic.u_differentiator.count[2] ),
    .B(_0359_),
    .Y(_0360_));
 sg13g2_nor2_1 _1984_ (.A(_0343_),
    .B(_0360_),
    .Y(_0169_));
 sg13g2_nor2_1 _1985_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[0] ),
    .B(net57),
    .Y(_0361_));
 sg13g2_a22oi_1 _1986_ (.Y(_0362_),
    .B1(_0359_),
    .B2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[0] ),
    .A2(_0348_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[0] ));
 sg13g2_nand2_1 _1987_ (.Y(_0363_),
    .A(\u_top_module.u_cic.u_differentiator.temp[0] ),
    .B(_0362_));
 sg13g2_xor2_1 _1988_ (.B(_0362_),
    .A(\u_top_module.u_cic.u_differentiator.temp[0] ),
    .X(_0364_));
 sg13g2_a21oi_1 _1989_ (.A1(net57),
    .A2(_0364_),
    .Y(_0171_),
    .B1(_0361_));
 sg13g2_nor2_1 _1990_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[1] ),
    .B(net56),
    .Y(_0365_));
 sg13g2_nand2_1 _1991_ (.Y(_0366_),
    .A(net94),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[1] ));
 sg13g2_o21ai_1 _1992_ (.B1(net85),
    .Y(_0367_),
    .A1(net94),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[1] ));
 sg13g2_a22oi_1 _1993_ (.Y(_0368_),
    .B1(_0366_),
    .B2(_0367_),
    .A2(net73),
    .A1(_0699_));
 sg13g2_nor2b_1 _1994_ (.A(\u_top_module.u_cic.u_differentiator.temp[1] ),
    .B_N(_0368_),
    .Y(_0369_));
 sg13g2_xnor2_1 _1995_ (.Y(_0370_),
    .A(\u_top_module.u_cic.u_differentiator.temp[1] ),
    .B(_0368_));
 sg13g2_xnor2_1 _1996_ (.Y(_0371_),
    .A(_0363_),
    .B(_0370_));
 sg13g2_a21oi_1 _1997_ (.A1(net56),
    .A2(_0371_),
    .Y(_0172_),
    .B1(_0365_));
 sg13g2_nor2_1 _1998_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[2] ),
    .B(net55),
    .Y(_0372_));
 sg13g2_a21o_1 _1999_ (.A2(_0370_),
    .A1(_0363_),
    .B1(_0369_),
    .X(_0373_));
 sg13g2_nand2_1 _2000_ (.Y(_0374_),
    .A(net93),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[2] ));
 sg13g2_o21ai_1 _2001_ (.B1(net85),
    .Y(_0375_),
    .A1(net94),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[2] ));
 sg13g2_a22oi_1 _2002_ (.Y(_0376_),
    .B1(_0374_),
    .B2(_0375_),
    .A2(net73),
    .A1(_0701_));
 sg13g2_nor2b_1 _2003_ (.A(\u_top_module.u_cic.u_differentiator.temp[2] ),
    .B_N(_0376_),
    .Y(_0377_));
 sg13g2_xnor2_1 _2004_ (.Y(_0378_),
    .A(\u_top_module.u_cic.u_differentiator.temp[2] ),
    .B(_0376_));
 sg13g2_xnor2_1 _2005_ (.Y(_0379_),
    .A(_0373_),
    .B(_0378_));
 sg13g2_a21oi_1 _2006_ (.A1(net56),
    .A2(_0379_),
    .Y(_0173_),
    .B1(_0372_));
 sg13g2_nor2_1 _2007_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[3] ),
    .B(net56),
    .Y(_0380_));
 sg13g2_a21oi_2 _2008_ (.B1(_0377_),
    .Y(_0381_),
    .A2(_0378_),
    .A1(_0373_));
 sg13g2_nand2_1 _2009_ (.Y(_0382_),
    .A(net93),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[3] ));
 sg13g2_o21ai_1 _2010_ (.B1(net85),
    .Y(_0383_),
    .A1(net94),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[3] ));
 sg13g2_a22oi_1 _2011_ (.Y(_0384_),
    .B1(_0382_),
    .B2(_0383_),
    .A2(net73),
    .A1(_0702_));
 sg13g2_nand2b_1 _2012_ (.Y(_0385_),
    .B(_0384_),
    .A_N(\u_top_module.u_cic.u_differentiator.temp[3] ));
 sg13g2_xor2_1 _2013_ (.B(_0384_),
    .A(\u_top_module.u_cic.u_differentiator.temp[3] ),
    .X(_0386_));
 sg13g2_xnor2_1 _2014_ (.Y(_0387_),
    .A(_0381_),
    .B(_0386_));
 sg13g2_a21oi_1 _2015_ (.A1(net55),
    .A2(_0387_),
    .Y(_0174_),
    .B1(_0380_));
 sg13g2_nor2_1 _2016_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[4] ),
    .B(net55),
    .Y(_0388_));
 sg13g2_o21ai_1 _2017_ (.B1(_0385_),
    .Y(_0389_),
    .A1(_0381_),
    .A2(_0386_));
 sg13g2_nand2_1 _2018_ (.Y(_0390_),
    .A(net93),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[4] ));
 sg13g2_o21ai_1 _2019_ (.B1(net85),
    .Y(_0391_),
    .A1(net93),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[4] ));
 sg13g2_a22oi_1 _2020_ (.Y(_0392_),
    .B1(_0390_),
    .B2(_0391_),
    .A2(net73),
    .A1(_0704_));
 sg13g2_nor2b_1 _2021_ (.A(\u_top_module.u_cic.u_differentiator.temp[4] ),
    .B_N(_0392_),
    .Y(_0393_));
 sg13g2_xnor2_1 _2022_ (.Y(_0394_),
    .A(\u_top_module.u_cic.u_differentiator.temp[4] ),
    .B(_0392_));
 sg13g2_xnor2_1 _2023_ (.Y(_0395_),
    .A(_0389_),
    .B(_0394_));
 sg13g2_a21oi_1 _2024_ (.A1(net55),
    .A2(_0395_),
    .Y(_0175_),
    .B1(_0388_));
 sg13g2_nor2_1 _2025_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[5] ),
    .B(net55),
    .Y(_0396_));
 sg13g2_a21oi_1 _2026_ (.A1(_0389_),
    .A2(_0394_),
    .Y(_0397_),
    .B1(_0393_));
 sg13g2_nand2_1 _2027_ (.Y(_0398_),
    .A(net93),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[5] ));
 sg13g2_o21ai_1 _2028_ (.B1(net85),
    .Y(_0399_),
    .A1(net93),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[5] ));
 sg13g2_a22oi_1 _2029_ (.Y(_0400_),
    .B1(_0398_),
    .B2(_0399_),
    .A2(net72),
    .A1(_0705_));
 sg13g2_nand2b_1 _2030_ (.Y(_0401_),
    .B(_0400_),
    .A_N(\u_top_module.u_cic.u_differentiator.temp[5] ));
 sg13g2_xor2_1 _2031_ (.B(_0400_),
    .A(\u_top_module.u_cic.u_differentiator.temp[5] ),
    .X(_0402_));
 sg13g2_xnor2_1 _2032_ (.Y(_0403_),
    .A(_0397_),
    .B(_0402_));
 sg13g2_a21oi_1 _2033_ (.A1(net55),
    .A2(_0403_),
    .Y(_0176_),
    .B1(_0396_));
 sg13g2_nor2_1 _2034_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[6] ),
    .B(net55),
    .Y(_0404_));
 sg13g2_o21ai_1 _2035_ (.B1(_0401_),
    .Y(_0405_),
    .A1(_0397_),
    .A2(_0402_));
 sg13g2_nand2_1 _2036_ (.Y(_0406_),
    .A(net93),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[6] ));
 sg13g2_o21ai_1 _2037_ (.B1(net85),
    .Y(_0407_),
    .A1(net93),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[6] ));
 sg13g2_a22oi_1 _2038_ (.Y(_0408_),
    .B1(_0406_),
    .B2(_0407_),
    .A2(net72),
    .A1(_0707_));
 sg13g2_nor2b_1 _2039_ (.A(\u_top_module.u_cic.u_differentiator.temp[6] ),
    .B_N(_0408_),
    .Y(_0409_));
 sg13g2_xnor2_1 _2040_ (.Y(_0410_),
    .A(\u_top_module.u_cic.u_differentiator.temp[6] ),
    .B(_0408_));
 sg13g2_xnor2_1 _2041_ (.Y(_0411_),
    .A(_0405_),
    .B(_0410_));
 sg13g2_a21oi_1 _2042_ (.A1(net55),
    .A2(_0411_),
    .Y(_0177_),
    .B1(_0404_));
 sg13g2_nor2_1 _2043_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[7] ),
    .B(net56),
    .Y(_0412_));
 sg13g2_a21oi_2 _2044_ (.B1(_0409_),
    .Y(_0413_),
    .A2(_0410_),
    .A1(_0405_));
 sg13g2_nand2_1 _2045_ (.Y(_0414_),
    .A(net94),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[7] ));
 sg13g2_o21ai_1 _2046_ (.B1(net84),
    .Y(_0415_),
    .A1(net94),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[7] ));
 sg13g2_a22oi_1 _2047_ (.Y(_0416_),
    .B1(_0414_),
    .B2(_0415_),
    .A2(net72),
    .A1(_0708_));
 sg13g2_nand2b_1 _2048_ (.Y(_0417_),
    .B(_0416_),
    .A_N(\u_top_module.u_cic.u_differentiator.temp[7] ));
 sg13g2_xor2_1 _2049_ (.B(_0416_),
    .A(\u_top_module.u_cic.u_differentiator.temp[7] ),
    .X(_0418_));
 sg13g2_xnor2_1 _2050_ (.Y(_0419_),
    .A(_0413_),
    .B(_0418_));
 sg13g2_a21oi_1 _2051_ (.A1(net56),
    .A2(_0419_),
    .Y(_0178_),
    .B1(_0412_));
 sg13g2_nor2_1 _2052_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[8] ),
    .B(net54),
    .Y(_0420_));
 sg13g2_o21ai_1 _2053_ (.B1(_0417_),
    .Y(_0421_),
    .A1(_0413_),
    .A2(_0418_));
 sg13g2_nand2_1 _2054_ (.Y(_0422_),
    .A(net91),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[8] ));
 sg13g2_o21ai_1 _2055_ (.B1(net84),
    .Y(_0423_),
    .A1(net92),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[8] ));
 sg13g2_a22oi_1 _2056_ (.Y(_0424_),
    .B1(_0422_),
    .B2(_0423_),
    .A2(net72),
    .A1(_0710_));
 sg13g2_nor2b_1 _2057_ (.A(\u_top_module.u_cic.u_differentiator.temp[8] ),
    .B_N(_0424_),
    .Y(_0425_));
 sg13g2_xnor2_1 _2058_ (.Y(_0426_),
    .A(\u_top_module.u_cic.u_differentiator.temp[8] ),
    .B(_0424_));
 sg13g2_xnor2_1 _2059_ (.Y(_0427_),
    .A(_0421_),
    .B(_0426_));
 sg13g2_a21oi_1 _2060_ (.A1(net54),
    .A2(_0427_),
    .Y(_0179_),
    .B1(_0420_));
 sg13g2_nor2_1 _2061_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[9] ),
    .B(net54),
    .Y(_0428_));
 sg13g2_a21oi_1 _2062_ (.A1(_0421_),
    .A2(_0426_),
    .Y(_0429_),
    .B1(_0425_));
 sg13g2_nand2_1 _2063_ (.Y(_0430_),
    .A(net91),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[9] ));
 sg13g2_o21ai_1 _2064_ (.B1(net84),
    .Y(_0431_),
    .A1(net91),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[9] ));
 sg13g2_a22oi_1 _2065_ (.Y(_0432_),
    .B1(_0430_),
    .B2(_0431_),
    .A2(net72),
    .A1(_0711_));
 sg13g2_nor2_1 _2066_ (.A(_0734_),
    .B(_0432_),
    .Y(_0433_));
 sg13g2_xnor2_1 _2067_ (.Y(_0434_),
    .A(_0734_),
    .B(_0432_));
 sg13g2_xnor2_1 _2068_ (.Y(_0435_),
    .A(_0429_),
    .B(_0434_));
 sg13g2_a21oi_1 _2069_ (.A1(net54),
    .A2(_0435_),
    .Y(_0180_),
    .B1(_0428_));
 sg13g2_nor2_1 _2070_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[10] ),
    .B(net54),
    .Y(_0436_));
 sg13g2_nand2_1 _2071_ (.Y(_0437_),
    .A(net91),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[10] ));
 sg13g2_o21ai_1 _2072_ (.B1(net84),
    .Y(_0438_),
    .A1(net91),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[10] ));
 sg13g2_a22oi_1 _2073_ (.Y(_0439_),
    .B1(_0437_),
    .B2(_0438_),
    .A2(net72),
    .A1(_0713_));
 sg13g2_nor2b_1 _2074_ (.A(\u_top_module.u_cic.u_differentiator.temp[10] ),
    .B_N(_0439_),
    .Y(_0440_));
 sg13g2_xnor2_1 _2075_ (.Y(_0441_),
    .A(\u_top_module.u_cic.u_differentiator.temp[10] ),
    .B(_0439_));
 sg13g2_a221oi_1 _2076_ (.B2(_0734_),
    .C1(_0425_),
    .B1(_0432_),
    .A1(_0421_),
    .Y(_0442_),
    .A2(_0426_));
 sg13g2_nor2_1 _2077_ (.A(_0433_),
    .B(_0442_),
    .Y(_0443_));
 sg13g2_xnor2_1 _2078_ (.Y(_0444_),
    .A(_0441_),
    .B(_0443_));
 sg13g2_a21oi_1 _2079_ (.A1(net54),
    .A2(_0444_),
    .Y(_0181_),
    .B1(_0436_));
 sg13g2_nor2_1 _2080_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[11] ),
    .B(net54),
    .Y(_0445_));
 sg13g2_nand2_1 _2081_ (.Y(_0446_),
    .A(net91),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[11] ));
 sg13g2_o21ai_1 _2082_ (.B1(net84),
    .Y(_0447_),
    .A1(net91),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[11] ));
 sg13g2_a22oi_1 _2083_ (.Y(_0448_),
    .B1(_0446_),
    .B2(_0447_),
    .A2(net72),
    .A1(_0714_));
 sg13g2_nor2b_1 _2084_ (.A(\u_top_module.u_cic.u_differentiator.temp[11] ),
    .B_N(_0448_),
    .Y(_0449_));
 sg13g2_nand2b_1 _2085_ (.Y(_0450_),
    .B(\u_top_module.u_cic.u_differentiator.temp[11] ),
    .A_N(_0448_));
 sg13g2_nor2b_1 _2086_ (.A(_0449_),
    .B_N(_0450_),
    .Y(_0451_));
 sg13g2_a21oi_1 _2087_ (.A1(_0441_),
    .A2(_0443_),
    .Y(_0452_),
    .B1(_0440_));
 sg13g2_xor2_1 _2088_ (.B(_0452_),
    .A(_0451_),
    .X(_0453_));
 sg13g2_a21oi_1 _2089_ (.A1(net54),
    .A2(_0453_),
    .Y(_0182_),
    .B1(_0445_));
 sg13g2_nor2_1 _2090_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[12] ),
    .B(net51),
    .Y(_0454_));
 sg13g2_nand2_1 _2091_ (.Y(_0455_),
    .A(net90),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[12] ));
 sg13g2_o21ai_1 _2092_ (.B1(net83),
    .Y(_0456_),
    .A1(net89),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[12] ));
 sg13g2_a22oi_1 _2093_ (.Y(_0457_),
    .B1(_0455_),
    .B2(_0456_),
    .A2(net71),
    .A1(_0716_));
 sg13g2_nor2b_1 _2094_ (.A(\u_top_module.u_cic.u_differentiator.temp[12] ),
    .B_N(_0457_),
    .Y(_0458_));
 sg13g2_xnor2_1 _2095_ (.Y(_0459_),
    .A(\u_top_module.u_cic.u_differentiator.temp[12] ),
    .B(_0457_));
 sg13g2_and2_1 _2096_ (.A(_0440_),
    .B(_0450_),
    .X(_0460_));
 sg13g2_nand2_1 _2097_ (.Y(_0461_),
    .A(_0441_),
    .B(_0451_));
 sg13g2_nor3_1 _2098_ (.A(_0433_),
    .B(_0442_),
    .C(_0461_),
    .Y(_0462_));
 sg13g2_or3_1 _2099_ (.A(_0449_),
    .B(_0460_),
    .C(_0462_),
    .X(_0463_));
 sg13g2_xnor2_1 _2100_ (.Y(_0464_),
    .A(_0459_),
    .B(_0463_));
 sg13g2_a21oi_1 _2101_ (.A1(net52),
    .A2(_0464_),
    .Y(_0183_),
    .B1(_0454_));
 sg13g2_nor2_1 _2102_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[13] ),
    .B(net51),
    .Y(_0465_));
 sg13g2_or2_1 _2103_ (.X(_0466_),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[13] ),
    .A(net90));
 sg13g2_a21oi_1 _2104_ (.A1(net90),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[13] ),
    .Y(_0467_),
    .B1(net83));
 sg13g2_o21ai_1 _2105_ (.B1(_0466_),
    .Y(_0468_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[13] ),
    .A2(_0351_));
 sg13g2_nor3_1 _2106_ (.A(\u_top_module.u_cic.u_differentiator.temp[13] ),
    .B(_0467_),
    .C(_0468_),
    .Y(_0469_));
 sg13g2_o21ai_1 _2107_ (.B1(\u_top_module.u_cic.u_differentiator.temp[13] ),
    .Y(_0470_),
    .A1(_0467_),
    .A2(_0468_));
 sg13g2_nor2b_1 _2108_ (.A(_0469_),
    .B_N(_0470_),
    .Y(_0471_));
 sg13g2_a21o_1 _2109_ (.A2(_0463_),
    .A1(_0459_),
    .B1(_0458_),
    .X(_0472_));
 sg13g2_xnor2_1 _2110_ (.Y(_0473_),
    .A(_0471_),
    .B(_0472_));
 sg13g2_a21oi_1 _2111_ (.A1(net52),
    .A2(_0473_),
    .Y(_0184_),
    .B1(_0465_));
 sg13g2_nor2_1 _2112_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[14] ),
    .B(net52),
    .Y(_0474_));
 sg13g2_nand2_1 _2113_ (.Y(_0475_),
    .A(net89),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[14] ));
 sg13g2_o21ai_1 _2114_ (.B1(net83),
    .Y(_0476_),
    .A1(net89),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[14] ));
 sg13g2_a22oi_1 _2115_ (.Y(_0477_),
    .B1(_0475_),
    .B2(_0476_),
    .A2(net74),
    .A1(_0718_));
 sg13g2_nor2b_1 _2116_ (.A(\u_top_module.u_cic.u_differentiator.temp[14] ),
    .B_N(_0477_),
    .Y(_0478_));
 sg13g2_xnor2_1 _2117_ (.Y(_0479_),
    .A(\u_top_module.u_cic.u_differentiator.temp[14] ),
    .B(_0477_));
 sg13g2_and2_1 _2118_ (.A(_0459_),
    .B(_0471_),
    .X(_0480_));
 sg13g2_a221oi_1 _2119_ (.B2(_0463_),
    .C1(_0469_),
    .B1(_0480_),
    .A1(_0458_),
    .Y(_0481_),
    .A2(_0470_));
 sg13g2_nor2b_1 _2120_ (.A(_0481_),
    .B_N(_0479_),
    .Y(_0482_));
 sg13g2_xor2_1 _2121_ (.B(_0481_),
    .A(_0479_),
    .X(_0483_));
 sg13g2_a21oi_1 _2122_ (.A1(net52),
    .A2(_0483_),
    .Y(_0185_),
    .B1(_0474_));
 sg13g2_nor2_1 _2123_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[15] ),
    .B(net51),
    .Y(_0484_));
 sg13g2_or2_1 _2124_ (.X(_0485_),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[15] ),
    .A(net89));
 sg13g2_a21oi_1 _2125_ (.A1(net89),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[15] ),
    .Y(_0486_),
    .B1(net83));
 sg13g2_o21ai_1 _2126_ (.B1(_0485_),
    .Y(_0487_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[15] ),
    .A2(_0351_));
 sg13g2_nor3_1 _2127_ (.A(\u_top_module.u_cic.u_differentiator.temp[15] ),
    .B(_0486_),
    .C(_0487_),
    .Y(_0488_));
 sg13g2_o21ai_1 _2128_ (.B1(\u_top_module.u_cic.u_differentiator.temp[15] ),
    .Y(_0489_),
    .A1(_0486_),
    .A2(_0487_));
 sg13g2_nor2b_1 _2129_ (.A(_0488_),
    .B_N(_0489_),
    .Y(_0490_));
 sg13g2_nor2_1 _2130_ (.A(_0478_),
    .B(_0482_),
    .Y(_0491_));
 sg13g2_xor2_1 _2131_ (.B(_0491_),
    .A(_0490_),
    .X(_0492_));
 sg13g2_a21oi_1 _2132_ (.A1(net51),
    .A2(_0492_),
    .Y(_0186_),
    .B1(_0484_));
 sg13g2_nor2_1 _2133_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[16] ),
    .B(net50),
    .Y(_0493_));
 sg13g2_nand2_1 _2134_ (.Y(_0494_),
    .A(net88),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[16] ));
 sg13g2_o21ai_1 _2135_ (.B1(net82),
    .Y(_0495_),
    .A1(net87),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[16] ));
 sg13g2_a22oi_1 _2136_ (.Y(_0496_),
    .B1(_0494_),
    .B2(_0495_),
    .A2(net71),
    .A1(_0720_));
 sg13g2_nor2b_1 _2137_ (.A(\u_top_module.u_cic.u_differentiator.temp[16] ),
    .B_N(_0496_),
    .Y(_0497_));
 sg13g2_xnor2_1 _2138_ (.Y(_0498_),
    .A(\u_top_module.u_cic.u_differentiator.temp[16] ),
    .B(_0496_));
 sg13g2_nand2_1 _2139_ (.Y(_0499_),
    .A(_0479_),
    .B(_0490_));
 sg13g2_a21oi_1 _2140_ (.A1(_0478_),
    .A2(_0489_),
    .Y(_0500_),
    .B1(_0488_));
 sg13g2_o21ai_1 _2141_ (.B1(_0500_),
    .Y(_0501_),
    .A1(_0481_),
    .A2(_0499_));
 sg13g2_nand2_1 _2142_ (.Y(_0502_),
    .A(_0498_),
    .B(_0501_));
 sg13g2_xnor2_1 _2143_ (.Y(_0503_),
    .A(_0498_),
    .B(_0501_));
 sg13g2_a21oi_1 _2144_ (.A1(net50),
    .A2(_0503_),
    .Y(_0187_),
    .B1(_0493_));
 sg13g2_nor2_1 _2145_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[17] ),
    .B(net51),
    .Y(_0504_));
 sg13g2_nand2_1 _2146_ (.Y(_0505_),
    .A(net88),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[17] ));
 sg13g2_o21ai_1 _2147_ (.B1(net82),
    .Y(_0506_),
    .A1(net88),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[17] ));
 sg13g2_a22oi_1 _2148_ (.Y(_0507_),
    .B1(_0505_),
    .B2(_0506_),
    .A2(net71),
    .A1(_0721_));
 sg13g2_nor2_1 _2149_ (.A(_0735_),
    .B(_0507_),
    .Y(_0508_));
 sg13g2_xnor2_1 _2150_ (.Y(_0509_),
    .A(_0735_),
    .B(_0507_));
 sg13g2_a21oi_1 _2151_ (.A1(_0498_),
    .A2(_0501_),
    .Y(_0510_),
    .B1(_0497_));
 sg13g2_xnor2_1 _2152_ (.Y(_0511_),
    .A(_0509_),
    .B(_0510_));
 sg13g2_a21oi_1 _2153_ (.A1(net51),
    .A2(_0511_),
    .Y(_0188_),
    .B1(_0504_));
 sg13g2_nor2_1 _2154_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[18] ),
    .B(net49),
    .Y(_0512_));
 sg13g2_a21oi_1 _2155_ (.A1(_0735_),
    .A2(_0507_),
    .Y(_0513_),
    .B1(_0497_));
 sg13g2_a21oi_2 _2156_ (.B1(_0508_),
    .Y(_0514_),
    .A2(_0513_),
    .A1(_0502_));
 sg13g2_nand2_1 _2157_ (.Y(_0515_),
    .A(net88),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[18] ));
 sg13g2_o21ai_1 _2158_ (.B1(net82),
    .Y(_0516_),
    .A1(net88),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[18] ));
 sg13g2_a22oi_1 _2159_ (.Y(_0517_),
    .B1(_0515_),
    .B2(_0516_),
    .A2(net71),
    .A1(_0723_));
 sg13g2_nor2b_1 _2160_ (.A(\u_top_module.u_cic.u_differentiator.temp[18] ),
    .B_N(_0517_),
    .Y(_0518_));
 sg13g2_xnor2_1 _2161_ (.Y(_0519_),
    .A(\u_top_module.u_cic.u_differentiator.temp[18] ),
    .B(_0517_));
 sg13g2_xnor2_1 _2162_ (.Y(_0520_),
    .A(_0514_),
    .B(_0519_));
 sg13g2_a21oi_1 _2163_ (.A1(net49),
    .A2(_0520_),
    .Y(_0189_),
    .B1(_0512_));
 sg13g2_nor2_1 _2164_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[19] ),
    .B(net50),
    .Y(_0521_));
 sg13g2_or2_1 _2165_ (.X(_0522_),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[19] ),
    .A(net87));
 sg13g2_a21oi_1 _2166_ (.A1(net87),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[19] ),
    .Y(_0523_),
    .B1(net82));
 sg13g2_o21ai_1 _2167_ (.B1(_0522_),
    .Y(_0524_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[19] ),
    .A2(_0351_));
 sg13g2_nor3_1 _2168_ (.A(\u_top_module.u_cic.u_differentiator.temp[19] ),
    .B(_0523_),
    .C(_0524_),
    .Y(_0525_));
 sg13g2_o21ai_1 _2169_ (.B1(\u_top_module.u_cic.u_differentiator.temp[19] ),
    .Y(_0526_),
    .A1(_0523_),
    .A2(_0524_));
 sg13g2_nor2b_1 _2170_ (.A(_0525_),
    .B_N(_0526_),
    .Y(_0527_));
 sg13g2_a21oi_1 _2171_ (.A1(_0514_),
    .A2(_0519_),
    .Y(_0528_),
    .B1(_0518_));
 sg13g2_xor2_1 _2172_ (.B(_0528_),
    .A(_0527_),
    .X(_0529_));
 sg13g2_a21oi_1 _2173_ (.A1(net50),
    .A2(_0529_),
    .Y(_0190_),
    .B1(_0521_));
 sg13g2_nor2_1 _2174_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[20] ),
    .B(net49),
    .Y(_0530_));
 sg13g2_nand2_1 _2175_ (.Y(_0531_),
    .A(net87),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[20] ));
 sg13g2_o21ai_1 _2176_ (.B1(net82),
    .Y(_0532_),
    .A1(net88),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[20] ));
 sg13g2_a22oi_1 _2177_ (.Y(_0533_),
    .B1(_0531_),
    .B2(_0532_),
    .A2(net71),
    .A1(_0725_));
 sg13g2_nor2b_1 _2178_ (.A(\u_top_module.u_cic.u_differentiator.temp[20] ),
    .B_N(_0533_),
    .Y(_0534_));
 sg13g2_inv_1 _2179_ (.Y(_0535_),
    .A(_0534_));
 sg13g2_xnor2_1 _2180_ (.Y(_0536_),
    .A(\u_top_module.u_cic.u_differentiator.temp[20] ),
    .B(_0533_));
 sg13g2_inv_1 _2181_ (.Y(_0537_),
    .A(_0536_));
 sg13g2_and2_1 _2182_ (.A(_0519_),
    .B(_0527_),
    .X(_0538_));
 sg13g2_a221oi_1 _2183_ (.B2(_0514_),
    .C1(_0525_),
    .B1(_0538_),
    .A1(_0518_),
    .Y(_0539_),
    .A2(_0526_));
 sg13g2_xnor2_1 _2184_ (.Y(_0540_),
    .A(_0537_),
    .B(_0539_));
 sg13g2_a21oi_1 _2185_ (.A1(net49),
    .A2(_0540_),
    .Y(_0191_),
    .B1(_0530_));
 sg13g2_nor2_1 _2186_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[21] ),
    .B(net49),
    .Y(_0541_));
 sg13g2_o21ai_1 _2187_ (.B1(_0535_),
    .Y(_0542_),
    .A1(_0537_),
    .A2(_0539_));
 sg13g2_nand2_1 _2188_ (.Y(_0543_),
    .A(net87),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[21] ));
 sg13g2_o21ai_1 _2189_ (.B1(net82),
    .Y(_0544_),
    .A1(net87),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[21] ));
 sg13g2_a22oi_1 _2190_ (.Y(_0545_),
    .B1(_0543_),
    .B2(_0544_),
    .A2(net71),
    .A1(_0726_));
 sg13g2_nand2b_1 _2191_ (.Y(_0546_),
    .B(\u_top_module.u_cic.u_differentiator.temp[21] ),
    .A_N(_0545_));
 sg13g2_nor2b_1 _2192_ (.A(\u_top_module.u_cic.u_differentiator.temp[21] ),
    .B_N(_0545_),
    .Y(_0547_));
 sg13g2_xnor2_1 _2193_ (.Y(_0548_),
    .A(\u_top_module.u_cic.u_differentiator.temp[21] ),
    .B(_0545_));
 sg13g2_xnor2_1 _2194_ (.Y(_0549_),
    .A(_0542_),
    .B(_0548_));
 sg13g2_a21oi_1 _2195_ (.A1(net49),
    .A2(_0549_),
    .Y(_0192_),
    .B1(_0541_));
 sg13g2_nor2_1 _2196_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[22] ),
    .B(net49),
    .Y(_0550_));
 sg13g2_nand2_1 _2197_ (.Y(_0551_),
    .A(net87),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[22] ));
 sg13g2_o21ai_1 _2198_ (.B1(net82),
    .Y(_0552_),
    .A1(net87),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[22] ));
 sg13g2_a22oi_1 _2199_ (.Y(_0553_),
    .B1(_0551_),
    .B2(_0552_),
    .A2(net71),
    .A1(_0727_));
 sg13g2_nor2b_1 _2200_ (.A(\u_top_module.u_cic.u_differentiator.temp[22] ),
    .B_N(_0553_),
    .Y(_0554_));
 sg13g2_xnor2_1 _2201_ (.Y(_0555_),
    .A(\u_top_module.u_cic.u_differentiator.temp[22] ),
    .B(_0553_));
 sg13g2_a21o_1 _2202_ (.A2(_0546_),
    .A1(_0542_),
    .B1(_0547_),
    .X(_0556_));
 sg13g2_xnor2_1 _2203_ (.Y(_0557_),
    .A(_0555_),
    .B(_0556_));
 sg13g2_a21oi_1 _2204_ (.A1(net49),
    .A2(_0557_),
    .Y(_0193_),
    .B1(_0550_));
 sg13g2_nor2_1 _2205_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[23] ),
    .B(net51),
    .Y(_0558_));
 sg13g2_a21oi_1 _2206_ (.A1(_0555_),
    .A2(_0556_),
    .Y(_0559_),
    .B1(_0554_));
 sg13g2_nand2_1 _2207_ (.Y(_0560_),
    .A(net89),
    .B(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[23] ));
 sg13g2_o21ai_1 _2208_ (.B1(net83),
    .Y(_0561_),
    .A1(net89),
    .A2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[23] ));
 sg13g2_a22oi_1 _2209_ (.Y(_0562_),
    .B1(_0560_),
    .B2(_0561_),
    .A2(net71),
    .A1(_0728_));
 sg13g2_xnor2_1 _2210_ (.Y(_0563_),
    .A(\u_top_module.u_cic.u_differentiator.temp[23] ),
    .B(_0562_));
 sg13g2_xor2_1 _2211_ (.B(_0563_),
    .A(_0559_),
    .X(_0564_));
 sg13g2_a21oi_1 _2212_ (.A1(net51),
    .A2(_0564_),
    .Y(_0194_),
    .B1(_0558_));
 sg13g2_nor2_1 _2213_ (.A(_0344_),
    .B(_0359_),
    .Y(_0565_));
 sg13g2_or2_1 _2214_ (.X(_0566_),
    .B(_0359_),
    .A(_0344_));
 sg13g2_a22oi_1 _2215_ (.Y(_0567_),
    .B1(net67),
    .B2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[0] ),
    .A2(net68),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[0] ));
 sg13g2_nor2_1 _2216_ (.A(\u_top_module.u_cic.u_differentiator.temp[0] ),
    .B(net37),
    .Y(_0568_));
 sg13g2_a21oi_1 _2217_ (.A1(net37),
    .A2(_0567_),
    .Y(_0195_),
    .B1(_0568_));
 sg13g2_o21ai_1 _2218_ (.B1(net62),
    .Y(_0569_),
    .A1(_0036_),
    .A2(_0349_));
 sg13g2_a21oi_1 _2219_ (.A1(_0700_),
    .A2(net69),
    .Y(_0570_),
    .B1(_0569_));
 sg13g2_o21ai_1 _2220_ (.B1(net38),
    .Y(_0571_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[1] ),
    .A2(net62));
 sg13g2_nand2_1 _2221_ (.Y(_0572_),
    .A(\u_top_module.u_cic.u_differentiator.temp[1] ),
    .B(net34));
 sg13g2_o21ai_1 _2222_ (.B1(_0572_),
    .Y(_0196_),
    .A1(_0570_),
    .A2(_0571_));
 sg13g2_a221oi_1 _2223_ (.B2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[2] ),
    .C1(net59),
    .B1(net68),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[2] ),
    .Y(_0573_),
    .A2(_0348_));
 sg13g2_o21ai_1 _2224_ (.B1(net38),
    .Y(_0574_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[2] ),
    .A2(net64));
 sg13g2_nand2_1 _2225_ (.Y(_0575_),
    .A(\u_top_module.u_cic.u_differentiator.temp[2] ),
    .B(net34));
 sg13g2_o21ai_1 _2226_ (.B1(_0575_),
    .Y(_0197_),
    .A1(_0573_),
    .A2(_0574_));
 sg13g2_o21ai_1 _2227_ (.B1(net63),
    .Y(_0576_),
    .A1(_0038_),
    .A2(_0354_));
 sg13g2_a21oi_1 _2228_ (.A1(_0703_),
    .A2(net68),
    .Y(_0577_),
    .B1(_0576_));
 sg13g2_o21ai_1 _2229_ (.B1(net38),
    .Y(_0578_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[3] ),
    .A2(net62));
 sg13g2_nand2_1 _2230_ (.Y(_0579_),
    .A(\u_top_module.u_cic.u_differentiator.temp[3] ),
    .B(net34));
 sg13g2_o21ai_1 _2231_ (.B1(_0579_),
    .Y(_0198_),
    .A1(_0577_),
    .A2(_0578_));
 sg13g2_a221oi_1 _2232_ (.B2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[4] ),
    .C1(net59),
    .B1(net67),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[4] ),
    .Y(_0580_),
    .A2(net76));
 sg13g2_o21ai_1 _2233_ (.B1(net38),
    .Y(_0581_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[4] ),
    .A2(net62));
 sg13g2_nand2_1 _2234_ (.Y(_0582_),
    .A(\u_top_module.u_cic.u_differentiator.temp[4] ),
    .B(net33));
 sg13g2_o21ai_1 _2235_ (.B1(_0582_),
    .Y(_0199_),
    .A1(_0580_),
    .A2(_0581_));
 sg13g2_o21ai_1 _2236_ (.B1(net64),
    .Y(_0583_),
    .A1(_0040_),
    .A2(net65));
 sg13g2_a21oi_1 _2237_ (.A1(_0706_),
    .A2(net68),
    .Y(_0584_),
    .B1(_0583_));
 sg13g2_o21ai_1 _2238_ (.B1(net38),
    .Y(_0585_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[5] ),
    .A2(net62));
 sg13g2_nand2_1 _2239_ (.Y(_0586_),
    .A(\u_top_module.u_cic.u_differentiator.temp[5] ),
    .B(net33));
 sg13g2_o21ai_1 _2240_ (.B1(_0586_),
    .Y(_0200_),
    .A1(_0584_),
    .A2(_0585_));
 sg13g2_a221oi_1 _2241_ (.B2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[6] ),
    .C1(net59),
    .B1(net67),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[6] ),
    .Y(_0587_),
    .A2(net76));
 sg13g2_o21ai_1 _2242_ (.B1(net37),
    .Y(_0588_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[6] ),
    .A2(net62));
 sg13g2_nand2_1 _2243_ (.Y(_0589_),
    .A(\u_top_module.u_cic.u_differentiator.temp[6] ),
    .B(net33));
 sg13g2_o21ai_1 _2244_ (.B1(_0589_),
    .Y(_0201_),
    .A1(_0587_),
    .A2(_0588_));
 sg13g2_o21ai_1 _2245_ (.B1(net62),
    .Y(_0590_),
    .A1(_0042_),
    .A2(net65));
 sg13g2_a21oi_1 _2246_ (.A1(_0709_),
    .A2(net68),
    .Y(_0591_),
    .B1(_0590_));
 sg13g2_o21ai_1 _2247_ (.B1(net37),
    .Y(_0592_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[7] ),
    .A2(net62));
 sg13g2_nand2_1 _2248_ (.Y(_0593_),
    .A(\u_top_module.u_cic.u_differentiator.temp[7] ),
    .B(net33));
 sg13g2_o21ai_1 _2249_ (.B1(_0593_),
    .Y(_0202_),
    .A1(_0591_),
    .A2(_0592_));
 sg13g2_a221oi_1 _2250_ (.B2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[8] ),
    .C1(net58),
    .B1(net67),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[8] ),
    .Y(_0594_),
    .A2(net76));
 sg13g2_o21ai_1 _2251_ (.B1(net37),
    .Y(_0595_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[8] ),
    .A2(net63));
 sg13g2_nand2_1 _2252_ (.Y(_0596_),
    .A(\u_top_module.u_cic.u_differentiator.temp[8] ),
    .B(net33));
 sg13g2_o21ai_1 _2253_ (.B1(_0596_),
    .Y(_0203_),
    .A1(_0594_),
    .A2(_0595_));
 sg13g2_o21ai_1 _2254_ (.B1(net63),
    .Y(_0597_),
    .A1(_0044_),
    .A2(net65));
 sg13g2_a21oi_1 _2255_ (.A1(_0712_),
    .A2(net68),
    .Y(_0598_),
    .B1(_0597_));
 sg13g2_o21ai_1 _2256_ (.B1(net37),
    .Y(_0599_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[9] ),
    .A2(net63));
 sg13g2_nand2_1 _2257_ (.Y(_0600_),
    .A(\u_top_module.u_cic.u_differentiator.temp[9] ),
    .B(net33));
 sg13g2_o21ai_1 _2258_ (.B1(_0600_),
    .Y(_0204_),
    .A1(_0598_),
    .A2(_0599_));
 sg13g2_a221oi_1 _2259_ (.B2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[10] ),
    .C1(net59),
    .B1(net67),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[10] ),
    .Y(_0601_),
    .A2(net75));
 sg13g2_o21ai_1 _2260_ (.B1(net37),
    .Y(_0602_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[10] ),
    .A2(net63));
 sg13g2_nand2_1 _2261_ (.Y(_0603_),
    .A(\u_top_module.u_cic.u_differentiator.temp[10] ),
    .B(net33));
 sg13g2_o21ai_1 _2262_ (.B1(_0603_),
    .Y(_0205_),
    .A1(_0601_),
    .A2(_0602_));
 sg13g2_o21ai_1 _2263_ (.B1(net63),
    .Y(_0604_),
    .A1(_0046_),
    .A2(net65));
 sg13g2_a21oi_1 _2264_ (.A1(_0715_),
    .A2(net68),
    .Y(_0605_),
    .B1(_0604_));
 sg13g2_o21ai_1 _2265_ (.B1(net37),
    .Y(_0606_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[11] ),
    .A2(net63));
 sg13g2_nand2_1 _2266_ (.Y(_0607_),
    .A(\u_top_module.u_cic.u_differentiator.temp[11] ),
    .B(net33));
 sg13g2_o21ai_1 _2267_ (.B1(_0607_),
    .Y(_0206_),
    .A1(_0605_),
    .A2(_0606_));
 sg13g2_a221oi_1 _2268_ (.B2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[12] ),
    .C1(net59),
    .B1(net67),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[12] ),
    .Y(_0608_),
    .A2(net76));
 sg13g2_o21ai_1 _2269_ (.B1(net36),
    .Y(_0609_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[12] ),
    .A2(net64));
 sg13g2_nand2_1 _2270_ (.Y(_0610_),
    .A(\u_top_module.u_cic.u_differentiator.temp[12] ),
    .B(net32));
 sg13g2_o21ai_1 _2271_ (.B1(_0610_),
    .Y(_0207_),
    .A1(_0608_),
    .A2(_0609_));
 sg13g2_o21ai_1 _2272_ (.B1(net61),
    .Y(_0611_),
    .A1(_0048_),
    .A2(net65));
 sg13g2_a21oi_1 _2273_ (.A1(_0717_),
    .A2(net69),
    .Y(_0612_),
    .B1(_0611_));
 sg13g2_o21ai_1 _2274_ (.B1(net36),
    .Y(_0613_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[13] ),
    .A2(net61));
 sg13g2_nand2_1 _2275_ (.Y(_0614_),
    .A(\u_top_module.u_cic.u_differentiator.temp[13] ),
    .B(net31));
 sg13g2_o21ai_1 _2276_ (.B1(_0614_),
    .Y(_0208_),
    .A1(_0612_),
    .A2(_0613_));
 sg13g2_a221oi_1 _2277_ (.B2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[14] ),
    .C1(net58),
    .B1(net66),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[14] ),
    .Y(_0615_),
    .A2(net75));
 sg13g2_o21ai_1 _2278_ (.B1(net36),
    .Y(_0616_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[14] ),
    .A2(net61));
 sg13g2_nand2_1 _2279_ (.Y(_0617_),
    .A(\u_top_module.u_cic.u_differentiator.temp[14] ),
    .B(net32));
 sg13g2_o21ai_1 _2280_ (.B1(_0617_),
    .Y(_0209_),
    .A1(_0615_),
    .A2(_0616_));
 sg13g2_o21ai_1 _2281_ (.B1(net61),
    .Y(_0618_),
    .A1(_0050_),
    .A2(net65));
 sg13g2_a21oi_1 _2282_ (.A1(_0719_),
    .A2(net69),
    .Y(_0619_),
    .B1(_0618_));
 sg13g2_o21ai_1 _2283_ (.B1(net36),
    .Y(_0620_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[15] ),
    .A2(net61));
 sg13g2_nand2_1 _2284_ (.Y(_0621_),
    .A(\u_top_module.u_cic.u_differentiator.temp[15] ),
    .B(net32));
 sg13g2_o21ai_1 _2285_ (.B1(_0621_),
    .Y(_0210_),
    .A1(_0619_),
    .A2(_0620_));
 sg13g2_a221oi_1 _2286_ (.B2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[16] ),
    .C1(net58),
    .B1(net66),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[16] ),
    .Y(_0622_),
    .A2(net75));
 sg13g2_o21ai_1 _2287_ (.B1(net35),
    .Y(_0623_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[16] ),
    .A2(net61));
 sg13g2_nand2_1 _2288_ (.Y(_0624_),
    .A(\u_top_module.u_cic.u_differentiator.temp[16] ),
    .B(net31));
 sg13g2_o21ai_1 _2289_ (.B1(_0624_),
    .Y(_0211_),
    .A1(_0622_),
    .A2(_0623_));
 sg13g2_o21ai_1 _2290_ (.B1(net60),
    .Y(_0625_),
    .A1(_0052_),
    .A2(net65));
 sg13g2_a21oi_1 _2291_ (.A1(_0722_),
    .A2(net69),
    .Y(_0626_),
    .B1(_0625_));
 sg13g2_o21ai_1 _2292_ (.B1(net35),
    .Y(_0627_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[17] ),
    .A2(net60));
 sg13g2_nand2_1 _2293_ (.Y(_0628_),
    .A(\u_top_module.u_cic.u_differentiator.temp[17] ),
    .B(net31));
 sg13g2_o21ai_1 _2294_ (.B1(_0628_),
    .Y(_0212_),
    .A1(_0626_),
    .A2(_0627_));
 sg13g2_a221oi_1 _2295_ (.B2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[18] ),
    .C1(net58),
    .B1(net66),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[18] ),
    .Y(_0629_),
    .A2(net75));
 sg13g2_o21ai_1 _2296_ (.B1(net35),
    .Y(_0630_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[18] ),
    .A2(net60));
 sg13g2_nand2_1 _2297_ (.Y(_0631_),
    .A(\u_top_module.u_cic.u_differentiator.temp[18] ),
    .B(net31));
 sg13g2_o21ai_1 _2298_ (.B1(_0631_),
    .Y(_0213_),
    .A1(_0629_),
    .A2(_0630_));
 sg13g2_o21ai_1 _2299_ (.B1(net60),
    .Y(_0632_),
    .A1(_0054_),
    .A2(net65));
 sg13g2_a21oi_1 _2300_ (.A1(_0724_),
    .A2(net69),
    .Y(_0633_),
    .B1(_0632_));
 sg13g2_o21ai_1 _2301_ (.B1(net35),
    .Y(_0634_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[19] ),
    .A2(net60));
 sg13g2_nand2_1 _2302_ (.Y(_0635_),
    .A(\u_top_module.u_cic.u_differentiator.temp[19] ),
    .B(net31));
 sg13g2_o21ai_1 _2303_ (.B1(_0635_),
    .Y(_0214_),
    .A1(_0633_),
    .A2(_0634_));
 sg13g2_a221oi_1 _2304_ (.B2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[20] ),
    .C1(net58),
    .B1(net66),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[20] ),
    .Y(_0636_),
    .A2(net75));
 sg13g2_o21ai_1 _2305_ (.B1(net35),
    .Y(_0637_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[20] ),
    .A2(net60));
 sg13g2_nand2_1 _2306_ (.Y(_0638_),
    .A(\u_top_module.u_cic.u_differentiator.temp[20] ),
    .B(net31));
 sg13g2_o21ai_1 _2307_ (.B1(_0638_),
    .Y(_0215_),
    .A1(_0636_),
    .A2(_0637_));
 sg13g2_a221oi_1 _2308_ (.B2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[21] ),
    .C1(net58),
    .B1(net66),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[21] ),
    .Y(_0639_),
    .A2(net75));
 sg13g2_o21ai_1 _2309_ (.B1(net35),
    .Y(_0640_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[21] ),
    .A2(net60));
 sg13g2_nand2_1 _2310_ (.Y(_0641_),
    .A(\u_top_module.u_cic.u_differentiator.temp[21] ),
    .B(net31));
 sg13g2_o21ai_1 _2311_ (.B1(_0641_),
    .Y(_0216_),
    .A1(_0639_),
    .A2(_0640_));
 sg13g2_a221oi_1 _2312_ (.B2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[22] ),
    .C1(net58),
    .B1(net66),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[22] ),
    .Y(_0642_),
    .A2(net75));
 sg13g2_o21ai_1 _2313_ (.B1(net35),
    .Y(_0643_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[22] ),
    .A2(net60));
 sg13g2_nand2_1 _2314_ (.Y(_0644_),
    .A(\u_top_module.u_cic.u_differentiator.temp[22] ),
    .B(net31));
 sg13g2_o21ai_1 _2315_ (.B1(_0644_),
    .Y(_0217_),
    .A1(_0642_),
    .A2(_0643_));
 sg13g2_a221oi_1 _2316_ (.B2(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[23] ),
    .C1(net58),
    .B1(net66),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[23] ),
    .Y(_0645_),
    .A2(net75));
 sg13g2_o21ai_1 _2317_ (.B1(net35),
    .Y(_0646_),
    .A1(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[23] ),
    .A2(net61));
 sg13g2_nand2_1 _2318_ (.Y(_0647_),
    .A(\u_top_module.u_cic.u_differentiator.temp[23] ),
    .B(net32));
 sg13g2_o21ai_1 _2319_ (.B1(_0647_),
    .Y(_0218_),
    .A1(_0645_),
    .A2(_0646_));
 sg13g2_nor2_1 _2320_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[0] ),
    .B(net48),
    .Y(_0648_));
 sg13g2_a21oi_1 _2321_ (.A1(net48),
    .A2(_0364_),
    .Y(_0219_),
    .B1(_0648_));
 sg13g2_nor2_1 _2322_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[1] ),
    .B(net47),
    .Y(_0649_));
 sg13g2_a21oi_1 _2323_ (.A1(net47),
    .A2(_0371_),
    .Y(_0220_),
    .B1(_0649_));
 sg13g2_nor2_1 _2324_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[2] ),
    .B(net46),
    .Y(_0650_));
 sg13g2_a21oi_1 _2325_ (.A1(net46),
    .A2(_0379_),
    .Y(_0221_),
    .B1(_0650_));
 sg13g2_nor2_1 _2326_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[3] ),
    .B(net47),
    .Y(_0651_));
 sg13g2_a21oi_1 _2327_ (.A1(net47),
    .A2(_0387_),
    .Y(_0222_),
    .B1(_0651_));
 sg13g2_nor2_1 _2328_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[4] ),
    .B(net46),
    .Y(_0652_));
 sg13g2_a21oi_1 _2329_ (.A1(net46),
    .A2(_0395_),
    .Y(_0223_),
    .B1(_0652_));
 sg13g2_nor2_1 _2330_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[5] ),
    .B(net46),
    .Y(_0653_));
 sg13g2_a21oi_1 _2331_ (.A1(net46),
    .A2(_0403_),
    .Y(_0224_),
    .B1(_0653_));
 sg13g2_nor2_1 _2332_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[6] ),
    .B(net46),
    .Y(_0654_));
 sg13g2_a21oi_1 _2333_ (.A1(net46),
    .A2(_0411_),
    .Y(_0225_),
    .B1(_0654_));
 sg13g2_nor2_1 _2334_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[7] ),
    .B(net47),
    .Y(_0655_));
 sg13g2_a21oi_1 _2335_ (.A1(net47),
    .A2(_0419_),
    .Y(_0226_),
    .B1(_0655_));
 sg13g2_nor2_1 _2336_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[8] ),
    .B(net45),
    .Y(_0656_));
 sg13g2_a21oi_1 _2337_ (.A1(net45),
    .A2(_0427_),
    .Y(_0227_),
    .B1(_0656_));
 sg13g2_nor2_1 _2338_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[9] ),
    .B(net45),
    .Y(_0657_));
 sg13g2_a21oi_1 _2339_ (.A1(net45),
    .A2(_0435_),
    .Y(_0228_),
    .B1(_0657_));
 sg13g2_nor2_1 _2340_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[10] ),
    .B(net45),
    .Y(_0658_));
 sg13g2_a21oi_1 _2341_ (.A1(net45),
    .A2(_0444_),
    .Y(_0229_),
    .B1(_0658_));
 sg13g2_nor2_1 _2342_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[11] ),
    .B(net45),
    .Y(_0659_));
 sg13g2_a21oi_1 _2343_ (.A1(net45),
    .A2(_0453_),
    .Y(_0230_),
    .B1(_0659_));
 sg13g2_nor2_1 _2344_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[12] ),
    .B(net43),
    .Y(_0660_));
 sg13g2_a21oi_1 _2345_ (.A1(net43),
    .A2(_0464_),
    .Y(_0231_),
    .B1(_0660_));
 sg13g2_nor2_1 _2346_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[13] ),
    .B(net43),
    .Y(_0661_));
 sg13g2_a21oi_1 _2347_ (.A1(net43),
    .A2(_0473_),
    .Y(_0232_),
    .B1(_0661_));
 sg13g2_nor2_1 _2348_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[14] ),
    .B(net42),
    .Y(_0662_));
 sg13g2_a21oi_1 _2349_ (.A1(net42),
    .A2(_0483_),
    .Y(_0233_),
    .B1(_0662_));
 sg13g2_nor2_1 _2350_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[15] ),
    .B(net42),
    .Y(_0663_));
 sg13g2_a21oi_1 _2351_ (.A1(net42),
    .A2(_0492_),
    .Y(_0234_),
    .B1(_0663_));
 sg13g2_nor2_1 _2352_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[16] ),
    .B(net41),
    .Y(_0664_));
 sg13g2_a21oi_1 _2353_ (.A1(net41),
    .A2(_0503_),
    .Y(_0235_),
    .B1(_0664_));
 sg13g2_nor2_1 _2354_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[17] ),
    .B(net42),
    .Y(_0665_));
 sg13g2_a21oi_1 _2355_ (.A1(net42),
    .A2(_0511_),
    .Y(_0236_),
    .B1(_0665_));
 sg13g2_nor2_1 _2356_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[18] ),
    .B(net40),
    .Y(_0666_));
 sg13g2_a21oi_1 _2357_ (.A1(net40),
    .A2(_0520_),
    .Y(_0237_),
    .B1(_0666_));
 sg13g2_nor2_1 _2358_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[19] ),
    .B(net41),
    .Y(_0667_));
 sg13g2_a21oi_1 _2359_ (.A1(net41),
    .A2(_0529_),
    .Y(_0238_),
    .B1(_0667_));
 sg13g2_nor2_1 _2360_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[20] ),
    .B(net40),
    .Y(_0668_));
 sg13g2_a21oi_1 _2361_ (.A1(net40),
    .A2(_0540_),
    .Y(_0239_),
    .B1(_0668_));
 sg13g2_nor2_1 _2362_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[21] ),
    .B(net40),
    .Y(_0669_));
 sg13g2_a21oi_1 _2363_ (.A1(net40),
    .A2(_0549_),
    .Y(_0240_),
    .B1(_0669_));
 sg13g2_nor2_1 _2364_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[22] ),
    .B(net40),
    .Y(_0670_));
 sg13g2_a21oi_1 _2365_ (.A1(net40),
    .A2(_0557_),
    .Y(_0241_),
    .B1(_0670_));
 sg13g2_nor2_1 _2366_ (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[23] ),
    .B(net42),
    .Y(_0671_));
 sg13g2_a21oi_1 _2367_ (.A1(net42),
    .A2(_0564_),
    .Y(_0242_),
    .B1(_0671_));
 sg13g2_nand2_1 _2368_ (.Y(_0672_),
    .A(net166),
    .B(_0359_));
 sg13g2_nor2_1 _2369_ (.A(_0344_),
    .B(_0672_),
    .Y(_0673_));
 sg13g2_nor2_1 _2370_ (.A(\u_top_module.u_i2s_bus.u_mux_shift.sum_res ),
    .B(net26),
    .Y(_0674_));
 sg13g2_a21oi_1 _2371_ (.A1(_0364_),
    .A2(net26),
    .Y(_0243_),
    .B1(_0674_));
 sg13g2_nor2_1 _2372_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ),
    .B(net27),
    .Y(_0675_));
 sg13g2_a21oi_1 _2373_ (.A1(_0371_),
    .A2(net27),
    .Y(_0244_),
    .B1(_0675_));
 sg13g2_nor2_1 _2374_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ),
    .B(net27),
    .Y(_0676_));
 sg13g2_a21oi_1 _2375_ (.A1(_0379_),
    .A2(net27),
    .Y(_0245_),
    .B1(_0676_));
 sg13g2_nor2_1 _2376_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ),
    .B(net28),
    .Y(_0677_));
 sg13g2_a21oi_1 _2377_ (.A1(_0387_),
    .A2(net28),
    .Y(_0246_),
    .B1(_0677_));
 sg13g2_nor2_1 _2378_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ),
    .B(net27),
    .Y(_0678_));
 sg13g2_a21oi_1 _2379_ (.A1(_0395_),
    .A2(net27),
    .Y(_0247_),
    .B1(_0678_));
 sg13g2_nor2_1 _2380_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ),
    .B(net28),
    .Y(_0679_));
 sg13g2_a21oi_1 _2381_ (.A1(_0403_),
    .A2(net28),
    .Y(_0248_),
    .B1(_0679_));
 sg13g2_nor2_1 _2382_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ),
    .B(net27),
    .Y(_0680_));
 sg13g2_a21oi_1 _2383_ (.A1(_0411_),
    .A2(net27),
    .Y(_0249_),
    .B1(_0680_));
 sg13g2_nor2_1 _2384_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ),
    .B(net25),
    .Y(_0681_));
 sg13g2_a21oi_1 _2385_ (.A1(_0419_),
    .A2(net26),
    .Y(_0250_),
    .B1(_0681_));
 sg13g2_nor2_1 _2386_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ),
    .B(net26),
    .Y(_0682_));
 sg13g2_a21oi_1 _2387_ (.A1(_0427_),
    .A2(net25),
    .Y(_0251_),
    .B1(_0682_));
 sg13g2_nor2_1 _2388_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ),
    .B(net25),
    .Y(_0683_));
 sg13g2_a21oi_1 _2389_ (.A1(_0435_),
    .A2(net25),
    .Y(_0252_),
    .B1(_0683_));
 sg13g2_nor2_1 _2390_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ),
    .B(net25),
    .Y(_0684_));
 sg13g2_a21oi_1 _2391_ (.A1(_0444_),
    .A2(net25),
    .Y(_0253_),
    .B1(_0684_));
 sg13g2_nor2_1 _2392_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ),
    .B(net25),
    .Y(_0685_));
 sg13g2_a21oi_1 _2393_ (.A1(_0453_),
    .A2(net25),
    .Y(_0254_),
    .B1(_0685_));
 sg13g2_nor2_1 _2394_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ),
    .B(net24),
    .Y(_0686_));
 sg13g2_a21oi_1 _2395_ (.A1(_0464_),
    .A2(net30),
    .Y(_0255_),
    .B1(_0686_));
 sg13g2_nor2_1 _2396_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ),
    .B(net24),
    .Y(_0687_));
 sg13g2_a21oi_1 _2397_ (.A1(_0473_),
    .A2(net24),
    .Y(_0256_),
    .B1(_0687_));
 sg13g2_nor2_1 _2398_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ),
    .B(net24),
    .Y(_0688_));
 sg13g2_a21oi_1 _2399_ (.A1(_0483_),
    .A2(net24),
    .Y(_0257_),
    .B1(_0688_));
 sg13g2_nor2_1 _2400_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ),
    .B(net24),
    .Y(_0689_));
 sg13g2_a21oi_1 _2401_ (.A1(_0492_),
    .A2(net24),
    .Y(_0258_),
    .B1(_0689_));
 sg13g2_nor2_1 _2402_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ),
    .B(net22),
    .Y(_0690_));
 sg13g2_a21oi_1 _2403_ (.A1(_0503_),
    .A2(net23),
    .Y(_0259_),
    .B1(_0690_));
 sg13g2_nor2_1 _2404_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ),
    .B(net22),
    .Y(_0691_));
 sg13g2_a21oi_1 _2405_ (.A1(_0511_),
    .A2(net24),
    .Y(_0260_),
    .B1(_0691_));
 sg13g2_nor2_1 _2406_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ),
    .B(net22),
    .Y(_0692_));
 sg13g2_a21oi_1 _2407_ (.A1(_0520_),
    .A2(net22),
    .Y(_0261_),
    .B1(_0692_));
 sg13g2_nor2_1 _2408_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.sum_res ),
    .B(net22),
    .Y(_0693_));
 sg13g2_a21oi_1 _2409_ (.A1(_0529_),
    .A2(net22),
    .Y(_0262_),
    .B1(_0693_));
 sg13g2_nor2_1 _2410_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.sum_res ),
    .B(net22),
    .Y(_0694_));
 sg13g2_a21oi_1 _2411_ (.A1(_0540_),
    .A2(net22),
    .Y(_0263_),
    .B1(_0694_));
 sg13g2_nor2_1 _2412_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.sum_res ),
    .B(net23),
    .Y(_0695_));
 sg13g2_a21oi_1 _2413_ (.A1(_0549_),
    .A2(net23),
    .Y(_0264_),
    .B1(_0695_));
 sg13g2_nor2_1 _2414_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.sum_res ),
    .B(net23),
    .Y(_0696_));
 sg13g2_a21oi_1 _2415_ (.A1(_0557_),
    .A2(net23),
    .Y(_0265_),
    .B1(_0696_));
 sg13g2_nor2_1 _2416_ (.A(\u_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.sum_res ),
    .B(net28),
    .Y(_0697_));
 sg13g2_a21oi_1 _2417_ (.A1(_0564_),
    .A2(net29),
    .Y(_0266_),
    .B1(_0697_));
 sg13g2_nor3_1 _2418_ (.A(net91),
    .B(net84),
    .C(_0344_),
    .Y(_0698_));
 sg13g2_mux2_1 _2419_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[1] ),
    .A1(\u_top_module.u_cic.int_2_out[1] ),
    .S(net21),
    .X(_0267_));
 sg13g2_mux2_1 _2420_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[2] ),
    .A1(\u_top_module.u_cic.int_2_out[2] ),
    .S(net21),
    .X(_0268_));
 sg13g2_mux2_1 _2421_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[3] ),
    .A1(\u_top_module.u_cic.int_2_out[3] ),
    .S(net20),
    .X(_0269_));
 sg13g2_mux2_1 _2422_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[4] ),
    .A1(\u_top_module.u_cic.int_2_out[4] ),
    .S(net20),
    .X(_0270_));
 sg13g2_mux2_1 _2423_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[5] ),
    .A1(\u_top_module.u_cic.int_2_out[5] ),
    .S(net20),
    .X(_0271_));
 sg13g2_mux2_1 _2424_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[6] ),
    .A1(\u_top_module.u_cic.int_2_out[6] ),
    .S(net20),
    .X(_0272_));
 sg13g2_mux2_1 _2425_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[7] ),
    .A1(\u_top_module.u_cic.int_2_out[7] ),
    .S(net20),
    .X(_0273_));
 sg13g2_mux2_1 _2426_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[8] ),
    .A1(\u_top_module.u_cic.int_2_out[8] ),
    .S(net20),
    .X(_0274_));
 sg13g2_mux2_1 _2427_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[9] ),
    .A1(\u_top_module.u_cic.int_2_out[9] ),
    .S(net20),
    .X(_0275_));
 sg13g2_mux2_1 _2428_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[10] ),
    .A1(\u_top_module.u_cic.int_2_out[10] ),
    .S(net19),
    .X(_0276_));
 sg13g2_mux2_1 _2429_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[11] ),
    .A1(\u_top_module.u_cic.int_2_out[11] ),
    .S(net20),
    .X(_0277_));
 sg13g2_mux2_1 _2430_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[12] ),
    .A1(\u_top_module.u_cic.int_2_out[12] ),
    .S(net19),
    .X(_0278_));
 sg13g2_mux2_1 _2431_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[13] ),
    .A1(\u_top_module.u_cic.int_2_out[13] ),
    .S(net19),
    .X(_0279_));
 sg13g2_mux2_1 _2432_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[14] ),
    .A1(\u_top_module.u_cic.int_2_out[14] ),
    .S(net19),
    .X(_0280_));
 sg13g2_mux2_1 _2433_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[15] ),
    .A1(\u_top_module.u_cic.int_2_out[15] ),
    .S(net19),
    .X(_0281_));
 sg13g2_mux2_1 _2434_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[16] ),
    .A1(\u_top_module.u_cic.int_2_out[16] ),
    .S(net18),
    .X(_0282_));
 sg13g2_mux2_1 _2435_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[17] ),
    .A1(\u_top_module.u_cic.int_2_out[17] ),
    .S(net18),
    .X(_0283_));
 sg13g2_mux2_1 _2436_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[18] ),
    .A1(\u_top_module.u_cic.int_2_out[18] ),
    .S(net18),
    .X(_0284_));
 sg13g2_mux2_1 _2437_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[19] ),
    .A1(\u_top_module.u_cic.int_2_out[19] ),
    .S(net18),
    .X(_0285_));
 sg13g2_mux2_1 _2438_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[20] ),
    .A1(\u_top_module.u_cic.int_2_out[20] ),
    .S(net18),
    .X(_0286_));
 sg13g2_mux2_1 _2439_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[21] ),
    .A1(\u_top_module.u_cic.int_2_out[21] ),
    .S(net18),
    .X(_0287_));
 sg13g2_mux2_1 _2440_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[22] ),
    .A1(\u_top_module.u_cic.int_2_out[22] ),
    .S(net18),
    .X(_0288_));
 sg13g2_mux2_1 _2441_ (.A0(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[23] ),
    .A1(\u_top_module.u_cic.int_2_out[23] ),
    .S(net18),
    .X(_0289_));
 sg13g2_inv_1 _2442_ (.Y(_0126_),
    .A(net126));
 sg13g2_inv_1 _2443_ (.Y(_0127_),
    .A(net128));
 sg13g2_inv_1 _2444_ (.Y(_0128_),
    .A(net128));
 sg13g2_inv_1 _2445_ (.Y(_0129_),
    .A(net128));
 sg13g2_inv_1 _2446_ (.Y(_0130_),
    .A(net129));
 sg13g2_inv_1 _2447_ (.Y(_0131_),
    .A(net137));
 sg13g2_inv_1 _2448_ (.Y(_0132_),
    .A(net131));
 sg13g2_inv_1 _2449_ (.Y(_0133_),
    .A(net126));
 sg13g2_inv_1 _2450_ (.Y(_0134_),
    .A(net116));
 sg13g2_inv_1 _2451_ (.Y(_0135_),
    .A(net116));
 sg13g2_inv_1 _2452_ (.Y(_0136_),
    .A(net116));
 sg13g2_inv_1 _2453_ (.Y(_0137_),
    .A(net116));
 sg13g2_inv_1 _2454_ (.Y(_0138_),
    .A(net113));
 sg13g2_inv_1 _2455_ (.Y(_0139_),
    .A(net113));
 sg13g2_inv_1 _2456_ (.Y(_0140_),
    .A(net104));
 sg13g2_inv_1 _2457_ (.Y(_0141_),
    .A(net104));
 sg13g2_inv_1 _2458_ (.Y(_0142_),
    .A(net104));
 sg13g2_inv_1 _2459_ (.Y(_0143_),
    .A(net103));
 sg13g2_inv_1 _2460_ (.Y(_0144_),
    .A(net103));
 sg13g2_inv_1 _2461_ (.Y(_0145_),
    .A(net103));
 sg13g2_inv_1 _2462_ (.Y(_0146_),
    .A(net103));
 sg13g2_inv_1 _2463_ (.Y(_0147_),
    .A(net97));
 sg13g2_inv_1 _2464_ (.Y(_0148_),
    .A(net121));
 sg13g2_inv_1 _2465_ (.Y(_0149_),
    .A(net124));
 sg13g2_inv_1 _2466_ (.Y(_0150_),
    .A(net124));
 sg13g2_inv_1 _2467_ (.Y(_0151_),
    .A(net132));
 sg13g2_inv_1 _2468_ (.Y(_0152_),
    .A(net132));
 sg13g2_inv_1 _2469_ (.Y(_0153_),
    .A(net134));
 sg13g2_inv_1 _2470_ (.Y(_0154_),
    .A(net134));
 sg13g2_inv_1 _2471_ (.Y(_0155_),
    .A(net134));
 sg13g2_inv_1 _2472_ (.Y(_0156_),
    .A(net134));
 sg13g2_inv_1 _2473_ (.Y(_0157_),
    .A(net135));
 sg13g2_inv_1 _2474_ (.Y(_0158_),
    .A(net141));
 sg13g2_inv_1 _2475_ (.Y(_0159_),
    .A(net137));
 sg13g2_inv_1 _2476_ (.Y(_0160_),
    .A(net137));
 sg13g2_inv_1 _2477_ (.Y(_0161_),
    .A(net139));
 sg13g2_inv_1 _2478_ (.Y(_0162_),
    .A(net139));
 sg13g2_inv_1 _2479_ (.Y(_0163_),
    .A(net140));
 sg13g2_inv_1 _2480_ (.Y(_0164_),
    .A(net139));
 sg13g2_inv_1 _2481_ (.Y(_0165_),
    .A(net141));
 sg13g2_dfrbp_1 _2482_ (.CLK(net126),
    .RESET_B(net204),
    .D(_0166_),
    .Q_N(_1218_),
    .Q(\u_top_module.u_i2s_bus.u_mux_shift.data ));
 sg13g2_dfrbp_1 _2483_ (.CLK(net118),
    .RESET_B(net160),
    .D(_0167_),
    .Q_N(_1217_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.sel[0] ));
 sg13g2_dfrbp_1 _2484_ (.CLK(net127),
    .RESET_B(net166),
    .D(_0168_),
    .Q_N(_1216_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.sel[1] ));
 sg13g2_dfrbp_1 _2485_ (.CLK(net127),
    .RESET_B(net166),
    .D(_0169_),
    .Q_N(_1215_),
    .Q(\u_top_module.u_cic.u_differentiator.count[2] ));
 sg13g2_dfrbp_1 _2486_ (.CLK(_0125_),
    .RESET_B(net291),
    .D(_0170_),
    .Q_N(_1214_),
    .Q(out));
 sg13g2_dfrbp_1 _2487_ (.CLK(_0126_),
    .RESET_B(net206),
    .D(\u_top_module.u_i2s_bus.u_mux_shift.data ),
    .Q_N(_1219_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _2488_ (.CLK(net128),
    .RESET_B(net290),
    .D(_0010_),
    .Q_N(_1213_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2489_ (.CLK(_0127_),
    .RESET_B(net208),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.data ),
    .Q_N(_1220_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2490_ (.CLK(net128),
    .RESET_B(net289),
    .D(_0021_),
    .Q_N(_1212_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2491_ (.CLK(_0128_),
    .RESET_B(net210),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.data ),
    .Q_N(_1221_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2492_ (.CLK(net129),
    .RESET_B(net288),
    .D(_0024_),
    .Q_N(_1211_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2493_ (.CLK(_0129_),
    .RESET_B(net212),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.data ),
    .Q_N(_1222_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2494_ (.CLK(net129),
    .RESET_B(net287),
    .D(_0025_),
    .Q_N(_1210_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2495_ (.CLK(_0130_),
    .RESET_B(net214),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.data ),
    .Q_N(_1223_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2496_ (.CLK(net138),
    .RESET_B(net286),
    .D(_0026_),
    .Q_N(_1209_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2497_ (.CLK(_0131_),
    .RESET_B(net216),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.data ),
    .Q_N(_1224_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2498_ (.CLK(net131),
    .RESET_B(net285),
    .D(_0027_),
    .Q_N(_1208_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2499_ (.CLK(_0132_),
    .RESET_B(net218),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.data ),
    .Q_N(_1225_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2500_ (.CLK(net126),
    .RESET_B(net284),
    .D(_0028_),
    .Q_N(_1207_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2501_ (.CLK(_0133_),
    .RESET_B(net220),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.data ),
    .Q_N(_1226_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2502_ (.CLK(net117),
    .RESET_B(net283),
    .D(_0029_),
    .Q_N(_1206_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2503_ (.CLK(_0134_),
    .RESET_B(net222),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.data ),
    .Q_N(_1227_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2504_ (.CLK(net117),
    .RESET_B(net282),
    .D(_0030_),
    .Q_N(_1205_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[9].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2505_ (.CLK(_0135_),
    .RESET_B(net223),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[9].u_mux_shift.data ),
    .Q_N(_1228_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.last_shift ));
 sg13g2_dfrbp_1 _2506_ (.CLK(net116),
    .RESET_B(net225),
    .D(_0000_),
    .Q_N(_1229_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2507_ (.CLK(net133),
    .RESET_B(net281),
    .D(net11),
    .Q_N(_1204_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.prev_lr_clk ));
 sg13g2_dfrbp_1 _2508_ (.CLK(_0136_),
    .RESET_B(net227),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.data ),
    .Q_N(_1230_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2509_ (.CLK(net116),
    .RESET_B(net280),
    .D(_0001_),
    .Q_N(_1203_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2510_ (.CLK(_0137_),
    .RESET_B(net229),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.data ),
    .Q_N(_1231_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2511_ (.CLK(net113),
    .RESET_B(net279),
    .D(_0002_),
    .Q_N(_1202_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2512_ (.CLK(_0138_),
    .RESET_B(net231),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.data ),
    .Q_N(_1232_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2513_ (.CLK(net113),
    .RESET_B(net278),
    .D(_0003_),
    .Q_N(_1201_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2514_ (.CLK(_0139_),
    .RESET_B(net233),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.data ),
    .Q_N(_1233_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2515_ (.CLK(net113),
    .RESET_B(net277),
    .D(_0004_),
    .Q_N(_1200_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2516_ (.CLK(_0140_),
    .RESET_B(net235),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.data ),
    .Q_N(_1234_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2517_ (.CLK(net106),
    .RESET_B(net276),
    .D(_0005_),
    .Q_N(_1199_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2518_ (.CLK(_0141_),
    .RESET_B(net237),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.data ),
    .Q_N(_1235_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2519_ (.CLK(net104),
    .RESET_B(net275),
    .D(_0006_),
    .Q_N(_1198_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2520_ (.CLK(_0142_),
    .RESET_B(net239),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.data ),
    .Q_N(_1236_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2521_ (.CLK(net104),
    .RESET_B(net274),
    .D(_0007_),
    .Q_N(_1197_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2522_ (.CLK(_0143_),
    .RESET_B(net241),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.data ),
    .Q_N(_1237_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2523_ (.CLK(net103),
    .RESET_B(net273),
    .D(_0008_),
    .Q_N(_1196_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2524_ (.CLK(_0144_),
    .RESET_B(net243),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.data ),
    .Q_N(_1238_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2525_ (.CLK(net103),
    .RESET_B(net272),
    .D(_0009_),
    .Q_N(_1195_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2526_ (.CLK(_0145_),
    .RESET_B(net245),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.data ),
    .Q_N(_1239_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2527_ (.CLK(net102),
    .RESET_B(net271),
    .D(_0011_),
    .Q_N(_1194_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2528_ (.CLK(_0146_),
    .RESET_B(net247),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.data ),
    .Q_N(_1240_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2529_ (.CLK(net97),
    .RESET_B(net270),
    .D(_0012_),
    .Q_N(_1193_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2530_ (.CLK(_0147_),
    .RESET_B(net249),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.data ),
    .Q_N(_1241_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2531_ (.CLK(net121),
    .RESET_B(net269),
    .D(_0013_),
    .Q_N(_1192_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2532_ (.CLK(_0148_),
    .RESET_B(net250),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.data ),
    .Q_N(_1242_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2533_ (.CLK(net124),
    .RESET_B(net268),
    .D(_0014_),
    .Q_N(_1191_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2534_ (.CLK(_0149_),
    .RESET_B(net251),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.data ),
    .Q_N(_1243_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2535_ (.CLK(net124),
    .RESET_B(net267),
    .D(_0015_),
    .Q_N(_1190_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2536_ (.CLK(_0150_),
    .RESET_B(net252),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.data ),
    .Q_N(_1244_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[24].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2537_ (.CLK(net132),
    .RESET_B(net266),
    .D(_0016_),
    .Q_N(_1189_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2538_ (.CLK(_0151_),
    .RESET_B(net253),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.data ),
    .Q_N(_1245_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[25].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2539_ (.CLK(net132),
    .RESET_B(net265),
    .D(_0017_),
    .Q_N(_1188_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2540_ (.CLK(_0152_),
    .RESET_B(net254),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.data ),
    .Q_N(_1246_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[26].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2541_ (.CLK(net134),
    .RESET_B(net264),
    .D(_0018_),
    .Q_N(_1187_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2542_ (.CLK(_0153_),
    .RESET_B(net255),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.data ),
    .Q_N(_1247_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[27].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2543_ (.CLK(net134),
    .RESET_B(net263),
    .D(_0019_),
    .Q_N(_1186_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2544_ (.CLK(_0154_),
    .RESET_B(net256),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.data ),
    .Q_N(_1248_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[28].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2545_ (.CLK(net134),
    .RESET_B(net262),
    .D(_0020_),
    .Q_N(_1185_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2546_ (.CLK(_0155_),
    .RESET_B(net257),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.data ),
    .Q_N(_1249_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[29].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2547_ (.CLK(net135),
    .RESET_B(net261),
    .D(_0022_),
    .Q_N(_1184_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2548_ (.CLK(_0156_),
    .RESET_B(net258),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.data ),
    .Q_N(_1250_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[30].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2549_ (.CLK(net135),
    .RESET_B(net260),
    .D(_0023_),
    .Q_N(_1183_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.data ));
 sg13g2_dfrbp_1 _2550_ (.CLK(_0157_),
    .RESET_B(net259),
    .D(\u_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.data ),
    .Q_N(_1251_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[31].u_mux_shift.out ));
 sg13g2_dfrbp_1 _2551_ (.CLK(net135),
    .RESET_B(net171),
    .D(_0079_),
    .Q_N(_1252_),
    .Q(\u_top_module.u_cic.inc_out[1] ));
 sg13g2_dfrbp_1 _2552_ (.CLK(net133),
    .RESET_B(net170),
    .D(_0094_),
    .Q_N(_1253_),
    .Q(\u_top_module.u_cic.inc_out[2] ));
 sg13g2_dfrbp_1 _2553_ (.CLK(net133),
    .RESET_B(net170),
    .D(_0095_),
    .Q_N(_1254_),
    .Q(\u_top_module.u_cic.inc_out[3] ));
 sg13g2_dfrbp_1 _2554_ (.CLK(net132),
    .RESET_B(net170),
    .D(_0096_),
    .Q_N(_1255_),
    .Q(\u_top_module.u_cic.inc_out[4] ));
 sg13g2_dfrbp_1 _2555_ (.CLK(net132),
    .RESET_B(net170),
    .D(_0097_),
    .Q_N(_1256_),
    .Q(\u_top_module.u_cic.inc_out[5] ));
 sg13g2_dfrbp_1 _2556_ (.CLK(net132),
    .RESET_B(net170),
    .D(_0098_),
    .Q_N(_1257_),
    .Q(\u_top_module.u_cic.inc_out[6] ));
 sg13g2_dfrbp_1 _2557_ (.CLK(net132),
    .RESET_B(net170),
    .D(_0099_),
    .Q_N(_1258_),
    .Q(\u_top_module.u_cic.inc_out[7] ));
 sg13g2_dfrbp_1 _2558_ (.CLK(net121),
    .RESET_B(net162),
    .D(_0100_),
    .Q_N(_1259_),
    .Q(\u_top_module.u_cic.inc_out[8] ));
 sg13g2_dfrbp_1 _2559_ (.CLK(net121),
    .RESET_B(net162),
    .D(_0101_),
    .Q_N(_1260_),
    .Q(\u_top_module.u_cic.inc_out[9] ));
 sg13g2_dfrbp_1 _2560_ (.CLK(net111),
    .RESET_B(net156),
    .D(_0080_),
    .Q_N(_1261_),
    .Q(\u_top_module.u_cic.inc_out[10] ));
 sg13g2_dfrbp_1 _2561_ (.CLK(net111),
    .RESET_B(net156),
    .D(_0081_),
    .Q_N(_1262_),
    .Q(\u_top_module.u_cic.inc_out[11] ));
 sg13g2_dfrbp_1 _2562_ (.CLK(net111),
    .RESET_B(net156),
    .D(_0082_),
    .Q_N(_1263_),
    .Q(\u_top_module.u_cic.inc_out[12] ));
 sg13g2_dfrbp_1 _2563_ (.CLK(net111),
    .RESET_B(net156),
    .D(_0083_),
    .Q_N(_1264_),
    .Q(\u_top_module.u_cic.inc_out[13] ));
 sg13g2_dfrbp_1 _2564_ (.CLK(net108),
    .RESET_B(net153),
    .D(_0084_),
    .Q_N(_1265_),
    .Q(\u_top_module.u_cic.inc_out[14] ));
 sg13g2_dfrbp_1 _2565_ (.CLK(net108),
    .RESET_B(net153),
    .D(_0085_),
    .Q_N(_1266_),
    .Q(\u_top_module.u_cic.inc_out[15] ));
 sg13g2_dfrbp_1 _2566_ (.CLK(net108),
    .RESET_B(net153),
    .D(_0086_),
    .Q_N(_1267_),
    .Q(\u_top_module.u_cic.inc_out[16] ));
 sg13g2_dfrbp_1 _2567_ (.CLK(net100),
    .RESET_B(net148),
    .D(_0087_),
    .Q_N(_0035_),
    .Q(\u_top_module.u_cic.inc_out[17] ));
 sg13g2_dfrbp_1 _2568_ (.CLK(net100),
    .RESET_B(net148),
    .D(_0088_),
    .Q_N(_1268_),
    .Q(\u_top_module.u_cic.inc_out[18] ));
 sg13g2_dfrbp_1 _2569_ (.CLK(net100),
    .RESET_B(net148),
    .D(_0089_),
    .Q_N(_1269_),
    .Q(\u_top_module.u_cic.inc_out[19] ));
 sg13g2_dfrbp_1 _2570_ (.CLK(net96),
    .RESET_B(net145),
    .D(_0090_),
    .Q_N(_1270_),
    .Q(\u_top_module.u_cic.inc_out[20] ));
 sg13g2_dfrbp_1 _2571_ (.CLK(net96),
    .RESET_B(net145),
    .D(_0091_),
    .Q_N(_1271_),
    .Q(\u_top_module.u_cic.inc_out[21] ));
 sg13g2_dfrbp_1 _2572_ (.CLK(net96),
    .RESET_B(net144),
    .D(_0092_),
    .Q_N(_1272_),
    .Q(\u_top_module.u_cic.inc_out[22] ));
 sg13g2_dfrbp_1 _2573_ (.CLK(net96),
    .RESET_B(net144),
    .D(_0093_),
    .Q_N(_1273_),
    .Q(\u_top_module.u_cic.inc_out[23] ));
 sg13g2_dfrbp_1 _2574_ (.CLK(net135),
    .RESET_B(net171),
    .D(_0056_),
    .Q_N(_1274_),
    .Q(\u_top_module.u_cic.int_1_out[1] ));
 sg13g2_dfrbp_1 _2575_ (.CLK(net133),
    .RESET_B(net170),
    .D(_0071_),
    .Q_N(_1275_),
    .Q(\u_top_module.u_cic.int_1_out[2] ));
 sg13g2_dfrbp_1 _2576_ (.CLK(net133),
    .RESET_B(net170),
    .D(_0072_),
    .Q_N(_1276_),
    .Q(\u_top_module.u_cic.int_1_out[3] ));
 sg13g2_dfrbp_1 _2577_ (.CLK(net124),
    .RESET_B(net165),
    .D(_0073_),
    .Q_N(_1277_),
    .Q(\u_top_module.u_cic.int_1_out[4] ));
 sg13g2_dfrbp_1 _2578_ (.CLK(net124),
    .RESET_B(net165),
    .D(_0074_),
    .Q_N(_1278_),
    .Q(\u_top_module.u_cic.int_1_out[5] ));
 sg13g2_dfrbp_1 _2579_ (.CLK(net124),
    .RESET_B(net165),
    .D(_0075_),
    .Q_N(_1279_),
    .Q(\u_top_module.u_cic.int_1_out[6] ));
 sg13g2_dfrbp_1 _2580_ (.CLK(net122),
    .RESET_B(net162),
    .D(_0076_),
    .Q_N(_1280_),
    .Q(\u_top_module.u_cic.int_1_out[7] ));
 sg13g2_dfrbp_1 _2581_ (.CLK(net121),
    .RESET_B(net162),
    .D(_0077_),
    .Q_N(_1281_),
    .Q(\u_top_module.u_cic.int_1_out[8] ));
 sg13g2_dfrbp_1 _2582_ (.CLK(net121),
    .RESET_B(net162),
    .D(_0078_),
    .Q_N(_1282_),
    .Q(\u_top_module.u_cic.int_1_out[9] ));
 sg13g2_dfrbp_1 _2583_ (.CLK(net111),
    .RESET_B(net156),
    .D(_0057_),
    .Q_N(_1283_),
    .Q(\u_top_module.u_cic.int_1_out[10] ));
 sg13g2_dfrbp_1 _2584_ (.CLK(net111),
    .RESET_B(net156),
    .D(_0058_),
    .Q_N(_1284_),
    .Q(\u_top_module.u_cic.int_1_out[11] ));
 sg13g2_dfrbp_1 _2585_ (.CLK(net111),
    .RESET_B(net156),
    .D(_0059_),
    .Q_N(_1285_),
    .Q(\u_top_module.u_cic.int_1_out[12] ));
 sg13g2_dfrbp_1 _2586_ (.CLK(net108),
    .RESET_B(net153),
    .D(_0060_),
    .Q_N(_1286_),
    .Q(\u_top_module.u_cic.int_1_out[13] ));
 sg13g2_dfrbp_1 _2587_ (.CLK(net108),
    .RESET_B(net153),
    .D(_0061_),
    .Q_N(_1287_),
    .Q(\u_top_module.u_cic.int_1_out[14] ));
 sg13g2_dfrbp_1 _2588_ (.CLK(net108),
    .RESET_B(net153),
    .D(_0062_),
    .Q_N(_1288_),
    .Q(\u_top_module.u_cic.int_1_out[15] ));
 sg13g2_dfrbp_1 _2589_ (.CLK(net108),
    .RESET_B(net153),
    .D(_0063_),
    .Q_N(_1289_),
    .Q(\u_top_module.u_cic.int_1_out[16] ));
 sg13g2_dfrbp_1 _2590_ (.CLK(net100),
    .RESET_B(net148),
    .D(_0064_),
    .Q_N(_1290_),
    .Q(\u_top_module.u_cic.int_1_out[17] ));
 sg13g2_dfrbp_1 _2591_ (.CLK(net100),
    .RESET_B(net148),
    .D(_0065_),
    .Q_N(_1291_),
    .Q(\u_top_module.u_cic.int_1_out[18] ));
 sg13g2_dfrbp_1 _2592_ (.CLK(net100),
    .RESET_B(net148),
    .D(_0066_),
    .Q_N(_1292_),
    .Q(\u_top_module.u_cic.int_1_out[19] ));
 sg13g2_dfrbp_1 _2593_ (.CLK(net96),
    .RESET_B(net145),
    .D(_0067_),
    .Q_N(_1293_),
    .Q(\u_top_module.u_cic.int_1_out[20] ));
 sg13g2_dfrbp_1 _2594_ (.CLK(net98),
    .RESET_B(net144),
    .D(_0068_),
    .Q_N(_1294_),
    .Q(\u_top_module.u_cic.int_1_out[21] ));
 sg13g2_dfrbp_1 _2595_ (.CLK(net96),
    .RESET_B(net144),
    .D(_0069_),
    .Q_N(_1295_),
    .Q(\u_top_module.u_cic.int_1_out[22] ));
 sg13g2_dfrbp_1 _2596_ (.CLK(net96),
    .RESET_B(net144),
    .D(_0070_),
    .Q_N(_1296_),
    .Q(\u_top_module.u_cic.int_1_out[23] ));
 sg13g2_dfrbp_1 _2597_ (.CLK(net140),
    .RESET_B(net175),
    .D(_0112_),
    .Q_N(_1297_),
    .Q(\u_top_module.u_cic.int_2_out[1] ));
 sg13g2_dfrbp_1 _2598_ (.CLK(net138),
    .RESET_B(net172),
    .D(_0117_),
    .Q_N(_1298_),
    .Q(\u_top_module.u_cic.int_2_out[2] ));
 sg13g2_dfrbp_1 _2599_ (.CLK(net133),
    .RESET_B(net171),
    .D(_0118_),
    .Q_N(_1299_),
    .Q(\u_top_module.u_cic.int_2_out[3] ));
 sg13g2_dfrbp_1 _2600_ (.CLK(net123),
    .RESET_B(net164),
    .D(_0119_),
    .Q_N(_1300_),
    .Q(\u_top_module.u_cic.int_2_out[4] ));
 sg13g2_dfrbp_1 _2601_ (.CLK(net123),
    .RESET_B(net164),
    .D(_0120_),
    .Q_N(_1301_),
    .Q(\u_top_module.u_cic.int_2_out[5] ));
 sg13g2_dfrbp_1 _2602_ (.CLK(net123),
    .RESET_B(net164),
    .D(_0121_),
    .Q_N(_1302_),
    .Q(\u_top_module.u_cic.int_2_out[6] ));
 sg13g2_dfrbp_1 _2603_ (.CLK(net122),
    .RESET_B(net162),
    .D(_0122_),
    .Q_N(_1303_),
    .Q(\u_top_module.u_cic.int_2_out[7] ));
 sg13g2_dfrbp_1 _2604_ (.CLK(net121),
    .RESET_B(net162),
    .D(_0123_),
    .Q_N(_1304_),
    .Q(\u_top_module.u_cic.int_2_out[8] ));
 sg13g2_dfrbp_1 _2605_ (.CLK(net121),
    .RESET_B(net162),
    .D(_0124_),
    .Q_N(_1305_),
    .Q(\u_top_module.u_cic.int_2_out[9] ));
 sg13g2_dfrbp_1 _2606_ (.CLK(net109),
    .RESET_B(net155),
    .D(_0102_),
    .Q_N(_1306_),
    .Q(\u_top_module.u_cic.int_2_out[10] ));
 sg13g2_dfrbp_1 _2607_ (.CLK(net109),
    .RESET_B(net156),
    .D(_0103_),
    .Q_N(_1307_),
    .Q(\u_top_module.u_cic.int_2_out[11] ));
 sg13g2_dfrbp_1 _2608_ (.CLK(net109),
    .RESET_B(net155),
    .D(_0104_),
    .Q_N(_1308_),
    .Q(\u_top_module.u_cic.int_2_out[12] ));
 sg13g2_dfrbp_1 _2609_ (.CLK(net107),
    .RESET_B(net152),
    .D(_0105_),
    .Q_N(_1309_),
    .Q(\u_top_module.u_cic.int_2_out[13] ));
 sg13g2_dfrbp_1 _2610_ (.CLK(net107),
    .RESET_B(net152),
    .D(_0106_),
    .Q_N(_1310_),
    .Q(\u_top_module.u_cic.int_2_out[14] ));
 sg13g2_dfrbp_1 _2611_ (.CLK(net108),
    .RESET_B(net153),
    .D(_0107_),
    .Q_N(_1311_),
    .Q(\u_top_module.u_cic.int_2_out[15] ));
 sg13g2_dfrbp_1 _2612_ (.CLK(net107),
    .RESET_B(net147),
    .D(_0108_),
    .Q_N(_1312_),
    .Q(\u_top_module.u_cic.int_2_out[16] ));
 sg13g2_dfrbp_1 _2613_ (.CLK(net99),
    .RESET_B(net147),
    .D(_0109_),
    .Q_N(_1313_),
    .Q(\u_top_module.u_cic.int_2_out[17] ));
 sg13g2_dfrbp_1 _2614_ (.CLK(net100),
    .RESET_B(net148),
    .D(_0110_),
    .Q_N(_1314_),
    .Q(\u_top_module.u_cic.int_2_out[18] ));
 sg13g2_dfrbp_1 _2615_ (.CLK(net100),
    .RESET_B(net148),
    .D(_0111_),
    .Q_N(_1315_),
    .Q(\u_top_module.u_cic.int_2_out[19] ));
 sg13g2_dfrbp_1 _2616_ (.CLK(net98),
    .RESET_B(net145),
    .D(_0113_),
    .Q_N(_1316_),
    .Q(\u_top_module.u_cic.int_2_out[20] ));
 sg13g2_dfrbp_1 _2617_ (.CLK(net98),
    .RESET_B(net144),
    .D(_0114_),
    .Q_N(_1317_),
    .Q(\u_top_module.u_cic.int_2_out[21] ));
 sg13g2_dfrbp_1 _2618_ (.CLK(net97),
    .RESET_B(net144),
    .D(_0115_),
    .Q_N(_1318_),
    .Q(\u_top_module.u_cic.int_2_out[22] ));
 sg13g2_dfrbp_1 _2619_ (.CLK(net96),
    .RESET_B(net144),
    .D(_0116_),
    .Q_N(_1182_),
    .Q(\u_top_module.u_cic.int_2_out[23] ));
 sg13g2_dfrbp_1 _2620_ (.CLK(net126),
    .RESET_B(net166),
    .D(_0171_),
    .Q_N(_1181_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[0] ));
 sg13g2_dfrbp_1 _2621_ (.CLK(net127),
    .RESET_B(net166),
    .D(_0172_),
    .Q_N(_0037_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[1] ));
 sg13g2_dfrbp_1 _2622_ (.CLK(net128),
    .RESET_B(net167),
    .D(_0173_),
    .Q_N(_1180_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[2] ));
 sg13g2_dfrbp_1 _2623_ (.CLK(net130),
    .RESET_B(net167),
    .D(_0174_),
    .Q_N(_0039_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[3] ));
 sg13g2_dfrbp_1 _2624_ (.CLK(net130),
    .RESET_B(net167),
    .D(_0175_),
    .Q_N(_1179_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[4] ));
 sg13g2_dfrbp_1 _2625_ (.CLK(net123),
    .RESET_B(net164),
    .D(_0176_),
    .Q_N(_0041_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[5] ));
 sg13g2_dfrbp_1 _2626_ (.CLK(net123),
    .RESET_B(net164),
    .D(_0177_),
    .Q_N(_1178_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[6] ));
 sg13g2_dfrbp_1 _2627_ (.CLK(net122),
    .RESET_B(net163),
    .D(_0178_),
    .Q_N(_0043_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[7] ));
 sg13g2_dfrbp_1 _2628_ (.CLK(net109),
    .RESET_B(net155),
    .D(_0179_),
    .Q_N(_1177_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[8] ));
 sg13g2_dfrbp_1 _2629_ (.CLK(net110),
    .RESET_B(net155),
    .D(_0180_),
    .Q_N(_0045_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[9] ));
 sg13g2_dfrbp_1 _2630_ (.CLK(net109),
    .RESET_B(net152),
    .D(_0181_),
    .Q_N(_1176_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[10] ));
 sg13g2_dfrbp_1 _2631_ (.CLK(net118),
    .RESET_B(net160),
    .D(_0182_),
    .Q_N(_0047_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[11] ));
 sg13g2_dfrbp_1 _2632_ (.CLK(net114),
    .RESET_B(net158),
    .D(_0183_),
    .Q_N(_1175_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[12] ));
 sg13g2_dfrbp_1 _2633_ (.CLK(net115),
    .RESET_B(net158),
    .D(_0184_),
    .Q_N(_0049_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[13] ));
 sg13g2_dfrbp_1 _2634_ (.CLK(net113),
    .RESET_B(net159),
    .D(_0185_),
    .Q_N(_1174_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[14] ));
 sg13g2_dfrbp_1 _2635_ (.CLK(net115),
    .RESET_B(net158),
    .D(_0186_),
    .Q_N(_0051_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[15] ));
 sg13g2_dfrbp_1 _2636_ (.CLK(net104),
    .RESET_B(net150),
    .D(_0187_),
    .Q_N(_1173_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[16] ));
 sg13g2_dfrbp_1 _2637_ (.CLK(net105),
    .RESET_B(net150),
    .D(_0188_),
    .Q_N(_0053_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[17] ));
 sg13g2_dfrbp_1 _2638_ (.CLK(net102),
    .RESET_B(net151),
    .D(_0189_),
    .Q_N(_1172_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[18] ));
 sg13g2_dfrbp_1 _2639_ (.CLK(net105),
    .RESET_B(net150),
    .D(_0190_),
    .Q_N(_0055_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[19] ));
 sg13g2_dfrbp_1 _2640_ (.CLK(net102),
    .RESET_B(net151),
    .D(_0191_),
    .Q_N(_1171_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[20] ));
 sg13g2_dfrbp_1 _2641_ (.CLK(net97),
    .RESET_B(net146),
    .D(_0192_),
    .Q_N(_1170_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[21] ));
 sg13g2_dfrbp_1 _2642_ (.CLK(net99),
    .RESET_B(net147),
    .D(_0193_),
    .Q_N(_1169_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[22] ));
 sg13g2_dfrbp_1 _2643_ (.CLK(net107),
    .RESET_B(net152),
    .D(_0194_),
    .Q_N(_1168_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d2[23] ));
 sg13g2_dfrbp_1 _2644_ (.CLK(net127),
    .RESET_B(net166),
    .D(_0195_),
    .Q_N(_1167_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[0] ));
 sg13g2_dfrbp_1 _2645_ (.CLK(net127),
    .RESET_B(net166),
    .D(_0196_),
    .Q_N(_1166_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[1] ));
 sg13g2_dfrbp_1 _2646_ (.CLK(net130),
    .RESET_B(net167),
    .D(_0197_),
    .Q_N(_1165_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[2] ));
 sg13g2_dfrbp_1 _2647_ (.CLK(net130),
    .RESET_B(net167),
    .D(_0198_),
    .Q_N(_1164_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[3] ));
 sg13g2_dfrbp_1 _2648_ (.CLK(net130),
    .RESET_B(net167),
    .D(_0199_),
    .Q_N(_1163_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[4] ));
 sg13g2_dfrbp_1 _2649_ (.CLK(net125),
    .RESET_B(net165),
    .D(_0200_),
    .Q_N(_1162_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[5] ));
 sg13g2_dfrbp_1 _2650_ (.CLK(net123),
    .RESET_B(net164),
    .D(_0201_),
    .Q_N(_1161_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[6] ));
 sg13g2_dfrbp_1 _2651_ (.CLK(net122),
    .RESET_B(net163),
    .D(_0202_),
    .Q_N(_1160_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[7] ));
 sg13g2_dfrbp_1 _2652_ (.CLK(net122),
    .RESET_B(net163),
    .D(_0203_),
    .Q_N(_1159_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[8] ));
 sg13g2_dfrbp_1 _2653_ (.CLK(net118),
    .RESET_B(net160),
    .D(_0204_),
    .Q_N(_1158_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[9] ));
 sg13g2_dfrbp_1 _2654_ (.CLK(net118),
    .RESET_B(net160),
    .D(_0205_),
    .Q_N(_1157_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[10] ));
 sg13g2_dfrbp_1 _2655_ (.CLK(net118),
    .RESET_B(net160),
    .D(_0206_),
    .Q_N(_1156_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[11] ));
 sg13g2_dfrbp_1 _2656_ (.CLK(net115),
    .RESET_B(net159),
    .D(_0207_),
    .Q_N(_1155_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[12] ));
 sg13g2_dfrbp_1 _2657_ (.CLK(net115),
    .RESET_B(net158),
    .D(_0208_),
    .Q_N(_1154_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[13] ));
 sg13g2_dfrbp_1 _2658_ (.CLK(net115),
    .RESET_B(net158),
    .D(_0209_),
    .Q_N(_1153_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[14] ));
 sg13g2_dfrbp_1 _2659_ (.CLK(net115),
    .RESET_B(net158),
    .D(_0210_),
    .Q_N(_1152_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[15] ));
 sg13g2_dfrbp_1 _2660_ (.CLK(net105),
    .RESET_B(net150),
    .D(_0211_),
    .Q_N(_1151_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[16] ));
 sg13g2_dfrbp_1 _2661_ (.CLK(net105),
    .RESET_B(net150),
    .D(_0212_),
    .Q_N(_1150_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[17] ));
 sg13g2_dfrbp_1 _2662_ (.CLK(net102),
    .RESET_B(net151),
    .D(_0213_),
    .Q_N(_1149_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[18] ));
 sg13g2_dfrbp_1 _2663_ (.CLK(net105),
    .RESET_B(net150),
    .D(_0214_),
    .Q_N(_1148_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[19] ));
 sg13g2_dfrbp_1 _2664_ (.CLK(net102),
    .RESET_B(net151),
    .D(_0215_),
    .Q_N(_1147_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[20] ));
 sg13g2_dfrbp_1 _2665_ (.CLK(net98),
    .RESET_B(net146),
    .D(_0216_),
    .Q_N(_1146_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[21] ));
 sg13g2_dfrbp_1 _2666_ (.CLK(net99),
    .RESET_B(net147),
    .D(_0217_),
    .Q_N(_1145_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[22] ));
 sg13g2_dfrbp_1 _2667_ (.CLK(net107),
    .RESET_B(net152),
    .D(_0218_),
    .Q_N(_1144_),
    .Q(\u_top_module.u_cic.u_differentiator.temp[23] ));
 sg13g2_dfrbp_1 _2668_ (.CLK(net126),
    .RESET_B(net168),
    .D(_0219_),
    .Q_N(_1143_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[0] ));
 sg13g2_dfrbp_1 _2669_ (.CLK(net127),
    .RESET_B(net166),
    .D(_0220_),
    .Q_N(_0036_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[1] ));
 sg13g2_dfrbp_1 _2670_ (.CLK(net128),
    .RESET_B(net168),
    .D(_0221_),
    .Q_N(_1142_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[2] ));
 sg13g2_dfrbp_1 _2671_ (.CLK(net130),
    .RESET_B(net167),
    .D(_0222_),
    .Q_N(_0038_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[3] ));
 sg13g2_dfrbp_1 _2672_ (.CLK(net130),
    .RESET_B(net167),
    .D(_0223_),
    .Q_N(_1141_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[4] ));
 sg13g2_dfrbp_1 _2673_ (.CLK(net125),
    .RESET_B(net165),
    .D(_0224_),
    .Q_N(_0040_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[5] ));
 sg13g2_dfrbp_1 _2674_ (.CLK(net123),
    .RESET_B(net164),
    .D(_0225_),
    .Q_N(_1140_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[6] ));
 sg13g2_dfrbp_1 _2675_ (.CLK(net122),
    .RESET_B(net163),
    .D(_0226_),
    .Q_N(_0042_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[7] ));
 sg13g2_dfrbp_1 _2676_ (.CLK(net110),
    .RESET_B(net155),
    .D(_0227_),
    .Q_N(_1139_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[8] ));
 sg13g2_dfrbp_1 _2677_ (.CLK(net110),
    .RESET_B(net155),
    .D(_0228_),
    .Q_N(_0044_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[9] ));
 sg13g2_dfrbp_1 _2678_ (.CLK(net109),
    .RESET_B(net154),
    .D(_0229_),
    .Q_N(_1138_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[10] ));
 sg13g2_dfrbp_1 _2679_ (.CLK(net118),
    .RESET_B(net160),
    .D(_0230_),
    .Q_N(_0046_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[11] ));
 sg13g2_dfrbp_1 _2680_ (.CLK(net114),
    .RESET_B(net159),
    .D(_0231_),
    .Q_N(_1137_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[12] ));
 sg13g2_dfrbp_1 _2681_ (.CLK(net115),
    .RESET_B(net158),
    .D(_0232_),
    .Q_N(_0048_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[13] ));
 sg13g2_dfrbp_1 _2682_ (.CLK(net113),
    .RESET_B(net159),
    .D(_0233_),
    .Q_N(_1136_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[14] ));
 sg13g2_dfrbp_1 _2683_ (.CLK(net115),
    .RESET_B(net158),
    .D(_0234_),
    .Q_N(_0050_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[15] ));
 sg13g2_dfrbp_1 _2684_ (.CLK(net104),
    .RESET_B(net151),
    .D(_0235_),
    .Q_N(_1135_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[16] ));
 sg13g2_dfrbp_1 _2685_ (.CLK(net105),
    .RESET_B(net150),
    .D(_0236_),
    .Q_N(_0052_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[17] ));
 sg13g2_dfrbp_1 _2686_ (.CLK(net103),
    .RESET_B(net151),
    .D(_0237_),
    .Q_N(_1134_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[18] ));
 sg13g2_dfrbp_1 _2687_ (.CLK(net105),
    .RESET_B(net150),
    .D(_0238_),
    .Q_N(_0054_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[19] ));
 sg13g2_dfrbp_1 _2688_ (.CLK(net102),
    .RESET_B(net151),
    .D(_0239_),
    .Q_N(_1133_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[20] ));
 sg13g2_dfrbp_1 _2689_ (.CLK(net97),
    .RESET_B(net146),
    .D(_0240_),
    .Q_N(_1132_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[21] ));
 sg13g2_dfrbp_1 _2690_ (.CLK(net99),
    .RESET_B(net147),
    .D(_0241_),
    .Q_N(_1131_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[22] ));
 sg13g2_dfrbp_1 _2691_ (.CLK(net107),
    .RESET_B(net152),
    .D(_0242_),
    .Q_N(_1130_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d3[23] ));
 sg13g2_dfrbp_1 _2692_ (.CLK(net126),
    .RESET_B(net248),
    .D(_0243_),
    .Q_N(_1129_),
    .Q(\u_top_module.u_i2s_bus.u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2693_ (.CLK(net127),
    .RESET_B(net246),
    .D(_0244_),
    .Q_N(_1128_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[1].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2694_ (.CLK(net128),
    .RESET_B(net244),
    .D(_0245_),
    .Q_N(_1127_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[2].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2695_ (.CLK(net129),
    .RESET_B(net242),
    .D(_0246_),
    .Q_N(_1126_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[3].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2696_ (.CLK(net129),
    .RESET_B(net240),
    .D(_0247_),
    .Q_N(_1125_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[4].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2697_ (.CLK(net130),
    .RESET_B(net238),
    .D(_0248_),
    .Q_N(_1124_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[5].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2698_ (.CLK(net137),
    .RESET_B(net236),
    .D(_0249_),
    .Q_N(_1123_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[6].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2699_ (.CLK(net126),
    .RESET_B(net234),
    .D(_0250_),
    .Q_N(_1122_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[7].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2700_ (.CLK(net117),
    .RESET_B(net232),
    .D(_0251_),
    .Q_N(_1121_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[8].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2701_ (.CLK(net117),
    .RESET_B(net230),
    .D(_0252_),
    .Q_N(_1120_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[9].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2702_ (.CLK(net116),
    .RESET_B(net228),
    .D(_0253_),
    .Q_N(_1119_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[10].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2703_ (.CLK(net116),
    .RESET_B(net226),
    .D(_0254_),
    .Q_N(_1118_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[11].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2704_ (.CLK(net114),
    .RESET_B(net224),
    .D(_0255_),
    .Q_N(_1117_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[12].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2705_ (.CLK(net114),
    .RESET_B(net221),
    .D(_0256_),
    .Q_N(_1116_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[13].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2706_ (.CLK(net113),
    .RESET_B(net219),
    .D(_0257_),
    .Q_N(_1115_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[14].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2707_ (.CLK(net106),
    .RESET_B(net217),
    .D(_0258_),
    .Q_N(_1114_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[15].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2708_ (.CLK(net104),
    .RESET_B(net215),
    .D(_0259_),
    .Q_N(_1113_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[16].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2709_ (.CLK(net106),
    .RESET_B(net213),
    .D(_0260_),
    .Q_N(_1112_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[17].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2710_ (.CLK(net103),
    .RESET_B(net211),
    .D(_0261_),
    .Q_N(_1111_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[18].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2711_ (.CLK(net102),
    .RESET_B(net209),
    .D(_0262_),
    .Q_N(_1110_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[19].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2712_ (.CLK(net102),
    .RESET_B(net207),
    .D(_0263_),
    .Q_N(_1109_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[20].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2713_ (.CLK(net97),
    .RESET_B(net205),
    .D(_0264_),
    .Q_N(_1108_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[21].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2714_ (.CLK(net99),
    .RESET_B(net203),
    .D(_0265_),
    .Q_N(_1107_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[22].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2715_ (.CLK(net122),
    .RESET_B(net202),
    .D(_0266_),
    .Q_N(_1106_),
    .Q(\u_top_module.u_i2s_bus.mux_shift_inst[23].u_mux_shift.sum_res ));
 sg13g2_dfrbp_1 _2716_ (.CLK(net138),
    .RESET_B(net172),
    .D(_0267_),
    .Q_N(_1105_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[1] ));
 sg13g2_dfrbp_1 _2717_ (.CLK(net138),
    .RESET_B(net172),
    .D(_0268_),
    .Q_N(_1104_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[2] ));
 sg13g2_dfrbp_1 _2718_ (.CLK(net138),
    .RESET_B(net172),
    .D(_0269_),
    .Q_N(_1103_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[3] ));
 sg13g2_dfrbp_1 _2719_ (.CLK(net133),
    .RESET_B(net171),
    .D(_0270_),
    .Q_N(_1102_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[4] ));
 sg13g2_dfrbp_1 _2720_ (.CLK(net125),
    .RESET_B(net165),
    .D(_0271_),
    .Q_N(_1101_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[5] ));
 sg13g2_dfrbp_1 _2721_ (.CLK(net123),
    .RESET_B(net164),
    .D(_0272_),
    .Q_N(_1100_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[6] ));
 sg13g2_dfrbp_1 _2722_ (.CLK(net125),
    .RESET_B(net163),
    .D(_0273_),
    .Q_N(_1099_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[7] ));
 sg13g2_dfrbp_1 _2723_ (.CLK(net125),
    .RESET_B(net163),
    .D(_0274_),
    .Q_N(_1098_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[8] ));
 sg13g2_dfrbp_1 _2724_ (.CLK(net110),
    .RESET_B(net157),
    .D(_0275_),
    .Q_N(_1097_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[9] ));
 sg13g2_dfrbp_1 _2725_ (.CLK(net109),
    .RESET_B(net155),
    .D(_0276_),
    .Q_N(_1096_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[10] ));
 sg13g2_dfrbp_1 _2726_ (.CLK(net109),
    .RESET_B(net155),
    .D(_0277_),
    .Q_N(_1095_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[11] ));
 sg13g2_dfrbp_1 _2727_ (.CLK(net107),
    .RESET_B(net154),
    .D(_0278_),
    .Q_N(_1094_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[12] ));
 sg13g2_dfrbp_1 _2728_ (.CLK(net112),
    .RESET_B(net154),
    .D(_0279_),
    .Q_N(_1093_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[13] ));
 sg13g2_dfrbp_1 _2729_ (.CLK(net112),
    .RESET_B(net152),
    .D(_0280_),
    .Q_N(_1092_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[14] ));
 sg13g2_dfrbp_1 _2730_ (.CLK(net107),
    .RESET_B(net152),
    .D(_0281_),
    .Q_N(_1091_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[15] ));
 sg13g2_dfrbp_1 _2731_ (.CLK(net99),
    .RESET_B(net147),
    .D(_0282_),
    .Q_N(_1090_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[16] ));
 sg13g2_dfrbp_1 _2732_ (.CLK(net99),
    .RESET_B(net147),
    .D(_0283_),
    .Q_N(_1089_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[17] ));
 sg13g2_dfrbp_1 _2733_ (.CLK(net98),
    .RESET_B(net146),
    .D(_0284_),
    .Q_N(_1088_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[18] ));
 sg13g2_dfrbp_1 _2734_ (.CLK(net99),
    .RESET_B(net147),
    .D(_0285_),
    .Q_N(_1087_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[19] ));
 sg13g2_dfrbp_1 _2735_ (.CLK(net98),
    .RESET_B(net146),
    .D(_0286_),
    .Q_N(_1086_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[20] ));
 sg13g2_dfrbp_1 _2736_ (.CLK(net97),
    .RESET_B(net146),
    .D(_0287_),
    .Q_N(_1085_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[21] ));
 sg13g2_dfrbp_1 _2737_ (.CLK(net97),
    .RESET_B(net149),
    .D(_0288_),
    .Q_N(_1084_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[22] ));
 sg13g2_dfrbp_1 _2738_ (.CLK(net101),
    .RESET_B(net149),
    .D(_0289_),
    .Q_N(_1319_),
    .Q(\u_top_module.u_cic.u_differentiator.a_mux4to1.d1[23] ));
 sg13g2_dfrbp_1 _2739_ (.CLK(net133),
    .RESET_B(net171),
    .D(net11),
    .Q_N(_1083_),
    .Q(\u_top_module.u_cic.u_differentiator.prev_lr_clk ));
 sg13g2_dfrbp_1 _2740_ (.CLK(_0158_),
    .RESET_B(net176),
    .D(net3),
    .Q_N(_1082_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[1].u_ddr_to_sdr.ddr_data_falling ));
 sg13g2_dfrbp_1 _2741_ (.CLK(_0159_),
    .RESET_B(net172),
    .D(net4),
    .Q_N(_1081_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[2].u_ddr_to_sdr.ddr_data_falling ));
 sg13g2_dfrbp_1 _2742_ (.CLK(_0160_),
    .RESET_B(net172),
    .D(net5),
    .Q_N(_1080_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[3].u_ddr_to_sdr.ddr_data_falling ));
 sg13g2_dfrbp_1 _2743_ (.CLK(_0161_),
    .RESET_B(net174),
    .D(net6),
    .Q_N(_1079_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[4].u_ddr_to_sdr.ddr_data_falling ));
 sg13g2_dfrbp_1 _2744_ (.CLK(_0162_),
    .RESET_B(net174),
    .D(net7),
    .Q_N(_1078_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.ddr_data_falling ));
 sg13g2_dfrbp_1 _2745_ (.CLK(_0163_),
    .RESET_B(net175),
    .D(net8),
    .Q_N(_1077_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[6].u_ddr_to_sdr.ddr_data_falling ));
 sg13g2_dfrbp_1 _2746_ (.CLK(_0164_),
    .RESET_B(net176),
    .D(net9),
    .Q_N(_1320_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[7].u_ddr_to_sdr.ddr_data_falling ));
 sg13g2_dfrbp_1 _2747_ (.CLK(net141),
    .RESET_B(net176),
    .D(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.ddr_data_falling ),
    .Q_N(_1321_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.sdr_data_1 ));
 sg13g2_dfrbp_1 _2748_ (.CLK(net141),
    .RESET_B(net176),
    .D(net2),
    .Q_N(_1322_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.ddr_data_rising ));
 sg13g2_dfrbp_1 _2749_ (.CLK(net141),
    .RESET_B(net176),
    .D(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.ddr_data_rising ),
    .Q_N(_1323_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.sdr_data_0 ));
 sg13g2_dfrbp_1 _2750_ (.CLK(net141),
    .RESET_B(net176),
    .D(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[1].u_ddr_to_sdr.ddr_data_falling ),
    .Q_N(_1324_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[1].u_ddr_to_sdr.sdr_data_1 ));
 sg13g2_dfrbp_1 _2751_ (.CLK(net141),
    .RESET_B(net176),
    .D(net3),
    .Q_N(_1325_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[1].u_ddr_to_sdr.ddr_data_rising ));
 sg13g2_dfrbp_1 _2752_ (.CLK(net141),
    .RESET_B(net176),
    .D(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[1].u_ddr_to_sdr.ddr_data_rising ),
    .Q_N(_1326_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[1].u_ddr_to_sdr.sdr_data_0 ));
 sg13g2_dfrbp_1 _2753_ (.CLK(net137),
    .RESET_B(net172),
    .D(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[2].u_ddr_to_sdr.ddr_data_falling ),
    .Q_N(_1327_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[2].u_ddr_to_sdr.sdr_data_1 ));
 sg13g2_dfrbp_1 _2754_ (.CLK(net137),
    .RESET_B(net172),
    .D(net4),
    .Q_N(_1328_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[2].u_ddr_to_sdr.ddr_data_rising ));
 sg13g2_dfrbp_1 _2755_ (.CLK(net138),
    .RESET_B(net173),
    .D(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[2].u_ddr_to_sdr.ddr_data_rising ),
    .Q_N(_0032_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[2].u_ddr_to_sdr.sdr_data_0 ));
 sg13g2_dfrbp_1 _2756_ (.CLK(net138),
    .RESET_B(net173),
    .D(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[3].u_ddr_to_sdr.ddr_data_falling ),
    .Q_N(_0033_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[3].u_ddr_to_sdr.sdr_data_1 ));
 sg13g2_dfrbp_1 _2757_ (.CLK(net137),
    .RESET_B(net173),
    .D(net5),
    .Q_N(_1329_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[3].u_ddr_to_sdr.ddr_data_rising ));
 sg13g2_dfrbp_1 _2758_ (.CLK(net137),
    .RESET_B(net173),
    .D(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[3].u_ddr_to_sdr.ddr_data_rising ),
    .Q_N(_1330_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[3].u_ddr_to_sdr.sdr_data_0 ));
 sg13g2_dfrbp_1 _2759_ (.CLK(net139),
    .RESET_B(net174),
    .D(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[4].u_ddr_to_sdr.ddr_data_falling ),
    .Q_N(_1331_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[4].u_ddr_to_sdr.sdr_data_1 ));
 sg13g2_dfrbp_1 _2760_ (.CLK(net139),
    .RESET_B(net174),
    .D(net6),
    .Q_N(_1332_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[4].u_ddr_to_sdr.ddr_data_rising ));
 sg13g2_dfrbp_1 _2761_ (.CLK(net139),
    .RESET_B(net174),
    .D(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[4].u_ddr_to_sdr.ddr_data_rising ),
    .Q_N(_1333_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[4].u_ddr_to_sdr.sdr_data_0 ));
 sg13g2_dfrbp_1 _2762_ (.CLK(net140),
    .RESET_B(net174),
    .D(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.ddr_data_falling ),
    .Q_N(_1334_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.sdr_data_1 ));
 sg13g2_dfrbp_1 _2763_ (.CLK(net139),
    .RESET_B(net174),
    .D(net7),
    .Q_N(_1335_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.ddr_data_rising ));
 sg13g2_dfrbp_1 _2764_ (.CLK(net140),
    .RESET_B(net175),
    .D(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.ddr_data_rising ),
    .Q_N(_1336_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[5].u_ddr_to_sdr.sdr_data_0 ));
 sg13g2_dfrbp_1 _2765_ (.CLK(net140),
    .RESET_B(net175),
    .D(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[6].u_ddr_to_sdr.ddr_data_falling ),
    .Q_N(_0034_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[6].u_ddr_to_sdr.sdr_data_1 ));
 sg13g2_dfrbp_1 _2766_ (.CLK(net139),
    .RESET_B(net174),
    .D(net8),
    .Q_N(_1337_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[6].u_ddr_to_sdr.ddr_data_rising ));
 sg13g2_dfrbp_1 _2767_ (.CLK(net140),
    .RESET_B(net175),
    .D(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[6].u_ddr_to_sdr.ddr_data_rising ),
    .Q_N(_1338_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[6].u_ddr_to_sdr.sdr_data_0 ));
 sg13g2_dfrbp_1 _2768_ (.CLK(net142),
    .RESET_B(net177),
    .D(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[7].u_ddr_to_sdr.ddr_data_falling ),
    .Q_N(_1339_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[7].u_ddr_to_sdr.sdr_data_1 ));
 sg13g2_dfrbp_1 _2769_ (.CLK(net135),
    .RESET_B(net171),
    .D(net9),
    .Q_N(_1340_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[7].u_ddr_to_sdr.ddr_data_rising ));
 sg13g2_dfrbp_1 _2770_ (.CLK(net140),
    .RESET_B(net175),
    .D(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[7].u_ddr_to_sdr.ddr_data_rising ),
    .Q_N(_0031_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[7].u_ddr_to_sdr.sdr_data_0 ));
 sg13g2_dfrbp_1 _2771_ (.CLK(_0165_),
    .RESET_B(net177),
    .D(net2),
    .Q_N(_1076_),
    .Q(\u_top_module.u_multi_ddr_to_sdr.ddr_to_sdr_inst[0].u_ddr_to_sdr.ddr_data_falling ));
 sg13g2_tiehi _2714__203 (.L_HI(net203));
 sg13g2_tiehi _2482__204 (.L_HI(net204));
 sg13g2_tiehi _2713__205 (.L_HI(net205));
 sg13g2_tiehi _2487__206 (.L_HI(net206));
 sg13g2_tiehi _2712__207 (.L_HI(net207));
 sg13g2_tiehi _2489__208 (.L_HI(net208));
 sg13g2_tiehi _2711__209 (.L_HI(net209));
 sg13g2_tiehi _2491__210 (.L_HI(net210));
 sg13g2_tiehi _2710__211 (.L_HI(net211));
 sg13g2_tiehi _2493__212 (.L_HI(net212));
 sg13g2_tiehi _2709__213 (.L_HI(net213));
 sg13g2_tiehi _2495__214 (.L_HI(net214));
 sg13g2_tiehi _2708__215 (.L_HI(net215));
 sg13g2_tiehi _2497__216 (.L_HI(net216));
 sg13g2_tiehi _2707__217 (.L_HI(net217));
 sg13g2_tiehi _2499__218 (.L_HI(net218));
 sg13g2_tiehi _2706__219 (.L_HI(net219));
 sg13g2_tiehi _2501__220 (.L_HI(net220));
 sg13g2_tiehi _2705__221 (.L_HI(net221));
 sg13g2_tiehi _2503__222 (.L_HI(net222));
 sg13g2_tiehi _2505__223 (.L_HI(net223));
 sg13g2_tiehi _2704__224 (.L_HI(net224));
 sg13g2_tiehi _2506__225 (.L_HI(net225));
 sg13g2_tiehi _2703__226 (.L_HI(net226));
 sg13g2_tiehi _2508__227 (.L_HI(net227));
 sg13g2_tiehi _2702__228 (.L_HI(net228));
 sg13g2_tiehi _2510__229 (.L_HI(net229));
 sg13g2_tiehi _2701__230 (.L_HI(net230));
 sg13g2_tiehi _2512__231 (.L_HI(net231));
 sg13g2_tiehi _2700__232 (.L_HI(net232));
 sg13g2_tiehi _2514__233 (.L_HI(net233));
 sg13g2_tiehi _2699__234 (.L_HI(net234));
 sg13g2_tiehi _2516__235 (.L_HI(net235));
 sg13g2_tiehi _2698__236 (.L_HI(net236));
 sg13g2_tiehi _2518__237 (.L_HI(net237));
 sg13g2_tiehi _2697__238 (.L_HI(net238));
 sg13g2_tiehi _2520__239 (.L_HI(net239));
 sg13g2_tiehi _2696__240 (.L_HI(net240));
 sg13g2_tiehi _2522__241 (.L_HI(net241));
 sg13g2_tiehi _2695__242 (.L_HI(net242));
 sg13g2_tiehi _2524__243 (.L_HI(net243));
 sg13g2_tiehi _2694__244 (.L_HI(net244));
 sg13g2_tiehi _2526__245 (.L_HI(net245));
 sg13g2_tiehi _2693__246 (.L_HI(net246));
 sg13g2_tiehi _2528__247 (.L_HI(net247));
 sg13g2_tiehi _2692__248 (.L_HI(net248));
 sg13g2_tiehi _2530__249 (.L_HI(net249));
 sg13g2_tiehi _2532__250 (.L_HI(net250));
 sg13g2_tiehi _2534__251 (.L_HI(net251));
 sg13g2_tiehi _2536__252 (.L_HI(net252));
 sg13g2_tiehi _2538__253 (.L_HI(net253));
 sg13g2_tiehi _2540__254 (.L_HI(net254));
 sg13g2_tiehi _2542__255 (.L_HI(net255));
 sg13g2_tiehi _2544__256 (.L_HI(net256));
 sg13g2_tiehi _2546__257 (.L_HI(net257));
 sg13g2_tiehi _2548__258 (.L_HI(net258));
 sg13g2_tiehi _2550__259 (.L_HI(net259));
 sg13g2_tiehi _2549__260 (.L_HI(net260));
 sg13g2_tiehi _2547__261 (.L_HI(net261));
 sg13g2_tiehi _2545__262 (.L_HI(net262));
 sg13g2_tiehi _2543__263 (.L_HI(net263));
 sg13g2_tiehi _2541__264 (.L_HI(net264));
 sg13g2_tiehi _2539__265 (.L_HI(net265));
 sg13g2_tiehi _2537__266 (.L_HI(net266));
 sg13g2_tiehi _2535__267 (.L_HI(net267));
 sg13g2_tiehi _2533__268 (.L_HI(net268));
 sg13g2_tiehi _2531__269 (.L_HI(net269));
 sg13g2_tiehi _2529__270 (.L_HI(net270));
 sg13g2_tiehi _2527__271 (.L_HI(net271));
 sg13g2_tiehi _2525__272 (.L_HI(net272));
 sg13g2_tiehi _2523__273 (.L_HI(net273));
 sg13g2_tiehi _2521__274 (.L_HI(net274));
 sg13g2_tiehi _2519__275 (.L_HI(net275));
 sg13g2_tiehi _2517__276 (.L_HI(net276));
 sg13g2_tiehi _2515__277 (.L_HI(net277));
 sg13g2_tiehi _2513__278 (.L_HI(net278));
 sg13g2_tiehi _2511__279 (.L_HI(net279));
 sg13g2_tiehi _2509__280 (.L_HI(net280));
 sg13g2_tiehi _2507__281 (.L_HI(net281));
 sg13g2_tiehi _2504__282 (.L_HI(net282));
 sg13g2_tiehi _2502__283 (.L_HI(net283));
 sg13g2_tiehi _2500__284 (.L_HI(net284));
 sg13g2_tiehi _2498__285 (.L_HI(net285));
 sg13g2_tiehi _2496__286 (.L_HI(net286));
 sg13g2_tiehi _2494__287 (.L_HI(net287));
 sg13g2_tiehi _2492__288 (.L_HI(net288));
 sg13g2_tiehi _2490__289 (.L_HI(net289));
 sg13g2_tiehi _2488__290 (.L_HI(net290));
 sg13g2_tiehi _2486__291 (.L_HI(net291));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_180 (.L_LO(net180));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_181 (.L_LO(net181));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_182 (.L_LO(net182));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_183 (.L_LO(net183));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_184 (.L_LO(net184));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_185 (.L_LO(net185));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_186 (.L_LO(net186));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_187 (.L_LO(net187));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_188 (.L_LO(net188));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_189 (.L_LO(net189));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_190 (.L_LO(net190));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_191 (.L_LO(net191));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_192 (.L_LO(net192));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_193 (.L_LO(net193));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_194 (.L_LO(net194));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_195 (.L_LO(net195));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_196 (.L_LO(net196));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_197 (.L_LO(net197));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_198 (.L_LO(net198));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_199 (.L_LO(net199));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_200 (.L_LO(net200));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_201 (.L_LO(net201));
 sg13g2_tiehi _2715__202 (.L_HI(net202));
 sg13g2_buf_1 _2885_ (.A(out),
    .X(uo_out[0]));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[1]),
    .X(net11));
 sg13g2_buf_4 fanout12 (.X(net12),
    .A(net15));
 sg13g2_buf_1 fanout13 (.A(net15),
    .X(net13));
 sg13g2_buf_4 fanout14 (.X(net14),
    .A(net15));
 sg13g2_buf_2 fanout15 (.A(net17),
    .X(net15));
 sg13g2_buf_4 fanout16 (.X(net16),
    .A(net17));
 sg13g2_buf_4 fanout17 (.X(net17),
    .A(_1048_));
 sg13g2_buf_4 fanout18 (.X(net18),
    .A(net21));
 sg13g2_buf_2 fanout19 (.A(net21),
    .X(net19));
 sg13g2_buf_4 fanout20 (.X(net20),
    .A(net21));
 sg13g2_buf_4 fanout21 (.X(net21),
    .A(_0698_));
 sg13g2_buf_2 fanout22 (.A(net23),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(net30),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(net30),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(net29),
    .X(net25));
 sg13g2_buf_1 fanout26 (.A(net29),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(net28),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(net29),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(net30),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0673_),
    .X(net30));
 sg13g2_buf_4 fanout31 (.X(net31),
    .A(net34));
 sg13g2_buf_1 fanout32 (.A(net34),
    .X(net32));
 sg13g2_buf_4 fanout33 (.X(net33),
    .A(net34));
 sg13g2_buf_4 fanout34 (.X(net34),
    .A(_0566_));
 sg13g2_buf_4 fanout35 (.X(net35),
    .A(net39));
 sg13g2_buf_1 fanout36 (.A(net39),
    .X(net36));
 sg13g2_buf_4 fanout37 (.X(net37),
    .A(net39));
 sg13g2_buf_2 fanout38 (.A(net39),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0565_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(net44),
    .X(net40));
 sg13g2_buf_1 fanout41 (.A(net44),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(net44),
    .X(net42));
 sg13g2_buf_1 fanout43 (.A(net44),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0358_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(net48),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(net47),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(net48),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0358_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(net53),
    .X(net49));
 sg13g2_buf_1 fanout50 (.A(net53),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(net53),
    .X(net51));
 sg13g2_buf_1 fanout52 (.A(net53),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0357_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(net57),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(net56),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(net57),
    .X(net56));
 sg13g2_buf_1 fanout57 (.A(_0357_),
    .X(net57));
 sg13g2_buf_4 fanout58 (.X(net58),
    .A(_0356_));
 sg13g2_buf_2 fanout59 (.A(_0356_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(net61),
    .X(net60));
 sg13g2_buf_4 fanout61 (.X(net61),
    .A(net64));
 sg13g2_buf_4 fanout62 (.X(net62),
    .A(net63));
 sg13g2_buf_4 fanout63 (.X(net63),
    .A(net64));
 sg13g2_buf_2 fanout64 (.A(_0355_),
    .X(net64));
 sg13g2_buf_4 fanout65 (.X(net65),
    .A(_0354_));
 sg13g2_buf_4 fanout66 (.X(net66),
    .A(_0353_));
 sg13g2_buf_4 fanout67 (.X(net67),
    .A(_0353_));
 sg13g2_buf_4 fanout68 (.X(net68),
    .A(net69));
 sg13g2_buf_4 fanout69 (.X(net69),
    .A(_0352_));
 sg13g2_buf_2 fanout70 (.A(_0740_),
    .X(net70));
 sg13g2_buf_4 fanout71 (.X(net71),
    .A(net74));
 sg13g2_buf_4 fanout72 (.X(net72),
    .A(net74));
 sg13g2_buf_1 fanout73 (.A(net74),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0350_),
    .X(net74));
 sg13g2_buf_4 fanout75 (.X(net75),
    .A(_0347_));
 sg13g2_buf_2 fanout76 (.A(_0347_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0739_),
    .X(net77));
 sg13g2_buf_4 fanout78 (.X(net78),
    .A(net81));
 sg13g2_buf_4 fanout79 (.X(net79),
    .A(net81));
 sg13g2_buf_2 fanout80 (.A(net81),
    .X(net80));
 sg13g2_buf_4 fanout81 (.X(net81),
    .A(_0738_));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(net86));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(net86));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(net86));
 sg13g2_buf_2 fanout85 (.A(net86),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.sel[1] ),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(net88),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(net95),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(net95),
    .X(net89));
 sg13g2_buf_1 fanout90 (.A(net95),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(net95),
    .X(net91));
 sg13g2_buf_1 fanout92 (.A(net95),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(net94),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(net95),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(\u_top_module.u_cic.u_differentiator.a_mux4to1.sel[0] ),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(net98),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(net98),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(net101),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(net101),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(net101),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(net120),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(net106),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(net106),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(net105),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(net106),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(net120),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(net112),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(net112),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(net112),
    .X(net109));
 sg13g2_buf_1 fanout110 (.A(net111),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(net112),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(net120),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(net119),
    .X(net113));
 sg13g2_buf_1 fanout114 (.A(net119),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(net119),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(net118),
    .X(net116));
 sg13g2_buf_1 fanout117 (.A(net118),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(net119),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(net120),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(net10),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(net122),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(net125),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(net124),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(net125),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(net143),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(net127),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(net131),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(net131),
    .X(net128));
 sg13g2_buf_1 fanout129 (.A(net131),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(net131),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(net143),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(net136),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(net136),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(net136),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(net136),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(net143),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(net138),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(net142),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(net142),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(net142),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(net143),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(net10),
    .X(net143));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(net146));
 sg13g2_buf_2 fanout145 (.A(net146),
    .X(net145));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(net149));
 sg13g2_buf_4 fanout147 (.X(net147),
    .A(net149));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(net149));
 sg13g2_buf_2 fanout149 (.A(net161),
    .X(net149));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(net151));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(net161));
 sg13g2_buf_4 fanout152 (.X(net152),
    .A(net154));
 sg13g2_buf_4 fanout153 (.X(net153),
    .A(net157));
 sg13g2_buf_2 fanout154 (.A(net157),
    .X(net154));
 sg13g2_buf_4 fanout155 (.X(net155),
    .A(net157));
 sg13g2_buf_4 fanout156 (.X(net156),
    .A(net157));
 sg13g2_buf_2 fanout157 (.A(net161),
    .X(net157));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(net160));
 sg13g2_buf_2 fanout159 (.A(net160),
    .X(net159));
 sg13g2_buf_4 fanout160 (.X(net160),
    .A(net161));
 sg13g2_buf_2 fanout161 (.A(net1),
    .X(net161));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(net169));
 sg13g2_buf_4 fanout163 (.X(net163),
    .A(net169));
 sg13g2_buf_4 fanout164 (.X(net164),
    .A(net165));
 sg13g2_buf_4 fanout165 (.X(net165),
    .A(net169));
 sg13g2_buf_4 fanout166 (.X(net166),
    .A(net168));
 sg13g2_buf_4 fanout167 (.X(net167),
    .A(net168));
 sg13g2_buf_2 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(net1),
    .X(net169));
 sg13g2_buf_4 fanout170 (.X(net170),
    .A(net171));
 sg13g2_buf_4 fanout171 (.X(net171),
    .A(net178));
 sg13g2_buf_4 fanout172 (.X(net172),
    .A(net178));
 sg13g2_buf_2 fanout173 (.A(net178),
    .X(net173));
 sg13g2_buf_4 fanout174 (.X(net174),
    .A(net175));
 sg13g2_buf_4 fanout175 (.X(net175),
    .A(net177));
 sg13g2_buf_4 fanout176 (.X(net176),
    .A(net177));
 sg13g2_buf_2 fanout177 (.A(net178),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(net1),
    .X(net178));
 sg13g2_tielo tt_um_16_mic_beamformer_arghunter_179 (.L_LO(net179));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_4 FILLER_0_147 ();
 sg13g2_fill_1 FILLER_0_151 ();
 sg13g2_decap_8 FILLER_0_165 ();
 sg13g2_decap_8 FILLER_0_172 ();
 sg13g2_decap_4 FILLER_0_179 ();
 sg13g2_fill_1 FILLER_0_183 ();
 sg13g2_decap_8 FILLER_0_192 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_decap_8 FILLER_0_206 ();
 sg13g2_decap_8 FILLER_0_213 ();
 sg13g2_decap_8 FILLER_0_220 ();
 sg13g2_decap_8 FILLER_0_227 ();
 sg13g2_decap_8 FILLER_0_234 ();
 sg13g2_decap_4 FILLER_0_245 ();
 sg13g2_fill_1 FILLER_0_254 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_4 FILLER_1_126 ();
 sg13g2_fill_2 FILLER_1_156 ();
 sg13g2_fill_1 FILLER_1_158 ();
 sg13g2_decap_8 FILLER_1_193 ();
 sg13g2_decap_8 FILLER_1_226 ();
 sg13g2_decap_4 FILLER_1_233 ();
 sg13g2_fill_2 FILLER_1_242 ();
 sg13g2_fill_2 FILLER_1_270 ();
 sg13g2_fill_1 FILLER_1_272 ();
 sg13g2_fill_2 FILLER_1_282 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_fill_2 FILLER_2_119 ();
 sg13g2_fill_2 FILLER_2_155 ();
 sg13g2_fill_1 FILLER_2_157 ();
 sg13g2_fill_1 FILLER_2_184 ();
 sg13g2_fill_2 FILLER_2_263 ();
 sg13g2_fill_2 FILLER_2_310 ();
 sg13g2_fill_1 FILLER_2_312 ();
 sg13g2_fill_1 FILLER_2_317 ();
 sg13g2_decap_4 FILLER_2_350 ();
 sg13g2_fill_2 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_360 ();
 sg13g2_decap_8 FILLER_2_367 ();
 sg13g2_decap_8 FILLER_2_374 ();
 sg13g2_decap_8 FILLER_2_381 ();
 sg13g2_decap_8 FILLER_2_388 ();
 sg13g2_decap_8 FILLER_2_395 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_fill_2 FILLER_3_119 ();
 sg13g2_fill_1 FILLER_3_121 ();
 sg13g2_fill_2 FILLER_3_146 ();
 sg13g2_fill_1 FILLER_3_148 ();
 sg13g2_fill_2 FILLER_3_170 ();
 sg13g2_fill_1 FILLER_3_172 ();
 sg13g2_fill_2 FILLER_3_219 ();
 sg13g2_fill_1 FILLER_3_225 ();
 sg13g2_fill_1 FILLER_3_266 ();
 sg13g2_fill_2 FILLER_3_293 ();
 sg13g2_decap_8 FILLER_3_299 ();
 sg13g2_decap_8 FILLER_3_306 ();
 sg13g2_decap_4 FILLER_3_321 ();
 sg13g2_fill_2 FILLER_3_339 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_4 FILLER_4_126 ();
 sg13g2_fill_2 FILLER_4_130 ();
 sg13g2_decap_8 FILLER_4_141 ();
 sg13g2_decap_8 FILLER_4_148 ();
 sg13g2_decap_4 FILLER_4_168 ();
 sg13g2_fill_2 FILLER_4_172 ();
 sg13g2_decap_8 FILLER_4_192 ();
 sg13g2_decap_8 FILLER_4_199 ();
 sg13g2_decap_8 FILLER_4_206 ();
 sg13g2_decap_4 FILLER_4_213 ();
 sg13g2_fill_1 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_223 ();
 sg13g2_decap_4 FILLER_4_230 ();
 sg13g2_fill_2 FILLER_4_234 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_fill_1 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_286 ();
 sg13g2_decap_4 FILLER_4_293 ();
 sg13g2_fill_2 FILLER_4_328 ();
 sg13g2_decap_8 FILLER_4_356 ();
 sg13g2_decap_8 FILLER_4_363 ();
 sg13g2_decap_8 FILLER_4_370 ();
 sg13g2_decap_8 FILLER_4_377 ();
 sg13g2_decap_8 FILLER_4_384 ();
 sg13g2_decap_8 FILLER_4_391 ();
 sg13g2_decap_8 FILLER_4_398 ();
 sg13g2_decap_4 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_fill_1 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_164 ();
 sg13g2_fill_2 FILLER_5_171 ();
 sg13g2_decap_8 FILLER_5_190 ();
 sg13g2_decap_4 FILLER_5_197 ();
 sg13g2_fill_2 FILLER_5_201 ();
 sg13g2_decap_4 FILLER_5_239 ();
 sg13g2_fill_2 FILLER_5_243 ();
 sg13g2_fill_2 FILLER_5_248 ();
 sg13g2_fill_1 FILLER_5_250 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_4 FILLER_5_266 ();
 sg13g2_fill_2 FILLER_5_275 ();
 sg13g2_decap_4 FILLER_5_293 ();
 sg13g2_fill_2 FILLER_5_297 ();
 sg13g2_decap_8 FILLER_5_303 ();
 sg13g2_decap_4 FILLER_5_310 ();
 sg13g2_decap_8 FILLER_5_319 ();
 sg13g2_decap_8 FILLER_5_326 ();
 sg13g2_decap_8 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_340 ();
 sg13g2_decap_8 FILLER_5_347 ();
 sg13g2_decap_8 FILLER_5_354 ();
 sg13g2_decap_4 FILLER_5_361 ();
 sg13g2_decap_8 FILLER_5_369 ();
 sg13g2_decap_8 FILLER_5_376 ();
 sg13g2_decap_8 FILLER_5_383 ();
 sg13g2_decap_8 FILLER_5_390 ();
 sg13g2_decap_8 FILLER_5_397 ();
 sg13g2_decap_4 FILLER_5_404 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_fill_2 FILLER_6_126 ();
 sg13g2_fill_1 FILLER_6_146 ();
 sg13g2_fill_2 FILLER_6_207 ();
 sg13g2_fill_1 FILLER_6_209 ();
 sg13g2_fill_1 FILLER_6_236 ();
 sg13g2_decap_8 FILLER_6_328 ();
 sg13g2_decap_8 FILLER_6_335 ();
 sg13g2_decap_8 FILLER_6_342 ();
 sg13g2_fill_2 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_fill_1 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_163 ();
 sg13g2_decap_8 FILLER_7_170 ();
 sg13g2_fill_2 FILLER_7_186 ();
 sg13g2_fill_1 FILLER_7_188 ();
 sg13g2_fill_1 FILLER_7_233 ();
 sg13g2_fill_2 FILLER_7_340 ();
 sg13g2_decap_8 FILLER_7_368 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_4 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_4 FILLER_8_126 ();
 sg13g2_fill_2 FILLER_8_130 ();
 sg13g2_fill_2 FILLER_8_145 ();
 sg13g2_fill_1 FILLER_8_147 ();
 sg13g2_decap_4 FILLER_8_166 ();
 sg13g2_fill_2 FILLER_8_170 ();
 sg13g2_decap_8 FILLER_8_193 ();
 sg13g2_decap_8 FILLER_8_220 ();
 sg13g2_decap_8 FILLER_8_227 ();
 sg13g2_fill_2 FILLER_8_248 ();
 sg13g2_decap_4 FILLER_8_285 ();
 sg13g2_fill_1 FILLER_8_298 ();
 sg13g2_fill_1 FILLER_8_313 ();
 sg13g2_decap_8 FILLER_8_362 ();
 sg13g2_decap_8 FILLER_8_369 ();
 sg13g2_decap_8 FILLER_8_376 ();
 sg13g2_decap_8 FILLER_8_383 ();
 sg13g2_decap_8 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_decap_4 FILLER_8_404 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_230 ();
 sg13g2_fill_2 FILLER_9_237 ();
 sg13g2_fill_1 FILLER_9_239 ();
 sg13g2_fill_2 FILLER_9_244 ();
 sg13g2_fill_1 FILLER_9_246 ();
 sg13g2_decap_8 FILLER_9_256 ();
 sg13g2_decap_4 FILLER_9_263 ();
 sg13g2_fill_1 FILLER_9_267 ();
 sg13g2_fill_2 FILLER_9_272 ();
 sg13g2_decap_8 FILLER_9_278 ();
 sg13g2_decap_4 FILLER_9_285 ();
 sg13g2_fill_2 FILLER_9_289 ();
 sg13g2_fill_2 FILLER_9_301 ();
 sg13g2_fill_1 FILLER_9_303 ();
 sg13g2_fill_1 FILLER_9_329 ();
 sg13g2_fill_1 FILLER_9_356 ();
 sg13g2_decap_8 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_fill_2 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_145 ();
 sg13g2_decap_8 FILLER_10_164 ();
 sg13g2_decap_8 FILLER_10_171 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_fill_2 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_4 FILLER_10_224 ();
 sg13g2_fill_2 FILLER_10_228 ();
 sg13g2_fill_1 FILLER_10_239 ();
 sg13g2_decap_4 FILLER_10_258 ();
 sg13g2_fill_2 FILLER_10_262 ();
 sg13g2_fill_2 FILLER_10_274 ();
 sg13g2_decap_8 FILLER_10_285 ();
 sg13g2_fill_1 FILLER_10_292 ();
 sg13g2_decap_8 FILLER_10_314 ();
 sg13g2_fill_2 FILLER_10_321 ();
 sg13g2_fill_1 FILLER_10_323 ();
 sg13g2_decap_8 FILLER_10_328 ();
 sg13g2_decap_8 FILLER_10_335 ();
 sg13g2_decap_8 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_363 ();
 sg13g2_fill_1 FILLER_10_370 ();
 sg13g2_decap_8 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_4 FILLER_10_403 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_4 FILLER_11_154 ();
 sg13g2_fill_1 FILLER_11_158 ();
 sg13g2_fill_1 FILLER_11_163 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_4 FILLER_11_175 ();
 sg13g2_fill_1 FILLER_11_179 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_4 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_299 ();
 sg13g2_decap_4 FILLER_11_306 ();
 sg13g2_fill_2 FILLER_11_317 ();
 sg13g2_decap_8 FILLER_11_376 ();
 sg13g2_decap_8 FILLER_11_383 ();
 sg13g2_decap_8 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_4 FILLER_12_126 ();
 sg13g2_fill_1 FILLER_12_130 ();
 sg13g2_fill_1 FILLER_12_157 ();
 sg13g2_decap_4 FILLER_12_210 ();
 sg13g2_fill_2 FILLER_12_240 ();
 sg13g2_fill_1 FILLER_12_305 ();
 sg13g2_decap_4 FILLER_12_350 ();
 sg13g2_fill_1 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_366 ();
 sg13g2_decap_8 FILLER_12_373 ();
 sg13g2_decap_8 FILLER_12_380 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_fill_2 FILLER_13_126 ();
 sg13g2_fill_2 FILLER_13_173 ();
 sg13g2_fill_1 FILLER_13_190 ();
 sg13g2_fill_1 FILLER_13_232 ();
 sg13g2_fill_2 FILLER_13_269 ();
 sg13g2_fill_1 FILLER_13_296 ();
 sg13g2_decap_8 FILLER_13_339 ();
 sg13g2_decap_8 FILLER_13_346 ();
 sg13g2_decap_8 FILLER_13_353 ();
 sg13g2_decap_8 FILLER_13_360 ();
 sg13g2_decap_8 FILLER_13_367 ();
 sg13g2_decap_8 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_13_388 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_fill_2 FILLER_14_119 ();
 sg13g2_fill_1 FILLER_14_121 ();
 sg13g2_fill_1 FILLER_14_151 ();
 sg13g2_fill_2 FILLER_14_170 ();
 sg13g2_fill_1 FILLER_14_172 ();
 sg13g2_fill_2 FILLER_14_209 ();
 sg13g2_fill_1 FILLER_14_211 ();
 sg13g2_decap_8 FILLER_14_216 ();
 sg13g2_fill_1 FILLER_14_223 ();
 sg13g2_fill_1 FILLER_14_237 ();
 sg13g2_fill_1 FILLER_14_243 ();
 sg13g2_decap_8 FILLER_14_261 ();
 sg13g2_fill_1 FILLER_14_268 ();
 sg13g2_decap_4 FILLER_14_284 ();
 sg13g2_fill_1 FILLER_14_288 ();
 sg13g2_decap_8 FILLER_14_292 ();
 sg13g2_fill_2 FILLER_14_299 ();
 sg13g2_fill_1 FILLER_14_301 ();
 sg13g2_decap_4 FILLER_14_328 ();
 sg13g2_fill_1 FILLER_14_332 ();
 sg13g2_fill_1 FILLER_14_338 ();
 sg13g2_decap_8 FILLER_14_353 ();
 sg13g2_decap_8 FILLER_14_360 ();
 sg13g2_fill_2 FILLER_14_367 ();
 sg13g2_fill_1 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_fill_2 FILLER_15_126 ();
 sg13g2_fill_1 FILLER_15_128 ();
 sg13g2_decap_8 FILLER_15_146 ();
 sg13g2_decap_4 FILLER_15_153 ();
 sg13g2_fill_1 FILLER_15_157 ();
 sg13g2_decap_8 FILLER_15_166 ();
 sg13g2_decap_8 FILLER_15_173 ();
 sg13g2_fill_2 FILLER_15_180 ();
 sg13g2_fill_1 FILLER_15_182 ();
 sg13g2_decap_4 FILLER_15_196 ();
 sg13g2_fill_1 FILLER_15_200 ();
 sg13g2_decap_4 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_247 ();
 sg13g2_decap_8 FILLER_15_254 ();
 sg13g2_decap_8 FILLER_15_261 ();
 sg13g2_decap_8 FILLER_15_268 ();
 sg13g2_decap_8 FILLER_15_275 ();
 sg13g2_fill_2 FILLER_15_282 ();
 sg13g2_fill_2 FILLER_15_304 ();
 sg13g2_fill_1 FILLER_15_306 ();
 sg13g2_fill_1 FILLER_15_315 ();
 sg13g2_fill_1 FILLER_15_324 ();
 sg13g2_fill_1 FILLER_15_330 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_fill_1 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_146 ();
 sg13g2_fill_1 FILLER_16_153 ();
 sg13g2_decap_8 FILLER_16_198 ();
 sg13g2_decap_8 FILLER_16_205 ();
 sg13g2_decap_8 FILLER_16_212 ();
 sg13g2_decap_4 FILLER_16_219 ();
 sg13g2_fill_1 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_258 ();
 sg13g2_fill_2 FILLER_16_265 ();
 sg13g2_fill_1 FILLER_16_293 ();
 sg13g2_fill_2 FILLER_16_322 ();
 sg13g2_fill_1 FILLER_16_350 ();
 sg13g2_fill_2 FILLER_16_361 ();
 sg13g2_fill_1 FILLER_16_363 ();
 sg13g2_decap_4 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_4 FILLER_17_112 ();
 sg13g2_fill_2 FILLER_17_116 ();
 sg13g2_decap_8 FILLER_17_177 ();
 sg13g2_decap_8 FILLER_17_197 ();
 sg13g2_decap_8 FILLER_17_204 ();
 sg13g2_decap_8 FILLER_17_211 ();
 sg13g2_decap_8 FILLER_17_218 ();
 sg13g2_fill_1 FILLER_17_225 ();
 sg13g2_fill_2 FILLER_17_252 ();
 sg13g2_fill_1 FILLER_17_254 ();
 sg13g2_fill_1 FILLER_17_262 ();
 sg13g2_fill_1 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_352 ();
 sg13g2_fill_2 FILLER_17_359 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_fill_1 FILLER_18_152 ();
 sg13g2_fill_1 FILLER_18_163 ();
 sg13g2_fill_1 FILLER_18_169 ();
 sg13g2_fill_2 FILLER_18_178 ();
 sg13g2_fill_2 FILLER_18_189 ();
 sg13g2_fill_1 FILLER_18_191 ();
 sg13g2_fill_2 FILLER_18_254 ();
 sg13g2_decap_8 FILLER_18_262 ();
 sg13g2_decap_4 FILLER_18_269 ();
 sg13g2_fill_1 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_321 ();
 sg13g2_decap_8 FILLER_18_328 ();
 sg13g2_fill_2 FILLER_18_335 ();
 sg13g2_decap_8 FILLER_18_341 ();
 sg13g2_fill_2 FILLER_18_348 ();
 sg13g2_decap_8 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_128 ();
 sg13g2_fill_2 FILLER_19_149 ();
 sg13g2_fill_1 FILLER_19_151 ();
 sg13g2_fill_2 FILLER_19_194 ();
 sg13g2_fill_1 FILLER_19_196 ();
 sg13g2_decap_4 FILLER_19_233 ();
 sg13g2_fill_2 FILLER_19_247 ();
 sg13g2_decap_8 FILLER_19_254 ();
 sg13g2_fill_1 FILLER_19_261 ();
 sg13g2_fill_1 FILLER_19_267 ();
 sg13g2_fill_2 FILLER_19_276 ();
 sg13g2_fill_1 FILLER_19_278 ();
 sg13g2_fill_2 FILLER_19_306 ();
 sg13g2_decap_8 FILLER_19_316 ();
 sg13g2_fill_2 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_4 FILLER_20_126 ();
 sg13g2_fill_2 FILLER_20_130 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_fill_2 FILLER_20_147 ();
 sg13g2_fill_1 FILLER_20_149 ();
 sg13g2_decap_8 FILLER_20_166 ();
 sg13g2_decap_4 FILLER_20_173 ();
 sg13g2_fill_2 FILLER_20_177 ();
 sg13g2_decap_8 FILLER_20_199 ();
 sg13g2_decap_8 FILLER_20_206 ();
 sg13g2_decap_8 FILLER_20_213 ();
 sg13g2_decap_8 FILLER_20_220 ();
 sg13g2_fill_1 FILLER_20_227 ();
 sg13g2_decap_8 FILLER_20_282 ();
 sg13g2_fill_2 FILLER_20_289 ();
 sg13g2_decap_4 FILLER_20_296 ();
 sg13g2_fill_1 FILLER_20_300 ();
 sg13g2_fill_1 FILLER_20_320 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_decap_8 FILLER_20_354 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_decap_4 FILLER_20_368 ();
 sg13g2_fill_2 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_383 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_fill_1 FILLER_21_119 ();
 sg13g2_decap_4 FILLER_21_154 ();
 sg13g2_fill_2 FILLER_21_158 ();
 sg13g2_fill_1 FILLER_21_186 ();
 sg13g2_decap_4 FILLER_21_218 ();
 sg13g2_fill_2 FILLER_21_231 ();
 sg13g2_fill_2 FILLER_21_303 ();
 sg13g2_fill_1 FILLER_21_305 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_fill_2 FILLER_21_361 ();
 sg13g2_fill_2 FILLER_21_367 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_fill_2 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_173 ();
 sg13g2_decap_4 FILLER_22_180 ();
 sg13g2_fill_1 FILLER_22_184 ();
 sg13g2_decap_8 FILLER_22_197 ();
 sg13g2_decap_8 FILLER_22_204 ();
 sg13g2_decap_4 FILLER_22_211 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_4 FILLER_23_147 ();
 sg13g2_fill_1 FILLER_23_151 ();
 sg13g2_decap_8 FILLER_23_169 ();
 sg13g2_fill_1 FILLER_23_176 ();
 sg13g2_fill_2 FILLER_23_195 ();
 sg13g2_fill_1 FILLER_23_197 ();
 sg13g2_fill_1 FILLER_23_234 ();
 sg13g2_fill_2 FILLER_23_329 ();
 sg13g2_fill_1 FILLER_23_331 ();
 sg13g2_decap_8 FILLER_23_358 ();
 sg13g2_fill_2 FILLER_23_365 ();
 sg13g2_fill_1 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_fill_2 FILLER_24_126 ();
 sg13g2_fill_1 FILLER_24_184 ();
 sg13g2_decap_8 FILLER_24_211 ();
 sg13g2_decap_8 FILLER_24_218 ();
 sg13g2_decap_8 FILLER_24_225 ();
 sg13g2_fill_2 FILLER_24_232 ();
 sg13g2_fill_2 FILLER_24_243 ();
 sg13g2_decap_8 FILLER_24_254 ();
 sg13g2_decap_8 FILLER_24_261 ();
 sg13g2_decap_4 FILLER_24_268 ();
 sg13g2_fill_2 FILLER_24_272 ();
 sg13g2_fill_1 FILLER_24_277 ();
 sg13g2_decap_8 FILLER_24_282 ();
 sg13g2_fill_1 FILLER_24_289 ();
 sg13g2_fill_1 FILLER_24_299 ();
 sg13g2_fill_2 FILLER_24_319 ();
 sg13g2_decap_8 FILLER_24_330 ();
 sg13g2_decap_4 FILLER_24_337 ();
 sg13g2_fill_2 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_347 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_4 FILLER_25_119 ();
 sg13g2_fill_1 FILLER_25_123 ();
 sg13g2_decap_8 FILLER_25_145 ();
 sg13g2_fill_2 FILLER_25_152 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_fill_1 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_198 ();
 sg13g2_decap_4 FILLER_25_205 ();
 sg13g2_fill_1 FILLER_25_209 ();
 sg13g2_decap_8 FILLER_25_220 ();
 sg13g2_fill_2 FILLER_25_227 ();
 sg13g2_decap_8 FILLER_25_255 ();
 sg13g2_decap_8 FILLER_25_262 ();
 sg13g2_fill_1 FILLER_25_277 ();
 sg13g2_decap_8 FILLER_25_281 ();
 sg13g2_decap_8 FILLER_25_288 ();
 sg13g2_decap_8 FILLER_25_295 ();
 sg13g2_decap_8 FILLER_25_309 ();
 sg13g2_decap_4 FILLER_25_316 ();
 sg13g2_fill_1 FILLER_25_324 ();
 sg13g2_decap_4 FILLER_25_329 ();
 sg13g2_fill_1 FILLER_25_333 ();
 sg13g2_decap_4 FILLER_25_339 ();
 sg13g2_fill_2 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_353 ();
 sg13g2_decap_4 FILLER_25_360 ();
 sg13g2_fill_1 FILLER_25_364 ();
 sg13g2_fill_1 FILLER_25_369 ();
 sg13g2_decap_8 FILLER_25_376 ();
 sg13g2_decap_8 FILLER_25_383 ();
 sg13g2_decap_8 FILLER_25_390 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_4 FILLER_26_119 ();
 sg13g2_fill_2 FILLER_26_123 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_4 FILLER_26_175 ();
 sg13g2_fill_1 FILLER_26_179 ();
 sg13g2_decap_4 FILLER_26_240 ();
 sg13g2_fill_1 FILLER_26_244 ();
 sg13g2_fill_2 FILLER_26_299 ();
 sg13g2_fill_1 FILLER_26_301 ();
 sg13g2_fill_2 FILLER_26_324 ();
 sg13g2_fill_2 FILLER_26_331 ();
 sg13g2_fill_1 FILLER_26_333 ();
 sg13g2_fill_1 FILLER_26_370 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_119 ();
 sg13g2_fill_1 FILLER_27_121 ();
 sg13g2_decap_4 FILLER_27_148 ();
 sg13g2_fill_1 FILLER_27_186 ();
 sg13g2_decap_8 FILLER_27_199 ();
 sg13g2_decap_8 FILLER_27_206 ();
 sg13g2_decap_8 FILLER_27_213 ();
 sg13g2_decap_8 FILLER_27_220 ();
 sg13g2_decap_8 FILLER_27_227 ();
 sg13g2_decap_8 FILLER_27_234 ();
 sg13g2_decap_8 FILLER_27_241 ();
 sg13g2_decap_8 FILLER_27_248 ();
 sg13g2_fill_2 FILLER_27_312 ();
 sg13g2_fill_2 FILLER_27_322 ();
 sg13g2_fill_1 FILLER_27_324 ();
 sg13g2_decap_8 FILLER_27_351 ();
 sg13g2_fill_2 FILLER_27_358 ();
 sg13g2_fill_1 FILLER_27_360 ();
 sg13g2_fill_1 FILLER_27_366 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_4 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_fill_1 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_144 ();
 sg13g2_fill_1 FILLER_28_151 ();
 sg13g2_decap_8 FILLER_28_167 ();
 sg13g2_decap_8 FILLER_28_174 ();
 sg13g2_fill_2 FILLER_28_181 ();
 sg13g2_fill_1 FILLER_28_183 ();
 sg13g2_decap_4 FILLER_28_200 ();
 sg13g2_decap_8 FILLER_28_240 ();
 sg13g2_decap_8 FILLER_28_247 ();
 sg13g2_decap_8 FILLER_28_254 ();
 sg13g2_fill_1 FILLER_28_275 ();
 sg13g2_fill_2 FILLER_28_302 ();
 sg13g2_decap_8 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_4 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_123 ();
 sg13g2_fill_1 FILLER_29_146 ();
 sg13g2_fill_1 FILLER_29_150 ();
 sg13g2_fill_2 FILLER_29_218 ();
 sg13g2_fill_1 FILLER_29_220 ();
 sg13g2_decap_4 FILLER_29_226 ();
 sg13g2_fill_1 FILLER_29_256 ();
 sg13g2_fill_2 FILLER_29_262 ();
 sg13g2_fill_1 FILLER_29_264 ();
 sg13g2_fill_2 FILLER_29_279 ();
 sg13g2_decap_8 FILLER_29_369 ();
 sg13g2_decap_8 FILLER_29_376 ();
 sg13g2_decap_8 FILLER_29_383 ();
 sg13g2_decap_8 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_166 ();
 sg13g2_fill_1 FILLER_30_172 ();
 sg13g2_fill_2 FILLER_30_181 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_198 ();
 sg13g2_fill_1 FILLER_30_205 ();
 sg13g2_decap_8 FILLER_30_268 ();
 sg13g2_fill_1 FILLER_30_275 ();
 sg13g2_fill_1 FILLER_30_281 ();
 sg13g2_fill_2 FILLER_30_305 ();
 sg13g2_fill_2 FILLER_30_323 ();
 sg13g2_fill_1 FILLER_30_325 ();
 sg13g2_fill_2 FILLER_30_353 ();
 sg13g2_decap_4 FILLER_30_365 ();
 sg13g2_decap_4 FILLER_30_372 ();
 sg13g2_fill_1 FILLER_30_376 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_4 FILLER_31_119 ();
 sg13g2_fill_1 FILLER_31_123 ();
 sg13g2_decap_8 FILLER_31_166 ();
 sg13g2_decap_8 FILLER_31_173 ();
 sg13g2_decap_4 FILLER_31_180 ();
 sg13g2_fill_2 FILLER_31_184 ();
 sg13g2_decap_8 FILLER_31_220 ();
 sg13g2_fill_2 FILLER_31_227 ();
 sg13g2_fill_1 FILLER_31_229 ();
 sg13g2_decap_4 FILLER_31_280 ();
 sg13g2_fill_1 FILLER_31_284 ();
 sg13g2_fill_2 FILLER_31_301 ();
 sg13g2_fill_2 FILLER_31_307 ();
 sg13g2_fill_1 FILLER_31_309 ();
 sg13g2_decap_4 FILLER_31_323 ();
 sg13g2_fill_2 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_31_333 ();
 sg13g2_decap_8 FILLER_31_340 ();
 sg13g2_fill_2 FILLER_31_347 ();
 sg13g2_fill_1 FILLER_31_349 ();
 sg13g2_decap_8 FILLER_31_354 ();
 sg13g2_fill_1 FILLER_31_365 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_fill_2 FILLER_32_119 ();
 sg13g2_fill_1 FILLER_32_121 ();
 sg13g2_fill_2 FILLER_32_156 ();
 sg13g2_decap_8 FILLER_32_201 ();
 sg13g2_fill_2 FILLER_32_208 ();
 sg13g2_fill_1 FILLER_32_210 ();
 sg13g2_decap_4 FILLER_32_237 ();
 sg13g2_fill_1 FILLER_32_241 ();
 sg13g2_fill_2 FILLER_32_293 ();
 sg13g2_fill_1 FILLER_32_295 ();
 sg13g2_fill_1 FILLER_32_305 ();
 sg13g2_decap_8 FILLER_32_319 ();
 sg13g2_fill_2 FILLER_32_326 ();
 sg13g2_decap_8 FILLER_32_380 ();
 sg13g2_decap_8 FILLER_32_387 ();
 sg13g2_decap_8 FILLER_32_394 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_4 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_171 ();
 sg13g2_decap_8 FILLER_33_178 ();
 sg13g2_fill_2 FILLER_33_185 ();
 sg13g2_fill_2 FILLER_33_197 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_fill_1 FILLER_33_252 ();
 sg13g2_fill_1 FILLER_33_271 ();
 sg13g2_fill_2 FILLER_33_316 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_fill_2 FILLER_33_364 ();
 sg13g2_fill_1 FILLER_33_366 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_fill_2 FILLER_34_154 ();
 sg13g2_fill_1 FILLER_34_156 ();
 sg13g2_decap_8 FILLER_34_166 ();
 sg13g2_decap_4 FILLER_34_173 ();
 sg13g2_decap_4 FILLER_34_234 ();
 sg13g2_decap_8 FILLER_34_254 ();
 sg13g2_decap_4 FILLER_34_261 ();
 sg13g2_fill_1 FILLER_34_265 ();
 sg13g2_decap_4 FILLER_34_270 ();
 sg13g2_fill_1 FILLER_34_283 ();
 sg13g2_fill_2 FILLER_34_292 ();
 sg13g2_fill_1 FILLER_34_299 ();
 sg13g2_fill_2 FILLER_34_306 ();
 sg13g2_fill_2 FILLER_34_339 ();
 sg13g2_fill_1 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_fill_2 FILLER_35_133 ();
 sg13g2_decap_4 FILLER_35_143 ();
 sg13g2_fill_2 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_204 ();
 sg13g2_decap_8 FILLER_35_211 ();
 sg13g2_decap_4 FILLER_35_218 ();
 sg13g2_fill_2 FILLER_35_222 ();
 sg13g2_fill_1 FILLER_35_250 ();
 sg13g2_decap_8 FILLER_35_274 ();
 sg13g2_fill_1 FILLER_35_344 ();
 sg13g2_decap_8 FILLER_35_355 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_4 FILLER_36_119 ();
 sg13g2_fill_2 FILLER_36_123 ();
 sg13g2_decap_8 FILLER_36_172 ();
 sg13g2_decap_8 FILLER_36_179 ();
 sg13g2_fill_1 FILLER_36_186 ();
 sg13g2_decap_8 FILLER_36_195 ();
 sg13g2_decap_8 FILLER_36_202 ();
 sg13g2_decap_8 FILLER_36_209 ();
 sg13g2_decap_8 FILLER_36_216 ();
 sg13g2_fill_2 FILLER_36_223 ();
 sg13g2_fill_1 FILLER_36_251 ();
 sg13g2_decap_8 FILLER_36_282 ();
 sg13g2_fill_2 FILLER_36_289 ();
 sg13g2_fill_1 FILLER_36_296 ();
 sg13g2_decap_8 FILLER_36_326 ();
 sg13g2_fill_2 FILLER_36_333 ();
 sg13g2_fill_1 FILLER_36_343 ();
 sg13g2_decap_4 FILLER_36_354 ();
 sg13g2_fill_2 FILLER_36_358 ();
 sg13g2_decap_4 FILLER_36_364 ();
 sg13g2_decap_4 FILLER_36_371 ();
 sg13g2_fill_2 FILLER_36_375 ();
 sg13g2_decap_8 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_decap_8 FILLER_36_395 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_fill_1 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_166 ();
 sg13g2_decap_8 FILLER_37_173 ();
 sg13g2_decap_4 FILLER_37_180 ();
 sg13g2_decap_8 FILLER_37_192 ();
 sg13g2_decap_4 FILLER_37_199 ();
 sg13g2_fill_1 FILLER_37_203 ();
 sg13g2_decap_4 FILLER_37_230 ();
 sg13g2_fill_1 FILLER_37_258 ();
 sg13g2_decap_8 FILLER_37_283 ();
 sg13g2_decap_4 FILLER_37_290 ();
 sg13g2_fill_2 FILLER_37_294 ();
 sg13g2_fill_1 FILLER_37_300 ();
 sg13g2_fill_2 FILLER_37_304 ();
 sg13g2_fill_1 FILLER_37_306 ();
 sg13g2_fill_1 FILLER_37_316 ();
 sg13g2_fill_1 FILLER_37_348 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_4 FILLER_38_119 ();
 sg13g2_fill_2 FILLER_38_123 ();
 sg13g2_fill_2 FILLER_38_151 ();
 sg13g2_decap_8 FILLER_38_213 ();
 sg13g2_decap_8 FILLER_38_220 ();
 sg13g2_fill_2 FILLER_38_227 ();
 sg13g2_fill_2 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_253 ();
 sg13g2_fill_2 FILLER_38_265 ();
 sg13g2_decap_8 FILLER_38_272 ();
 sg13g2_decap_8 FILLER_38_279 ();
 sg13g2_decap_4 FILLER_38_286 ();
 sg13g2_fill_1 FILLER_38_290 ();
 sg13g2_fill_1 FILLER_38_296 ();
 sg13g2_decap_8 FILLER_38_310 ();
 sg13g2_decap_8 FILLER_38_317 ();
 sg13g2_decap_8 FILLER_38_324 ();
 sg13g2_fill_2 FILLER_38_331 ();
 sg13g2_decap_8 FILLER_38_337 ();
 sg13g2_fill_1 FILLER_38_344 ();
 sg13g2_decap_8 FILLER_38_349 ();
 sg13g2_decap_8 FILLER_38_356 ();
 sg13g2_decap_4 FILLER_38_363 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_fill_2 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_149 ();
 sg13g2_decap_4 FILLER_39_156 ();
 sg13g2_fill_1 FILLER_39_160 ();
 sg13g2_fill_2 FILLER_39_170 ();
 sg13g2_decap_4 FILLER_39_197 ();
 sg13g2_fill_1 FILLER_39_201 ();
 sg13g2_decap_4 FILLER_39_212 ();
 sg13g2_fill_2 FILLER_39_252 ();
 sg13g2_fill_1 FILLER_39_254 ();
 sg13g2_fill_2 FILLER_39_279 ();
 sg13g2_fill_1 FILLER_39_281 ();
 sg13g2_fill_2 FILLER_39_327 ();
 sg13g2_decap_8 FILLER_39_390 ();
 sg13g2_decap_8 FILLER_39_397 ();
 sg13g2_decap_4 FILLER_39_404 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_4 FILLER_40_126 ();
 sg13g2_decap_4 FILLER_40_151 ();
 sg13g2_fill_1 FILLER_40_155 ();
 sg13g2_fill_1 FILLER_40_173 ();
 sg13g2_decap_8 FILLER_40_200 ();
 sg13g2_decap_4 FILLER_40_207 ();
 sg13g2_fill_1 FILLER_40_275 ();
 sg13g2_fill_1 FILLER_40_306 ();
 sg13g2_fill_1 FILLER_40_338 ();
 sg13g2_decap_4 FILLER_40_362 ();
 sg13g2_decap_8 FILLER_40_370 ();
 sg13g2_decap_8 FILLER_40_377 ();
 sg13g2_decap_8 FILLER_40_384 ();
 sg13g2_decap_8 FILLER_40_391 ();
 sg13g2_decap_8 FILLER_40_398 ();
 sg13g2_decap_4 FILLER_40_405 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_4 FILLER_41_119 ();
 sg13g2_fill_2 FILLER_41_123 ();
 sg13g2_decap_4 FILLER_41_211 ();
 sg13g2_fill_2 FILLER_41_215 ();
 sg13g2_fill_1 FILLER_41_226 ();
 sg13g2_fill_1 FILLER_41_240 ();
 sg13g2_fill_2 FILLER_41_259 ();
 sg13g2_fill_1 FILLER_41_269 ();
 sg13g2_fill_2 FILLER_41_298 ();
 sg13g2_fill_1 FILLER_41_300 ();
 sg13g2_fill_2 FILLER_41_309 ();
 sg13g2_fill_1 FILLER_41_311 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_400 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_fill_2 FILLER_42_133 ();
 sg13g2_fill_1 FILLER_42_138 ();
 sg13g2_decap_4 FILLER_42_149 ();
 sg13g2_fill_2 FILLER_42_153 ();
 sg13g2_decap_8 FILLER_42_173 ();
 sg13g2_decap_4 FILLER_42_180 ();
 sg13g2_fill_2 FILLER_42_184 ();
 sg13g2_decap_4 FILLER_42_229 ();
 sg13g2_decap_8 FILLER_42_250 ();
 sg13g2_decap_4 FILLER_42_257 ();
 sg13g2_fill_2 FILLER_42_261 ();
 sg13g2_fill_2 FILLER_42_327 ();
 sg13g2_fill_1 FILLER_42_329 ();
 sg13g2_decap_4 FILLER_42_356 ();
 sg13g2_decap_8 FILLER_42_390 ();
 sg13g2_decap_8 FILLER_42_397 ();
 sg13g2_decap_4 FILLER_42_404 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_4 FILLER_43_126 ();
 sg13g2_fill_2 FILLER_43_130 ();
 sg13g2_decap_8 FILLER_43_148 ();
 sg13g2_decap_8 FILLER_43_155 ();
 sg13g2_decap_8 FILLER_43_162 ();
 sg13g2_decap_8 FILLER_43_169 ();
 sg13g2_decap_8 FILLER_43_176 ();
 sg13g2_decap_4 FILLER_43_183 ();
 sg13g2_decap_8 FILLER_43_192 ();
 sg13g2_fill_2 FILLER_43_199 ();
 sg13g2_fill_1 FILLER_43_201 ();
 sg13g2_decap_8 FILLER_43_220 ();
 sg13g2_decap_8 FILLER_43_227 ();
 sg13g2_decap_4 FILLER_43_234 ();
 sg13g2_fill_1 FILLER_43_238 ();
 sg13g2_fill_2 FILLER_43_260 ();
 sg13g2_decap_4 FILLER_43_267 ();
 sg13g2_fill_1 FILLER_43_271 ();
 sg13g2_decap_8 FILLER_43_381 ();
 sg13g2_decap_8 FILLER_43_388 ();
 sg13g2_decap_8 FILLER_43_395 ();
 sg13g2_decap_8 FILLER_43_402 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_fill_2 FILLER_44_133 ();
 sg13g2_fill_1 FILLER_44_161 ();
 sg13g2_fill_2 FILLER_44_175 ();
 sg13g2_decap_8 FILLER_44_211 ();
 sg13g2_fill_2 FILLER_44_218 ();
 sg13g2_fill_1 FILLER_44_220 ();
 sg13g2_fill_1 FILLER_44_257 ();
 sg13g2_fill_1 FILLER_44_271 ();
 sg13g2_decap_4 FILLER_44_283 ();
 sg13g2_fill_1 FILLER_44_287 ();
 sg13g2_fill_2 FILLER_44_296 ();
 sg13g2_fill_1 FILLER_44_298 ();
 sg13g2_fill_1 FILLER_44_303 ();
 sg13g2_decap_4 FILLER_44_334 ();
 sg13g2_fill_2 FILLER_44_338 ();
 sg13g2_fill_2 FILLER_44_345 ();
 sg13g2_fill_1 FILLER_44_347 ();
 sg13g2_decap_4 FILLER_44_357 ();
 sg13g2_fill_1 FILLER_44_361 ();
 sg13g2_decap_8 FILLER_44_366 ();
 sg13g2_decap_8 FILLER_44_373 ();
 sg13g2_decap_8 FILLER_44_380 ();
 sg13g2_decap_8 FILLER_44_387 ();
 sg13g2_decap_8 FILLER_44_394 ();
 sg13g2_decap_8 FILLER_44_401 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_fill_2 FILLER_45_154 ();
 sg13g2_fill_1 FILLER_45_156 ();
 sg13g2_fill_2 FILLER_45_293 ();
 sg13g2_fill_2 FILLER_45_313 ();
 sg13g2_decap_4 FILLER_45_327 ();
 sg13g2_decap_8 FILLER_45_372 ();
 sg13g2_decap_8 FILLER_45_383 ();
 sg13g2_decap_8 FILLER_45_390 ();
 sg13g2_decap_8 FILLER_45_397 ();
 sg13g2_decap_4 FILLER_45_404 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_4 FILLER_46_161 ();
 sg13g2_fill_2 FILLER_46_165 ();
 sg13g2_decap_8 FILLER_46_174 ();
 sg13g2_decap_8 FILLER_46_181 ();
 sg13g2_decap_8 FILLER_46_193 ();
 sg13g2_fill_2 FILLER_46_200 ();
 sg13g2_decap_4 FILLER_46_268 ();
 sg13g2_decap_4 FILLER_46_337 ();
 sg13g2_fill_2 FILLER_46_350 ();
 sg13g2_fill_1 FILLER_46_352 ();
 sg13g2_fill_2 FILLER_46_363 ();
 sg13g2_decap_8 FILLER_46_394 ();
 sg13g2_decap_8 FILLER_46_401 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_fill_2 FILLER_47_175 ();
 sg13g2_decap_4 FILLER_47_182 ();
 sg13g2_fill_1 FILLER_47_186 ();
 sg13g2_decap_8 FILLER_47_228 ();
 sg13g2_fill_2 FILLER_47_235 ();
 sg13g2_fill_1 FILLER_47_237 ();
 sg13g2_fill_1 FILLER_47_247 ();
 sg13g2_decap_8 FILLER_47_258 ();
 sg13g2_decap_4 FILLER_47_265 ();
 sg13g2_fill_2 FILLER_47_269 ();
 sg13g2_fill_1 FILLER_47_300 ();
 sg13g2_fill_2 FILLER_47_329 ();
 sg13g2_fill_1 FILLER_47_331 ();
 sg13g2_decap_8 FILLER_47_387 ();
 sg13g2_decap_8 FILLER_47_394 ();
 sg13g2_decap_8 FILLER_47_401 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_4 FILLER_48_126 ();
 sg13g2_fill_1 FILLER_48_130 ();
 sg13g2_decap_8 FILLER_48_157 ();
 sg13g2_decap_4 FILLER_48_164 ();
 sg13g2_decap_4 FILLER_48_173 ();
 sg13g2_fill_1 FILLER_48_177 ();
 sg13g2_decap_8 FILLER_48_212 ();
 sg13g2_decap_8 FILLER_48_219 ();
 sg13g2_decap_4 FILLER_48_226 ();
 sg13g2_fill_2 FILLER_48_230 ();
 sg13g2_decap_8 FILLER_48_236 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_4 FILLER_48_273 ();
 sg13g2_fill_1 FILLER_48_277 ();
 sg13g2_fill_2 FILLER_48_331 ();
 sg13g2_decap_8 FILLER_48_356 ();
 sg13g2_decap_8 FILLER_48_363 ();
 sg13g2_fill_2 FILLER_48_370 ();
 sg13g2_decap_8 FILLER_48_376 ();
 sg13g2_decap_8 FILLER_48_383 ();
 sg13g2_decap_8 FILLER_48_390 ();
 sg13g2_decap_8 FILLER_48_397 ();
 sg13g2_decap_4 FILLER_48_404 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_fill_1 FILLER_49_140 ();
 sg13g2_fill_2 FILLER_49_145 ();
 sg13g2_fill_1 FILLER_49_147 ();
 sg13g2_fill_2 FILLER_49_153 ();
 sg13g2_fill_1 FILLER_49_155 ();
 sg13g2_fill_2 FILLER_49_160 ();
 sg13g2_fill_1 FILLER_49_162 ();
 sg13g2_decap_8 FILLER_49_202 ();
 sg13g2_decap_8 FILLER_49_209 ();
 sg13g2_fill_2 FILLER_49_251 ();
 sg13g2_decap_8 FILLER_49_266 ();
 sg13g2_fill_2 FILLER_49_273 ();
 sg13g2_fill_1 FILLER_49_275 ();
 sg13g2_fill_2 FILLER_49_285 ();
 sg13g2_fill_1 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_331 ();
 sg13g2_decap_4 FILLER_49_338 ();
 sg13g2_decap_8 FILLER_49_368 ();
 sg13g2_decap_8 FILLER_49_375 ();
 sg13g2_decap_8 FILLER_49_382 ();
 sg13g2_decap_8 FILLER_49_389 ();
 sg13g2_decap_8 FILLER_49_396 ();
 sg13g2_decap_4 FILLER_49_403 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_8 FILLER_50_126 ();
 sg13g2_decap_8 FILLER_50_133 ();
 sg13g2_fill_2 FILLER_50_140 ();
 sg13g2_decap_4 FILLER_50_187 ();
 sg13g2_decap_4 FILLER_50_199 ();
 sg13g2_fill_1 FILLER_50_203 ();
 sg13g2_decap_4 FILLER_50_291 ();
 sg13g2_fill_1 FILLER_50_295 ();
 sg13g2_fill_2 FILLER_50_313 ();
 sg13g2_fill_1 FILLER_50_352 ();
 sg13g2_fill_1 FILLER_50_357 ();
 sg13g2_decap_8 FILLER_50_384 ();
 sg13g2_decap_8 FILLER_50_391 ();
 sg13g2_decap_8 FILLER_50_398 ();
 sg13g2_decap_4 FILLER_50_405 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_8 FILLER_51_119 ();
 sg13g2_decap_8 FILLER_51_126 ();
 sg13g2_decap_8 FILLER_51_133 ();
 sg13g2_decap_8 FILLER_51_140 ();
 sg13g2_decap_8 FILLER_51_147 ();
 sg13g2_decap_8 FILLER_51_154 ();
 sg13g2_decap_8 FILLER_51_161 ();
 sg13g2_decap_4 FILLER_51_168 ();
 sg13g2_fill_2 FILLER_51_172 ();
 sg13g2_fill_2 FILLER_51_182 ();
 sg13g2_fill_2 FILLER_51_201 ();
 sg13g2_fill_1 FILLER_51_203 ();
 sg13g2_fill_2 FILLER_51_253 ();
 sg13g2_fill_2 FILLER_51_299 ();
 sg13g2_fill_2 FILLER_51_353 ();
 sg13g2_fill_2 FILLER_51_365 ();
 sg13g2_fill_1 FILLER_51_367 ();
 sg13g2_decap_8 FILLER_51_398 ();
 sg13g2_decap_4 FILLER_51_405 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_119 ();
 sg13g2_decap_8 FILLER_52_126 ();
 sg13g2_decap_8 FILLER_52_133 ();
 sg13g2_decap_8 FILLER_52_140 ();
 sg13g2_decap_8 FILLER_52_147 ();
 sg13g2_decap_8 FILLER_52_154 ();
 sg13g2_decap_8 FILLER_52_161 ();
 sg13g2_decap_8 FILLER_52_168 ();
 sg13g2_fill_2 FILLER_52_175 ();
 sg13g2_fill_1 FILLER_52_189 ();
 sg13g2_decap_8 FILLER_52_216 ();
 sg13g2_decap_8 FILLER_52_223 ();
 sg13g2_decap_4 FILLER_52_230 ();
 sg13g2_decap_4 FILLER_52_238 ();
 sg13g2_fill_2 FILLER_52_242 ();
 sg13g2_fill_1 FILLER_52_249 ();
 sg13g2_decap_8 FILLER_52_254 ();
 sg13g2_decap_4 FILLER_52_261 ();
 sg13g2_decap_4 FILLER_52_294 ();
 sg13g2_decap_8 FILLER_52_365 ();
 sg13g2_fill_2 FILLER_52_372 ();
 sg13g2_decap_4 FILLER_52_377 ();
 sg13g2_fill_2 FILLER_52_381 ();
 sg13g2_decap_8 FILLER_52_387 ();
 sg13g2_decap_8 FILLER_52_394 ();
 sg13g2_decap_8 FILLER_52_401 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_decap_8 FILLER_53_133 ();
 sg13g2_decap_8 FILLER_53_140 ();
 sg13g2_decap_8 FILLER_53_147 ();
 sg13g2_decap_8 FILLER_53_154 ();
 sg13g2_decap_4 FILLER_53_161 ();
 sg13g2_fill_2 FILLER_53_165 ();
 sg13g2_decap_8 FILLER_53_210 ();
 sg13g2_decap_8 FILLER_53_217 ();
 sg13g2_decap_8 FILLER_53_224 ();
 sg13g2_decap_8 FILLER_53_231 ();
 sg13g2_decap_8 FILLER_53_238 ();
 sg13g2_decap_8 FILLER_53_245 ();
 sg13g2_decap_8 FILLER_53_252 ();
 sg13g2_decap_8 FILLER_53_259 ();
 sg13g2_fill_2 FILLER_53_266 ();
 sg13g2_fill_1 FILLER_53_268 ();
 sg13g2_decap_8 FILLER_53_285 ();
 sg13g2_decap_8 FILLER_53_292 ();
 sg13g2_fill_1 FILLER_53_299 ();
 sg13g2_fill_1 FILLER_53_304 ();
 sg13g2_fill_2 FILLER_53_324 ();
 sg13g2_decap_8 FILLER_53_330 ();
 sg13g2_fill_2 FILLER_53_337 ();
 sg13g2_decap_4 FILLER_53_344 ();
 sg13g2_decap_8 FILLER_53_356 ();
 sg13g2_decap_4 FILLER_53_363 ();
 sg13g2_fill_2 FILLER_53_367 ();
 sg13g2_decap_8 FILLER_53_373 ();
 sg13g2_decap_8 FILLER_53_380 ();
 sg13g2_decap_8 FILLER_53_387 ();
 sg13g2_decap_8 FILLER_53_394 ();
 sg13g2_decap_8 FILLER_53_401 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_decap_8 FILLER_54_119 ();
 sg13g2_decap_8 FILLER_54_126 ();
 sg13g2_decap_4 FILLER_54_171 ();
 sg13g2_decap_8 FILLER_54_187 ();
 sg13g2_decap_8 FILLER_54_194 ();
 sg13g2_decap_8 FILLER_54_201 ();
 sg13g2_decap_8 FILLER_54_208 ();
 sg13g2_decap_8 FILLER_54_215 ();
 sg13g2_decap_8 FILLER_54_222 ();
 sg13g2_decap_4 FILLER_54_229 ();
 sg13g2_fill_2 FILLER_54_259 ();
 sg13g2_fill_1 FILLER_54_334 ();
 sg13g2_fill_1 FILLER_54_339 ();
 sg13g2_decap_8 FILLER_54_350 ();
 sg13g2_fill_1 FILLER_54_357 ();
 sg13g2_decap_8 FILLER_54_388 ();
 sg13g2_decap_8 FILLER_54_395 ();
 sg13g2_decap_8 FILLER_54_402 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_decap_8 FILLER_55_126 ();
 sg13g2_decap_8 FILLER_55_133 ();
 sg13g2_decap_4 FILLER_55_140 ();
 sg13g2_decap_8 FILLER_55_174 ();
 sg13g2_decap_8 FILLER_55_181 ();
 sg13g2_decap_8 FILLER_55_188 ();
 sg13g2_fill_2 FILLER_55_195 ();
 sg13g2_decap_8 FILLER_55_201 ();
 sg13g2_fill_2 FILLER_55_208 ();
 sg13g2_fill_2 FILLER_55_322 ();
 sg13g2_fill_2 FILLER_55_350 ();
 sg13g2_fill_1 FILLER_55_352 ();
 sg13g2_decap_4 FILLER_55_357 ();
 sg13g2_decap_4 FILLER_55_364 ();
 sg13g2_fill_2 FILLER_55_368 ();
 sg13g2_decap_8 FILLER_55_399 ();
 sg13g2_fill_2 FILLER_55_406 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_decap_8 FILLER_56_119 ();
 sg13g2_decap_8 FILLER_56_126 ();
 sg13g2_fill_2 FILLER_56_133 ();
 sg13g2_fill_1 FILLER_56_135 ();
 sg13g2_decap_8 FILLER_56_140 ();
 sg13g2_fill_2 FILLER_56_147 ();
 sg13g2_fill_1 FILLER_56_149 ();
 sg13g2_decap_4 FILLER_56_153 ();
 sg13g2_fill_2 FILLER_56_157 ();
 sg13g2_fill_2 FILLER_56_170 ();
 sg13g2_fill_1 FILLER_56_172 ();
 sg13g2_decap_8 FILLER_56_185 ();
 sg13g2_fill_2 FILLER_56_192 ();
 sg13g2_fill_1 FILLER_56_220 ();
 sg13g2_fill_1 FILLER_56_286 ();
 sg13g2_fill_2 FILLER_56_339 ();
 sg13g2_fill_1 FILLER_56_341 ();
 sg13g2_decap_8 FILLER_56_373 ();
 sg13g2_decap_8 FILLER_56_380 ();
 sg13g2_decap_8 FILLER_56_387 ();
 sg13g2_decap_8 FILLER_56_394 ();
 sg13g2_decap_8 FILLER_56_401 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_4 FILLER_57_119 ();
 sg13g2_fill_2 FILLER_57_123 ();
 sg13g2_decap_4 FILLER_57_151 ();
 sg13g2_fill_1 FILLER_57_155 ();
 sg13g2_fill_2 FILLER_57_163 ();
 sg13g2_fill_2 FILLER_57_207 ();
 sg13g2_fill_2 FILLER_57_219 ();
 sg13g2_decap_4 FILLER_57_271 ();
 sg13g2_fill_1 FILLER_57_275 ();
 sg13g2_decap_8 FILLER_57_281 ();
 sg13g2_decap_8 FILLER_57_288 ();
 sg13g2_fill_2 FILLER_57_295 ();
 sg13g2_fill_2 FILLER_57_331 ();
 sg13g2_fill_1 FILLER_57_333 ();
 sg13g2_decap_8 FILLER_57_386 ();
 sg13g2_decap_8 FILLER_57_393 ();
 sg13g2_decap_8 FILLER_57_400 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_4 FILLER_58_133 ();
 sg13g2_fill_2 FILLER_58_137 ();
 sg13g2_fill_2 FILLER_58_168 ();
 sg13g2_decap_4 FILLER_58_191 ();
 sg13g2_decap_8 FILLER_58_221 ();
 sg13g2_decap_8 FILLER_58_228 ();
 sg13g2_decap_8 FILLER_58_235 ();
 sg13g2_fill_2 FILLER_58_242 ();
 sg13g2_decap_8 FILLER_58_255 ();
 sg13g2_decap_8 FILLER_58_262 ();
 sg13g2_decap_8 FILLER_58_269 ();
 sg13g2_fill_2 FILLER_58_276 ();
 sg13g2_decap_8 FILLER_58_282 ();
 sg13g2_decap_8 FILLER_58_289 ();
 sg13g2_decap_4 FILLER_58_296 ();
 sg13g2_fill_2 FILLER_58_319 ();
 sg13g2_decap_4 FILLER_58_331 ();
 sg13g2_decap_8 FILLER_58_384 ();
 sg13g2_decap_8 FILLER_58_391 ();
 sg13g2_decap_8 FILLER_58_398 ();
 sg13g2_decap_4 FILLER_58_405 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_8 FILLER_59_126 ();
 sg13g2_fill_1 FILLER_59_133 ();
 sg13g2_decap_8 FILLER_59_138 ();
 sg13g2_decap_8 FILLER_59_145 ();
 sg13g2_fill_1 FILLER_59_152 ();
 sg13g2_decap_8 FILLER_59_157 ();
 sg13g2_decap_4 FILLER_59_164 ();
 sg13g2_fill_2 FILLER_59_202 ();
 sg13g2_fill_1 FILLER_59_204 ();
 sg13g2_decap_8 FILLER_59_241 ();
 sg13g2_fill_2 FILLER_59_248 ();
 sg13g2_fill_1 FILLER_59_250 ();
 sg13g2_fill_1 FILLER_59_292 ();
 sg13g2_decap_4 FILLER_59_308 ();
 sg13g2_decap_4 FILLER_59_317 ();
 sg13g2_fill_2 FILLER_59_321 ();
 sg13g2_decap_8 FILLER_59_327 ();
 sg13g2_decap_8 FILLER_59_334 ();
 sg13g2_decap_4 FILLER_59_341 ();
 sg13g2_decap_8 FILLER_59_353 ();
 sg13g2_decap_4 FILLER_59_360 ();
 sg13g2_fill_1 FILLER_59_364 ();
 sg13g2_fill_2 FILLER_59_373 ();
 sg13g2_decap_8 FILLER_59_401 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_112 ();
 sg13g2_decap_4 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_153 ();
 sg13g2_decap_8 FILLER_60_160 ();
 sg13g2_decap_8 FILLER_60_167 ();
 sg13g2_decap_8 FILLER_60_179 ();
 sg13g2_decap_8 FILLER_60_186 ();
 sg13g2_fill_2 FILLER_60_214 ();
 sg13g2_fill_1 FILLER_60_262 ();
 sg13g2_fill_1 FILLER_60_284 ();
 sg13g2_decap_8 FILLER_60_347 ();
 sg13g2_decap_8 FILLER_60_354 ();
 sg13g2_decap_8 FILLER_60_361 ();
 sg13g2_decap_8 FILLER_60_368 ();
 sg13g2_fill_1 FILLER_60_375 ();
 sg13g2_decap_8 FILLER_60_379 ();
 sg13g2_decap_8 FILLER_60_390 ();
 sg13g2_decap_8 FILLER_60_397 ();
 sg13g2_decap_4 FILLER_60_404 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_decap_8 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_126 ();
 sg13g2_fill_2 FILLER_61_179 ();
 sg13g2_fill_1 FILLER_61_181 ();
 sg13g2_fill_1 FILLER_61_186 ();
 sg13g2_decap_8 FILLER_61_191 ();
 sg13g2_decap_4 FILLER_61_198 ();
 sg13g2_fill_1 FILLER_61_202 ();
 sg13g2_fill_1 FILLER_61_229 ();
 sg13g2_fill_2 FILLER_61_342 ();
 sg13g2_fill_1 FILLER_61_344 ();
 sg13g2_decap_8 FILLER_61_348 ();
 sg13g2_fill_2 FILLER_61_355 ();
 sg13g2_fill_1 FILLER_61_357 ();
 sg13g2_decap_8 FILLER_61_384 ();
 sg13g2_decap_8 FILLER_61_391 ();
 sg13g2_decap_8 FILLER_61_398 ();
 sg13g2_decap_4 FILLER_61_405 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_decap_8 FILLER_62_126 ();
 sg13g2_decap_8 FILLER_62_133 ();
 sg13g2_decap_4 FILLER_62_140 ();
 sg13g2_fill_2 FILLER_62_187 ();
 sg13g2_fill_1 FILLER_62_189 ();
 sg13g2_fill_2 FILLER_62_203 ();
 sg13g2_decap_4 FILLER_62_224 ();
 sg13g2_decap_4 FILLER_62_241 ();
 sg13g2_fill_2 FILLER_62_245 ();
 sg13g2_fill_2 FILLER_62_273 ();
 sg13g2_fill_1 FILLER_62_275 ();
 sg13g2_decap_8 FILLER_62_286 ();
 sg13g2_decap_4 FILLER_62_293 ();
 sg13g2_fill_2 FILLER_62_297 ();
 sg13g2_decap_4 FILLER_62_307 ();
 sg13g2_fill_1 FILLER_62_315 ();
 sg13g2_decap_8 FILLER_62_397 ();
 sg13g2_decap_4 FILLER_62_404 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_8 FILLER_63_126 ();
 sg13g2_decap_8 FILLER_63_133 ();
 sg13g2_fill_2 FILLER_63_140 ();
 sg13g2_fill_1 FILLER_63_142 ();
 sg13g2_fill_1 FILLER_63_177 ();
 sg13g2_decap_4 FILLER_63_209 ();
 sg13g2_decap_8 FILLER_63_230 ();
 sg13g2_decap_8 FILLER_63_237 ();
 sg13g2_decap_8 FILLER_63_244 ();
 sg13g2_decap_8 FILLER_63_251 ();
 sg13g2_decap_8 FILLER_63_258 ();
 sg13g2_decap_8 FILLER_63_265 ();
 sg13g2_decap_8 FILLER_63_272 ();
 sg13g2_decap_8 FILLER_63_279 ();
 sg13g2_fill_1 FILLER_63_286 ();
 sg13g2_decap_8 FILLER_63_291 ();
 sg13g2_decap_8 FILLER_63_298 ();
 sg13g2_decap_8 FILLER_63_305 ();
 sg13g2_decap_8 FILLER_63_312 ();
 sg13g2_decap_8 FILLER_63_319 ();
 sg13g2_decap_8 FILLER_63_326 ();
 sg13g2_decap_8 FILLER_63_359 ();
 sg13g2_decap_8 FILLER_63_366 ();
 sg13g2_decap_8 FILLER_63_373 ();
 sg13g2_decap_8 FILLER_63_380 ();
 sg13g2_decap_8 FILLER_63_387 ();
 sg13g2_decap_8 FILLER_63_394 ();
 sg13g2_decap_8 FILLER_63_401 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_fill_2 FILLER_64_147 ();
 sg13g2_fill_1 FILLER_64_149 ();
 sg13g2_decap_8 FILLER_64_237 ();
 sg13g2_decap_8 FILLER_64_244 ();
 sg13g2_fill_1 FILLER_64_251 ();
 sg13g2_decap_8 FILLER_64_265 ();
 sg13g2_decap_8 FILLER_64_272 ();
 sg13g2_fill_1 FILLER_64_279 ();
 sg13g2_decap_8 FILLER_64_299 ();
 sg13g2_decap_8 FILLER_64_306 ();
 sg13g2_decap_8 FILLER_64_313 ();
 sg13g2_decap_4 FILLER_64_320 ();
 sg13g2_fill_1 FILLER_64_324 ();
 sg13g2_decap_8 FILLER_64_356 ();
 sg13g2_decap_8 FILLER_64_363 ();
 sg13g2_decap_8 FILLER_64_370 ();
 sg13g2_fill_2 FILLER_64_377 ();
 sg13g2_fill_1 FILLER_64_379 ();
 sg13g2_decap_8 FILLER_64_392 ();
 sg13g2_decap_8 FILLER_64_399 ();
 sg13g2_fill_2 FILLER_64_406 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_decap_8 FILLER_65_140 ();
 sg13g2_decap_8 FILLER_65_147 ();
 sg13g2_decap_4 FILLER_65_154 ();
 sg13g2_fill_2 FILLER_65_158 ();
 sg13g2_fill_2 FILLER_65_168 ();
 sg13g2_fill_1 FILLER_65_170 ();
 sg13g2_decap_8 FILLER_65_210 ();
 sg13g2_fill_2 FILLER_65_230 ();
 sg13g2_decap_4 FILLER_65_271 ();
 sg13g2_fill_2 FILLER_65_301 ();
 sg13g2_fill_1 FILLER_65_303 ();
 sg13g2_decap_8 FILLER_65_324 ();
 sg13g2_fill_2 FILLER_65_334 ();
 sg13g2_fill_1 FILLER_65_341 ();
 sg13g2_decap_8 FILLER_65_368 ();
 sg13g2_fill_2 FILLER_65_375 ();
 sg13g2_fill_1 FILLER_65_377 ();
 sg13g2_decap_8 FILLER_65_386 ();
 sg13g2_decap_8 FILLER_65_393 ();
 sg13g2_decap_8 FILLER_65_400 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_126 ();
 sg13g2_decap_8 FILLER_66_133 ();
 sg13g2_decap_8 FILLER_66_140 ();
 sg13g2_fill_2 FILLER_66_147 ();
 sg13g2_fill_1 FILLER_66_149 ();
 sg13g2_decap_8 FILLER_66_154 ();
 sg13g2_decap_8 FILLER_66_161 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_fill_2 FILLER_66_175 ();
 sg13g2_fill_1 FILLER_66_177 ();
 sg13g2_decap_8 FILLER_66_208 ();
 sg13g2_fill_2 FILLER_66_215 ();
 sg13g2_decap_4 FILLER_66_233 ();
 sg13g2_fill_1 FILLER_66_237 ();
 sg13g2_fill_1 FILLER_66_251 ();
 sg13g2_decap_8 FILLER_66_334 ();
 sg13g2_decap_8 FILLER_66_341 ();
 sg13g2_decap_4 FILLER_66_348 ();
 sg13g2_fill_1 FILLER_66_352 ();
 sg13g2_decap_8 FILLER_66_392 ();
 sg13g2_decap_8 FILLER_66_399 ();
 sg13g2_fill_2 FILLER_66_406 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_4 FILLER_67_133 ();
 sg13g2_fill_2 FILLER_67_137 ();
 sg13g2_decap_8 FILLER_67_169 ();
 sg13g2_decap_8 FILLER_67_176 ();
 sg13g2_fill_2 FILLER_67_183 ();
 sg13g2_fill_1 FILLER_67_185 ();
 sg13g2_decap_8 FILLER_67_191 ();
 sg13g2_decap_4 FILLER_67_198 ();
 sg13g2_fill_1 FILLER_67_202 ();
 sg13g2_fill_2 FILLER_67_229 ();
 sg13g2_fill_2 FILLER_67_249 ();
 sg13g2_fill_1 FILLER_67_251 ();
 sg13g2_decap_8 FILLER_67_260 ();
 sg13g2_fill_1 FILLER_67_284 ();
 sg13g2_fill_1 FILLER_67_320 ();
 sg13g2_fill_2 FILLER_67_351 ();
 sg13g2_fill_2 FILLER_67_361 ();
 sg13g2_decap_8 FILLER_67_397 ();
 sg13g2_decap_4 FILLER_67_404 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_decap_8 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_decap_4 FILLER_68_147 ();
 sg13g2_decap_8 FILLER_68_180 ();
 sg13g2_decap_8 FILLER_68_187 ();
 sg13g2_decap_8 FILLER_68_194 ();
 sg13g2_decap_8 FILLER_68_201 ();
 sg13g2_decap_4 FILLER_68_208 ();
 sg13g2_fill_1 FILLER_68_225 ();
 sg13g2_fill_1 FILLER_68_252 ();
 sg13g2_decap_4 FILLER_68_270 ();
 sg13g2_fill_2 FILLER_68_282 ();
 sg13g2_fill_2 FILLER_68_314 ();
 sg13g2_fill_2 FILLER_68_360 ();
 sg13g2_decap_8 FILLER_68_389 ();
 sg13g2_decap_8 FILLER_68_396 ();
 sg13g2_decap_4 FILLER_68_403 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_fill_2 FILLER_69_126 ();
 sg13g2_fill_1 FILLER_69_128 ();
 sg13g2_decap_8 FILLER_69_155 ();
 sg13g2_fill_2 FILLER_69_162 ();
 sg13g2_fill_1 FILLER_69_164 ();
 sg13g2_decap_8 FILLER_69_172 ();
 sg13g2_decap_4 FILLER_69_179 ();
 sg13g2_fill_2 FILLER_69_183 ();
 sg13g2_decap_4 FILLER_69_188 ();
 sg13g2_fill_1 FILLER_69_192 ();
 sg13g2_decap_8 FILLER_69_201 ();
 sg13g2_decap_8 FILLER_69_208 ();
 sg13g2_decap_8 FILLER_69_215 ();
 sg13g2_fill_1 FILLER_69_222 ();
 sg13g2_fill_1 FILLER_69_252 ();
 sg13g2_decap_8 FILLER_69_279 ();
 sg13g2_decap_8 FILLER_69_286 ();
 sg13g2_fill_1 FILLER_69_293 ();
 sg13g2_fill_2 FILLER_69_301 ();
 sg13g2_fill_1 FILLER_69_303 ();
 sg13g2_fill_1 FILLER_69_308 ();
 sg13g2_decap_4 FILLER_69_313 ();
 sg13g2_fill_2 FILLER_69_317 ();
 sg13g2_fill_1 FILLER_69_329 ();
 sg13g2_decap_8 FILLER_69_385 ();
 sg13g2_decap_8 FILLER_69_392 ();
 sg13g2_decap_8 FILLER_69_399 ();
 sg13g2_fill_2 FILLER_69_406 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_4 FILLER_70_133 ();
 sg13g2_fill_2 FILLER_70_137 ();
 sg13g2_decap_4 FILLER_70_169 ();
 sg13g2_fill_2 FILLER_70_173 ();
 sg13g2_decap_8 FILLER_70_215 ();
 sg13g2_fill_2 FILLER_70_222 ();
 sg13g2_fill_1 FILLER_70_239 ();
 sg13g2_decap_8 FILLER_70_266 ();
 sg13g2_decap_4 FILLER_70_273 ();
 sg13g2_fill_1 FILLER_70_277 ();
 sg13g2_fill_2 FILLER_70_290 ();
 sg13g2_decap_4 FILLER_70_331 ();
 sg13g2_fill_1 FILLER_70_335 ();
 sg13g2_fill_2 FILLER_70_352 ();
 sg13g2_fill_1 FILLER_70_384 ();
 sg13g2_decap_8 FILLER_70_389 ();
 sg13g2_decap_8 FILLER_70_396 ();
 sg13g2_decap_4 FILLER_70_403 ();
 sg13g2_fill_2 FILLER_70_407 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_4 FILLER_71_140 ();
 sg13g2_fill_1 FILLER_71_144 ();
 sg13g2_decap_4 FILLER_71_148 ();
 sg13g2_fill_1 FILLER_71_152 ();
 sg13g2_decap_8 FILLER_71_252 ();
 sg13g2_decap_8 FILLER_71_259 ();
 sg13g2_decap_8 FILLER_71_266 ();
 sg13g2_decap_8 FILLER_71_273 ();
 sg13g2_decap_8 FILLER_71_280 ();
 sg13g2_decap_8 FILLER_71_287 ();
 sg13g2_decap_8 FILLER_71_294 ();
 sg13g2_fill_2 FILLER_71_301 ();
 sg13g2_decap_8 FILLER_71_336 ();
 sg13g2_fill_1 FILLER_71_343 ();
 sg13g2_fill_1 FILLER_71_375 ();
 sg13g2_decap_8 FILLER_71_395 ();
 sg13g2_decap_8 FILLER_71_402 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_4 FILLER_72_147 ();
 sg13g2_fill_2 FILLER_72_151 ();
 sg13g2_fill_1 FILLER_72_209 ();
 sg13g2_decap_8 FILLER_72_221 ();
 sg13g2_decap_8 FILLER_72_228 ();
 sg13g2_decap_4 FILLER_72_235 ();
 sg13g2_decap_8 FILLER_72_247 ();
 sg13g2_decap_8 FILLER_72_254 ();
 sg13g2_decap_4 FILLER_72_261 ();
 sg13g2_fill_1 FILLER_72_329 ();
 sg13g2_fill_2 FILLER_72_367 ();
 sg13g2_fill_2 FILLER_72_407 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_4 FILLER_73_140 ();
 sg13g2_fill_2 FILLER_73_144 ();
 sg13g2_fill_1 FILLER_73_172 ();
 sg13g2_decap_8 FILLER_73_177 ();
 sg13g2_decap_8 FILLER_73_184 ();
 sg13g2_decap_8 FILLER_73_191 ();
 sg13g2_decap_8 FILLER_73_198 ();
 sg13g2_decap_8 FILLER_73_231 ();
 sg13g2_decap_8 FILLER_73_238 ();
 sg13g2_decap_8 FILLER_73_245 ();
 sg13g2_fill_2 FILLER_73_252 ();
 sg13g2_decap_8 FILLER_73_283 ();
 sg13g2_decap_8 FILLER_73_290 ();
 sg13g2_decap_4 FILLER_73_297 ();
 sg13g2_fill_2 FILLER_73_301 ();
 sg13g2_fill_1 FILLER_73_315 ();
 sg13g2_fill_1 FILLER_73_341 ();
 sg13g2_decap_8 FILLER_73_402 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_168 ();
 sg13g2_decap_8 FILLER_74_175 ();
 sg13g2_decap_8 FILLER_74_182 ();
 sg13g2_decap_8 FILLER_74_189 ();
 sg13g2_decap_8 FILLER_74_196 ();
 sg13g2_decap_8 FILLER_74_203 ();
 sg13g2_decap_4 FILLER_74_210 ();
 sg13g2_fill_2 FILLER_74_214 ();
 sg13g2_fill_2 FILLER_74_220 ();
 sg13g2_decap_8 FILLER_74_248 ();
 sg13g2_decap_8 FILLER_74_307 ();
 sg13g2_fill_1 FILLER_74_314 ();
 sg13g2_decap_8 FILLER_74_338 ();
 sg13g2_fill_2 FILLER_74_345 ();
 sg13g2_decap_8 FILLER_74_376 ();
 sg13g2_decap_8 FILLER_74_383 ();
 sg13g2_decap_8 FILLER_74_390 ();
 sg13g2_decap_8 FILLER_74_397 ();
 sg13g2_decap_4 FILLER_74_404 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_8 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_182 ();
 sg13g2_decap_8 FILLER_75_189 ();
 sg13g2_decap_8 FILLER_75_196 ();
 sg13g2_decap_8 FILLER_75_203 ();
 sg13g2_decap_8 FILLER_75_210 ();
 sg13g2_decap_8 FILLER_75_217 ();
 sg13g2_decap_4 FILLER_75_227 ();
 sg13g2_fill_2 FILLER_75_231 ();
 sg13g2_decap_8 FILLER_75_237 ();
 sg13g2_decap_8 FILLER_75_244 ();
 sg13g2_decap_8 FILLER_75_251 ();
 sg13g2_decap_8 FILLER_75_258 ();
 sg13g2_decap_8 FILLER_75_265 ();
 sg13g2_decap_8 FILLER_75_272 ();
 sg13g2_decap_8 FILLER_75_279 ();
 sg13g2_decap_8 FILLER_75_286 ();
 sg13g2_fill_2 FILLER_75_293 ();
 sg13g2_decap_4 FILLER_75_321 ();
 sg13g2_decap_8 FILLER_75_333 ();
 sg13g2_decap_8 FILLER_75_340 ();
 sg13g2_decap_8 FILLER_75_347 ();
 sg13g2_decap_8 FILLER_75_354 ();
 sg13g2_decap_8 FILLER_75_361 ();
 sg13g2_decap_8 FILLER_75_368 ();
 sg13g2_decap_8 FILLER_75_375 ();
 sg13g2_decap_8 FILLER_75_382 ();
 sg13g2_decap_8 FILLER_75_389 ();
 sg13g2_decap_8 FILLER_75_396 ();
 sg13g2_decap_4 FILLER_75_403 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_8 FILLER_76_189 ();
 sg13g2_decap_8 FILLER_76_196 ();
 sg13g2_decap_8 FILLER_76_203 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_decap_8 FILLER_76_217 ();
 sg13g2_decap_8 FILLER_76_224 ();
 sg13g2_decap_4 FILLER_76_231 ();
 sg13g2_decap_8 FILLER_76_240 ();
 sg13g2_decap_4 FILLER_76_247 ();
 sg13g2_fill_1 FILLER_76_251 ();
 sg13g2_decap_4 FILLER_76_257 ();
 sg13g2_fill_1 FILLER_76_261 ();
 sg13g2_fill_1 FILLER_76_314 ();
 sg13g2_decap_4 FILLER_76_324 ();
 sg13g2_fill_1 FILLER_76_335 ();
 sg13g2_decap_4 FILLER_76_340 ();
 sg13g2_decap_8 FILLER_76_348 ();
 sg13g2_decap_8 FILLER_76_355 ();
 sg13g2_decap_4 FILLER_76_362 ();
 sg13g2_decap_8 FILLER_76_375 ();
 sg13g2_decap_8 FILLER_76_382 ();
 sg13g2_decap_8 FILLER_76_389 ();
 sg13g2_decap_8 FILLER_76_396 ();
 sg13g2_decap_4 FILLER_76_403 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_8 FILLER_77_217 ();
 sg13g2_fill_1 FILLER_77_224 ();
 sg13g2_decap_8 FILLER_77_283 ();
 sg13g2_decap_8 FILLER_77_290 ();
 sg13g2_decap_8 FILLER_77_297 ();
 sg13g2_decap_8 FILLER_77_381 ();
 sg13g2_decap_8 FILLER_77_388 ();
 sg13g2_decap_8 FILLER_77_395 ();
 sg13g2_decap_8 FILLER_77_402 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_203 ();
 sg13g2_decap_8 FILLER_78_210 ();
 sg13g2_decap_8 FILLER_78_217 ();
 sg13g2_decap_8 FILLER_78_224 ();
 sg13g2_fill_1 FILLER_78_231 ();
 sg13g2_fill_2 FILLER_78_237 ();
 sg13g2_decap_8 FILLER_78_243 ();
 sg13g2_fill_2 FILLER_78_250 ();
 sg13g2_fill_1 FILLER_78_252 ();
 sg13g2_fill_1 FILLER_78_266 ();
 sg13g2_decap_8 FILLER_78_293 ();
 sg13g2_fill_1 FILLER_78_300 ();
 sg13g2_fill_1 FILLER_78_350 ();
 sg13g2_decap_8 FILLER_78_381 ();
 sg13g2_decap_8 FILLER_78_388 ();
 sg13g2_decap_8 FILLER_78_395 ();
 sg13g2_decap_8 FILLER_78_402 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_decap_8 FILLER_79_231 ();
 sg13g2_decap_4 FILLER_79_238 ();
 sg13g2_fill_2 FILLER_79_242 ();
 sg13g2_decap_8 FILLER_79_248 ();
 sg13g2_decap_8 FILLER_79_255 ();
 sg13g2_decap_8 FILLER_79_262 ();
 sg13g2_decap_8 FILLER_79_269 ();
 sg13g2_decap_4 FILLER_79_276 ();
 sg13g2_decap_8 FILLER_79_387 ();
 sg13g2_decap_8 FILLER_79_394 ();
 sg13g2_decap_8 FILLER_79_401 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_4 FILLER_80_180 ();
 sg13g2_decap_4 FILLER_80_188 ();
 sg13g2_decap_4 FILLER_80_196 ();
 sg13g2_decap_4 FILLER_80_204 ();
 sg13g2_decap_4 FILLER_80_212 ();
 sg13g2_decap_4 FILLER_80_220 ();
 sg13g2_decap_4 FILLER_80_228 ();
 sg13g2_decap_8 FILLER_80_236 ();
 sg13g2_decap_8 FILLER_80_243 ();
 sg13g2_decap_8 FILLER_80_250 ();
 sg13g2_decap_8 FILLER_80_257 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_decap_8 FILLER_80_271 ();
 sg13g2_decap_4 FILLER_80_278 ();
 sg13g2_fill_1 FILLER_80_282 ();
 sg13g2_fill_2 FILLER_80_314 ();
 sg13g2_fill_1 FILLER_80_316 ();
 sg13g2_fill_2 FILLER_80_361 ();
 sg13g2_fill_1 FILLER_80_363 ();
 sg13g2_decap_8 FILLER_80_395 ();
 sg13g2_decap_8 FILLER_80_402 ();
 assign uio_oe[0] = net179;
 assign uio_oe[1] = net180;
 assign uio_oe[2] = net181;
 assign uio_oe[3] = net182;
 assign uio_oe[4] = net183;
 assign uio_oe[5] = net184;
 assign uio_oe[6] = net185;
 assign uio_oe[7] = net186;
 assign uio_out[0] = net187;
 assign uio_out[1] = net188;
 assign uio_out[2] = net189;
 assign uio_out[3] = net190;
 assign uio_out[4] = net191;
 assign uio_out[5] = net192;
 assign uio_out[6] = net193;
 assign uio_out[7] = net194;
 assign uo_out[1] = net195;
 assign uo_out[2] = net196;
 assign uo_out[3] = net197;
 assign uo_out[4] = net198;
 assign uo_out[5] = net199;
 assign uo_out[6] = net200;
 assign uo_out[7] = net201;
endmodule
